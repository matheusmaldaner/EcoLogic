library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs : in std_logic_vector(255 downto 0);
        outputs : out std_logic_vector(7679 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs : std_logic_vector(7679 downto 0);
    signal layer1_outputs : std_logic_vector(7679 downto 0);
    signal layer2_outputs : std_logic_vector(7679 downto 0);
    signal layer3_outputs : std_logic_vector(7679 downto 0);
    signal layer4_outputs : std_logic_vector(7679 downto 0);
    signal layer5_outputs : std_logic_vector(7679 downto 0);
    signal layer6_outputs : std_logic_vector(7679 downto 0);

begin

    layer0_outputs(0) <= not((inputs(223)) or (inputs(155)));
    layer0_outputs(1) <= not(inputs(67)) or (inputs(69));
    layer0_outputs(2) <= inputs(70);
    layer0_outputs(3) <= not(inputs(114));
    layer0_outputs(4) <= not(inputs(140));
    layer0_outputs(5) <= (inputs(172)) and not (inputs(17));
    layer0_outputs(6) <= (inputs(250)) or (inputs(235));
    layer0_outputs(7) <= not((inputs(238)) and (inputs(132)));
    layer0_outputs(8) <= not((inputs(85)) xor (inputs(160)));
    layer0_outputs(9) <= not((inputs(169)) or (inputs(47)));
    layer0_outputs(10) <= inputs(102);
    layer0_outputs(11) <= not((inputs(35)) and (inputs(116)));
    layer0_outputs(12) <= '0';
    layer0_outputs(13) <= not(inputs(16));
    layer0_outputs(14) <= (inputs(26)) or (inputs(49));
    layer0_outputs(15) <= (inputs(150)) or (inputs(146));
    layer0_outputs(16) <= not((inputs(31)) or (inputs(35)));
    layer0_outputs(17) <= not(inputs(62));
    layer0_outputs(18) <= not(inputs(152)) or (inputs(236));
    layer0_outputs(19) <= (inputs(85)) and not (inputs(205));
    layer0_outputs(20) <= not((inputs(198)) and (inputs(216)));
    layer0_outputs(21) <= '1';
    layer0_outputs(22) <= not((inputs(127)) or (inputs(6)));
    layer0_outputs(23) <= (inputs(223)) and not (inputs(22));
    layer0_outputs(24) <= not((inputs(51)) xor (inputs(4)));
    layer0_outputs(25) <= '1';
    layer0_outputs(26) <= '0';
    layer0_outputs(27) <= not(inputs(17)) or (inputs(1));
    layer0_outputs(28) <= not(inputs(37));
    layer0_outputs(29) <= inputs(118);
    layer0_outputs(30) <= inputs(31);
    layer0_outputs(31) <= not(inputs(7));
    layer0_outputs(32) <= (inputs(20)) and (inputs(119));
    layer0_outputs(33) <= not((inputs(57)) or (inputs(249)));
    layer0_outputs(34) <= '1';
    layer0_outputs(35) <= (inputs(209)) or (inputs(99));
    layer0_outputs(36) <= (inputs(66)) and (inputs(8));
    layer0_outputs(37) <= '0';
    layer0_outputs(38) <= not(inputs(169)) or (inputs(50));
    layer0_outputs(39) <= not(inputs(106));
    layer0_outputs(40) <= not(inputs(181)) or (inputs(62));
    layer0_outputs(41) <= not(inputs(66));
    layer0_outputs(42) <= not((inputs(74)) xor (inputs(121)));
    layer0_outputs(43) <= inputs(88);
    layer0_outputs(44) <= '1';
    layer0_outputs(45) <= not(inputs(89));
    layer0_outputs(46) <= not(inputs(110));
    layer0_outputs(47) <= not(inputs(8));
    layer0_outputs(48) <= inputs(182);
    layer0_outputs(49) <= not(inputs(149)) or (inputs(204));
    layer0_outputs(50) <= not(inputs(156));
    layer0_outputs(51) <= not((inputs(124)) xor (inputs(53)));
    layer0_outputs(52) <= inputs(114);
    layer0_outputs(53) <= (inputs(15)) and (inputs(210));
    layer0_outputs(54) <= not((inputs(144)) and (inputs(238)));
    layer0_outputs(55) <= inputs(105);
    layer0_outputs(56) <= inputs(199);
    layer0_outputs(57) <= inputs(119);
    layer0_outputs(58) <= not(inputs(159));
    layer0_outputs(59) <= not(inputs(223));
    layer0_outputs(60) <= (inputs(125)) or (inputs(231));
    layer0_outputs(61) <= not(inputs(252)) or (inputs(72));
    layer0_outputs(62) <= inputs(25);
    layer0_outputs(63) <= not(inputs(10));
    layer0_outputs(64) <= not(inputs(2));
    layer0_outputs(65) <= '1';
    layer0_outputs(66) <= inputs(20);
    layer0_outputs(67) <= not(inputs(235));
    layer0_outputs(68) <= not(inputs(212));
    layer0_outputs(69) <= inputs(142);
    layer0_outputs(70) <= '1';
    layer0_outputs(71) <= not(inputs(80));
    layer0_outputs(72) <= not(inputs(89));
    layer0_outputs(73) <= (inputs(140)) xor (inputs(188));
    layer0_outputs(74) <= not((inputs(17)) or (inputs(9)));
    layer0_outputs(75) <= '0';
    layer0_outputs(76) <= not((inputs(49)) or (inputs(117)));
    layer0_outputs(77) <= not(inputs(113));
    layer0_outputs(78) <= not(inputs(228));
    layer0_outputs(79) <= (inputs(164)) xor (inputs(181));
    layer0_outputs(80) <= '1';
    layer0_outputs(81) <= inputs(147);
    layer0_outputs(82) <= inputs(222);
    layer0_outputs(83) <= inputs(53);
    layer0_outputs(84) <= inputs(151);
    layer0_outputs(85) <= not(inputs(237)) or (inputs(158));
    layer0_outputs(86) <= not((inputs(26)) or (inputs(77)));
    layer0_outputs(87) <= (inputs(63)) and not (inputs(110));
    layer0_outputs(88) <= '0';
    layer0_outputs(89) <= '0';
    layer0_outputs(90) <= (inputs(219)) or (inputs(230));
    layer0_outputs(91) <= not((inputs(56)) or (inputs(243)));
    layer0_outputs(92) <= inputs(10);
    layer0_outputs(93) <= (inputs(83)) or (inputs(252));
    layer0_outputs(94) <= (inputs(104)) and not (inputs(205));
    layer0_outputs(95) <= not(inputs(110)) or (inputs(134));
    layer0_outputs(96) <= not((inputs(253)) or (inputs(122)));
    layer0_outputs(97) <= not(inputs(129)) or (inputs(180));
    layer0_outputs(98) <= inputs(32);
    layer0_outputs(99) <= inputs(12);
    layer0_outputs(100) <= inputs(172);
    layer0_outputs(101) <= not((inputs(2)) and (inputs(11)));
    layer0_outputs(102) <= (inputs(190)) or (inputs(160));
    layer0_outputs(103) <= not((inputs(84)) or (inputs(114)));
    layer0_outputs(104) <= not(inputs(181)) or (inputs(71));
    layer0_outputs(105) <= inputs(74);
    layer0_outputs(106) <= '1';
    layer0_outputs(107) <= '0';
    layer0_outputs(108) <= not(inputs(229)) or (inputs(229));
    layer0_outputs(109) <= not(inputs(23)) or (inputs(200));
    layer0_outputs(110) <= (inputs(196)) and not (inputs(119));
    layer0_outputs(111) <= (inputs(208)) xor (inputs(218));
    layer0_outputs(112) <= not((inputs(157)) and (inputs(58)));
    layer0_outputs(113) <= '1';
    layer0_outputs(114) <= inputs(119);
    layer0_outputs(115) <= not((inputs(93)) and (inputs(133)));
    layer0_outputs(116) <= not(inputs(22)) or (inputs(138));
    layer0_outputs(117) <= not(inputs(105));
    layer0_outputs(118) <= (inputs(205)) or (inputs(233));
    layer0_outputs(119) <= not(inputs(24)) or (inputs(109));
    layer0_outputs(120) <= not(inputs(188)) or (inputs(181));
    layer0_outputs(121) <= inputs(14);
    layer0_outputs(122) <= inputs(140);
    layer0_outputs(123) <= (inputs(173)) and not (inputs(205));
    layer0_outputs(124) <= inputs(242);
    layer0_outputs(125) <= '0';
    layer0_outputs(126) <= '0';
    layer0_outputs(127) <= not(inputs(145));
    layer0_outputs(128) <= not((inputs(83)) and (inputs(104)));
    layer0_outputs(129) <= (inputs(9)) and (inputs(51));
    layer0_outputs(130) <= not(inputs(115));
    layer0_outputs(131) <= inputs(71);
    layer0_outputs(132) <= not(inputs(138));
    layer0_outputs(133) <= inputs(194);
    layer0_outputs(134) <= not((inputs(92)) and (inputs(166)));
    layer0_outputs(135) <= inputs(245);
    layer0_outputs(136) <= (inputs(39)) and not (inputs(147));
    layer0_outputs(137) <= (inputs(86)) and not (inputs(4));
    layer0_outputs(138) <= not(inputs(191));
    layer0_outputs(139) <= not((inputs(147)) or (inputs(195)));
    layer0_outputs(140) <= inputs(72);
    layer0_outputs(141) <= not(inputs(87)) or (inputs(66));
    layer0_outputs(142) <= (inputs(132)) and not (inputs(34));
    layer0_outputs(143) <= not((inputs(69)) or (inputs(117)));
    layer0_outputs(144) <= inputs(99);
    layer0_outputs(145) <= (inputs(251)) or (inputs(234));
    layer0_outputs(146) <= not(inputs(68));
    layer0_outputs(147) <= not((inputs(88)) xor (inputs(29)));
    layer0_outputs(148) <= not((inputs(52)) and (inputs(15)));
    layer0_outputs(149) <= not(inputs(53));
    layer0_outputs(150) <= '1';
    layer0_outputs(151) <= (inputs(121)) and not (inputs(100));
    layer0_outputs(152) <= not(inputs(194));
    layer0_outputs(153) <= (inputs(92)) or (inputs(122));
    layer0_outputs(154) <= not(inputs(59));
    layer0_outputs(155) <= (inputs(130)) and not (inputs(102));
    layer0_outputs(156) <= (inputs(241)) and not (inputs(174));
    layer0_outputs(157) <= (inputs(119)) and (inputs(92));
    layer0_outputs(158) <= (inputs(71)) and not (inputs(150));
    layer0_outputs(159) <= '1';
    layer0_outputs(160) <= not(inputs(239));
    layer0_outputs(161) <= inputs(247);
    layer0_outputs(162) <= (inputs(28)) xor (inputs(241));
    layer0_outputs(163) <= inputs(177);
    layer0_outputs(164) <= not(inputs(197));
    layer0_outputs(165) <= (inputs(193)) or (inputs(71));
    layer0_outputs(166) <= '1';
    layer0_outputs(167) <= not(inputs(166));
    layer0_outputs(168) <= (inputs(16)) or (inputs(70));
    layer0_outputs(169) <= (inputs(216)) or (inputs(197));
    layer0_outputs(170) <= not(inputs(28)) or (inputs(5));
    layer0_outputs(171) <= not(inputs(43));
    layer0_outputs(172) <= inputs(234);
    layer0_outputs(173) <= not(inputs(217));
    layer0_outputs(174) <= (inputs(83)) or (inputs(238));
    layer0_outputs(175) <= '1';
    layer0_outputs(176) <= not((inputs(175)) and (inputs(82)));
    layer0_outputs(177) <= not(inputs(224));
    layer0_outputs(178) <= '1';
    layer0_outputs(179) <= not(inputs(127)) or (inputs(119));
    layer0_outputs(180) <= '0';
    layer0_outputs(181) <= '1';
    layer0_outputs(182) <= (inputs(203)) and not (inputs(152));
    layer0_outputs(183) <= '1';
    layer0_outputs(184) <= not(inputs(129));
    layer0_outputs(185) <= (inputs(101)) and not (inputs(222));
    layer0_outputs(186) <= not(inputs(6));
    layer0_outputs(187) <= inputs(212);
    layer0_outputs(188) <= '0';
    layer0_outputs(189) <= inputs(44);
    layer0_outputs(190) <= inputs(28);
    layer0_outputs(191) <= (inputs(184)) or (inputs(1));
    layer0_outputs(192) <= (inputs(168)) or (inputs(56));
    layer0_outputs(193) <= inputs(29);
    layer0_outputs(194) <= not(inputs(134));
    layer0_outputs(195) <= inputs(118);
    layer0_outputs(196) <= (inputs(5)) or (inputs(220));
    layer0_outputs(197) <= inputs(230);
    layer0_outputs(198) <= (inputs(8)) xor (inputs(191));
    layer0_outputs(199) <= (inputs(147)) and not (inputs(228));
    layer0_outputs(200) <= not(inputs(193));
    layer0_outputs(201) <= inputs(16);
    layer0_outputs(202) <= not(inputs(211));
    layer0_outputs(203) <= not(inputs(36));
    layer0_outputs(204) <= (inputs(214)) and not (inputs(137));
    layer0_outputs(205) <= not(inputs(122));
    layer0_outputs(206) <= not(inputs(80)) or (inputs(231));
    layer0_outputs(207) <= '1';
    layer0_outputs(208) <= (inputs(204)) and not (inputs(135));
    layer0_outputs(209) <= (inputs(253)) or (inputs(157));
    layer0_outputs(210) <= not((inputs(158)) or (inputs(248)));
    layer0_outputs(211) <= not((inputs(223)) or (inputs(188)));
    layer0_outputs(212) <= not((inputs(213)) and (inputs(138)));
    layer0_outputs(213) <= not(inputs(138)) or (inputs(46));
    layer0_outputs(214) <= inputs(116);
    layer0_outputs(215) <= not(inputs(234)) or (inputs(112));
    layer0_outputs(216) <= (inputs(67)) and not (inputs(13));
    layer0_outputs(217) <= inputs(86);
    layer0_outputs(218) <= (inputs(253)) and (inputs(203));
    layer0_outputs(219) <= not((inputs(161)) or (inputs(102)));
    layer0_outputs(220) <= not(inputs(33));
    layer0_outputs(221) <= '1';
    layer0_outputs(222) <= not(inputs(255));
    layer0_outputs(223) <= inputs(201);
    layer0_outputs(224) <= (inputs(200)) and not (inputs(184));
    layer0_outputs(225) <= (inputs(22)) or (inputs(108));
    layer0_outputs(226) <= not(inputs(154)) or (inputs(215));
    layer0_outputs(227) <= not(inputs(190));
    layer0_outputs(228) <= inputs(21);
    layer0_outputs(229) <= (inputs(124)) and not (inputs(151));
    layer0_outputs(230) <= not(inputs(197)) or (inputs(28));
    layer0_outputs(231) <= not(inputs(115));
    layer0_outputs(232) <= inputs(161);
    layer0_outputs(233) <= not((inputs(130)) or (inputs(85)));
    layer0_outputs(234) <= (inputs(159)) and not (inputs(233));
    layer0_outputs(235) <= (inputs(192)) and not (inputs(0));
    layer0_outputs(236) <= not(inputs(65));
    layer0_outputs(237) <= inputs(76);
    layer0_outputs(238) <= (inputs(13)) and (inputs(0));
    layer0_outputs(239) <= (inputs(193)) or (inputs(229));
    layer0_outputs(240) <= not((inputs(13)) or (inputs(113)));
    layer0_outputs(241) <= '1';
    layer0_outputs(242) <= '1';
    layer0_outputs(243) <= (inputs(172)) and (inputs(122));
    layer0_outputs(244) <= not((inputs(7)) or (inputs(121)));
    layer0_outputs(245) <= not(inputs(57));
    layer0_outputs(246) <= '0';
    layer0_outputs(247) <= '0';
    layer0_outputs(248) <= not(inputs(43));
    layer0_outputs(249) <= '1';
    layer0_outputs(250) <= inputs(114);
    layer0_outputs(251) <= (inputs(17)) and not (inputs(24));
    layer0_outputs(252) <= not(inputs(153)) or (inputs(210));
    layer0_outputs(253) <= not(inputs(170)) or (inputs(163));
    layer0_outputs(254) <= '0';
    layer0_outputs(255) <= (inputs(232)) and (inputs(88));
    layer0_outputs(256) <= not(inputs(231)) or (inputs(125));
    layer0_outputs(257) <= (inputs(207)) or (inputs(174));
    layer0_outputs(258) <= (inputs(232)) or (inputs(251));
    layer0_outputs(259) <= not(inputs(72)) or (inputs(213));
    layer0_outputs(260) <= (inputs(140)) or (inputs(143));
    layer0_outputs(261) <= not(inputs(188)) or (inputs(242));
    layer0_outputs(262) <= (inputs(164)) or (inputs(236));
    layer0_outputs(263) <= (inputs(82)) and (inputs(14));
    layer0_outputs(264) <= not((inputs(202)) or (inputs(103)));
    layer0_outputs(265) <= not((inputs(162)) and (inputs(172)));
    layer0_outputs(266) <= '1';
    layer0_outputs(267) <= not(inputs(102));
    layer0_outputs(268) <= '1';
    layer0_outputs(269) <= not((inputs(81)) and (inputs(213)));
    layer0_outputs(270) <= (inputs(158)) and not (inputs(69));
    layer0_outputs(271) <= '0';
    layer0_outputs(272) <= (inputs(147)) or (inputs(110));
    layer0_outputs(273) <= not(inputs(114));
    layer0_outputs(274) <= not((inputs(240)) and (inputs(167)));
    layer0_outputs(275) <= (inputs(52)) or (inputs(8));
    layer0_outputs(276) <= not(inputs(15));
    layer0_outputs(277) <= (inputs(191)) xor (inputs(165));
    layer0_outputs(278) <= inputs(148);
    layer0_outputs(279) <= (inputs(30)) or (inputs(102));
    layer0_outputs(280) <= not(inputs(160));
    layer0_outputs(281) <= (inputs(52)) and not (inputs(159));
    layer0_outputs(282) <= (inputs(12)) and not (inputs(101));
    layer0_outputs(283) <= not((inputs(197)) or (inputs(48)));
    layer0_outputs(284) <= inputs(185);
    layer0_outputs(285) <= inputs(201);
    layer0_outputs(286) <= '1';
    layer0_outputs(287) <= not(inputs(128)) or (inputs(88));
    layer0_outputs(288) <= (inputs(107)) or (inputs(250));
    layer0_outputs(289) <= (inputs(189)) and not (inputs(8));
    layer0_outputs(290) <= (inputs(64)) and (inputs(201));
    layer0_outputs(291) <= not(inputs(219));
    layer0_outputs(292) <= (inputs(53)) and not (inputs(45));
    layer0_outputs(293) <= not(inputs(63)) or (inputs(148));
    layer0_outputs(294) <= not(inputs(95)) or (inputs(72));
    layer0_outputs(295) <= (inputs(6)) or (inputs(189));
    layer0_outputs(296) <= not(inputs(177));
    layer0_outputs(297) <= (inputs(35)) and not (inputs(7));
    layer0_outputs(298) <= (inputs(64)) or (inputs(239));
    layer0_outputs(299) <= inputs(130);
    layer0_outputs(300) <= '1';
    layer0_outputs(301) <= (inputs(21)) or (inputs(169));
    layer0_outputs(302) <= (inputs(4)) and not (inputs(79));
    layer0_outputs(303) <= inputs(229);
    layer0_outputs(304) <= '1';
    layer0_outputs(305) <= not(inputs(112)) or (inputs(18));
    layer0_outputs(306) <= not(inputs(135)) or (inputs(29));
    layer0_outputs(307) <= not(inputs(112)) or (inputs(97));
    layer0_outputs(308) <= (inputs(246)) or (inputs(195));
    layer0_outputs(309) <= not(inputs(22));
    layer0_outputs(310) <= not(inputs(44));
    layer0_outputs(311) <= (inputs(122)) or (inputs(19));
    layer0_outputs(312) <= '1';
    layer0_outputs(313) <= inputs(132);
    layer0_outputs(314) <= not(inputs(187)) or (inputs(87));
    layer0_outputs(315) <= (inputs(126)) and not (inputs(214));
    layer0_outputs(316) <= (inputs(67)) or (inputs(109));
    layer0_outputs(317) <= not(inputs(40)) or (inputs(230));
    layer0_outputs(318) <= (inputs(37)) and (inputs(48));
    layer0_outputs(319) <= not(inputs(124));
    layer0_outputs(320) <= inputs(15);
    layer0_outputs(321) <= not((inputs(96)) and (inputs(72)));
    layer0_outputs(322) <= '0';
    layer0_outputs(323) <= inputs(122);
    layer0_outputs(324) <= inputs(195);
    layer0_outputs(325) <= not((inputs(219)) and (inputs(86)));
    layer0_outputs(326) <= inputs(120);
    layer0_outputs(327) <= not(inputs(62)) or (inputs(35));
    layer0_outputs(328) <= '1';
    layer0_outputs(329) <= inputs(27);
    layer0_outputs(330) <= (inputs(192)) and not (inputs(193));
    layer0_outputs(331) <= '1';
    layer0_outputs(332) <= not(inputs(33));
    layer0_outputs(333) <= (inputs(0)) or (inputs(223));
    layer0_outputs(334) <= inputs(190);
    layer0_outputs(335) <= not((inputs(41)) and (inputs(192)));
    layer0_outputs(336) <= not(inputs(227));
    layer0_outputs(337) <= not(inputs(178)) or (inputs(31));
    layer0_outputs(338) <= not(inputs(48));
    layer0_outputs(339) <= (inputs(203)) xor (inputs(236));
    layer0_outputs(340) <= '0';
    layer0_outputs(341) <= not(inputs(15));
    layer0_outputs(342) <= not(inputs(185));
    layer0_outputs(343) <= (inputs(156)) and not (inputs(80));
    layer0_outputs(344) <= (inputs(132)) and (inputs(151));
    layer0_outputs(345) <= not((inputs(234)) xor (inputs(33)));
    layer0_outputs(346) <= inputs(21);
    layer0_outputs(347) <= not(inputs(203));
    layer0_outputs(348) <= not((inputs(116)) xor (inputs(127)));
    layer0_outputs(349) <= not(inputs(98));
    layer0_outputs(350) <= (inputs(154)) and not (inputs(15));
    layer0_outputs(351) <= '0';
    layer0_outputs(352) <= not((inputs(237)) or (inputs(221)));
    layer0_outputs(353) <= (inputs(127)) and (inputs(198));
    layer0_outputs(354) <= (inputs(53)) and not (inputs(102));
    layer0_outputs(355) <= not(inputs(164)) or (inputs(202));
    layer0_outputs(356) <= (inputs(98)) and not (inputs(155));
    layer0_outputs(357) <= inputs(1);
    layer0_outputs(358) <= (inputs(156)) or (inputs(29));
    layer0_outputs(359) <= '1';
    layer0_outputs(360) <= inputs(160);
    layer0_outputs(361) <= '0';
    layer0_outputs(362) <= not(inputs(203)) or (inputs(211));
    layer0_outputs(363) <= inputs(181);
    layer0_outputs(364) <= '0';
    layer0_outputs(365) <= not(inputs(198)) or (inputs(98));
    layer0_outputs(366) <= '1';
    layer0_outputs(367) <= not((inputs(43)) or (inputs(8)));
    layer0_outputs(368) <= (inputs(105)) and not (inputs(86));
    layer0_outputs(369) <= (inputs(202)) and not (inputs(108));
    layer0_outputs(370) <= (inputs(154)) and (inputs(77));
    layer0_outputs(371) <= '0';
    layer0_outputs(372) <= (inputs(112)) and (inputs(146));
    layer0_outputs(373) <= inputs(73);
    layer0_outputs(374) <= not(inputs(205)) or (inputs(185));
    layer0_outputs(375) <= (inputs(206)) and (inputs(63));
    layer0_outputs(376) <= (inputs(40)) and not (inputs(173));
    layer0_outputs(377) <= (inputs(119)) or (inputs(14));
    layer0_outputs(378) <= inputs(77);
    layer0_outputs(379) <= not((inputs(254)) and (inputs(149)));
    layer0_outputs(380) <= not(inputs(70));
    layer0_outputs(381) <= not(inputs(194));
    layer0_outputs(382) <= (inputs(20)) and not (inputs(234));
    layer0_outputs(383) <= not(inputs(224)) or (inputs(169));
    layer0_outputs(384) <= not(inputs(166));
    layer0_outputs(385) <= not(inputs(149)) or (inputs(142));
    layer0_outputs(386) <= not(inputs(203)) or (inputs(203));
    layer0_outputs(387) <= not(inputs(131));
    layer0_outputs(388) <= not(inputs(202)) or (inputs(235));
    layer0_outputs(389) <= not((inputs(155)) and (inputs(236)));
    layer0_outputs(390) <= not((inputs(18)) and (inputs(68)));
    layer0_outputs(391) <= inputs(136);
    layer0_outputs(392) <= inputs(92);
    layer0_outputs(393) <= (inputs(143)) or (inputs(37));
    layer0_outputs(394) <= not(inputs(11)) or (inputs(143));
    layer0_outputs(395) <= (inputs(110)) and not (inputs(23));
    layer0_outputs(396) <= not((inputs(70)) xor (inputs(90)));
    layer0_outputs(397) <= not((inputs(186)) or (inputs(211)));
    layer0_outputs(398) <= not((inputs(164)) or (inputs(77)));
    layer0_outputs(399) <= not((inputs(126)) or (inputs(93)));
    layer0_outputs(400) <= not(inputs(210));
    layer0_outputs(401) <= (inputs(160)) and (inputs(68));
    layer0_outputs(402) <= not(inputs(77));
    layer0_outputs(403) <= '1';
    layer0_outputs(404) <= (inputs(120)) or (inputs(151));
    layer0_outputs(405) <= '0';
    layer0_outputs(406) <= inputs(93);
    layer0_outputs(407) <= '1';
    layer0_outputs(408) <= not((inputs(186)) or (inputs(219)));
    layer0_outputs(409) <= (inputs(229)) or (inputs(173));
    layer0_outputs(410) <= not((inputs(186)) and (inputs(22)));
    layer0_outputs(411) <= (inputs(47)) and (inputs(142));
    layer0_outputs(412) <= (inputs(94)) or (inputs(216));
    layer0_outputs(413) <= not((inputs(131)) or (inputs(53)));
    layer0_outputs(414) <= '1';
    layer0_outputs(415) <= (inputs(11)) and not (inputs(207));
    layer0_outputs(416) <= not(inputs(161));
    layer0_outputs(417) <= (inputs(1)) or (inputs(225));
    layer0_outputs(418) <= not(inputs(2));
    layer0_outputs(419) <= not((inputs(199)) or (inputs(231)));
    layer0_outputs(420) <= not((inputs(176)) xor (inputs(96)));
    layer0_outputs(421) <= inputs(79);
    layer0_outputs(422) <= (inputs(202)) and (inputs(244));
    layer0_outputs(423) <= inputs(72);
    layer0_outputs(424) <= not((inputs(172)) xor (inputs(21)));
    layer0_outputs(425) <= not((inputs(52)) or (inputs(137)));
    layer0_outputs(426) <= not(inputs(1)) or (inputs(138));
    layer0_outputs(427) <= '0';
    layer0_outputs(428) <= not(inputs(126)) or (inputs(213));
    layer0_outputs(429) <= (inputs(234)) xor (inputs(11));
    layer0_outputs(430) <= inputs(232);
    layer0_outputs(431) <= (inputs(127)) and (inputs(183));
    layer0_outputs(432) <= inputs(164);
    layer0_outputs(433) <= (inputs(51)) xor (inputs(48));
    layer0_outputs(434) <= not((inputs(96)) or (inputs(128)));
    layer0_outputs(435) <= not(inputs(216)) or (inputs(183));
    layer0_outputs(436) <= not((inputs(51)) xor (inputs(65)));
    layer0_outputs(437) <= '0';
    layer0_outputs(438) <= '0';
    layer0_outputs(439) <= (inputs(196)) and not (inputs(230));
    layer0_outputs(440) <= not(inputs(231)) or (inputs(20));
    layer0_outputs(441) <= (inputs(114)) and not (inputs(245));
    layer0_outputs(442) <= not((inputs(170)) and (inputs(66)));
    layer0_outputs(443) <= not(inputs(34));
    layer0_outputs(444) <= not(inputs(156)) or (inputs(37));
    layer0_outputs(445) <= inputs(212);
    layer0_outputs(446) <= (inputs(165)) and not (inputs(142));
    layer0_outputs(447) <= inputs(59);
    layer0_outputs(448) <= (inputs(47)) and (inputs(48));
    layer0_outputs(449) <= '1';
    layer0_outputs(450) <= not((inputs(14)) or (inputs(242)));
    layer0_outputs(451) <= (inputs(248)) or (inputs(20));
    layer0_outputs(452) <= not((inputs(160)) or (inputs(67)));
    layer0_outputs(453) <= (inputs(185)) or (inputs(206));
    layer0_outputs(454) <= inputs(131);
    layer0_outputs(455) <= '1';
    layer0_outputs(456) <= (inputs(81)) or (inputs(115));
    layer0_outputs(457) <= (inputs(87)) and not (inputs(14));
    layer0_outputs(458) <= not(inputs(196)) or (inputs(45));
    layer0_outputs(459) <= not((inputs(129)) or (inputs(130)));
    layer0_outputs(460) <= not(inputs(229)) or (inputs(98));
    layer0_outputs(461) <= '1';
    layer0_outputs(462) <= '0';
    layer0_outputs(463) <= not(inputs(233)) or (inputs(74));
    layer0_outputs(464) <= inputs(54);
    layer0_outputs(465) <= not(inputs(11)) or (inputs(63));
    layer0_outputs(466) <= '1';
    layer0_outputs(467) <= '1';
    layer0_outputs(468) <= (inputs(137)) or (inputs(223));
    layer0_outputs(469) <= (inputs(239)) and not (inputs(150));
    layer0_outputs(470) <= (inputs(146)) and not (inputs(236));
    layer0_outputs(471) <= (inputs(8)) and not (inputs(199));
    layer0_outputs(472) <= (inputs(31)) or (inputs(35));
    layer0_outputs(473) <= not((inputs(34)) or (inputs(150)));
    layer0_outputs(474) <= not(inputs(17)) or (inputs(241));
    layer0_outputs(475) <= inputs(85);
    layer0_outputs(476) <= not((inputs(74)) xor (inputs(79)));
    layer0_outputs(477) <= inputs(182);
    layer0_outputs(478) <= '1';
    layer0_outputs(479) <= (inputs(86)) or (inputs(222));
    layer0_outputs(480) <= (inputs(111)) and not (inputs(126));
    layer0_outputs(481) <= not(inputs(118));
    layer0_outputs(482) <= (inputs(79)) and not (inputs(89));
    layer0_outputs(483) <= (inputs(38)) and (inputs(226));
    layer0_outputs(484) <= inputs(161);
    layer0_outputs(485) <= (inputs(29)) and not (inputs(91));
    layer0_outputs(486) <= '1';
    layer0_outputs(487) <= not((inputs(243)) or (inputs(7)));
    layer0_outputs(488) <= '1';
    layer0_outputs(489) <= not(inputs(63));
    layer0_outputs(490) <= (inputs(50)) and (inputs(86));
    layer0_outputs(491) <= (inputs(236)) or (inputs(206));
    layer0_outputs(492) <= inputs(110);
    layer0_outputs(493) <= not((inputs(108)) xor (inputs(70)));
    layer0_outputs(494) <= inputs(1);
    layer0_outputs(495) <= not(inputs(240));
    layer0_outputs(496) <= not(inputs(14));
    layer0_outputs(497) <= '1';
    layer0_outputs(498) <= not((inputs(147)) or (inputs(196)));
    layer0_outputs(499) <= '0';
    layer0_outputs(500) <= inputs(246);
    layer0_outputs(501) <= (inputs(114)) and not (inputs(116));
    layer0_outputs(502) <= inputs(38);
    layer0_outputs(503) <= not(inputs(181));
    layer0_outputs(504) <= (inputs(20)) xor (inputs(119));
    layer0_outputs(505) <= not(inputs(120));
    layer0_outputs(506) <= (inputs(104)) xor (inputs(138));
    layer0_outputs(507) <= not((inputs(36)) or (inputs(45)));
    layer0_outputs(508) <= not(inputs(168));
    layer0_outputs(509) <= inputs(205);
    layer0_outputs(510) <= not((inputs(139)) xor (inputs(131)));
    layer0_outputs(511) <= inputs(142);
    layer0_outputs(512) <= not(inputs(195)) or (inputs(75));
    layer0_outputs(513) <= not(inputs(159)) or (inputs(163));
    layer0_outputs(514) <= not(inputs(58));
    layer0_outputs(515) <= inputs(168);
    layer0_outputs(516) <= inputs(73);
    layer0_outputs(517) <= not(inputs(162));
    layer0_outputs(518) <= not(inputs(19)) or (inputs(158));
    layer0_outputs(519) <= (inputs(65)) or (inputs(192));
    layer0_outputs(520) <= '0';
    layer0_outputs(521) <= not(inputs(229));
    layer0_outputs(522) <= '1';
    layer0_outputs(523) <= not(inputs(133));
    layer0_outputs(524) <= not(inputs(148));
    layer0_outputs(525) <= not((inputs(133)) or (inputs(70)));
    layer0_outputs(526) <= (inputs(115)) and (inputs(64));
    layer0_outputs(527) <= (inputs(153)) and (inputs(13));
    layer0_outputs(528) <= not((inputs(119)) xor (inputs(75)));
    layer0_outputs(529) <= inputs(19);
    layer0_outputs(530) <= not(inputs(216));
    layer0_outputs(531) <= not((inputs(58)) and (inputs(23)));
    layer0_outputs(532) <= not(inputs(203));
    layer0_outputs(533) <= not(inputs(228)) or (inputs(167));
    layer0_outputs(534) <= not(inputs(35));
    layer0_outputs(535) <= inputs(4);
    layer0_outputs(536) <= (inputs(188)) and (inputs(224));
    layer0_outputs(537) <= inputs(229);
    layer0_outputs(538) <= not((inputs(147)) or (inputs(18)));
    layer0_outputs(539) <= inputs(157);
    layer0_outputs(540) <= (inputs(142)) and (inputs(153));
    layer0_outputs(541) <= not((inputs(24)) and (inputs(89)));
    layer0_outputs(542) <= inputs(9);
    layer0_outputs(543) <= not(inputs(68)) or (inputs(191));
    layer0_outputs(544) <= (inputs(105)) and not (inputs(233));
    layer0_outputs(545) <= (inputs(197)) and (inputs(32));
    layer0_outputs(546) <= '1';
    layer0_outputs(547) <= inputs(56);
    layer0_outputs(548) <= inputs(221);
    layer0_outputs(549) <= not((inputs(173)) and (inputs(214)));
    layer0_outputs(550) <= '0';
    layer0_outputs(551) <= not(inputs(163)) or (inputs(24));
    layer0_outputs(552) <= not((inputs(96)) and (inputs(23)));
    layer0_outputs(553) <= not((inputs(67)) and (inputs(129)));
    layer0_outputs(554) <= (inputs(248)) and not (inputs(253));
    layer0_outputs(555) <= not((inputs(246)) xor (inputs(231)));
    layer0_outputs(556) <= '1';
    layer0_outputs(557) <= (inputs(168)) or (inputs(32));
    layer0_outputs(558) <= not((inputs(25)) and (inputs(58)));
    layer0_outputs(559) <= not((inputs(7)) and (inputs(81)));
    layer0_outputs(560) <= not((inputs(24)) xor (inputs(70)));
    layer0_outputs(561) <= '1';
    layer0_outputs(562) <= not((inputs(150)) and (inputs(161)));
    layer0_outputs(563) <= '1';
    layer0_outputs(564) <= not(inputs(69)) or (inputs(148));
    layer0_outputs(565) <= '1';
    layer0_outputs(566) <= inputs(233);
    layer0_outputs(567) <= '1';
    layer0_outputs(568) <= '1';
    layer0_outputs(569) <= inputs(72);
    layer0_outputs(570) <= '1';
    layer0_outputs(571) <= (inputs(144)) and not (inputs(121));
    layer0_outputs(572) <= not(inputs(177));
    layer0_outputs(573) <= '0';
    layer0_outputs(574) <= (inputs(218)) or (inputs(224));
    layer0_outputs(575) <= (inputs(134)) or (inputs(86));
    layer0_outputs(576) <= not(inputs(209));
    layer0_outputs(577) <= inputs(179);
    layer0_outputs(578) <= not(inputs(145)) or (inputs(94));
    layer0_outputs(579) <= inputs(68);
    layer0_outputs(580) <= inputs(127);
    layer0_outputs(581) <= inputs(145);
    layer0_outputs(582) <= (inputs(69)) and (inputs(150));
    layer0_outputs(583) <= '1';
    layer0_outputs(584) <= not(inputs(233)) or (inputs(113));
    layer0_outputs(585) <= inputs(52);
    layer0_outputs(586) <= '0';
    layer0_outputs(587) <= (inputs(156)) and not (inputs(193));
    layer0_outputs(588) <= (inputs(201)) or (inputs(34));
    layer0_outputs(589) <= (inputs(18)) and not (inputs(65));
    layer0_outputs(590) <= inputs(8);
    layer0_outputs(591) <= not(inputs(55)) or (inputs(176));
    layer0_outputs(592) <= inputs(188);
    layer0_outputs(593) <= '1';
    layer0_outputs(594) <= (inputs(239)) and not (inputs(10));
    layer0_outputs(595) <= (inputs(19)) or (inputs(171));
    layer0_outputs(596) <= inputs(50);
    layer0_outputs(597) <= (inputs(6)) and not (inputs(97));
    layer0_outputs(598) <= (inputs(31)) or (inputs(237));
    layer0_outputs(599) <= not(inputs(211)) or (inputs(14));
    layer0_outputs(600) <= not(inputs(192)) or (inputs(114));
    layer0_outputs(601) <= not(inputs(213));
    layer0_outputs(602) <= not(inputs(73));
    layer0_outputs(603) <= inputs(103);
    layer0_outputs(604) <= (inputs(132)) and not (inputs(65));
    layer0_outputs(605) <= (inputs(201)) and not (inputs(69));
    layer0_outputs(606) <= not(inputs(181));
    layer0_outputs(607) <= not((inputs(31)) and (inputs(134)));
    layer0_outputs(608) <= not(inputs(191)) or (inputs(22));
    layer0_outputs(609) <= not((inputs(27)) and (inputs(25)));
    layer0_outputs(610) <= not((inputs(228)) or (inputs(227)));
    layer0_outputs(611) <= inputs(111);
    layer0_outputs(612) <= inputs(206);
    layer0_outputs(613) <= (inputs(205)) or (inputs(252));
    layer0_outputs(614) <= not(inputs(201)) or (inputs(70));
    layer0_outputs(615) <= '0';
    layer0_outputs(616) <= not(inputs(249)) or (inputs(188));
    layer0_outputs(617) <= (inputs(218)) or (inputs(178));
    layer0_outputs(618) <= inputs(25);
    layer0_outputs(619) <= (inputs(228)) or (inputs(43));
    layer0_outputs(620) <= inputs(169);
    layer0_outputs(621) <= '0';
    layer0_outputs(622) <= not(inputs(99));
    layer0_outputs(623) <= not((inputs(10)) and (inputs(236)));
    layer0_outputs(624) <= (inputs(130)) or (inputs(14));
    layer0_outputs(625) <= (inputs(183)) and not (inputs(190));
    layer0_outputs(626) <= (inputs(1)) and not (inputs(157));
    layer0_outputs(627) <= not((inputs(107)) xor (inputs(16)));
    layer0_outputs(628) <= inputs(92);
    layer0_outputs(629) <= (inputs(222)) and (inputs(64));
    layer0_outputs(630) <= inputs(146);
    layer0_outputs(631) <= '1';
    layer0_outputs(632) <= not(inputs(26)) or (inputs(191));
    layer0_outputs(633) <= (inputs(132)) and not (inputs(194));
    layer0_outputs(634) <= (inputs(190)) and not (inputs(185));
    layer0_outputs(635) <= not((inputs(151)) xor (inputs(111)));
    layer0_outputs(636) <= '0';
    layer0_outputs(637) <= (inputs(134)) or (inputs(109));
    layer0_outputs(638) <= not(inputs(231)) or (inputs(209));
    layer0_outputs(639) <= inputs(213);
    layer0_outputs(640) <= (inputs(29)) and (inputs(190));
    layer0_outputs(641) <= not((inputs(19)) or (inputs(228)));
    layer0_outputs(642) <= (inputs(244)) and not (inputs(120));
    layer0_outputs(643) <= '0';
    layer0_outputs(644) <= not(inputs(54));
    layer0_outputs(645) <= not((inputs(180)) or (inputs(139)));
    layer0_outputs(646) <= (inputs(113)) and not (inputs(118));
    layer0_outputs(647) <= not((inputs(23)) or (inputs(191)));
    layer0_outputs(648) <= not(inputs(78));
    layer0_outputs(649) <= '1';
    layer0_outputs(650) <= not(inputs(98)) or (inputs(145));
    layer0_outputs(651) <= (inputs(3)) or (inputs(188));
    layer0_outputs(652) <= (inputs(21)) and (inputs(179));
    layer0_outputs(653) <= inputs(29);
    layer0_outputs(654) <= not((inputs(9)) xor (inputs(49)));
    layer0_outputs(655) <= inputs(111);
    layer0_outputs(656) <= inputs(29);
    layer0_outputs(657) <= (inputs(144)) and not (inputs(114));
    layer0_outputs(658) <= inputs(254);
    layer0_outputs(659) <= not(inputs(191));
    layer0_outputs(660) <= inputs(182);
    layer0_outputs(661) <= '0';
    layer0_outputs(662) <= not((inputs(220)) and (inputs(142)));
    layer0_outputs(663) <= inputs(195);
    layer0_outputs(664) <= (inputs(33)) and not (inputs(128));
    layer0_outputs(665) <= inputs(132);
    layer0_outputs(666) <= not((inputs(183)) or (inputs(112)));
    layer0_outputs(667) <= not(inputs(5));
    layer0_outputs(668) <= not((inputs(226)) or (inputs(208)));
    layer0_outputs(669) <= inputs(188);
    layer0_outputs(670) <= inputs(25);
    layer0_outputs(671) <= (inputs(0)) and not (inputs(159));
    layer0_outputs(672) <= not((inputs(15)) xor (inputs(254)));
    layer0_outputs(673) <= not(inputs(158));
    layer0_outputs(674) <= not(inputs(217));
    layer0_outputs(675) <= inputs(249);
    layer0_outputs(676) <= not(inputs(24)) or (inputs(152));
    layer0_outputs(677) <= not(inputs(196)) or (inputs(14));
    layer0_outputs(678) <= not((inputs(73)) and (inputs(45)));
    layer0_outputs(679) <= '1';
    layer0_outputs(680) <= inputs(103);
    layer0_outputs(681) <= (inputs(76)) and not (inputs(1));
    layer0_outputs(682) <= not(inputs(16));
    layer0_outputs(683) <= '1';
    layer0_outputs(684) <= (inputs(134)) or (inputs(15));
    layer0_outputs(685) <= inputs(202);
    layer0_outputs(686) <= not((inputs(187)) xor (inputs(218)));
    layer0_outputs(687) <= not(inputs(97));
    layer0_outputs(688) <= inputs(252);
    layer0_outputs(689) <= inputs(6);
    layer0_outputs(690) <= not((inputs(93)) or (inputs(172)));
    layer0_outputs(691) <= '1';
    layer0_outputs(692) <= '0';
    layer0_outputs(693) <= inputs(211);
    layer0_outputs(694) <= not(inputs(136)) or (inputs(161));
    layer0_outputs(695) <= '0';
    layer0_outputs(696) <= not((inputs(248)) and (inputs(204)));
    layer0_outputs(697) <= inputs(19);
    layer0_outputs(698) <= inputs(79);
    layer0_outputs(699) <= (inputs(23)) and not (inputs(31));
    layer0_outputs(700) <= inputs(238);
    layer0_outputs(701) <= '0';
    layer0_outputs(702) <= inputs(117);
    layer0_outputs(703) <= not(inputs(182)) or (inputs(157));
    layer0_outputs(704) <= not(inputs(83));
    layer0_outputs(705) <= inputs(119);
    layer0_outputs(706) <= (inputs(184)) and (inputs(4));
    layer0_outputs(707) <= (inputs(111)) and (inputs(212));
    layer0_outputs(708) <= not(inputs(83));
    layer0_outputs(709) <= inputs(35);
    layer0_outputs(710) <= '0';
    layer0_outputs(711) <= '0';
    layer0_outputs(712) <= not((inputs(132)) or (inputs(62)));
    layer0_outputs(713) <= not((inputs(40)) xor (inputs(152)));
    layer0_outputs(714) <= not(inputs(52));
    layer0_outputs(715) <= (inputs(129)) or (inputs(110));
    layer0_outputs(716) <= (inputs(61)) or (inputs(23));
    layer0_outputs(717) <= not(inputs(78));
    layer0_outputs(718) <= (inputs(202)) xor (inputs(171));
    layer0_outputs(719) <= not(inputs(40));
    layer0_outputs(720) <= '1';
    layer0_outputs(721) <= not(inputs(199)) or (inputs(81));
    layer0_outputs(722) <= '1';
    layer0_outputs(723) <= (inputs(69)) and not (inputs(55));
    layer0_outputs(724) <= inputs(113);
    layer0_outputs(725) <= not(inputs(118)) or (inputs(218));
    layer0_outputs(726) <= inputs(183);
    layer0_outputs(727) <= not((inputs(53)) or (inputs(248)));
    layer0_outputs(728) <= not(inputs(124));
    layer0_outputs(729) <= '0';
    layer0_outputs(730) <= (inputs(155)) or (inputs(228));
    layer0_outputs(731) <= not(inputs(87));
    layer0_outputs(732) <= '0';
    layer0_outputs(733) <= '0';
    layer0_outputs(734) <= not(inputs(237));
    layer0_outputs(735) <= not((inputs(14)) and (inputs(147)));
    layer0_outputs(736) <= (inputs(170)) and not (inputs(179));
    layer0_outputs(737) <= not(inputs(2));
    layer0_outputs(738) <= not(inputs(168));
    layer0_outputs(739) <= not(inputs(49));
    layer0_outputs(740) <= (inputs(239)) or (inputs(204));
    layer0_outputs(741) <= not(inputs(233));
    layer0_outputs(742) <= '0';
    layer0_outputs(743) <= (inputs(217)) and (inputs(180));
    layer0_outputs(744) <= inputs(23);
    layer0_outputs(745) <= not((inputs(171)) xor (inputs(217)));
    layer0_outputs(746) <= (inputs(244)) or (inputs(59));
    layer0_outputs(747) <= '0';
    layer0_outputs(748) <= (inputs(182)) or (inputs(83));
    layer0_outputs(749) <= not(inputs(133)) or (inputs(17));
    layer0_outputs(750) <= (inputs(180)) and not (inputs(123));
    layer0_outputs(751) <= not(inputs(189)) or (inputs(141));
    layer0_outputs(752) <= not(inputs(16));
    layer0_outputs(753) <= not((inputs(253)) or (inputs(7)));
    layer0_outputs(754) <= inputs(106);
    layer0_outputs(755) <= inputs(113);
    layer0_outputs(756) <= (inputs(127)) or (inputs(128));
    layer0_outputs(757) <= not(inputs(133)) or (inputs(224));
    layer0_outputs(758) <= not(inputs(254)) or (inputs(133));
    layer0_outputs(759) <= (inputs(176)) and (inputs(192));
    layer0_outputs(760) <= '0';
    layer0_outputs(761) <= inputs(82);
    layer0_outputs(762) <= (inputs(224)) and not (inputs(158));
    layer0_outputs(763) <= not((inputs(243)) or (inputs(79)));
    layer0_outputs(764) <= '0';
    layer0_outputs(765) <= not(inputs(104)) or (inputs(186));
    layer0_outputs(766) <= not(inputs(211));
    layer0_outputs(767) <= not(inputs(199));
    layer0_outputs(768) <= (inputs(112)) and not (inputs(248));
    layer0_outputs(769) <= not(inputs(160)) or (inputs(111));
    layer0_outputs(770) <= not((inputs(95)) and (inputs(139)));
    layer0_outputs(771) <= not((inputs(69)) or (inputs(93)));
    layer0_outputs(772) <= inputs(31);
    layer0_outputs(773) <= not((inputs(147)) or (inputs(88)));
    layer0_outputs(774) <= inputs(27);
    layer0_outputs(775) <= not((inputs(237)) and (inputs(118)));
    layer0_outputs(776) <= (inputs(14)) or (inputs(68));
    layer0_outputs(777) <= inputs(21);
    layer0_outputs(778) <= inputs(201);
    layer0_outputs(779) <= inputs(197);
    layer0_outputs(780) <= not((inputs(111)) or (inputs(88)));
    layer0_outputs(781) <= (inputs(32)) or (inputs(21));
    layer0_outputs(782) <= inputs(5);
    layer0_outputs(783) <= (inputs(222)) and (inputs(210));
    layer0_outputs(784) <= not((inputs(146)) or (inputs(206)));
    layer0_outputs(785) <= '1';
    layer0_outputs(786) <= '0';
    layer0_outputs(787) <= (inputs(180)) and not (inputs(166));
    layer0_outputs(788) <= not(inputs(169));
    layer0_outputs(789) <= '1';
    layer0_outputs(790) <= not(inputs(160));
    layer0_outputs(791) <= (inputs(168)) or (inputs(240));
    layer0_outputs(792) <= inputs(235);
    layer0_outputs(793) <= (inputs(68)) and (inputs(150));
    layer0_outputs(794) <= (inputs(61)) or (inputs(77));
    layer0_outputs(795) <= not(inputs(99));
    layer0_outputs(796) <= not((inputs(182)) and (inputs(172)));
    layer0_outputs(797) <= (inputs(222)) and not (inputs(66));
    layer0_outputs(798) <= not(inputs(41)) or (inputs(82));
    layer0_outputs(799) <= not((inputs(215)) and (inputs(87)));
    layer0_outputs(800) <= (inputs(88)) and not (inputs(95));
    layer0_outputs(801) <= not((inputs(120)) or (inputs(82)));
    layer0_outputs(802) <= inputs(48);
    layer0_outputs(803) <= (inputs(10)) or (inputs(246));
    layer0_outputs(804) <= not((inputs(49)) or (inputs(166)));
    layer0_outputs(805) <= not((inputs(174)) and (inputs(12)));
    layer0_outputs(806) <= not((inputs(51)) or (inputs(155)));
    layer0_outputs(807) <= not(inputs(68));
    layer0_outputs(808) <= (inputs(225)) and (inputs(12));
    layer0_outputs(809) <= (inputs(155)) and not (inputs(189));
    layer0_outputs(810) <= not((inputs(251)) or (inputs(66)));
    layer0_outputs(811) <= not(inputs(27));
    layer0_outputs(812) <= not(inputs(104));
    layer0_outputs(813) <= inputs(97);
    layer0_outputs(814) <= not(inputs(104));
    layer0_outputs(815) <= not(inputs(205)) or (inputs(236));
    layer0_outputs(816) <= not(inputs(104)) or (inputs(121));
    layer0_outputs(817) <= not(inputs(249));
    layer0_outputs(818) <= not((inputs(80)) or (inputs(135)));
    layer0_outputs(819) <= inputs(177);
    layer0_outputs(820) <= not(inputs(187));
    layer0_outputs(821) <= (inputs(90)) and not (inputs(133));
    layer0_outputs(822) <= inputs(246);
    layer0_outputs(823) <= not((inputs(232)) and (inputs(41)));
    layer0_outputs(824) <= (inputs(9)) xor (inputs(198));
    layer0_outputs(825) <= not((inputs(118)) or (inputs(162)));
    layer0_outputs(826) <= not((inputs(252)) and (inputs(182)));
    layer0_outputs(827) <= not(inputs(19));
    layer0_outputs(828) <= not(inputs(70));
    layer0_outputs(829) <= '1';
    layer0_outputs(830) <= not(inputs(96)) or (inputs(32));
    layer0_outputs(831) <= not(inputs(142));
    layer0_outputs(832) <= not((inputs(196)) and (inputs(178)));
    layer0_outputs(833) <= not(inputs(151));
    layer0_outputs(834) <= not((inputs(57)) xor (inputs(190)));
    layer0_outputs(835) <= not((inputs(100)) and (inputs(156)));
    layer0_outputs(836) <= '0';
    layer0_outputs(837) <= not((inputs(95)) or (inputs(210)));
    layer0_outputs(838) <= (inputs(194)) or (inputs(223));
    layer0_outputs(839) <= inputs(104);
    layer0_outputs(840) <= (inputs(15)) and not (inputs(184));
    layer0_outputs(841) <= '1';
    layer0_outputs(842) <= (inputs(172)) xor (inputs(222));
    layer0_outputs(843) <= '1';
    layer0_outputs(844) <= '0';
    layer0_outputs(845) <= not(inputs(29));
    layer0_outputs(846) <= not(inputs(51)) or (inputs(205));
    layer0_outputs(847) <= inputs(30);
    layer0_outputs(848) <= '0';
    layer0_outputs(849) <= not(inputs(139)) or (inputs(243));
    layer0_outputs(850) <= not(inputs(5));
    layer0_outputs(851) <= inputs(241);
    layer0_outputs(852) <= '1';
    layer0_outputs(853) <= not(inputs(18)) or (inputs(146));
    layer0_outputs(854) <= '0';
    layer0_outputs(855) <= inputs(243);
    layer0_outputs(856) <= '0';
    layer0_outputs(857) <= not((inputs(46)) xor (inputs(179)));
    layer0_outputs(858) <= (inputs(161)) and not (inputs(150));
    layer0_outputs(859) <= not((inputs(12)) and (inputs(0)));
    layer0_outputs(860) <= '0';
    layer0_outputs(861) <= not((inputs(20)) or (inputs(63)));
    layer0_outputs(862) <= '0';
    layer0_outputs(863) <= (inputs(125)) or (inputs(95));
    layer0_outputs(864) <= (inputs(116)) or (inputs(162));
    layer0_outputs(865) <= (inputs(193)) or (inputs(97));
    layer0_outputs(866) <= (inputs(114)) or (inputs(164));
    layer0_outputs(867) <= (inputs(160)) and not (inputs(216));
    layer0_outputs(868) <= not(inputs(133)) or (inputs(245));
    layer0_outputs(869) <= inputs(78);
    layer0_outputs(870) <= '0';
    layer0_outputs(871) <= not(inputs(10));
    layer0_outputs(872) <= inputs(37);
    layer0_outputs(873) <= inputs(215);
    layer0_outputs(874) <= (inputs(228)) and (inputs(108));
    layer0_outputs(875) <= not(inputs(104));
    layer0_outputs(876) <= inputs(137);
    layer0_outputs(877) <= '0';
    layer0_outputs(878) <= inputs(255);
    layer0_outputs(879) <= not(inputs(63)) or (inputs(234));
    layer0_outputs(880) <= not(inputs(208));
    layer0_outputs(881) <= not((inputs(29)) xor (inputs(33)));
    layer0_outputs(882) <= not(inputs(98));
    layer0_outputs(883) <= not((inputs(251)) and (inputs(132)));
    layer0_outputs(884) <= (inputs(144)) and (inputs(165));
    layer0_outputs(885) <= not((inputs(88)) and (inputs(156)));
    layer0_outputs(886) <= not(inputs(161));
    layer0_outputs(887) <= '1';
    layer0_outputs(888) <= (inputs(174)) or (inputs(222));
    layer0_outputs(889) <= not(inputs(158));
    layer0_outputs(890) <= not(inputs(61));
    layer0_outputs(891) <= (inputs(242)) and not (inputs(91));
    layer0_outputs(892) <= not((inputs(226)) xor (inputs(165)));
    layer0_outputs(893) <= inputs(137);
    layer0_outputs(894) <= (inputs(68)) and not (inputs(61));
    layer0_outputs(895) <= inputs(62);
    layer0_outputs(896) <= not((inputs(205)) or (inputs(175)));
    layer0_outputs(897) <= (inputs(181)) or (inputs(167));
    layer0_outputs(898) <= '1';
    layer0_outputs(899) <= not(inputs(56)) or (inputs(78));
    layer0_outputs(900) <= (inputs(233)) and (inputs(202));
    layer0_outputs(901) <= (inputs(229)) or (inputs(236));
    layer0_outputs(902) <= not((inputs(78)) and (inputs(123)));
    layer0_outputs(903) <= (inputs(55)) and not (inputs(150));
    layer0_outputs(904) <= '1';
    layer0_outputs(905) <= (inputs(44)) and not (inputs(188));
    layer0_outputs(906) <= not((inputs(12)) or (inputs(172)));
    layer0_outputs(907) <= not(inputs(116)) or (inputs(41));
    layer0_outputs(908) <= '1';
    layer0_outputs(909) <= (inputs(227)) and not (inputs(225));
    layer0_outputs(910) <= not((inputs(91)) or (inputs(18)));
    layer0_outputs(911) <= inputs(253);
    layer0_outputs(912) <= not(inputs(229));
    layer0_outputs(913) <= not(inputs(193));
    layer0_outputs(914) <= (inputs(116)) and not (inputs(167));
    layer0_outputs(915) <= (inputs(119)) and not (inputs(20));
    layer0_outputs(916) <= not(inputs(103));
    layer0_outputs(917) <= (inputs(108)) and (inputs(28));
    layer0_outputs(918) <= not(inputs(213));
    layer0_outputs(919) <= not(inputs(255));
    layer0_outputs(920) <= not(inputs(210));
    layer0_outputs(921) <= not(inputs(183)) or (inputs(111));
    layer0_outputs(922) <= '1';
    layer0_outputs(923) <= inputs(99);
    layer0_outputs(924) <= inputs(222);
    layer0_outputs(925) <= '0';
    layer0_outputs(926) <= not(inputs(246));
    layer0_outputs(927) <= (inputs(22)) and not (inputs(196));
    layer0_outputs(928) <= (inputs(188)) or (inputs(225));
    layer0_outputs(929) <= not(inputs(221)) or (inputs(156));
    layer0_outputs(930) <= not(inputs(69));
    layer0_outputs(931) <= (inputs(106)) xor (inputs(38));
    layer0_outputs(932) <= (inputs(42)) and not (inputs(151));
    layer0_outputs(933) <= not((inputs(242)) xor (inputs(114)));
    layer0_outputs(934) <= inputs(161);
    layer0_outputs(935) <= '0';
    layer0_outputs(936) <= inputs(193);
    layer0_outputs(937) <= (inputs(3)) and not (inputs(22));
    layer0_outputs(938) <= (inputs(251)) xor (inputs(125));
    layer0_outputs(939) <= '0';
    layer0_outputs(940) <= inputs(22);
    layer0_outputs(941) <= (inputs(124)) or (inputs(159));
    layer0_outputs(942) <= inputs(11);
    layer0_outputs(943) <= not((inputs(100)) or (inputs(250)));
    layer0_outputs(944) <= '1';
    layer0_outputs(945) <= not(inputs(56)) or (inputs(105));
    layer0_outputs(946) <= '0';
    layer0_outputs(947) <= not(inputs(114));
    layer0_outputs(948) <= not((inputs(44)) or (inputs(88)));
    layer0_outputs(949) <= (inputs(119)) or (inputs(50));
    layer0_outputs(950) <= not((inputs(78)) and (inputs(117)));
    layer0_outputs(951) <= (inputs(177)) or (inputs(96));
    layer0_outputs(952) <= not(inputs(44));
    layer0_outputs(953) <= (inputs(211)) and not (inputs(230));
    layer0_outputs(954) <= inputs(229);
    layer0_outputs(955) <= not((inputs(7)) or (inputs(120)));
    layer0_outputs(956) <= not(inputs(197));
    layer0_outputs(957) <= inputs(242);
    layer0_outputs(958) <= inputs(135);
    layer0_outputs(959) <= not(inputs(93));
    layer0_outputs(960) <= (inputs(126)) or (inputs(146));
    layer0_outputs(961) <= (inputs(190)) or (inputs(171));
    layer0_outputs(962) <= (inputs(146)) and not (inputs(120));
    layer0_outputs(963) <= not(inputs(147)) or (inputs(114));
    layer0_outputs(964) <= inputs(65);
    layer0_outputs(965) <= not(inputs(196));
    layer0_outputs(966) <= inputs(182);
    layer0_outputs(967) <= not((inputs(236)) and (inputs(228)));
    layer0_outputs(968) <= not(inputs(188));
    layer0_outputs(969) <= inputs(147);
    layer0_outputs(970) <= inputs(61);
    layer0_outputs(971) <= not(inputs(93)) or (inputs(174));
    layer0_outputs(972) <= (inputs(172)) and (inputs(183));
    layer0_outputs(973) <= not((inputs(252)) and (inputs(205)));
    layer0_outputs(974) <= (inputs(30)) or (inputs(182));
    layer0_outputs(975) <= (inputs(148)) and not (inputs(190));
    layer0_outputs(976) <= '0';
    layer0_outputs(977) <= (inputs(145)) or (inputs(231));
    layer0_outputs(978) <= (inputs(229)) and not (inputs(163));
    layer0_outputs(979) <= not((inputs(131)) or (inputs(239)));
    layer0_outputs(980) <= (inputs(230)) and not (inputs(135));
    layer0_outputs(981) <= inputs(30);
    layer0_outputs(982) <= not((inputs(48)) or (inputs(29)));
    layer0_outputs(983) <= not(inputs(225));
    layer0_outputs(984) <= not((inputs(124)) xor (inputs(89)));
    layer0_outputs(985) <= not(inputs(75));
    layer0_outputs(986) <= not((inputs(148)) or (inputs(25)));
    layer0_outputs(987) <= (inputs(112)) or (inputs(178));
    layer0_outputs(988) <= not(inputs(182)) or (inputs(44));
    layer0_outputs(989) <= not(inputs(11)) or (inputs(235));
    layer0_outputs(990) <= not(inputs(16)) or (inputs(174));
    layer0_outputs(991) <= not(inputs(220)) or (inputs(253));
    layer0_outputs(992) <= (inputs(79)) or (inputs(26));
    layer0_outputs(993) <= not((inputs(112)) or (inputs(222)));
    layer0_outputs(994) <= '1';
    layer0_outputs(995) <= '1';
    layer0_outputs(996) <= not((inputs(232)) or (inputs(220)));
    layer0_outputs(997) <= inputs(93);
    layer0_outputs(998) <= not(inputs(29));
    layer0_outputs(999) <= not(inputs(45));
    layer0_outputs(1000) <= not((inputs(103)) xor (inputs(243)));
    layer0_outputs(1001) <= not((inputs(11)) or (inputs(60)));
    layer0_outputs(1002) <= (inputs(63)) and not (inputs(172));
    layer0_outputs(1003) <= not((inputs(31)) or (inputs(74)));
    layer0_outputs(1004) <= '1';
    layer0_outputs(1005) <= (inputs(61)) xor (inputs(90));
    layer0_outputs(1006) <= inputs(235);
    layer0_outputs(1007) <= (inputs(19)) and not (inputs(255));
    layer0_outputs(1008) <= not(inputs(70)) or (inputs(41));
    layer0_outputs(1009) <= (inputs(13)) xor (inputs(80));
    layer0_outputs(1010) <= (inputs(23)) and not (inputs(124));
    layer0_outputs(1011) <= (inputs(111)) or (inputs(99));
    layer0_outputs(1012) <= not((inputs(96)) and (inputs(190)));
    layer0_outputs(1013) <= (inputs(46)) and not (inputs(94));
    layer0_outputs(1014) <= (inputs(54)) and (inputs(178));
    layer0_outputs(1015) <= '0';
    layer0_outputs(1016) <= '0';
    layer0_outputs(1017) <= not(inputs(163));
    layer0_outputs(1018) <= '1';
    layer0_outputs(1019) <= (inputs(168)) and (inputs(218));
    layer0_outputs(1020) <= '0';
    layer0_outputs(1021) <= not(inputs(80));
    layer0_outputs(1022) <= not(inputs(159)) or (inputs(155));
    layer0_outputs(1023) <= not((inputs(196)) or (inputs(88)));
    layer0_outputs(1024) <= not(inputs(42));
    layer0_outputs(1025) <= (inputs(220)) and (inputs(82));
    layer0_outputs(1026) <= inputs(108);
    layer0_outputs(1027) <= inputs(80);
    layer0_outputs(1028) <= not(inputs(158)) or (inputs(178));
    layer0_outputs(1029) <= not((inputs(146)) or (inputs(147)));
    layer0_outputs(1030) <= not(inputs(23));
    layer0_outputs(1031) <= '0';
    layer0_outputs(1032) <= not(inputs(146));
    layer0_outputs(1033) <= '1';
    layer0_outputs(1034) <= (inputs(13)) or (inputs(15));
    layer0_outputs(1035) <= (inputs(161)) or (inputs(170));
    layer0_outputs(1036) <= not((inputs(11)) and (inputs(104)));
    layer0_outputs(1037) <= '0';
    layer0_outputs(1038) <= not(inputs(231));
    layer0_outputs(1039) <= not((inputs(103)) or (inputs(240)));
    layer0_outputs(1040) <= (inputs(199)) and not (inputs(210));
    layer0_outputs(1041) <= '1';
    layer0_outputs(1042) <= (inputs(152)) or (inputs(149));
    layer0_outputs(1043) <= not((inputs(173)) or (inputs(11)));
    layer0_outputs(1044) <= not((inputs(154)) xor (inputs(130)));
    layer0_outputs(1045) <= inputs(250);
    layer0_outputs(1046) <= not(inputs(48)) or (inputs(32));
    layer0_outputs(1047) <= (inputs(217)) or (inputs(212));
    layer0_outputs(1048) <= '0';
    layer0_outputs(1049) <= '1';
    layer0_outputs(1050) <= not(inputs(44));
    layer0_outputs(1051) <= not((inputs(217)) or (inputs(47)));
    layer0_outputs(1052) <= not(inputs(248)) or (inputs(195));
    layer0_outputs(1053) <= (inputs(144)) and not (inputs(172));
    layer0_outputs(1054) <= (inputs(203)) or (inputs(17));
    layer0_outputs(1055) <= (inputs(240)) and (inputs(37));
    layer0_outputs(1056) <= inputs(70);
    layer0_outputs(1057) <= not((inputs(206)) xor (inputs(210)));
    layer0_outputs(1058) <= not(inputs(216)) or (inputs(159));
    layer0_outputs(1059) <= (inputs(57)) and not (inputs(152));
    layer0_outputs(1060) <= (inputs(204)) and not (inputs(104));
    layer0_outputs(1061) <= not(inputs(28)) or (inputs(216));
    layer0_outputs(1062) <= not((inputs(123)) and (inputs(36)));
    layer0_outputs(1063) <= not(inputs(23));
    layer0_outputs(1064) <= not((inputs(240)) or (inputs(156)));
    layer0_outputs(1065) <= not(inputs(240));
    layer0_outputs(1066) <= not(inputs(153));
    layer0_outputs(1067) <= '0';
    layer0_outputs(1068) <= inputs(75);
    layer0_outputs(1069) <= not((inputs(245)) xor (inputs(148)));
    layer0_outputs(1070) <= not(inputs(95));
    layer0_outputs(1071) <= inputs(0);
    layer0_outputs(1072) <= not((inputs(182)) or (inputs(211)));
    layer0_outputs(1073) <= '0';
    layer0_outputs(1074) <= not((inputs(8)) or (inputs(11)));
    layer0_outputs(1075) <= '0';
    layer0_outputs(1076) <= not(inputs(102));
    layer0_outputs(1077) <= inputs(83);
    layer0_outputs(1078) <= not(inputs(200)) or (inputs(75));
    layer0_outputs(1079) <= inputs(103);
    layer0_outputs(1080) <= (inputs(206)) or (inputs(104));
    layer0_outputs(1081) <= (inputs(97)) or (inputs(96));
    layer0_outputs(1082) <= (inputs(120)) and not (inputs(69));
    layer0_outputs(1083) <= '1';
    layer0_outputs(1084) <= not(inputs(62)) or (inputs(147));
    layer0_outputs(1085) <= (inputs(243)) and not (inputs(0));
    layer0_outputs(1086) <= (inputs(155)) and not (inputs(176));
    layer0_outputs(1087) <= (inputs(67)) or (inputs(29));
    layer0_outputs(1088) <= inputs(195);
    layer0_outputs(1089) <= (inputs(73)) and not (inputs(38));
    layer0_outputs(1090) <= not((inputs(171)) or (inputs(65)));
    layer0_outputs(1091) <= not(inputs(10));
    layer0_outputs(1092) <= '1';
    layer0_outputs(1093) <= (inputs(116)) and (inputs(240));
    layer0_outputs(1094) <= not(inputs(19));
    layer0_outputs(1095) <= not(inputs(10)) or (inputs(240));
    layer0_outputs(1096) <= '1';
    layer0_outputs(1097) <= not((inputs(63)) or (inputs(30)));
    layer0_outputs(1098) <= (inputs(158)) and (inputs(51));
    layer0_outputs(1099) <= (inputs(151)) and (inputs(216));
    layer0_outputs(1100) <= '1';
    layer0_outputs(1101) <= not(inputs(194));
    layer0_outputs(1102) <= not((inputs(246)) or (inputs(121)));
    layer0_outputs(1103) <= not(inputs(13));
    layer0_outputs(1104) <= (inputs(180)) xor (inputs(129));
    layer0_outputs(1105) <= not(inputs(61)) or (inputs(50));
    layer0_outputs(1106) <= '1';
    layer0_outputs(1107) <= inputs(61);
    layer0_outputs(1108) <= '0';
    layer0_outputs(1109) <= inputs(158);
    layer0_outputs(1110) <= (inputs(119)) and (inputs(41));
    layer0_outputs(1111) <= (inputs(140)) or (inputs(131));
    layer0_outputs(1112) <= (inputs(227)) or (inputs(220));
    layer0_outputs(1113) <= not(inputs(187));
    layer0_outputs(1114) <= inputs(59);
    layer0_outputs(1115) <= not(inputs(218)) or (inputs(58));
    layer0_outputs(1116) <= inputs(155);
    layer0_outputs(1117) <= (inputs(53)) and not (inputs(169));
    layer0_outputs(1118) <= not(inputs(41));
    layer0_outputs(1119) <= '1';
    layer0_outputs(1120) <= '1';
    layer0_outputs(1121) <= inputs(10);
    layer0_outputs(1122) <= inputs(14);
    layer0_outputs(1123) <= inputs(118);
    layer0_outputs(1124) <= '0';
    layer0_outputs(1125) <= '1';
    layer0_outputs(1126) <= inputs(123);
    layer0_outputs(1127) <= not(inputs(188));
    layer0_outputs(1128) <= (inputs(117)) and not (inputs(57));
    layer0_outputs(1129) <= '1';
    layer0_outputs(1130) <= (inputs(209)) or (inputs(80));
    layer0_outputs(1131) <= '1';
    layer0_outputs(1132) <= not((inputs(254)) or (inputs(129)));
    layer0_outputs(1133) <= not(inputs(134)) or (inputs(153));
    layer0_outputs(1134) <= inputs(225);
    layer0_outputs(1135) <= (inputs(125)) or (inputs(177));
    layer0_outputs(1136) <= '1';
    layer0_outputs(1137) <= '0';
    layer0_outputs(1138) <= '1';
    layer0_outputs(1139) <= (inputs(138)) and not (inputs(159));
    layer0_outputs(1140) <= (inputs(183)) xor (inputs(66));
    layer0_outputs(1141) <= '0';
    layer0_outputs(1142) <= not(inputs(30));
    layer0_outputs(1143) <= not((inputs(132)) and (inputs(108)));
    layer0_outputs(1144) <= (inputs(3)) or (inputs(1));
    layer0_outputs(1145) <= inputs(129);
    layer0_outputs(1146) <= not(inputs(208)) or (inputs(231));
    layer0_outputs(1147) <= not(inputs(235)) or (inputs(194));
    layer0_outputs(1148) <= not((inputs(53)) or (inputs(129)));
    layer0_outputs(1149) <= '0';
    layer0_outputs(1150) <= '1';
    layer0_outputs(1151) <= not(inputs(63));
    layer0_outputs(1152) <= not((inputs(141)) or (inputs(84)));
    layer0_outputs(1153) <= not(inputs(58));
    layer0_outputs(1154) <= inputs(157);
    layer0_outputs(1155) <= not((inputs(207)) or (inputs(175)));
    layer0_outputs(1156) <= not(inputs(153)) or (inputs(41));
    layer0_outputs(1157) <= (inputs(29)) and not (inputs(27));
    layer0_outputs(1158) <= not(inputs(165));
    layer0_outputs(1159) <= (inputs(141)) or (inputs(177));
    layer0_outputs(1160) <= not(inputs(228));
    layer0_outputs(1161) <= (inputs(191)) or (inputs(238));
    layer0_outputs(1162) <= not(inputs(210)) or (inputs(3));
    layer0_outputs(1163) <= inputs(96);
    layer0_outputs(1164) <= not(inputs(86));
    layer0_outputs(1165) <= (inputs(207)) and not (inputs(231));
    layer0_outputs(1166) <= (inputs(100)) and (inputs(100));
    layer0_outputs(1167) <= not(inputs(130));
    layer0_outputs(1168) <= not((inputs(105)) or (inputs(4)));
    layer0_outputs(1169) <= not((inputs(178)) and (inputs(250)));
    layer0_outputs(1170) <= not((inputs(54)) and (inputs(55)));
    layer0_outputs(1171) <= '0';
    layer0_outputs(1172) <= (inputs(182)) or (inputs(25));
    layer0_outputs(1173) <= (inputs(168)) and not (inputs(44));
    layer0_outputs(1174) <= inputs(89);
    layer0_outputs(1175) <= not(inputs(240));
    layer0_outputs(1176) <= inputs(57);
    layer0_outputs(1177) <= '0';
    layer0_outputs(1178) <= (inputs(85)) or (inputs(205));
    layer0_outputs(1179) <= '0';
    layer0_outputs(1180) <= (inputs(251)) and not (inputs(232));
    layer0_outputs(1181) <= '1';
    layer0_outputs(1182) <= (inputs(196)) and (inputs(233));
    layer0_outputs(1183) <= not((inputs(199)) and (inputs(187)));
    layer0_outputs(1184) <= not(inputs(32)) or (inputs(140));
    layer0_outputs(1185) <= (inputs(223)) or (inputs(237));
    layer0_outputs(1186) <= not((inputs(117)) and (inputs(102)));
    layer0_outputs(1187) <= not(inputs(7));
    layer0_outputs(1188) <= '1';
    layer0_outputs(1189) <= (inputs(180)) or (inputs(249));
    layer0_outputs(1190) <= not(inputs(238));
    layer0_outputs(1191) <= not((inputs(188)) or (inputs(12)));
    layer0_outputs(1192) <= not((inputs(144)) or (inputs(145)));
    layer0_outputs(1193) <= not((inputs(221)) or (inputs(17)));
    layer0_outputs(1194) <= not(inputs(79));
    layer0_outputs(1195) <= (inputs(74)) and (inputs(96));
    layer0_outputs(1196) <= not(inputs(169));
    layer0_outputs(1197) <= (inputs(117)) and not (inputs(191));
    layer0_outputs(1198) <= inputs(130);
    layer0_outputs(1199) <= not(inputs(93));
    layer0_outputs(1200) <= (inputs(65)) xor (inputs(190));
    layer0_outputs(1201) <= (inputs(83)) or (inputs(81));
    layer0_outputs(1202) <= not((inputs(134)) or (inputs(234)));
    layer0_outputs(1203) <= (inputs(113)) and not (inputs(153));
    layer0_outputs(1204) <= not(inputs(28));
    layer0_outputs(1205) <= inputs(239);
    layer0_outputs(1206) <= not(inputs(79)) or (inputs(176));
    layer0_outputs(1207) <= not((inputs(28)) or (inputs(87)));
    layer0_outputs(1208) <= not(inputs(100)) or (inputs(143));
    layer0_outputs(1209) <= (inputs(87)) and not (inputs(223));
    layer0_outputs(1210) <= '1';
    layer0_outputs(1211) <= '1';
    layer0_outputs(1212) <= inputs(114);
    layer0_outputs(1213) <= not(inputs(35)) or (inputs(130));
    layer0_outputs(1214) <= not(inputs(1));
    layer0_outputs(1215) <= inputs(232);
    layer0_outputs(1216) <= not(inputs(173)) or (inputs(153));
    layer0_outputs(1217) <= '0';
    layer0_outputs(1218) <= not(inputs(172));
    layer0_outputs(1219) <= not(inputs(121));
    layer0_outputs(1220) <= inputs(67);
    layer0_outputs(1221) <= not((inputs(33)) or (inputs(152)));
    layer0_outputs(1222) <= '0';
    layer0_outputs(1223) <= (inputs(172)) and not (inputs(230));
    layer0_outputs(1224) <= not(inputs(200));
    layer0_outputs(1225) <= '0';
    layer0_outputs(1226) <= (inputs(113)) or (inputs(173));
    layer0_outputs(1227) <= (inputs(102)) and (inputs(157));
    layer0_outputs(1228) <= not(inputs(71)) or (inputs(14));
    layer0_outputs(1229) <= not(inputs(146));
    layer0_outputs(1230) <= not((inputs(207)) xor (inputs(193)));
    layer0_outputs(1231) <= not(inputs(52));
    layer0_outputs(1232) <= not((inputs(201)) or (inputs(36)));
    layer0_outputs(1233) <= '1';
    layer0_outputs(1234) <= not(inputs(40));
    layer0_outputs(1235) <= not(inputs(134));
    layer0_outputs(1236) <= not((inputs(42)) xor (inputs(188)));
    layer0_outputs(1237) <= inputs(141);
    layer0_outputs(1238) <= inputs(239);
    layer0_outputs(1239) <= not((inputs(226)) xor (inputs(211)));
    layer0_outputs(1240) <= (inputs(165)) or (inputs(53));
    layer0_outputs(1241) <= not((inputs(110)) or (inputs(84)));
    layer0_outputs(1242) <= (inputs(255)) and not (inputs(112));
    layer0_outputs(1243) <= not(inputs(189));
    layer0_outputs(1244) <= (inputs(114)) and not (inputs(122));
    layer0_outputs(1245) <= not(inputs(246));
    layer0_outputs(1246) <= inputs(239);
    layer0_outputs(1247) <= (inputs(184)) and not (inputs(124));
    layer0_outputs(1248) <= not(inputs(241)) or (inputs(104));
    layer0_outputs(1249) <= '1';
    layer0_outputs(1250) <= (inputs(237)) or (inputs(180));
    layer0_outputs(1251) <= inputs(15);
    layer0_outputs(1252) <= '0';
    layer0_outputs(1253) <= (inputs(77)) or (inputs(99));
    layer0_outputs(1254) <= (inputs(21)) and (inputs(251));
    layer0_outputs(1255) <= (inputs(202)) and not (inputs(127));
    layer0_outputs(1256) <= not((inputs(20)) and (inputs(237)));
    layer0_outputs(1257) <= inputs(193);
    layer0_outputs(1258) <= not(inputs(123)) or (inputs(60));
    layer0_outputs(1259) <= not((inputs(254)) and (inputs(61)));
    layer0_outputs(1260) <= inputs(56);
    layer0_outputs(1261) <= not(inputs(199));
    layer0_outputs(1262) <= not((inputs(102)) or (inputs(44)));
    layer0_outputs(1263) <= inputs(213);
    layer0_outputs(1264) <= inputs(205);
    layer0_outputs(1265) <= not((inputs(90)) or (inputs(98)));
    layer0_outputs(1266) <= not(inputs(1));
    layer0_outputs(1267) <= '1';
    layer0_outputs(1268) <= not((inputs(178)) xor (inputs(6)));
    layer0_outputs(1269) <= (inputs(235)) or (inputs(6));
    layer0_outputs(1270) <= (inputs(173)) and not (inputs(71));
    layer0_outputs(1271) <= not(inputs(220)) or (inputs(73));
    layer0_outputs(1272) <= inputs(249);
    layer0_outputs(1273) <= (inputs(31)) or (inputs(210));
    layer0_outputs(1274) <= (inputs(133)) and not (inputs(133));
    layer0_outputs(1275) <= inputs(165);
    layer0_outputs(1276) <= (inputs(116)) or (inputs(146));
    layer0_outputs(1277) <= not(inputs(88));
    layer0_outputs(1278) <= '0';
    layer0_outputs(1279) <= not((inputs(94)) or (inputs(90)));
    layer0_outputs(1280) <= '1';
    layer0_outputs(1281) <= (inputs(182)) and (inputs(42));
    layer0_outputs(1282) <= not(inputs(177)) or (inputs(157));
    layer0_outputs(1283) <= '0';
    layer0_outputs(1284) <= (inputs(208)) and (inputs(112));
    layer0_outputs(1285) <= inputs(229);
    layer0_outputs(1286) <= not(inputs(18)) or (inputs(40));
    layer0_outputs(1287) <= (inputs(247)) and not (inputs(18));
    layer0_outputs(1288) <= not((inputs(100)) and (inputs(16)));
    layer0_outputs(1289) <= inputs(69);
    layer0_outputs(1290) <= not(inputs(60)) or (inputs(235));
    layer0_outputs(1291) <= not(inputs(150)) or (inputs(179));
    layer0_outputs(1292) <= not(inputs(247));
    layer0_outputs(1293) <= not((inputs(27)) and (inputs(230)));
    layer0_outputs(1294) <= not(inputs(136));
    layer0_outputs(1295) <= '0';
    layer0_outputs(1296) <= (inputs(165)) and not (inputs(47));
    layer0_outputs(1297) <= '1';
    layer0_outputs(1298) <= '1';
    layer0_outputs(1299) <= inputs(50);
    layer0_outputs(1300) <= '0';
    layer0_outputs(1301) <= (inputs(204)) and not (inputs(148));
    layer0_outputs(1302) <= not((inputs(232)) or (inputs(196)));
    layer0_outputs(1303) <= '0';
    layer0_outputs(1304) <= inputs(63);
    layer0_outputs(1305) <= (inputs(253)) and (inputs(184));
    layer0_outputs(1306) <= not(inputs(1)) or (inputs(247));
    layer0_outputs(1307) <= '0';
    layer0_outputs(1308) <= '1';
    layer0_outputs(1309) <= inputs(71);
    layer0_outputs(1310) <= inputs(18);
    layer0_outputs(1311) <= not((inputs(216)) or (inputs(170)));
    layer0_outputs(1312) <= not(inputs(219));
    layer0_outputs(1313) <= (inputs(245)) and not (inputs(27));
    layer0_outputs(1314) <= '0';
    layer0_outputs(1315) <= not(inputs(193)) or (inputs(138));
    layer0_outputs(1316) <= not((inputs(15)) and (inputs(166)));
    layer0_outputs(1317) <= '0';
    layer0_outputs(1318) <= (inputs(228)) or (inputs(243));
    layer0_outputs(1319) <= (inputs(21)) or (inputs(142));
    layer0_outputs(1320) <= not(inputs(108));
    layer0_outputs(1321) <= not(inputs(165));
    layer0_outputs(1322) <= (inputs(15)) and not (inputs(163));
    layer0_outputs(1323) <= not((inputs(223)) xor (inputs(234)));
    layer0_outputs(1324) <= (inputs(220)) and not (inputs(0));
    layer0_outputs(1325) <= not(inputs(65)) or (inputs(30));
    layer0_outputs(1326) <= '1';
    layer0_outputs(1327) <= '0';
    layer0_outputs(1328) <= '1';
    layer0_outputs(1329) <= '0';
    layer0_outputs(1330) <= (inputs(215)) or (inputs(7));
    layer0_outputs(1331) <= not((inputs(33)) xor (inputs(222)));
    layer0_outputs(1332) <= not(inputs(233));
    layer0_outputs(1333) <= '1';
    layer0_outputs(1334) <= not(inputs(21)) or (inputs(0));
    layer0_outputs(1335) <= not((inputs(175)) or (inputs(144)));
    layer0_outputs(1336) <= not(inputs(119)) or (inputs(19));
    layer0_outputs(1337) <= not(inputs(148));
    layer0_outputs(1338) <= not(inputs(167)) or (inputs(15));
    layer0_outputs(1339) <= inputs(182);
    layer0_outputs(1340) <= not((inputs(126)) xor (inputs(153)));
    layer0_outputs(1341) <= not(inputs(152));
    layer0_outputs(1342) <= (inputs(144)) xor (inputs(118));
    layer0_outputs(1343) <= inputs(193);
    layer0_outputs(1344) <= inputs(149);
    layer0_outputs(1345) <= '0';
    layer0_outputs(1346) <= not((inputs(221)) or (inputs(146)));
    layer0_outputs(1347) <= not(inputs(101));
    layer0_outputs(1348) <= not((inputs(110)) and (inputs(197)));
    layer0_outputs(1349) <= '1';
    layer0_outputs(1350) <= '1';
    layer0_outputs(1351) <= '1';
    layer0_outputs(1352) <= '0';
    layer0_outputs(1353) <= '0';
    layer0_outputs(1354) <= '1';
    layer0_outputs(1355) <= '1';
    layer0_outputs(1356) <= not((inputs(46)) and (inputs(78)));
    layer0_outputs(1357) <= '0';
    layer0_outputs(1358) <= inputs(107);
    layer0_outputs(1359) <= inputs(133);
    layer0_outputs(1360) <= not((inputs(4)) or (inputs(155)));
    layer0_outputs(1361) <= inputs(118);
    layer0_outputs(1362) <= '0';
    layer0_outputs(1363) <= not(inputs(99)) or (inputs(196));
    layer0_outputs(1364) <= (inputs(66)) and not (inputs(184));
    layer0_outputs(1365) <= (inputs(241)) and not (inputs(21));
    layer0_outputs(1366) <= (inputs(99)) or (inputs(133));
    layer0_outputs(1367) <= not(inputs(221));
    layer0_outputs(1368) <= '1';
    layer0_outputs(1369) <= '0';
    layer0_outputs(1370) <= not(inputs(35));
    layer0_outputs(1371) <= inputs(20);
    layer0_outputs(1372) <= not(inputs(39));
    layer0_outputs(1373) <= inputs(192);
    layer0_outputs(1374) <= (inputs(207)) and (inputs(225));
    layer0_outputs(1375) <= not(inputs(208)) or (inputs(91));
    layer0_outputs(1376) <= '0';
    layer0_outputs(1377) <= (inputs(117)) and not (inputs(157));
    layer0_outputs(1378) <= (inputs(59)) and (inputs(123));
    layer0_outputs(1379) <= not(inputs(173));
    layer0_outputs(1380) <= '1';
    layer0_outputs(1381) <= (inputs(130)) and not (inputs(239));
    layer0_outputs(1382) <= (inputs(2)) or (inputs(111));
    layer0_outputs(1383) <= not(inputs(40));
    layer0_outputs(1384) <= inputs(95);
    layer0_outputs(1385) <= '0';
    layer0_outputs(1386) <= not((inputs(138)) xor (inputs(160)));
    layer0_outputs(1387) <= (inputs(42)) and not (inputs(68));
    layer0_outputs(1388) <= '0';
    layer0_outputs(1389) <= '0';
    layer0_outputs(1390) <= not(inputs(56)) or (inputs(219));
    layer0_outputs(1391) <= not(inputs(134));
    layer0_outputs(1392) <= not(inputs(59)) or (inputs(200));
    layer0_outputs(1393) <= not(inputs(139));
    layer0_outputs(1394) <= not((inputs(176)) and (inputs(241)));
    layer0_outputs(1395) <= not(inputs(42));
    layer0_outputs(1396) <= '1';
    layer0_outputs(1397) <= not(inputs(90));
    layer0_outputs(1398) <= not(inputs(74));
    layer0_outputs(1399) <= not(inputs(93));
    layer0_outputs(1400) <= inputs(133);
    layer0_outputs(1401) <= '0';
    layer0_outputs(1402) <= (inputs(92)) or (inputs(138));
    layer0_outputs(1403) <= '0';
    layer0_outputs(1404) <= not(inputs(111)) or (inputs(242));
    layer0_outputs(1405) <= '0';
    layer0_outputs(1406) <= (inputs(208)) or (inputs(117));
    layer0_outputs(1407) <= (inputs(30)) or (inputs(12));
    layer0_outputs(1408) <= (inputs(30)) and (inputs(57));
    layer0_outputs(1409) <= not((inputs(21)) or (inputs(142)));
    layer0_outputs(1410) <= not(inputs(56));
    layer0_outputs(1411) <= not((inputs(65)) and (inputs(224)));
    layer0_outputs(1412) <= not((inputs(1)) and (inputs(76)));
    layer0_outputs(1413) <= inputs(193);
    layer0_outputs(1414) <= '1';
    layer0_outputs(1415) <= (inputs(242)) and (inputs(255));
    layer0_outputs(1416) <= not(inputs(239));
    layer0_outputs(1417) <= not((inputs(225)) and (inputs(1)));
    layer0_outputs(1418) <= '1';
    layer0_outputs(1419) <= (inputs(63)) and not (inputs(248));
    layer0_outputs(1420) <= '0';
    layer0_outputs(1421) <= '0';
    layer0_outputs(1422) <= inputs(154);
    layer0_outputs(1423) <= not(inputs(164));
    layer0_outputs(1424) <= (inputs(203)) and not (inputs(99));
    layer0_outputs(1425) <= '0';
    layer0_outputs(1426) <= not(inputs(84)) or (inputs(184));
    layer0_outputs(1427) <= not((inputs(196)) and (inputs(26)));
    layer0_outputs(1428) <= not(inputs(70)) or (inputs(206));
    layer0_outputs(1429) <= not((inputs(226)) and (inputs(72)));
    layer0_outputs(1430) <= (inputs(156)) or (inputs(190));
    layer0_outputs(1431) <= not(inputs(182)) or (inputs(227));
    layer0_outputs(1432) <= not(inputs(52)) or (inputs(112));
    layer0_outputs(1433) <= not(inputs(7)) or (inputs(145));
    layer0_outputs(1434) <= not(inputs(19));
    layer0_outputs(1435) <= inputs(200);
    layer0_outputs(1436) <= inputs(100);
    layer0_outputs(1437) <= '1';
    layer0_outputs(1438) <= not(inputs(139));
    layer0_outputs(1439) <= not(inputs(88)) or (inputs(136));
    layer0_outputs(1440) <= (inputs(42)) or (inputs(117));
    layer0_outputs(1441) <= not(inputs(227));
    layer0_outputs(1442) <= '1';
    layer0_outputs(1443) <= not(inputs(239));
    layer0_outputs(1444) <= inputs(165);
    layer0_outputs(1445) <= (inputs(147)) or (inputs(154));
    layer0_outputs(1446) <= '0';
    layer0_outputs(1447) <= inputs(103);
    layer0_outputs(1448) <= not((inputs(44)) or (inputs(63)));
    layer0_outputs(1449) <= not(inputs(18));
    layer0_outputs(1450) <= (inputs(41)) or (inputs(0));
    layer0_outputs(1451) <= '0';
    layer0_outputs(1452) <= '0';
    layer0_outputs(1453) <= (inputs(155)) and (inputs(166));
    layer0_outputs(1454) <= not(inputs(214));
    layer0_outputs(1455) <= not(inputs(72));
    layer0_outputs(1456) <= inputs(92);
    layer0_outputs(1457) <= not(inputs(211)) or (inputs(44));
    layer0_outputs(1458) <= not(inputs(211));
    layer0_outputs(1459) <= not(inputs(43)) or (inputs(101));
    layer0_outputs(1460) <= not(inputs(63));
    layer0_outputs(1461) <= not(inputs(85));
    layer0_outputs(1462) <= not(inputs(119)) or (inputs(4));
    layer0_outputs(1463) <= not(inputs(235));
    layer0_outputs(1464) <= '0';
    layer0_outputs(1465) <= (inputs(113)) and (inputs(215));
    layer0_outputs(1466) <= (inputs(248)) and (inputs(213));
    layer0_outputs(1467) <= (inputs(42)) or (inputs(87));
    layer0_outputs(1468) <= (inputs(174)) or (inputs(0));
    layer0_outputs(1469) <= not(inputs(246)) or (inputs(80));
    layer0_outputs(1470) <= not(inputs(141)) or (inputs(64));
    layer0_outputs(1471) <= not(inputs(136));
    layer0_outputs(1472) <= not(inputs(143)) or (inputs(61));
    layer0_outputs(1473) <= not((inputs(76)) and (inputs(63)));
    layer0_outputs(1474) <= inputs(203);
    layer0_outputs(1475) <= (inputs(54)) and (inputs(224));
    layer0_outputs(1476) <= inputs(98);
    layer0_outputs(1477) <= not(inputs(61));
    layer0_outputs(1478) <= not(inputs(191)) or (inputs(188));
    layer0_outputs(1479) <= not(inputs(25));
    layer0_outputs(1480) <= (inputs(6)) and (inputs(129));
    layer0_outputs(1481) <= not((inputs(122)) or (inputs(110)));
    layer0_outputs(1482) <= not((inputs(140)) or (inputs(26)));
    layer0_outputs(1483) <= inputs(102);
    layer0_outputs(1484) <= (inputs(236)) and (inputs(200));
    layer0_outputs(1485) <= inputs(114);
    layer0_outputs(1486) <= (inputs(250)) or (inputs(65));
    layer0_outputs(1487) <= '1';
    layer0_outputs(1488) <= (inputs(146)) and not (inputs(45));
    layer0_outputs(1489) <= not(inputs(126));
    layer0_outputs(1490) <= '0';
    layer0_outputs(1491) <= (inputs(176)) and (inputs(111));
    layer0_outputs(1492) <= (inputs(104)) and not (inputs(50));
    layer0_outputs(1493) <= inputs(49);
    layer0_outputs(1494) <= (inputs(142)) and (inputs(81));
    layer0_outputs(1495) <= '1';
    layer0_outputs(1496) <= not(inputs(77));
    layer0_outputs(1497) <= inputs(194);
    layer0_outputs(1498) <= '1';
    layer0_outputs(1499) <= inputs(146);
    layer0_outputs(1500) <= not((inputs(15)) xor (inputs(85)));
    layer0_outputs(1501) <= inputs(231);
    layer0_outputs(1502) <= not(inputs(48));
    layer0_outputs(1503) <= not(inputs(126));
    layer0_outputs(1504) <= not(inputs(163));
    layer0_outputs(1505) <= (inputs(146)) and not (inputs(209));
    layer0_outputs(1506) <= (inputs(17)) or (inputs(140));
    layer0_outputs(1507) <= (inputs(134)) and not (inputs(223));
    layer0_outputs(1508) <= (inputs(211)) and not (inputs(78));
    layer0_outputs(1509) <= not(inputs(53)) or (inputs(27));
    layer0_outputs(1510) <= (inputs(170)) or (inputs(155));
    layer0_outputs(1511) <= (inputs(226)) or (inputs(147));
    layer0_outputs(1512) <= inputs(74);
    layer0_outputs(1513) <= not(inputs(89)) or (inputs(50));
    layer0_outputs(1514) <= not(inputs(54));
    layer0_outputs(1515) <= (inputs(112)) and not (inputs(66));
    layer0_outputs(1516) <= (inputs(188)) or (inputs(204));
    layer0_outputs(1517) <= (inputs(103)) and not (inputs(98));
    layer0_outputs(1518) <= (inputs(67)) xor (inputs(176));
    layer0_outputs(1519) <= not((inputs(179)) or (inputs(225)));
    layer0_outputs(1520) <= (inputs(26)) or (inputs(251));
    layer0_outputs(1521) <= not(inputs(74));
    layer0_outputs(1522) <= inputs(221);
    layer0_outputs(1523) <= (inputs(245)) or (inputs(193));
    layer0_outputs(1524) <= (inputs(194)) and not (inputs(15));
    layer0_outputs(1525) <= not(inputs(194));
    layer0_outputs(1526) <= inputs(227);
    layer0_outputs(1527) <= not(inputs(239));
    layer0_outputs(1528) <= not((inputs(24)) or (inputs(65)));
    layer0_outputs(1529) <= inputs(131);
    layer0_outputs(1530) <= '1';
    layer0_outputs(1531) <= (inputs(254)) xor (inputs(59));
    layer0_outputs(1532) <= not(inputs(75));
    layer0_outputs(1533) <= (inputs(41)) and not (inputs(0));
    layer0_outputs(1534) <= inputs(87);
    layer0_outputs(1535) <= not((inputs(198)) or (inputs(87)));
    layer0_outputs(1536) <= not(inputs(39));
    layer0_outputs(1537) <= inputs(191);
    layer0_outputs(1538) <= not((inputs(14)) and (inputs(96)));
    layer0_outputs(1539) <= (inputs(109)) and not (inputs(133));
    layer0_outputs(1540) <= not(inputs(171)) or (inputs(64));
    layer0_outputs(1541) <= inputs(120);
    layer0_outputs(1542) <= (inputs(186)) and (inputs(124));
    layer0_outputs(1543) <= (inputs(217)) and not (inputs(29));
    layer0_outputs(1544) <= (inputs(210)) or (inputs(210));
    layer0_outputs(1545) <= (inputs(88)) and (inputs(242));
    layer0_outputs(1546) <= not(inputs(72)) or (inputs(0));
    layer0_outputs(1547) <= not(inputs(31)) or (inputs(31));
    layer0_outputs(1548) <= not((inputs(109)) or (inputs(177)));
    layer0_outputs(1549) <= not((inputs(155)) xor (inputs(185)));
    layer0_outputs(1550) <= (inputs(177)) or (inputs(204));
    layer0_outputs(1551) <= not(inputs(57));
    layer0_outputs(1552) <= '1';
    layer0_outputs(1553) <= not((inputs(94)) or (inputs(100)));
    layer0_outputs(1554) <= (inputs(15)) and not (inputs(149));
    layer0_outputs(1555) <= not(inputs(53));
    layer0_outputs(1556) <= '1';
    layer0_outputs(1557) <= (inputs(98)) and not (inputs(51));
    layer0_outputs(1558) <= '1';
    layer0_outputs(1559) <= (inputs(255)) and (inputs(42));
    layer0_outputs(1560) <= not(inputs(172)) or (inputs(85));
    layer0_outputs(1561) <= (inputs(45)) xor (inputs(11));
    layer0_outputs(1562) <= not((inputs(175)) and (inputs(208)));
    layer0_outputs(1563) <= not(inputs(207)) or (inputs(127));
    layer0_outputs(1564) <= inputs(114);
    layer0_outputs(1565) <= (inputs(97)) or (inputs(141));
    layer0_outputs(1566) <= '0';
    layer0_outputs(1567) <= not(inputs(158)) or (inputs(57));
    layer0_outputs(1568) <= (inputs(74)) or (inputs(77));
    layer0_outputs(1569) <= (inputs(106)) and (inputs(115));
    layer0_outputs(1570) <= not(inputs(223)) or (inputs(140));
    layer0_outputs(1571) <= (inputs(99)) and not (inputs(220));
    layer0_outputs(1572) <= '0';
    layer0_outputs(1573) <= not(inputs(84));
    layer0_outputs(1574) <= not((inputs(223)) or (inputs(196)));
    layer0_outputs(1575) <= (inputs(3)) and (inputs(140));
    layer0_outputs(1576) <= not(inputs(190));
    layer0_outputs(1577) <= not((inputs(197)) and (inputs(247)));
    layer0_outputs(1578) <= not((inputs(126)) or (inputs(207)));
    layer0_outputs(1579) <= '0';
    layer0_outputs(1580) <= not(inputs(132));
    layer0_outputs(1581) <= inputs(158);
    layer0_outputs(1582) <= not((inputs(211)) and (inputs(92)));
    layer0_outputs(1583) <= not(inputs(98));
    layer0_outputs(1584) <= '1';
    layer0_outputs(1585) <= not(inputs(75)) or (inputs(160));
    layer0_outputs(1586) <= not((inputs(85)) and (inputs(49)));
    layer0_outputs(1587) <= (inputs(170)) or (inputs(148));
    layer0_outputs(1588) <= not((inputs(187)) or (inputs(229)));
    layer0_outputs(1589) <= not(inputs(60));
    layer0_outputs(1590) <= (inputs(161)) and not (inputs(184));
    layer0_outputs(1591) <= (inputs(153)) and not (inputs(10));
    layer0_outputs(1592) <= '0';
    layer0_outputs(1593) <= inputs(243);
    layer0_outputs(1594) <= not(inputs(24)) or (inputs(17));
    layer0_outputs(1595) <= not(inputs(89)) or (inputs(170));
    layer0_outputs(1596) <= not((inputs(192)) or (inputs(37)));
    layer0_outputs(1597) <= not(inputs(35));
    layer0_outputs(1598) <= '1';
    layer0_outputs(1599) <= inputs(23);
    layer0_outputs(1600) <= not((inputs(36)) and (inputs(13)));
    layer0_outputs(1601) <= '1';
    layer0_outputs(1602) <= not((inputs(105)) or (inputs(97)));
    layer0_outputs(1603) <= not(inputs(234));
    layer0_outputs(1604) <= not(inputs(61)) or (inputs(192));
    layer0_outputs(1605) <= not((inputs(112)) or (inputs(15)));
    layer0_outputs(1606) <= not(inputs(105)) or (inputs(55));
    layer0_outputs(1607) <= not(inputs(75));
    layer0_outputs(1608) <= (inputs(241)) and not (inputs(153));
    layer0_outputs(1609) <= (inputs(108)) and not (inputs(128));
    layer0_outputs(1610) <= not(inputs(21));
    layer0_outputs(1611) <= not(inputs(100));
    layer0_outputs(1612) <= not(inputs(37));
    layer0_outputs(1613) <= inputs(240);
    layer0_outputs(1614) <= (inputs(7)) and not (inputs(200));
    layer0_outputs(1615) <= not((inputs(23)) or (inputs(84)));
    layer0_outputs(1616) <= inputs(58);
    layer0_outputs(1617) <= not(inputs(123));
    layer0_outputs(1618) <= (inputs(23)) and (inputs(150));
    layer0_outputs(1619) <= not(inputs(137));
    layer0_outputs(1620) <= '1';
    layer0_outputs(1621) <= not(inputs(145));
    layer0_outputs(1622) <= not(inputs(38)) or (inputs(192));
    layer0_outputs(1623) <= '1';
    layer0_outputs(1624) <= not(inputs(94));
    layer0_outputs(1625) <= '1';
    layer0_outputs(1626) <= (inputs(211)) and not (inputs(121));
    layer0_outputs(1627) <= inputs(66);
    layer0_outputs(1628) <= not((inputs(160)) and (inputs(217)));
    layer0_outputs(1629) <= not(inputs(22));
    layer0_outputs(1630) <= not(inputs(192));
    layer0_outputs(1631) <= (inputs(131)) or (inputs(81));
    layer0_outputs(1632) <= '1';
    layer0_outputs(1633) <= not(inputs(33));
    layer0_outputs(1634) <= not(inputs(151)) or (inputs(209));
    layer0_outputs(1635) <= '0';
    layer0_outputs(1636) <= '1';
    layer0_outputs(1637) <= (inputs(254)) and (inputs(79));
    layer0_outputs(1638) <= inputs(204);
    layer0_outputs(1639) <= not(inputs(24)) or (inputs(109));
    layer0_outputs(1640) <= not((inputs(180)) and (inputs(119)));
    layer0_outputs(1641) <= (inputs(35)) and not (inputs(186));
    layer0_outputs(1642) <= not(inputs(14)) or (inputs(94));
    layer0_outputs(1643) <= (inputs(106)) and (inputs(189));
    layer0_outputs(1644) <= not(inputs(204)) or (inputs(74));
    layer0_outputs(1645) <= not(inputs(161));
    layer0_outputs(1646) <= '1';
    layer0_outputs(1647) <= not((inputs(139)) or (inputs(93)));
    layer0_outputs(1648) <= not((inputs(233)) and (inputs(147)));
    layer0_outputs(1649) <= (inputs(206)) and not (inputs(246));
    layer0_outputs(1650) <= inputs(170);
    layer0_outputs(1651) <= (inputs(29)) or (inputs(83));
    layer0_outputs(1652) <= (inputs(119)) and not (inputs(94));
    layer0_outputs(1653) <= (inputs(176)) and not (inputs(61));
    layer0_outputs(1654) <= not((inputs(187)) or (inputs(113)));
    layer0_outputs(1655) <= not((inputs(76)) or (inputs(92)));
    layer0_outputs(1656) <= '0';
    layer0_outputs(1657) <= not((inputs(71)) xor (inputs(206)));
    layer0_outputs(1658) <= not((inputs(49)) or (inputs(26)));
    layer0_outputs(1659) <= (inputs(85)) and not (inputs(47));
    layer0_outputs(1660) <= '0';
    layer0_outputs(1661) <= not((inputs(108)) and (inputs(166)));
    layer0_outputs(1662) <= not(inputs(142)) or (inputs(28));
    layer0_outputs(1663) <= inputs(32);
    layer0_outputs(1664) <= not(inputs(111)) or (inputs(228));
    layer0_outputs(1665) <= not(inputs(175)) or (inputs(142));
    layer0_outputs(1666) <= not(inputs(83));
    layer0_outputs(1667) <= not(inputs(212)) or (inputs(36));
    layer0_outputs(1668) <= (inputs(51)) and not (inputs(109));
    layer0_outputs(1669) <= not((inputs(244)) or (inputs(248)));
    layer0_outputs(1670) <= inputs(188);
    layer0_outputs(1671) <= not((inputs(81)) and (inputs(10)));
    layer0_outputs(1672) <= not(inputs(33));
    layer0_outputs(1673) <= not(inputs(164));
    layer0_outputs(1674) <= not(inputs(78));
    layer0_outputs(1675) <= '1';
    layer0_outputs(1676) <= '1';
    layer0_outputs(1677) <= not(inputs(119));
    layer0_outputs(1678) <= inputs(25);
    layer0_outputs(1679) <= inputs(253);
    layer0_outputs(1680) <= inputs(187);
    layer0_outputs(1681) <= not((inputs(145)) xor (inputs(216)));
    layer0_outputs(1682) <= (inputs(86)) or (inputs(141));
    layer0_outputs(1683) <= (inputs(225)) or (inputs(220));
    layer0_outputs(1684) <= (inputs(86)) and (inputs(80));
    layer0_outputs(1685) <= inputs(139);
    layer0_outputs(1686) <= not((inputs(84)) and (inputs(247)));
    layer0_outputs(1687) <= (inputs(129)) and not (inputs(45));
    layer0_outputs(1688) <= not(inputs(5)) or (inputs(5));
    layer0_outputs(1689) <= not(inputs(220));
    layer0_outputs(1690) <= not(inputs(248));
    layer0_outputs(1691) <= (inputs(45)) and (inputs(59));
    layer0_outputs(1692) <= not(inputs(242));
    layer0_outputs(1693) <= '1';
    layer0_outputs(1694) <= not(inputs(71)) or (inputs(163));
    layer0_outputs(1695) <= (inputs(162)) and (inputs(189));
    layer0_outputs(1696) <= (inputs(97)) and not (inputs(134));
    layer0_outputs(1697) <= not((inputs(178)) and (inputs(50)));
    layer0_outputs(1698) <= (inputs(43)) or (inputs(175));
    layer0_outputs(1699) <= (inputs(92)) or (inputs(47));
    layer0_outputs(1700) <= (inputs(147)) and not (inputs(61));
    layer0_outputs(1701) <= not(inputs(42));
    layer0_outputs(1702) <= inputs(149);
    layer0_outputs(1703) <= '1';
    layer0_outputs(1704) <= '1';
    layer0_outputs(1705) <= not((inputs(92)) xor (inputs(11)));
    layer0_outputs(1706) <= not((inputs(40)) and (inputs(146)));
    layer0_outputs(1707) <= not((inputs(118)) or (inputs(131)));
    layer0_outputs(1708) <= not(inputs(71)) or (inputs(56));
    layer0_outputs(1709) <= not((inputs(161)) xor (inputs(140)));
    layer0_outputs(1710) <= inputs(151);
    layer0_outputs(1711) <= not(inputs(159));
    layer0_outputs(1712) <= not(inputs(20)) or (inputs(99));
    layer0_outputs(1713) <= inputs(121);
    layer0_outputs(1714) <= not((inputs(86)) and (inputs(27)));
    layer0_outputs(1715) <= (inputs(244)) or (inputs(245));
    layer0_outputs(1716) <= '1';
    layer0_outputs(1717) <= (inputs(78)) or (inputs(79));
    layer0_outputs(1718) <= not((inputs(230)) or (inputs(194)));
    layer0_outputs(1719) <= not(inputs(231)) or (inputs(23));
    layer0_outputs(1720) <= (inputs(211)) or (inputs(185));
    layer0_outputs(1721) <= (inputs(243)) or (inputs(42));
    layer0_outputs(1722) <= not(inputs(97));
    layer0_outputs(1723) <= (inputs(127)) and (inputs(157));
    layer0_outputs(1724) <= not(inputs(17)) or (inputs(26));
    layer0_outputs(1725) <= '0';
    layer0_outputs(1726) <= not((inputs(47)) or (inputs(209)));
    layer0_outputs(1727) <= not(inputs(167));
    layer0_outputs(1728) <= not(inputs(125));
    layer0_outputs(1729) <= inputs(223);
    layer0_outputs(1730) <= not((inputs(155)) or (inputs(139)));
    layer0_outputs(1731) <= '0';
    layer0_outputs(1732) <= not(inputs(135));
    layer0_outputs(1733) <= not((inputs(139)) or (inputs(201)));
    layer0_outputs(1734) <= (inputs(115)) and not (inputs(19));
    layer0_outputs(1735) <= inputs(183);
    layer0_outputs(1736) <= not(inputs(207));
    layer0_outputs(1737) <= '0';
    layer0_outputs(1738) <= inputs(169);
    layer0_outputs(1739) <= (inputs(215)) and (inputs(166));
    layer0_outputs(1740) <= not(inputs(3));
    layer0_outputs(1741) <= (inputs(32)) and not (inputs(22));
    layer0_outputs(1742) <= not(inputs(160));
    layer0_outputs(1743) <= '1';
    layer0_outputs(1744) <= (inputs(238)) or (inputs(156));
    layer0_outputs(1745) <= not(inputs(49)) or (inputs(154));
    layer0_outputs(1746) <= not(inputs(144)) or (inputs(120));
    layer0_outputs(1747) <= (inputs(232)) or (inputs(192));
    layer0_outputs(1748) <= inputs(21);
    layer0_outputs(1749) <= not(inputs(161)) or (inputs(163));
    layer0_outputs(1750) <= not(inputs(148));
    layer0_outputs(1751) <= (inputs(171)) and (inputs(25));
    layer0_outputs(1752) <= not((inputs(244)) or (inputs(240)));
    layer0_outputs(1753) <= inputs(196);
    layer0_outputs(1754) <= '0';
    layer0_outputs(1755) <= (inputs(163)) and not (inputs(76));
    layer0_outputs(1756) <= not((inputs(245)) and (inputs(2)));
    layer0_outputs(1757) <= '1';
    layer0_outputs(1758) <= not((inputs(216)) and (inputs(161)));
    layer0_outputs(1759) <= not((inputs(251)) or (inputs(253)));
    layer0_outputs(1760) <= not(inputs(52));
    layer0_outputs(1761) <= not((inputs(217)) or (inputs(20)));
    layer0_outputs(1762) <= not(inputs(80)) or (inputs(208));
    layer0_outputs(1763) <= inputs(72);
    layer0_outputs(1764) <= inputs(227);
    layer0_outputs(1765) <= (inputs(133)) or (inputs(227));
    layer0_outputs(1766) <= (inputs(162)) and not (inputs(64));
    layer0_outputs(1767) <= (inputs(84)) xor (inputs(16));
    layer0_outputs(1768) <= '0';
    layer0_outputs(1769) <= not(inputs(151));
    layer0_outputs(1770) <= (inputs(139)) or (inputs(93));
    layer0_outputs(1771) <= '1';
    layer0_outputs(1772) <= inputs(201);
    layer0_outputs(1773) <= (inputs(108)) and not (inputs(185));
    layer0_outputs(1774) <= inputs(0);
    layer0_outputs(1775) <= '0';
    layer0_outputs(1776) <= not((inputs(232)) xor (inputs(169)));
    layer0_outputs(1777) <= (inputs(104)) or (inputs(101));
    layer0_outputs(1778) <= not(inputs(203));
    layer0_outputs(1779) <= (inputs(122)) or (inputs(44));
    layer0_outputs(1780) <= '1';
    layer0_outputs(1781) <= (inputs(216)) and (inputs(214));
    layer0_outputs(1782) <= not(inputs(120));
    layer0_outputs(1783) <= (inputs(244)) and not (inputs(133));
    layer0_outputs(1784) <= (inputs(151)) and not (inputs(156));
    layer0_outputs(1785) <= not(inputs(166));
    layer0_outputs(1786) <= (inputs(161)) xor (inputs(37));
    layer0_outputs(1787) <= inputs(87);
    layer0_outputs(1788) <= inputs(45);
    layer0_outputs(1789) <= not(inputs(34));
    layer0_outputs(1790) <= inputs(231);
    layer0_outputs(1791) <= (inputs(141)) or (inputs(158));
    layer0_outputs(1792) <= inputs(210);
    layer0_outputs(1793) <= '1';
    layer0_outputs(1794) <= '0';
    layer0_outputs(1795) <= not(inputs(152));
    layer0_outputs(1796) <= not((inputs(170)) and (inputs(244)));
    layer0_outputs(1797) <= (inputs(111)) or (inputs(173));
    layer0_outputs(1798) <= (inputs(231)) and not (inputs(107));
    layer0_outputs(1799) <= (inputs(116)) and not (inputs(194));
    layer0_outputs(1800) <= (inputs(186)) xor (inputs(221));
    layer0_outputs(1801) <= '1';
    layer0_outputs(1802) <= not(inputs(109));
    layer0_outputs(1803) <= inputs(184);
    layer0_outputs(1804) <= not(inputs(103)) or (inputs(180));
    layer0_outputs(1805) <= (inputs(113)) or (inputs(44));
    layer0_outputs(1806) <= (inputs(95)) or (inputs(192));
    layer0_outputs(1807) <= (inputs(138)) and not (inputs(47));
    layer0_outputs(1808) <= not((inputs(98)) xor (inputs(191)));
    layer0_outputs(1809) <= '0';
    layer0_outputs(1810) <= '0';
    layer0_outputs(1811) <= not((inputs(19)) or (inputs(253)));
    layer0_outputs(1812) <= (inputs(227)) and not (inputs(252));
    layer0_outputs(1813) <= not((inputs(8)) or (inputs(40)));
    layer0_outputs(1814) <= inputs(92);
    layer0_outputs(1815) <= '0';
    layer0_outputs(1816) <= not((inputs(151)) or (inputs(198)));
    layer0_outputs(1817) <= (inputs(212)) xor (inputs(44));
    layer0_outputs(1818) <= not((inputs(251)) or (inputs(170)));
    layer0_outputs(1819) <= '0';
    layer0_outputs(1820) <= (inputs(94)) xor (inputs(90));
    layer0_outputs(1821) <= not(inputs(242));
    layer0_outputs(1822) <= not(inputs(216));
    layer0_outputs(1823) <= (inputs(50)) and not (inputs(79));
    layer0_outputs(1824) <= not((inputs(196)) and (inputs(240)));
    layer0_outputs(1825) <= '0';
    layer0_outputs(1826) <= '0';
    layer0_outputs(1827) <= (inputs(58)) and not (inputs(190));
    layer0_outputs(1828) <= not((inputs(77)) or (inputs(65)));
    layer0_outputs(1829) <= not(inputs(163));
    layer0_outputs(1830) <= (inputs(112)) or (inputs(143));
    layer0_outputs(1831) <= '0';
    layer0_outputs(1832) <= (inputs(110)) or (inputs(243));
    layer0_outputs(1833) <= not(inputs(222)) or (inputs(154));
    layer0_outputs(1834) <= not(inputs(29));
    layer0_outputs(1835) <= inputs(84);
    layer0_outputs(1836) <= (inputs(95)) or (inputs(74));
    layer0_outputs(1837) <= (inputs(48)) and (inputs(41));
    layer0_outputs(1838) <= not((inputs(111)) or (inputs(227)));
    layer0_outputs(1839) <= (inputs(217)) and (inputs(223));
    layer0_outputs(1840) <= not(inputs(82)) or (inputs(24));
    layer0_outputs(1841) <= '0';
    layer0_outputs(1842) <= '1';
    layer0_outputs(1843) <= (inputs(46)) xor (inputs(120));
    layer0_outputs(1844) <= not(inputs(126));
    layer0_outputs(1845) <= not((inputs(115)) and (inputs(172)));
    layer0_outputs(1846) <= (inputs(182)) or (inputs(34));
    layer0_outputs(1847) <= '0';
    layer0_outputs(1848) <= '1';
    layer0_outputs(1849) <= '1';
    layer0_outputs(1850) <= (inputs(223)) or (inputs(53));
    layer0_outputs(1851) <= not(inputs(150));
    layer0_outputs(1852) <= inputs(35);
    layer0_outputs(1853) <= (inputs(228)) and not (inputs(59));
    layer0_outputs(1854) <= (inputs(128)) xor (inputs(180));
    layer0_outputs(1855) <= not(inputs(11)) or (inputs(177));
    layer0_outputs(1856) <= '1';
    layer0_outputs(1857) <= not(inputs(127));
    layer0_outputs(1858) <= '0';
    layer0_outputs(1859) <= not((inputs(43)) or (inputs(114)));
    layer0_outputs(1860) <= not(inputs(168));
    layer0_outputs(1861) <= '0';
    layer0_outputs(1862) <= inputs(145);
    layer0_outputs(1863) <= not((inputs(57)) or (inputs(140)));
    layer0_outputs(1864) <= inputs(144);
    layer0_outputs(1865) <= '0';
    layer0_outputs(1866) <= not(inputs(126)) or (inputs(247));
    layer0_outputs(1867) <= not(inputs(78));
    layer0_outputs(1868) <= not(inputs(180)) or (inputs(24));
    layer0_outputs(1869) <= not((inputs(163)) or (inputs(180)));
    layer0_outputs(1870) <= '0';
    layer0_outputs(1871) <= inputs(6);
    layer0_outputs(1872) <= '0';
    layer0_outputs(1873) <= '0';
    layer0_outputs(1874) <= '1';
    layer0_outputs(1875) <= inputs(239);
    layer0_outputs(1876) <= (inputs(1)) xor (inputs(3));
    layer0_outputs(1877) <= (inputs(233)) and not (inputs(193));
    layer0_outputs(1878) <= inputs(132);
    layer0_outputs(1879) <= '1';
    layer0_outputs(1880) <= (inputs(221)) and not (inputs(126));
    layer0_outputs(1881) <= not((inputs(230)) and (inputs(8)));
    layer0_outputs(1882) <= not(inputs(218)) or (inputs(151));
    layer0_outputs(1883) <= (inputs(177)) or (inputs(158));
    layer0_outputs(1884) <= not(inputs(157));
    layer0_outputs(1885) <= inputs(128);
    layer0_outputs(1886) <= not((inputs(159)) or (inputs(132)));
    layer0_outputs(1887) <= (inputs(165)) or (inputs(207));
    layer0_outputs(1888) <= not((inputs(213)) and (inputs(201)));
    layer0_outputs(1889) <= not(inputs(244)) or (inputs(237));
    layer0_outputs(1890) <= inputs(129);
    layer0_outputs(1891) <= (inputs(62)) or (inputs(140));
    layer0_outputs(1892) <= not(inputs(131)) or (inputs(32));
    layer0_outputs(1893) <= inputs(128);
    layer0_outputs(1894) <= inputs(246);
    layer0_outputs(1895) <= inputs(151);
    layer0_outputs(1896) <= (inputs(229)) or (inputs(9));
    layer0_outputs(1897) <= (inputs(208)) and not (inputs(216));
    layer0_outputs(1898) <= (inputs(180)) and (inputs(64));
    layer0_outputs(1899) <= (inputs(201)) and not (inputs(122));
    layer0_outputs(1900) <= (inputs(7)) or (inputs(187));
    layer0_outputs(1901) <= (inputs(161)) and not (inputs(31));
    layer0_outputs(1902) <= inputs(145);
    layer0_outputs(1903) <= not((inputs(232)) or (inputs(164)));
    layer0_outputs(1904) <= not(inputs(179));
    layer0_outputs(1905) <= not(inputs(80)) or (inputs(218));
    layer0_outputs(1906) <= '0';
    layer0_outputs(1907) <= inputs(129);
    layer0_outputs(1908) <= (inputs(244)) and not (inputs(238));
    layer0_outputs(1909) <= (inputs(108)) or (inputs(83));
    layer0_outputs(1910) <= inputs(93);
    layer0_outputs(1911) <= not(inputs(236)) or (inputs(191));
    layer0_outputs(1912) <= (inputs(54)) and not (inputs(103));
    layer0_outputs(1913) <= inputs(118);
    layer0_outputs(1914) <= (inputs(102)) and not (inputs(2));
    layer0_outputs(1915) <= not(inputs(182));
    layer0_outputs(1916) <= inputs(88);
    layer0_outputs(1917) <= (inputs(169)) and not (inputs(83));
    layer0_outputs(1918) <= '0';
    layer0_outputs(1919) <= not(inputs(179));
    layer0_outputs(1920) <= (inputs(162)) or (inputs(253));
    layer0_outputs(1921) <= (inputs(83)) or (inputs(138));
    layer0_outputs(1922) <= not((inputs(61)) and (inputs(224)));
    layer0_outputs(1923) <= not(inputs(46));
    layer0_outputs(1924) <= (inputs(197)) and not (inputs(232));
    layer0_outputs(1925) <= (inputs(88)) and not (inputs(202));
    layer0_outputs(1926) <= not((inputs(33)) or (inputs(174)));
    layer0_outputs(1927) <= not(inputs(33)) or (inputs(112));
    layer0_outputs(1928) <= not((inputs(63)) or (inputs(170)));
    layer0_outputs(1929) <= inputs(182);
    layer0_outputs(1930) <= not((inputs(63)) and (inputs(206)));
    layer0_outputs(1931) <= (inputs(234)) and not (inputs(25));
    layer0_outputs(1932) <= not(inputs(111)) or (inputs(155));
    layer0_outputs(1933) <= not(inputs(64)) or (inputs(46));
    layer0_outputs(1934) <= inputs(118);
    layer0_outputs(1935) <= not(inputs(57)) or (inputs(156));
    layer0_outputs(1936) <= not((inputs(247)) or (inputs(59)));
    layer0_outputs(1937) <= not(inputs(87));
    layer0_outputs(1938) <= not(inputs(33));
    layer0_outputs(1939) <= inputs(43);
    layer0_outputs(1940) <= inputs(156);
    layer0_outputs(1941) <= (inputs(48)) and not (inputs(106));
    layer0_outputs(1942) <= (inputs(166)) and (inputs(151));
    layer0_outputs(1943) <= (inputs(222)) and not (inputs(157));
    layer0_outputs(1944) <= not(inputs(22));
    layer0_outputs(1945) <= (inputs(120)) and not (inputs(111));
    layer0_outputs(1946) <= (inputs(77)) or (inputs(187));
    layer0_outputs(1947) <= (inputs(93)) or (inputs(95));
    layer0_outputs(1948) <= inputs(107);
    layer0_outputs(1949) <= '0';
    layer0_outputs(1950) <= not(inputs(25));
    layer0_outputs(1951) <= (inputs(47)) and (inputs(59));
    layer0_outputs(1952) <= inputs(147);
    layer0_outputs(1953) <= not((inputs(172)) or (inputs(221)));
    layer0_outputs(1954) <= not((inputs(228)) or (inputs(167)));
    layer0_outputs(1955) <= not((inputs(69)) or (inputs(138)));
    layer0_outputs(1956) <= (inputs(160)) or (inputs(25));
    layer0_outputs(1957) <= (inputs(100)) or (inputs(90));
    layer0_outputs(1958) <= not(inputs(207));
    layer0_outputs(1959) <= inputs(253);
    layer0_outputs(1960) <= (inputs(24)) and not (inputs(67));
    layer0_outputs(1961) <= (inputs(159)) or (inputs(193));
    layer0_outputs(1962) <= inputs(163);
    layer0_outputs(1963) <= (inputs(195)) and not (inputs(191));
    layer0_outputs(1964) <= not((inputs(152)) or (inputs(103)));
    layer0_outputs(1965) <= not((inputs(37)) and (inputs(36)));
    layer0_outputs(1966) <= (inputs(50)) and not (inputs(12));
    layer0_outputs(1967) <= not((inputs(1)) or (inputs(90)));
    layer0_outputs(1968) <= (inputs(6)) and not (inputs(240));
    layer0_outputs(1969) <= '1';
    layer0_outputs(1970) <= (inputs(241)) and (inputs(154));
    layer0_outputs(1971) <= not(inputs(61));
    layer0_outputs(1972) <= (inputs(85)) and not (inputs(62));
    layer0_outputs(1973) <= (inputs(139)) and not (inputs(37));
    layer0_outputs(1974) <= '1';
    layer0_outputs(1975) <= '1';
    layer0_outputs(1976) <= not(inputs(190)) or (inputs(81));
    layer0_outputs(1977) <= '1';
    layer0_outputs(1978) <= (inputs(57)) and not (inputs(251));
    layer0_outputs(1979) <= (inputs(219)) or (inputs(86));
    layer0_outputs(1980) <= '0';
    layer0_outputs(1981) <= not((inputs(60)) xor (inputs(171)));
    layer0_outputs(1982) <= inputs(157);
    layer0_outputs(1983) <= not(inputs(1));
    layer0_outputs(1984) <= not((inputs(27)) or (inputs(188)));
    layer0_outputs(1985) <= (inputs(106)) and not (inputs(34));
    layer0_outputs(1986) <= '1';
    layer0_outputs(1987) <= (inputs(134)) and not (inputs(190));
    layer0_outputs(1988) <= '1';
    layer0_outputs(1989) <= (inputs(28)) or (inputs(46));
    layer0_outputs(1990) <= inputs(206);
    layer0_outputs(1991) <= '1';
    layer0_outputs(1992) <= '1';
    layer0_outputs(1993) <= (inputs(56)) and (inputs(220));
    layer0_outputs(1994) <= (inputs(67)) or (inputs(84));
    layer0_outputs(1995) <= (inputs(191)) and not (inputs(20));
    layer0_outputs(1996) <= (inputs(155)) and not (inputs(188));
    layer0_outputs(1997) <= not((inputs(64)) and (inputs(203)));
    layer0_outputs(1998) <= not((inputs(115)) or (inputs(98)));
    layer0_outputs(1999) <= not(inputs(59)) or (inputs(245));
    layer0_outputs(2000) <= not((inputs(45)) and (inputs(58)));
    layer0_outputs(2001) <= '0';
    layer0_outputs(2002) <= inputs(10);
    layer0_outputs(2003) <= (inputs(231)) and not (inputs(64));
    layer0_outputs(2004) <= '1';
    layer0_outputs(2005) <= not(inputs(214));
    layer0_outputs(2006) <= not((inputs(218)) and (inputs(181)));
    layer0_outputs(2007) <= not(inputs(28)) or (inputs(114));
    layer0_outputs(2008) <= (inputs(139)) and not (inputs(243));
    layer0_outputs(2009) <= not(inputs(130)) or (inputs(56));
    layer0_outputs(2010) <= not(inputs(231)) or (inputs(252));
    layer0_outputs(2011) <= (inputs(169)) and not (inputs(95));
    layer0_outputs(2012) <= not(inputs(245));
    layer0_outputs(2013) <= inputs(235);
    layer0_outputs(2014) <= not(inputs(3)) or (inputs(247));
    layer0_outputs(2015) <= not(inputs(69));
    layer0_outputs(2016) <= (inputs(91)) and not (inputs(176));
    layer0_outputs(2017) <= not(inputs(107));
    layer0_outputs(2018) <= (inputs(127)) and (inputs(186));
    layer0_outputs(2019) <= inputs(0);
    layer0_outputs(2020) <= not(inputs(88));
    layer0_outputs(2021) <= not(inputs(136)) or (inputs(139));
    layer0_outputs(2022) <= not(inputs(145));
    layer0_outputs(2023) <= '0';
    layer0_outputs(2024) <= inputs(233);
    layer0_outputs(2025) <= '1';
    layer0_outputs(2026) <= not(inputs(167));
    layer0_outputs(2027) <= (inputs(119)) and not (inputs(123));
    layer0_outputs(2028) <= not(inputs(168)) or (inputs(60));
    layer0_outputs(2029) <= (inputs(18)) and (inputs(151));
    layer0_outputs(2030) <= not(inputs(8));
    layer0_outputs(2031) <= inputs(188);
    layer0_outputs(2032) <= not((inputs(200)) xor (inputs(170)));
    layer0_outputs(2033) <= (inputs(60)) xor (inputs(73));
    layer0_outputs(2034) <= not(inputs(59));
    layer0_outputs(2035) <= not(inputs(25));
    layer0_outputs(2036) <= '1';
    layer0_outputs(2037) <= not(inputs(133)) or (inputs(42));
    layer0_outputs(2038) <= not((inputs(98)) and (inputs(11)));
    layer0_outputs(2039) <= (inputs(244)) and (inputs(30));
    layer0_outputs(2040) <= (inputs(15)) and not (inputs(62));
    layer0_outputs(2041) <= '0';
    layer0_outputs(2042) <= not((inputs(235)) or (inputs(187)));
    layer0_outputs(2043) <= not(inputs(237));
    layer0_outputs(2044) <= (inputs(53)) or (inputs(2));
    layer0_outputs(2045) <= not(inputs(64)) or (inputs(244));
    layer0_outputs(2046) <= (inputs(73)) xor (inputs(67));
    layer0_outputs(2047) <= inputs(95);
    layer0_outputs(2048) <= not(inputs(253)) or (inputs(152));
    layer0_outputs(2049) <= '1';
    layer0_outputs(2050) <= (inputs(133)) and not (inputs(229));
    layer0_outputs(2051) <= inputs(55);
    layer0_outputs(2052) <= not((inputs(32)) or (inputs(142)));
    layer0_outputs(2053) <= not(inputs(101)) or (inputs(52));
    layer0_outputs(2054) <= inputs(77);
    layer0_outputs(2055) <= inputs(138);
    layer0_outputs(2056) <= '0';
    layer0_outputs(2057) <= (inputs(113)) and (inputs(42));
    layer0_outputs(2058) <= inputs(41);
    layer0_outputs(2059) <= inputs(76);
    layer0_outputs(2060) <= not((inputs(38)) and (inputs(208)));
    layer0_outputs(2061) <= not((inputs(206)) and (inputs(88)));
    layer0_outputs(2062) <= (inputs(188)) or (inputs(89));
    layer0_outputs(2063) <= (inputs(157)) and not (inputs(51));
    layer0_outputs(2064) <= not(inputs(61));
    layer0_outputs(2065) <= inputs(197);
    layer0_outputs(2066) <= (inputs(90)) xor (inputs(91));
    layer0_outputs(2067) <= (inputs(226)) and not (inputs(200));
    layer0_outputs(2068) <= '0';
    layer0_outputs(2069) <= not(inputs(240)) or (inputs(68));
    layer0_outputs(2070) <= (inputs(239)) and not (inputs(117));
    layer0_outputs(2071) <= (inputs(67)) and (inputs(23));
    layer0_outputs(2072) <= not((inputs(214)) or (inputs(205)));
    layer0_outputs(2073) <= inputs(64);
    layer0_outputs(2074) <= not((inputs(225)) or (inputs(250)));
    layer0_outputs(2075) <= '1';
    layer0_outputs(2076) <= '0';
    layer0_outputs(2077) <= not((inputs(102)) or (inputs(116)));
    layer0_outputs(2078) <= (inputs(175)) xor (inputs(176));
    layer0_outputs(2079) <= not((inputs(116)) or (inputs(223)));
    layer0_outputs(2080) <= inputs(147);
    layer0_outputs(2081) <= (inputs(193)) and not (inputs(184));
    layer0_outputs(2082) <= (inputs(122)) and not (inputs(116));
    layer0_outputs(2083) <= not(inputs(49)) or (inputs(73));
    layer0_outputs(2084) <= (inputs(208)) or (inputs(123));
    layer0_outputs(2085) <= (inputs(238)) and not (inputs(178));
    layer0_outputs(2086) <= (inputs(77)) and not (inputs(203));
    layer0_outputs(2087) <= '1';
    layer0_outputs(2088) <= (inputs(202)) or (inputs(137));
    layer0_outputs(2089) <= '1';
    layer0_outputs(2090) <= (inputs(216)) and (inputs(19));
    layer0_outputs(2091) <= (inputs(197)) and not (inputs(3));
    layer0_outputs(2092) <= '0';
    layer0_outputs(2093) <= (inputs(46)) or (inputs(61));
    layer0_outputs(2094) <= (inputs(156)) and not (inputs(34));
    layer0_outputs(2095) <= inputs(198);
    layer0_outputs(2096) <= not((inputs(234)) or (inputs(192)));
    layer0_outputs(2097) <= inputs(60);
    layer0_outputs(2098) <= not((inputs(80)) and (inputs(69)));
    layer0_outputs(2099) <= (inputs(78)) and not (inputs(186));
    layer0_outputs(2100) <= not((inputs(208)) or (inputs(171)));
    layer0_outputs(2101) <= '1';
    layer0_outputs(2102) <= '0';
    layer0_outputs(2103) <= '1';
    layer0_outputs(2104) <= '0';
    layer0_outputs(2105) <= not((inputs(84)) or (inputs(245)));
    layer0_outputs(2106) <= not(inputs(58));
    layer0_outputs(2107) <= inputs(174);
    layer0_outputs(2108) <= '1';
    layer0_outputs(2109) <= not((inputs(119)) xor (inputs(84)));
    layer0_outputs(2110) <= not((inputs(169)) and (inputs(236)));
    layer0_outputs(2111) <= (inputs(28)) and not (inputs(193));
    layer0_outputs(2112) <= (inputs(237)) or (inputs(48));
    layer0_outputs(2113) <= not(inputs(242)) or (inputs(203));
    layer0_outputs(2114) <= (inputs(25)) and not (inputs(205));
    layer0_outputs(2115) <= not(inputs(62));
    layer0_outputs(2116) <= inputs(41);
    layer0_outputs(2117) <= not(inputs(125)) or (inputs(233));
    layer0_outputs(2118) <= (inputs(36)) and (inputs(101));
    layer0_outputs(2119) <= '1';
    layer0_outputs(2120) <= (inputs(91)) or (inputs(36));
    layer0_outputs(2121) <= not((inputs(80)) and (inputs(142)));
    layer0_outputs(2122) <= (inputs(220)) or (inputs(143));
    layer0_outputs(2123) <= not((inputs(73)) xor (inputs(75)));
    layer0_outputs(2124) <= (inputs(24)) and not (inputs(180));
    layer0_outputs(2125) <= not((inputs(90)) or (inputs(162)));
    layer0_outputs(2126) <= inputs(240);
    layer0_outputs(2127) <= '0';
    layer0_outputs(2128) <= '1';
    layer0_outputs(2129) <= not((inputs(129)) or (inputs(72)));
    layer0_outputs(2130) <= '0';
    layer0_outputs(2131) <= '0';
    layer0_outputs(2132) <= (inputs(89)) and (inputs(2));
    layer0_outputs(2133) <= inputs(225);
    layer0_outputs(2134) <= not(inputs(117)) or (inputs(211));
    layer0_outputs(2135) <= inputs(192);
    layer0_outputs(2136) <= '0';
    layer0_outputs(2137) <= (inputs(47)) and not (inputs(170));
    layer0_outputs(2138) <= (inputs(81)) or (inputs(123));
    layer0_outputs(2139) <= inputs(78);
    layer0_outputs(2140) <= (inputs(86)) and not (inputs(45));
    layer0_outputs(2141) <= '0';
    layer0_outputs(2142) <= '0';
    layer0_outputs(2143) <= (inputs(61)) or (inputs(12));
    layer0_outputs(2144) <= '0';
    layer0_outputs(2145) <= inputs(193);
    layer0_outputs(2146) <= inputs(47);
    layer0_outputs(2147) <= (inputs(192)) and (inputs(44));
    layer0_outputs(2148) <= not((inputs(127)) xor (inputs(15)));
    layer0_outputs(2149) <= not((inputs(230)) xor (inputs(96)));
    layer0_outputs(2150) <= (inputs(220)) and not (inputs(20));
    layer0_outputs(2151) <= '0';
    layer0_outputs(2152) <= (inputs(232)) and (inputs(110));
    layer0_outputs(2153) <= (inputs(25)) and not (inputs(255));
    layer0_outputs(2154) <= (inputs(103)) or (inputs(253));
    layer0_outputs(2155) <= inputs(143);
    layer0_outputs(2156) <= (inputs(35)) or (inputs(65));
    layer0_outputs(2157) <= '0';
    layer0_outputs(2158) <= not((inputs(10)) and (inputs(21)));
    layer0_outputs(2159) <= (inputs(55)) and not (inputs(164));
    layer0_outputs(2160) <= not(inputs(233)) or (inputs(89));
    layer0_outputs(2161) <= (inputs(116)) and (inputs(101));
    layer0_outputs(2162) <= (inputs(139)) and not (inputs(181));
    layer0_outputs(2163) <= inputs(231);
    layer0_outputs(2164) <= (inputs(199)) and (inputs(91));
    layer0_outputs(2165) <= (inputs(164)) or (inputs(81));
    layer0_outputs(2166) <= (inputs(139)) xor (inputs(250));
    layer0_outputs(2167) <= (inputs(206)) and (inputs(184));
    layer0_outputs(2168) <= '0';
    layer0_outputs(2169) <= '1';
    layer0_outputs(2170) <= (inputs(84)) and (inputs(203));
    layer0_outputs(2171) <= '0';
    layer0_outputs(2172) <= not(inputs(250)) or (inputs(203));
    layer0_outputs(2173) <= not((inputs(225)) xor (inputs(255)));
    layer0_outputs(2174) <= not(inputs(47));
    layer0_outputs(2175) <= not(inputs(69)) or (inputs(234));
    layer0_outputs(2176) <= '0';
    layer0_outputs(2177) <= not((inputs(103)) and (inputs(251)));
    layer0_outputs(2178) <= not((inputs(87)) or (inputs(183)));
    layer0_outputs(2179) <= not((inputs(145)) and (inputs(83)));
    layer0_outputs(2180) <= not(inputs(108)) or (inputs(195));
    layer0_outputs(2181) <= inputs(255);
    layer0_outputs(2182) <= not((inputs(154)) or (inputs(190)));
    layer0_outputs(2183) <= (inputs(179)) or (inputs(166));
    layer0_outputs(2184) <= not((inputs(51)) and (inputs(72)));
    layer0_outputs(2185) <= not(inputs(189));
    layer0_outputs(2186) <= (inputs(100)) and not (inputs(63));
    layer0_outputs(2187) <= not(inputs(212)) or (inputs(167));
    layer0_outputs(2188) <= not(inputs(212));
    layer0_outputs(2189) <= '0';
    layer0_outputs(2190) <= '0';
    layer0_outputs(2191) <= not(inputs(163));
    layer0_outputs(2192) <= inputs(252);
    layer0_outputs(2193) <= '0';
    layer0_outputs(2194) <= not(inputs(64));
    layer0_outputs(2195) <= (inputs(197)) or (inputs(236));
    layer0_outputs(2196) <= '1';
    layer0_outputs(2197) <= (inputs(125)) and not (inputs(2));
    layer0_outputs(2198) <= not(inputs(126)) or (inputs(71));
    layer0_outputs(2199) <= not(inputs(199));
    layer0_outputs(2200) <= not(inputs(23));
    layer0_outputs(2201) <= (inputs(106)) xor (inputs(153));
    layer0_outputs(2202) <= inputs(99);
    layer0_outputs(2203) <= '1';
    layer0_outputs(2204) <= (inputs(116)) xor (inputs(112));
    layer0_outputs(2205) <= not((inputs(236)) or (inputs(164)));
    layer0_outputs(2206) <= not(inputs(157));
    layer0_outputs(2207) <= inputs(37);
    layer0_outputs(2208) <= inputs(230);
    layer0_outputs(2209) <= '0';
    layer0_outputs(2210) <= (inputs(53)) and not (inputs(198));
    layer0_outputs(2211) <= not((inputs(53)) and (inputs(19)));
    layer0_outputs(2212) <= (inputs(35)) and not (inputs(148));
    layer0_outputs(2213) <= not(inputs(92));
    layer0_outputs(2214) <= '0';
    layer0_outputs(2215) <= inputs(112);
    layer0_outputs(2216) <= (inputs(24)) and not (inputs(97));
    layer0_outputs(2217) <= inputs(87);
    layer0_outputs(2218) <= not((inputs(218)) or (inputs(204)));
    layer0_outputs(2219) <= (inputs(144)) or (inputs(33));
    layer0_outputs(2220) <= '1';
    layer0_outputs(2221) <= not((inputs(115)) or (inputs(156)));
    layer0_outputs(2222) <= (inputs(13)) or (inputs(105));
    layer0_outputs(2223) <= not(inputs(188));
    layer0_outputs(2224) <= '1';
    layer0_outputs(2225) <= '1';
    layer0_outputs(2226) <= inputs(209);
    layer0_outputs(2227) <= not(inputs(53));
    layer0_outputs(2228) <= not(inputs(107));
    layer0_outputs(2229) <= '1';
    layer0_outputs(2230) <= inputs(18);
    layer0_outputs(2231) <= (inputs(8)) and (inputs(117));
    layer0_outputs(2232) <= not(inputs(128)) or (inputs(28));
    layer0_outputs(2233) <= not(inputs(20));
    layer0_outputs(2234) <= not((inputs(95)) or (inputs(151)));
    layer0_outputs(2235) <= not(inputs(186)) or (inputs(16));
    layer0_outputs(2236) <= not(inputs(255)) or (inputs(133));
    layer0_outputs(2237) <= inputs(37);
    layer0_outputs(2238) <= '1';
    layer0_outputs(2239) <= not((inputs(107)) xor (inputs(113)));
    layer0_outputs(2240) <= not((inputs(189)) or (inputs(127)));
    layer0_outputs(2241) <= (inputs(207)) and (inputs(160));
    layer0_outputs(2242) <= not(inputs(204)) or (inputs(241));
    layer0_outputs(2243) <= not((inputs(145)) or (inputs(0)));
    layer0_outputs(2244) <= not(inputs(248)) or (inputs(137));
    layer0_outputs(2245) <= not(inputs(184));
    layer0_outputs(2246) <= '1';
    layer0_outputs(2247) <= inputs(89);
    layer0_outputs(2248) <= not(inputs(138)) or (inputs(207));
    layer0_outputs(2249) <= inputs(95);
    layer0_outputs(2250) <= not(inputs(71));
    layer0_outputs(2251) <= inputs(186);
    layer0_outputs(2252) <= (inputs(52)) or (inputs(33));
    layer0_outputs(2253) <= not(inputs(56)) or (inputs(2));
    layer0_outputs(2254) <= (inputs(13)) and not (inputs(185));
    layer0_outputs(2255) <= (inputs(3)) and not (inputs(220));
    layer0_outputs(2256) <= (inputs(87)) and not (inputs(141));
    layer0_outputs(2257) <= '1';
    layer0_outputs(2258) <= not((inputs(145)) or (inputs(159)));
    layer0_outputs(2259) <= inputs(184);
    layer0_outputs(2260) <= (inputs(249)) and not (inputs(14));
    layer0_outputs(2261) <= not(inputs(14));
    layer0_outputs(2262) <= '1';
    layer0_outputs(2263) <= not(inputs(97)) or (inputs(191));
    layer0_outputs(2264) <= inputs(39);
    layer0_outputs(2265) <= '1';
    layer0_outputs(2266) <= not(inputs(103));
    layer0_outputs(2267) <= not((inputs(210)) or (inputs(204)));
    layer0_outputs(2268) <= not((inputs(176)) xor (inputs(64)));
    layer0_outputs(2269) <= not((inputs(220)) or (inputs(2)));
    layer0_outputs(2270) <= (inputs(243)) or (inputs(33));
    layer0_outputs(2271) <= (inputs(91)) and not (inputs(224));
    layer0_outputs(2272) <= not((inputs(1)) or (inputs(6)));
    layer0_outputs(2273) <= '0';
    layer0_outputs(2274) <= not((inputs(162)) xor (inputs(160)));
    layer0_outputs(2275) <= not((inputs(222)) xor (inputs(252)));
    layer0_outputs(2276) <= '0';
    layer0_outputs(2277) <= (inputs(41)) and (inputs(247));
    layer0_outputs(2278) <= (inputs(117)) or (inputs(14));
    layer0_outputs(2279) <= not(inputs(125));
    layer0_outputs(2280) <= not(inputs(100));
    layer0_outputs(2281) <= not(inputs(87));
    layer0_outputs(2282) <= not(inputs(87)) or (inputs(108));
    layer0_outputs(2283) <= inputs(211);
    layer0_outputs(2284) <= '1';
    layer0_outputs(2285) <= not(inputs(219)) or (inputs(206));
    layer0_outputs(2286) <= inputs(134);
    layer0_outputs(2287) <= not((inputs(43)) or (inputs(46)));
    layer0_outputs(2288) <= not((inputs(123)) or (inputs(236)));
    layer0_outputs(2289) <= (inputs(141)) and not (inputs(61));
    layer0_outputs(2290) <= not(inputs(46));
    layer0_outputs(2291) <= inputs(115);
    layer0_outputs(2292) <= not(inputs(217));
    layer0_outputs(2293) <= not(inputs(230));
    layer0_outputs(2294) <= not((inputs(223)) or (inputs(166)));
    layer0_outputs(2295) <= not(inputs(52));
    layer0_outputs(2296) <= not((inputs(168)) and (inputs(29)));
    layer0_outputs(2297) <= not(inputs(41));
    layer0_outputs(2298) <= not((inputs(122)) and (inputs(210)));
    layer0_outputs(2299) <= (inputs(68)) or (inputs(54));
    layer0_outputs(2300) <= inputs(162);
    layer0_outputs(2301) <= not((inputs(196)) or (inputs(159)));
    layer0_outputs(2302) <= not((inputs(193)) or (inputs(219)));
    layer0_outputs(2303) <= (inputs(107)) or (inputs(112));
    layer0_outputs(2304) <= not((inputs(231)) or (inputs(15)));
    layer0_outputs(2305) <= '0';
    layer0_outputs(2306) <= not((inputs(92)) or (inputs(2)));
    layer0_outputs(2307) <= not(inputs(39)) or (inputs(100));
    layer0_outputs(2308) <= '1';
    layer0_outputs(2309) <= (inputs(95)) or (inputs(101));
    layer0_outputs(2310) <= (inputs(198)) and (inputs(119));
    layer0_outputs(2311) <= not(inputs(135));
    layer0_outputs(2312) <= not(inputs(86));
    layer0_outputs(2313) <= not(inputs(70)) or (inputs(63));
    layer0_outputs(2314) <= (inputs(179)) or (inputs(2));
    layer0_outputs(2315) <= inputs(242);
    layer0_outputs(2316) <= not((inputs(39)) xor (inputs(70)));
    layer0_outputs(2317) <= not((inputs(56)) and (inputs(64)));
    layer0_outputs(2318) <= not(inputs(242));
    layer0_outputs(2319) <= not((inputs(136)) or (inputs(190)));
    layer0_outputs(2320) <= not((inputs(204)) or (inputs(221)));
    layer0_outputs(2321) <= inputs(149);
    layer0_outputs(2322) <= not(inputs(85));
    layer0_outputs(2323) <= not(inputs(240)) or (inputs(59));
    layer0_outputs(2324) <= not((inputs(24)) and (inputs(31)));
    layer0_outputs(2325) <= not(inputs(192));
    layer0_outputs(2326) <= not(inputs(162));
    layer0_outputs(2327) <= (inputs(180)) or (inputs(238));
    layer0_outputs(2328) <= not(inputs(46));
    layer0_outputs(2329) <= not((inputs(86)) and (inputs(80)));
    layer0_outputs(2330) <= (inputs(253)) and (inputs(92));
    layer0_outputs(2331) <= (inputs(227)) and not (inputs(0));
    layer0_outputs(2332) <= '0';
    layer0_outputs(2333) <= not(inputs(230));
    layer0_outputs(2334) <= inputs(144);
    layer0_outputs(2335) <= '0';
    layer0_outputs(2336) <= not(inputs(102));
    layer0_outputs(2337) <= '0';
    layer0_outputs(2338) <= not(inputs(78));
    layer0_outputs(2339) <= (inputs(1)) and not (inputs(189));
    layer0_outputs(2340) <= '0';
    layer0_outputs(2341) <= inputs(102);
    layer0_outputs(2342) <= '0';
    layer0_outputs(2343) <= (inputs(135)) or (inputs(92));
    layer0_outputs(2344) <= not(inputs(143));
    layer0_outputs(2345) <= inputs(117);
    layer0_outputs(2346) <= (inputs(255)) and not (inputs(15));
    layer0_outputs(2347) <= not(inputs(33));
    layer0_outputs(2348) <= inputs(229);
    layer0_outputs(2349) <= '0';
    layer0_outputs(2350) <= '1';
    layer0_outputs(2351) <= (inputs(225)) or (inputs(0));
    layer0_outputs(2352) <= inputs(161);
    layer0_outputs(2353) <= '0';
    layer0_outputs(2354) <= inputs(128);
    layer0_outputs(2355) <= (inputs(18)) or (inputs(52));
    layer0_outputs(2356) <= (inputs(239)) and not (inputs(123));
    layer0_outputs(2357) <= (inputs(69)) xor (inputs(239));
    layer0_outputs(2358) <= (inputs(10)) and (inputs(207));
    layer0_outputs(2359) <= '1';
    layer0_outputs(2360) <= not(inputs(166));
    layer0_outputs(2361) <= (inputs(103)) and not (inputs(255));
    layer0_outputs(2362) <= inputs(96);
    layer0_outputs(2363) <= (inputs(27)) and not (inputs(149));
    layer0_outputs(2364) <= inputs(154);
    layer0_outputs(2365) <= not((inputs(194)) or (inputs(216)));
    layer0_outputs(2366) <= not(inputs(167)) or (inputs(51));
    layer0_outputs(2367) <= not(inputs(131));
    layer0_outputs(2368) <= (inputs(136)) and not (inputs(183));
    layer0_outputs(2369) <= (inputs(116)) and not (inputs(9));
    layer0_outputs(2370) <= not(inputs(106));
    layer0_outputs(2371) <= (inputs(168)) and not (inputs(183));
    layer0_outputs(2372) <= not(inputs(228)) or (inputs(34));
    layer0_outputs(2373) <= (inputs(83)) and not (inputs(18));
    layer0_outputs(2374) <= not((inputs(152)) or (inputs(98)));
    layer0_outputs(2375) <= (inputs(99)) and not (inputs(221));
    layer0_outputs(2376) <= not(inputs(114));
    layer0_outputs(2377) <= not(inputs(151)) or (inputs(50));
    layer0_outputs(2378) <= not(inputs(192)) or (inputs(203));
    layer0_outputs(2379) <= '1';
    layer0_outputs(2380) <= '1';
    layer0_outputs(2381) <= not(inputs(198)) or (inputs(1));
    layer0_outputs(2382) <= not((inputs(163)) or (inputs(66)));
    layer0_outputs(2383) <= not(inputs(126));
    layer0_outputs(2384) <= (inputs(179)) or (inputs(38));
    layer0_outputs(2385) <= inputs(101);
    layer0_outputs(2386) <= not(inputs(65)) or (inputs(127));
    layer0_outputs(2387) <= (inputs(70)) and not (inputs(157));
    layer0_outputs(2388) <= '0';
    layer0_outputs(2389) <= inputs(127);
    layer0_outputs(2390) <= (inputs(108)) and not (inputs(62));
    layer0_outputs(2391) <= (inputs(0)) and not (inputs(29));
    layer0_outputs(2392) <= not((inputs(165)) or (inputs(161)));
    layer0_outputs(2393) <= not(inputs(41));
    layer0_outputs(2394) <= (inputs(85)) and not (inputs(191));
    layer0_outputs(2395) <= not(inputs(240)) or (inputs(2));
    layer0_outputs(2396) <= inputs(124);
    layer0_outputs(2397) <= not((inputs(82)) or (inputs(179)));
    layer0_outputs(2398) <= (inputs(34)) and (inputs(60));
    layer0_outputs(2399) <= (inputs(176)) and not (inputs(96));
    layer0_outputs(2400) <= not(inputs(160));
    layer0_outputs(2401) <= not(inputs(138)) or (inputs(118));
    layer0_outputs(2402) <= '1';
    layer0_outputs(2403) <= not((inputs(167)) and (inputs(221)));
    layer0_outputs(2404) <= inputs(111);
    layer0_outputs(2405) <= inputs(132);
    layer0_outputs(2406) <= '0';
    layer0_outputs(2407) <= (inputs(74)) and not (inputs(227));
    layer0_outputs(2408) <= not(inputs(182));
    layer0_outputs(2409) <= not(inputs(31)) or (inputs(104));
    layer0_outputs(2410) <= '1';
    layer0_outputs(2411) <= '0';
    layer0_outputs(2412) <= (inputs(32)) and not (inputs(151));
    layer0_outputs(2413) <= not(inputs(190));
    layer0_outputs(2414) <= (inputs(2)) or (inputs(253));
    layer0_outputs(2415) <= not(inputs(159));
    layer0_outputs(2416) <= not(inputs(173));
    layer0_outputs(2417) <= (inputs(177)) xor (inputs(15));
    layer0_outputs(2418) <= not(inputs(151));
    layer0_outputs(2419) <= (inputs(92)) and not (inputs(152));
    layer0_outputs(2420) <= (inputs(69)) or (inputs(160));
    layer0_outputs(2421) <= inputs(129);
    layer0_outputs(2422) <= (inputs(24)) and not (inputs(64));
    layer0_outputs(2423) <= inputs(218);
    layer0_outputs(2424) <= not(inputs(203)) or (inputs(129));
    layer0_outputs(2425) <= (inputs(44)) and not (inputs(195));
    layer0_outputs(2426) <= inputs(148);
    layer0_outputs(2427) <= not((inputs(82)) xor (inputs(186)));
    layer0_outputs(2428) <= (inputs(11)) and (inputs(219));
    layer0_outputs(2429) <= not(inputs(76)) or (inputs(112));
    layer0_outputs(2430) <= (inputs(134)) and not (inputs(109));
    layer0_outputs(2431) <= inputs(98);
    layer0_outputs(2432) <= not(inputs(113));
    layer0_outputs(2433) <= inputs(205);
    layer0_outputs(2434) <= (inputs(115)) and (inputs(121));
    layer0_outputs(2435) <= inputs(67);
    layer0_outputs(2436) <= '1';
    layer0_outputs(2437) <= inputs(27);
    layer0_outputs(2438) <= (inputs(17)) and not (inputs(140));
    layer0_outputs(2439) <= (inputs(13)) or (inputs(207));
    layer0_outputs(2440) <= (inputs(209)) or (inputs(224));
    layer0_outputs(2441) <= not(inputs(165));
    layer0_outputs(2442) <= inputs(165);
    layer0_outputs(2443) <= (inputs(193)) or (inputs(251));
    layer0_outputs(2444) <= (inputs(194)) and not (inputs(48));
    layer0_outputs(2445) <= (inputs(81)) and (inputs(28));
    layer0_outputs(2446) <= '1';
    layer0_outputs(2447) <= (inputs(84)) and not (inputs(205));
    layer0_outputs(2448) <= (inputs(125)) and not (inputs(13));
    layer0_outputs(2449) <= '1';
    layer0_outputs(2450) <= (inputs(110)) and (inputs(31));
    layer0_outputs(2451) <= not(inputs(105));
    layer0_outputs(2452) <= not(inputs(128));
    layer0_outputs(2453) <= '1';
    layer0_outputs(2454) <= '1';
    layer0_outputs(2455) <= inputs(134);
    layer0_outputs(2456) <= not((inputs(110)) and (inputs(54)));
    layer0_outputs(2457) <= inputs(255);
    layer0_outputs(2458) <= '1';
    layer0_outputs(2459) <= (inputs(253)) and (inputs(76));
    layer0_outputs(2460) <= not(inputs(139));
    layer0_outputs(2461) <= '0';
    layer0_outputs(2462) <= not((inputs(146)) or (inputs(201)));
    layer0_outputs(2463) <= (inputs(199)) and (inputs(242));
    layer0_outputs(2464) <= inputs(170);
    layer0_outputs(2465) <= not(inputs(45));
    layer0_outputs(2466) <= (inputs(138)) and not (inputs(228));
    layer0_outputs(2467) <= not(inputs(206)) or (inputs(49));
    layer0_outputs(2468) <= '1';
    layer0_outputs(2469) <= not((inputs(178)) or (inputs(246)));
    layer0_outputs(2470) <= not((inputs(42)) or (inputs(195)));
    layer0_outputs(2471) <= '1';
    layer0_outputs(2472) <= not((inputs(191)) or (inputs(225)));
    layer0_outputs(2473) <= not((inputs(225)) or (inputs(159)));
    layer0_outputs(2474) <= not((inputs(87)) and (inputs(17)));
    layer0_outputs(2475) <= (inputs(20)) or (inputs(18));
    layer0_outputs(2476) <= (inputs(160)) or (inputs(220));
    layer0_outputs(2477) <= not(inputs(110));
    layer0_outputs(2478) <= (inputs(140)) or (inputs(233));
    layer0_outputs(2479) <= not(inputs(2));
    layer0_outputs(2480) <= not(inputs(219)) or (inputs(39));
    layer0_outputs(2481) <= (inputs(12)) and not (inputs(245));
    layer0_outputs(2482) <= not(inputs(157));
    layer0_outputs(2483) <= not((inputs(213)) xor (inputs(209)));
    layer0_outputs(2484) <= not(inputs(168));
    layer0_outputs(2485) <= not((inputs(193)) or (inputs(54)));
    layer0_outputs(2486) <= (inputs(6)) or (inputs(213));
    layer0_outputs(2487) <= '0';
    layer0_outputs(2488) <= (inputs(157)) and not (inputs(179));
    layer0_outputs(2489) <= (inputs(151)) and not (inputs(90));
    layer0_outputs(2490) <= (inputs(130)) or (inputs(160));
    layer0_outputs(2491) <= (inputs(175)) or (inputs(146));
    layer0_outputs(2492) <= not(inputs(230));
    layer0_outputs(2493) <= '0';
    layer0_outputs(2494) <= '0';
    layer0_outputs(2495) <= inputs(39);
    layer0_outputs(2496) <= (inputs(127)) and not (inputs(8));
    layer0_outputs(2497) <= '0';
    layer0_outputs(2498) <= (inputs(175)) and not (inputs(142));
    layer0_outputs(2499) <= '1';
    layer0_outputs(2500) <= inputs(243);
    layer0_outputs(2501) <= '1';
    layer0_outputs(2502) <= (inputs(203)) and not (inputs(171));
    layer0_outputs(2503) <= not(inputs(215)) or (inputs(59));
    layer0_outputs(2504) <= not((inputs(197)) and (inputs(96)));
    layer0_outputs(2505) <= (inputs(161)) and (inputs(70));
    layer0_outputs(2506) <= '1';
    layer0_outputs(2507) <= '1';
    layer0_outputs(2508) <= '1';
    layer0_outputs(2509) <= inputs(105);
    layer0_outputs(2510) <= not(inputs(234));
    layer0_outputs(2511) <= (inputs(208)) or (inputs(157));
    layer0_outputs(2512) <= inputs(33);
    layer0_outputs(2513) <= not(inputs(253));
    layer0_outputs(2514) <= not(inputs(96)) or (inputs(27));
    layer0_outputs(2515) <= inputs(167);
    layer0_outputs(2516) <= not(inputs(192));
    layer0_outputs(2517) <= (inputs(157)) and not (inputs(133));
    layer0_outputs(2518) <= not((inputs(236)) xor (inputs(159)));
    layer0_outputs(2519) <= inputs(156);
    layer0_outputs(2520) <= not((inputs(159)) xor (inputs(243)));
    layer0_outputs(2521) <= not(inputs(55));
    layer0_outputs(2522) <= (inputs(254)) or (inputs(105));
    layer0_outputs(2523) <= not((inputs(71)) or (inputs(159)));
    layer0_outputs(2524) <= '0';
    layer0_outputs(2525) <= not(inputs(82)) or (inputs(64));
    layer0_outputs(2526) <= '0';
    layer0_outputs(2527) <= (inputs(70)) and not (inputs(49));
    layer0_outputs(2528) <= '1';
    layer0_outputs(2529) <= not(inputs(231)) or (inputs(234));
    layer0_outputs(2530) <= inputs(214);
    layer0_outputs(2531) <= not(inputs(164)) or (inputs(25));
    layer0_outputs(2532) <= inputs(165);
    layer0_outputs(2533) <= not(inputs(98)) or (inputs(162));
    layer0_outputs(2534) <= not(inputs(90));
    layer0_outputs(2535) <= '1';
    layer0_outputs(2536) <= not((inputs(218)) or (inputs(138)));
    layer0_outputs(2537) <= (inputs(139)) and not (inputs(146));
    layer0_outputs(2538) <= '0';
    layer0_outputs(2539) <= not(inputs(26)) or (inputs(183));
    layer0_outputs(2540) <= (inputs(94)) and (inputs(148));
    layer0_outputs(2541) <= not(inputs(57));
    layer0_outputs(2542) <= not(inputs(230));
    layer0_outputs(2543) <= (inputs(187)) or (inputs(190));
    layer0_outputs(2544) <= not(inputs(141));
    layer0_outputs(2545) <= (inputs(76)) or (inputs(162));
    layer0_outputs(2546) <= not(inputs(183)) or (inputs(62));
    layer0_outputs(2547) <= not(inputs(128));
    layer0_outputs(2548) <= '0';
    layer0_outputs(2549) <= not(inputs(165));
    layer0_outputs(2550) <= not(inputs(9));
    layer0_outputs(2551) <= not((inputs(82)) or (inputs(81)));
    layer0_outputs(2552) <= not(inputs(221)) or (inputs(62));
    layer0_outputs(2553) <= (inputs(36)) and not (inputs(250));
    layer0_outputs(2554) <= '0';
    layer0_outputs(2555) <= not(inputs(176));
    layer0_outputs(2556) <= not((inputs(252)) and (inputs(141)));
    layer0_outputs(2557) <= (inputs(164)) and not (inputs(138));
    layer0_outputs(2558) <= (inputs(199)) and not (inputs(159));
    layer0_outputs(2559) <= not(inputs(64));
    layer0_outputs(2560) <= (inputs(121)) or (inputs(230));
    layer0_outputs(2561) <= (inputs(30)) and not (inputs(191));
    layer0_outputs(2562) <= not(inputs(71)) or (inputs(251));
    layer0_outputs(2563) <= (inputs(23)) xor (inputs(114));
    layer0_outputs(2564) <= not(inputs(241));
    layer0_outputs(2565) <= not((inputs(100)) xor (inputs(163)));
    layer0_outputs(2566) <= '1';
    layer0_outputs(2567) <= '0';
    layer0_outputs(2568) <= not(inputs(7));
    layer0_outputs(2569) <= not((inputs(119)) or (inputs(48)));
    layer0_outputs(2570) <= not(inputs(37));
    layer0_outputs(2571) <= not(inputs(123));
    layer0_outputs(2572) <= '0';
    layer0_outputs(2573) <= inputs(221);
    layer0_outputs(2574) <= not((inputs(245)) and (inputs(192)));
    layer0_outputs(2575) <= inputs(150);
    layer0_outputs(2576) <= (inputs(112)) and not (inputs(7));
    layer0_outputs(2577) <= '1';
    layer0_outputs(2578) <= inputs(114);
    layer0_outputs(2579) <= not(inputs(252));
    layer0_outputs(2580) <= inputs(195);
    layer0_outputs(2581) <= (inputs(227)) and not (inputs(124));
    layer0_outputs(2582) <= (inputs(105)) or (inputs(197));
    layer0_outputs(2583) <= not(inputs(211)) or (inputs(48));
    layer0_outputs(2584) <= inputs(252);
    layer0_outputs(2585) <= not(inputs(15));
    layer0_outputs(2586) <= not(inputs(56)) or (inputs(29));
    layer0_outputs(2587) <= not((inputs(242)) and (inputs(241)));
    layer0_outputs(2588) <= inputs(86);
    layer0_outputs(2589) <= (inputs(212)) and (inputs(167));
    layer0_outputs(2590) <= '0';
    layer0_outputs(2591) <= '1';
    layer0_outputs(2592) <= not(inputs(252)) or (inputs(191));
    layer0_outputs(2593) <= not((inputs(146)) or (inputs(151)));
    layer0_outputs(2594) <= (inputs(157)) and not (inputs(59));
    layer0_outputs(2595) <= inputs(109);
    layer0_outputs(2596) <= '1';
    layer0_outputs(2597) <= not((inputs(141)) and (inputs(42)));
    layer0_outputs(2598) <= (inputs(89)) and not (inputs(31));
    layer0_outputs(2599) <= '1';
    layer0_outputs(2600) <= not(inputs(32));
    layer0_outputs(2601) <= inputs(117);
    layer0_outputs(2602) <= (inputs(64)) xor (inputs(131));
    layer0_outputs(2603) <= not(inputs(132));
    layer0_outputs(2604) <= inputs(33);
    layer0_outputs(2605) <= '1';
    layer0_outputs(2606) <= not(inputs(197));
    layer0_outputs(2607) <= not(inputs(79));
    layer0_outputs(2608) <= inputs(206);
    layer0_outputs(2609) <= (inputs(119)) and not (inputs(205));
    layer0_outputs(2610) <= inputs(105);
    layer0_outputs(2611) <= inputs(161);
    layer0_outputs(2612) <= not(inputs(64)) or (inputs(74));
    layer0_outputs(2613) <= (inputs(194)) and (inputs(229));
    layer0_outputs(2614) <= (inputs(107)) and not (inputs(195));
    layer0_outputs(2615) <= not((inputs(43)) or (inputs(125)));
    layer0_outputs(2616) <= not(inputs(63));
    layer0_outputs(2617) <= (inputs(94)) and (inputs(58));
    layer0_outputs(2618) <= not((inputs(76)) or (inputs(12)));
    layer0_outputs(2619) <= (inputs(250)) and not (inputs(221));
    layer0_outputs(2620) <= inputs(145);
    layer0_outputs(2621) <= not(inputs(210)) or (inputs(237));
    layer0_outputs(2622) <= (inputs(222)) and not (inputs(81));
    layer0_outputs(2623) <= inputs(231);
    layer0_outputs(2624) <= '1';
    layer0_outputs(2625) <= '0';
    layer0_outputs(2626) <= (inputs(33)) and not (inputs(185));
    layer0_outputs(2627) <= (inputs(188)) and not (inputs(148));
    layer0_outputs(2628) <= not(inputs(135)) or (inputs(101));
    layer0_outputs(2629) <= inputs(163);
    layer0_outputs(2630) <= not((inputs(91)) xor (inputs(15)));
    layer0_outputs(2631) <= '0';
    layer0_outputs(2632) <= inputs(64);
    layer0_outputs(2633) <= '0';
    layer0_outputs(2634) <= '0';
    layer0_outputs(2635) <= not(inputs(227)) or (inputs(88));
    layer0_outputs(2636) <= not((inputs(19)) xor (inputs(50)));
    layer0_outputs(2637) <= not(inputs(44)) or (inputs(16));
    layer0_outputs(2638) <= not(inputs(226));
    layer0_outputs(2639) <= not(inputs(235));
    layer0_outputs(2640) <= inputs(26);
    layer0_outputs(2641) <= inputs(104);
    layer0_outputs(2642) <= not((inputs(157)) or (inputs(100)));
    layer0_outputs(2643) <= inputs(180);
    layer0_outputs(2644) <= not(inputs(157));
    layer0_outputs(2645) <= not(inputs(205));
    layer0_outputs(2646) <= '1';
    layer0_outputs(2647) <= not(inputs(79)) or (inputs(4));
    layer0_outputs(2648) <= '0';
    layer0_outputs(2649) <= not(inputs(8)) or (inputs(184));
    layer0_outputs(2650) <= not((inputs(135)) and (inputs(188)));
    layer0_outputs(2651) <= not(inputs(227)) or (inputs(40));
    layer0_outputs(2652) <= not((inputs(206)) xor (inputs(159)));
    layer0_outputs(2653) <= (inputs(251)) and (inputs(97));
    layer0_outputs(2654) <= not(inputs(178));
    layer0_outputs(2655) <= (inputs(133)) xor (inputs(114));
    layer0_outputs(2656) <= (inputs(120)) or (inputs(46));
    layer0_outputs(2657) <= inputs(158);
    layer0_outputs(2658) <= not(inputs(100)) or (inputs(217));
    layer0_outputs(2659) <= (inputs(140)) and (inputs(221));
    layer0_outputs(2660) <= not(inputs(90)) or (inputs(144));
    layer0_outputs(2661) <= not((inputs(216)) xor (inputs(176)));
    layer0_outputs(2662) <= not(inputs(1)) or (inputs(176));
    layer0_outputs(2663) <= '0';
    layer0_outputs(2664) <= not(inputs(96));
    layer0_outputs(2665) <= inputs(38);
    layer0_outputs(2666) <= not((inputs(68)) and (inputs(170)));
    layer0_outputs(2667) <= not((inputs(7)) or (inputs(123)));
    layer0_outputs(2668) <= '1';
    layer0_outputs(2669) <= (inputs(255)) xor (inputs(115));
    layer0_outputs(2670) <= not((inputs(235)) or (inputs(30)));
    layer0_outputs(2671) <= '0';
    layer0_outputs(2672) <= not(inputs(8));
    layer0_outputs(2673) <= (inputs(141)) and not (inputs(249));
    layer0_outputs(2674) <= not((inputs(217)) or (inputs(210)));
    layer0_outputs(2675) <= not((inputs(148)) or (inputs(98)));
    layer0_outputs(2676) <= not(inputs(180)) or (inputs(89));
    layer0_outputs(2677) <= (inputs(148)) xor (inputs(117));
    layer0_outputs(2678) <= (inputs(19)) xor (inputs(18));
    layer0_outputs(2679) <= inputs(124);
    layer0_outputs(2680) <= (inputs(158)) and (inputs(201));
    layer0_outputs(2681) <= not(inputs(100));
    layer0_outputs(2682) <= not(inputs(74)) or (inputs(0));
    layer0_outputs(2683) <= (inputs(125)) and not (inputs(48));
    layer0_outputs(2684) <= '1';
    layer0_outputs(2685) <= (inputs(22)) xor (inputs(231));
    layer0_outputs(2686) <= (inputs(67)) and not (inputs(93));
    layer0_outputs(2687) <= '1';
    layer0_outputs(2688) <= not(inputs(65));
    layer0_outputs(2689) <= not(inputs(43));
    layer0_outputs(2690) <= (inputs(30)) and not (inputs(178));
    layer0_outputs(2691) <= not(inputs(67));
    layer0_outputs(2692) <= inputs(31);
    layer0_outputs(2693) <= not((inputs(128)) or (inputs(134)));
    layer0_outputs(2694) <= (inputs(208)) or (inputs(108));
    layer0_outputs(2695) <= (inputs(37)) and not (inputs(114));
    layer0_outputs(2696) <= inputs(168);
    layer0_outputs(2697) <= not(inputs(71));
    layer0_outputs(2698) <= (inputs(229)) or (inputs(162));
    layer0_outputs(2699) <= not(inputs(124));
    layer0_outputs(2700) <= inputs(26);
    layer0_outputs(2701) <= '1';
    layer0_outputs(2702) <= inputs(86);
    layer0_outputs(2703) <= (inputs(123)) or (inputs(5));
    layer0_outputs(2704) <= inputs(57);
    layer0_outputs(2705) <= inputs(120);
    layer0_outputs(2706) <= (inputs(252)) or (inputs(9));
    layer0_outputs(2707) <= (inputs(209)) or (inputs(172));
    layer0_outputs(2708) <= '0';
    layer0_outputs(2709) <= inputs(93);
    layer0_outputs(2710) <= not(inputs(240)) or (inputs(19));
    layer0_outputs(2711) <= (inputs(73)) or (inputs(89));
    layer0_outputs(2712) <= '0';
    layer0_outputs(2713) <= (inputs(58)) or (inputs(232));
    layer0_outputs(2714) <= not(inputs(225));
    layer0_outputs(2715) <= not(inputs(188));
    layer0_outputs(2716) <= '0';
    layer0_outputs(2717) <= inputs(195);
    layer0_outputs(2718) <= (inputs(20)) and not (inputs(14));
    layer0_outputs(2719) <= (inputs(217)) or (inputs(173));
    layer0_outputs(2720) <= not(inputs(0));
    layer0_outputs(2721) <= (inputs(99)) or (inputs(32));
    layer0_outputs(2722) <= '1';
    layer0_outputs(2723) <= not(inputs(4));
    layer0_outputs(2724) <= not((inputs(28)) or (inputs(5)));
    layer0_outputs(2725) <= '0';
    layer0_outputs(2726) <= not(inputs(242));
    layer0_outputs(2727) <= not(inputs(120));
    layer0_outputs(2728) <= not((inputs(250)) and (inputs(163)));
    layer0_outputs(2729) <= not(inputs(104)) or (inputs(168));
    layer0_outputs(2730) <= not(inputs(25));
    layer0_outputs(2731) <= not(inputs(155)) or (inputs(214));
    layer0_outputs(2732) <= (inputs(27)) and (inputs(11));
    layer0_outputs(2733) <= (inputs(227)) and not (inputs(95));
    layer0_outputs(2734) <= not(inputs(124));
    layer0_outputs(2735) <= (inputs(170)) and not (inputs(71));
    layer0_outputs(2736) <= '1';
    layer0_outputs(2737) <= (inputs(66)) or (inputs(217));
    layer0_outputs(2738) <= '1';
    layer0_outputs(2739) <= not(inputs(63));
    layer0_outputs(2740) <= not(inputs(24));
    layer0_outputs(2741) <= not(inputs(227));
    layer0_outputs(2742) <= not(inputs(131)) or (inputs(30));
    layer0_outputs(2743) <= '0';
    layer0_outputs(2744) <= not((inputs(111)) xor (inputs(103)));
    layer0_outputs(2745) <= inputs(160);
    layer0_outputs(2746) <= not(inputs(42)) or (inputs(172));
    layer0_outputs(2747) <= (inputs(189)) and not (inputs(75));
    layer0_outputs(2748) <= '0';
    layer0_outputs(2749) <= not(inputs(180));
    layer0_outputs(2750) <= not((inputs(41)) and (inputs(255)));
    layer0_outputs(2751) <= inputs(199);
    layer0_outputs(2752) <= not(inputs(194));
    layer0_outputs(2753) <= not(inputs(135)) or (inputs(189));
    layer0_outputs(2754) <= '1';
    layer0_outputs(2755) <= not(inputs(78)) or (inputs(220));
    layer0_outputs(2756) <= not(inputs(57)) or (inputs(34));
    layer0_outputs(2757) <= not(inputs(113));
    layer0_outputs(2758) <= not(inputs(189));
    layer0_outputs(2759) <= inputs(196);
    layer0_outputs(2760) <= (inputs(158)) or (inputs(96));
    layer0_outputs(2761) <= '1';
    layer0_outputs(2762) <= not(inputs(224)) or (inputs(93));
    layer0_outputs(2763) <= (inputs(70)) and not (inputs(79));
    layer0_outputs(2764) <= (inputs(54)) and not (inputs(123));
    layer0_outputs(2765) <= inputs(189);
    layer0_outputs(2766) <= not(inputs(254));
    layer0_outputs(2767) <= '1';
    layer0_outputs(2768) <= '1';
    layer0_outputs(2769) <= (inputs(187)) and (inputs(166));
    layer0_outputs(2770) <= not(inputs(89));
    layer0_outputs(2771) <= inputs(160);
    layer0_outputs(2772) <= '0';
    layer0_outputs(2773) <= not(inputs(100));
    layer0_outputs(2774) <= (inputs(149)) and not (inputs(3));
    layer0_outputs(2775) <= inputs(92);
    layer0_outputs(2776) <= '0';
    layer0_outputs(2777) <= not(inputs(232));
    layer0_outputs(2778) <= (inputs(69)) and not (inputs(137));
    layer0_outputs(2779) <= inputs(145);
    layer0_outputs(2780) <= (inputs(65)) or (inputs(170));
    layer0_outputs(2781) <= inputs(108);
    layer0_outputs(2782) <= inputs(108);
    layer0_outputs(2783) <= (inputs(189)) and not (inputs(91));
    layer0_outputs(2784) <= (inputs(142)) xor (inputs(105));
    layer0_outputs(2785) <= (inputs(176)) and not (inputs(110));
    layer0_outputs(2786) <= not((inputs(148)) or (inputs(212)));
    layer0_outputs(2787) <= '1';
    layer0_outputs(2788) <= not(inputs(93)) or (inputs(2));
    layer0_outputs(2789) <= inputs(65);
    layer0_outputs(2790) <= not(inputs(33)) or (inputs(112));
    layer0_outputs(2791) <= not((inputs(217)) or (inputs(189)));
    layer0_outputs(2792) <= not((inputs(68)) and (inputs(155)));
    layer0_outputs(2793) <= (inputs(14)) or (inputs(210));
    layer0_outputs(2794) <= inputs(143);
    layer0_outputs(2795) <= (inputs(143)) and (inputs(196));
    layer0_outputs(2796) <= (inputs(107)) and not (inputs(156));
    layer0_outputs(2797) <= '1';
    layer0_outputs(2798) <= not((inputs(87)) and (inputs(203)));
    layer0_outputs(2799) <= inputs(222);
    layer0_outputs(2800) <= not((inputs(222)) and (inputs(174)));
    layer0_outputs(2801) <= not((inputs(48)) or (inputs(59)));
    layer0_outputs(2802) <= not(inputs(25));
    layer0_outputs(2803) <= not(inputs(80)) or (inputs(227));
    layer0_outputs(2804) <= '0';
    layer0_outputs(2805) <= not((inputs(5)) or (inputs(90)));
    layer0_outputs(2806) <= inputs(6);
    layer0_outputs(2807) <= (inputs(164)) and not (inputs(208));
    layer0_outputs(2808) <= (inputs(189)) or (inputs(18));
    layer0_outputs(2809) <= (inputs(229)) and not (inputs(0));
    layer0_outputs(2810) <= (inputs(234)) or (inputs(145));
    layer0_outputs(2811) <= (inputs(133)) and (inputs(14));
    layer0_outputs(2812) <= (inputs(211)) or (inputs(229));
    layer0_outputs(2813) <= inputs(229);
    layer0_outputs(2814) <= '0';
    layer0_outputs(2815) <= (inputs(82)) xor (inputs(123));
    layer0_outputs(2816) <= inputs(67);
    layer0_outputs(2817) <= not(inputs(91)) or (inputs(38));
    layer0_outputs(2818) <= (inputs(176)) and not (inputs(236));
    layer0_outputs(2819) <= inputs(101);
    layer0_outputs(2820) <= '0';
    layer0_outputs(2821) <= not(inputs(232));
    layer0_outputs(2822) <= not(inputs(64));
    layer0_outputs(2823) <= inputs(95);
    layer0_outputs(2824) <= not((inputs(237)) or (inputs(51)));
    layer0_outputs(2825) <= not((inputs(116)) or (inputs(115)));
    layer0_outputs(2826) <= (inputs(255)) or (inputs(63));
    layer0_outputs(2827) <= inputs(127);
    layer0_outputs(2828) <= (inputs(226)) and not (inputs(211));
    layer0_outputs(2829) <= (inputs(199)) xor (inputs(247));
    layer0_outputs(2830) <= (inputs(195)) and not (inputs(21));
    layer0_outputs(2831) <= (inputs(169)) and not (inputs(161));
    layer0_outputs(2832) <= not((inputs(167)) or (inputs(92)));
    layer0_outputs(2833) <= not(inputs(180)) or (inputs(172));
    layer0_outputs(2834) <= (inputs(99)) and (inputs(117));
    layer0_outputs(2835) <= (inputs(166)) or (inputs(252));
    layer0_outputs(2836) <= not(inputs(151));
    layer0_outputs(2837) <= (inputs(23)) xor (inputs(207));
    layer0_outputs(2838) <= not((inputs(148)) or (inputs(185)));
    layer0_outputs(2839) <= (inputs(91)) xor (inputs(48));
    layer0_outputs(2840) <= not((inputs(212)) or (inputs(144)));
    layer0_outputs(2841) <= (inputs(69)) and not (inputs(204));
    layer0_outputs(2842) <= not(inputs(22)) or (inputs(65));
    layer0_outputs(2843) <= '1';
    layer0_outputs(2844) <= not(inputs(121));
    layer0_outputs(2845) <= not(inputs(222));
    layer0_outputs(2846) <= '1';
    layer0_outputs(2847) <= not(inputs(159));
    layer0_outputs(2848) <= not(inputs(212));
    layer0_outputs(2849) <= not(inputs(105)) or (inputs(79));
    layer0_outputs(2850) <= (inputs(231)) and not (inputs(14));
    layer0_outputs(2851) <= (inputs(246)) and not (inputs(146));
    layer0_outputs(2852) <= (inputs(64)) and (inputs(189));
    layer0_outputs(2853) <= (inputs(173)) xor (inputs(95));
    layer0_outputs(2854) <= not(inputs(72));
    layer0_outputs(2855) <= not((inputs(136)) or (inputs(32)));
    layer0_outputs(2856) <= '1';
    layer0_outputs(2857) <= '1';
    layer0_outputs(2858) <= (inputs(210)) and not (inputs(114));
    layer0_outputs(2859) <= (inputs(123)) and not (inputs(9));
    layer0_outputs(2860) <= not((inputs(56)) and (inputs(156)));
    layer0_outputs(2861) <= not((inputs(52)) and (inputs(157)));
    layer0_outputs(2862) <= '0';
    layer0_outputs(2863) <= not(inputs(171)) or (inputs(181));
    layer0_outputs(2864) <= not((inputs(51)) xor (inputs(77)));
    layer0_outputs(2865) <= '0';
    layer0_outputs(2866) <= '1';
    layer0_outputs(2867) <= inputs(118);
    layer0_outputs(2868) <= inputs(84);
    layer0_outputs(2869) <= inputs(55);
    layer0_outputs(2870) <= not(inputs(137)) or (inputs(75));
    layer0_outputs(2871) <= (inputs(64)) or (inputs(49));
    layer0_outputs(2872) <= (inputs(225)) xor (inputs(209));
    layer0_outputs(2873) <= inputs(11);
    layer0_outputs(2874) <= (inputs(162)) or (inputs(161));
    layer0_outputs(2875) <= not(inputs(226)) or (inputs(127));
    layer0_outputs(2876) <= (inputs(189)) and (inputs(217));
    layer0_outputs(2877) <= inputs(39);
    layer0_outputs(2878) <= inputs(8);
    layer0_outputs(2879) <= not(inputs(15)) or (inputs(215));
    layer0_outputs(2880) <= not((inputs(3)) or (inputs(131)));
    layer0_outputs(2881) <= not((inputs(66)) and (inputs(29)));
    layer0_outputs(2882) <= not(inputs(5)) or (inputs(150));
    layer0_outputs(2883) <= not((inputs(38)) or (inputs(41)));
    layer0_outputs(2884) <= inputs(38);
    layer0_outputs(2885) <= not(inputs(247));
    layer0_outputs(2886) <= inputs(55);
    layer0_outputs(2887) <= (inputs(2)) or (inputs(63));
    layer0_outputs(2888) <= (inputs(21)) and (inputs(134));
    layer0_outputs(2889) <= inputs(9);
    layer0_outputs(2890) <= inputs(230);
    layer0_outputs(2891) <= (inputs(198)) or (inputs(165));
    layer0_outputs(2892) <= not(inputs(167));
    layer0_outputs(2893) <= inputs(112);
    layer0_outputs(2894) <= (inputs(48)) or (inputs(159));
    layer0_outputs(2895) <= inputs(67);
    layer0_outputs(2896) <= not(inputs(218));
    layer0_outputs(2897) <= (inputs(35)) or (inputs(48));
    layer0_outputs(2898) <= not((inputs(61)) or (inputs(108)));
    layer0_outputs(2899) <= (inputs(125)) or (inputs(32));
    layer0_outputs(2900) <= (inputs(5)) or (inputs(255));
    layer0_outputs(2901) <= not(inputs(2));
    layer0_outputs(2902) <= not(inputs(244));
    layer0_outputs(2903) <= inputs(99);
    layer0_outputs(2904) <= (inputs(193)) and not (inputs(52));
    layer0_outputs(2905) <= not(inputs(97)) or (inputs(73));
    layer0_outputs(2906) <= (inputs(50)) and (inputs(26));
    layer0_outputs(2907) <= inputs(200);
    layer0_outputs(2908) <= inputs(18);
    layer0_outputs(2909) <= inputs(71);
    layer0_outputs(2910) <= (inputs(248)) and not (inputs(241));
    layer0_outputs(2911) <= inputs(111);
    layer0_outputs(2912) <= '0';
    layer0_outputs(2913) <= (inputs(247)) xor (inputs(143));
    layer0_outputs(2914) <= (inputs(18)) or (inputs(150));
    layer0_outputs(2915) <= not((inputs(26)) and (inputs(40)));
    layer0_outputs(2916) <= not((inputs(106)) or (inputs(147)));
    layer0_outputs(2917) <= '0';
    layer0_outputs(2918) <= '1';
    layer0_outputs(2919) <= not(inputs(124));
    layer0_outputs(2920) <= not(inputs(186));
    layer0_outputs(2921) <= (inputs(17)) and (inputs(60));
    layer0_outputs(2922) <= inputs(148);
    layer0_outputs(2923) <= not(inputs(147));
    layer0_outputs(2924) <= not((inputs(169)) or (inputs(132)));
    layer0_outputs(2925) <= not(inputs(207)) or (inputs(150));
    layer0_outputs(2926) <= not(inputs(115)) or (inputs(81));
    layer0_outputs(2927) <= (inputs(229)) and not (inputs(251));
    layer0_outputs(2928) <= (inputs(186)) xor (inputs(54));
    layer0_outputs(2929) <= not((inputs(27)) and (inputs(45)));
    layer0_outputs(2930) <= (inputs(81)) and (inputs(159));
    layer0_outputs(2931) <= not(inputs(116));
    layer0_outputs(2932) <= not(inputs(22));
    layer0_outputs(2933) <= not(inputs(170));
    layer0_outputs(2934) <= (inputs(170)) and (inputs(251));
    layer0_outputs(2935) <= '0';
    layer0_outputs(2936) <= not(inputs(143)) or (inputs(34));
    layer0_outputs(2937) <= not((inputs(161)) or (inputs(60)));
    layer0_outputs(2938) <= (inputs(137)) or (inputs(7));
    layer0_outputs(2939) <= not(inputs(76)) or (inputs(196));
    layer0_outputs(2940) <= not(inputs(181));
    layer0_outputs(2941) <= inputs(75);
    layer0_outputs(2942) <= (inputs(208)) and not (inputs(138));
    layer0_outputs(2943) <= inputs(66);
    layer0_outputs(2944) <= (inputs(103)) or (inputs(13));
    layer0_outputs(2945) <= (inputs(205)) or (inputs(213));
    layer0_outputs(2946) <= not((inputs(117)) or (inputs(96)));
    layer0_outputs(2947) <= not(inputs(158));
    layer0_outputs(2948) <= (inputs(79)) and not (inputs(217));
    layer0_outputs(2949) <= '1';
    layer0_outputs(2950) <= (inputs(17)) and not (inputs(155));
    layer0_outputs(2951) <= not(inputs(114));
    layer0_outputs(2952) <= not(inputs(155)) or (inputs(59));
    layer0_outputs(2953) <= '1';
    layer0_outputs(2954) <= inputs(163);
    layer0_outputs(2955) <= '0';
    layer0_outputs(2956) <= (inputs(198)) and (inputs(117));
    layer0_outputs(2957) <= inputs(132);
    layer0_outputs(2958) <= not((inputs(227)) or (inputs(106)));
    layer0_outputs(2959) <= inputs(246);
    layer0_outputs(2960) <= inputs(125);
    layer0_outputs(2961) <= (inputs(198)) and not (inputs(112));
    layer0_outputs(2962) <= inputs(156);
    layer0_outputs(2963) <= (inputs(246)) or (inputs(181));
    layer0_outputs(2964) <= not(inputs(103));
    layer0_outputs(2965) <= not(inputs(177));
    layer0_outputs(2966) <= '0';
    layer0_outputs(2967) <= not(inputs(247)) or (inputs(47));
    layer0_outputs(2968) <= '1';
    layer0_outputs(2969) <= not((inputs(118)) and (inputs(226)));
    layer0_outputs(2970) <= not((inputs(93)) xor (inputs(146)));
    layer0_outputs(2971) <= '1';
    layer0_outputs(2972) <= not(inputs(241));
    layer0_outputs(2973) <= not(inputs(239)) or (inputs(193));
    layer0_outputs(2974) <= (inputs(91)) or (inputs(93));
    layer0_outputs(2975) <= '1';
    layer0_outputs(2976) <= not(inputs(59)) or (inputs(87));
    layer0_outputs(2977) <= (inputs(162)) or (inputs(239));
    layer0_outputs(2978) <= '0';
    layer0_outputs(2979) <= '0';
    layer0_outputs(2980) <= '1';
    layer0_outputs(2981) <= (inputs(21)) and not (inputs(14));
    layer0_outputs(2982) <= not((inputs(23)) and (inputs(173)));
    layer0_outputs(2983) <= '0';
    layer0_outputs(2984) <= '1';
    layer0_outputs(2985) <= '0';
    layer0_outputs(2986) <= not(inputs(204)) or (inputs(44));
    layer0_outputs(2987) <= (inputs(32)) or (inputs(148));
    layer0_outputs(2988) <= (inputs(69)) and not (inputs(18));
    layer0_outputs(2989) <= (inputs(237)) or (inputs(165));
    layer0_outputs(2990) <= not((inputs(33)) xor (inputs(85)));
    layer0_outputs(2991) <= not(inputs(148));
    layer0_outputs(2992) <= not(inputs(181));
    layer0_outputs(2993) <= (inputs(117)) or (inputs(140));
    layer0_outputs(2994) <= not((inputs(233)) or (inputs(126)));
    layer0_outputs(2995) <= inputs(39);
    layer0_outputs(2996) <= not(inputs(38));
    layer0_outputs(2997) <= not((inputs(113)) or (inputs(230)));
    layer0_outputs(2998) <= (inputs(121)) and not (inputs(211));
    layer0_outputs(2999) <= '0';
    layer0_outputs(3000) <= not(inputs(0));
    layer0_outputs(3001) <= (inputs(222)) or (inputs(169));
    layer0_outputs(3002) <= not(inputs(109));
    layer0_outputs(3003) <= not(inputs(144));
    layer0_outputs(3004) <= not(inputs(234)) or (inputs(139));
    layer0_outputs(3005) <= '0';
    layer0_outputs(3006) <= not(inputs(27));
    layer0_outputs(3007) <= inputs(168);
    layer0_outputs(3008) <= inputs(15);
    layer0_outputs(3009) <= not(inputs(145));
    layer0_outputs(3010) <= not(inputs(81));
    layer0_outputs(3011) <= '0';
    layer0_outputs(3012) <= not((inputs(46)) and (inputs(232)));
    layer0_outputs(3013) <= (inputs(108)) and not (inputs(254));
    layer0_outputs(3014) <= '0';
    layer0_outputs(3015) <= inputs(27);
    layer0_outputs(3016) <= not(inputs(126));
    layer0_outputs(3017) <= '1';
    layer0_outputs(3018) <= '1';
    layer0_outputs(3019) <= inputs(166);
    layer0_outputs(3020) <= inputs(37);
    layer0_outputs(3021) <= (inputs(105)) and not (inputs(30));
    layer0_outputs(3022) <= (inputs(225)) and not (inputs(91));
    layer0_outputs(3023) <= not(inputs(85));
    layer0_outputs(3024) <= '1';
    layer0_outputs(3025) <= '0';
    layer0_outputs(3026) <= (inputs(123)) or (inputs(91));
    layer0_outputs(3027) <= '0';
    layer0_outputs(3028) <= inputs(37);
    layer0_outputs(3029) <= '0';
    layer0_outputs(3030) <= '1';
    layer0_outputs(3031) <= not(inputs(201)) or (inputs(246));
    layer0_outputs(3032) <= (inputs(120)) and not (inputs(83));
    layer0_outputs(3033) <= not((inputs(217)) or (inputs(57)));
    layer0_outputs(3034) <= not(inputs(249)) or (inputs(143));
    layer0_outputs(3035) <= not((inputs(158)) or (inputs(180)));
    layer0_outputs(3036) <= inputs(1);
    layer0_outputs(3037) <= (inputs(96)) and (inputs(1));
    layer0_outputs(3038) <= not(inputs(209));
    layer0_outputs(3039) <= (inputs(4)) or (inputs(44));
    layer0_outputs(3040) <= '0';
    layer0_outputs(3041) <= inputs(106);
    layer0_outputs(3042) <= inputs(97);
    layer0_outputs(3043) <= '0';
    layer0_outputs(3044) <= not((inputs(141)) or (inputs(123)));
    layer0_outputs(3045) <= not(inputs(47)) or (inputs(149));
    layer0_outputs(3046) <= (inputs(136)) and not (inputs(154));
    layer0_outputs(3047) <= (inputs(6)) and (inputs(50));
    layer0_outputs(3048) <= not((inputs(53)) xor (inputs(54)));
    layer0_outputs(3049) <= not((inputs(214)) xor (inputs(93)));
    layer0_outputs(3050) <= not(inputs(186));
    layer0_outputs(3051) <= (inputs(95)) or (inputs(216));
    layer0_outputs(3052) <= not(inputs(24)) or (inputs(233));
    layer0_outputs(3053) <= not(inputs(71)) or (inputs(157));
    layer0_outputs(3054) <= (inputs(133)) or (inputs(65));
    layer0_outputs(3055) <= (inputs(46)) and not (inputs(147));
    layer0_outputs(3056) <= inputs(100);
    layer0_outputs(3057) <= (inputs(126)) or (inputs(37));
    layer0_outputs(3058) <= inputs(26);
    layer0_outputs(3059) <= inputs(122);
    layer0_outputs(3060) <= (inputs(138)) or (inputs(146));
    layer0_outputs(3061) <= '0';
    layer0_outputs(3062) <= inputs(40);
    layer0_outputs(3063) <= not((inputs(223)) xor (inputs(79)));
    layer0_outputs(3064) <= not((inputs(162)) xor (inputs(35)));
    layer0_outputs(3065) <= not(inputs(178)) or (inputs(78));
    layer0_outputs(3066) <= '1';
    layer0_outputs(3067) <= inputs(107);
    layer0_outputs(3068) <= (inputs(184)) and (inputs(66));
    layer0_outputs(3069) <= not((inputs(80)) or (inputs(175)));
    layer0_outputs(3070) <= not((inputs(127)) or (inputs(82)));
    layer0_outputs(3071) <= not(inputs(148)) or (inputs(31));
    layer0_outputs(3072) <= not((inputs(17)) or (inputs(146)));
    layer0_outputs(3073) <= '0';
    layer0_outputs(3074) <= not(inputs(245));
    layer0_outputs(3075) <= not(inputs(136));
    layer0_outputs(3076) <= not(inputs(40)) or (inputs(171));
    layer0_outputs(3077) <= not(inputs(224)) or (inputs(219));
    layer0_outputs(3078) <= (inputs(67)) and not (inputs(238));
    layer0_outputs(3079) <= not((inputs(223)) or (inputs(210)));
    layer0_outputs(3080) <= not(inputs(175)) or (inputs(15));
    layer0_outputs(3081) <= not((inputs(237)) or (inputs(1)));
    layer0_outputs(3082) <= '1';
    layer0_outputs(3083) <= '1';
    layer0_outputs(3084) <= not(inputs(12)) or (inputs(85));
    layer0_outputs(3085) <= not((inputs(192)) or (inputs(133)));
    layer0_outputs(3086) <= (inputs(64)) and (inputs(62));
    layer0_outputs(3087) <= (inputs(171)) or (inputs(45));
    layer0_outputs(3088) <= (inputs(199)) and not (inputs(111));
    layer0_outputs(3089) <= (inputs(50)) or (inputs(38));
    layer0_outputs(3090) <= (inputs(182)) and not (inputs(83));
    layer0_outputs(3091) <= (inputs(120)) and not (inputs(5));
    layer0_outputs(3092) <= '1';
    layer0_outputs(3093) <= not(inputs(115));
    layer0_outputs(3094) <= not(inputs(84));
    layer0_outputs(3095) <= not((inputs(235)) or (inputs(222)));
    layer0_outputs(3096) <= not(inputs(70)) or (inputs(146));
    layer0_outputs(3097) <= (inputs(10)) and (inputs(39));
    layer0_outputs(3098) <= (inputs(91)) and (inputs(219));
    layer0_outputs(3099) <= (inputs(113)) xor (inputs(50));
    layer0_outputs(3100) <= (inputs(76)) and not (inputs(50));
    layer0_outputs(3101) <= not(inputs(165)) or (inputs(31));
    layer0_outputs(3102) <= not((inputs(189)) and (inputs(202)));
    layer0_outputs(3103) <= not(inputs(99));
    layer0_outputs(3104) <= not(inputs(51));
    layer0_outputs(3105) <= not((inputs(41)) or (inputs(34)));
    layer0_outputs(3106) <= inputs(241);
    layer0_outputs(3107) <= not(inputs(90));
    layer0_outputs(3108) <= '0';
    layer0_outputs(3109) <= inputs(122);
    layer0_outputs(3110) <= inputs(86);
    layer0_outputs(3111) <= not((inputs(179)) or (inputs(197)));
    layer0_outputs(3112) <= '1';
    layer0_outputs(3113) <= '1';
    layer0_outputs(3114) <= not(inputs(50));
    layer0_outputs(3115) <= not(inputs(54)) or (inputs(230));
    layer0_outputs(3116) <= inputs(127);
    layer0_outputs(3117) <= not((inputs(219)) or (inputs(31)));
    layer0_outputs(3118) <= not(inputs(117)) or (inputs(40));
    layer0_outputs(3119) <= '0';
    layer0_outputs(3120) <= not(inputs(132)) or (inputs(126));
    layer0_outputs(3121) <= '0';
    layer0_outputs(3122) <= not(inputs(82));
    layer0_outputs(3123) <= not((inputs(80)) and (inputs(89)));
    layer0_outputs(3124) <= not(inputs(106)) or (inputs(226));
    layer0_outputs(3125) <= not(inputs(105));
    layer0_outputs(3126) <= (inputs(150)) and not (inputs(13));
    layer0_outputs(3127) <= (inputs(172)) and not (inputs(87));
    layer0_outputs(3128) <= not((inputs(212)) or (inputs(221)));
    layer0_outputs(3129) <= '1';
    layer0_outputs(3130) <= not((inputs(154)) xor (inputs(93)));
    layer0_outputs(3131) <= not((inputs(79)) xor (inputs(143)));
    layer0_outputs(3132) <= '1';
    layer0_outputs(3133) <= not(inputs(4));
    layer0_outputs(3134) <= (inputs(99)) and not (inputs(104));
    layer0_outputs(3135) <= (inputs(255)) and (inputs(6));
    layer0_outputs(3136) <= inputs(158);
    layer0_outputs(3137) <= not((inputs(221)) or (inputs(162)));
    layer0_outputs(3138) <= inputs(149);
    layer0_outputs(3139) <= not((inputs(241)) and (inputs(92)));
    layer0_outputs(3140) <= '0';
    layer0_outputs(3141) <= (inputs(255)) and not (inputs(101));
    layer0_outputs(3142) <= '1';
    layer0_outputs(3143) <= not((inputs(162)) or (inputs(36)));
    layer0_outputs(3144) <= (inputs(180)) or (inputs(183));
    layer0_outputs(3145) <= (inputs(79)) and not (inputs(225));
    layer0_outputs(3146) <= (inputs(122)) and not (inputs(200));
    layer0_outputs(3147) <= '0';
    layer0_outputs(3148) <= not(inputs(197)) or (inputs(42));
    layer0_outputs(3149) <= not(inputs(68)) or (inputs(77));
    layer0_outputs(3150) <= (inputs(125)) and (inputs(252));
    layer0_outputs(3151) <= inputs(214);
    layer0_outputs(3152) <= (inputs(98)) xor (inputs(172));
    layer0_outputs(3153) <= inputs(85);
    layer0_outputs(3154) <= '0';
    layer0_outputs(3155) <= (inputs(62)) and not (inputs(11));
    layer0_outputs(3156) <= not(inputs(95)) or (inputs(49));
    layer0_outputs(3157) <= inputs(223);
    layer0_outputs(3158) <= (inputs(189)) and not (inputs(14));
    layer0_outputs(3159) <= not((inputs(213)) xor (inputs(32)));
    layer0_outputs(3160) <= '1';
    layer0_outputs(3161) <= (inputs(111)) or (inputs(144));
    layer0_outputs(3162) <= inputs(65);
    layer0_outputs(3163) <= not(inputs(94));
    layer0_outputs(3164) <= '1';
    layer0_outputs(3165) <= not(inputs(84)) or (inputs(143));
    layer0_outputs(3166) <= inputs(106);
    layer0_outputs(3167) <= not(inputs(237));
    layer0_outputs(3168) <= (inputs(79)) xor (inputs(19));
    layer0_outputs(3169) <= '0';
    layer0_outputs(3170) <= inputs(165);
    layer0_outputs(3171) <= not((inputs(192)) or (inputs(93)));
    layer0_outputs(3172) <= not(inputs(56));
    layer0_outputs(3173) <= inputs(148);
    layer0_outputs(3174) <= inputs(218);
    layer0_outputs(3175) <= (inputs(192)) and not (inputs(15));
    layer0_outputs(3176) <= not(inputs(15));
    layer0_outputs(3177) <= not((inputs(36)) and (inputs(166)));
    layer0_outputs(3178) <= not(inputs(209)) or (inputs(168));
    layer0_outputs(3179) <= not(inputs(226)) or (inputs(97));
    layer0_outputs(3180) <= not(inputs(224)) or (inputs(180));
    layer0_outputs(3181) <= inputs(3);
    layer0_outputs(3182) <= not(inputs(177));
    layer0_outputs(3183) <= inputs(212);
    layer0_outputs(3184) <= not(inputs(119));
    layer0_outputs(3185) <= not((inputs(32)) or (inputs(129)));
    layer0_outputs(3186) <= (inputs(234)) and not (inputs(19));
    layer0_outputs(3187) <= (inputs(186)) xor (inputs(135));
    layer0_outputs(3188) <= not(inputs(24)) or (inputs(25));
    layer0_outputs(3189) <= (inputs(101)) or (inputs(126));
    layer0_outputs(3190) <= '1';
    layer0_outputs(3191) <= (inputs(133)) or (inputs(118));
    layer0_outputs(3192) <= (inputs(177)) and (inputs(6));
    layer0_outputs(3193) <= not((inputs(249)) and (inputs(181)));
    layer0_outputs(3194) <= not(inputs(89)) or (inputs(26));
    layer0_outputs(3195) <= not(inputs(234));
    layer0_outputs(3196) <= '1';
    layer0_outputs(3197) <= '1';
    layer0_outputs(3198) <= (inputs(179)) and not (inputs(238));
    layer0_outputs(3199) <= not((inputs(29)) or (inputs(124)));
    layer0_outputs(3200) <= (inputs(192)) or (inputs(175));
    layer0_outputs(3201) <= not(inputs(53));
    layer0_outputs(3202) <= not((inputs(255)) or (inputs(181)));
    layer0_outputs(3203) <= (inputs(73)) and (inputs(154));
    layer0_outputs(3204) <= not(inputs(3));
    layer0_outputs(3205) <= (inputs(179)) and not (inputs(159));
    layer0_outputs(3206) <= inputs(100);
    layer0_outputs(3207) <= inputs(71);
    layer0_outputs(3208) <= (inputs(209)) or (inputs(233));
    layer0_outputs(3209) <= '1';
    layer0_outputs(3210) <= '1';
    layer0_outputs(3211) <= not(inputs(178)) or (inputs(21));
    layer0_outputs(3212) <= not((inputs(83)) and (inputs(154)));
    layer0_outputs(3213) <= '0';
    layer0_outputs(3214) <= (inputs(150)) and not (inputs(108));
    layer0_outputs(3215) <= (inputs(84)) or (inputs(183));
    layer0_outputs(3216) <= inputs(149);
    layer0_outputs(3217) <= inputs(178);
    layer0_outputs(3218) <= (inputs(24)) and not (inputs(81));
    layer0_outputs(3219) <= (inputs(250)) and not (inputs(247));
    layer0_outputs(3220) <= '1';
    layer0_outputs(3221) <= not(inputs(119)) or (inputs(148));
    layer0_outputs(3222) <= inputs(223);
    layer0_outputs(3223) <= not((inputs(159)) xor (inputs(182)));
    layer0_outputs(3224) <= not((inputs(181)) or (inputs(115)));
    layer0_outputs(3225) <= '0';
    layer0_outputs(3226) <= '1';
    layer0_outputs(3227) <= (inputs(114)) and not (inputs(238));
    layer0_outputs(3228) <= not(inputs(39)) or (inputs(204));
    layer0_outputs(3229) <= '1';
    layer0_outputs(3230) <= not((inputs(236)) xor (inputs(157)));
    layer0_outputs(3231) <= (inputs(155)) and (inputs(191));
    layer0_outputs(3232) <= inputs(153);
    layer0_outputs(3233) <= not(inputs(22)) or (inputs(238));
    layer0_outputs(3234) <= '1';
    layer0_outputs(3235) <= not(inputs(226)) or (inputs(23));
    layer0_outputs(3236) <= inputs(30);
    layer0_outputs(3237) <= not((inputs(53)) and (inputs(24)));
    layer0_outputs(3238) <= not((inputs(4)) or (inputs(246)));
    layer0_outputs(3239) <= '0';
    layer0_outputs(3240) <= '1';
    layer0_outputs(3241) <= (inputs(238)) or (inputs(38));
    layer0_outputs(3242) <= '1';
    layer0_outputs(3243) <= '1';
    layer0_outputs(3244) <= not((inputs(239)) and (inputs(216)));
    layer0_outputs(3245) <= '1';
    layer0_outputs(3246) <= not(inputs(121));
    layer0_outputs(3247) <= inputs(32);
    layer0_outputs(3248) <= '1';
    layer0_outputs(3249) <= (inputs(163)) and not (inputs(253));
    layer0_outputs(3250) <= not(inputs(123)) or (inputs(168));
    layer0_outputs(3251) <= not((inputs(183)) or (inputs(49)));
    layer0_outputs(3252) <= (inputs(184)) and (inputs(50));
    layer0_outputs(3253) <= (inputs(61)) and (inputs(113));
    layer0_outputs(3254) <= '1';
    layer0_outputs(3255) <= '1';
    layer0_outputs(3256) <= not(inputs(116)) or (inputs(200));
    layer0_outputs(3257) <= not(inputs(136));
    layer0_outputs(3258) <= '1';
    layer0_outputs(3259) <= not((inputs(237)) or (inputs(20)));
    layer0_outputs(3260) <= (inputs(133)) and not (inputs(18));
    layer0_outputs(3261) <= (inputs(198)) and (inputs(211));
    layer0_outputs(3262) <= (inputs(47)) or (inputs(190));
    layer0_outputs(3263) <= '0';
    layer0_outputs(3264) <= inputs(14);
    layer0_outputs(3265) <= not(inputs(190));
    layer0_outputs(3266) <= (inputs(245)) and (inputs(129));
    layer0_outputs(3267) <= not((inputs(59)) and (inputs(189)));
    layer0_outputs(3268) <= inputs(198);
    layer0_outputs(3269) <= not(inputs(214)) or (inputs(90));
    layer0_outputs(3270) <= not(inputs(149)) or (inputs(141));
    layer0_outputs(3271) <= not(inputs(151)) or (inputs(111));
    layer0_outputs(3272) <= not((inputs(145)) or (inputs(86)));
    layer0_outputs(3273) <= not(inputs(125));
    layer0_outputs(3274) <= not(inputs(207));
    layer0_outputs(3275) <= inputs(178);
    layer0_outputs(3276) <= (inputs(125)) and not (inputs(215));
    layer0_outputs(3277) <= (inputs(107)) and not (inputs(117));
    layer0_outputs(3278) <= inputs(113);
    layer0_outputs(3279) <= '1';
    layer0_outputs(3280) <= inputs(254);
    layer0_outputs(3281) <= not(inputs(143));
    layer0_outputs(3282) <= (inputs(118)) and not (inputs(85));
    layer0_outputs(3283) <= (inputs(75)) and not (inputs(24));
    layer0_outputs(3284) <= not((inputs(143)) and (inputs(78)));
    layer0_outputs(3285) <= inputs(3);
    layer0_outputs(3286) <= not(inputs(46));
    layer0_outputs(3287) <= inputs(108);
    layer0_outputs(3288) <= not(inputs(217)) or (inputs(109));
    layer0_outputs(3289) <= not(inputs(43));
    layer0_outputs(3290) <= not(inputs(93)) or (inputs(124));
    layer0_outputs(3291) <= not((inputs(174)) and (inputs(185)));
    layer0_outputs(3292) <= not(inputs(252)) or (inputs(109));
    layer0_outputs(3293) <= (inputs(190)) and not (inputs(228));
    layer0_outputs(3294) <= not((inputs(126)) or (inputs(22)));
    layer0_outputs(3295) <= (inputs(119)) and not (inputs(66));
    layer0_outputs(3296) <= '1';
    layer0_outputs(3297) <= '0';
    layer0_outputs(3298) <= '1';
    layer0_outputs(3299) <= inputs(90);
    layer0_outputs(3300) <= (inputs(141)) and (inputs(198));
    layer0_outputs(3301) <= not((inputs(240)) or (inputs(224)));
    layer0_outputs(3302) <= not((inputs(181)) xor (inputs(119)));
    layer0_outputs(3303) <= (inputs(137)) and not (inputs(5));
    layer0_outputs(3304) <= not((inputs(51)) and (inputs(155)));
    layer0_outputs(3305) <= not(inputs(152)) or (inputs(113));
    layer0_outputs(3306) <= inputs(65);
    layer0_outputs(3307) <= '1';
    layer0_outputs(3308) <= not(inputs(73));
    layer0_outputs(3309) <= not(inputs(107)) or (inputs(210));
    layer0_outputs(3310) <= not(inputs(45)) or (inputs(2));
    layer0_outputs(3311) <= '0';
    layer0_outputs(3312) <= not(inputs(197)) or (inputs(97));
    layer0_outputs(3313) <= '0';
    layer0_outputs(3314) <= not(inputs(112));
    layer0_outputs(3315) <= not(inputs(130)) or (inputs(208));
    layer0_outputs(3316) <= not((inputs(102)) or (inputs(189)));
    layer0_outputs(3317) <= not(inputs(185));
    layer0_outputs(3318) <= '0';
    layer0_outputs(3319) <= (inputs(20)) and not (inputs(76));
    layer0_outputs(3320) <= '1';
    layer0_outputs(3321) <= not((inputs(96)) and (inputs(103)));
    layer0_outputs(3322) <= inputs(196);
    layer0_outputs(3323) <= not(inputs(75));
    layer0_outputs(3324) <= '1';
    layer0_outputs(3325) <= not(inputs(122));
    layer0_outputs(3326) <= not(inputs(115)) or (inputs(207));
    layer0_outputs(3327) <= (inputs(166)) and (inputs(140));
    layer0_outputs(3328) <= inputs(128);
    layer0_outputs(3329) <= not(inputs(80));
    layer0_outputs(3330) <= inputs(23);
    layer0_outputs(3331) <= not((inputs(34)) and (inputs(6)));
    layer0_outputs(3332) <= not(inputs(101)) or (inputs(123));
    layer0_outputs(3333) <= not((inputs(215)) or (inputs(87)));
    layer0_outputs(3334) <= not((inputs(139)) or (inputs(156)));
    layer0_outputs(3335) <= '0';
    layer0_outputs(3336) <= not(inputs(73));
    layer0_outputs(3337) <= not((inputs(2)) and (inputs(49)));
    layer0_outputs(3338) <= not(inputs(14));
    layer0_outputs(3339) <= '1';
    layer0_outputs(3340) <= not(inputs(129)) or (inputs(224));
    layer0_outputs(3341) <= not((inputs(48)) xor (inputs(18)));
    layer0_outputs(3342) <= '0';
    layer0_outputs(3343) <= not(inputs(115));
    layer0_outputs(3344) <= not((inputs(93)) and (inputs(1)));
    layer0_outputs(3345) <= not(inputs(218));
    layer0_outputs(3346) <= inputs(193);
    layer0_outputs(3347) <= not(inputs(224));
    layer0_outputs(3348) <= '1';
    layer0_outputs(3349) <= inputs(231);
    layer0_outputs(3350) <= (inputs(17)) or (inputs(43));
    layer0_outputs(3351) <= inputs(213);
    layer0_outputs(3352) <= not(inputs(120)) or (inputs(192));
    layer0_outputs(3353) <= inputs(243);
    layer0_outputs(3354) <= inputs(121);
    layer0_outputs(3355) <= not((inputs(22)) or (inputs(58)));
    layer0_outputs(3356) <= not(inputs(221));
    layer0_outputs(3357) <= (inputs(168)) or (inputs(126));
    layer0_outputs(3358) <= '1';
    layer0_outputs(3359) <= not(inputs(192)) or (inputs(197));
    layer0_outputs(3360) <= '1';
    layer0_outputs(3361) <= not((inputs(33)) or (inputs(72)));
    layer0_outputs(3362) <= not(inputs(107)) or (inputs(41));
    layer0_outputs(3363) <= '1';
    layer0_outputs(3364) <= (inputs(144)) or (inputs(214));
    layer0_outputs(3365) <= inputs(227);
    layer0_outputs(3366) <= not(inputs(32)) or (inputs(153));
    layer0_outputs(3367) <= not((inputs(13)) or (inputs(60)));
    layer0_outputs(3368) <= not(inputs(204));
    layer0_outputs(3369) <= '0';
    layer0_outputs(3370) <= '1';
    layer0_outputs(3371) <= inputs(238);
    layer0_outputs(3372) <= '0';
    layer0_outputs(3373) <= not(inputs(143));
    layer0_outputs(3374) <= inputs(180);
    layer0_outputs(3375) <= not((inputs(227)) xor (inputs(238)));
    layer0_outputs(3376) <= not((inputs(63)) and (inputs(59)));
    layer0_outputs(3377) <= inputs(57);
    layer0_outputs(3378) <= inputs(177);
    layer0_outputs(3379) <= not(inputs(78));
    layer0_outputs(3380) <= (inputs(86)) or (inputs(201));
    layer0_outputs(3381) <= not(inputs(43));
    layer0_outputs(3382) <= (inputs(11)) and (inputs(194));
    layer0_outputs(3383) <= inputs(85);
    layer0_outputs(3384) <= '1';
    layer0_outputs(3385) <= (inputs(53)) and not (inputs(187));
    layer0_outputs(3386) <= not((inputs(27)) and (inputs(40)));
    layer0_outputs(3387) <= not((inputs(115)) and (inputs(26)));
    layer0_outputs(3388) <= not(inputs(24));
    layer0_outputs(3389) <= not(inputs(158)) or (inputs(115));
    layer0_outputs(3390) <= (inputs(105)) and not (inputs(24));
    layer0_outputs(3391) <= inputs(38);
    layer0_outputs(3392) <= not(inputs(8));
    layer0_outputs(3393) <= not(inputs(68));
    layer0_outputs(3394) <= not(inputs(101));
    layer0_outputs(3395) <= (inputs(202)) or (inputs(212));
    layer0_outputs(3396) <= inputs(61);
    layer0_outputs(3397) <= inputs(140);
    layer0_outputs(3398) <= not(inputs(88)) or (inputs(241));
    layer0_outputs(3399) <= '1';
    layer0_outputs(3400) <= not(inputs(120));
    layer0_outputs(3401) <= (inputs(47)) xor (inputs(230));
    layer0_outputs(3402) <= (inputs(207)) and not (inputs(32));
    layer0_outputs(3403) <= '1';
    layer0_outputs(3404) <= (inputs(227)) and not (inputs(251));
    layer0_outputs(3405) <= inputs(101);
    layer0_outputs(3406) <= inputs(179);
    layer0_outputs(3407) <= (inputs(71)) and not (inputs(254));
    layer0_outputs(3408) <= not(inputs(216));
    layer0_outputs(3409) <= not((inputs(157)) or (inputs(7)));
    layer0_outputs(3410) <= inputs(36);
    layer0_outputs(3411) <= '0';
    layer0_outputs(3412) <= (inputs(185)) and (inputs(179));
    layer0_outputs(3413) <= not((inputs(140)) or (inputs(59)));
    layer0_outputs(3414) <= (inputs(247)) and not (inputs(7));
    layer0_outputs(3415) <= '1';
    layer0_outputs(3416) <= inputs(131);
    layer0_outputs(3417) <= (inputs(8)) xor (inputs(128));
    layer0_outputs(3418) <= (inputs(157)) or (inputs(219));
    layer0_outputs(3419) <= not(inputs(136));
    layer0_outputs(3420) <= inputs(7);
    layer0_outputs(3421) <= not(inputs(127)) or (inputs(165));
    layer0_outputs(3422) <= inputs(73);
    layer0_outputs(3423) <= not((inputs(204)) and (inputs(14)));
    layer0_outputs(3424) <= (inputs(55)) or (inputs(196));
    layer0_outputs(3425) <= not((inputs(174)) and (inputs(174)));
    layer0_outputs(3426) <= inputs(227);
    layer0_outputs(3427) <= not(inputs(9));
    layer0_outputs(3428) <= not(inputs(5));
    layer0_outputs(3429) <= not((inputs(3)) or (inputs(22)));
    layer0_outputs(3430) <= '0';
    layer0_outputs(3431) <= not(inputs(117));
    layer0_outputs(3432) <= '0';
    layer0_outputs(3433) <= '1';
    layer0_outputs(3434) <= inputs(26);
    layer0_outputs(3435) <= (inputs(231)) and not (inputs(101));
    layer0_outputs(3436) <= not(inputs(32));
    layer0_outputs(3437) <= '0';
    layer0_outputs(3438) <= not((inputs(164)) or (inputs(217)));
    layer0_outputs(3439) <= inputs(28);
    layer0_outputs(3440) <= inputs(157);
    layer0_outputs(3441) <= not(inputs(198));
    layer0_outputs(3442) <= not(inputs(135)) or (inputs(192));
    layer0_outputs(3443) <= (inputs(125)) and not (inputs(138));
    layer0_outputs(3444) <= not(inputs(63));
    layer0_outputs(3445) <= (inputs(206)) or (inputs(193));
    layer0_outputs(3446) <= not((inputs(227)) or (inputs(224)));
    layer0_outputs(3447) <= not(inputs(194));
    layer0_outputs(3448) <= not((inputs(194)) xor (inputs(150)));
    layer0_outputs(3449) <= (inputs(144)) and not (inputs(130));
    layer0_outputs(3450) <= not((inputs(79)) xor (inputs(47)));
    layer0_outputs(3451) <= inputs(155);
    layer0_outputs(3452) <= not(inputs(175)) or (inputs(23));
    layer0_outputs(3453) <= (inputs(144)) or (inputs(130));
    layer0_outputs(3454) <= (inputs(65)) xor (inputs(239));
    layer0_outputs(3455) <= inputs(24);
    layer0_outputs(3456) <= not(inputs(83));
    layer0_outputs(3457) <= not(inputs(148)) or (inputs(40));
    layer0_outputs(3458) <= not(inputs(106));
    layer0_outputs(3459) <= (inputs(21)) and not (inputs(241));
    layer0_outputs(3460) <= inputs(68);
    layer0_outputs(3461) <= (inputs(162)) and (inputs(177));
    layer0_outputs(3462) <= '0';
    layer0_outputs(3463) <= (inputs(216)) or (inputs(33));
    layer0_outputs(3464) <= (inputs(139)) and not (inputs(254));
    layer0_outputs(3465) <= '1';
    layer0_outputs(3466) <= not(inputs(14));
    layer0_outputs(3467) <= not(inputs(177));
    layer0_outputs(3468) <= not(inputs(56));
    layer0_outputs(3469) <= not(inputs(197)) or (inputs(135));
    layer0_outputs(3470) <= not((inputs(137)) xor (inputs(137)));
    layer0_outputs(3471) <= not(inputs(31));
    layer0_outputs(3472) <= not(inputs(18));
    layer0_outputs(3473) <= inputs(104);
    layer0_outputs(3474) <= not((inputs(55)) or (inputs(160)));
    layer0_outputs(3475) <= inputs(8);
    layer0_outputs(3476) <= inputs(113);
    layer0_outputs(3477) <= inputs(13);
    layer0_outputs(3478) <= (inputs(21)) and not (inputs(52));
    layer0_outputs(3479) <= inputs(245);
    layer0_outputs(3480) <= not(inputs(35));
    layer0_outputs(3481) <= inputs(226);
    layer0_outputs(3482) <= '1';
    layer0_outputs(3483) <= inputs(41);
    layer0_outputs(3484) <= not(inputs(208)) or (inputs(116));
    layer0_outputs(3485) <= (inputs(196)) and (inputs(185));
    layer0_outputs(3486) <= not((inputs(157)) or (inputs(4)));
    layer0_outputs(3487) <= (inputs(243)) and (inputs(189));
    layer0_outputs(3488) <= '1';
    layer0_outputs(3489) <= not((inputs(71)) xor (inputs(83)));
    layer0_outputs(3490) <= '1';
    layer0_outputs(3491) <= inputs(219);
    layer0_outputs(3492) <= (inputs(165)) and (inputs(35));
    layer0_outputs(3493) <= '1';
    layer0_outputs(3494) <= not((inputs(219)) or (inputs(238)));
    layer0_outputs(3495) <= (inputs(156)) and not (inputs(120));
    layer0_outputs(3496) <= not(inputs(1)) or (inputs(163));
    layer0_outputs(3497) <= (inputs(112)) and not (inputs(143));
    layer0_outputs(3498) <= (inputs(81)) and (inputs(5));
    layer0_outputs(3499) <= not(inputs(160));
    layer0_outputs(3500) <= not((inputs(145)) and (inputs(71)));
    layer0_outputs(3501) <= not(inputs(198)) or (inputs(28));
    layer0_outputs(3502) <= not((inputs(235)) and (inputs(41)));
    layer0_outputs(3503) <= '1';
    layer0_outputs(3504) <= not(inputs(164));
    layer0_outputs(3505) <= '0';
    layer0_outputs(3506) <= inputs(75);
    layer0_outputs(3507) <= (inputs(163)) or (inputs(209));
    layer0_outputs(3508) <= '0';
    layer0_outputs(3509) <= '0';
    layer0_outputs(3510) <= not(inputs(24)) or (inputs(87));
    layer0_outputs(3511) <= not((inputs(106)) or (inputs(93)));
    layer0_outputs(3512) <= inputs(182);
    layer0_outputs(3513) <= not(inputs(146));
    layer0_outputs(3514) <= not(inputs(100)) or (inputs(178));
    layer0_outputs(3515) <= '0';
    layer0_outputs(3516) <= (inputs(219)) and not (inputs(55));
    layer0_outputs(3517) <= inputs(130);
    layer0_outputs(3518) <= inputs(215);
    layer0_outputs(3519) <= (inputs(241)) and not (inputs(57));
    layer0_outputs(3520) <= not((inputs(179)) or (inputs(252)));
    layer0_outputs(3521) <= not(inputs(118));
    layer0_outputs(3522) <= not(inputs(137));
    layer0_outputs(3523) <= not((inputs(140)) and (inputs(186)));
    layer0_outputs(3524) <= not(inputs(254));
    layer0_outputs(3525) <= (inputs(59)) and not (inputs(244));
    layer0_outputs(3526) <= not(inputs(111)) or (inputs(224));
    layer0_outputs(3527) <= not(inputs(159));
    layer0_outputs(3528) <= not((inputs(88)) and (inputs(86)));
    layer0_outputs(3529) <= inputs(223);
    layer0_outputs(3530) <= not(inputs(252));
    layer0_outputs(3531) <= '0';
    layer0_outputs(3532) <= (inputs(59)) and (inputs(136));
    layer0_outputs(3533) <= (inputs(6)) and not (inputs(164));
    layer0_outputs(3534) <= inputs(38);
    layer0_outputs(3535) <= not(inputs(90));
    layer0_outputs(3536) <= '0';
    layer0_outputs(3537) <= inputs(106);
    layer0_outputs(3538) <= not(inputs(37)) or (inputs(115));
    layer0_outputs(3539) <= (inputs(213)) and not (inputs(107));
    layer0_outputs(3540) <= inputs(97);
    layer0_outputs(3541) <= '0';
    layer0_outputs(3542) <= not((inputs(151)) or (inputs(196)));
    layer0_outputs(3543) <= not((inputs(80)) or (inputs(94)));
    layer0_outputs(3544) <= not((inputs(53)) or (inputs(22)));
    layer0_outputs(3545) <= not((inputs(212)) or (inputs(221)));
    layer0_outputs(3546) <= not(inputs(211));
    layer0_outputs(3547) <= not((inputs(104)) or (inputs(58)));
    layer0_outputs(3548) <= inputs(24);
    layer0_outputs(3549) <= (inputs(219)) or (inputs(122));
    layer0_outputs(3550) <= inputs(161);
    layer0_outputs(3551) <= '0';
    layer0_outputs(3552) <= '0';
    layer0_outputs(3553) <= inputs(136);
    layer0_outputs(3554) <= inputs(237);
    layer0_outputs(3555) <= not((inputs(216)) and (inputs(91)));
    layer0_outputs(3556) <= '0';
    layer0_outputs(3557) <= not(inputs(39)) or (inputs(189));
    layer0_outputs(3558) <= '0';
    layer0_outputs(3559) <= inputs(129);
    layer0_outputs(3560) <= (inputs(187)) xor (inputs(252));
    layer0_outputs(3561) <= (inputs(63)) and not (inputs(188));
    layer0_outputs(3562) <= inputs(241);
    layer0_outputs(3563) <= '1';
    layer0_outputs(3564) <= inputs(141);
    layer0_outputs(3565) <= not((inputs(80)) or (inputs(82)));
    layer0_outputs(3566) <= inputs(43);
    layer0_outputs(3567) <= (inputs(240)) xor (inputs(169));
    layer0_outputs(3568) <= (inputs(7)) and not (inputs(45));
    layer0_outputs(3569) <= not(inputs(138)) or (inputs(226));
    layer0_outputs(3570) <= (inputs(67)) xor (inputs(18));
    layer0_outputs(3571) <= inputs(88);
    layer0_outputs(3572) <= not((inputs(149)) or (inputs(184)));
    layer0_outputs(3573) <= not(inputs(88)) or (inputs(73));
    layer0_outputs(3574) <= (inputs(4)) or (inputs(192));
    layer0_outputs(3575) <= not(inputs(102));
    layer0_outputs(3576) <= not((inputs(1)) and (inputs(186)));
    layer0_outputs(3577) <= not(inputs(124));
    layer0_outputs(3578) <= inputs(203);
    layer0_outputs(3579) <= not(inputs(171));
    layer0_outputs(3580) <= '0';
    layer0_outputs(3581) <= not(inputs(169));
    layer0_outputs(3582) <= inputs(212);
    layer0_outputs(3583) <= not(inputs(21)) or (inputs(218));
    layer0_outputs(3584) <= not(inputs(7));
    layer0_outputs(3585) <= (inputs(196)) xor (inputs(3));
    layer0_outputs(3586) <= not(inputs(120));
    layer0_outputs(3587) <= not((inputs(187)) or (inputs(170)));
    layer0_outputs(3588) <= not(inputs(110));
    layer0_outputs(3589) <= '0';
    layer0_outputs(3590) <= (inputs(121)) and not (inputs(219));
    layer0_outputs(3591) <= '0';
    layer0_outputs(3592) <= not(inputs(50)) or (inputs(113));
    layer0_outputs(3593) <= not((inputs(144)) or (inputs(177)));
    layer0_outputs(3594) <= '0';
    layer0_outputs(3595) <= not(inputs(231));
    layer0_outputs(3596) <= '0';
    layer0_outputs(3597) <= (inputs(195)) or (inputs(237));
    layer0_outputs(3598) <= not(inputs(194)) or (inputs(47));
    layer0_outputs(3599) <= inputs(133);
    layer0_outputs(3600) <= not(inputs(245)) or (inputs(8));
    layer0_outputs(3601) <= not(inputs(55)) or (inputs(210));
    layer0_outputs(3602) <= not(inputs(85));
    layer0_outputs(3603) <= inputs(151);
    layer0_outputs(3604) <= '1';
    layer0_outputs(3605) <= (inputs(102)) and (inputs(253));
    layer0_outputs(3606) <= (inputs(58)) and (inputs(201));
    layer0_outputs(3607) <= '0';
    layer0_outputs(3608) <= (inputs(90)) and not (inputs(31));
    layer0_outputs(3609) <= not((inputs(96)) or (inputs(89)));
    layer0_outputs(3610) <= not(inputs(101)) or (inputs(175));
    layer0_outputs(3611) <= not((inputs(128)) and (inputs(39)));
    layer0_outputs(3612) <= not(inputs(99));
    layer0_outputs(3613) <= not(inputs(15)) or (inputs(1));
    layer0_outputs(3614) <= not(inputs(252)) or (inputs(204));
    layer0_outputs(3615) <= (inputs(26)) or (inputs(107));
    layer0_outputs(3616) <= inputs(3);
    layer0_outputs(3617) <= not((inputs(217)) or (inputs(170)));
    layer0_outputs(3618) <= not(inputs(51));
    layer0_outputs(3619) <= (inputs(149)) and not (inputs(154));
    layer0_outputs(3620) <= '1';
    layer0_outputs(3621) <= not((inputs(140)) or (inputs(24)));
    layer0_outputs(3622) <= not(inputs(140)) or (inputs(5));
    layer0_outputs(3623) <= '1';
    layer0_outputs(3624) <= inputs(89);
    layer0_outputs(3625) <= (inputs(47)) and not (inputs(255));
    layer0_outputs(3626) <= not((inputs(78)) and (inputs(185)));
    layer0_outputs(3627) <= (inputs(229)) and not (inputs(73));
    layer0_outputs(3628) <= (inputs(73)) and not (inputs(251));
    layer0_outputs(3629) <= (inputs(50)) and (inputs(4));
    layer0_outputs(3630) <= not(inputs(112));
    layer0_outputs(3631) <= not(inputs(217));
    layer0_outputs(3632) <= not(inputs(126));
    layer0_outputs(3633) <= '0';
    layer0_outputs(3634) <= '0';
    layer0_outputs(3635) <= (inputs(234)) and not (inputs(94));
    layer0_outputs(3636) <= (inputs(195)) and not (inputs(208));
    layer0_outputs(3637) <= not((inputs(178)) or (inputs(70)));
    layer0_outputs(3638) <= not(inputs(156));
    layer0_outputs(3639) <= '1';
    layer0_outputs(3640) <= inputs(233);
    layer0_outputs(3641) <= (inputs(179)) and not (inputs(56));
    layer0_outputs(3642) <= (inputs(204)) and not (inputs(12));
    layer0_outputs(3643) <= (inputs(121)) and not (inputs(7));
    layer0_outputs(3644) <= '0';
    layer0_outputs(3645) <= (inputs(36)) or (inputs(125));
    layer0_outputs(3646) <= not(inputs(63)) or (inputs(37));
    layer0_outputs(3647) <= '0';
    layer0_outputs(3648) <= '0';
    layer0_outputs(3649) <= inputs(83);
    layer0_outputs(3650) <= '1';
    layer0_outputs(3651) <= not(inputs(199)) or (inputs(74));
    layer0_outputs(3652) <= '0';
    layer0_outputs(3653) <= '0';
    layer0_outputs(3654) <= not(inputs(153));
    layer0_outputs(3655) <= not(inputs(146));
    layer0_outputs(3656) <= not((inputs(171)) or (inputs(47)));
    layer0_outputs(3657) <= not(inputs(8));
    layer0_outputs(3658) <= '1';
    layer0_outputs(3659) <= not(inputs(80));
    layer0_outputs(3660) <= not(inputs(88)) or (inputs(127));
    layer0_outputs(3661) <= (inputs(17)) and (inputs(143));
    layer0_outputs(3662) <= (inputs(199)) and (inputs(39));
    layer0_outputs(3663) <= not(inputs(51)) or (inputs(55));
    layer0_outputs(3664) <= (inputs(126)) or (inputs(78));
    layer0_outputs(3665) <= not(inputs(105)) or (inputs(177));
    layer0_outputs(3666) <= (inputs(167)) and not (inputs(69));
    layer0_outputs(3667) <= (inputs(149)) or (inputs(240));
    layer0_outputs(3668) <= inputs(199);
    layer0_outputs(3669) <= '0';
    layer0_outputs(3670) <= not((inputs(227)) or (inputs(222)));
    layer0_outputs(3671) <= (inputs(234)) and (inputs(198));
    layer0_outputs(3672) <= not(inputs(54));
    layer0_outputs(3673) <= '0';
    layer0_outputs(3674) <= (inputs(197)) and not (inputs(74));
    layer0_outputs(3675) <= (inputs(105)) and (inputs(220));
    layer0_outputs(3676) <= (inputs(246)) xor (inputs(196));
    layer0_outputs(3677) <= (inputs(229)) or (inputs(212));
    layer0_outputs(3678) <= not(inputs(190)) or (inputs(81));
    layer0_outputs(3679) <= (inputs(179)) or (inputs(221));
    layer0_outputs(3680) <= (inputs(235)) or (inputs(189));
    layer0_outputs(3681) <= not((inputs(19)) or (inputs(249)));
    layer0_outputs(3682) <= not(inputs(0)) or (inputs(238));
    layer0_outputs(3683) <= not((inputs(47)) or (inputs(83)));
    layer0_outputs(3684) <= (inputs(143)) and (inputs(144));
    layer0_outputs(3685) <= (inputs(14)) and not (inputs(87));
    layer0_outputs(3686) <= inputs(27);
    layer0_outputs(3687) <= inputs(192);
    layer0_outputs(3688) <= inputs(51);
    layer0_outputs(3689) <= not(inputs(132));
    layer0_outputs(3690) <= (inputs(238)) and not (inputs(4));
    layer0_outputs(3691) <= not(inputs(223)) or (inputs(142));
    layer0_outputs(3692) <= (inputs(35)) and not (inputs(128));
    layer0_outputs(3693) <= not(inputs(75));
    layer0_outputs(3694) <= not((inputs(120)) or (inputs(89)));
    layer0_outputs(3695) <= '1';
    layer0_outputs(3696) <= (inputs(225)) and not (inputs(95));
    layer0_outputs(3697) <= (inputs(244)) or (inputs(193));
    layer0_outputs(3698) <= inputs(68);
    layer0_outputs(3699) <= not(inputs(173)) or (inputs(65));
    layer0_outputs(3700) <= '0';
    layer0_outputs(3701) <= (inputs(175)) and not (inputs(229));
    layer0_outputs(3702) <= '0';
    layer0_outputs(3703) <= not(inputs(105)) or (inputs(84));
    layer0_outputs(3704) <= (inputs(19)) and not (inputs(252));
    layer0_outputs(3705) <= '1';
    layer0_outputs(3706) <= '1';
    layer0_outputs(3707) <= not(inputs(251));
    layer0_outputs(3708) <= (inputs(98)) and not (inputs(235));
    layer0_outputs(3709) <= not((inputs(164)) or (inputs(222)));
    layer0_outputs(3710) <= not((inputs(158)) xor (inputs(163)));
    layer0_outputs(3711) <= inputs(208);
    layer0_outputs(3712) <= not(inputs(141));
    layer0_outputs(3713) <= (inputs(16)) or (inputs(178));
    layer0_outputs(3714) <= inputs(85);
    layer0_outputs(3715) <= (inputs(237)) and (inputs(202));
    layer0_outputs(3716) <= not((inputs(195)) or (inputs(199)));
    layer0_outputs(3717) <= not(inputs(93)) or (inputs(193));
    layer0_outputs(3718) <= not((inputs(252)) xor (inputs(188)));
    layer0_outputs(3719) <= not(inputs(184)) or (inputs(142));
    layer0_outputs(3720) <= '0';
    layer0_outputs(3721) <= inputs(169);
    layer0_outputs(3722) <= '0';
    layer0_outputs(3723) <= not(inputs(29));
    layer0_outputs(3724) <= not(inputs(110)) or (inputs(238));
    layer0_outputs(3725) <= not(inputs(130));
    layer0_outputs(3726) <= '1';
    layer0_outputs(3727) <= inputs(99);
    layer0_outputs(3728) <= inputs(98);
    layer0_outputs(3729) <= not(inputs(232));
    layer0_outputs(3730) <= not(inputs(20));
    layer0_outputs(3731) <= (inputs(171)) and not (inputs(58));
    layer0_outputs(3732) <= (inputs(176)) or (inputs(169));
    layer0_outputs(3733) <= not(inputs(135));
    layer0_outputs(3734) <= inputs(18);
    layer0_outputs(3735) <= (inputs(222)) or (inputs(219));
    layer0_outputs(3736) <= '1';
    layer0_outputs(3737) <= not((inputs(157)) and (inputs(145)));
    layer0_outputs(3738) <= not((inputs(160)) xor (inputs(208)));
    layer0_outputs(3739) <= not((inputs(215)) or (inputs(249)));
    layer0_outputs(3740) <= not((inputs(3)) and (inputs(45)));
    layer0_outputs(3741) <= not((inputs(162)) or (inputs(242)));
    layer0_outputs(3742) <= not((inputs(45)) or (inputs(35)));
    layer0_outputs(3743) <= not(inputs(254));
    layer0_outputs(3744) <= inputs(249);
    layer0_outputs(3745) <= not((inputs(240)) or (inputs(80)));
    layer0_outputs(3746) <= not(inputs(242));
    layer0_outputs(3747) <= not(inputs(36));
    layer0_outputs(3748) <= not(inputs(112)) or (inputs(218));
    layer0_outputs(3749) <= '1';
    layer0_outputs(3750) <= '0';
    layer0_outputs(3751) <= not(inputs(97));
    layer0_outputs(3752) <= not((inputs(219)) xor (inputs(253)));
    layer0_outputs(3753) <= inputs(135);
    layer0_outputs(3754) <= '0';
    layer0_outputs(3755) <= '1';
    layer0_outputs(3756) <= (inputs(30)) and not (inputs(249));
    layer0_outputs(3757) <= inputs(235);
    layer0_outputs(3758) <= inputs(20);
    layer0_outputs(3759) <= (inputs(26)) and not (inputs(178));
    layer0_outputs(3760) <= not(inputs(160));
    layer0_outputs(3761) <= not(inputs(224)) or (inputs(205));
    layer0_outputs(3762) <= not((inputs(234)) xor (inputs(174)));
    layer0_outputs(3763) <= not(inputs(128)) or (inputs(159));
    layer0_outputs(3764) <= not((inputs(230)) and (inputs(116)));
    layer0_outputs(3765) <= inputs(116);
    layer0_outputs(3766) <= '0';
    layer0_outputs(3767) <= not((inputs(123)) and (inputs(217)));
    layer0_outputs(3768) <= inputs(49);
    layer0_outputs(3769) <= '1';
    layer0_outputs(3770) <= '1';
    layer0_outputs(3771) <= not(inputs(226));
    layer0_outputs(3772) <= '1';
    layer0_outputs(3773) <= '0';
    layer0_outputs(3774) <= (inputs(0)) and not (inputs(226));
    layer0_outputs(3775) <= inputs(23);
    layer0_outputs(3776) <= not(inputs(81)) or (inputs(50));
    layer0_outputs(3777) <= inputs(209);
    layer0_outputs(3778) <= inputs(26);
    layer0_outputs(3779) <= '0';
    layer0_outputs(3780) <= (inputs(17)) and not (inputs(81));
    layer0_outputs(3781) <= not((inputs(223)) or (inputs(64)));
    layer0_outputs(3782) <= not(inputs(41)) or (inputs(31));
    layer0_outputs(3783) <= (inputs(152)) or (inputs(100));
    layer0_outputs(3784) <= (inputs(139)) or (inputs(31));
    layer0_outputs(3785) <= inputs(253);
    layer0_outputs(3786) <= (inputs(151)) and not (inputs(106));
    layer0_outputs(3787) <= '0';
    layer0_outputs(3788) <= not(inputs(97)) or (inputs(155));
    layer0_outputs(3789) <= '1';
    layer0_outputs(3790) <= (inputs(27)) xor (inputs(71));
    layer0_outputs(3791) <= not(inputs(131));
    layer0_outputs(3792) <= not((inputs(91)) or (inputs(69)));
    layer0_outputs(3793) <= not((inputs(182)) or (inputs(17)));
    layer0_outputs(3794) <= not(inputs(174));
    layer0_outputs(3795) <= '1';
    layer0_outputs(3796) <= not(inputs(86)) or (inputs(70));
    layer0_outputs(3797) <= (inputs(133)) and not (inputs(200));
    layer0_outputs(3798) <= (inputs(138)) and not (inputs(208));
    layer0_outputs(3799) <= (inputs(160)) and not (inputs(145));
    layer0_outputs(3800) <= not((inputs(34)) or (inputs(191)));
    layer0_outputs(3801) <= (inputs(180)) xor (inputs(128));
    layer0_outputs(3802) <= inputs(68);
    layer0_outputs(3803) <= not(inputs(103));
    layer0_outputs(3804) <= inputs(230);
    layer0_outputs(3805) <= '1';
    layer0_outputs(3806) <= not(inputs(71)) or (inputs(211));
    layer0_outputs(3807) <= inputs(104);
    layer0_outputs(3808) <= '0';
    layer0_outputs(3809) <= (inputs(231)) and not (inputs(121));
    layer0_outputs(3810) <= not(inputs(22)) or (inputs(144));
    layer0_outputs(3811) <= '1';
    layer0_outputs(3812) <= not((inputs(183)) and (inputs(153)));
    layer0_outputs(3813) <= not(inputs(184)) or (inputs(215));
    layer0_outputs(3814) <= '1';
    layer0_outputs(3815) <= '0';
    layer0_outputs(3816) <= not((inputs(80)) and (inputs(6)));
    layer0_outputs(3817) <= (inputs(219)) or (inputs(36));
    layer0_outputs(3818) <= not((inputs(30)) or (inputs(169)));
    layer0_outputs(3819) <= not(inputs(189)) or (inputs(103));
    layer0_outputs(3820) <= inputs(84);
    layer0_outputs(3821) <= not((inputs(225)) or (inputs(229)));
    layer0_outputs(3822) <= not(inputs(145));
    layer0_outputs(3823) <= not(inputs(143));
    layer0_outputs(3824) <= (inputs(172)) and not (inputs(65));
    layer0_outputs(3825) <= (inputs(255)) and (inputs(250));
    layer0_outputs(3826) <= (inputs(219)) or (inputs(162));
    layer0_outputs(3827) <= '0';
    layer0_outputs(3828) <= not(inputs(182));
    layer0_outputs(3829) <= not(inputs(121)) or (inputs(195));
    layer0_outputs(3830) <= (inputs(147)) and (inputs(5));
    layer0_outputs(3831) <= '0';
    layer0_outputs(3832) <= not(inputs(148)) or (inputs(196));
    layer0_outputs(3833) <= '0';
    layer0_outputs(3834) <= (inputs(176)) and not (inputs(176));
    layer0_outputs(3835) <= not(inputs(160));
    layer0_outputs(3836) <= inputs(67);
    layer0_outputs(3837) <= '1';
    layer0_outputs(3838) <= not(inputs(17));
    layer0_outputs(3839) <= (inputs(223)) and not (inputs(187));
    layer0_outputs(3840) <= not((inputs(154)) or (inputs(153)));
    layer0_outputs(3841) <= not(inputs(48)) or (inputs(188));
    layer0_outputs(3842) <= inputs(87);
    layer0_outputs(3843) <= not(inputs(21)) or (inputs(84));
    layer0_outputs(3844) <= inputs(193);
    layer0_outputs(3845) <= (inputs(149)) and not (inputs(221));
    layer0_outputs(3846) <= (inputs(152)) and (inputs(152));
    layer0_outputs(3847) <= (inputs(4)) and not (inputs(114));
    layer0_outputs(3848) <= inputs(179);
    layer0_outputs(3849) <= not(inputs(89));
    layer0_outputs(3850) <= not(inputs(211));
    layer0_outputs(3851) <= not((inputs(1)) or (inputs(2)));
    layer0_outputs(3852) <= inputs(222);
    layer0_outputs(3853) <= inputs(90);
    layer0_outputs(3854) <= inputs(222);
    layer0_outputs(3855) <= not((inputs(246)) or (inputs(22)));
    layer0_outputs(3856) <= not(inputs(136));
    layer0_outputs(3857) <= not((inputs(84)) or (inputs(186)));
    layer0_outputs(3858) <= inputs(211);
    layer0_outputs(3859) <= inputs(106);
    layer0_outputs(3860) <= '1';
    layer0_outputs(3861) <= (inputs(159)) or (inputs(190));
    layer0_outputs(3862) <= not(inputs(26));
    layer0_outputs(3863) <= '1';
    layer0_outputs(3864) <= '1';
    layer0_outputs(3865) <= inputs(25);
    layer0_outputs(3866) <= not(inputs(197));
    layer0_outputs(3867) <= inputs(152);
    layer0_outputs(3868) <= not(inputs(130));
    layer0_outputs(3869) <= (inputs(3)) xor (inputs(18));
    layer0_outputs(3870) <= not((inputs(205)) or (inputs(220)));
    layer0_outputs(3871) <= not(inputs(18));
    layer0_outputs(3872) <= '1';
    layer0_outputs(3873) <= not((inputs(145)) or (inputs(39)));
    layer0_outputs(3874) <= (inputs(226)) or (inputs(60));
    layer0_outputs(3875) <= not(inputs(105));
    layer0_outputs(3876) <= not((inputs(202)) or (inputs(49)));
    layer0_outputs(3877) <= inputs(42);
    layer0_outputs(3878) <= not(inputs(211)) or (inputs(240));
    layer0_outputs(3879) <= (inputs(238)) or (inputs(31));
    layer0_outputs(3880) <= inputs(236);
    layer0_outputs(3881) <= '1';
    layer0_outputs(3882) <= not(inputs(94)) or (inputs(26));
    layer0_outputs(3883) <= (inputs(126)) or (inputs(105));
    layer0_outputs(3884) <= (inputs(186)) xor (inputs(29));
    layer0_outputs(3885) <= '0';
    layer0_outputs(3886) <= '0';
    layer0_outputs(3887) <= '1';
    layer0_outputs(3888) <= not(inputs(42));
    layer0_outputs(3889) <= not(inputs(141));
    layer0_outputs(3890) <= inputs(138);
    layer0_outputs(3891) <= not(inputs(178));
    layer0_outputs(3892) <= '1';
    layer0_outputs(3893) <= not(inputs(115));
    layer0_outputs(3894) <= not(inputs(177));
    layer0_outputs(3895) <= '1';
    layer0_outputs(3896) <= inputs(167);
    layer0_outputs(3897) <= not(inputs(167));
    layer0_outputs(3898) <= (inputs(202)) or (inputs(238));
    layer0_outputs(3899) <= (inputs(153)) or (inputs(9));
    layer0_outputs(3900) <= not((inputs(27)) or (inputs(106)));
    layer0_outputs(3901) <= (inputs(64)) and not (inputs(36));
    layer0_outputs(3902) <= not(inputs(147));
    layer0_outputs(3903) <= not(inputs(152));
    layer0_outputs(3904) <= not(inputs(181)) or (inputs(30));
    layer0_outputs(3905) <= '1';
    layer0_outputs(3906) <= not(inputs(81));
    layer0_outputs(3907) <= inputs(19);
    layer0_outputs(3908) <= inputs(191);
    layer0_outputs(3909) <= not(inputs(228)) or (inputs(98));
    layer0_outputs(3910) <= inputs(68);
    layer0_outputs(3911) <= (inputs(69)) or (inputs(128));
    layer0_outputs(3912) <= not(inputs(204)) or (inputs(65));
    layer0_outputs(3913) <= '0';
    layer0_outputs(3914) <= inputs(17);
    layer0_outputs(3915) <= not(inputs(90)) or (inputs(218));
    layer0_outputs(3916) <= inputs(69);
    layer0_outputs(3917) <= '1';
    layer0_outputs(3918) <= inputs(85);
    layer0_outputs(3919) <= not(inputs(40)) or (inputs(67));
    layer0_outputs(3920) <= inputs(40);
    layer0_outputs(3921) <= not((inputs(188)) or (inputs(209)));
    layer0_outputs(3922) <= (inputs(180)) xor (inputs(209));
    layer0_outputs(3923) <= inputs(172);
    layer0_outputs(3924) <= not(inputs(153)) or (inputs(10));
    layer0_outputs(3925) <= not(inputs(166));
    layer0_outputs(3926) <= (inputs(241)) or (inputs(125));
    layer0_outputs(3927) <= (inputs(137)) and not (inputs(70));
    layer0_outputs(3928) <= '1';
    layer0_outputs(3929) <= not(inputs(222)) or (inputs(200));
    layer0_outputs(3930) <= not((inputs(164)) xor (inputs(126)));
    layer0_outputs(3931) <= (inputs(198)) and not (inputs(100));
    layer0_outputs(3932) <= not((inputs(50)) and (inputs(86)));
    layer0_outputs(3933) <= inputs(159);
    layer0_outputs(3934) <= '0';
    layer0_outputs(3935) <= '0';
    layer0_outputs(3936) <= inputs(230);
    layer0_outputs(3937) <= inputs(72);
    layer0_outputs(3938) <= not((inputs(222)) or (inputs(203)));
    layer0_outputs(3939) <= '1';
    layer0_outputs(3940) <= not(inputs(194)) or (inputs(18));
    layer0_outputs(3941) <= inputs(255);
    layer0_outputs(3942) <= inputs(168);
    layer0_outputs(3943) <= not((inputs(169)) or (inputs(236)));
    layer0_outputs(3944) <= not(inputs(60)) or (inputs(55));
    layer0_outputs(3945) <= not((inputs(255)) xor (inputs(56)));
    layer0_outputs(3946) <= not(inputs(68)) or (inputs(149));
    layer0_outputs(3947) <= inputs(163);
    layer0_outputs(3948) <= (inputs(205)) or (inputs(178));
    layer0_outputs(3949) <= (inputs(222)) and (inputs(144));
    layer0_outputs(3950) <= not(inputs(23)) or (inputs(45));
    layer0_outputs(3951) <= not((inputs(242)) or (inputs(196)));
    layer0_outputs(3952) <= not(inputs(153)) or (inputs(55));
    layer0_outputs(3953) <= inputs(67);
    layer0_outputs(3954) <= (inputs(12)) and not (inputs(251));
    layer0_outputs(3955) <= inputs(225);
    layer0_outputs(3956) <= (inputs(115)) or (inputs(113));
    layer0_outputs(3957) <= (inputs(157)) and (inputs(72));
    layer0_outputs(3958) <= not(inputs(63));
    layer0_outputs(3959) <= (inputs(250)) and not (inputs(119));
    layer0_outputs(3960) <= (inputs(120)) and not (inputs(35));
    layer0_outputs(3961) <= inputs(182);
    layer0_outputs(3962) <= '1';
    layer0_outputs(3963) <= not((inputs(215)) and (inputs(79)));
    layer0_outputs(3964) <= not((inputs(11)) xor (inputs(50)));
    layer0_outputs(3965) <= '0';
    layer0_outputs(3966) <= (inputs(195)) and not (inputs(113));
    layer0_outputs(3967) <= not(inputs(110));
    layer0_outputs(3968) <= (inputs(69)) or (inputs(200));
    layer0_outputs(3969) <= inputs(230);
    layer0_outputs(3970) <= not((inputs(176)) xor (inputs(180)));
    layer0_outputs(3971) <= '1';
    layer0_outputs(3972) <= inputs(197);
    layer0_outputs(3973) <= inputs(237);
    layer0_outputs(3974) <= not(inputs(120));
    layer0_outputs(3975) <= (inputs(222)) or (inputs(232));
    layer0_outputs(3976) <= (inputs(128)) and (inputs(161));
    layer0_outputs(3977) <= (inputs(112)) and (inputs(81));
    layer0_outputs(3978) <= not(inputs(30)) or (inputs(105));
    layer0_outputs(3979) <= not(inputs(86)) or (inputs(74));
    layer0_outputs(3980) <= (inputs(3)) and not (inputs(153));
    layer0_outputs(3981) <= inputs(83);
    layer0_outputs(3982) <= not(inputs(255));
    layer0_outputs(3983) <= not(inputs(39));
    layer0_outputs(3984) <= (inputs(148)) and not (inputs(238));
    layer0_outputs(3985) <= '1';
    layer0_outputs(3986) <= (inputs(60)) or (inputs(48));
    layer0_outputs(3987) <= (inputs(250)) and (inputs(61));
    layer0_outputs(3988) <= inputs(86);
    layer0_outputs(3989) <= not((inputs(36)) or (inputs(10)));
    layer0_outputs(3990) <= inputs(223);
    layer0_outputs(3991) <= not(inputs(55));
    layer0_outputs(3992) <= '0';
    layer0_outputs(3993) <= inputs(130);
    layer0_outputs(3994) <= not((inputs(9)) or (inputs(140)));
    layer0_outputs(3995) <= not(inputs(132)) or (inputs(163));
    layer0_outputs(3996) <= (inputs(176)) and not (inputs(75));
    layer0_outputs(3997) <= (inputs(119)) or (inputs(253));
    layer0_outputs(3998) <= '1';
    layer0_outputs(3999) <= (inputs(9)) and not (inputs(210));
    layer0_outputs(4000) <= not((inputs(162)) xor (inputs(88)));
    layer0_outputs(4001) <= '0';
    layer0_outputs(4002) <= not((inputs(10)) or (inputs(25)));
    layer0_outputs(4003) <= (inputs(77)) and (inputs(118));
    layer0_outputs(4004) <= inputs(190);
    layer0_outputs(4005) <= (inputs(208)) and not (inputs(126));
    layer0_outputs(4006) <= '1';
    layer0_outputs(4007) <= inputs(91);
    layer0_outputs(4008) <= not(inputs(133));
    layer0_outputs(4009) <= '1';
    layer0_outputs(4010) <= (inputs(146)) or (inputs(83));
    layer0_outputs(4011) <= inputs(238);
    layer0_outputs(4012) <= not(inputs(88)) or (inputs(221));
    layer0_outputs(4013) <= not(inputs(35));
    layer0_outputs(4014) <= (inputs(54)) and (inputs(176));
    layer0_outputs(4015) <= (inputs(177)) and (inputs(84));
    layer0_outputs(4016) <= not((inputs(97)) and (inputs(222)));
    layer0_outputs(4017) <= (inputs(27)) and (inputs(39));
    layer0_outputs(4018) <= (inputs(198)) or (inputs(222));
    layer0_outputs(4019) <= '1';
    layer0_outputs(4020) <= (inputs(0)) or (inputs(43));
    layer0_outputs(4021) <= (inputs(144)) and not (inputs(240));
    layer0_outputs(4022) <= not(inputs(2));
    layer0_outputs(4023) <= inputs(122);
    layer0_outputs(4024) <= not((inputs(4)) or (inputs(109)));
    layer0_outputs(4025) <= inputs(36);
    layer0_outputs(4026) <= (inputs(211)) or (inputs(147));
    layer0_outputs(4027) <= not((inputs(80)) or (inputs(137)));
    layer0_outputs(4028) <= inputs(210);
    layer0_outputs(4029) <= '1';
    layer0_outputs(4030) <= '0';
    layer0_outputs(4031) <= not(inputs(104));
    layer0_outputs(4032) <= '0';
    layer0_outputs(4033) <= inputs(27);
    layer0_outputs(4034) <= (inputs(167)) xor (inputs(166));
    layer0_outputs(4035) <= (inputs(250)) and (inputs(66));
    layer0_outputs(4036) <= '0';
    layer0_outputs(4037) <= not(inputs(209));
    layer0_outputs(4038) <= '0';
    layer0_outputs(4039) <= not((inputs(176)) xor (inputs(3)));
    layer0_outputs(4040) <= inputs(211);
    layer0_outputs(4041) <= inputs(40);
    layer0_outputs(4042) <= not(inputs(105));
    layer0_outputs(4043) <= inputs(185);
    layer0_outputs(4044) <= (inputs(237)) and (inputs(176));
    layer0_outputs(4045) <= not(inputs(194));
    layer0_outputs(4046) <= (inputs(52)) and not (inputs(228));
    layer0_outputs(4047) <= (inputs(228)) and (inputs(112));
    layer0_outputs(4048) <= (inputs(251)) and not (inputs(233));
    layer0_outputs(4049) <= not((inputs(137)) and (inputs(201)));
    layer0_outputs(4050) <= (inputs(3)) xor (inputs(85));
    layer0_outputs(4051) <= inputs(166);
    layer0_outputs(4052) <= not(inputs(89)) or (inputs(174));
    layer0_outputs(4053) <= (inputs(56)) or (inputs(22));
    layer0_outputs(4054) <= inputs(157);
    layer0_outputs(4055) <= (inputs(135)) or (inputs(46));
    layer0_outputs(4056) <= '1';
    layer0_outputs(4057) <= inputs(25);
    layer0_outputs(4058) <= '0';
    layer0_outputs(4059) <= not(inputs(253)) or (inputs(241));
    layer0_outputs(4060) <= not((inputs(113)) or (inputs(11)));
    layer0_outputs(4061) <= not((inputs(49)) or (inputs(156)));
    layer0_outputs(4062) <= not((inputs(24)) or (inputs(196)));
    layer0_outputs(4063) <= (inputs(180)) or (inputs(8));
    layer0_outputs(4064) <= not(inputs(70)) or (inputs(220));
    layer0_outputs(4065) <= not((inputs(46)) or (inputs(144)));
    layer0_outputs(4066) <= not((inputs(19)) and (inputs(93)));
    layer0_outputs(4067) <= '1';
    layer0_outputs(4068) <= not(inputs(122)) or (inputs(196));
    layer0_outputs(4069) <= (inputs(220)) or (inputs(129));
    layer0_outputs(4070) <= not((inputs(20)) and (inputs(217)));
    layer0_outputs(4071) <= not(inputs(84)) or (inputs(220));
    layer0_outputs(4072) <= (inputs(39)) and not (inputs(110));
    layer0_outputs(4073) <= not(inputs(157));
    layer0_outputs(4074) <= not(inputs(233)) or (inputs(236));
    layer0_outputs(4075) <= not(inputs(91)) or (inputs(169));
    layer0_outputs(4076) <= not(inputs(193));
    layer0_outputs(4077) <= (inputs(195)) or (inputs(167));
    layer0_outputs(4078) <= (inputs(125)) or (inputs(8));
    layer0_outputs(4079) <= not(inputs(67)) or (inputs(115));
    layer0_outputs(4080) <= '0';
    layer0_outputs(4081) <= (inputs(104)) and not (inputs(242));
    layer0_outputs(4082) <= (inputs(225)) or (inputs(169));
    layer0_outputs(4083) <= (inputs(1)) and (inputs(63));
    layer0_outputs(4084) <= inputs(66);
    layer0_outputs(4085) <= (inputs(53)) and not (inputs(92));
    layer0_outputs(4086) <= (inputs(183)) and not (inputs(94));
    layer0_outputs(4087) <= '0';
    layer0_outputs(4088) <= (inputs(178)) or (inputs(177));
    layer0_outputs(4089) <= not((inputs(198)) or (inputs(149)));
    layer0_outputs(4090) <= not(inputs(235));
    layer0_outputs(4091) <= '0';
    layer0_outputs(4092) <= (inputs(191)) or (inputs(211));
    layer0_outputs(4093) <= '0';
    layer0_outputs(4094) <= (inputs(235)) and not (inputs(116));
    layer0_outputs(4095) <= '0';
    layer0_outputs(4096) <= inputs(99);
    layer0_outputs(4097) <= '1';
    layer0_outputs(4098) <= '1';
    layer0_outputs(4099) <= not((inputs(33)) xor (inputs(249)));
    layer0_outputs(4100) <= (inputs(115)) and not (inputs(72));
    layer0_outputs(4101) <= not(inputs(224));
    layer0_outputs(4102) <= not(inputs(147));
    layer0_outputs(4103) <= not((inputs(84)) or (inputs(209)));
    layer0_outputs(4104) <= '1';
    layer0_outputs(4105) <= (inputs(210)) and not (inputs(46));
    layer0_outputs(4106) <= not(inputs(92));
    layer0_outputs(4107) <= not(inputs(50)) or (inputs(120));
    layer0_outputs(4108) <= not(inputs(231));
    layer0_outputs(4109) <= (inputs(11)) and (inputs(177));
    layer0_outputs(4110) <= '0';
    layer0_outputs(4111) <= not((inputs(69)) or (inputs(68)));
    layer0_outputs(4112) <= not(inputs(215)) or (inputs(63));
    layer0_outputs(4113) <= inputs(102);
    layer0_outputs(4114) <= not(inputs(153));
    layer0_outputs(4115) <= inputs(98);
    layer0_outputs(4116) <= (inputs(101)) and not (inputs(143));
    layer0_outputs(4117) <= '0';
    layer0_outputs(4118) <= (inputs(220)) and not (inputs(226));
    layer0_outputs(4119) <= (inputs(102)) and not (inputs(109));
    layer0_outputs(4120) <= inputs(224);
    layer0_outputs(4121) <= (inputs(194)) or (inputs(212));
    layer0_outputs(4122) <= not((inputs(183)) or (inputs(57)));
    layer0_outputs(4123) <= '1';
    layer0_outputs(4124) <= not(inputs(120));
    layer0_outputs(4125) <= (inputs(54)) or (inputs(125));
    layer0_outputs(4126) <= inputs(123);
    layer0_outputs(4127) <= not(inputs(85)) or (inputs(101));
    layer0_outputs(4128) <= not(inputs(146)) or (inputs(171));
    layer0_outputs(4129) <= not((inputs(87)) and (inputs(90)));
    layer0_outputs(4130) <= (inputs(49)) and not (inputs(247));
    layer0_outputs(4131) <= not((inputs(96)) or (inputs(120)));
    layer0_outputs(4132) <= not(inputs(206));
    layer0_outputs(4133) <= not(inputs(35)) or (inputs(177));
    layer0_outputs(4134) <= (inputs(75)) and (inputs(31));
    layer0_outputs(4135) <= inputs(128);
    layer0_outputs(4136) <= inputs(209);
    layer0_outputs(4137) <= '1';
    layer0_outputs(4138) <= '0';
    layer0_outputs(4139) <= (inputs(110)) or (inputs(60));
    layer0_outputs(4140) <= (inputs(142)) and not (inputs(199));
    layer0_outputs(4141) <= (inputs(111)) xor (inputs(123));
    layer0_outputs(4142) <= not(inputs(58));
    layer0_outputs(4143) <= not((inputs(182)) and (inputs(195)));
    layer0_outputs(4144) <= not((inputs(229)) or (inputs(203)));
    layer0_outputs(4145) <= (inputs(50)) and not (inputs(67));
    layer0_outputs(4146) <= (inputs(130)) or (inputs(133));
    layer0_outputs(4147) <= '0';
    layer0_outputs(4148) <= not((inputs(105)) or (inputs(216)));
    layer0_outputs(4149) <= inputs(95);
    layer0_outputs(4150) <= (inputs(7)) and not (inputs(228));
    layer0_outputs(4151) <= not(inputs(137)) or (inputs(212));
    layer0_outputs(4152) <= (inputs(14)) and (inputs(117));
    layer0_outputs(4153) <= not((inputs(108)) and (inputs(10)));
    layer0_outputs(4154) <= (inputs(170)) and not (inputs(239));
    layer0_outputs(4155) <= not(inputs(245)) or (inputs(36));
    layer0_outputs(4156) <= '1';
    layer0_outputs(4157) <= not(inputs(125)) or (inputs(10));
    layer0_outputs(4158) <= (inputs(9)) and not (inputs(56));
    layer0_outputs(4159) <= not((inputs(67)) or (inputs(76)));
    layer0_outputs(4160) <= '0';
    layer0_outputs(4161) <= not(inputs(101));
    layer0_outputs(4162) <= not((inputs(128)) or (inputs(134)));
    layer0_outputs(4163) <= '1';
    layer0_outputs(4164) <= inputs(76);
    layer0_outputs(4165) <= (inputs(38)) and not (inputs(152));
    layer0_outputs(4166) <= '0';
    layer0_outputs(4167) <= '0';
    layer0_outputs(4168) <= not(inputs(208));
    layer0_outputs(4169) <= (inputs(25)) and not (inputs(126));
    layer0_outputs(4170) <= (inputs(158)) and not (inputs(178));
    layer0_outputs(4171) <= not(inputs(98));
    layer0_outputs(4172) <= not(inputs(84)) or (inputs(207));
    layer0_outputs(4173) <= not(inputs(129)) or (inputs(209));
    layer0_outputs(4174) <= (inputs(165)) and not (inputs(5));
    layer0_outputs(4175) <= not(inputs(233)) or (inputs(34));
    layer0_outputs(4176) <= inputs(110);
    layer0_outputs(4177) <= (inputs(94)) xor (inputs(197));
    layer0_outputs(4178) <= inputs(39);
    layer0_outputs(4179) <= '0';
    layer0_outputs(4180) <= (inputs(197)) and not (inputs(244));
    layer0_outputs(4181) <= not(inputs(162));
    layer0_outputs(4182) <= (inputs(15)) or (inputs(56));
    layer0_outputs(4183) <= not((inputs(204)) or (inputs(165)));
    layer0_outputs(4184) <= '1';
    layer0_outputs(4185) <= not(inputs(42));
    layer0_outputs(4186) <= not(inputs(43)) or (inputs(102));
    layer0_outputs(4187) <= '0';
    layer0_outputs(4188) <= inputs(39);
    layer0_outputs(4189) <= (inputs(155)) and not (inputs(57));
    layer0_outputs(4190) <= not(inputs(71));
    layer0_outputs(4191) <= '0';
    layer0_outputs(4192) <= (inputs(18)) xor (inputs(45));
    layer0_outputs(4193) <= not((inputs(106)) or (inputs(254)));
    layer0_outputs(4194) <= not((inputs(1)) xor (inputs(249)));
    layer0_outputs(4195) <= not((inputs(246)) and (inputs(91)));
    layer0_outputs(4196) <= (inputs(93)) or (inputs(167));
    layer0_outputs(4197) <= not((inputs(252)) or (inputs(141)));
    layer0_outputs(4198) <= not((inputs(100)) or (inputs(81)));
    layer0_outputs(4199) <= (inputs(7)) or (inputs(230));
    layer0_outputs(4200) <= not((inputs(81)) and (inputs(149)));
    layer0_outputs(4201) <= inputs(233);
    layer0_outputs(4202) <= inputs(41);
    layer0_outputs(4203) <= inputs(66);
    layer0_outputs(4204) <= inputs(103);
    layer0_outputs(4205) <= inputs(5);
    layer0_outputs(4206) <= inputs(8);
    layer0_outputs(4207) <= not(inputs(94)) or (inputs(186));
    layer0_outputs(4208) <= not((inputs(94)) xor (inputs(48)));
    layer0_outputs(4209) <= '0';
    layer0_outputs(4210) <= not((inputs(197)) or (inputs(119)));
    layer0_outputs(4211) <= (inputs(27)) and not (inputs(40));
    layer0_outputs(4212) <= (inputs(169)) and not (inputs(58));
    layer0_outputs(4213) <= not((inputs(98)) or (inputs(100)));
    layer0_outputs(4214) <= '1';
    layer0_outputs(4215) <= inputs(96);
    layer0_outputs(4216) <= '0';
    layer0_outputs(4217) <= inputs(97);
    layer0_outputs(4218) <= (inputs(137)) and not (inputs(90));
    layer0_outputs(4219) <= (inputs(156)) and not (inputs(159));
    layer0_outputs(4220) <= not(inputs(206)) or (inputs(9));
    layer0_outputs(4221) <= not((inputs(158)) and (inputs(174)));
    layer0_outputs(4222) <= not(inputs(145));
    layer0_outputs(4223) <= not(inputs(162));
    layer0_outputs(4224) <= (inputs(88)) or (inputs(162));
    layer0_outputs(4225) <= (inputs(62)) xor (inputs(142));
    layer0_outputs(4226) <= (inputs(10)) and not (inputs(72));
    layer0_outputs(4227) <= (inputs(137)) and not (inputs(177));
    layer0_outputs(4228) <= not((inputs(107)) or (inputs(252)));
    layer0_outputs(4229) <= not((inputs(78)) xor (inputs(131)));
    layer0_outputs(4230) <= (inputs(225)) or (inputs(212));
    layer0_outputs(4231) <= not(inputs(40));
    layer0_outputs(4232) <= not((inputs(187)) or (inputs(226)));
    layer0_outputs(4233) <= inputs(112);
    layer0_outputs(4234) <= not((inputs(105)) or (inputs(158)));
    layer0_outputs(4235) <= inputs(83);
    layer0_outputs(4236) <= inputs(82);
    layer0_outputs(4237) <= (inputs(66)) and not (inputs(249));
    layer0_outputs(4238) <= (inputs(148)) and not (inputs(223));
    layer0_outputs(4239) <= (inputs(21)) and not (inputs(214));
    layer0_outputs(4240) <= inputs(81);
    layer0_outputs(4241) <= not(inputs(230)) or (inputs(88));
    layer0_outputs(4242) <= (inputs(99)) or (inputs(247));
    layer0_outputs(4243) <= not((inputs(149)) and (inputs(204)));
    layer0_outputs(4244) <= '1';
    layer0_outputs(4245) <= not((inputs(36)) xor (inputs(125)));
    layer0_outputs(4246) <= (inputs(75)) or (inputs(75));
    layer0_outputs(4247) <= not(inputs(245));
    layer0_outputs(4248) <= not(inputs(154));
    layer0_outputs(4249) <= (inputs(89)) and not (inputs(191));
    layer0_outputs(4250) <= not(inputs(118));
    layer0_outputs(4251) <= not((inputs(130)) xor (inputs(152)));
    layer0_outputs(4252) <= '0';
    layer0_outputs(4253) <= not(inputs(122));
    layer0_outputs(4254) <= not((inputs(237)) or (inputs(221)));
    layer0_outputs(4255) <= (inputs(115)) and not (inputs(53));
    layer0_outputs(4256) <= inputs(230);
    layer0_outputs(4257) <= not((inputs(91)) xor (inputs(212)));
    layer0_outputs(4258) <= not(inputs(211)) or (inputs(176));
    layer0_outputs(4259) <= (inputs(81)) xor (inputs(34));
    layer0_outputs(4260) <= not((inputs(68)) or (inputs(129)));
    layer0_outputs(4261) <= (inputs(0)) and not (inputs(1));
    layer0_outputs(4262) <= not(inputs(146));
    layer0_outputs(4263) <= '0';
    layer0_outputs(4264) <= '0';
    layer0_outputs(4265) <= not(inputs(166));
    layer0_outputs(4266) <= inputs(26);
    layer0_outputs(4267) <= inputs(248);
    layer0_outputs(4268) <= not((inputs(178)) or (inputs(182)));
    layer0_outputs(4269) <= not(inputs(180));
    layer0_outputs(4270) <= not(inputs(22));
    layer0_outputs(4271) <= not((inputs(181)) or (inputs(183)));
    layer0_outputs(4272) <= not((inputs(77)) or (inputs(108)));
    layer0_outputs(4273) <= (inputs(245)) or (inputs(230));
    layer0_outputs(4274) <= not((inputs(50)) or (inputs(132)));
    layer0_outputs(4275) <= (inputs(206)) and not (inputs(80));
    layer0_outputs(4276) <= '0';
    layer0_outputs(4277) <= inputs(238);
    layer0_outputs(4278) <= inputs(234);
    layer0_outputs(4279) <= (inputs(66)) xor (inputs(199));
    layer0_outputs(4280) <= not((inputs(202)) and (inputs(90)));
    layer0_outputs(4281) <= not((inputs(254)) or (inputs(193)));
    layer0_outputs(4282) <= not(inputs(129));
    layer0_outputs(4283) <= not((inputs(109)) xor (inputs(228)));
    layer0_outputs(4284) <= not((inputs(131)) xor (inputs(222)));
    layer0_outputs(4285) <= not(inputs(108));
    layer0_outputs(4286) <= not(inputs(156)) or (inputs(201));
    layer0_outputs(4287) <= (inputs(2)) or (inputs(47));
    layer0_outputs(4288) <= (inputs(35)) and not (inputs(75));
    layer0_outputs(4289) <= (inputs(51)) and not (inputs(246));
    layer0_outputs(4290) <= not(inputs(107));
    layer0_outputs(4291) <= inputs(254);
    layer0_outputs(4292) <= '0';
    layer0_outputs(4293) <= not((inputs(29)) or (inputs(51)));
    layer0_outputs(4294) <= (inputs(139)) and not (inputs(72));
    layer0_outputs(4295) <= not(inputs(94)) or (inputs(176));
    layer0_outputs(4296) <= not((inputs(107)) xor (inputs(183)));
    layer0_outputs(4297) <= inputs(46);
    layer0_outputs(4298) <= '0';
    layer0_outputs(4299) <= '0';
    layer0_outputs(4300) <= '0';
    layer0_outputs(4301) <= (inputs(30)) and not (inputs(167));
    layer0_outputs(4302) <= not(inputs(107));
    layer0_outputs(4303) <= not(inputs(109)) or (inputs(51));
    layer0_outputs(4304) <= (inputs(215)) xor (inputs(130));
    layer0_outputs(4305) <= (inputs(196)) or (inputs(172));
    layer0_outputs(4306) <= not(inputs(59)) or (inputs(175));
    layer0_outputs(4307) <= inputs(80);
    layer0_outputs(4308) <= not(inputs(45));
    layer0_outputs(4309) <= not(inputs(48)) or (inputs(206));
    layer0_outputs(4310) <= (inputs(5)) and (inputs(99));
    layer0_outputs(4311) <= (inputs(62)) and not (inputs(108));
    layer0_outputs(4312) <= (inputs(178)) or (inputs(188));
    layer0_outputs(4313) <= not(inputs(179));
    layer0_outputs(4314) <= '0';
    layer0_outputs(4315) <= inputs(199);
    layer0_outputs(4316) <= (inputs(103)) or (inputs(109));
    layer0_outputs(4317) <= inputs(255);
    layer0_outputs(4318) <= not(inputs(31)) or (inputs(6));
    layer0_outputs(4319) <= (inputs(159)) and not (inputs(65));
    layer0_outputs(4320) <= '0';
    layer0_outputs(4321) <= inputs(0);
    layer0_outputs(4322) <= not(inputs(211)) or (inputs(28));
    layer0_outputs(4323) <= inputs(117);
    layer0_outputs(4324) <= not(inputs(34));
    layer0_outputs(4325) <= inputs(134);
    layer0_outputs(4326) <= not(inputs(176));
    layer0_outputs(4327) <= not(inputs(239));
    layer0_outputs(4328) <= not(inputs(187));
    layer0_outputs(4329) <= (inputs(128)) and not (inputs(27));
    layer0_outputs(4330) <= inputs(167);
    layer0_outputs(4331) <= (inputs(234)) and not (inputs(193));
    layer0_outputs(4332) <= inputs(128);
    layer0_outputs(4333) <= (inputs(20)) xor (inputs(239));
    layer0_outputs(4334) <= inputs(65);
    layer0_outputs(4335) <= not(inputs(4)) or (inputs(84));
    layer0_outputs(4336) <= not((inputs(250)) xor (inputs(21)));
    layer0_outputs(4337) <= not((inputs(70)) or (inputs(148)));
    layer0_outputs(4338) <= not((inputs(72)) and (inputs(128)));
    layer0_outputs(4339) <= not(inputs(160)) or (inputs(221));
    layer0_outputs(4340) <= not(inputs(215)) or (inputs(16));
    layer0_outputs(4341) <= not(inputs(6));
    layer0_outputs(4342) <= '0';
    layer0_outputs(4343) <= (inputs(0)) or (inputs(77));
    layer0_outputs(4344) <= not(inputs(21));
    layer0_outputs(4345) <= '1';
    layer0_outputs(4346) <= inputs(119);
    layer0_outputs(4347) <= (inputs(196)) or (inputs(198));
    layer0_outputs(4348) <= inputs(209);
    layer0_outputs(4349) <= (inputs(40)) or (inputs(244));
    layer0_outputs(4350) <= inputs(29);
    layer0_outputs(4351) <= not(inputs(136));
    layer0_outputs(4352) <= not((inputs(24)) xor (inputs(69)));
    layer0_outputs(4353) <= (inputs(128)) and not (inputs(72));
    layer0_outputs(4354) <= not(inputs(211));
    layer0_outputs(4355) <= not((inputs(75)) or (inputs(7)));
    layer0_outputs(4356) <= (inputs(165)) or (inputs(110));
    layer0_outputs(4357) <= not(inputs(81)) or (inputs(107));
    layer0_outputs(4358) <= not((inputs(2)) and (inputs(245)));
    layer0_outputs(4359) <= not((inputs(127)) and (inputs(30)));
    layer0_outputs(4360) <= not(inputs(60)) or (inputs(83));
    layer0_outputs(4361) <= '1';
    layer0_outputs(4362) <= not(inputs(202));
    layer0_outputs(4363) <= not((inputs(132)) and (inputs(164)));
    layer0_outputs(4364) <= not(inputs(122));
    layer0_outputs(4365) <= (inputs(155)) xor (inputs(94));
    layer0_outputs(4366) <= not(inputs(43));
    layer0_outputs(4367) <= '1';
    layer0_outputs(4368) <= '1';
    layer0_outputs(4369) <= '0';
    layer0_outputs(4370) <= not(inputs(34));
    layer0_outputs(4371) <= '1';
    layer0_outputs(4372) <= inputs(163);
    layer0_outputs(4373) <= not((inputs(46)) or (inputs(20)));
    layer0_outputs(4374) <= (inputs(51)) and not (inputs(162));
    layer0_outputs(4375) <= (inputs(70)) and not (inputs(109));
    layer0_outputs(4376) <= (inputs(209)) and not (inputs(87));
    layer0_outputs(4377) <= not((inputs(144)) or (inputs(233)));
    layer0_outputs(4378) <= inputs(223);
    layer0_outputs(4379) <= not((inputs(147)) and (inputs(150)));
    layer0_outputs(4380) <= inputs(160);
    layer0_outputs(4381) <= inputs(12);
    layer0_outputs(4382) <= (inputs(231)) and (inputs(63));
    layer0_outputs(4383) <= (inputs(49)) and not (inputs(60));
    layer0_outputs(4384) <= (inputs(112)) or (inputs(67));
    layer0_outputs(4385) <= inputs(98);
    layer0_outputs(4386) <= not((inputs(38)) or (inputs(155)));
    layer0_outputs(4387) <= (inputs(109)) and not (inputs(44));
    layer0_outputs(4388) <= inputs(134);
    layer0_outputs(4389) <= (inputs(74)) and (inputs(25));
    layer0_outputs(4390) <= not((inputs(145)) or (inputs(124)));
    layer0_outputs(4391) <= inputs(11);
    layer0_outputs(4392) <= not((inputs(64)) xor (inputs(170)));
    layer0_outputs(4393) <= inputs(168);
    layer0_outputs(4394) <= not(inputs(139));
    layer0_outputs(4395) <= not(inputs(112));
    layer0_outputs(4396) <= inputs(213);
    layer0_outputs(4397) <= not(inputs(163));
    layer0_outputs(4398) <= not(inputs(39));
    layer0_outputs(4399) <= (inputs(232)) xor (inputs(92));
    layer0_outputs(4400) <= not(inputs(21));
    layer0_outputs(4401) <= '0';
    layer0_outputs(4402) <= not((inputs(73)) and (inputs(242)));
    layer0_outputs(4403) <= '0';
    layer0_outputs(4404) <= not((inputs(173)) or (inputs(100)));
    layer0_outputs(4405) <= not((inputs(183)) or (inputs(162)));
    layer0_outputs(4406) <= inputs(193);
    layer0_outputs(4407) <= not(inputs(88));
    layer0_outputs(4408) <= not(inputs(152));
    layer0_outputs(4409) <= not(inputs(248)) or (inputs(238));
    layer0_outputs(4410) <= not(inputs(174)) or (inputs(216));
    layer0_outputs(4411) <= '1';
    layer0_outputs(4412) <= inputs(89);
    layer0_outputs(4413) <= not(inputs(21));
    layer0_outputs(4414) <= not(inputs(85)) or (inputs(191));
    layer0_outputs(4415) <= not(inputs(189));
    layer0_outputs(4416) <= (inputs(230)) and not (inputs(72));
    layer0_outputs(4417) <= inputs(59);
    layer0_outputs(4418) <= not(inputs(246)) or (inputs(246));
    layer0_outputs(4419) <= '0';
    layer0_outputs(4420) <= (inputs(211)) xor (inputs(5));
    layer0_outputs(4421) <= inputs(170);
    layer0_outputs(4422) <= not(inputs(118));
    layer0_outputs(4423) <= not(inputs(151));
    layer0_outputs(4424) <= inputs(14);
    layer0_outputs(4425) <= not(inputs(235));
    layer0_outputs(4426) <= (inputs(155)) and not (inputs(185));
    layer0_outputs(4427) <= not(inputs(194));
    layer0_outputs(4428) <= inputs(164);
    layer0_outputs(4429) <= not((inputs(167)) and (inputs(35)));
    layer0_outputs(4430) <= (inputs(36)) and not (inputs(191));
    layer0_outputs(4431) <= inputs(207);
    layer0_outputs(4432) <= (inputs(157)) and not (inputs(246));
    layer0_outputs(4433) <= not((inputs(40)) or (inputs(9)));
    layer0_outputs(4434) <= '1';
    layer0_outputs(4435) <= not(inputs(34));
    layer0_outputs(4436) <= '0';
    layer0_outputs(4437) <= (inputs(108)) and not (inputs(254));
    layer0_outputs(4438) <= inputs(152);
    layer0_outputs(4439) <= '0';
    layer0_outputs(4440) <= '0';
    layer0_outputs(4441) <= not(inputs(183));
    layer0_outputs(4442) <= inputs(99);
    layer0_outputs(4443) <= inputs(235);
    layer0_outputs(4444) <= (inputs(169)) or (inputs(192));
    layer0_outputs(4445) <= (inputs(59)) or (inputs(91));
    layer0_outputs(4446) <= not(inputs(75));
    layer0_outputs(4447) <= '0';
    layer0_outputs(4448) <= inputs(110);
    layer0_outputs(4449) <= (inputs(254)) and not (inputs(86));
    layer0_outputs(4450) <= not(inputs(159));
    layer0_outputs(4451) <= not(inputs(220));
    layer0_outputs(4452) <= not((inputs(82)) xor (inputs(139)));
    layer0_outputs(4453) <= not(inputs(80));
    layer0_outputs(4454) <= '0';
    layer0_outputs(4455) <= inputs(199);
    layer0_outputs(4456) <= '0';
    layer0_outputs(4457) <= not((inputs(179)) and (inputs(27)));
    layer0_outputs(4458) <= not((inputs(80)) or (inputs(154)));
    layer0_outputs(4459) <= not((inputs(244)) and (inputs(165)));
    layer0_outputs(4460) <= inputs(239);
    layer0_outputs(4461) <= inputs(146);
    layer0_outputs(4462) <= not(inputs(165));
    layer0_outputs(4463) <= not(inputs(22));
    layer0_outputs(4464) <= (inputs(74)) or (inputs(6));
    layer0_outputs(4465) <= (inputs(89)) and not (inputs(110));
    layer0_outputs(4466) <= inputs(132);
    layer0_outputs(4467) <= not(inputs(122));
    layer0_outputs(4468) <= inputs(119);
    layer0_outputs(4469) <= not(inputs(187)) or (inputs(165));
    layer0_outputs(4470) <= not(inputs(21)) or (inputs(72));
    layer0_outputs(4471) <= '1';
    layer0_outputs(4472) <= inputs(200);
    layer0_outputs(4473) <= not(inputs(184)) or (inputs(28));
    layer0_outputs(4474) <= not(inputs(41));
    layer0_outputs(4475) <= not(inputs(142)) or (inputs(81));
    layer0_outputs(4476) <= (inputs(149)) and not (inputs(196));
    layer0_outputs(4477) <= not(inputs(102));
    layer0_outputs(4478) <= '1';
    layer0_outputs(4479) <= not(inputs(255));
    layer0_outputs(4480) <= not(inputs(38));
    layer0_outputs(4481) <= not((inputs(236)) and (inputs(93)));
    layer0_outputs(4482) <= (inputs(38)) or (inputs(21));
    layer0_outputs(4483) <= inputs(48);
    layer0_outputs(4484) <= '0';
    layer0_outputs(4485) <= inputs(28);
    layer0_outputs(4486) <= '0';
    layer0_outputs(4487) <= (inputs(152)) and not (inputs(145));
    layer0_outputs(4488) <= (inputs(237)) or (inputs(68));
    layer0_outputs(4489) <= (inputs(241)) and (inputs(32));
    layer0_outputs(4490) <= not((inputs(12)) xor (inputs(144)));
    layer0_outputs(4491) <= (inputs(165)) and not (inputs(76));
    layer0_outputs(4492) <= not(inputs(196));
    layer0_outputs(4493) <= not((inputs(18)) or (inputs(31)));
    layer0_outputs(4494) <= inputs(247);
    layer0_outputs(4495) <= '1';
    layer0_outputs(4496) <= not(inputs(89));
    layer0_outputs(4497) <= (inputs(232)) or (inputs(169));
    layer0_outputs(4498) <= '1';
    layer0_outputs(4499) <= not(inputs(152));
    layer0_outputs(4500) <= (inputs(57)) and (inputs(165));
    layer0_outputs(4501) <= inputs(10);
    layer0_outputs(4502) <= (inputs(182)) or (inputs(235));
    layer0_outputs(4503) <= (inputs(209)) and (inputs(139));
    layer0_outputs(4504) <= not(inputs(208)) or (inputs(236));
    layer0_outputs(4505) <= inputs(204);
    layer0_outputs(4506) <= '0';
    layer0_outputs(4507) <= inputs(186);
    layer0_outputs(4508) <= not((inputs(152)) xor (inputs(32)));
    layer0_outputs(4509) <= '0';
    layer0_outputs(4510) <= (inputs(195)) and not (inputs(16));
    layer0_outputs(4511) <= not(inputs(158)) or (inputs(30));
    layer0_outputs(4512) <= not(inputs(247));
    layer0_outputs(4513) <= not(inputs(148));
    layer0_outputs(4514) <= (inputs(37)) or (inputs(63));
    layer0_outputs(4515) <= not((inputs(91)) xor (inputs(109)));
    layer0_outputs(4516) <= not(inputs(222));
    layer0_outputs(4517) <= not((inputs(45)) and (inputs(249)));
    layer0_outputs(4518) <= not(inputs(175));
    layer0_outputs(4519) <= not(inputs(102));
    layer0_outputs(4520) <= not(inputs(205)) or (inputs(77));
    layer0_outputs(4521) <= not(inputs(127));
    layer0_outputs(4522) <= not(inputs(119));
    layer0_outputs(4523) <= '0';
    layer0_outputs(4524) <= not((inputs(241)) xor (inputs(50)));
    layer0_outputs(4525) <= (inputs(56)) and (inputs(243));
    layer0_outputs(4526) <= not((inputs(141)) or (inputs(205)));
    layer0_outputs(4527) <= not(inputs(67));
    layer0_outputs(4528) <= not(inputs(194));
    layer0_outputs(4529) <= not((inputs(15)) or (inputs(86)));
    layer0_outputs(4530) <= '1';
    layer0_outputs(4531) <= inputs(172);
    layer0_outputs(4532) <= (inputs(70)) and (inputs(72));
    layer0_outputs(4533) <= (inputs(97)) and not (inputs(164));
    layer0_outputs(4534) <= not(inputs(175)) or (inputs(158));
    layer0_outputs(4535) <= '1';
    layer0_outputs(4536) <= (inputs(235)) and not (inputs(48));
    layer0_outputs(4537) <= inputs(203);
    layer0_outputs(4538) <= (inputs(92)) and not (inputs(247));
    layer0_outputs(4539) <= (inputs(148)) and not (inputs(5));
    layer0_outputs(4540) <= (inputs(114)) and not (inputs(150));
    layer0_outputs(4541) <= inputs(128);
    layer0_outputs(4542) <= inputs(136);
    layer0_outputs(4543) <= not(inputs(176)) or (inputs(57));
    layer0_outputs(4544) <= '0';
    layer0_outputs(4545) <= not((inputs(221)) or (inputs(18)));
    layer0_outputs(4546) <= not(inputs(31));
    layer0_outputs(4547) <= (inputs(165)) xor (inputs(56));
    layer0_outputs(4548) <= (inputs(222)) xor (inputs(199));
    layer0_outputs(4549) <= (inputs(99)) and not (inputs(20));
    layer0_outputs(4550) <= inputs(3);
    layer0_outputs(4551) <= '1';
    layer0_outputs(4552) <= not(inputs(15)) or (inputs(234));
    layer0_outputs(4553) <= not(inputs(234)) or (inputs(151));
    layer0_outputs(4554) <= not(inputs(118)) or (inputs(75));
    layer0_outputs(4555) <= '0';
    layer0_outputs(4556) <= not((inputs(71)) or (inputs(89)));
    layer0_outputs(4557) <= '0';
    layer0_outputs(4558) <= '0';
    layer0_outputs(4559) <= '0';
    layer0_outputs(4560) <= not((inputs(52)) or (inputs(161)));
    layer0_outputs(4561) <= inputs(203);
    layer0_outputs(4562) <= (inputs(193)) and (inputs(5));
    layer0_outputs(4563) <= not(inputs(92)) or (inputs(41));
    layer0_outputs(4564) <= not((inputs(234)) or (inputs(69)));
    layer0_outputs(4565) <= inputs(97);
    layer0_outputs(4566) <= (inputs(202)) xor (inputs(5));
    layer0_outputs(4567) <= (inputs(24)) or (inputs(39));
    layer0_outputs(4568) <= '0';
    layer0_outputs(4569) <= inputs(162);
    layer0_outputs(4570) <= (inputs(145)) xor (inputs(198));
    layer0_outputs(4571) <= '0';
    layer0_outputs(4572) <= (inputs(92)) and not (inputs(34));
    layer0_outputs(4573) <= not(inputs(238)) or (inputs(123));
    layer0_outputs(4574) <= '0';
    layer0_outputs(4575) <= inputs(253);
    layer0_outputs(4576) <= not(inputs(232));
    layer0_outputs(4577) <= not(inputs(220));
    layer0_outputs(4578) <= (inputs(51)) and (inputs(164));
    layer0_outputs(4579) <= (inputs(195)) xor (inputs(237));
    layer0_outputs(4580) <= (inputs(30)) and not (inputs(219));
    layer0_outputs(4581) <= not((inputs(150)) and (inputs(54)));
    layer0_outputs(4582) <= not(inputs(222)) or (inputs(75));
    layer0_outputs(4583) <= not((inputs(11)) and (inputs(79)));
    layer0_outputs(4584) <= '1';
    layer0_outputs(4585) <= (inputs(92)) and not (inputs(125));
    layer0_outputs(4586) <= '1';
    layer0_outputs(4587) <= inputs(210);
    layer0_outputs(4588) <= inputs(134);
    layer0_outputs(4589) <= not((inputs(15)) or (inputs(45)));
    layer0_outputs(4590) <= (inputs(131)) and not (inputs(254));
    layer0_outputs(4591) <= '1';
    layer0_outputs(4592) <= not((inputs(210)) or (inputs(210)));
    layer0_outputs(4593) <= (inputs(154)) or (inputs(20));
    layer0_outputs(4594) <= inputs(252);
    layer0_outputs(4595) <= not(inputs(137));
    layer0_outputs(4596) <= not(inputs(236));
    layer0_outputs(4597) <= not(inputs(235));
    layer0_outputs(4598) <= not((inputs(134)) xor (inputs(128)));
    layer0_outputs(4599) <= inputs(141);
    layer0_outputs(4600) <= not((inputs(132)) or (inputs(181)));
    layer0_outputs(4601) <= not(inputs(125));
    layer0_outputs(4602) <= (inputs(189)) and not (inputs(111));
    layer0_outputs(4603) <= not((inputs(175)) and (inputs(67)));
    layer0_outputs(4604) <= (inputs(59)) and not (inputs(233));
    layer0_outputs(4605) <= (inputs(118)) and not (inputs(34));
    layer0_outputs(4606) <= not(inputs(135));
    layer0_outputs(4607) <= not(inputs(72));
    layer0_outputs(4608) <= not((inputs(94)) and (inputs(158)));
    layer0_outputs(4609) <= not((inputs(193)) xor (inputs(144)));
    layer0_outputs(4610) <= not(inputs(82));
    layer0_outputs(4611) <= inputs(65);
    layer0_outputs(4612) <= (inputs(215)) or (inputs(114));
    layer0_outputs(4613) <= inputs(215);
    layer0_outputs(4614) <= (inputs(143)) and not (inputs(124));
    layer0_outputs(4615) <= (inputs(79)) and (inputs(167));
    layer0_outputs(4616) <= not(inputs(74));
    layer0_outputs(4617) <= not((inputs(231)) or (inputs(61)));
    layer0_outputs(4618) <= not(inputs(32));
    layer0_outputs(4619) <= (inputs(10)) and not (inputs(181));
    layer0_outputs(4620) <= not((inputs(131)) or (inputs(20)));
    layer0_outputs(4621) <= not(inputs(195));
    layer0_outputs(4622) <= '1';
    layer0_outputs(4623) <= inputs(165);
    layer0_outputs(4624) <= not((inputs(109)) or (inputs(23)));
    layer0_outputs(4625) <= '0';
    layer0_outputs(4626) <= inputs(233);
    layer0_outputs(4627) <= inputs(76);
    layer0_outputs(4628) <= not(inputs(78)) or (inputs(166));
    layer0_outputs(4629) <= inputs(215);
    layer0_outputs(4630) <= not(inputs(229)) or (inputs(29));
    layer0_outputs(4631) <= not((inputs(16)) and (inputs(44)));
    layer0_outputs(4632) <= not((inputs(73)) xor (inputs(173)));
    layer0_outputs(4633) <= (inputs(203)) or (inputs(75));
    layer0_outputs(4634) <= '1';
    layer0_outputs(4635) <= not(inputs(243)) or (inputs(203));
    layer0_outputs(4636) <= not(inputs(210));
    layer0_outputs(4637) <= inputs(171);
    layer0_outputs(4638) <= inputs(224);
    layer0_outputs(4639) <= not(inputs(226));
    layer0_outputs(4640) <= inputs(87);
    layer0_outputs(4641) <= (inputs(70)) and (inputs(0));
    layer0_outputs(4642) <= not(inputs(131));
    layer0_outputs(4643) <= not(inputs(3));
    layer0_outputs(4644) <= (inputs(10)) and (inputs(82));
    layer0_outputs(4645) <= (inputs(212)) and (inputs(222));
    layer0_outputs(4646) <= not(inputs(56));
    layer0_outputs(4647) <= inputs(180);
    layer0_outputs(4648) <= inputs(159);
    layer0_outputs(4649) <= not((inputs(108)) xor (inputs(158)));
    layer0_outputs(4650) <= (inputs(67)) or (inputs(17));
    layer0_outputs(4651) <= (inputs(173)) and not (inputs(133));
    layer0_outputs(4652) <= not((inputs(229)) or (inputs(28)));
    layer0_outputs(4653) <= '0';
    layer0_outputs(4654) <= '1';
    layer0_outputs(4655) <= inputs(183);
    layer0_outputs(4656) <= '0';
    layer0_outputs(4657) <= not(inputs(163)) or (inputs(110));
    layer0_outputs(4658) <= not(inputs(18)) or (inputs(173));
    layer0_outputs(4659) <= not((inputs(189)) and (inputs(195)));
    layer0_outputs(4660) <= not(inputs(230));
    layer0_outputs(4661) <= (inputs(78)) and not (inputs(249));
    layer0_outputs(4662) <= not((inputs(182)) and (inputs(249)));
    layer0_outputs(4663) <= not(inputs(90));
    layer0_outputs(4664) <= '0';
    layer0_outputs(4665) <= (inputs(84)) or (inputs(119));
    layer0_outputs(4666) <= (inputs(102)) and not (inputs(106));
    layer0_outputs(4667) <= not((inputs(251)) and (inputs(144)));
    layer0_outputs(4668) <= inputs(197);
    layer0_outputs(4669) <= (inputs(128)) xor (inputs(223));
    layer0_outputs(4670) <= not((inputs(246)) and (inputs(106)));
    layer0_outputs(4671) <= not(inputs(112));
    layer0_outputs(4672) <= inputs(235);
    layer0_outputs(4673) <= (inputs(245)) and not (inputs(60));
    layer0_outputs(4674) <= '0';
    layer0_outputs(4675) <= not(inputs(141)) or (inputs(184));
    layer0_outputs(4676) <= not(inputs(140));
    layer0_outputs(4677) <= inputs(165);
    layer0_outputs(4678) <= '0';
    layer0_outputs(4679) <= (inputs(108)) and not (inputs(183));
    layer0_outputs(4680) <= not(inputs(121)) or (inputs(1));
    layer0_outputs(4681) <= (inputs(162)) and not (inputs(159));
    layer0_outputs(4682) <= '1';
    layer0_outputs(4683) <= not((inputs(216)) or (inputs(208)));
    layer0_outputs(4684) <= '0';
    layer0_outputs(4685) <= not(inputs(221)) or (inputs(148));
    layer0_outputs(4686) <= (inputs(83)) or (inputs(243));
    layer0_outputs(4687) <= not(inputs(158));
    layer0_outputs(4688) <= not(inputs(98)) or (inputs(144));
    layer0_outputs(4689) <= not((inputs(72)) and (inputs(19)));
    layer0_outputs(4690) <= not((inputs(145)) and (inputs(75)));
    layer0_outputs(4691) <= inputs(205);
    layer0_outputs(4692) <= not((inputs(30)) or (inputs(76)));
    layer0_outputs(4693) <= not((inputs(113)) or (inputs(147)));
    layer0_outputs(4694) <= '1';
    layer0_outputs(4695) <= not(inputs(214));
    layer0_outputs(4696) <= (inputs(232)) or (inputs(141));
    layer0_outputs(4697) <= (inputs(13)) and not (inputs(169));
    layer0_outputs(4698) <= inputs(105);
    layer0_outputs(4699) <= (inputs(229)) and not (inputs(187));
    layer0_outputs(4700) <= not((inputs(205)) and (inputs(55)));
    layer0_outputs(4701) <= not(inputs(94));
    layer0_outputs(4702) <= not(inputs(181));
    layer0_outputs(4703) <= not((inputs(202)) or (inputs(240)));
    layer0_outputs(4704) <= (inputs(111)) or (inputs(37));
    layer0_outputs(4705) <= not((inputs(6)) and (inputs(13)));
    layer0_outputs(4706) <= (inputs(130)) or (inputs(37));
    layer0_outputs(4707) <= not((inputs(210)) and (inputs(204)));
    layer0_outputs(4708) <= (inputs(153)) and not (inputs(178));
    layer0_outputs(4709) <= (inputs(215)) and not (inputs(23));
    layer0_outputs(4710) <= not(inputs(184));
    layer0_outputs(4711) <= not(inputs(73)) or (inputs(223));
    layer0_outputs(4712) <= inputs(219);
    layer0_outputs(4713) <= not((inputs(161)) xor (inputs(236)));
    layer0_outputs(4714) <= not((inputs(152)) or (inputs(45)));
    layer0_outputs(4715) <= (inputs(244)) and not (inputs(130));
    layer0_outputs(4716) <= (inputs(225)) and (inputs(183));
    layer0_outputs(4717) <= inputs(177);
    layer0_outputs(4718) <= (inputs(8)) and (inputs(76));
    layer0_outputs(4719) <= '1';
    layer0_outputs(4720) <= inputs(63);
    layer0_outputs(4721) <= (inputs(157)) or (inputs(188));
    layer0_outputs(4722) <= '0';
    layer0_outputs(4723) <= not(inputs(64));
    layer0_outputs(4724) <= not(inputs(109)) or (inputs(213));
    layer0_outputs(4725) <= (inputs(6)) and (inputs(49));
    layer0_outputs(4726) <= '0';
    layer0_outputs(4727) <= not(inputs(155));
    layer0_outputs(4728) <= '1';
    layer0_outputs(4729) <= (inputs(26)) or (inputs(172));
    layer0_outputs(4730) <= not(inputs(13));
    layer0_outputs(4731) <= (inputs(228)) or (inputs(31));
    layer0_outputs(4732) <= (inputs(131)) or (inputs(110));
    layer0_outputs(4733) <= not(inputs(5)) or (inputs(220));
    layer0_outputs(4734) <= (inputs(104)) and not (inputs(182));
    layer0_outputs(4735) <= (inputs(211)) or (inputs(193));
    layer0_outputs(4736) <= '0';
    layer0_outputs(4737) <= not((inputs(179)) or (inputs(168)));
    layer0_outputs(4738) <= not(inputs(85));
    layer0_outputs(4739) <= not(inputs(3));
    layer0_outputs(4740) <= not((inputs(251)) xor (inputs(222)));
    layer0_outputs(4741) <= '0';
    layer0_outputs(4742) <= not(inputs(179));
    layer0_outputs(4743) <= '0';
    layer0_outputs(4744) <= (inputs(43)) and not (inputs(91));
    layer0_outputs(4745) <= not((inputs(35)) or (inputs(248)));
    layer0_outputs(4746) <= '1';
    layer0_outputs(4747) <= '1';
    layer0_outputs(4748) <= inputs(152);
    layer0_outputs(4749) <= not((inputs(95)) or (inputs(22)));
    layer0_outputs(4750) <= not(inputs(119)) or (inputs(130));
    layer0_outputs(4751) <= '1';
    layer0_outputs(4752) <= (inputs(216)) and not (inputs(60));
    layer0_outputs(4753) <= not((inputs(1)) or (inputs(90)));
    layer0_outputs(4754) <= not(inputs(98)) or (inputs(106));
    layer0_outputs(4755) <= '0';
    layer0_outputs(4756) <= (inputs(220)) or (inputs(53));
    layer0_outputs(4757) <= not(inputs(175));
    layer0_outputs(4758) <= not(inputs(162));
    layer0_outputs(4759) <= '0';
    layer0_outputs(4760) <= inputs(2);
    layer0_outputs(4761) <= not(inputs(124));
    layer0_outputs(4762) <= '1';
    layer0_outputs(4763) <= (inputs(0)) and (inputs(102));
    layer0_outputs(4764) <= inputs(134);
    layer0_outputs(4765) <= inputs(149);
    layer0_outputs(4766) <= not(inputs(45)) or (inputs(74));
    layer0_outputs(4767) <= not((inputs(132)) or (inputs(31)));
    layer0_outputs(4768) <= inputs(215);
    layer0_outputs(4769) <= inputs(198);
    layer0_outputs(4770) <= not(inputs(198));
    layer0_outputs(4771) <= not((inputs(176)) and (inputs(237)));
    layer0_outputs(4772) <= (inputs(152)) or (inputs(34));
    layer0_outputs(4773) <= not(inputs(228)) or (inputs(240));
    layer0_outputs(4774) <= (inputs(206)) and not (inputs(23));
    layer0_outputs(4775) <= inputs(108);
    layer0_outputs(4776) <= '0';
    layer0_outputs(4777) <= inputs(65);
    layer0_outputs(4778) <= inputs(0);
    layer0_outputs(4779) <= (inputs(3)) and not (inputs(1));
    layer0_outputs(4780) <= not((inputs(71)) xor (inputs(69)));
    layer0_outputs(4781) <= not(inputs(188)) or (inputs(40));
    layer0_outputs(4782) <= not((inputs(18)) xor (inputs(54)));
    layer0_outputs(4783) <= inputs(228);
    layer0_outputs(4784) <= not(inputs(26));
    layer0_outputs(4785) <= (inputs(60)) xor (inputs(94));
    layer0_outputs(4786) <= (inputs(64)) or (inputs(150));
    layer0_outputs(4787) <= '0';
    layer0_outputs(4788) <= (inputs(156)) and not (inputs(2));
    layer0_outputs(4789) <= (inputs(176)) or (inputs(206));
    layer0_outputs(4790) <= inputs(100);
    layer0_outputs(4791) <= inputs(127);
    layer0_outputs(4792) <= '0';
    layer0_outputs(4793) <= '1';
    layer0_outputs(4794) <= not(inputs(100));
    layer0_outputs(4795) <= inputs(86);
    layer0_outputs(4796) <= (inputs(145)) and not (inputs(142));
    layer0_outputs(4797) <= not(inputs(125)) or (inputs(24));
    layer0_outputs(4798) <= not(inputs(103)) or (inputs(4));
    layer0_outputs(4799) <= not(inputs(107)) or (inputs(238));
    layer0_outputs(4800) <= not(inputs(13)) or (inputs(232));
    layer0_outputs(4801) <= not((inputs(161)) and (inputs(106)));
    layer0_outputs(4802) <= (inputs(105)) and not (inputs(112));
    layer0_outputs(4803) <= inputs(52);
    layer0_outputs(4804) <= not(inputs(96)) or (inputs(198));
    layer0_outputs(4805) <= (inputs(60)) xor (inputs(28));
    layer0_outputs(4806) <= not((inputs(236)) or (inputs(178)));
    layer0_outputs(4807) <= inputs(248);
    layer0_outputs(4808) <= '0';
    layer0_outputs(4809) <= not(inputs(74));
    layer0_outputs(4810) <= not((inputs(252)) xor (inputs(71)));
    layer0_outputs(4811) <= not((inputs(208)) or (inputs(135)));
    layer0_outputs(4812) <= inputs(177);
    layer0_outputs(4813) <= not(inputs(187)) or (inputs(154));
    layer0_outputs(4814) <= '1';
    layer0_outputs(4815) <= '1';
    layer0_outputs(4816) <= (inputs(120)) and not (inputs(197));
    layer0_outputs(4817) <= (inputs(23)) and not (inputs(212));
    layer0_outputs(4818) <= not(inputs(150));
    layer0_outputs(4819) <= (inputs(69)) and not (inputs(209));
    layer0_outputs(4820) <= inputs(166);
    layer0_outputs(4821) <= not((inputs(132)) or (inputs(190)));
    layer0_outputs(4822) <= '1';
    layer0_outputs(4823) <= (inputs(85)) and not (inputs(254));
    layer0_outputs(4824) <= '0';
    layer0_outputs(4825) <= inputs(116);
    layer0_outputs(4826) <= not((inputs(185)) and (inputs(179)));
    layer0_outputs(4827) <= not(inputs(129));
    layer0_outputs(4828) <= '0';
    layer0_outputs(4829) <= not(inputs(247));
    layer0_outputs(4830) <= '0';
    layer0_outputs(4831) <= (inputs(164)) or (inputs(165));
    layer0_outputs(4832) <= '1';
    layer0_outputs(4833) <= (inputs(104)) xor (inputs(251));
    layer0_outputs(4834) <= not(inputs(233)) or (inputs(209));
    layer0_outputs(4835) <= not(inputs(171)) or (inputs(230));
    layer0_outputs(4836) <= not(inputs(234)) or (inputs(247));
    layer0_outputs(4837) <= not(inputs(210)) or (inputs(122));
    layer0_outputs(4838) <= (inputs(172)) xor (inputs(196));
    layer0_outputs(4839) <= not(inputs(46));
    layer0_outputs(4840) <= inputs(51);
    layer0_outputs(4841) <= not(inputs(27));
    layer0_outputs(4842) <= not(inputs(193)) or (inputs(6));
    layer0_outputs(4843) <= (inputs(230)) and (inputs(78));
    layer0_outputs(4844) <= not(inputs(212)) or (inputs(181));
    layer0_outputs(4845) <= not(inputs(94));
    layer0_outputs(4846) <= (inputs(167)) or (inputs(227));
    layer0_outputs(4847) <= inputs(109);
    layer0_outputs(4848) <= (inputs(71)) and not (inputs(133));
    layer0_outputs(4849) <= not((inputs(232)) or (inputs(199)));
    layer0_outputs(4850) <= (inputs(0)) or (inputs(207));
    layer0_outputs(4851) <= (inputs(196)) or (inputs(212));
    layer0_outputs(4852) <= (inputs(4)) xor (inputs(246));
    layer0_outputs(4853) <= '0';
    layer0_outputs(4854) <= (inputs(218)) and not (inputs(155));
    layer0_outputs(4855) <= not(inputs(10));
    layer0_outputs(4856) <= not(inputs(237));
    layer0_outputs(4857) <= (inputs(26)) and not (inputs(235));
    layer0_outputs(4858) <= not(inputs(146));
    layer0_outputs(4859) <= (inputs(48)) and not (inputs(170));
    layer0_outputs(4860) <= not(inputs(188));
    layer0_outputs(4861) <= inputs(239);
    layer0_outputs(4862) <= inputs(34);
    layer0_outputs(4863) <= not(inputs(4));
    layer0_outputs(4864) <= (inputs(135)) and not (inputs(54));
    layer0_outputs(4865) <= not(inputs(124)) or (inputs(253));
    layer0_outputs(4866) <= '0';
    layer0_outputs(4867) <= (inputs(11)) and (inputs(15));
    layer0_outputs(4868) <= not((inputs(2)) and (inputs(148)));
    layer0_outputs(4869) <= inputs(155);
    layer0_outputs(4870) <= (inputs(144)) or (inputs(111));
    layer0_outputs(4871) <= not((inputs(186)) xor (inputs(113)));
    layer0_outputs(4872) <= '0';
    layer0_outputs(4873) <= '1';
    layer0_outputs(4874) <= not(inputs(111));
    layer0_outputs(4875) <= '1';
    layer0_outputs(4876) <= inputs(152);
    layer0_outputs(4877) <= (inputs(39)) or (inputs(150));
    layer0_outputs(4878) <= not((inputs(5)) or (inputs(73)));
    layer0_outputs(4879) <= not(inputs(88));
    layer0_outputs(4880) <= (inputs(94)) and not (inputs(255));
    layer0_outputs(4881) <= inputs(68);
    layer0_outputs(4882) <= inputs(62);
    layer0_outputs(4883) <= '0';
    layer0_outputs(4884) <= '0';
    layer0_outputs(4885) <= (inputs(53)) xor (inputs(62));
    layer0_outputs(4886) <= inputs(91);
    layer0_outputs(4887) <= not(inputs(93)) or (inputs(140));
    layer0_outputs(4888) <= '0';
    layer0_outputs(4889) <= not(inputs(60));
    layer0_outputs(4890) <= '0';
    layer0_outputs(4891) <= not(inputs(179));
    layer0_outputs(4892) <= not((inputs(207)) and (inputs(109)));
    layer0_outputs(4893) <= (inputs(223)) xor (inputs(28));
    layer0_outputs(4894) <= not((inputs(79)) or (inputs(70)));
    layer0_outputs(4895) <= (inputs(231)) and not (inputs(163));
    layer0_outputs(4896) <= (inputs(182)) and not (inputs(62));
    layer0_outputs(4897) <= not((inputs(86)) and (inputs(54)));
    layer0_outputs(4898) <= '0';
    layer0_outputs(4899) <= (inputs(224)) or (inputs(101));
    layer0_outputs(4900) <= inputs(52);
    layer0_outputs(4901) <= inputs(115);
    layer0_outputs(4902) <= inputs(44);
    layer0_outputs(4903) <= (inputs(165)) and not (inputs(68));
    layer0_outputs(4904) <= not(inputs(11));
    layer0_outputs(4905) <= (inputs(153)) and not (inputs(202));
    layer0_outputs(4906) <= '0';
    layer0_outputs(4907) <= (inputs(231)) and not (inputs(121));
    layer0_outputs(4908) <= not((inputs(183)) xor (inputs(254)));
    layer0_outputs(4909) <= inputs(203);
    layer0_outputs(4910) <= not(inputs(123)) or (inputs(160));
    layer0_outputs(4911) <= not(inputs(189));
    layer0_outputs(4912) <= inputs(104);
    layer0_outputs(4913) <= not((inputs(90)) or (inputs(110)));
    layer0_outputs(4914) <= inputs(208);
    layer0_outputs(4915) <= inputs(59);
    layer0_outputs(4916) <= inputs(152);
    layer0_outputs(4917) <= (inputs(41)) or (inputs(58));
    layer0_outputs(4918) <= '0';
    layer0_outputs(4919) <= inputs(71);
    layer0_outputs(4920) <= (inputs(174)) and not (inputs(129));
    layer0_outputs(4921) <= not(inputs(228));
    layer0_outputs(4922) <= inputs(136);
    layer0_outputs(4923) <= inputs(20);
    layer0_outputs(4924) <= not((inputs(182)) and (inputs(220)));
    layer0_outputs(4925) <= '1';
    layer0_outputs(4926) <= not((inputs(98)) or (inputs(163)));
    layer0_outputs(4927) <= '1';
    layer0_outputs(4928) <= not(inputs(158)) or (inputs(184));
    layer0_outputs(4929) <= '1';
    layer0_outputs(4930) <= '0';
    layer0_outputs(4931) <= (inputs(135)) and not (inputs(46));
    layer0_outputs(4932) <= not(inputs(223)) or (inputs(18));
    layer0_outputs(4933) <= '1';
    layer0_outputs(4934) <= (inputs(148)) and (inputs(65));
    layer0_outputs(4935) <= (inputs(196)) and not (inputs(136));
    layer0_outputs(4936) <= (inputs(203)) xor (inputs(228));
    layer0_outputs(4937) <= (inputs(124)) and (inputs(11));
    layer0_outputs(4938) <= '1';
    layer0_outputs(4939) <= (inputs(231)) and not (inputs(110));
    layer0_outputs(4940) <= not(inputs(89));
    layer0_outputs(4941) <= not(inputs(100));
    layer0_outputs(4942) <= not(inputs(100)) or (inputs(74));
    layer0_outputs(4943) <= (inputs(74)) and not (inputs(73));
    layer0_outputs(4944) <= not(inputs(237));
    layer0_outputs(4945) <= inputs(58);
    layer0_outputs(4946) <= not(inputs(3));
    layer0_outputs(4947) <= not((inputs(213)) and (inputs(208)));
    layer0_outputs(4948) <= inputs(75);
    layer0_outputs(4949) <= not((inputs(180)) or (inputs(117)));
    layer0_outputs(4950) <= '0';
    layer0_outputs(4951) <= not(inputs(248));
    layer0_outputs(4952) <= not((inputs(188)) or (inputs(187)));
    layer0_outputs(4953) <= (inputs(186)) and (inputs(120));
    layer0_outputs(4954) <= (inputs(132)) and not (inputs(246));
    layer0_outputs(4955) <= not(inputs(80));
    layer0_outputs(4956) <= (inputs(104)) and not (inputs(4));
    layer0_outputs(4957) <= '0';
    layer0_outputs(4958) <= not(inputs(249)) or (inputs(148));
    layer0_outputs(4959) <= inputs(79);
    layer0_outputs(4960) <= inputs(213);
    layer0_outputs(4961) <= (inputs(100)) or (inputs(90));
    layer0_outputs(4962) <= not(inputs(171));
    layer0_outputs(4963) <= (inputs(126)) and not (inputs(65));
    layer0_outputs(4964) <= not((inputs(122)) and (inputs(224)));
    layer0_outputs(4965) <= inputs(17);
    layer0_outputs(4966) <= (inputs(172)) or (inputs(96));
    layer0_outputs(4967) <= not(inputs(116)) or (inputs(233));
    layer0_outputs(4968) <= not((inputs(132)) or (inputs(219)));
    layer0_outputs(4969) <= not(inputs(227));
    layer0_outputs(4970) <= (inputs(140)) and not (inputs(150));
    layer0_outputs(4971) <= (inputs(166)) and not (inputs(76));
    layer0_outputs(4972) <= inputs(59);
    layer0_outputs(4973) <= not((inputs(212)) or (inputs(191)));
    layer0_outputs(4974) <= not(inputs(186)) or (inputs(82));
    layer0_outputs(4975) <= not(inputs(115));
    layer0_outputs(4976) <= not((inputs(97)) or (inputs(124)));
    layer0_outputs(4977) <= not(inputs(197));
    layer0_outputs(4978) <= (inputs(143)) and not (inputs(112));
    layer0_outputs(4979) <= not(inputs(60)) or (inputs(48));
    layer0_outputs(4980) <= inputs(223);
    layer0_outputs(4981) <= (inputs(203)) or (inputs(82));
    layer0_outputs(4982) <= '0';
    layer0_outputs(4983) <= '1';
    layer0_outputs(4984) <= '1';
    layer0_outputs(4985) <= '1';
    layer0_outputs(4986) <= '1';
    layer0_outputs(4987) <= '0';
    layer0_outputs(4988) <= (inputs(27)) or (inputs(154));
    layer0_outputs(4989) <= inputs(232);
    layer0_outputs(4990) <= inputs(24);
    layer0_outputs(4991) <= inputs(177);
    layer0_outputs(4992) <= (inputs(214)) and not (inputs(108));
    layer0_outputs(4993) <= not(inputs(159)) or (inputs(87));
    layer0_outputs(4994) <= '1';
    layer0_outputs(4995) <= (inputs(95)) and not (inputs(43));
    layer0_outputs(4996) <= not(inputs(158));
    layer0_outputs(4997) <= inputs(94);
    layer0_outputs(4998) <= '1';
    layer0_outputs(4999) <= not(inputs(205));
    layer0_outputs(5000) <= inputs(141);
    layer0_outputs(5001) <= (inputs(163)) and not (inputs(14));
    layer0_outputs(5002) <= not(inputs(186));
    layer0_outputs(5003) <= (inputs(197)) or (inputs(175));
    layer0_outputs(5004) <= (inputs(21)) xor (inputs(22));
    layer0_outputs(5005) <= '0';
    layer0_outputs(5006) <= not((inputs(18)) or (inputs(192)));
    layer0_outputs(5007) <= not((inputs(226)) and (inputs(65)));
    layer0_outputs(5008) <= (inputs(57)) and (inputs(171));
    layer0_outputs(5009) <= not((inputs(249)) and (inputs(87)));
    layer0_outputs(5010) <= not(inputs(36)) or (inputs(130));
    layer0_outputs(5011) <= (inputs(123)) or (inputs(62));
    layer0_outputs(5012) <= inputs(109);
    layer0_outputs(5013) <= '1';
    layer0_outputs(5014) <= inputs(230);
    layer0_outputs(5015) <= (inputs(21)) or (inputs(254));
    layer0_outputs(5016) <= not(inputs(206)) or (inputs(16));
    layer0_outputs(5017) <= (inputs(221)) and not (inputs(64));
    layer0_outputs(5018) <= not(inputs(172)) or (inputs(114));
    layer0_outputs(5019) <= inputs(94);
    layer0_outputs(5020) <= not(inputs(21)) or (inputs(189));
    layer0_outputs(5021) <= not(inputs(88));
    layer0_outputs(5022) <= not(inputs(166)) or (inputs(249));
    layer0_outputs(5023) <= inputs(23);
    layer0_outputs(5024) <= '0';
    layer0_outputs(5025) <= not(inputs(168)) or (inputs(170));
    layer0_outputs(5026) <= '1';
    layer0_outputs(5027) <= not(inputs(2));
    layer0_outputs(5028) <= not(inputs(64)) or (inputs(150));
    layer0_outputs(5029) <= '1';
    layer0_outputs(5030) <= (inputs(68)) xor (inputs(229));
    layer0_outputs(5031) <= (inputs(215)) and (inputs(254));
    layer0_outputs(5032) <= (inputs(12)) and not (inputs(200));
    layer0_outputs(5033) <= (inputs(7)) and not (inputs(113));
    layer0_outputs(5034) <= (inputs(153)) and not (inputs(123));
    layer0_outputs(5035) <= '0';
    layer0_outputs(5036) <= inputs(110);
    layer0_outputs(5037) <= (inputs(201)) and (inputs(197));
    layer0_outputs(5038) <= inputs(120);
    layer0_outputs(5039) <= inputs(93);
    layer0_outputs(5040) <= not(inputs(93)) or (inputs(132));
    layer0_outputs(5041) <= (inputs(113)) or (inputs(163));
    layer0_outputs(5042) <= '0';
    layer0_outputs(5043) <= not(inputs(6)) or (inputs(13));
    layer0_outputs(5044) <= not(inputs(183)) or (inputs(62));
    layer0_outputs(5045) <= not((inputs(105)) xor (inputs(156)));
    layer0_outputs(5046) <= not(inputs(202)) or (inputs(66));
    layer0_outputs(5047) <= '1';
    layer0_outputs(5048) <= inputs(224);
    layer0_outputs(5049) <= not(inputs(144));
    layer0_outputs(5050) <= '1';
    layer0_outputs(5051) <= '1';
    layer0_outputs(5052) <= (inputs(49)) and not (inputs(153));
    layer0_outputs(5053) <= not((inputs(161)) and (inputs(210)));
    layer0_outputs(5054) <= not(inputs(38));
    layer0_outputs(5055) <= not(inputs(148));
    layer0_outputs(5056) <= (inputs(5)) and not (inputs(232));
    layer0_outputs(5057) <= inputs(232);
    layer0_outputs(5058) <= (inputs(113)) and (inputs(23));
    layer0_outputs(5059) <= (inputs(88)) xor (inputs(90));
    layer0_outputs(5060) <= '0';
    layer0_outputs(5061) <= not(inputs(25));
    layer0_outputs(5062) <= not(inputs(15)) or (inputs(242));
    layer0_outputs(5063) <= inputs(32);
    layer0_outputs(5064) <= (inputs(175)) or (inputs(107));
    layer0_outputs(5065) <= not(inputs(150));
    layer0_outputs(5066) <= not((inputs(175)) or (inputs(251)));
    layer0_outputs(5067) <= not((inputs(3)) xor (inputs(29)));
    layer0_outputs(5068) <= (inputs(238)) and (inputs(42));
    layer0_outputs(5069) <= not(inputs(199));
    layer0_outputs(5070) <= not((inputs(201)) or (inputs(45)));
    layer0_outputs(5071) <= inputs(86);
    layer0_outputs(5072) <= inputs(95);
    layer0_outputs(5073) <= not(inputs(124)) or (inputs(34));
    layer0_outputs(5074) <= not((inputs(233)) and (inputs(32)));
    layer0_outputs(5075) <= not(inputs(151));
    layer0_outputs(5076) <= (inputs(43)) xor (inputs(9));
    layer0_outputs(5077) <= not(inputs(255));
    layer0_outputs(5078) <= inputs(164);
    layer0_outputs(5079) <= not((inputs(223)) or (inputs(56)));
    layer0_outputs(5080) <= (inputs(60)) or (inputs(47));
    layer0_outputs(5081) <= not(inputs(201)) or (inputs(245));
    layer0_outputs(5082) <= (inputs(253)) xor (inputs(221));
    layer0_outputs(5083) <= not(inputs(117)) or (inputs(191));
    layer0_outputs(5084) <= '1';
    layer0_outputs(5085) <= not(inputs(64)) or (inputs(85));
    layer0_outputs(5086) <= '0';
    layer0_outputs(5087) <= inputs(173);
    layer0_outputs(5088) <= not((inputs(151)) and (inputs(254)));
    layer0_outputs(5089) <= (inputs(57)) and (inputs(76));
    layer0_outputs(5090) <= '0';
    layer0_outputs(5091) <= '0';
    layer0_outputs(5092) <= (inputs(179)) or (inputs(46));
    layer0_outputs(5093) <= inputs(136);
    layer0_outputs(5094) <= not(inputs(114)) or (inputs(166));
    layer0_outputs(5095) <= '1';
    layer0_outputs(5096) <= not(inputs(90));
    layer0_outputs(5097) <= (inputs(76)) and (inputs(120));
    layer0_outputs(5098) <= not((inputs(237)) and (inputs(16)));
    layer0_outputs(5099) <= '1';
    layer0_outputs(5100) <= inputs(128);
    layer0_outputs(5101) <= not(inputs(229));
    layer0_outputs(5102) <= '0';
    layer0_outputs(5103) <= not(inputs(218)) or (inputs(164));
    layer0_outputs(5104) <= inputs(151);
    layer0_outputs(5105) <= '0';
    layer0_outputs(5106) <= (inputs(74)) and (inputs(104));
    layer0_outputs(5107) <= (inputs(61)) and not (inputs(107));
    layer0_outputs(5108) <= not((inputs(255)) or (inputs(143)));
    layer0_outputs(5109) <= not(inputs(175));
    layer0_outputs(5110) <= not(inputs(202));
    layer0_outputs(5111) <= not(inputs(66));
    layer0_outputs(5112) <= inputs(51);
    layer0_outputs(5113) <= not((inputs(145)) and (inputs(65)));
    layer0_outputs(5114) <= not(inputs(88)) or (inputs(221));
    layer0_outputs(5115) <= not((inputs(231)) and (inputs(169)));
    layer0_outputs(5116) <= (inputs(130)) or (inputs(173));
    layer0_outputs(5117) <= (inputs(49)) and (inputs(26));
    layer0_outputs(5118) <= (inputs(255)) and (inputs(238));
    layer0_outputs(5119) <= inputs(79);
    layer0_outputs(5120) <= not((inputs(140)) or (inputs(108)));
    layer0_outputs(5121) <= not(inputs(198)) or (inputs(176));
    layer0_outputs(5122) <= '0';
    layer0_outputs(5123) <= inputs(179);
    layer0_outputs(5124) <= inputs(59);
    layer0_outputs(5125) <= (inputs(254)) or (inputs(177));
    layer0_outputs(5126) <= (inputs(241)) xor (inputs(42));
    layer0_outputs(5127) <= not(inputs(230));
    layer0_outputs(5128) <= (inputs(54)) or (inputs(126));
    layer0_outputs(5129) <= (inputs(129)) or (inputs(4));
    layer0_outputs(5130) <= not((inputs(16)) or (inputs(81)));
    layer0_outputs(5131) <= not((inputs(33)) or (inputs(217)));
    layer0_outputs(5132) <= inputs(105);
    layer0_outputs(5133) <= not((inputs(50)) or (inputs(152)));
    layer0_outputs(5134) <= inputs(183);
    layer0_outputs(5135) <= '1';
    layer0_outputs(5136) <= (inputs(29)) and not (inputs(185));
    layer0_outputs(5137) <= not(inputs(4)) or (inputs(198));
    layer0_outputs(5138) <= not(inputs(230));
    layer0_outputs(5139) <= (inputs(186)) and not (inputs(253));
    layer0_outputs(5140) <= not(inputs(213)) or (inputs(30));
    layer0_outputs(5141) <= (inputs(62)) and (inputs(61));
    layer0_outputs(5142) <= '0';
    layer0_outputs(5143) <= inputs(189);
    layer0_outputs(5144) <= not(inputs(126));
    layer0_outputs(5145) <= not(inputs(162)) or (inputs(204));
    layer0_outputs(5146) <= (inputs(46)) and not (inputs(230));
    layer0_outputs(5147) <= not(inputs(73));
    layer0_outputs(5148) <= '1';
    layer0_outputs(5149) <= (inputs(243)) xor (inputs(180));
    layer0_outputs(5150) <= not((inputs(90)) and (inputs(106)));
    layer0_outputs(5151) <= '1';
    layer0_outputs(5152) <= not(inputs(10)) or (inputs(235));
    layer0_outputs(5153) <= (inputs(218)) or (inputs(122));
    layer0_outputs(5154) <= not((inputs(26)) and (inputs(54)));
    layer0_outputs(5155) <= not((inputs(162)) or (inputs(57)));
    layer0_outputs(5156) <= '1';
    layer0_outputs(5157) <= not((inputs(204)) or (inputs(176)));
    layer0_outputs(5158) <= '1';
    layer0_outputs(5159) <= '1';
    layer0_outputs(5160) <= not(inputs(19));
    layer0_outputs(5161) <= (inputs(241)) and not (inputs(102));
    layer0_outputs(5162) <= (inputs(255)) or (inputs(134));
    layer0_outputs(5163) <= (inputs(26)) or (inputs(252));
    layer0_outputs(5164) <= not(inputs(41));
    layer0_outputs(5165) <= '1';
    layer0_outputs(5166) <= (inputs(239)) and (inputs(190));
    layer0_outputs(5167) <= inputs(141);
    layer0_outputs(5168) <= (inputs(193)) and (inputs(164));
    layer0_outputs(5169) <= not((inputs(143)) or (inputs(94)));
    layer0_outputs(5170) <= not(inputs(122));
    layer0_outputs(5171) <= (inputs(23)) xor (inputs(1));
    layer0_outputs(5172) <= (inputs(73)) and not (inputs(83));
    layer0_outputs(5173) <= not((inputs(75)) and (inputs(179)));
    layer0_outputs(5174) <= inputs(254);
    layer0_outputs(5175) <= (inputs(92)) and not (inputs(58));
    layer0_outputs(5176) <= inputs(4);
    layer0_outputs(5177) <= (inputs(221)) or (inputs(239));
    layer0_outputs(5178) <= (inputs(226)) and not (inputs(92));
    layer0_outputs(5179) <= inputs(76);
    layer0_outputs(5180) <= '1';
    layer0_outputs(5181) <= not(inputs(189));
    layer0_outputs(5182) <= (inputs(228)) and not (inputs(166));
    layer0_outputs(5183) <= not((inputs(194)) and (inputs(225)));
    layer0_outputs(5184) <= not((inputs(206)) and (inputs(138)));
    layer0_outputs(5185) <= (inputs(207)) or (inputs(142));
    layer0_outputs(5186) <= not(inputs(248));
    layer0_outputs(5187) <= not(inputs(45)) or (inputs(201));
    layer0_outputs(5188) <= not(inputs(85)) or (inputs(221));
    layer0_outputs(5189) <= (inputs(90)) and (inputs(238));
    layer0_outputs(5190) <= '0';
    layer0_outputs(5191) <= inputs(214);
    layer0_outputs(5192) <= not(inputs(161)) or (inputs(108));
    layer0_outputs(5193) <= not(inputs(96));
    layer0_outputs(5194) <= not(inputs(162)) or (inputs(33));
    layer0_outputs(5195) <= (inputs(219)) or (inputs(132));
    layer0_outputs(5196) <= inputs(88);
    layer0_outputs(5197) <= '0';
    layer0_outputs(5198) <= '1';
    layer0_outputs(5199) <= inputs(185);
    layer0_outputs(5200) <= (inputs(254)) or (inputs(123));
    layer0_outputs(5201) <= not(inputs(184));
    layer0_outputs(5202) <= not(inputs(90));
    layer0_outputs(5203) <= not(inputs(97)) or (inputs(42));
    layer0_outputs(5204) <= not((inputs(14)) or (inputs(214)));
    layer0_outputs(5205) <= (inputs(175)) and (inputs(188));
    layer0_outputs(5206) <= '0';
    layer0_outputs(5207) <= not(inputs(196)) or (inputs(44));
    layer0_outputs(5208) <= not((inputs(68)) xor (inputs(81)));
    layer0_outputs(5209) <= '1';
    layer0_outputs(5210) <= (inputs(97)) and not (inputs(22));
    layer0_outputs(5211) <= not(inputs(120));
    layer0_outputs(5212) <= not(inputs(207)) or (inputs(35));
    layer0_outputs(5213) <= inputs(33);
    layer0_outputs(5214) <= not(inputs(209));
    layer0_outputs(5215) <= inputs(211);
    layer0_outputs(5216) <= (inputs(173)) and not (inputs(172));
    layer0_outputs(5217) <= not(inputs(23));
    layer0_outputs(5218) <= (inputs(154)) and not (inputs(199));
    layer0_outputs(5219) <= not(inputs(90)) or (inputs(163));
    layer0_outputs(5220) <= not((inputs(228)) or (inputs(162)));
    layer0_outputs(5221) <= '1';
    layer0_outputs(5222) <= inputs(129);
    layer0_outputs(5223) <= not(inputs(80));
    layer0_outputs(5224) <= not((inputs(37)) or (inputs(94)));
    layer0_outputs(5225) <= not(inputs(241));
    layer0_outputs(5226) <= (inputs(166)) and not (inputs(54));
    layer0_outputs(5227) <= not((inputs(161)) or (inputs(145)));
    layer0_outputs(5228) <= inputs(164);
    layer0_outputs(5229) <= (inputs(8)) and not (inputs(231));
    layer0_outputs(5230) <= not(inputs(228));
    layer0_outputs(5231) <= (inputs(30)) and (inputs(191));
    layer0_outputs(5232) <= not((inputs(156)) or (inputs(85)));
    layer0_outputs(5233) <= inputs(149);
    layer0_outputs(5234) <= '0';
    layer0_outputs(5235) <= not(inputs(254)) or (inputs(32));
    layer0_outputs(5236) <= (inputs(70)) or (inputs(18));
    layer0_outputs(5237) <= not((inputs(224)) xor (inputs(7)));
    layer0_outputs(5238) <= inputs(247);
    layer0_outputs(5239) <= (inputs(225)) or (inputs(136));
    layer0_outputs(5240) <= inputs(20);
    layer0_outputs(5241) <= (inputs(128)) or (inputs(20));
    layer0_outputs(5242) <= (inputs(85)) or (inputs(115));
    layer0_outputs(5243) <= not((inputs(114)) or (inputs(34)));
    layer0_outputs(5244) <= (inputs(129)) and (inputs(125));
    layer0_outputs(5245) <= not(inputs(29));
    layer0_outputs(5246) <= '0';
    layer0_outputs(5247) <= (inputs(92)) and (inputs(239));
    layer0_outputs(5248) <= not((inputs(238)) and (inputs(226)));
    layer0_outputs(5249) <= not(inputs(140));
    layer0_outputs(5250) <= inputs(123);
    layer0_outputs(5251) <= '1';
    layer0_outputs(5252) <= inputs(144);
    layer0_outputs(5253) <= (inputs(230)) or (inputs(157));
    layer0_outputs(5254) <= (inputs(244)) and (inputs(122));
    layer0_outputs(5255) <= (inputs(39)) or (inputs(190));
    layer0_outputs(5256) <= not((inputs(138)) or (inputs(112)));
    layer0_outputs(5257) <= '1';
    layer0_outputs(5258) <= not((inputs(204)) xor (inputs(186)));
    layer0_outputs(5259) <= inputs(44);
    layer0_outputs(5260) <= '1';
    layer0_outputs(5261) <= (inputs(20)) xor (inputs(210));
    layer0_outputs(5262) <= not((inputs(87)) or (inputs(1)));
    layer0_outputs(5263) <= not(inputs(94)) or (inputs(242));
    layer0_outputs(5264) <= (inputs(235)) and (inputs(9));
    layer0_outputs(5265) <= '0';
    layer0_outputs(5266) <= not(inputs(165));
    layer0_outputs(5267) <= '1';
    layer0_outputs(5268) <= (inputs(144)) or (inputs(188));
    layer0_outputs(5269) <= (inputs(143)) and not (inputs(99));
    layer0_outputs(5270) <= not((inputs(84)) xor (inputs(254)));
    layer0_outputs(5271) <= not(inputs(223)) or (inputs(135));
    layer0_outputs(5272) <= not((inputs(165)) or (inputs(199)));
    layer0_outputs(5273) <= (inputs(93)) and not (inputs(38));
    layer0_outputs(5274) <= not(inputs(168));
    layer0_outputs(5275) <= (inputs(217)) and (inputs(54));
    layer0_outputs(5276) <= (inputs(190)) or (inputs(127));
    layer0_outputs(5277) <= inputs(169);
    layer0_outputs(5278) <= inputs(77);
    layer0_outputs(5279) <= (inputs(223)) xor (inputs(70));
    layer0_outputs(5280) <= inputs(92);
    layer0_outputs(5281) <= '0';
    layer0_outputs(5282) <= not((inputs(201)) and (inputs(61)));
    layer0_outputs(5283) <= (inputs(192)) or (inputs(129));
    layer0_outputs(5284) <= not(inputs(215)) or (inputs(30));
    layer0_outputs(5285) <= not((inputs(145)) and (inputs(145)));
    layer0_outputs(5286) <= (inputs(7)) or (inputs(221));
    layer0_outputs(5287) <= not((inputs(67)) and (inputs(123)));
    layer0_outputs(5288) <= '0';
    layer0_outputs(5289) <= not(inputs(166));
    layer0_outputs(5290) <= (inputs(253)) or (inputs(218));
    layer0_outputs(5291) <= (inputs(242)) and (inputs(192));
    layer0_outputs(5292) <= not((inputs(97)) or (inputs(85)));
    layer0_outputs(5293) <= not(inputs(185));
    layer0_outputs(5294) <= '0';
    layer0_outputs(5295) <= (inputs(247)) and not (inputs(240));
    layer0_outputs(5296) <= not((inputs(218)) and (inputs(173)));
    layer0_outputs(5297) <= (inputs(72)) and not (inputs(13));
    layer0_outputs(5298) <= (inputs(120)) and not (inputs(98));
    layer0_outputs(5299) <= not((inputs(178)) or (inputs(183)));
    layer0_outputs(5300) <= not(inputs(252));
    layer0_outputs(5301) <= '1';
    layer0_outputs(5302) <= (inputs(214)) and (inputs(24));
    layer0_outputs(5303) <= inputs(179);
    layer0_outputs(5304) <= '0';
    layer0_outputs(5305) <= (inputs(161)) and not (inputs(197));
    layer0_outputs(5306) <= inputs(56);
    layer0_outputs(5307) <= not(inputs(173));
    layer0_outputs(5308) <= '1';
    layer0_outputs(5309) <= not((inputs(175)) and (inputs(144)));
    layer0_outputs(5310) <= not((inputs(167)) or (inputs(162)));
    layer0_outputs(5311) <= not(inputs(109));
    layer0_outputs(5312) <= inputs(230);
    layer0_outputs(5313) <= '0';
    layer0_outputs(5314) <= not(inputs(183));
    layer0_outputs(5315) <= (inputs(7)) and (inputs(18));
    layer0_outputs(5316) <= '0';
    layer0_outputs(5317) <= '1';
    layer0_outputs(5318) <= (inputs(164)) or (inputs(116));
    layer0_outputs(5319) <= not(inputs(79)) or (inputs(154));
    layer0_outputs(5320) <= (inputs(225)) and not (inputs(154));
    layer0_outputs(5321) <= not((inputs(163)) and (inputs(34)));
    layer0_outputs(5322) <= inputs(20);
    layer0_outputs(5323) <= not(inputs(177)) or (inputs(219));
    layer0_outputs(5324) <= inputs(191);
    layer0_outputs(5325) <= not(inputs(114));
    layer0_outputs(5326) <= not(inputs(25));
    layer0_outputs(5327) <= '1';
    layer0_outputs(5328) <= not(inputs(203));
    layer0_outputs(5329) <= inputs(24);
    layer0_outputs(5330) <= (inputs(174)) or (inputs(142));
    layer0_outputs(5331) <= not(inputs(40));
    layer0_outputs(5332) <= not((inputs(32)) or (inputs(75)));
    layer0_outputs(5333) <= inputs(221);
    layer0_outputs(5334) <= '0';
    layer0_outputs(5335) <= (inputs(241)) and not (inputs(81));
    layer0_outputs(5336) <= inputs(160);
    layer0_outputs(5337) <= (inputs(154)) xor (inputs(109));
    layer0_outputs(5338) <= (inputs(162)) and (inputs(247));
    layer0_outputs(5339) <= inputs(233);
    layer0_outputs(5340) <= not(inputs(95)) or (inputs(16));
    layer0_outputs(5341) <= not((inputs(160)) or (inputs(9)));
    layer0_outputs(5342) <= not(inputs(26)) or (inputs(163));
    layer0_outputs(5343) <= (inputs(177)) xor (inputs(145));
    layer0_outputs(5344) <= inputs(19);
    layer0_outputs(5345) <= not(inputs(123));
    layer0_outputs(5346) <= (inputs(255)) xor (inputs(153));
    layer0_outputs(5347) <= not((inputs(41)) and (inputs(150)));
    layer0_outputs(5348) <= '0';
    layer0_outputs(5349) <= '0';
    layer0_outputs(5350) <= (inputs(247)) or (inputs(226));
    layer0_outputs(5351) <= not((inputs(43)) or (inputs(251)));
    layer0_outputs(5352) <= (inputs(233)) and not (inputs(29));
    layer0_outputs(5353) <= (inputs(246)) or (inputs(227));
    layer0_outputs(5354) <= not(inputs(234)) or (inputs(85));
    layer0_outputs(5355) <= not(inputs(46));
    layer0_outputs(5356) <= not(inputs(104));
    layer0_outputs(5357) <= not(inputs(74)) or (inputs(240));
    layer0_outputs(5358) <= (inputs(70)) and (inputs(254));
    layer0_outputs(5359) <= not(inputs(93)) or (inputs(14));
    layer0_outputs(5360) <= (inputs(237)) and not (inputs(53));
    layer0_outputs(5361) <= '0';
    layer0_outputs(5362) <= '1';
    layer0_outputs(5363) <= '0';
    layer0_outputs(5364) <= not((inputs(160)) xor (inputs(219)));
    layer0_outputs(5365) <= inputs(201);
    layer0_outputs(5366) <= '0';
    layer0_outputs(5367) <= '0';
    layer0_outputs(5368) <= (inputs(125)) or (inputs(99));
    layer0_outputs(5369) <= not((inputs(255)) and (inputs(108)));
    layer0_outputs(5370) <= inputs(160);
    layer0_outputs(5371) <= inputs(199);
    layer0_outputs(5372) <= (inputs(169)) and not (inputs(227));
    layer0_outputs(5373) <= (inputs(200)) or (inputs(103));
    layer0_outputs(5374) <= (inputs(12)) or (inputs(133));
    layer0_outputs(5375) <= not(inputs(237));
    layer0_outputs(5376) <= '1';
    layer0_outputs(5377) <= inputs(247);
    layer0_outputs(5378) <= inputs(26);
    layer0_outputs(5379) <= not(inputs(100)) or (inputs(158));
    layer0_outputs(5380) <= (inputs(67)) and (inputs(26));
    layer0_outputs(5381) <= inputs(24);
    layer0_outputs(5382) <= not((inputs(137)) or (inputs(252)));
    layer0_outputs(5383) <= inputs(235);
    layer0_outputs(5384) <= not((inputs(145)) or (inputs(217)));
    layer0_outputs(5385) <= not((inputs(103)) or (inputs(142)));
    layer0_outputs(5386) <= not(inputs(34));
    layer0_outputs(5387) <= (inputs(192)) and not (inputs(162));
    layer0_outputs(5388) <= not(inputs(194));
    layer0_outputs(5389) <= '1';
    layer0_outputs(5390) <= not((inputs(216)) or (inputs(255)));
    layer0_outputs(5391) <= '0';
    layer0_outputs(5392) <= not(inputs(165));
    layer0_outputs(5393) <= not(inputs(84)) or (inputs(79));
    layer0_outputs(5394) <= not((inputs(204)) or (inputs(188)));
    layer0_outputs(5395) <= inputs(254);
    layer0_outputs(5396) <= '0';
    layer0_outputs(5397) <= '0';
    layer0_outputs(5398) <= (inputs(131)) and not (inputs(28));
    layer0_outputs(5399) <= (inputs(52)) and not (inputs(82));
    layer0_outputs(5400) <= inputs(175);
    layer0_outputs(5401) <= not((inputs(203)) or (inputs(106)));
    layer0_outputs(5402) <= '1';
    layer0_outputs(5403) <= inputs(53);
    layer0_outputs(5404) <= not(inputs(204));
    layer0_outputs(5405) <= not(inputs(207));
    layer0_outputs(5406) <= not(inputs(204)) or (inputs(248));
    layer0_outputs(5407) <= inputs(78);
    layer0_outputs(5408) <= not(inputs(178));
    layer0_outputs(5409) <= '1';
    layer0_outputs(5410) <= not(inputs(13));
    layer0_outputs(5411) <= not((inputs(239)) xor (inputs(18)));
    layer0_outputs(5412) <= inputs(24);
    layer0_outputs(5413) <= not((inputs(191)) xor (inputs(9)));
    layer0_outputs(5414) <= not((inputs(74)) and (inputs(236)));
    layer0_outputs(5415) <= not(inputs(114)) or (inputs(53));
    layer0_outputs(5416) <= inputs(152);
    layer0_outputs(5417) <= inputs(223);
    layer0_outputs(5418) <= (inputs(130)) or (inputs(206));
    layer0_outputs(5419) <= not((inputs(143)) and (inputs(121)));
    layer0_outputs(5420) <= (inputs(40)) and not (inputs(25));
    layer0_outputs(5421) <= not(inputs(170));
    layer0_outputs(5422) <= not(inputs(23));
    layer0_outputs(5423) <= '1';
    layer0_outputs(5424) <= not(inputs(41));
    layer0_outputs(5425) <= (inputs(134)) xor (inputs(112));
    layer0_outputs(5426) <= not((inputs(117)) or (inputs(4)));
    layer0_outputs(5427) <= '0';
    layer0_outputs(5428) <= not((inputs(197)) or (inputs(76)));
    layer0_outputs(5429) <= not((inputs(95)) and (inputs(249)));
    layer0_outputs(5430) <= (inputs(110)) and not (inputs(31));
    layer0_outputs(5431) <= inputs(119);
    layer0_outputs(5432) <= (inputs(142)) and not (inputs(252));
    layer0_outputs(5433) <= not(inputs(194));
    layer0_outputs(5434) <= not(inputs(27)) or (inputs(15));
    layer0_outputs(5435) <= '1';
    layer0_outputs(5436) <= inputs(60);
    layer0_outputs(5437) <= '1';
    layer0_outputs(5438) <= not(inputs(220));
    layer0_outputs(5439) <= inputs(181);
    layer0_outputs(5440) <= inputs(94);
    layer0_outputs(5441) <= not(inputs(151));
    layer0_outputs(5442) <= (inputs(98)) and not (inputs(40));
    layer0_outputs(5443) <= not((inputs(75)) or (inputs(128)));
    layer0_outputs(5444) <= '0';
    layer0_outputs(5445) <= not(inputs(71)) or (inputs(134));
    layer0_outputs(5446) <= (inputs(213)) and not (inputs(135));
    layer0_outputs(5447) <= not(inputs(130)) or (inputs(152));
    layer0_outputs(5448) <= (inputs(195)) and not (inputs(243));
    layer0_outputs(5449) <= (inputs(23)) or (inputs(61));
    layer0_outputs(5450) <= not(inputs(230));
    layer0_outputs(5451) <= '1';
    layer0_outputs(5452) <= not(inputs(152));
    layer0_outputs(5453) <= inputs(77);
    layer0_outputs(5454) <= not((inputs(190)) or (inputs(126)));
    layer0_outputs(5455) <= not((inputs(139)) xor (inputs(173)));
    layer0_outputs(5456) <= (inputs(165)) and (inputs(105));
    layer0_outputs(5457) <= not(inputs(26));
    layer0_outputs(5458) <= (inputs(234)) xor (inputs(79));
    layer0_outputs(5459) <= not(inputs(207));
    layer0_outputs(5460) <= (inputs(146)) and not (inputs(225));
    layer0_outputs(5461) <= inputs(234);
    layer0_outputs(5462) <= (inputs(9)) and not (inputs(218));
    layer0_outputs(5463) <= not((inputs(74)) or (inputs(116)));
    layer0_outputs(5464) <= not(inputs(50));
    layer0_outputs(5465) <= not(inputs(254)) or (inputs(12));
    layer0_outputs(5466) <= (inputs(73)) or (inputs(28));
    layer0_outputs(5467) <= (inputs(78)) and not (inputs(220));
    layer0_outputs(5468) <= '0';
    layer0_outputs(5469) <= (inputs(124)) and not (inputs(67));
    layer0_outputs(5470) <= '0';
    layer0_outputs(5471) <= (inputs(83)) or (inputs(96));
    layer0_outputs(5472) <= (inputs(14)) or (inputs(247));
    layer0_outputs(5473) <= (inputs(226)) or (inputs(206));
    layer0_outputs(5474) <= not(inputs(192));
    layer0_outputs(5475) <= not(inputs(249));
    layer0_outputs(5476) <= not(inputs(91));
    layer0_outputs(5477) <= (inputs(6)) xor (inputs(10));
    layer0_outputs(5478) <= (inputs(193)) and (inputs(125));
    layer0_outputs(5479) <= '0';
    layer0_outputs(5480) <= (inputs(91)) and not (inputs(213));
    layer0_outputs(5481) <= not((inputs(93)) or (inputs(112)));
    layer0_outputs(5482) <= inputs(226);
    layer0_outputs(5483) <= not(inputs(199)) or (inputs(43));
    layer0_outputs(5484) <= not(inputs(254)) or (inputs(49));
    layer0_outputs(5485) <= '1';
    layer0_outputs(5486) <= not((inputs(150)) and (inputs(198)));
    layer0_outputs(5487) <= '0';
    layer0_outputs(5488) <= inputs(211);
    layer0_outputs(5489) <= (inputs(203)) xor (inputs(250));
    layer0_outputs(5490) <= not((inputs(201)) or (inputs(48)));
    layer0_outputs(5491) <= not(inputs(9)) or (inputs(6));
    layer0_outputs(5492) <= not(inputs(220));
    layer0_outputs(5493) <= inputs(190);
    layer0_outputs(5494) <= (inputs(141)) and not (inputs(183));
    layer0_outputs(5495) <= '1';
    layer0_outputs(5496) <= (inputs(12)) and not (inputs(12));
    layer0_outputs(5497) <= inputs(56);
    layer0_outputs(5498) <= not(inputs(106)) or (inputs(59));
    layer0_outputs(5499) <= '0';
    layer0_outputs(5500) <= '1';
    layer0_outputs(5501) <= not(inputs(235)) or (inputs(130));
    layer0_outputs(5502) <= not(inputs(122));
    layer0_outputs(5503) <= inputs(99);
    layer0_outputs(5504) <= inputs(47);
    layer0_outputs(5505) <= '0';
    layer0_outputs(5506) <= '0';
    layer0_outputs(5507) <= not((inputs(175)) xor (inputs(92)));
    layer0_outputs(5508) <= not(inputs(26));
    layer0_outputs(5509) <= (inputs(76)) or (inputs(220));
    layer0_outputs(5510) <= not((inputs(147)) xor (inputs(99)));
    layer0_outputs(5511) <= not(inputs(194));
    layer0_outputs(5512) <= inputs(206);
    layer0_outputs(5513) <= (inputs(87)) and not (inputs(142));
    layer0_outputs(5514) <= '1';
    layer0_outputs(5515) <= inputs(199);
    layer0_outputs(5516) <= not(inputs(94));
    layer0_outputs(5517) <= inputs(215);
    layer0_outputs(5518) <= '0';
    layer0_outputs(5519) <= inputs(121);
    layer0_outputs(5520) <= (inputs(40)) and not (inputs(10));
    layer0_outputs(5521) <= inputs(178);
    layer0_outputs(5522) <= (inputs(225)) and not (inputs(155));
    layer0_outputs(5523) <= not((inputs(77)) or (inputs(71)));
    layer0_outputs(5524) <= inputs(101);
    layer0_outputs(5525) <= not(inputs(85));
    layer0_outputs(5526) <= not((inputs(126)) and (inputs(174)));
    layer0_outputs(5527) <= not(inputs(207)) or (inputs(76));
    layer0_outputs(5528) <= not(inputs(156));
    layer0_outputs(5529) <= '0';
    layer0_outputs(5530) <= '0';
    layer0_outputs(5531) <= (inputs(215)) and (inputs(174));
    layer0_outputs(5532) <= not(inputs(45));
    layer0_outputs(5533) <= inputs(116);
    layer0_outputs(5534) <= not(inputs(83));
    layer0_outputs(5535) <= (inputs(32)) or (inputs(49));
    layer0_outputs(5536) <= not((inputs(225)) and (inputs(12)));
    layer0_outputs(5537) <= not((inputs(120)) or (inputs(157)));
    layer0_outputs(5538) <= inputs(229);
    layer0_outputs(5539) <= not((inputs(251)) xor (inputs(173)));
    layer0_outputs(5540) <= not((inputs(20)) and (inputs(206)));
    layer0_outputs(5541) <= not((inputs(166)) or (inputs(30)));
    layer0_outputs(5542) <= not(inputs(129));
    layer0_outputs(5543) <= (inputs(252)) and not (inputs(141));
    layer0_outputs(5544) <= inputs(49);
    layer0_outputs(5545) <= not(inputs(33)) or (inputs(50));
    layer0_outputs(5546) <= not(inputs(171)) or (inputs(151));
    layer0_outputs(5547) <= not(inputs(115)) or (inputs(137));
    layer0_outputs(5548) <= '0';
    layer0_outputs(5549) <= not(inputs(93)) or (inputs(19));
    layer0_outputs(5550) <= not((inputs(129)) and (inputs(88)));
    layer0_outputs(5551) <= not(inputs(69)) or (inputs(58));
    layer0_outputs(5552) <= (inputs(222)) and (inputs(126));
    layer0_outputs(5553) <= not(inputs(255));
    layer0_outputs(5554) <= '1';
    layer0_outputs(5555) <= (inputs(14)) xor (inputs(46));
    layer0_outputs(5556) <= (inputs(163)) xor (inputs(198));
    layer0_outputs(5557) <= not(inputs(22));
    layer0_outputs(5558) <= not(inputs(241));
    layer0_outputs(5559) <= not(inputs(21));
    layer0_outputs(5560) <= not((inputs(189)) or (inputs(92)));
    layer0_outputs(5561) <= not((inputs(146)) or (inputs(72)));
    layer0_outputs(5562) <= (inputs(241)) xor (inputs(6));
    layer0_outputs(5563) <= (inputs(9)) and not (inputs(15));
    layer0_outputs(5564) <= inputs(195);
    layer0_outputs(5565) <= (inputs(111)) or (inputs(202));
    layer0_outputs(5566) <= '1';
    layer0_outputs(5567) <= not((inputs(3)) or (inputs(229)));
    layer0_outputs(5568) <= '0';
    layer0_outputs(5569) <= (inputs(127)) and not (inputs(54));
    layer0_outputs(5570) <= not(inputs(247)) or (inputs(103));
    layer0_outputs(5571) <= (inputs(123)) or (inputs(78));
    layer0_outputs(5572) <= inputs(176);
    layer0_outputs(5573) <= inputs(136);
    layer0_outputs(5574) <= (inputs(48)) and (inputs(31));
    layer0_outputs(5575) <= not(inputs(229));
    layer0_outputs(5576) <= (inputs(91)) and not (inputs(96));
    layer0_outputs(5577) <= not(inputs(106)) or (inputs(175));
    layer0_outputs(5578) <= '1';
    layer0_outputs(5579) <= not(inputs(16)) or (inputs(213));
    layer0_outputs(5580) <= not(inputs(60));
    layer0_outputs(5581) <= not((inputs(117)) and (inputs(97)));
    layer0_outputs(5582) <= (inputs(217)) and not (inputs(148));
    layer0_outputs(5583) <= '1';
    layer0_outputs(5584) <= (inputs(63)) xor (inputs(59));
    layer0_outputs(5585) <= '1';
    layer0_outputs(5586) <= not(inputs(88));
    layer0_outputs(5587) <= not((inputs(114)) or (inputs(44)));
    layer0_outputs(5588) <= (inputs(237)) and (inputs(55));
    layer0_outputs(5589) <= not(inputs(168)) or (inputs(104));
    layer0_outputs(5590) <= not(inputs(99));
    layer0_outputs(5591) <= '1';
    layer0_outputs(5592) <= not(inputs(49)) or (inputs(135));
    layer0_outputs(5593) <= (inputs(9)) and not (inputs(58));
    layer0_outputs(5594) <= not((inputs(129)) or (inputs(27)));
    layer0_outputs(5595) <= not((inputs(171)) or (inputs(64)));
    layer0_outputs(5596) <= (inputs(77)) or (inputs(88));
    layer0_outputs(5597) <= not((inputs(131)) xor (inputs(129)));
    layer0_outputs(5598) <= not((inputs(100)) and (inputs(95)));
    layer0_outputs(5599) <= not(inputs(48));
    layer0_outputs(5600) <= (inputs(145)) or (inputs(114));
    layer0_outputs(5601) <= inputs(166);
    layer0_outputs(5602) <= (inputs(207)) and not (inputs(61));
    layer0_outputs(5603) <= not(inputs(111));
    layer0_outputs(5604) <= not((inputs(226)) and (inputs(22)));
    layer0_outputs(5605) <= not(inputs(10)) or (inputs(226));
    layer0_outputs(5606) <= not((inputs(89)) or (inputs(57)));
    layer0_outputs(5607) <= not((inputs(3)) and (inputs(13)));
    layer0_outputs(5608) <= inputs(54);
    layer0_outputs(5609) <= inputs(9);
    layer0_outputs(5610) <= '1';
    layer0_outputs(5611) <= inputs(16);
    layer0_outputs(5612) <= not(inputs(49));
    layer0_outputs(5613) <= not((inputs(219)) or (inputs(160)));
    layer0_outputs(5614) <= '0';
    layer0_outputs(5615) <= not(inputs(188));
    layer0_outputs(5616) <= (inputs(114)) and not (inputs(41));
    layer0_outputs(5617) <= not(inputs(167)) or (inputs(185));
    layer0_outputs(5618) <= not(inputs(10));
    layer0_outputs(5619) <= not((inputs(155)) or (inputs(165)));
    layer0_outputs(5620) <= not((inputs(141)) xor (inputs(252)));
    layer0_outputs(5621) <= not(inputs(127)) or (inputs(172));
    layer0_outputs(5622) <= inputs(173);
    layer0_outputs(5623) <= inputs(105);
    layer0_outputs(5624) <= (inputs(131)) or (inputs(187));
    layer0_outputs(5625) <= not(inputs(90));
    layer0_outputs(5626) <= (inputs(254)) xor (inputs(0));
    layer0_outputs(5627) <= (inputs(224)) and (inputs(142));
    layer0_outputs(5628) <= not((inputs(43)) or (inputs(194)));
    layer0_outputs(5629) <= (inputs(181)) and not (inputs(141));
    layer0_outputs(5630) <= (inputs(20)) and not (inputs(9));
    layer0_outputs(5631) <= not(inputs(74));
    layer0_outputs(5632) <= '0';
    layer0_outputs(5633) <= not(inputs(109));
    layer0_outputs(5634) <= not(inputs(126));
    layer0_outputs(5635) <= (inputs(105)) and not (inputs(116));
    layer0_outputs(5636) <= '1';
    layer0_outputs(5637) <= inputs(59);
    layer0_outputs(5638) <= (inputs(147)) and not (inputs(222));
    layer0_outputs(5639) <= '0';
    layer0_outputs(5640) <= not((inputs(237)) and (inputs(72)));
    layer0_outputs(5641) <= not(inputs(107));
    layer0_outputs(5642) <= (inputs(137)) or (inputs(13));
    layer0_outputs(5643) <= (inputs(8)) and not (inputs(72));
    layer0_outputs(5644) <= (inputs(107)) or (inputs(141));
    layer0_outputs(5645) <= not(inputs(180));
    layer0_outputs(5646) <= not(inputs(129)) or (inputs(85));
    layer0_outputs(5647) <= '0';
    layer0_outputs(5648) <= '1';
    layer0_outputs(5649) <= not(inputs(214));
    layer0_outputs(5650) <= not(inputs(54)) or (inputs(5));
    layer0_outputs(5651) <= inputs(52);
    layer0_outputs(5652) <= (inputs(111)) and not (inputs(170));
    layer0_outputs(5653) <= not(inputs(35)) or (inputs(95));
    layer0_outputs(5654) <= inputs(227);
    layer0_outputs(5655) <= (inputs(56)) or (inputs(19));
    layer0_outputs(5656) <= (inputs(158)) and not (inputs(121));
    layer0_outputs(5657) <= inputs(201);
    layer0_outputs(5658) <= not(inputs(25));
    layer0_outputs(5659) <= not((inputs(91)) or (inputs(173)));
    layer0_outputs(5660) <= (inputs(30)) or (inputs(139));
    layer0_outputs(5661) <= '0';
    layer0_outputs(5662) <= (inputs(194)) and not (inputs(237));
    layer0_outputs(5663) <= inputs(12);
    layer0_outputs(5664) <= not(inputs(103)) or (inputs(81));
    layer0_outputs(5665) <= not(inputs(5)) or (inputs(240));
    layer0_outputs(5666) <= inputs(244);
    layer0_outputs(5667) <= (inputs(224)) and not (inputs(39));
    layer0_outputs(5668) <= not((inputs(132)) xor (inputs(151)));
    layer0_outputs(5669) <= inputs(60);
    layer0_outputs(5670) <= not(inputs(181));
    layer0_outputs(5671) <= not(inputs(160)) or (inputs(104));
    layer0_outputs(5672) <= (inputs(221)) and not (inputs(13));
    layer0_outputs(5673) <= not((inputs(94)) xor (inputs(0)));
    layer0_outputs(5674) <= '1';
    layer0_outputs(5675) <= (inputs(17)) or (inputs(249));
    layer0_outputs(5676) <= not(inputs(81));
    layer0_outputs(5677) <= not(inputs(99)) or (inputs(155));
    layer0_outputs(5678) <= (inputs(85)) and not (inputs(105));
    layer0_outputs(5679) <= '0';
    layer0_outputs(5680) <= inputs(89);
    layer0_outputs(5681) <= '1';
    layer0_outputs(5682) <= '0';
    layer0_outputs(5683) <= not(inputs(57));
    layer0_outputs(5684) <= '0';
    layer0_outputs(5685) <= inputs(72);
    layer0_outputs(5686) <= (inputs(202)) and not (inputs(66));
    layer0_outputs(5687) <= not((inputs(178)) or (inputs(125)));
    layer0_outputs(5688) <= not(inputs(126));
    layer0_outputs(5689) <= not(inputs(86)) or (inputs(70));
    layer0_outputs(5690) <= not(inputs(112));
    layer0_outputs(5691) <= (inputs(190)) and not (inputs(53));
    layer0_outputs(5692) <= '1';
    layer0_outputs(5693) <= '0';
    layer0_outputs(5694) <= not((inputs(191)) or (inputs(131)));
    layer0_outputs(5695) <= (inputs(134)) and not (inputs(252));
    layer0_outputs(5696) <= not(inputs(219)) or (inputs(166));
    layer0_outputs(5697) <= not(inputs(205));
    layer0_outputs(5698) <= not(inputs(115));
    layer0_outputs(5699) <= inputs(234);
    layer0_outputs(5700) <= (inputs(98)) and not (inputs(48));
    layer0_outputs(5701) <= inputs(131);
    layer0_outputs(5702) <= not(inputs(101));
    layer0_outputs(5703) <= inputs(249);
    layer0_outputs(5704) <= (inputs(172)) and (inputs(8));
    layer0_outputs(5705) <= '1';
    layer0_outputs(5706) <= not((inputs(58)) and (inputs(12)));
    layer0_outputs(5707) <= not((inputs(189)) or (inputs(81)));
    layer0_outputs(5708) <= inputs(42);
    layer0_outputs(5709) <= not(inputs(254));
    layer0_outputs(5710) <= not(inputs(213));
    layer0_outputs(5711) <= '1';
    layer0_outputs(5712) <= not(inputs(58)) or (inputs(74));
    layer0_outputs(5713) <= (inputs(170)) or (inputs(236));
    layer0_outputs(5714) <= not(inputs(86));
    layer0_outputs(5715) <= not(inputs(170));
    layer0_outputs(5716) <= not((inputs(170)) xor (inputs(98)));
    layer0_outputs(5717) <= (inputs(223)) or (inputs(9));
    layer0_outputs(5718) <= not(inputs(8)) or (inputs(235));
    layer0_outputs(5719) <= (inputs(139)) and (inputs(83));
    layer0_outputs(5720) <= inputs(50);
    layer0_outputs(5721) <= not(inputs(19));
    layer0_outputs(5722) <= inputs(111);
    layer0_outputs(5723) <= not(inputs(158));
    layer0_outputs(5724) <= inputs(161);
    layer0_outputs(5725) <= (inputs(155)) or (inputs(216));
    layer0_outputs(5726) <= inputs(217);
    layer0_outputs(5727) <= not(inputs(145)) or (inputs(41));
    layer0_outputs(5728) <= (inputs(126)) and (inputs(229));
    layer0_outputs(5729) <= '1';
    layer0_outputs(5730) <= not((inputs(99)) or (inputs(78)));
    layer0_outputs(5731) <= not(inputs(148));
    layer0_outputs(5732) <= '1';
    layer0_outputs(5733) <= inputs(237);
    layer0_outputs(5734) <= not(inputs(101)) or (inputs(17));
    layer0_outputs(5735) <= not((inputs(226)) and (inputs(232)));
    layer0_outputs(5736) <= (inputs(127)) and (inputs(84));
    layer0_outputs(5737) <= not(inputs(60));
    layer0_outputs(5738) <= (inputs(221)) and not (inputs(64));
    layer0_outputs(5739) <= (inputs(105)) and not (inputs(62));
    layer0_outputs(5740) <= (inputs(118)) xor (inputs(147));
    layer0_outputs(5741) <= not(inputs(216)) or (inputs(59));
    layer0_outputs(5742) <= '1';
    layer0_outputs(5743) <= not(inputs(120));
    layer0_outputs(5744) <= (inputs(122)) xor (inputs(103));
    layer0_outputs(5745) <= '0';
    layer0_outputs(5746) <= inputs(94);
    layer0_outputs(5747) <= not((inputs(45)) or (inputs(69)));
    layer0_outputs(5748) <= (inputs(59)) and (inputs(182));
    layer0_outputs(5749) <= not((inputs(245)) xor (inputs(208)));
    layer0_outputs(5750) <= inputs(72);
    layer0_outputs(5751) <= (inputs(168)) and not (inputs(74));
    layer0_outputs(5752) <= not(inputs(184)) or (inputs(228));
    layer0_outputs(5753) <= (inputs(57)) and (inputs(71));
    layer0_outputs(5754) <= (inputs(144)) or (inputs(99));
    layer0_outputs(5755) <= not(inputs(21));
    layer0_outputs(5756) <= not(inputs(207));
    layer0_outputs(5757) <= inputs(184);
    layer0_outputs(5758) <= '0';
    layer0_outputs(5759) <= not(inputs(24));
    layer0_outputs(5760) <= '1';
    layer0_outputs(5761) <= '0';
    layer0_outputs(5762) <= not(inputs(169));
    layer0_outputs(5763) <= (inputs(185)) and not (inputs(135));
    layer0_outputs(5764) <= not(inputs(25)) or (inputs(86));
    layer0_outputs(5765) <= not(inputs(223));
    layer0_outputs(5766) <= '1';
    layer0_outputs(5767) <= not(inputs(238));
    layer0_outputs(5768) <= not(inputs(111)) or (inputs(182));
    layer0_outputs(5769) <= (inputs(89)) and not (inputs(182));
    layer0_outputs(5770) <= not(inputs(126)) or (inputs(136));
    layer0_outputs(5771) <= not((inputs(149)) xor (inputs(163)));
    layer0_outputs(5772) <= (inputs(236)) and (inputs(168));
    layer0_outputs(5773) <= not(inputs(115));
    layer0_outputs(5774) <= '1';
    layer0_outputs(5775) <= '0';
    layer0_outputs(5776) <= '1';
    layer0_outputs(5777) <= (inputs(197)) and not (inputs(131));
    layer0_outputs(5778) <= not((inputs(116)) or (inputs(177)));
    layer0_outputs(5779) <= inputs(41);
    layer0_outputs(5780) <= inputs(251);
    layer0_outputs(5781) <= (inputs(27)) and not (inputs(50));
    layer0_outputs(5782) <= '0';
    layer0_outputs(5783) <= not(inputs(104));
    layer0_outputs(5784) <= not(inputs(97));
    layer0_outputs(5785) <= not(inputs(130)) or (inputs(138));
    layer0_outputs(5786) <= inputs(97);
    layer0_outputs(5787) <= inputs(95);
    layer0_outputs(5788) <= '1';
    layer0_outputs(5789) <= '0';
    layer0_outputs(5790) <= (inputs(12)) or (inputs(255));
    layer0_outputs(5791) <= inputs(174);
    layer0_outputs(5792) <= not((inputs(207)) or (inputs(229)));
    layer0_outputs(5793) <= not(inputs(92)) or (inputs(29));
    layer0_outputs(5794) <= '1';
    layer0_outputs(5795) <= not((inputs(239)) and (inputs(87)));
    layer0_outputs(5796) <= inputs(173);
    layer0_outputs(5797) <= not((inputs(134)) or (inputs(13)));
    layer0_outputs(5798) <= inputs(135);
    layer0_outputs(5799) <= inputs(80);
    layer0_outputs(5800) <= not((inputs(74)) and (inputs(9)));
    layer0_outputs(5801) <= (inputs(34)) and (inputs(232));
    layer0_outputs(5802) <= not(inputs(105));
    layer0_outputs(5803) <= (inputs(69)) and not (inputs(32));
    layer0_outputs(5804) <= not(inputs(164));
    layer0_outputs(5805) <= not(inputs(50));
    layer0_outputs(5806) <= '1';
    layer0_outputs(5807) <= not((inputs(187)) or (inputs(217)));
    layer0_outputs(5808) <= (inputs(75)) or (inputs(60));
    layer0_outputs(5809) <= (inputs(238)) and (inputs(141));
    layer0_outputs(5810) <= inputs(25);
    layer0_outputs(5811) <= not(inputs(222));
    layer0_outputs(5812) <= (inputs(186)) or (inputs(217));
    layer0_outputs(5813) <= not(inputs(70));
    layer0_outputs(5814) <= (inputs(26)) xor (inputs(191));
    layer0_outputs(5815) <= (inputs(99)) and not (inputs(191));
    layer0_outputs(5816) <= (inputs(3)) or (inputs(209));
    layer0_outputs(5817) <= (inputs(31)) or (inputs(39));
    layer0_outputs(5818) <= not((inputs(175)) or (inputs(69)));
    layer0_outputs(5819) <= (inputs(106)) and not (inputs(1));
    layer0_outputs(5820) <= '0';
    layer0_outputs(5821) <= inputs(180);
    layer0_outputs(5822) <= not((inputs(77)) or (inputs(92)));
    layer0_outputs(5823) <= '0';
    layer0_outputs(5824) <= (inputs(119)) and (inputs(250));
    layer0_outputs(5825) <= not(inputs(62));
    layer0_outputs(5826) <= not(inputs(223));
    layer0_outputs(5827) <= not(inputs(224)) or (inputs(115));
    layer0_outputs(5828) <= '0';
    layer0_outputs(5829) <= inputs(173);
    layer0_outputs(5830) <= inputs(89);
    layer0_outputs(5831) <= (inputs(175)) or (inputs(229));
    layer0_outputs(5832) <= not((inputs(3)) or (inputs(77)));
    layer0_outputs(5833) <= inputs(42);
    layer0_outputs(5834) <= not((inputs(99)) or (inputs(51)));
    layer0_outputs(5835) <= (inputs(2)) or (inputs(23));
    layer0_outputs(5836) <= not((inputs(2)) or (inputs(92)));
    layer0_outputs(5837) <= '0';
    layer0_outputs(5838) <= '1';
    layer0_outputs(5839) <= not(inputs(62)) or (inputs(174));
    layer0_outputs(5840) <= not((inputs(38)) or (inputs(77)));
    layer0_outputs(5841) <= not(inputs(22));
    layer0_outputs(5842) <= not((inputs(212)) xor (inputs(175)));
    layer0_outputs(5843) <= inputs(121);
    layer0_outputs(5844) <= '0';
    layer0_outputs(5845) <= '0';
    layer0_outputs(5846) <= '1';
    layer0_outputs(5847) <= not(inputs(67));
    layer0_outputs(5848) <= (inputs(47)) and (inputs(244));
    layer0_outputs(5849) <= not(inputs(165)) or (inputs(251));
    layer0_outputs(5850) <= (inputs(112)) or (inputs(117));
    layer0_outputs(5851) <= not(inputs(64));
    layer0_outputs(5852) <= (inputs(170)) and not (inputs(14));
    layer0_outputs(5853) <= inputs(145);
    layer0_outputs(5854) <= '1';
    layer0_outputs(5855) <= inputs(138);
    layer0_outputs(5856) <= inputs(166);
    layer0_outputs(5857) <= not((inputs(115)) xor (inputs(100)));
    layer0_outputs(5858) <= inputs(82);
    layer0_outputs(5859) <= inputs(217);
    layer0_outputs(5860) <= inputs(250);
    layer0_outputs(5861) <= inputs(244);
    layer0_outputs(5862) <= (inputs(93)) and not (inputs(67));
    layer0_outputs(5863) <= '0';
    layer0_outputs(5864) <= not(inputs(244)) or (inputs(75));
    layer0_outputs(5865) <= '0';
    layer0_outputs(5866) <= (inputs(174)) and (inputs(7));
    layer0_outputs(5867) <= '0';
    layer0_outputs(5868) <= not(inputs(233)) or (inputs(244));
    layer0_outputs(5869) <= not((inputs(37)) or (inputs(239)));
    layer0_outputs(5870) <= inputs(218);
    layer0_outputs(5871) <= not(inputs(192));
    layer0_outputs(5872) <= not(inputs(23));
    layer0_outputs(5873) <= '1';
    layer0_outputs(5874) <= (inputs(159)) or (inputs(228));
    layer0_outputs(5875) <= inputs(157);
    layer0_outputs(5876) <= (inputs(16)) and not (inputs(96));
    layer0_outputs(5877) <= not(inputs(39));
    layer0_outputs(5878) <= not(inputs(85));
    layer0_outputs(5879) <= not(inputs(73)) or (inputs(139));
    layer0_outputs(5880) <= not((inputs(214)) or (inputs(254)));
    layer0_outputs(5881) <= (inputs(101)) and not (inputs(46));
    layer0_outputs(5882) <= not(inputs(244));
    layer0_outputs(5883) <= '1';
    layer0_outputs(5884) <= not(inputs(134)) or (inputs(47));
    layer0_outputs(5885) <= not(inputs(174));
    layer0_outputs(5886) <= inputs(178);
    layer0_outputs(5887) <= not(inputs(253)) or (inputs(198));
    layer0_outputs(5888) <= not(inputs(214));
    layer0_outputs(5889) <= (inputs(218)) and (inputs(228));
    layer0_outputs(5890) <= not(inputs(82));
    layer0_outputs(5891) <= inputs(95);
    layer0_outputs(5892) <= inputs(154);
    layer0_outputs(5893) <= '1';
    layer0_outputs(5894) <= '1';
    layer0_outputs(5895) <= inputs(173);
    layer0_outputs(5896) <= inputs(12);
    layer0_outputs(5897) <= not(inputs(142));
    layer0_outputs(5898) <= (inputs(92)) and (inputs(146));
    layer0_outputs(5899) <= inputs(234);
    layer0_outputs(5900) <= (inputs(18)) xor (inputs(236));
    layer0_outputs(5901) <= not(inputs(154));
    layer0_outputs(5902) <= not(inputs(236)) or (inputs(123));
    layer0_outputs(5903) <= inputs(110);
    layer0_outputs(5904) <= (inputs(117)) and not (inputs(11));
    layer0_outputs(5905) <= (inputs(195)) or (inputs(65));
    layer0_outputs(5906) <= not(inputs(109)) or (inputs(80));
    layer0_outputs(5907) <= inputs(101);
    layer0_outputs(5908) <= not((inputs(161)) xor (inputs(180)));
    layer0_outputs(5909) <= '1';
    layer0_outputs(5910) <= not(inputs(128)) or (inputs(153));
    layer0_outputs(5911) <= not(inputs(31)) or (inputs(250));
    layer0_outputs(5912) <= not((inputs(200)) or (inputs(221)));
    layer0_outputs(5913) <= not(inputs(76));
    layer0_outputs(5914) <= inputs(154);
    layer0_outputs(5915) <= not(inputs(93));
    layer0_outputs(5916) <= (inputs(191)) and not (inputs(250));
    layer0_outputs(5917) <= (inputs(37)) and not (inputs(175));
    layer0_outputs(5918) <= not(inputs(251)) or (inputs(203));
    layer0_outputs(5919) <= '1';
    layer0_outputs(5920) <= (inputs(90)) and not (inputs(143));
    layer0_outputs(5921) <= (inputs(141)) or (inputs(142));
    layer0_outputs(5922) <= '0';
    layer0_outputs(5923) <= not((inputs(68)) and (inputs(18)));
    layer0_outputs(5924) <= not(inputs(225)) or (inputs(217));
    layer0_outputs(5925) <= inputs(214);
    layer0_outputs(5926) <= not(inputs(177)) or (inputs(125));
    layer0_outputs(5927) <= not((inputs(120)) xor (inputs(123)));
    layer0_outputs(5928) <= (inputs(247)) or (inputs(23));
    layer0_outputs(5929) <= inputs(76);
    layer0_outputs(5930) <= '1';
    layer0_outputs(5931) <= not(inputs(222)) or (inputs(108));
    layer0_outputs(5932) <= inputs(100);
    layer0_outputs(5933) <= (inputs(97)) and not (inputs(75));
    layer0_outputs(5934) <= inputs(141);
    layer0_outputs(5935) <= '1';
    layer0_outputs(5936) <= not(inputs(35)) or (inputs(251));
    layer0_outputs(5937) <= inputs(146);
    layer0_outputs(5938) <= '1';
    layer0_outputs(5939) <= not(inputs(28));
    layer0_outputs(5940) <= not((inputs(60)) and (inputs(175)));
    layer0_outputs(5941) <= '0';
    layer0_outputs(5942) <= (inputs(249)) or (inputs(155));
    layer0_outputs(5943) <= not((inputs(43)) or (inputs(241)));
    layer0_outputs(5944) <= '1';
    layer0_outputs(5945) <= not(inputs(136)) or (inputs(211));
    layer0_outputs(5946) <= inputs(147);
    layer0_outputs(5947) <= inputs(90);
    layer0_outputs(5948) <= (inputs(30)) and not (inputs(60));
    layer0_outputs(5949) <= inputs(121);
    layer0_outputs(5950) <= not(inputs(62));
    layer0_outputs(5951) <= (inputs(131)) and not (inputs(122));
    layer0_outputs(5952) <= (inputs(29)) and not (inputs(130));
    layer0_outputs(5953) <= '1';
    layer0_outputs(5954) <= '0';
    layer0_outputs(5955) <= not((inputs(247)) or (inputs(190)));
    layer0_outputs(5956) <= not((inputs(187)) xor (inputs(2)));
    layer0_outputs(5957) <= inputs(197);
    layer0_outputs(5958) <= (inputs(246)) or (inputs(241));
    layer0_outputs(5959) <= not((inputs(213)) xor (inputs(79)));
    layer0_outputs(5960) <= not((inputs(222)) or (inputs(206)));
    layer0_outputs(5961) <= not(inputs(116)) or (inputs(16));
    layer0_outputs(5962) <= (inputs(33)) and not (inputs(145));
    layer0_outputs(5963) <= not(inputs(54)) or (inputs(191));
    layer0_outputs(5964) <= (inputs(18)) xor (inputs(129));
    layer0_outputs(5965) <= not(inputs(190)) or (inputs(38));
    layer0_outputs(5966) <= not((inputs(239)) or (inputs(187)));
    layer0_outputs(5967) <= '1';
    layer0_outputs(5968) <= not(inputs(194)) or (inputs(56));
    layer0_outputs(5969) <= '1';
    layer0_outputs(5970) <= not((inputs(217)) xor (inputs(170)));
    layer0_outputs(5971) <= not((inputs(208)) or (inputs(136)));
    layer0_outputs(5972) <= inputs(204);
    layer0_outputs(5973) <= (inputs(154)) or (inputs(111));
    layer0_outputs(5974) <= '0';
    layer0_outputs(5975) <= (inputs(146)) and (inputs(244));
    layer0_outputs(5976) <= (inputs(189)) and not (inputs(184));
    layer0_outputs(5977) <= not(inputs(117)) or (inputs(139));
    layer0_outputs(5978) <= not(inputs(105));
    layer0_outputs(5979) <= (inputs(111)) and not (inputs(34));
    layer0_outputs(5980) <= not(inputs(54)) or (inputs(251));
    layer0_outputs(5981) <= not(inputs(209));
    layer0_outputs(5982) <= (inputs(234)) and not (inputs(246));
    layer0_outputs(5983) <= inputs(168);
    layer0_outputs(5984) <= not((inputs(126)) and (inputs(19)));
    layer0_outputs(5985) <= inputs(149);
    layer0_outputs(5986) <= not(inputs(144)) or (inputs(57));
    layer0_outputs(5987) <= not(inputs(5)) or (inputs(10));
    layer0_outputs(5988) <= not(inputs(149)) or (inputs(79));
    layer0_outputs(5989) <= (inputs(171)) and (inputs(163));
    layer0_outputs(5990) <= (inputs(203)) xor (inputs(222));
    layer0_outputs(5991) <= not(inputs(107));
    layer0_outputs(5992) <= not(inputs(8));
    layer0_outputs(5993) <= not((inputs(192)) and (inputs(32)));
    layer0_outputs(5994) <= not((inputs(37)) or (inputs(20)));
    layer0_outputs(5995) <= not(inputs(33));
    layer0_outputs(5996) <= not((inputs(76)) xor (inputs(210)));
    layer0_outputs(5997) <= (inputs(55)) and not (inputs(237));
    layer0_outputs(5998) <= inputs(44);
    layer0_outputs(5999) <= not(inputs(21));
    layer0_outputs(6000) <= inputs(156);
    layer0_outputs(6001) <= not(inputs(34));
    layer0_outputs(6002) <= (inputs(248)) and not (inputs(208));
    layer0_outputs(6003) <= inputs(182);
    layer0_outputs(6004) <= not(inputs(136)) or (inputs(148));
    layer0_outputs(6005) <= inputs(58);
    layer0_outputs(6006) <= inputs(255);
    layer0_outputs(6007) <= not((inputs(246)) or (inputs(229)));
    layer0_outputs(6008) <= not((inputs(187)) or (inputs(27)));
    layer0_outputs(6009) <= (inputs(213)) and (inputs(253));
    layer0_outputs(6010) <= not((inputs(124)) and (inputs(112)));
    layer0_outputs(6011) <= not((inputs(127)) xor (inputs(3)));
    layer0_outputs(6012) <= inputs(141);
    layer0_outputs(6013) <= not((inputs(96)) and (inputs(22)));
    layer0_outputs(6014) <= inputs(21);
    layer0_outputs(6015) <= not(inputs(31)) or (inputs(214));
    layer0_outputs(6016) <= not(inputs(148));
    layer0_outputs(6017) <= '1';
    layer0_outputs(6018) <= (inputs(63)) xor (inputs(242));
    layer0_outputs(6019) <= (inputs(79)) and (inputs(150));
    layer0_outputs(6020) <= not((inputs(141)) or (inputs(14)));
    layer0_outputs(6021) <= not((inputs(109)) and (inputs(61)));
    layer0_outputs(6022) <= (inputs(52)) xor (inputs(49));
    layer0_outputs(6023) <= '0';
    layer0_outputs(6024) <= not(inputs(116));
    layer0_outputs(6025) <= not(inputs(175)) or (inputs(250));
    layer0_outputs(6026) <= (inputs(185)) or (inputs(186));
    layer0_outputs(6027) <= inputs(77);
    layer0_outputs(6028) <= (inputs(29)) or (inputs(90));
    layer0_outputs(6029) <= not(inputs(211)) or (inputs(205));
    layer0_outputs(6030) <= (inputs(1)) or (inputs(240));
    layer0_outputs(6031) <= (inputs(248)) or (inputs(70));
    layer0_outputs(6032) <= '0';
    layer0_outputs(6033) <= (inputs(190)) or (inputs(193));
    layer0_outputs(6034) <= '1';
    layer0_outputs(6035) <= '0';
    layer0_outputs(6036) <= not(inputs(254));
    layer0_outputs(6037) <= not(inputs(137));
    layer0_outputs(6038) <= not(inputs(140)) or (inputs(44));
    layer0_outputs(6039) <= (inputs(127)) and (inputs(34));
    layer0_outputs(6040) <= (inputs(174)) and not (inputs(251));
    layer0_outputs(6041) <= (inputs(91)) and not (inputs(57));
    layer0_outputs(6042) <= inputs(231);
    layer0_outputs(6043) <= '0';
    layer0_outputs(6044) <= not((inputs(142)) xor (inputs(35)));
    layer0_outputs(6045) <= not((inputs(166)) or (inputs(37)));
    layer0_outputs(6046) <= inputs(78);
    layer0_outputs(6047) <= (inputs(182)) and not (inputs(223));
    layer0_outputs(6048) <= inputs(156);
    layer0_outputs(6049) <= '1';
    layer0_outputs(6050) <= (inputs(233)) xor (inputs(63));
    layer0_outputs(6051) <= (inputs(228)) and not (inputs(41));
    layer0_outputs(6052) <= '0';
    layer0_outputs(6053) <= not((inputs(0)) and (inputs(73)));
    layer0_outputs(6054) <= not((inputs(16)) or (inputs(168)));
    layer0_outputs(6055) <= (inputs(118)) and not (inputs(226));
    layer0_outputs(6056) <= not((inputs(133)) and (inputs(179)));
    layer0_outputs(6057) <= not(inputs(52)) or (inputs(160));
    layer0_outputs(6058) <= not(inputs(189)) or (inputs(232));
    layer0_outputs(6059) <= (inputs(228)) or (inputs(48));
    layer0_outputs(6060) <= not((inputs(10)) and (inputs(212)));
    layer0_outputs(6061) <= (inputs(30)) and not (inputs(193));
    layer0_outputs(6062) <= '1';
    layer0_outputs(6063) <= not(inputs(138));
    layer0_outputs(6064) <= not(inputs(155)) or (inputs(70));
    layer0_outputs(6065) <= (inputs(75)) or (inputs(234));
    layer0_outputs(6066) <= not((inputs(143)) xor (inputs(219)));
    layer0_outputs(6067) <= (inputs(82)) or (inputs(38));
    layer0_outputs(6068) <= not((inputs(3)) or (inputs(205)));
    layer0_outputs(6069) <= '0';
    layer0_outputs(6070) <= (inputs(119)) xor (inputs(17));
    layer0_outputs(6071) <= inputs(134);
    layer0_outputs(6072) <= not(inputs(110)) or (inputs(254));
    layer0_outputs(6073) <= not((inputs(129)) and (inputs(246)));
    layer0_outputs(6074) <= not(inputs(35));
    layer0_outputs(6075) <= not((inputs(244)) xor (inputs(199)));
    layer0_outputs(6076) <= not((inputs(17)) or (inputs(120)));
    layer0_outputs(6077) <= '1';
    layer0_outputs(6078) <= not((inputs(190)) xor (inputs(237)));
    layer0_outputs(6079) <= inputs(121);
    layer0_outputs(6080) <= (inputs(103)) and not (inputs(237));
    layer0_outputs(6081) <= not(inputs(122)) or (inputs(173));
    layer0_outputs(6082) <= (inputs(177)) or (inputs(239));
    layer0_outputs(6083) <= not(inputs(82)) or (inputs(43));
    layer0_outputs(6084) <= (inputs(100)) xor (inputs(102));
    layer0_outputs(6085) <= inputs(77);
    layer0_outputs(6086) <= inputs(102);
    layer0_outputs(6087) <= not((inputs(205)) or (inputs(22)));
    layer0_outputs(6088) <= '0';
    layer0_outputs(6089) <= not((inputs(194)) or (inputs(145)));
    layer0_outputs(6090) <= (inputs(9)) and (inputs(102));
    layer0_outputs(6091) <= not(inputs(138)) or (inputs(133));
    layer0_outputs(6092) <= (inputs(253)) xor (inputs(114));
    layer0_outputs(6093) <= (inputs(243)) xor (inputs(227));
    layer0_outputs(6094) <= not(inputs(130));
    layer0_outputs(6095) <= inputs(233);
    layer0_outputs(6096) <= not((inputs(143)) or (inputs(87)));
    layer0_outputs(6097) <= (inputs(22)) and (inputs(128));
    layer0_outputs(6098) <= inputs(174);
    layer0_outputs(6099) <= not(inputs(33)) or (inputs(191));
    layer0_outputs(6100) <= not(inputs(126)) or (inputs(169));
    layer0_outputs(6101) <= not((inputs(226)) or (inputs(104)));
    layer0_outputs(6102) <= (inputs(129)) and (inputs(152));
    layer0_outputs(6103) <= inputs(187);
    layer0_outputs(6104) <= '1';
    layer0_outputs(6105) <= not(inputs(91)) or (inputs(56));
    layer0_outputs(6106) <= not(inputs(185)) or (inputs(20));
    layer0_outputs(6107) <= (inputs(37)) xor (inputs(34));
    layer0_outputs(6108) <= not(inputs(121)) or (inputs(253));
    layer0_outputs(6109) <= '0';
    layer0_outputs(6110) <= (inputs(167)) or (inputs(150));
    layer0_outputs(6111) <= inputs(116);
    layer0_outputs(6112) <= not(inputs(255)) or (inputs(89));
    layer0_outputs(6113) <= not(inputs(68));
    layer0_outputs(6114) <= not(inputs(50)) or (inputs(161));
    layer0_outputs(6115) <= not(inputs(243));
    layer0_outputs(6116) <= inputs(178);
    layer0_outputs(6117) <= not((inputs(16)) or (inputs(21)));
    layer0_outputs(6118) <= not(inputs(130));
    layer0_outputs(6119) <= not(inputs(147));
    layer0_outputs(6120) <= '1';
    layer0_outputs(6121) <= (inputs(180)) and (inputs(56));
    layer0_outputs(6122) <= not(inputs(94));
    layer0_outputs(6123) <= '0';
    layer0_outputs(6124) <= not(inputs(16)) or (inputs(199));
    layer0_outputs(6125) <= not((inputs(139)) or (inputs(217)));
    layer0_outputs(6126) <= '0';
    layer0_outputs(6127) <= not((inputs(116)) or (inputs(199)));
    layer0_outputs(6128) <= not((inputs(10)) xor (inputs(7)));
    layer0_outputs(6129) <= '0';
    layer0_outputs(6130) <= not((inputs(158)) and (inputs(125)));
    layer0_outputs(6131) <= (inputs(73)) and (inputs(94));
    layer0_outputs(6132) <= (inputs(215)) and (inputs(1));
    layer0_outputs(6133) <= '1';
    layer0_outputs(6134) <= '1';
    layer0_outputs(6135) <= (inputs(252)) or (inputs(202));
    layer0_outputs(6136) <= not(inputs(63));
    layer0_outputs(6137) <= '1';
    layer0_outputs(6138) <= not(inputs(201)) or (inputs(86));
    layer0_outputs(6139) <= inputs(106);
    layer0_outputs(6140) <= not(inputs(176)) or (inputs(59));
    layer0_outputs(6141) <= (inputs(228)) and not (inputs(103));
    layer0_outputs(6142) <= '1';
    layer0_outputs(6143) <= not(inputs(220));
    layer0_outputs(6144) <= (inputs(233)) and not (inputs(79));
    layer0_outputs(6145) <= not((inputs(143)) xor (inputs(142)));
    layer0_outputs(6146) <= not(inputs(40));
    layer0_outputs(6147) <= not(inputs(190));
    layer0_outputs(6148) <= inputs(95);
    layer0_outputs(6149) <= (inputs(33)) and (inputs(84));
    layer0_outputs(6150) <= not(inputs(235));
    layer0_outputs(6151) <= not(inputs(145));
    layer0_outputs(6152) <= (inputs(35)) and (inputs(6));
    layer0_outputs(6153) <= not(inputs(71));
    layer0_outputs(6154) <= (inputs(198)) and not (inputs(63));
    layer0_outputs(6155) <= (inputs(176)) xor (inputs(50));
    layer0_outputs(6156) <= '0';
    layer0_outputs(6157) <= not(inputs(253)) or (inputs(81));
    layer0_outputs(6158) <= (inputs(84)) and (inputs(121));
    layer0_outputs(6159) <= (inputs(46)) and (inputs(121));
    layer0_outputs(6160) <= (inputs(219)) and not (inputs(158));
    layer0_outputs(6161) <= '1';
    layer0_outputs(6162) <= (inputs(65)) and not (inputs(238));
    layer0_outputs(6163) <= '1';
    layer0_outputs(6164) <= not((inputs(116)) or (inputs(131)));
    layer0_outputs(6165) <= '1';
    layer0_outputs(6166) <= '1';
    layer0_outputs(6167) <= inputs(24);
    layer0_outputs(6168) <= not(inputs(21)) or (inputs(113));
    layer0_outputs(6169) <= not(inputs(128));
    layer0_outputs(6170) <= (inputs(47)) and not (inputs(123));
    layer0_outputs(6171) <= not(inputs(193));
    layer0_outputs(6172) <= inputs(247);
    layer0_outputs(6173) <= (inputs(25)) and not (inputs(193));
    layer0_outputs(6174) <= inputs(119);
    layer0_outputs(6175) <= (inputs(33)) and not (inputs(251));
    layer0_outputs(6176) <= (inputs(128)) or (inputs(148));
    layer0_outputs(6177) <= (inputs(90)) and not (inputs(96));
    layer0_outputs(6178) <= inputs(222);
    layer0_outputs(6179) <= (inputs(174)) or (inputs(229));
    layer0_outputs(6180) <= '0';
    layer0_outputs(6181) <= not((inputs(204)) or (inputs(2)));
    layer0_outputs(6182) <= (inputs(107)) or (inputs(126));
    layer0_outputs(6183) <= (inputs(152)) and not (inputs(160));
    layer0_outputs(6184) <= not(inputs(27));
    layer0_outputs(6185) <= inputs(181);
    layer0_outputs(6186) <= (inputs(119)) xor (inputs(12));
    layer0_outputs(6187) <= not((inputs(3)) or (inputs(190)));
    layer0_outputs(6188) <= '0';
    layer0_outputs(6189) <= not((inputs(240)) or (inputs(81)));
    layer0_outputs(6190) <= not(inputs(251)) or (inputs(169));
    layer0_outputs(6191) <= (inputs(146)) and not (inputs(149));
    layer0_outputs(6192) <= not(inputs(254)) or (inputs(121));
    layer0_outputs(6193) <= (inputs(112)) and not (inputs(152));
    layer0_outputs(6194) <= (inputs(134)) and not (inputs(143));
    layer0_outputs(6195) <= not(inputs(66)) or (inputs(176));
    layer0_outputs(6196) <= (inputs(206)) and not (inputs(110));
    layer0_outputs(6197) <= (inputs(197)) xor (inputs(19));
    layer0_outputs(6198) <= '1';
    layer0_outputs(6199) <= not(inputs(241)) or (inputs(204));
    layer0_outputs(6200) <= not(inputs(53));
    layer0_outputs(6201) <= not(inputs(31)) or (inputs(82));
    layer0_outputs(6202) <= not(inputs(120));
    layer0_outputs(6203) <= '0';
    layer0_outputs(6204) <= '0';
    layer0_outputs(6205) <= inputs(231);
    layer0_outputs(6206) <= not(inputs(104));
    layer0_outputs(6207) <= (inputs(217)) and (inputs(237));
    layer0_outputs(6208) <= (inputs(203)) and not (inputs(123));
    layer0_outputs(6209) <= not((inputs(209)) xor (inputs(158)));
    layer0_outputs(6210) <= not((inputs(156)) or (inputs(55)));
    layer0_outputs(6211) <= (inputs(111)) xor (inputs(221));
    layer0_outputs(6212) <= inputs(139);
    layer0_outputs(6213) <= '1';
    layer0_outputs(6214) <= not(inputs(16));
    layer0_outputs(6215) <= not(inputs(176)) or (inputs(158));
    layer0_outputs(6216) <= (inputs(111)) and (inputs(181));
    layer0_outputs(6217) <= not(inputs(203)) or (inputs(212));
    layer0_outputs(6218) <= not((inputs(78)) xor (inputs(175)));
    layer0_outputs(6219) <= inputs(188);
    layer0_outputs(6220) <= not((inputs(77)) or (inputs(9)));
    layer0_outputs(6221) <= inputs(132);
    layer0_outputs(6222) <= inputs(86);
    layer0_outputs(6223) <= inputs(78);
    layer0_outputs(6224) <= inputs(231);
    layer0_outputs(6225) <= not(inputs(80));
    layer0_outputs(6226) <= not((inputs(213)) or (inputs(35)));
    layer0_outputs(6227) <= (inputs(48)) and not (inputs(166));
    layer0_outputs(6228) <= (inputs(135)) and not (inputs(38));
    layer0_outputs(6229) <= inputs(43);
    layer0_outputs(6230) <= not(inputs(86)) or (inputs(253));
    layer0_outputs(6231) <= not(inputs(76));
    layer0_outputs(6232) <= (inputs(183)) and (inputs(92));
    layer0_outputs(6233) <= (inputs(159)) and not (inputs(129));
    layer0_outputs(6234) <= (inputs(58)) and (inputs(137));
    layer0_outputs(6235) <= not(inputs(229)) or (inputs(27));
    layer0_outputs(6236) <= not(inputs(194));
    layer0_outputs(6237) <= '0';
    layer0_outputs(6238) <= not(inputs(213)) or (inputs(237));
    layer0_outputs(6239) <= not(inputs(15)) or (inputs(137));
    layer0_outputs(6240) <= '0';
    layer0_outputs(6241) <= '1';
    layer0_outputs(6242) <= inputs(0);
    layer0_outputs(6243) <= '1';
    layer0_outputs(6244) <= inputs(0);
    layer0_outputs(6245) <= (inputs(4)) xor (inputs(16));
    layer0_outputs(6246) <= not(inputs(222)) or (inputs(234));
    layer0_outputs(6247) <= not((inputs(45)) or (inputs(107)));
    layer0_outputs(6248) <= inputs(205);
    layer0_outputs(6249) <= '1';
    layer0_outputs(6250) <= not(inputs(52));
    layer0_outputs(6251) <= '1';
    layer0_outputs(6252) <= '0';
    layer0_outputs(6253) <= not(inputs(118));
    layer0_outputs(6254) <= (inputs(21)) or (inputs(41));
    layer0_outputs(6255) <= (inputs(151)) and not (inputs(128));
    layer0_outputs(6256) <= '0';
    layer0_outputs(6257) <= '0';
    layer0_outputs(6258) <= not(inputs(81));
    layer0_outputs(6259) <= not(inputs(98)) or (inputs(198));
    layer0_outputs(6260) <= (inputs(1)) xor (inputs(90));
    layer0_outputs(6261) <= '1';
    layer0_outputs(6262) <= not((inputs(107)) or (inputs(35)));
    layer0_outputs(6263) <= (inputs(49)) and not (inputs(136));
    layer0_outputs(6264) <= inputs(23);
    layer0_outputs(6265) <= inputs(112);
    layer0_outputs(6266) <= inputs(144);
    layer0_outputs(6267) <= '0';
    layer0_outputs(6268) <= (inputs(43)) and (inputs(29));
    layer0_outputs(6269) <= not((inputs(244)) or (inputs(56)));
    layer0_outputs(6270) <= (inputs(23)) and not (inputs(178));
    layer0_outputs(6271) <= not(inputs(118));
    layer0_outputs(6272) <= inputs(195);
    layer0_outputs(6273) <= not(inputs(38));
    layer0_outputs(6274) <= '0';
    layer0_outputs(6275) <= inputs(167);
    layer0_outputs(6276) <= not(inputs(16));
    layer0_outputs(6277) <= (inputs(48)) and not (inputs(249));
    layer0_outputs(6278) <= (inputs(188)) and not (inputs(241));
    layer0_outputs(6279) <= not((inputs(18)) and (inputs(30)));
    layer0_outputs(6280) <= (inputs(95)) or (inputs(159));
    layer0_outputs(6281) <= not(inputs(235));
    layer0_outputs(6282) <= not(inputs(129));
    layer0_outputs(6283) <= not((inputs(50)) and (inputs(73)));
    layer0_outputs(6284) <= '0';
    layer0_outputs(6285) <= not(inputs(84));
    layer0_outputs(6286) <= '1';
    layer0_outputs(6287) <= '1';
    layer0_outputs(6288) <= (inputs(175)) and (inputs(57));
    layer0_outputs(6289) <= not((inputs(182)) and (inputs(202)));
    layer0_outputs(6290) <= (inputs(27)) or (inputs(4));
    layer0_outputs(6291) <= (inputs(194)) or (inputs(178));
    layer0_outputs(6292) <= not(inputs(189)) or (inputs(25));
    layer0_outputs(6293) <= inputs(37);
    layer0_outputs(6294) <= (inputs(131)) or (inputs(3));
    layer0_outputs(6295) <= '1';
    layer0_outputs(6296) <= '1';
    layer0_outputs(6297) <= (inputs(179)) and not (inputs(62));
    layer0_outputs(6298) <= (inputs(96)) and not (inputs(206));
    layer0_outputs(6299) <= inputs(99);
    layer0_outputs(6300) <= not(inputs(179));
    layer0_outputs(6301) <= '0';
    layer0_outputs(6302) <= inputs(163);
    layer0_outputs(6303) <= not(inputs(120)) or (inputs(65));
    layer0_outputs(6304) <= '0';
    layer0_outputs(6305) <= not(inputs(126)) or (inputs(27));
    layer0_outputs(6306) <= '0';
    layer0_outputs(6307) <= not(inputs(148)) or (inputs(30));
    layer0_outputs(6308) <= not(inputs(133));
    layer0_outputs(6309) <= (inputs(136)) and not (inputs(36));
    layer0_outputs(6310) <= (inputs(194)) and not (inputs(196));
    layer0_outputs(6311) <= (inputs(164)) and not (inputs(191));
    layer0_outputs(6312) <= inputs(255);
    layer0_outputs(6313) <= (inputs(78)) or (inputs(124));
    layer0_outputs(6314) <= (inputs(176)) and not (inputs(95));
    layer0_outputs(6315) <= '1';
    layer0_outputs(6316) <= (inputs(70)) and (inputs(195));
    layer0_outputs(6317) <= (inputs(9)) or (inputs(44));
    layer0_outputs(6318) <= inputs(172);
    layer0_outputs(6319) <= (inputs(174)) or (inputs(201));
    layer0_outputs(6320) <= (inputs(217)) or (inputs(77));
    layer0_outputs(6321) <= (inputs(3)) or (inputs(36));
    layer0_outputs(6322) <= not((inputs(209)) or (inputs(17)));
    layer0_outputs(6323) <= (inputs(108)) or (inputs(250));
    layer0_outputs(6324) <= (inputs(210)) and not (inputs(96));
    layer0_outputs(6325) <= (inputs(48)) xor (inputs(143));
    layer0_outputs(6326) <= (inputs(177)) or (inputs(223));
    layer0_outputs(6327) <= (inputs(173)) and not (inputs(67));
    layer0_outputs(6328) <= not(inputs(156)) or (inputs(235));
    layer0_outputs(6329) <= not((inputs(202)) or (inputs(243)));
    layer0_outputs(6330) <= not(inputs(141)) or (inputs(204));
    layer0_outputs(6331) <= inputs(202);
    layer0_outputs(6332) <= (inputs(106)) or (inputs(3));
    layer0_outputs(6333) <= '0';
    layer0_outputs(6334) <= (inputs(118)) and (inputs(227));
    layer0_outputs(6335) <= (inputs(72)) or (inputs(178));
    layer0_outputs(6336) <= not((inputs(24)) and (inputs(56)));
    layer0_outputs(6337) <= not((inputs(174)) xor (inputs(160)));
    layer0_outputs(6338) <= inputs(204);
    layer0_outputs(6339) <= not(inputs(30));
    layer0_outputs(6340) <= '0';
    layer0_outputs(6341) <= (inputs(80)) or (inputs(198));
    layer0_outputs(6342) <= not((inputs(251)) xor (inputs(33)));
    layer0_outputs(6343) <= inputs(175);
    layer0_outputs(6344) <= not(inputs(149));
    layer0_outputs(6345) <= not((inputs(71)) or (inputs(86)));
    layer0_outputs(6346) <= '1';
    layer0_outputs(6347) <= '0';
    layer0_outputs(6348) <= (inputs(146)) or (inputs(155));
    layer0_outputs(6349) <= not(inputs(226)) or (inputs(127));
    layer0_outputs(6350) <= (inputs(111)) and not (inputs(7));
    layer0_outputs(6351) <= (inputs(199)) and not (inputs(57));
    layer0_outputs(6352) <= '0';
    layer0_outputs(6353) <= (inputs(255)) xor (inputs(51));
    layer0_outputs(6354) <= '1';
    layer0_outputs(6355) <= not((inputs(112)) and (inputs(160)));
    layer0_outputs(6356) <= (inputs(179)) xor (inputs(207));
    layer0_outputs(6357) <= inputs(164);
    layer0_outputs(6358) <= inputs(246);
    layer0_outputs(6359) <= not((inputs(238)) xor (inputs(51)));
    layer0_outputs(6360) <= inputs(147);
    layer0_outputs(6361) <= not(inputs(226));
    layer0_outputs(6362) <= '0';
    layer0_outputs(6363) <= not(inputs(35)) or (inputs(251));
    layer0_outputs(6364) <= inputs(154);
    layer0_outputs(6365) <= not(inputs(103));
    layer0_outputs(6366) <= (inputs(28)) and not (inputs(243));
    layer0_outputs(6367) <= not((inputs(202)) or (inputs(7)));
    layer0_outputs(6368) <= inputs(180);
    layer0_outputs(6369) <= inputs(53);
    layer0_outputs(6370) <= '1';
    layer0_outputs(6371) <= inputs(46);
    layer0_outputs(6372) <= not(inputs(66));
    layer0_outputs(6373) <= '1';
    layer0_outputs(6374) <= not(inputs(135));
    layer0_outputs(6375) <= '0';
    layer0_outputs(6376) <= not((inputs(50)) xor (inputs(70)));
    layer0_outputs(6377) <= inputs(119);
    layer0_outputs(6378) <= (inputs(67)) and not (inputs(197));
    layer0_outputs(6379) <= not((inputs(54)) xor (inputs(239)));
    layer0_outputs(6380) <= inputs(247);
    layer0_outputs(6381) <= (inputs(31)) and not (inputs(111));
    layer0_outputs(6382) <= inputs(114);
    layer0_outputs(6383) <= not((inputs(228)) or (inputs(154)));
    layer0_outputs(6384) <= (inputs(217)) and not (inputs(107));
    layer0_outputs(6385) <= not(inputs(183)) or (inputs(185));
    layer0_outputs(6386) <= (inputs(192)) and not (inputs(57));
    layer0_outputs(6387) <= (inputs(48)) and not (inputs(78));
    layer0_outputs(6388) <= '0';
    layer0_outputs(6389) <= (inputs(162)) and not (inputs(31));
    layer0_outputs(6390) <= not((inputs(44)) and (inputs(72)));
    layer0_outputs(6391) <= not((inputs(43)) or (inputs(59)));
    layer0_outputs(6392) <= not((inputs(195)) or (inputs(142)));
    layer0_outputs(6393) <= (inputs(37)) and not (inputs(70));
    layer0_outputs(6394) <= not((inputs(208)) and (inputs(16)));
    layer0_outputs(6395) <= not((inputs(101)) or (inputs(167)));
    layer0_outputs(6396) <= not(inputs(161));
    layer0_outputs(6397) <= (inputs(183)) and (inputs(191));
    layer0_outputs(6398) <= (inputs(47)) and not (inputs(143));
    layer0_outputs(6399) <= not(inputs(165));
    layer0_outputs(6400) <= (inputs(131)) and (inputs(68));
    layer0_outputs(6401) <= not(inputs(66));
    layer0_outputs(6402) <= not((inputs(46)) and (inputs(67)));
    layer0_outputs(6403) <= not(inputs(89)) or (inputs(65));
    layer0_outputs(6404) <= not(inputs(182));
    layer0_outputs(6405) <= (inputs(183)) and (inputs(204));
    layer0_outputs(6406) <= (inputs(236)) and (inputs(137));
    layer0_outputs(6407) <= not((inputs(122)) or (inputs(208)));
    layer0_outputs(6408) <= inputs(7);
    layer0_outputs(6409) <= (inputs(232)) and not (inputs(14));
    layer0_outputs(6410) <= not(inputs(212));
    layer0_outputs(6411) <= not(inputs(86));
    layer0_outputs(6412) <= not((inputs(181)) or (inputs(248)));
    layer0_outputs(6413) <= (inputs(139)) and not (inputs(43));
    layer0_outputs(6414) <= inputs(45);
    layer0_outputs(6415) <= '0';
    layer0_outputs(6416) <= not(inputs(122));
    layer0_outputs(6417) <= (inputs(212)) or (inputs(94));
    layer0_outputs(6418) <= (inputs(10)) xor (inputs(175));
    layer0_outputs(6419) <= (inputs(232)) or (inputs(177));
    layer0_outputs(6420) <= (inputs(213)) and not (inputs(20));
    layer0_outputs(6421) <= not(inputs(14));
    layer0_outputs(6422) <= (inputs(215)) and not (inputs(162));
    layer0_outputs(6423) <= '1';
    layer0_outputs(6424) <= (inputs(189)) and (inputs(181));
    layer0_outputs(6425) <= '0';
    layer0_outputs(6426) <= not(inputs(189)) or (inputs(211));
    layer0_outputs(6427) <= not((inputs(144)) and (inputs(163)));
    layer0_outputs(6428) <= not((inputs(244)) or (inputs(30)));
    layer0_outputs(6429) <= '1';
    layer0_outputs(6430) <= not(inputs(189)) or (inputs(110));
    layer0_outputs(6431) <= inputs(230);
    layer0_outputs(6432) <= inputs(230);
    layer0_outputs(6433) <= not(inputs(198));
    layer0_outputs(6434) <= '1';
    layer0_outputs(6435) <= not((inputs(102)) or (inputs(84)));
    layer0_outputs(6436) <= inputs(103);
    layer0_outputs(6437) <= not((inputs(19)) or (inputs(227)));
    layer0_outputs(6438) <= '0';
    layer0_outputs(6439) <= not(inputs(22)) or (inputs(144));
    layer0_outputs(6440) <= not(inputs(109));
    layer0_outputs(6441) <= inputs(148);
    layer0_outputs(6442) <= inputs(63);
    layer0_outputs(6443) <= (inputs(61)) or (inputs(249));
    layer0_outputs(6444) <= '0';
    layer0_outputs(6445) <= not(inputs(82));
    layer0_outputs(6446) <= (inputs(95)) or (inputs(59));
    layer0_outputs(6447) <= not((inputs(92)) and (inputs(24)));
    layer0_outputs(6448) <= not(inputs(230)) or (inputs(25));
    layer0_outputs(6449) <= not((inputs(200)) or (inputs(210)));
    layer0_outputs(6450) <= inputs(114);
    layer0_outputs(6451) <= not((inputs(234)) or (inputs(122)));
    layer0_outputs(6452) <= inputs(150);
    layer0_outputs(6453) <= '1';
    layer0_outputs(6454) <= not((inputs(170)) and (inputs(250)));
    layer0_outputs(6455) <= not(inputs(121)) or (inputs(166));
    layer0_outputs(6456) <= not((inputs(30)) or (inputs(153)));
    layer0_outputs(6457) <= not(inputs(208)) or (inputs(212));
    layer0_outputs(6458) <= inputs(45);
    layer0_outputs(6459) <= not(inputs(22)) or (inputs(173));
    layer0_outputs(6460) <= not((inputs(24)) or (inputs(51)));
    layer0_outputs(6461) <= (inputs(219)) and not (inputs(32));
    layer0_outputs(6462) <= not(inputs(83)) or (inputs(144));
    layer0_outputs(6463) <= inputs(42);
    layer0_outputs(6464) <= '1';
    layer0_outputs(6465) <= not(inputs(226)) or (inputs(244));
    layer0_outputs(6466) <= '1';
    layer0_outputs(6467) <= not((inputs(98)) and (inputs(137)));
    layer0_outputs(6468) <= not((inputs(218)) or (inputs(173)));
    layer0_outputs(6469) <= not(inputs(36)) or (inputs(78));
    layer0_outputs(6470) <= not((inputs(230)) or (inputs(245)));
    layer0_outputs(6471) <= inputs(5);
    layer0_outputs(6472) <= not(inputs(153)) or (inputs(153));
    layer0_outputs(6473) <= not((inputs(197)) xor (inputs(239)));
    layer0_outputs(6474) <= (inputs(199)) or (inputs(232));
    layer0_outputs(6475) <= not((inputs(254)) or (inputs(111)));
    layer0_outputs(6476) <= not(inputs(42)) or (inputs(141));
    layer0_outputs(6477) <= (inputs(53)) and not (inputs(192));
    layer0_outputs(6478) <= (inputs(26)) and not (inputs(144));
    layer0_outputs(6479) <= '1';
    layer0_outputs(6480) <= (inputs(53)) xor (inputs(158));
    layer0_outputs(6481) <= '0';
    layer0_outputs(6482) <= (inputs(171)) xor (inputs(158));
    layer0_outputs(6483) <= inputs(230);
    layer0_outputs(6484) <= (inputs(172)) and not (inputs(13));
    layer0_outputs(6485) <= (inputs(255)) or (inputs(238));
    layer0_outputs(6486) <= not(inputs(207)) or (inputs(64));
    layer0_outputs(6487) <= '1';
    layer0_outputs(6488) <= inputs(58);
    layer0_outputs(6489) <= not(inputs(174)) or (inputs(127));
    layer0_outputs(6490) <= not((inputs(78)) or (inputs(66)));
    layer0_outputs(6491) <= '0';
    layer0_outputs(6492) <= not(inputs(80)) or (inputs(79));
    layer0_outputs(6493) <= (inputs(60)) and (inputs(17));
    layer0_outputs(6494) <= (inputs(140)) and not (inputs(57));
    layer0_outputs(6495) <= inputs(209);
    layer0_outputs(6496) <= not(inputs(114)) or (inputs(94));
    layer0_outputs(6497) <= not((inputs(201)) and (inputs(118)));
    layer0_outputs(6498) <= inputs(234);
    layer0_outputs(6499) <= not(inputs(78));
    layer0_outputs(6500) <= inputs(57);
    layer0_outputs(6501) <= '0';
    layer0_outputs(6502) <= not((inputs(238)) xor (inputs(181)));
    layer0_outputs(6503) <= inputs(120);
    layer0_outputs(6504) <= not(inputs(146)) or (inputs(107));
    layer0_outputs(6505) <= (inputs(54)) xor (inputs(104));
    layer0_outputs(6506) <= not(inputs(108)) or (inputs(55));
    layer0_outputs(6507) <= (inputs(22)) and (inputs(201));
    layer0_outputs(6508) <= inputs(239);
    layer0_outputs(6509) <= not((inputs(150)) or (inputs(225)));
    layer0_outputs(6510) <= not(inputs(98));
    layer0_outputs(6511) <= '0';
    layer0_outputs(6512) <= not((inputs(51)) or (inputs(218)));
    layer0_outputs(6513) <= not(inputs(156));
    layer0_outputs(6514) <= not((inputs(204)) and (inputs(139)));
    layer0_outputs(6515) <= not(inputs(251)) or (inputs(125));
    layer0_outputs(6516) <= not(inputs(184));
    layer0_outputs(6517) <= not(inputs(237));
    layer0_outputs(6518) <= '1';
    layer0_outputs(6519) <= (inputs(1)) and not (inputs(157));
    layer0_outputs(6520) <= '1';
    layer0_outputs(6521) <= not(inputs(133)) or (inputs(249));
    layer0_outputs(6522) <= not((inputs(218)) or (inputs(178)));
    layer0_outputs(6523) <= inputs(24);
    layer0_outputs(6524) <= '1';
    layer0_outputs(6525) <= '0';
    layer0_outputs(6526) <= not(inputs(218)) or (inputs(195));
    layer0_outputs(6527) <= (inputs(9)) and not (inputs(9));
    layer0_outputs(6528) <= not(inputs(15));
    layer0_outputs(6529) <= '0';
    layer0_outputs(6530) <= inputs(209);
    layer0_outputs(6531) <= (inputs(185)) and not (inputs(209));
    layer0_outputs(6532) <= '0';
    layer0_outputs(6533) <= (inputs(51)) and not (inputs(253));
    layer0_outputs(6534) <= inputs(200);
    layer0_outputs(6535) <= not(inputs(177));
    layer0_outputs(6536) <= not((inputs(166)) or (inputs(177)));
    layer0_outputs(6537) <= not((inputs(135)) or (inputs(168)));
    layer0_outputs(6538) <= not(inputs(243));
    layer0_outputs(6539) <= '1';
    layer0_outputs(6540) <= inputs(109);
    layer0_outputs(6541) <= '0';
    layer0_outputs(6542) <= not(inputs(97));
    layer0_outputs(6543) <= (inputs(2)) and not (inputs(251));
    layer0_outputs(6544) <= '1';
    layer0_outputs(6545) <= (inputs(249)) and not (inputs(137));
    layer0_outputs(6546) <= '1';
    layer0_outputs(6547) <= not(inputs(71)) or (inputs(17));
    layer0_outputs(6548) <= not(inputs(99)) or (inputs(241));
    layer0_outputs(6549) <= not(inputs(36));
    layer0_outputs(6550) <= not(inputs(71)) or (inputs(45));
    layer0_outputs(6551) <= (inputs(106)) and not (inputs(195));
    layer0_outputs(6552) <= (inputs(252)) and not (inputs(43));
    layer0_outputs(6553) <= (inputs(167)) and not (inputs(129));
    layer0_outputs(6554) <= (inputs(158)) and not (inputs(31));
    layer0_outputs(6555) <= not(inputs(150));
    layer0_outputs(6556) <= '1';
    layer0_outputs(6557) <= not(inputs(66));
    layer0_outputs(6558) <= not((inputs(97)) or (inputs(66)));
    layer0_outputs(6559) <= not(inputs(68)) or (inputs(43));
    layer0_outputs(6560) <= not((inputs(210)) or (inputs(46)));
    layer0_outputs(6561) <= (inputs(188)) and not (inputs(193));
    layer0_outputs(6562) <= '1';
    layer0_outputs(6563) <= '1';
    layer0_outputs(6564) <= not(inputs(207));
    layer0_outputs(6565) <= inputs(25);
    layer0_outputs(6566) <= not(inputs(228));
    layer0_outputs(6567) <= '0';
    layer0_outputs(6568) <= inputs(145);
    layer0_outputs(6569) <= not(inputs(45)) or (inputs(82));
    layer0_outputs(6570) <= (inputs(27)) or (inputs(242));
    layer0_outputs(6571) <= not((inputs(215)) or (inputs(230)));
    layer0_outputs(6572) <= not((inputs(110)) or (inputs(203)));
    layer0_outputs(6573) <= not((inputs(208)) and (inputs(149)));
    layer0_outputs(6574) <= not(inputs(206));
    layer0_outputs(6575) <= (inputs(244)) or (inputs(129));
    layer0_outputs(6576) <= not(inputs(227));
    layer0_outputs(6577) <= (inputs(169)) or (inputs(206));
    layer0_outputs(6578) <= not((inputs(49)) or (inputs(105)));
    layer0_outputs(6579) <= not((inputs(85)) xor (inputs(218)));
    layer0_outputs(6580) <= not(inputs(116)) or (inputs(50));
    layer0_outputs(6581) <= (inputs(140)) or (inputs(113));
    layer0_outputs(6582) <= (inputs(139)) and (inputs(208));
    layer0_outputs(6583) <= (inputs(147)) or (inputs(74));
    layer0_outputs(6584) <= '0';
    layer0_outputs(6585) <= (inputs(206)) and not (inputs(162));
    layer0_outputs(6586) <= '0';
    layer0_outputs(6587) <= inputs(130);
    layer0_outputs(6588) <= not((inputs(251)) and (inputs(244)));
    layer0_outputs(6589) <= '0';
    layer0_outputs(6590) <= inputs(79);
    layer0_outputs(6591) <= (inputs(243)) and not (inputs(186));
    layer0_outputs(6592) <= inputs(190);
    layer0_outputs(6593) <= '0';
    layer0_outputs(6594) <= '1';
    layer0_outputs(6595) <= '1';
    layer0_outputs(6596) <= inputs(251);
    layer0_outputs(6597) <= inputs(77);
    layer0_outputs(6598) <= not((inputs(9)) and (inputs(2)));
    layer0_outputs(6599) <= (inputs(125)) and (inputs(178));
    layer0_outputs(6600) <= (inputs(166)) and not (inputs(200));
    layer0_outputs(6601) <= not(inputs(135)) or (inputs(65));
    layer0_outputs(6602) <= '0';
    layer0_outputs(6603) <= '0';
    layer0_outputs(6604) <= not(inputs(51)) or (inputs(184));
    layer0_outputs(6605) <= not(inputs(67));
    layer0_outputs(6606) <= not(inputs(21));
    layer0_outputs(6607) <= (inputs(184)) and (inputs(188));
    layer0_outputs(6608) <= inputs(191);
    layer0_outputs(6609) <= inputs(176);
    layer0_outputs(6610) <= not((inputs(47)) or (inputs(219)));
    layer0_outputs(6611) <= inputs(159);
    layer0_outputs(6612) <= not((inputs(84)) or (inputs(6)));
    layer0_outputs(6613) <= not((inputs(10)) and (inputs(128)));
    layer0_outputs(6614) <= not(inputs(71)) or (inputs(36));
    layer0_outputs(6615) <= '0';
    layer0_outputs(6616) <= (inputs(31)) or (inputs(44));
    layer0_outputs(6617) <= not((inputs(240)) and (inputs(170)));
    layer0_outputs(6618) <= inputs(185);
    layer0_outputs(6619) <= not((inputs(168)) and (inputs(250)));
    layer0_outputs(6620) <= inputs(95);
    layer0_outputs(6621) <= (inputs(107)) and not (inputs(10));
    layer0_outputs(6622) <= '0';
    layer0_outputs(6623) <= not(inputs(224)) or (inputs(47));
    layer0_outputs(6624) <= (inputs(181)) or (inputs(193));
    layer0_outputs(6625) <= inputs(7);
    layer0_outputs(6626) <= not(inputs(194));
    layer0_outputs(6627) <= inputs(109);
    layer0_outputs(6628) <= not(inputs(22)) or (inputs(146));
    layer0_outputs(6629) <= not(inputs(219)) or (inputs(85));
    layer0_outputs(6630) <= not(inputs(137));
    layer0_outputs(6631) <= '1';
    layer0_outputs(6632) <= not((inputs(21)) or (inputs(32)));
    layer0_outputs(6633) <= not((inputs(101)) or (inputs(124)));
    layer0_outputs(6634) <= inputs(109);
    layer0_outputs(6635) <= (inputs(225)) and not (inputs(43));
    layer0_outputs(6636) <= (inputs(230)) and (inputs(165));
    layer0_outputs(6637) <= (inputs(115)) and not (inputs(106));
    layer0_outputs(6638) <= '1';
    layer0_outputs(6639) <= '0';
    layer0_outputs(6640) <= (inputs(247)) and not (inputs(248));
    layer0_outputs(6641) <= not(inputs(205)) or (inputs(185));
    layer0_outputs(6642) <= not(inputs(142)) or (inputs(44));
    layer0_outputs(6643) <= not((inputs(205)) xor (inputs(32)));
    layer0_outputs(6644) <= not(inputs(182));
    layer0_outputs(6645) <= not(inputs(60));
    layer0_outputs(6646) <= (inputs(158)) and not (inputs(80));
    layer0_outputs(6647) <= (inputs(213)) or (inputs(72));
    layer0_outputs(6648) <= not(inputs(19));
    layer0_outputs(6649) <= not(inputs(100)) or (inputs(101));
    layer0_outputs(6650) <= (inputs(165)) and not (inputs(207));
    layer0_outputs(6651) <= (inputs(216)) and not (inputs(2));
    layer0_outputs(6652) <= not(inputs(4)) or (inputs(44));
    layer0_outputs(6653) <= (inputs(184)) and (inputs(45));
    layer0_outputs(6654) <= (inputs(244)) or (inputs(247));
    layer0_outputs(6655) <= '0';
    layer0_outputs(6656) <= not((inputs(138)) and (inputs(108)));
    layer0_outputs(6657) <= '1';
    layer0_outputs(6658) <= inputs(137);
    layer0_outputs(6659) <= '1';
    layer0_outputs(6660) <= not(inputs(24)) or (inputs(145));
    layer0_outputs(6661) <= not((inputs(119)) and (inputs(26)));
    layer0_outputs(6662) <= (inputs(79)) and (inputs(4));
    layer0_outputs(6663) <= (inputs(171)) or (inputs(174));
    layer0_outputs(6664) <= not(inputs(62));
    layer0_outputs(6665) <= not(inputs(89));
    layer0_outputs(6666) <= not(inputs(104)) or (inputs(174));
    layer0_outputs(6667) <= '0';
    layer0_outputs(6668) <= (inputs(20)) xor (inputs(187));
    layer0_outputs(6669) <= '0';
    layer0_outputs(6670) <= not((inputs(116)) or (inputs(63)));
    layer0_outputs(6671) <= (inputs(93)) xor (inputs(224));
    layer0_outputs(6672) <= '1';
    layer0_outputs(6673) <= (inputs(131)) xor (inputs(206));
    layer0_outputs(6674) <= '0';
    layer0_outputs(6675) <= '0';
    layer0_outputs(6676) <= (inputs(36)) and not (inputs(66));
    layer0_outputs(6677) <= not((inputs(19)) or (inputs(93)));
    layer0_outputs(6678) <= inputs(83);
    layer0_outputs(6679) <= (inputs(220)) and not (inputs(77));
    layer0_outputs(6680) <= not((inputs(58)) and (inputs(111)));
    layer0_outputs(6681) <= inputs(108);
    layer0_outputs(6682) <= '0';
    layer0_outputs(6683) <= '1';
    layer0_outputs(6684) <= '0';
    layer0_outputs(6685) <= '0';
    layer0_outputs(6686) <= not(inputs(235));
    layer0_outputs(6687) <= inputs(81);
    layer0_outputs(6688) <= (inputs(198)) or (inputs(93));
    layer0_outputs(6689) <= '1';
    layer0_outputs(6690) <= not((inputs(253)) or (inputs(123)));
    layer0_outputs(6691) <= (inputs(155)) and (inputs(149));
    layer0_outputs(6692) <= not((inputs(142)) or (inputs(139)));
    layer0_outputs(6693) <= not(inputs(48)) or (inputs(20));
    layer0_outputs(6694) <= (inputs(232)) or (inputs(25));
    layer0_outputs(6695) <= inputs(5);
    layer0_outputs(6696) <= (inputs(2)) and not (inputs(154));
    layer0_outputs(6697) <= (inputs(103)) and not (inputs(202));
    layer0_outputs(6698) <= not(inputs(130));
    layer0_outputs(6699) <= '1';
    layer0_outputs(6700) <= not(inputs(98));
    layer0_outputs(6701) <= inputs(39);
    layer0_outputs(6702) <= inputs(107);
    layer0_outputs(6703) <= inputs(114);
    layer0_outputs(6704) <= inputs(48);
    layer0_outputs(6705) <= not(inputs(42));
    layer0_outputs(6706) <= '1';
    layer0_outputs(6707) <= not(inputs(32));
    layer0_outputs(6708) <= inputs(9);
    layer0_outputs(6709) <= not(inputs(107));
    layer0_outputs(6710) <= not(inputs(161)) or (inputs(67));
    layer0_outputs(6711) <= not(inputs(235)) or (inputs(118));
    layer0_outputs(6712) <= (inputs(135)) and (inputs(101));
    layer0_outputs(6713) <= (inputs(251)) and not (inputs(242));
    layer0_outputs(6714) <= not((inputs(97)) and (inputs(143)));
    layer0_outputs(6715) <= not(inputs(170));
    layer0_outputs(6716) <= inputs(217);
    layer0_outputs(6717) <= '0';
    layer0_outputs(6718) <= not(inputs(78)) or (inputs(175));
    layer0_outputs(6719) <= not(inputs(161));
    layer0_outputs(6720) <= inputs(75);
    layer0_outputs(6721) <= not(inputs(206));
    layer0_outputs(6722) <= (inputs(195)) and not (inputs(84));
    layer0_outputs(6723) <= '1';
    layer0_outputs(6724) <= not((inputs(147)) or (inputs(7)));
    layer0_outputs(6725) <= not(inputs(16)) or (inputs(240));
    layer0_outputs(6726) <= (inputs(190)) and not (inputs(109));
    layer0_outputs(6727) <= not((inputs(76)) or (inputs(131)));
    layer0_outputs(6728) <= not(inputs(35));
    layer0_outputs(6729) <= not(inputs(161));
    layer0_outputs(6730) <= not(inputs(241));
    layer0_outputs(6731) <= inputs(88);
    layer0_outputs(6732) <= (inputs(84)) and (inputs(27));
    layer0_outputs(6733) <= '1';
    layer0_outputs(6734) <= not(inputs(81));
    layer0_outputs(6735) <= (inputs(97)) and not (inputs(137));
    layer0_outputs(6736) <= '0';
    layer0_outputs(6737) <= (inputs(110)) and not (inputs(73));
    layer0_outputs(6738) <= '1';
    layer0_outputs(6739) <= not(inputs(207));
    layer0_outputs(6740) <= (inputs(153)) and not (inputs(32));
    layer0_outputs(6741) <= '0';
    layer0_outputs(6742) <= (inputs(30)) and (inputs(157));
    layer0_outputs(6743) <= not(inputs(18)) or (inputs(120));
    layer0_outputs(6744) <= not(inputs(131)) or (inputs(49));
    layer0_outputs(6745) <= inputs(24);
    layer0_outputs(6746) <= not(inputs(15)) or (inputs(211));
    layer0_outputs(6747) <= not(inputs(158)) or (inputs(249));
    layer0_outputs(6748) <= inputs(125);
    layer0_outputs(6749) <= (inputs(253)) and (inputs(211));
    layer0_outputs(6750) <= not(inputs(191));
    layer0_outputs(6751) <= inputs(42);
    layer0_outputs(6752) <= not(inputs(55));
    layer0_outputs(6753) <= (inputs(46)) or (inputs(61));
    layer0_outputs(6754) <= (inputs(106)) and (inputs(181));
    layer0_outputs(6755) <= not(inputs(67)) or (inputs(168));
    layer0_outputs(6756) <= not(inputs(137)) or (inputs(206));
    layer0_outputs(6757) <= not(inputs(189));
    layer0_outputs(6758) <= not(inputs(15));
    layer0_outputs(6759) <= (inputs(68)) and not (inputs(29));
    layer0_outputs(6760) <= not((inputs(216)) and (inputs(142)));
    layer0_outputs(6761) <= (inputs(108)) or (inputs(242));
    layer0_outputs(6762) <= not((inputs(194)) or (inputs(143)));
    layer0_outputs(6763) <= inputs(89);
    layer0_outputs(6764) <= not((inputs(115)) or (inputs(237)));
    layer0_outputs(6765) <= inputs(96);
    layer0_outputs(6766) <= not(inputs(133));
    layer0_outputs(6767) <= not((inputs(197)) or (inputs(202)));
    layer0_outputs(6768) <= not(inputs(20));
    layer0_outputs(6769) <= not(inputs(211)) or (inputs(32));
    layer0_outputs(6770) <= not(inputs(176)) or (inputs(230));
    layer0_outputs(6771) <= '1';
    layer0_outputs(6772) <= not(inputs(29));
    layer0_outputs(6773) <= '1';
    layer0_outputs(6774) <= not(inputs(23));
    layer0_outputs(6775) <= (inputs(6)) and not (inputs(129));
    layer0_outputs(6776) <= (inputs(16)) xor (inputs(64));
    layer0_outputs(6777) <= inputs(27);
    layer0_outputs(6778) <= not((inputs(8)) or (inputs(177)));
    layer0_outputs(6779) <= (inputs(173)) or (inputs(180));
    layer0_outputs(6780) <= not((inputs(90)) or (inputs(74)));
    layer0_outputs(6781) <= not(inputs(218)) or (inputs(238));
    layer0_outputs(6782) <= inputs(205);
    layer0_outputs(6783) <= (inputs(86)) xor (inputs(106));
    layer0_outputs(6784) <= '1';
    layer0_outputs(6785) <= not((inputs(4)) or (inputs(132)));
    layer0_outputs(6786) <= (inputs(139)) and not (inputs(194));
    layer0_outputs(6787) <= (inputs(117)) and not (inputs(206));
    layer0_outputs(6788) <= '0';
    layer0_outputs(6789) <= (inputs(240)) xor (inputs(168));
    layer0_outputs(6790) <= not(inputs(0));
    layer0_outputs(6791) <= inputs(26);
    layer0_outputs(6792) <= '0';
    layer0_outputs(6793) <= not(inputs(192));
    layer0_outputs(6794) <= '0';
    layer0_outputs(6795) <= not((inputs(40)) xor (inputs(33)));
    layer0_outputs(6796) <= inputs(2);
    layer0_outputs(6797) <= (inputs(181)) and (inputs(216));
    layer0_outputs(6798) <= not((inputs(119)) or (inputs(25)));
    layer0_outputs(6799) <= inputs(20);
    layer0_outputs(6800) <= inputs(110);
    layer0_outputs(6801) <= not((inputs(208)) or (inputs(198)));
    layer0_outputs(6802) <= (inputs(193)) and not (inputs(72));
    layer0_outputs(6803) <= (inputs(78)) or (inputs(227));
    layer0_outputs(6804) <= not(inputs(214));
    layer0_outputs(6805) <= not(inputs(227));
    layer0_outputs(6806) <= not(inputs(28));
    layer0_outputs(6807) <= not(inputs(249));
    layer0_outputs(6808) <= inputs(186);
    layer0_outputs(6809) <= (inputs(4)) xor (inputs(117));
    layer0_outputs(6810) <= '1';
    layer0_outputs(6811) <= not((inputs(225)) or (inputs(211)));
    layer0_outputs(6812) <= not(inputs(70)) or (inputs(207));
    layer0_outputs(6813) <= inputs(167);
    layer0_outputs(6814) <= not(inputs(174));
    layer0_outputs(6815) <= '0';
    layer0_outputs(6816) <= inputs(98);
    layer0_outputs(6817) <= not((inputs(136)) or (inputs(213)));
    layer0_outputs(6818) <= inputs(96);
    layer0_outputs(6819) <= (inputs(203)) and not (inputs(103));
    layer0_outputs(6820) <= not(inputs(110));
    layer0_outputs(6821) <= not(inputs(68));
    layer0_outputs(6822) <= inputs(51);
    layer0_outputs(6823) <= not(inputs(204)) or (inputs(133));
    layer0_outputs(6824) <= inputs(41);
    layer0_outputs(6825) <= (inputs(25)) and not (inputs(193));
    layer0_outputs(6826) <= inputs(165);
    layer0_outputs(6827) <= not(inputs(39)) or (inputs(155));
    layer0_outputs(6828) <= (inputs(244)) and not (inputs(143));
    layer0_outputs(6829) <= not(inputs(127));
    layer0_outputs(6830) <= not(inputs(76)) or (inputs(54));
    layer0_outputs(6831) <= (inputs(203)) and not (inputs(126));
    layer0_outputs(6832) <= inputs(239);
    layer0_outputs(6833) <= not(inputs(238)) or (inputs(14));
    layer0_outputs(6834) <= not(inputs(233));
    layer0_outputs(6835) <= inputs(222);
    layer0_outputs(6836) <= (inputs(28)) or (inputs(106));
    layer0_outputs(6837) <= inputs(38);
    layer0_outputs(6838) <= not(inputs(60));
    layer0_outputs(6839) <= (inputs(82)) or (inputs(97));
    layer0_outputs(6840) <= inputs(122);
    layer0_outputs(6841) <= (inputs(112)) and not (inputs(184));
    layer0_outputs(6842) <= (inputs(133)) or (inputs(173));
    layer0_outputs(6843) <= inputs(111);
    layer0_outputs(6844) <= not(inputs(136)) or (inputs(43));
    layer0_outputs(6845) <= not(inputs(110));
    layer0_outputs(6846) <= not(inputs(249));
    layer0_outputs(6847) <= '0';
    layer0_outputs(6848) <= not(inputs(57));
    layer0_outputs(6849) <= not(inputs(114));
    layer0_outputs(6850) <= '0';
    layer0_outputs(6851) <= not((inputs(105)) and (inputs(68)));
    layer0_outputs(6852) <= inputs(169);
    layer0_outputs(6853) <= '1';
    layer0_outputs(6854) <= inputs(57);
    layer0_outputs(6855) <= (inputs(113)) or (inputs(82));
    layer0_outputs(6856) <= inputs(146);
    layer0_outputs(6857) <= (inputs(156)) and (inputs(64));
    layer0_outputs(6858) <= not(inputs(243)) or (inputs(118));
    layer0_outputs(6859) <= (inputs(204)) and (inputs(93));
    layer0_outputs(6860) <= '1';
    layer0_outputs(6861) <= not((inputs(89)) and (inputs(247)));
    layer0_outputs(6862) <= not((inputs(182)) or (inputs(148)));
    layer0_outputs(6863) <= inputs(131);
    layer0_outputs(6864) <= not((inputs(32)) or (inputs(195)));
    layer0_outputs(6865) <= not(inputs(124));
    layer0_outputs(6866) <= '0';
    layer0_outputs(6867) <= '1';
    layer0_outputs(6868) <= (inputs(48)) or (inputs(156));
    layer0_outputs(6869) <= not((inputs(47)) and (inputs(128)));
    layer0_outputs(6870) <= inputs(121);
    layer0_outputs(6871) <= (inputs(201)) or (inputs(138));
    layer0_outputs(6872) <= '0';
    layer0_outputs(6873) <= (inputs(49)) and not (inputs(14));
    layer0_outputs(6874) <= (inputs(200)) or (inputs(28));
    layer0_outputs(6875) <= '0';
    layer0_outputs(6876) <= inputs(83);
    layer0_outputs(6877) <= '1';
    layer0_outputs(6878) <= not(inputs(85));
    layer0_outputs(6879) <= not(inputs(114)) or (inputs(163));
    layer0_outputs(6880) <= not(inputs(7)) or (inputs(52));
    layer0_outputs(6881) <= inputs(86);
    layer0_outputs(6882) <= '1';
    layer0_outputs(6883) <= (inputs(152)) and not (inputs(80));
    layer0_outputs(6884) <= (inputs(152)) and not (inputs(94));
    layer0_outputs(6885) <= (inputs(9)) and (inputs(118));
    layer0_outputs(6886) <= (inputs(68)) and (inputs(2));
    layer0_outputs(6887) <= (inputs(231)) or (inputs(164));
    layer0_outputs(6888) <= not(inputs(179));
    layer0_outputs(6889) <= inputs(119);
    layer0_outputs(6890) <= (inputs(48)) or (inputs(28));
    layer0_outputs(6891) <= (inputs(82)) xor (inputs(217));
    layer0_outputs(6892) <= '0';
    layer0_outputs(6893) <= (inputs(62)) or (inputs(33));
    layer0_outputs(6894) <= (inputs(72)) and (inputs(248));
    layer0_outputs(6895) <= inputs(181);
    layer0_outputs(6896) <= not(inputs(63));
    layer0_outputs(6897) <= not((inputs(12)) or (inputs(82)));
    layer0_outputs(6898) <= (inputs(226)) and (inputs(177));
    layer0_outputs(6899) <= '0';
    layer0_outputs(6900) <= not((inputs(52)) xor (inputs(21)));
    layer0_outputs(6901) <= not(inputs(0)) or (inputs(94));
    layer0_outputs(6902) <= not(inputs(39));
    layer0_outputs(6903) <= '1';
    layer0_outputs(6904) <= (inputs(192)) or (inputs(75));
    layer0_outputs(6905) <= not(inputs(6)) or (inputs(96));
    layer0_outputs(6906) <= '1';
    layer0_outputs(6907) <= not((inputs(20)) or (inputs(111)));
    layer0_outputs(6908) <= (inputs(11)) and not (inputs(131));
    layer0_outputs(6909) <= not(inputs(80)) or (inputs(41));
    layer0_outputs(6910) <= '0';
    layer0_outputs(6911) <= inputs(97);
    layer0_outputs(6912) <= not(inputs(26)) or (inputs(55));
    layer0_outputs(6913) <= (inputs(49)) and (inputs(71));
    layer0_outputs(6914) <= not(inputs(179));
    layer0_outputs(6915) <= not((inputs(66)) or (inputs(222)));
    layer0_outputs(6916) <= (inputs(65)) and (inputs(243));
    layer0_outputs(6917) <= inputs(88);
    layer0_outputs(6918) <= (inputs(246)) and (inputs(117));
    layer0_outputs(6919) <= not(inputs(121));
    layer0_outputs(6920) <= (inputs(148)) and not (inputs(27));
    layer0_outputs(6921) <= not(inputs(164));
    layer0_outputs(6922) <= '0';
    layer0_outputs(6923) <= (inputs(4)) and (inputs(156));
    layer0_outputs(6924) <= '0';
    layer0_outputs(6925) <= '1';
    layer0_outputs(6926) <= not(inputs(88)) or (inputs(104));
    layer0_outputs(6927) <= (inputs(139)) and (inputs(158));
    layer0_outputs(6928) <= inputs(43);
    layer0_outputs(6929) <= '0';
    layer0_outputs(6930) <= not(inputs(66));
    layer0_outputs(6931) <= inputs(151);
    layer0_outputs(6932) <= (inputs(238)) or (inputs(195));
    layer0_outputs(6933) <= not(inputs(113));
    layer0_outputs(6934) <= not(inputs(178));
    layer0_outputs(6935) <= (inputs(73)) and not (inputs(195));
    layer0_outputs(6936) <= not(inputs(179)) or (inputs(153));
    layer0_outputs(6937) <= not(inputs(0));
    layer0_outputs(6938) <= not(inputs(68));
    layer0_outputs(6939) <= (inputs(193)) and not (inputs(87));
    layer0_outputs(6940) <= not(inputs(1));
    layer0_outputs(6941) <= '1';
    layer0_outputs(6942) <= not(inputs(0)) or (inputs(225));
    layer0_outputs(6943) <= inputs(176);
    layer0_outputs(6944) <= (inputs(73)) or (inputs(132));
    layer0_outputs(6945) <= not((inputs(243)) or (inputs(152)));
    layer0_outputs(6946) <= not(inputs(19));
    layer0_outputs(6947) <= (inputs(249)) or (inputs(20));
    layer0_outputs(6948) <= not((inputs(46)) or (inputs(224)));
    layer0_outputs(6949) <= (inputs(21)) and (inputs(10));
    layer0_outputs(6950) <= not((inputs(229)) or (inputs(45)));
    layer0_outputs(6951) <= not(inputs(128));
    layer0_outputs(6952) <= not((inputs(14)) or (inputs(167)));
    layer0_outputs(6953) <= not((inputs(125)) and (inputs(15)));
    layer0_outputs(6954) <= (inputs(63)) and not (inputs(2));
    layer0_outputs(6955) <= inputs(3);
    layer0_outputs(6956) <= '1';
    layer0_outputs(6957) <= (inputs(44)) and (inputs(90));
    layer0_outputs(6958) <= not(inputs(244));
    layer0_outputs(6959) <= not((inputs(88)) and (inputs(149)));
    layer0_outputs(6960) <= not((inputs(36)) or (inputs(124)));
    layer0_outputs(6961) <= (inputs(61)) or (inputs(1));
    layer0_outputs(6962) <= not(inputs(38));
    layer0_outputs(6963) <= inputs(74);
    layer0_outputs(6964) <= not((inputs(89)) or (inputs(172)));
    layer0_outputs(6965) <= (inputs(198)) and not (inputs(46));
    layer0_outputs(6966) <= not((inputs(209)) xor (inputs(170)));
    layer0_outputs(6967) <= '0';
    layer0_outputs(6968) <= not((inputs(91)) or (inputs(2)));
    layer0_outputs(6969) <= (inputs(60)) and not (inputs(102));
    layer0_outputs(6970) <= '0';
    layer0_outputs(6971) <= not(inputs(2)) or (inputs(144));
    layer0_outputs(6972) <= not(inputs(38));
    layer0_outputs(6973) <= not((inputs(130)) or (inputs(14)));
    layer0_outputs(6974) <= not(inputs(121)) or (inputs(195));
    layer0_outputs(6975) <= (inputs(178)) and not (inputs(234));
    layer0_outputs(6976) <= '0';
    layer0_outputs(6977) <= (inputs(75)) and not (inputs(37));
    layer0_outputs(6978) <= not((inputs(116)) or (inputs(98)));
    layer0_outputs(6979) <= inputs(103);
    layer0_outputs(6980) <= not(inputs(112)) or (inputs(77));
    layer0_outputs(6981) <= not(inputs(40)) or (inputs(19));
    layer0_outputs(6982) <= (inputs(24)) and not (inputs(112));
    layer0_outputs(6983) <= not(inputs(138)) or (inputs(219));
    layer0_outputs(6984) <= '0';
    layer0_outputs(6985) <= not(inputs(222)) or (inputs(157));
    layer0_outputs(6986) <= inputs(178);
    layer0_outputs(6987) <= (inputs(100)) or (inputs(113));
    layer0_outputs(6988) <= not(inputs(234)) or (inputs(107));
    layer0_outputs(6989) <= not(inputs(14));
    layer0_outputs(6990) <= inputs(151);
    layer0_outputs(6991) <= (inputs(136)) and not (inputs(204));
    layer0_outputs(6992) <= '1';
    layer0_outputs(6993) <= '1';
    layer0_outputs(6994) <= '1';
    layer0_outputs(6995) <= (inputs(202)) and not (inputs(67));
    layer0_outputs(6996) <= inputs(51);
    layer0_outputs(6997) <= (inputs(252)) and not (inputs(54));
    layer0_outputs(6998) <= inputs(212);
    layer0_outputs(6999) <= inputs(230);
    layer0_outputs(7000) <= (inputs(84)) and not (inputs(167));
    layer0_outputs(7001) <= not((inputs(140)) and (inputs(10)));
    layer0_outputs(7002) <= '0';
    layer0_outputs(7003) <= '0';
    layer0_outputs(7004) <= inputs(85);
    layer0_outputs(7005) <= not(inputs(88)) or (inputs(232));
    layer0_outputs(7006) <= not(inputs(84));
    layer0_outputs(7007) <= not(inputs(93));
    layer0_outputs(7008) <= (inputs(104)) and not (inputs(127));
    layer0_outputs(7009) <= inputs(183);
    layer0_outputs(7010) <= (inputs(191)) and (inputs(32));
    layer0_outputs(7011) <= inputs(215);
    layer0_outputs(7012) <= not(inputs(138));
    layer0_outputs(7013) <= inputs(88);
    layer0_outputs(7014) <= '0';
    layer0_outputs(7015) <= not(inputs(169));
    layer0_outputs(7016) <= (inputs(191)) or (inputs(62));
    layer0_outputs(7017) <= not((inputs(12)) xor (inputs(46)));
    layer0_outputs(7018) <= '0';
    layer0_outputs(7019) <= inputs(104);
    layer0_outputs(7020) <= not((inputs(91)) and (inputs(62)));
    layer0_outputs(7021) <= not(inputs(97)) or (inputs(19));
    layer0_outputs(7022) <= inputs(10);
    layer0_outputs(7023) <= not((inputs(228)) or (inputs(52)));
    layer0_outputs(7024) <= '0';
    layer0_outputs(7025) <= not(inputs(194)) or (inputs(182));
    layer0_outputs(7026) <= not(inputs(180)) or (inputs(79));
    layer0_outputs(7027) <= not(inputs(187));
    layer0_outputs(7028) <= '1';
    layer0_outputs(7029) <= '0';
    layer0_outputs(7030) <= not(inputs(85));
    layer0_outputs(7031) <= inputs(88);
    layer0_outputs(7032) <= (inputs(37)) and not (inputs(243));
    layer0_outputs(7033) <= inputs(187);
    layer0_outputs(7034) <= (inputs(248)) or (inputs(129));
    layer0_outputs(7035) <= '0';
    layer0_outputs(7036) <= (inputs(229)) and (inputs(24));
    layer0_outputs(7037) <= (inputs(54)) and not (inputs(234));
    layer0_outputs(7038) <= not(inputs(100)) or (inputs(147));
    layer0_outputs(7039) <= inputs(231);
    layer0_outputs(7040) <= not(inputs(99));
    layer0_outputs(7041) <= (inputs(239)) xor (inputs(164));
    layer0_outputs(7042) <= (inputs(118)) or (inputs(60));
    layer0_outputs(7043) <= (inputs(0)) or (inputs(143));
    layer0_outputs(7044) <= not(inputs(179));
    layer0_outputs(7045) <= not(inputs(216)) or (inputs(169));
    layer0_outputs(7046) <= not(inputs(122));
    layer0_outputs(7047) <= '1';
    layer0_outputs(7048) <= inputs(232);
    layer0_outputs(7049) <= not(inputs(60)) or (inputs(239));
    layer0_outputs(7050) <= not(inputs(246)) or (inputs(98));
    layer0_outputs(7051) <= not(inputs(100));
    layer0_outputs(7052) <= '0';
    layer0_outputs(7053) <= not(inputs(80)) or (inputs(0));
    layer0_outputs(7054) <= not(inputs(37));
    layer0_outputs(7055) <= (inputs(242)) or (inputs(209));
    layer0_outputs(7056) <= inputs(105);
    layer0_outputs(7057) <= not(inputs(239));
    layer0_outputs(7058) <= inputs(118);
    layer0_outputs(7059) <= not(inputs(86));
    layer0_outputs(7060) <= '1';
    layer0_outputs(7061) <= inputs(74);
    layer0_outputs(7062) <= not(inputs(215));
    layer0_outputs(7063) <= not(inputs(226));
    layer0_outputs(7064) <= (inputs(59)) or (inputs(63));
    layer0_outputs(7065) <= not(inputs(232));
    layer0_outputs(7066) <= not((inputs(186)) or (inputs(228)));
    layer0_outputs(7067) <= not(inputs(159));
    layer0_outputs(7068) <= (inputs(7)) or (inputs(101));
    layer0_outputs(7069) <= not(inputs(118));
    layer0_outputs(7070) <= not(inputs(127)) or (inputs(55));
    layer0_outputs(7071) <= inputs(173);
    layer0_outputs(7072) <= (inputs(131)) and not (inputs(150));
    layer0_outputs(7073) <= (inputs(122)) and not (inputs(199));
    layer0_outputs(7074) <= (inputs(190)) or (inputs(126));
    layer0_outputs(7075) <= not((inputs(196)) and (inputs(203)));
    layer0_outputs(7076) <= inputs(84);
    layer0_outputs(7077) <= (inputs(37)) and not (inputs(161));
    layer0_outputs(7078) <= not((inputs(199)) and (inputs(16)));
    layer0_outputs(7079) <= not(inputs(163));
    layer0_outputs(7080) <= (inputs(20)) or (inputs(28));
    layer0_outputs(7081) <= not((inputs(247)) xor (inputs(216)));
    layer0_outputs(7082) <= (inputs(151)) xor (inputs(186));
    layer0_outputs(7083) <= not(inputs(105));
    layer0_outputs(7084) <= (inputs(111)) or (inputs(69));
    layer0_outputs(7085) <= not((inputs(104)) or (inputs(188)));
    layer0_outputs(7086) <= '0';
    layer0_outputs(7087) <= not(inputs(30)) or (inputs(55));
    layer0_outputs(7088) <= (inputs(206)) xor (inputs(238));
    layer0_outputs(7089) <= not(inputs(177));
    layer0_outputs(7090) <= not((inputs(86)) and (inputs(92)));
    layer0_outputs(7091) <= '1';
    layer0_outputs(7092) <= '1';
    layer0_outputs(7093) <= '0';
    layer0_outputs(7094) <= inputs(245);
    layer0_outputs(7095) <= inputs(34);
    layer0_outputs(7096) <= not(inputs(70)) or (inputs(18));
    layer0_outputs(7097) <= not((inputs(87)) or (inputs(183)));
    layer0_outputs(7098) <= (inputs(207)) or (inputs(179));
    layer0_outputs(7099) <= '0';
    layer0_outputs(7100) <= '0';
    layer0_outputs(7101) <= (inputs(23)) xor (inputs(55));
    layer0_outputs(7102) <= (inputs(223)) and (inputs(11));
    layer0_outputs(7103) <= not((inputs(110)) and (inputs(250)));
    layer0_outputs(7104) <= not(inputs(133));
    layer0_outputs(7105) <= not((inputs(8)) xor (inputs(55)));
    layer0_outputs(7106) <= not(inputs(170));
    layer0_outputs(7107) <= (inputs(175)) or (inputs(210));
    layer0_outputs(7108) <= not(inputs(24));
    layer0_outputs(7109) <= '1';
    layer0_outputs(7110) <= not((inputs(139)) or (inputs(2)));
    layer0_outputs(7111) <= not(inputs(73)) or (inputs(42));
    layer0_outputs(7112) <= (inputs(253)) and not (inputs(18));
    layer0_outputs(7113) <= not(inputs(107)) or (inputs(46));
    layer0_outputs(7114) <= not(inputs(136));
    layer0_outputs(7115) <= '0';
    layer0_outputs(7116) <= not(inputs(35));
    layer0_outputs(7117) <= inputs(23);
    layer0_outputs(7118) <= not(inputs(212)) or (inputs(48));
    layer0_outputs(7119) <= not(inputs(149));
    layer0_outputs(7120) <= (inputs(107)) or (inputs(108));
    layer0_outputs(7121) <= not(inputs(94));
    layer0_outputs(7122) <= '1';
    layer0_outputs(7123) <= inputs(230);
    layer0_outputs(7124) <= (inputs(112)) and not (inputs(204));
    layer0_outputs(7125) <= not(inputs(96));
    layer0_outputs(7126) <= '1';
    layer0_outputs(7127) <= '0';
    layer0_outputs(7128) <= not(inputs(115)) or (inputs(238));
    layer0_outputs(7129) <= inputs(230);
    layer0_outputs(7130) <= (inputs(12)) xor (inputs(255));
    layer0_outputs(7131) <= (inputs(220)) and not (inputs(36));
    layer0_outputs(7132) <= not(inputs(232)) or (inputs(47));
    layer0_outputs(7133) <= '0';
    layer0_outputs(7134) <= not((inputs(195)) and (inputs(88)));
    layer0_outputs(7135) <= not(inputs(199));
    layer0_outputs(7136) <= not(inputs(162)) or (inputs(91));
    layer0_outputs(7137) <= inputs(160);
    layer0_outputs(7138) <= (inputs(71)) or (inputs(43));
    layer0_outputs(7139) <= inputs(160);
    layer0_outputs(7140) <= not(inputs(138)) or (inputs(145));
    layer0_outputs(7141) <= not(inputs(220));
    layer0_outputs(7142) <= (inputs(24)) or (inputs(39));
    layer0_outputs(7143) <= '1';
    layer0_outputs(7144) <= not(inputs(225));
    layer0_outputs(7145) <= inputs(114);
    layer0_outputs(7146) <= not(inputs(16)) or (inputs(160));
    layer0_outputs(7147) <= inputs(37);
    layer0_outputs(7148) <= (inputs(153)) and (inputs(78));
    layer0_outputs(7149) <= not(inputs(223)) or (inputs(133));
    layer0_outputs(7150) <= (inputs(92)) or (inputs(88));
    layer0_outputs(7151) <= not(inputs(13)) or (inputs(178));
    layer0_outputs(7152) <= not((inputs(69)) or (inputs(79)));
    layer0_outputs(7153) <= (inputs(74)) and not (inputs(132));
    layer0_outputs(7154) <= (inputs(34)) or (inputs(242));
    layer0_outputs(7155) <= '1';
    layer0_outputs(7156) <= not((inputs(21)) or (inputs(248)));
    layer0_outputs(7157) <= (inputs(210)) and not (inputs(97));
    layer0_outputs(7158) <= '0';
    layer0_outputs(7159) <= (inputs(226)) and not (inputs(240));
    layer0_outputs(7160) <= (inputs(213)) or (inputs(166));
    layer0_outputs(7161) <= '0';
    layer0_outputs(7162) <= (inputs(106)) and not (inputs(101));
    layer0_outputs(7163) <= (inputs(175)) and (inputs(240));
    layer0_outputs(7164) <= not(inputs(147));
    layer0_outputs(7165) <= not(inputs(206));
    layer0_outputs(7166) <= (inputs(133)) and not (inputs(73));
    layer0_outputs(7167) <= not((inputs(233)) or (inputs(79)));
    layer0_outputs(7168) <= '1';
    layer0_outputs(7169) <= '1';
    layer0_outputs(7170) <= '0';
    layer0_outputs(7171) <= (inputs(94)) and not (inputs(50));
    layer0_outputs(7172) <= inputs(61);
    layer0_outputs(7173) <= '1';
    layer0_outputs(7174) <= not(inputs(181)) or (inputs(78));
    layer0_outputs(7175) <= (inputs(5)) and not (inputs(205));
    layer0_outputs(7176) <= inputs(215);
    layer0_outputs(7177) <= not(inputs(183));
    layer0_outputs(7178) <= '0';
    layer0_outputs(7179) <= (inputs(253)) and not (inputs(76));
    layer0_outputs(7180) <= inputs(174);
    layer0_outputs(7181) <= inputs(242);
    layer0_outputs(7182) <= inputs(106);
    layer0_outputs(7183) <= not(inputs(168)) or (inputs(231));
    layer0_outputs(7184) <= not(inputs(38));
    layer0_outputs(7185) <= not(inputs(131)) or (inputs(28));
    layer0_outputs(7186) <= '1';
    layer0_outputs(7187) <= not((inputs(54)) or (inputs(68)));
    layer0_outputs(7188) <= (inputs(141)) and not (inputs(35));
    layer0_outputs(7189) <= '0';
    layer0_outputs(7190) <= not(inputs(147)) or (inputs(199));
    layer0_outputs(7191) <= '0';
    layer0_outputs(7192) <= (inputs(34)) and not (inputs(249));
    layer0_outputs(7193) <= not(inputs(62));
    layer0_outputs(7194) <= not(inputs(42)) or (inputs(252));
    layer0_outputs(7195) <= not(inputs(160));
    layer0_outputs(7196) <= (inputs(149)) and not (inputs(11));
    layer0_outputs(7197) <= (inputs(22)) and not (inputs(205));
    layer0_outputs(7198) <= inputs(136);
    layer0_outputs(7199) <= (inputs(51)) and not (inputs(82));
    layer0_outputs(7200) <= '0';
    layer0_outputs(7201) <= (inputs(5)) or (inputs(1));
    layer0_outputs(7202) <= not(inputs(102));
    layer0_outputs(7203) <= inputs(238);
    layer0_outputs(7204) <= '1';
    layer0_outputs(7205) <= not(inputs(122));
    layer0_outputs(7206) <= inputs(39);
    layer0_outputs(7207) <= not(inputs(76));
    layer0_outputs(7208) <= '1';
    layer0_outputs(7209) <= '0';
    layer0_outputs(7210) <= (inputs(163)) or (inputs(89));
    layer0_outputs(7211) <= '1';
    layer0_outputs(7212) <= not(inputs(132)) or (inputs(225));
    layer0_outputs(7213) <= (inputs(60)) and not (inputs(180));
    layer0_outputs(7214) <= (inputs(116)) and not (inputs(171));
    layer0_outputs(7215) <= not((inputs(122)) and (inputs(194)));
    layer0_outputs(7216) <= not(inputs(104));
    layer0_outputs(7217) <= inputs(120);
    layer0_outputs(7218) <= (inputs(144)) xor (inputs(240));
    layer0_outputs(7219) <= not((inputs(97)) or (inputs(101)));
    layer0_outputs(7220) <= (inputs(225)) or (inputs(128));
    layer0_outputs(7221) <= '1';
    layer0_outputs(7222) <= '0';
    layer0_outputs(7223) <= not(inputs(16));
    layer0_outputs(7224) <= not((inputs(110)) and (inputs(93)));
    layer0_outputs(7225) <= (inputs(212)) or (inputs(242));
    layer0_outputs(7226) <= not(inputs(62)) or (inputs(110));
    layer0_outputs(7227) <= inputs(148);
    layer0_outputs(7228) <= not((inputs(178)) and (inputs(59)));
    layer0_outputs(7229) <= inputs(1);
    layer0_outputs(7230) <= '0';
    layer0_outputs(7231) <= not(inputs(118)) or (inputs(148));
    layer0_outputs(7232) <= inputs(223);
    layer0_outputs(7233) <= (inputs(248)) xor (inputs(125));
    layer0_outputs(7234) <= not((inputs(221)) and (inputs(16)));
    layer0_outputs(7235) <= inputs(23);
    layer0_outputs(7236) <= inputs(149);
    layer0_outputs(7237) <= not(inputs(120));
    layer0_outputs(7238) <= (inputs(236)) and not (inputs(38));
    layer0_outputs(7239) <= not(inputs(225)) or (inputs(78));
    layer0_outputs(7240) <= not(inputs(245));
    layer0_outputs(7241) <= not(inputs(17));
    layer0_outputs(7242) <= not((inputs(33)) and (inputs(94)));
    layer0_outputs(7243) <= not(inputs(98));
    layer0_outputs(7244) <= not(inputs(199));
    layer0_outputs(7245) <= not((inputs(233)) or (inputs(219)));
    layer0_outputs(7246) <= '1';
    layer0_outputs(7247) <= not((inputs(106)) or (inputs(123)));
    layer0_outputs(7248) <= not(inputs(157)) or (inputs(168));
    layer0_outputs(7249) <= inputs(114);
    layer0_outputs(7250) <= (inputs(192)) or (inputs(194));
    layer0_outputs(7251) <= not((inputs(13)) or (inputs(3)));
    layer0_outputs(7252) <= not(inputs(112));
    layer0_outputs(7253) <= not(inputs(229));
    layer0_outputs(7254) <= inputs(151);
    layer0_outputs(7255) <= '0';
    layer0_outputs(7256) <= (inputs(15)) and (inputs(15));
    layer0_outputs(7257) <= '0';
    layer0_outputs(7258) <= inputs(8);
    layer0_outputs(7259) <= not(inputs(168));
    layer0_outputs(7260) <= '1';
    layer0_outputs(7261) <= inputs(230);
    layer0_outputs(7262) <= (inputs(80)) and not (inputs(172));
    layer0_outputs(7263) <= '0';
    layer0_outputs(7264) <= '0';
    layer0_outputs(7265) <= inputs(63);
    layer0_outputs(7266) <= (inputs(12)) and not (inputs(117));
    layer0_outputs(7267) <= not(inputs(248)) or (inputs(33));
    layer0_outputs(7268) <= inputs(140);
    layer0_outputs(7269) <= not((inputs(226)) and (inputs(169)));
    layer0_outputs(7270) <= not(inputs(51));
    layer0_outputs(7271) <= inputs(62);
    layer0_outputs(7272) <= (inputs(190)) or (inputs(63));
    layer0_outputs(7273) <= (inputs(145)) or (inputs(225));
    layer0_outputs(7274) <= inputs(78);
    layer0_outputs(7275) <= not(inputs(49)) or (inputs(160));
    layer0_outputs(7276) <= inputs(248);
    layer0_outputs(7277) <= not(inputs(168)) or (inputs(76));
    layer0_outputs(7278) <= not(inputs(79));
    layer0_outputs(7279) <= '0';
    layer0_outputs(7280) <= (inputs(55)) and not (inputs(136));
    layer0_outputs(7281) <= inputs(83);
    layer0_outputs(7282) <= not(inputs(130)) or (inputs(142));
    layer0_outputs(7283) <= (inputs(27)) and not (inputs(194));
    layer0_outputs(7284) <= not((inputs(150)) or (inputs(199)));
    layer0_outputs(7285) <= '1';
    layer0_outputs(7286) <= not(inputs(41));
    layer0_outputs(7287) <= inputs(164);
    layer0_outputs(7288) <= not((inputs(88)) or (inputs(47)));
    layer0_outputs(7289) <= not(inputs(185));
    layer0_outputs(7290) <= not((inputs(240)) or (inputs(20)));
    layer0_outputs(7291) <= (inputs(188)) or (inputs(187));
    layer0_outputs(7292) <= not((inputs(5)) xor (inputs(142)));
    layer0_outputs(7293) <= (inputs(18)) and not (inputs(76));
    layer0_outputs(7294) <= '0';
    layer0_outputs(7295) <= not(inputs(198)) or (inputs(62));
    layer0_outputs(7296) <= (inputs(130)) and (inputs(13));
    layer0_outputs(7297) <= '0';
    layer0_outputs(7298) <= not(inputs(130));
    layer0_outputs(7299) <= inputs(127);
    layer0_outputs(7300) <= not((inputs(135)) and (inputs(180)));
    layer0_outputs(7301) <= '1';
    layer0_outputs(7302) <= '1';
    layer0_outputs(7303) <= not(inputs(196)) or (inputs(213));
    layer0_outputs(7304) <= (inputs(32)) and (inputs(42));
    layer0_outputs(7305) <= (inputs(215)) or (inputs(220));
    layer0_outputs(7306) <= inputs(171);
    layer0_outputs(7307) <= '1';
    layer0_outputs(7308) <= not((inputs(197)) or (inputs(132)));
    layer0_outputs(7309) <= not(inputs(178)) or (inputs(40));
    layer0_outputs(7310) <= (inputs(28)) and not (inputs(131));
    layer0_outputs(7311) <= not(inputs(22)) or (inputs(83));
    layer0_outputs(7312) <= '0';
    layer0_outputs(7313) <= (inputs(186)) and not (inputs(139));
    layer0_outputs(7314) <= (inputs(33)) and not (inputs(224));
    layer0_outputs(7315) <= inputs(88);
    layer0_outputs(7316) <= (inputs(221)) and (inputs(165));
    layer0_outputs(7317) <= inputs(201);
    layer0_outputs(7318) <= inputs(207);
    layer0_outputs(7319) <= (inputs(189)) and not (inputs(88));
    layer0_outputs(7320) <= not((inputs(196)) or (inputs(227)));
    layer0_outputs(7321) <= not((inputs(243)) or (inputs(246)));
    layer0_outputs(7322) <= '1';
    layer0_outputs(7323) <= not((inputs(161)) xor (inputs(37)));
    layer0_outputs(7324) <= not(inputs(81));
    layer0_outputs(7325) <= (inputs(202)) xor (inputs(17));
    layer0_outputs(7326) <= '1';
    layer0_outputs(7327) <= not((inputs(94)) xor (inputs(207)));
    layer0_outputs(7328) <= inputs(52);
    layer0_outputs(7329) <= '0';
    layer0_outputs(7330) <= not(inputs(233)) or (inputs(94));
    layer0_outputs(7331) <= (inputs(175)) or (inputs(212));
    layer0_outputs(7332) <= not((inputs(63)) xor (inputs(77)));
    layer0_outputs(7333) <= inputs(74);
    layer0_outputs(7334) <= (inputs(42)) or (inputs(46));
    layer0_outputs(7335) <= (inputs(148)) and not (inputs(224));
    layer0_outputs(7336) <= not(inputs(172));
    layer0_outputs(7337) <= not((inputs(114)) or (inputs(52)));
    layer0_outputs(7338) <= not(inputs(157)) or (inputs(249));
    layer0_outputs(7339) <= not((inputs(65)) and (inputs(69)));
    layer0_outputs(7340) <= (inputs(226)) or (inputs(83));
    layer0_outputs(7341) <= not(inputs(118));
    layer0_outputs(7342) <= inputs(241);
    layer0_outputs(7343) <= '0';
    layer0_outputs(7344) <= inputs(8);
    layer0_outputs(7345) <= '1';
    layer0_outputs(7346) <= not(inputs(158));
    layer0_outputs(7347) <= inputs(163);
    layer0_outputs(7348) <= not(inputs(57)) or (inputs(64));
    layer0_outputs(7349) <= inputs(76);
    layer0_outputs(7350) <= inputs(244);
    layer0_outputs(7351) <= inputs(62);
    layer0_outputs(7352) <= not(inputs(230)) or (inputs(91));
    layer0_outputs(7353) <= not(inputs(180));
    layer0_outputs(7354) <= inputs(246);
    layer0_outputs(7355) <= inputs(51);
    layer0_outputs(7356) <= not(inputs(178));
    layer0_outputs(7357) <= (inputs(92)) and not (inputs(37));
    layer0_outputs(7358) <= not((inputs(60)) xor (inputs(193)));
    layer0_outputs(7359) <= '0';
    layer0_outputs(7360) <= not(inputs(227));
    layer0_outputs(7361) <= not(inputs(228));
    layer0_outputs(7362) <= (inputs(52)) or (inputs(26));
    layer0_outputs(7363) <= not(inputs(16));
    layer0_outputs(7364) <= not((inputs(121)) and (inputs(5)));
    layer0_outputs(7365) <= '1';
    layer0_outputs(7366) <= not(inputs(150));
    layer0_outputs(7367) <= not((inputs(18)) and (inputs(24)));
    layer0_outputs(7368) <= (inputs(192)) or (inputs(230));
    layer0_outputs(7369) <= not((inputs(188)) and (inputs(133)));
    layer0_outputs(7370) <= '0';
    layer0_outputs(7371) <= inputs(171);
    layer0_outputs(7372) <= (inputs(69)) and (inputs(75));
    layer0_outputs(7373) <= not(inputs(242));
    layer0_outputs(7374) <= not((inputs(167)) or (inputs(34)));
    layer0_outputs(7375) <= not((inputs(68)) or (inputs(127)));
    layer0_outputs(7376) <= not(inputs(101)) or (inputs(62));
    layer0_outputs(7377) <= not(inputs(25)) or (inputs(181));
    layer0_outputs(7378) <= not((inputs(126)) and (inputs(154)));
    layer0_outputs(7379) <= '0';
    layer0_outputs(7380) <= not((inputs(192)) and (inputs(4)));
    layer0_outputs(7381) <= '1';
    layer0_outputs(7382) <= inputs(87);
    layer0_outputs(7383) <= not((inputs(177)) or (inputs(127)));
    layer0_outputs(7384) <= not(inputs(85));
    layer0_outputs(7385) <= not(inputs(113));
    layer0_outputs(7386) <= '1';
    layer0_outputs(7387) <= '1';
    layer0_outputs(7388) <= (inputs(58)) and not (inputs(47));
    layer0_outputs(7389) <= not((inputs(174)) xor (inputs(153)));
    layer0_outputs(7390) <= (inputs(62)) xor (inputs(15));
    layer0_outputs(7391) <= not(inputs(192));
    layer0_outputs(7392) <= not(inputs(26));
    layer0_outputs(7393) <= inputs(124);
    layer0_outputs(7394) <= not((inputs(24)) or (inputs(174)));
    layer0_outputs(7395) <= not(inputs(151)) or (inputs(45));
    layer0_outputs(7396) <= not((inputs(5)) and (inputs(128)));
    layer0_outputs(7397) <= (inputs(22)) and (inputs(243));
    layer0_outputs(7398) <= not(inputs(29)) or (inputs(98));
    layer0_outputs(7399) <= not(inputs(5)) or (inputs(216));
    layer0_outputs(7400) <= not(inputs(212)) or (inputs(40));
    layer0_outputs(7401) <= not(inputs(188));
    layer0_outputs(7402) <= not(inputs(19));
    layer0_outputs(7403) <= not((inputs(239)) xor (inputs(194)));
    layer0_outputs(7404) <= not(inputs(51));
    layer0_outputs(7405) <= (inputs(174)) and (inputs(12));
    layer0_outputs(7406) <= inputs(185);
    layer0_outputs(7407) <= inputs(72);
    layer0_outputs(7408) <= not(inputs(61));
    layer0_outputs(7409) <= '1';
    layer0_outputs(7410) <= not(inputs(64)) or (inputs(49));
    layer0_outputs(7411) <= not(inputs(221));
    layer0_outputs(7412) <= not((inputs(145)) or (inputs(90)));
    layer0_outputs(7413) <= not((inputs(29)) or (inputs(188)));
    layer0_outputs(7414) <= '0';
    layer0_outputs(7415) <= '1';
    layer0_outputs(7416) <= '1';
    layer0_outputs(7417) <= not(inputs(252)) or (inputs(26));
    layer0_outputs(7418) <= not(inputs(79));
    layer0_outputs(7419) <= not(inputs(246));
    layer0_outputs(7420) <= not(inputs(151)) or (inputs(191));
    layer0_outputs(7421) <= (inputs(51)) or (inputs(97));
    layer0_outputs(7422) <= not(inputs(255));
    layer0_outputs(7423) <= (inputs(23)) and not (inputs(218));
    layer0_outputs(7424) <= not(inputs(247));
    layer0_outputs(7425) <= inputs(195);
    layer0_outputs(7426) <= not((inputs(56)) and (inputs(241)));
    layer0_outputs(7427) <= not((inputs(38)) xor (inputs(143)));
    layer0_outputs(7428) <= not((inputs(109)) or (inputs(140)));
    layer0_outputs(7429) <= (inputs(213)) and not (inputs(68));
    layer0_outputs(7430) <= not((inputs(35)) or (inputs(131)));
    layer0_outputs(7431) <= not((inputs(1)) or (inputs(166)));
    layer0_outputs(7432) <= not(inputs(134));
    layer0_outputs(7433) <= (inputs(1)) or (inputs(16));
    layer0_outputs(7434) <= inputs(62);
    layer0_outputs(7435) <= (inputs(105)) and (inputs(76));
    layer0_outputs(7436) <= inputs(156);
    layer0_outputs(7437) <= not(inputs(102)) or (inputs(121));
    layer0_outputs(7438) <= '1';
    layer0_outputs(7439) <= inputs(58);
    layer0_outputs(7440) <= inputs(207);
    layer0_outputs(7441) <= inputs(39);
    layer0_outputs(7442) <= (inputs(25)) and not (inputs(147));
    layer0_outputs(7443) <= not((inputs(46)) xor (inputs(194)));
    layer0_outputs(7444) <= not((inputs(134)) and (inputs(216)));
    layer0_outputs(7445) <= not((inputs(20)) and (inputs(69)));
    layer0_outputs(7446) <= not(inputs(224));
    layer0_outputs(7447) <= '1';
    layer0_outputs(7448) <= not((inputs(51)) or (inputs(201)));
    layer0_outputs(7449) <= not(inputs(4)) or (inputs(100));
    layer0_outputs(7450) <= inputs(181);
    layer0_outputs(7451) <= not(inputs(247));
    layer0_outputs(7452) <= '0';
    layer0_outputs(7453) <= (inputs(127)) and not (inputs(138));
    layer0_outputs(7454) <= (inputs(207)) xor (inputs(238));
    layer0_outputs(7455) <= inputs(239);
    layer0_outputs(7456) <= not(inputs(66));
    layer0_outputs(7457) <= '0';
    layer0_outputs(7458) <= (inputs(241)) and not (inputs(87));
    layer0_outputs(7459) <= (inputs(125)) or (inputs(157));
    layer0_outputs(7460) <= not(inputs(205));
    layer0_outputs(7461) <= not(inputs(252)) or (inputs(184));
    layer0_outputs(7462) <= not(inputs(215)) or (inputs(236));
    layer0_outputs(7463) <= (inputs(181)) and not (inputs(73));
    layer0_outputs(7464) <= not(inputs(26));
    layer0_outputs(7465) <= '1';
    layer0_outputs(7466) <= (inputs(216)) and (inputs(171));
    layer0_outputs(7467) <= '0';
    layer0_outputs(7468) <= inputs(121);
    layer0_outputs(7469) <= (inputs(40)) and not (inputs(179));
    layer0_outputs(7470) <= not(inputs(168));
    layer0_outputs(7471) <= not(inputs(109));
    layer0_outputs(7472) <= (inputs(193)) and not (inputs(145));
    layer0_outputs(7473) <= not((inputs(11)) or (inputs(33)));
    layer0_outputs(7474) <= (inputs(202)) and (inputs(30));
    layer0_outputs(7475) <= '0';
    layer0_outputs(7476) <= not(inputs(254)) or (inputs(130));
    layer0_outputs(7477) <= inputs(172);
    layer0_outputs(7478) <= (inputs(221)) and not (inputs(138));
    layer0_outputs(7479) <= not((inputs(211)) and (inputs(40)));
    layer0_outputs(7480) <= (inputs(208)) and (inputs(3));
    layer0_outputs(7481) <= (inputs(106)) and not (inputs(22));
    layer0_outputs(7482) <= (inputs(115)) or (inputs(216));
    layer0_outputs(7483) <= '0';
    layer0_outputs(7484) <= '1';
    layer0_outputs(7485) <= '1';
    layer0_outputs(7486) <= '1';
    layer0_outputs(7487) <= inputs(183);
    layer0_outputs(7488) <= not(inputs(155));
    layer0_outputs(7489) <= not((inputs(212)) xor (inputs(32)));
    layer0_outputs(7490) <= inputs(228);
    layer0_outputs(7491) <= '1';
    layer0_outputs(7492) <= '0';
    layer0_outputs(7493) <= not(inputs(31));
    layer0_outputs(7494) <= (inputs(207)) and not (inputs(186));
    layer0_outputs(7495) <= not(inputs(171));
    layer0_outputs(7496) <= '1';
    layer0_outputs(7497) <= '0';
    layer0_outputs(7498) <= not(inputs(13)) or (inputs(115));
    layer0_outputs(7499) <= not(inputs(143));
    layer0_outputs(7500) <= not(inputs(111));
    layer0_outputs(7501) <= not((inputs(220)) or (inputs(178)));
    layer0_outputs(7502) <= inputs(86);
    layer0_outputs(7503) <= not(inputs(63)) or (inputs(139));
    layer0_outputs(7504) <= inputs(229);
    layer0_outputs(7505) <= not((inputs(173)) and (inputs(41)));
    layer0_outputs(7506) <= (inputs(60)) xor (inputs(58));
    layer0_outputs(7507) <= (inputs(28)) and not (inputs(199));
    layer0_outputs(7508) <= not(inputs(45)) or (inputs(200));
    layer0_outputs(7509) <= not(inputs(106));
    layer0_outputs(7510) <= not(inputs(84)) or (inputs(142));
    layer0_outputs(7511) <= not((inputs(138)) and (inputs(190)));
    layer0_outputs(7512) <= (inputs(190)) and not (inputs(124));
    layer0_outputs(7513) <= '1';
    layer0_outputs(7514) <= not(inputs(110));
    layer0_outputs(7515) <= not(inputs(243)) or (inputs(146));
    layer0_outputs(7516) <= (inputs(36)) or (inputs(45));
    layer0_outputs(7517) <= (inputs(144)) and (inputs(236));
    layer0_outputs(7518) <= not((inputs(68)) or (inputs(79)));
    layer0_outputs(7519) <= not(inputs(151));
    layer0_outputs(7520) <= not((inputs(69)) or (inputs(207)));
    layer0_outputs(7521) <= (inputs(111)) xor (inputs(152));
    layer0_outputs(7522) <= inputs(159);
    layer0_outputs(7523) <= not(inputs(205));
    layer0_outputs(7524) <= not(inputs(94));
    layer0_outputs(7525) <= not((inputs(221)) and (inputs(75)));
    layer0_outputs(7526) <= (inputs(99)) and not (inputs(203));
    layer0_outputs(7527) <= '1';
    layer0_outputs(7528) <= inputs(177);
    layer0_outputs(7529) <= not(inputs(49));
    layer0_outputs(7530) <= (inputs(209)) and not (inputs(10));
    layer0_outputs(7531) <= (inputs(157)) or (inputs(100));
    layer0_outputs(7532) <= not((inputs(12)) xor (inputs(236)));
    layer0_outputs(7533) <= inputs(212);
    layer0_outputs(7534) <= (inputs(212)) and not (inputs(246));
    layer0_outputs(7535) <= (inputs(161)) or (inputs(185));
    layer0_outputs(7536) <= not(inputs(232));
    layer0_outputs(7537) <= (inputs(247)) and not (inputs(29));
    layer0_outputs(7538) <= not(inputs(248)) or (inputs(217));
    layer0_outputs(7539) <= inputs(105);
    layer0_outputs(7540) <= not(inputs(196));
    layer0_outputs(7541) <= not(inputs(64)) or (inputs(93));
    layer0_outputs(7542) <= not((inputs(27)) or (inputs(85)));
    layer0_outputs(7543) <= (inputs(68)) and (inputs(13));
    layer0_outputs(7544) <= not(inputs(187)) or (inputs(2));
    layer0_outputs(7545) <= inputs(104);
    layer0_outputs(7546) <= (inputs(54)) or (inputs(63));
    layer0_outputs(7547) <= not(inputs(7)) or (inputs(113));
    layer0_outputs(7548) <= not((inputs(176)) or (inputs(161)));
    layer0_outputs(7549) <= '1';
    layer0_outputs(7550) <= not((inputs(224)) or (inputs(3)));
    layer0_outputs(7551) <= not(inputs(56));
    layer0_outputs(7552) <= (inputs(145)) and (inputs(167));
    layer0_outputs(7553) <= (inputs(120)) and not (inputs(138));
    layer0_outputs(7554) <= (inputs(103)) and (inputs(194));
    layer0_outputs(7555) <= inputs(93);
    layer0_outputs(7556) <= not(inputs(115));
    layer0_outputs(7557) <= '1';
    layer0_outputs(7558) <= (inputs(39)) or (inputs(80));
    layer0_outputs(7559) <= (inputs(255)) and not (inputs(29));
    layer0_outputs(7560) <= not((inputs(224)) or (inputs(114)));
    layer0_outputs(7561) <= inputs(135);
    layer0_outputs(7562) <= not((inputs(135)) and (inputs(67)));
    layer0_outputs(7563) <= not((inputs(240)) and (inputs(102)));
    layer0_outputs(7564) <= not(inputs(86));
    layer0_outputs(7565) <= not(inputs(139)) or (inputs(224));
    layer0_outputs(7566) <= (inputs(161)) or (inputs(146));
    layer0_outputs(7567) <= not(inputs(23));
    layer0_outputs(7568) <= not((inputs(161)) and (inputs(210)));
    layer0_outputs(7569) <= not(inputs(52));
    layer0_outputs(7570) <= not(inputs(49));
    layer0_outputs(7571) <= not((inputs(233)) and (inputs(132)));
    layer0_outputs(7572) <= inputs(195);
    layer0_outputs(7573) <= (inputs(247)) or (inputs(129));
    layer0_outputs(7574) <= inputs(177);
    layer0_outputs(7575) <= not((inputs(178)) or (inputs(251)));
    layer0_outputs(7576) <= not((inputs(123)) or (inputs(32)));
    layer0_outputs(7577) <= (inputs(191)) and not (inputs(170));
    layer0_outputs(7578) <= inputs(136);
    layer0_outputs(7579) <= inputs(198);
    layer0_outputs(7580) <= (inputs(58)) and (inputs(45));
    layer0_outputs(7581) <= not((inputs(189)) or (inputs(198)));
    layer0_outputs(7582) <= '1';
    layer0_outputs(7583) <= not(inputs(131));
    layer0_outputs(7584) <= not(inputs(183));
    layer0_outputs(7585) <= not(inputs(195)) or (inputs(36));
    layer0_outputs(7586) <= (inputs(67)) and not (inputs(8));
    layer0_outputs(7587) <= not(inputs(249));
    layer0_outputs(7588) <= (inputs(194)) and (inputs(45));
    layer0_outputs(7589) <= not(inputs(107)) or (inputs(248));
    layer0_outputs(7590) <= (inputs(202)) or (inputs(146));
    layer0_outputs(7591) <= (inputs(179)) or (inputs(194));
    layer0_outputs(7592) <= '0';
    layer0_outputs(7593) <= not((inputs(44)) and (inputs(48)));
    layer0_outputs(7594) <= not(inputs(180)) or (inputs(207));
    layer0_outputs(7595) <= (inputs(214)) and not (inputs(216));
    layer0_outputs(7596) <= not(inputs(111));
    layer0_outputs(7597) <= not(inputs(205));
    layer0_outputs(7598) <= not((inputs(103)) xor (inputs(26)));
    layer0_outputs(7599) <= inputs(17);
    layer0_outputs(7600) <= not((inputs(113)) xor (inputs(152)));
    layer0_outputs(7601) <= not((inputs(134)) or (inputs(19)));
    layer0_outputs(7602) <= not((inputs(161)) xor (inputs(25)));
    layer0_outputs(7603) <= '0';
    layer0_outputs(7604) <= (inputs(227)) or (inputs(81));
    layer0_outputs(7605) <= (inputs(125)) and not (inputs(37));
    layer0_outputs(7606) <= (inputs(243)) and not (inputs(238));
    layer0_outputs(7607) <= not(inputs(149));
    layer0_outputs(7608) <= not((inputs(192)) or (inputs(248)));
    layer0_outputs(7609) <= not((inputs(168)) xor (inputs(240)));
    layer0_outputs(7610) <= inputs(207);
    layer0_outputs(7611) <= inputs(136);
    layer0_outputs(7612) <= inputs(179);
    layer0_outputs(7613) <= '0';
    layer0_outputs(7614) <= (inputs(225)) or (inputs(109));
    layer0_outputs(7615) <= (inputs(28)) and not (inputs(226));
    layer0_outputs(7616) <= not((inputs(235)) or (inputs(240)));
    layer0_outputs(7617) <= not(inputs(159));
    layer0_outputs(7618) <= not(inputs(107)) or (inputs(186));
    layer0_outputs(7619) <= (inputs(94)) xor (inputs(223));
    layer0_outputs(7620) <= not(inputs(199)) or (inputs(179));
    layer0_outputs(7621) <= (inputs(67)) or (inputs(181));
    layer0_outputs(7622) <= not(inputs(162));
    layer0_outputs(7623) <= '0';
    layer0_outputs(7624) <= '0';
    layer0_outputs(7625) <= (inputs(221)) and not (inputs(210));
    layer0_outputs(7626) <= not(inputs(76)) or (inputs(214));
    layer0_outputs(7627) <= not(inputs(66)) or (inputs(41));
    layer0_outputs(7628) <= (inputs(154)) or (inputs(138));
    layer0_outputs(7629) <= inputs(15);
    layer0_outputs(7630) <= (inputs(224)) or (inputs(248));
    layer0_outputs(7631) <= not(inputs(62));
    layer0_outputs(7632) <= not((inputs(102)) xor (inputs(231)));
    layer0_outputs(7633) <= inputs(100);
    layer0_outputs(7634) <= inputs(92);
    layer0_outputs(7635) <= not((inputs(208)) xor (inputs(145)));
    layer0_outputs(7636) <= not(inputs(94));
    layer0_outputs(7637) <= inputs(125);
    layer0_outputs(7638) <= not((inputs(90)) or (inputs(12)));
    layer0_outputs(7639) <= not(inputs(115));
    layer0_outputs(7640) <= not((inputs(53)) or (inputs(208)));
    layer0_outputs(7641) <= not(inputs(77));
    layer0_outputs(7642) <= '0';
    layer0_outputs(7643) <= not(inputs(135)) or (inputs(21));
    layer0_outputs(7644) <= not(inputs(246));
    layer0_outputs(7645) <= not(inputs(236)) or (inputs(138));
    layer0_outputs(7646) <= not((inputs(148)) or (inputs(237)));
    layer0_outputs(7647) <= (inputs(25)) or (inputs(129));
    layer0_outputs(7648) <= not(inputs(13)) or (inputs(168));
    layer0_outputs(7649) <= (inputs(88)) and not (inputs(74));
    layer0_outputs(7650) <= (inputs(69)) or (inputs(171));
    layer0_outputs(7651) <= not((inputs(111)) or (inputs(224)));
    layer0_outputs(7652) <= (inputs(22)) or (inputs(124));
    layer0_outputs(7653) <= (inputs(16)) and not (inputs(94));
    layer0_outputs(7654) <= inputs(185);
    layer0_outputs(7655) <= not(inputs(234));
    layer0_outputs(7656) <= not((inputs(254)) xor (inputs(220)));
    layer0_outputs(7657) <= (inputs(19)) and not (inputs(124));
    layer0_outputs(7658) <= (inputs(234)) and not (inputs(62));
    layer0_outputs(7659) <= '1';
    layer0_outputs(7660) <= (inputs(247)) or (inputs(200));
    layer0_outputs(7661) <= not(inputs(100));
    layer0_outputs(7662) <= (inputs(213)) xor (inputs(179));
    layer0_outputs(7663) <= not(inputs(114));
    layer0_outputs(7664) <= not((inputs(19)) and (inputs(45)));
    layer0_outputs(7665) <= not(inputs(253));
    layer0_outputs(7666) <= not(inputs(61));
    layer0_outputs(7667) <= not(inputs(86));
    layer0_outputs(7668) <= (inputs(166)) or (inputs(193));
    layer0_outputs(7669) <= not((inputs(247)) or (inputs(87)));
    layer0_outputs(7670) <= inputs(170);
    layer0_outputs(7671) <= (inputs(25)) and not (inputs(181));
    layer0_outputs(7672) <= not(inputs(206));
    layer0_outputs(7673) <= inputs(211);
    layer0_outputs(7674) <= (inputs(58)) and not (inputs(171));
    layer0_outputs(7675) <= inputs(182);
    layer0_outputs(7676) <= '0';
    layer0_outputs(7677) <= not(inputs(116)) or (inputs(24));
    layer0_outputs(7678) <= (inputs(173)) and not (inputs(144));
    layer0_outputs(7679) <= not(inputs(99));
    layer1_outputs(0) <= not(layer0_outputs(4236));
    layer1_outputs(1) <= not(layer0_outputs(5512)) or (layer0_outputs(1906));
    layer1_outputs(2) <= '0';
    layer1_outputs(3) <= not((layer0_outputs(3167)) and (layer0_outputs(458)));
    layer1_outputs(4) <= '0';
    layer1_outputs(5) <= (layer0_outputs(5378)) and (layer0_outputs(5663));
    layer1_outputs(6) <= '0';
    layer1_outputs(7) <= layer0_outputs(5525);
    layer1_outputs(8) <= not(layer0_outputs(7081));
    layer1_outputs(9) <= not(layer0_outputs(5668)) or (layer0_outputs(5803));
    layer1_outputs(10) <= layer0_outputs(4703);
    layer1_outputs(11) <= not((layer0_outputs(1071)) xor (layer0_outputs(4346)));
    layer1_outputs(12) <= not(layer0_outputs(6347)) or (layer0_outputs(1813));
    layer1_outputs(13) <= not((layer0_outputs(3926)) and (layer0_outputs(3983)));
    layer1_outputs(14) <= layer0_outputs(2293);
    layer1_outputs(15) <= not(layer0_outputs(6353)) or (layer0_outputs(2404));
    layer1_outputs(16) <= not(layer0_outputs(7076));
    layer1_outputs(17) <= (layer0_outputs(1660)) and (layer0_outputs(165));
    layer1_outputs(18) <= not((layer0_outputs(2934)) or (layer0_outputs(7660)));
    layer1_outputs(19) <= (layer0_outputs(5889)) and not (layer0_outputs(2947));
    layer1_outputs(20) <= layer0_outputs(6504);
    layer1_outputs(21) <= (layer0_outputs(278)) or (layer0_outputs(5743));
    layer1_outputs(22) <= '1';
    layer1_outputs(23) <= layer0_outputs(3128);
    layer1_outputs(24) <= (layer0_outputs(3707)) and not (layer0_outputs(339));
    layer1_outputs(25) <= not(layer0_outputs(5908));
    layer1_outputs(26) <= not(layer0_outputs(1439)) or (layer0_outputs(6954));
    layer1_outputs(27) <= (layer0_outputs(5955)) or (layer0_outputs(5541));
    layer1_outputs(28) <= not(layer0_outputs(2068)) or (layer0_outputs(1051));
    layer1_outputs(29) <= (layer0_outputs(2366)) and (layer0_outputs(2704));
    layer1_outputs(30) <= (layer0_outputs(553)) and (layer0_outputs(4322));
    layer1_outputs(31) <= '1';
    layer1_outputs(32) <= '0';
    layer1_outputs(33) <= not((layer0_outputs(5440)) xor (layer0_outputs(7163)));
    layer1_outputs(34) <= not((layer0_outputs(4181)) or (layer0_outputs(2280)));
    layer1_outputs(35) <= not(layer0_outputs(4907));
    layer1_outputs(36) <= '1';
    layer1_outputs(37) <= '0';
    layer1_outputs(38) <= layer0_outputs(5216);
    layer1_outputs(39) <= '1';
    layer1_outputs(40) <= '1';
    layer1_outputs(41) <= not(layer0_outputs(7278));
    layer1_outputs(42) <= not(layer0_outputs(7605)) or (layer0_outputs(6313));
    layer1_outputs(43) <= '0';
    layer1_outputs(44) <= '0';
    layer1_outputs(45) <= not(layer0_outputs(3845)) or (layer0_outputs(2441));
    layer1_outputs(46) <= (layer0_outputs(7456)) and (layer0_outputs(5961));
    layer1_outputs(47) <= not((layer0_outputs(2254)) and (layer0_outputs(7238)));
    layer1_outputs(48) <= (layer0_outputs(3797)) and not (layer0_outputs(6433));
    layer1_outputs(49) <= not(layer0_outputs(1081));
    layer1_outputs(50) <= layer0_outputs(5298);
    layer1_outputs(51) <= layer0_outputs(4444);
    layer1_outputs(52) <= '0';
    layer1_outputs(53) <= not((layer0_outputs(918)) or (layer0_outputs(2553)));
    layer1_outputs(54) <= layer0_outputs(3714);
    layer1_outputs(55) <= not(layer0_outputs(537));
    layer1_outputs(56) <= not(layer0_outputs(2989));
    layer1_outputs(57) <= not(layer0_outputs(3217));
    layer1_outputs(58) <= not(layer0_outputs(2779));
    layer1_outputs(59) <= (layer0_outputs(5153)) or (layer0_outputs(7453));
    layer1_outputs(60) <= (layer0_outputs(5134)) and not (layer0_outputs(1717));
    layer1_outputs(61) <= not(layer0_outputs(3326)) or (layer0_outputs(7008));
    layer1_outputs(62) <= (layer0_outputs(4692)) and not (layer0_outputs(6868));
    layer1_outputs(63) <= not(layer0_outputs(3669)) or (layer0_outputs(2727));
    layer1_outputs(64) <= (layer0_outputs(1541)) and (layer0_outputs(4410));
    layer1_outputs(65) <= not((layer0_outputs(5860)) or (layer0_outputs(5919)));
    layer1_outputs(66) <= not((layer0_outputs(5190)) and (layer0_outputs(3486)));
    layer1_outputs(67) <= '0';
    layer1_outputs(68) <= not(layer0_outputs(290));
    layer1_outputs(69) <= '0';
    layer1_outputs(70) <= (layer0_outputs(7328)) or (layer0_outputs(7578));
    layer1_outputs(71) <= not(layer0_outputs(4831));
    layer1_outputs(72) <= not(layer0_outputs(5850));
    layer1_outputs(73) <= (layer0_outputs(5491)) and not (layer0_outputs(5821));
    layer1_outputs(74) <= '1';
    layer1_outputs(75) <= (layer0_outputs(3391)) xor (layer0_outputs(2737));
    layer1_outputs(76) <= layer0_outputs(399);
    layer1_outputs(77) <= (layer0_outputs(4074)) and not (layer0_outputs(6610));
    layer1_outputs(78) <= not((layer0_outputs(4600)) and (layer0_outputs(706)));
    layer1_outputs(79) <= not(layer0_outputs(2026)) or (layer0_outputs(4782));
    layer1_outputs(80) <= not((layer0_outputs(6036)) and (layer0_outputs(2757)));
    layer1_outputs(81) <= not(layer0_outputs(2376)) or (layer0_outputs(6620));
    layer1_outputs(82) <= not((layer0_outputs(927)) and (layer0_outputs(6793)));
    layer1_outputs(83) <= (layer0_outputs(5599)) and (layer0_outputs(5841));
    layer1_outputs(84) <= not(layer0_outputs(3791));
    layer1_outputs(85) <= not(layer0_outputs(5132)) or (layer0_outputs(3972));
    layer1_outputs(86) <= not((layer0_outputs(1803)) xor (layer0_outputs(5517)));
    layer1_outputs(87) <= layer0_outputs(7463);
    layer1_outputs(88) <= (layer0_outputs(571)) and (layer0_outputs(3532));
    layer1_outputs(89) <= not(layer0_outputs(2840));
    layer1_outputs(90) <= not(layer0_outputs(7158)) or (layer0_outputs(1334));
    layer1_outputs(91) <= not(layer0_outputs(1192));
    layer1_outputs(92) <= layer0_outputs(5822);
    layer1_outputs(93) <= layer0_outputs(4942);
    layer1_outputs(94) <= not(layer0_outputs(544));
    layer1_outputs(95) <= '0';
    layer1_outputs(96) <= not(layer0_outputs(6155)) or (layer0_outputs(273));
    layer1_outputs(97) <= not((layer0_outputs(6278)) or (layer0_outputs(3860)));
    layer1_outputs(98) <= not(layer0_outputs(6282)) or (layer0_outputs(6482));
    layer1_outputs(99) <= '1';
    layer1_outputs(100) <= '0';
    layer1_outputs(101) <= not(layer0_outputs(3964)) or (layer0_outputs(3016));
    layer1_outputs(102) <= (layer0_outputs(5553)) or (layer0_outputs(3106));
    layer1_outputs(103) <= not((layer0_outputs(7411)) and (layer0_outputs(3656)));
    layer1_outputs(104) <= layer0_outputs(505);
    layer1_outputs(105) <= not((layer0_outputs(1844)) and (layer0_outputs(882)));
    layer1_outputs(106) <= '1';
    layer1_outputs(107) <= (layer0_outputs(2420)) xor (layer0_outputs(1518));
    layer1_outputs(108) <= layer0_outputs(4280);
    layer1_outputs(109) <= layer0_outputs(1835);
    layer1_outputs(110) <= (layer0_outputs(4889)) and (layer0_outputs(4392));
    layer1_outputs(111) <= not((layer0_outputs(1879)) or (layer0_outputs(2918)));
    layer1_outputs(112) <= not(layer0_outputs(3110));
    layer1_outputs(113) <= (layer0_outputs(4497)) and (layer0_outputs(6447));
    layer1_outputs(114) <= '0';
    layer1_outputs(115) <= not(layer0_outputs(762));
    layer1_outputs(116) <= (layer0_outputs(1972)) or (layer0_outputs(4283));
    layer1_outputs(117) <= layer0_outputs(2961);
    layer1_outputs(118) <= (layer0_outputs(3713)) and not (layer0_outputs(1882));
    layer1_outputs(119) <= (layer0_outputs(177)) and not (layer0_outputs(5387));
    layer1_outputs(120) <= (layer0_outputs(3790)) or (layer0_outputs(1101));
    layer1_outputs(121) <= not(layer0_outputs(2629)) or (layer0_outputs(619));
    layer1_outputs(122) <= not(layer0_outputs(5519)) or (layer0_outputs(3098));
    layer1_outputs(123) <= (layer0_outputs(414)) and not (layer0_outputs(6961));
    layer1_outputs(124) <= (layer0_outputs(474)) and not (layer0_outputs(5807));
    layer1_outputs(125) <= '1';
    layer1_outputs(126) <= '0';
    layer1_outputs(127) <= not(layer0_outputs(3044));
    layer1_outputs(128) <= not(layer0_outputs(6746)) or (layer0_outputs(1510));
    layer1_outputs(129) <= layer0_outputs(5951);
    layer1_outputs(130) <= not(layer0_outputs(1517));
    layer1_outputs(131) <= (layer0_outputs(567)) or (layer0_outputs(3202));
    layer1_outputs(132) <= '0';
    layer1_outputs(133) <= (layer0_outputs(7487)) and not (layer0_outputs(526));
    layer1_outputs(134) <= (layer0_outputs(5049)) or (layer0_outputs(24));
    layer1_outputs(135) <= not(layer0_outputs(710));
    layer1_outputs(136) <= not(layer0_outputs(6639)) or (layer0_outputs(6937));
    layer1_outputs(137) <= (layer0_outputs(1777)) and not (layer0_outputs(1679));
    layer1_outputs(138) <= '1';
    layer1_outputs(139) <= not(layer0_outputs(5408));
    layer1_outputs(140) <= not((layer0_outputs(5894)) or (layer0_outputs(3772)));
    layer1_outputs(141) <= (layer0_outputs(3444)) and (layer0_outputs(5870));
    layer1_outputs(142) <= not(layer0_outputs(6130));
    layer1_outputs(143) <= (layer0_outputs(2425)) and not (layer0_outputs(693));
    layer1_outputs(144) <= not(layer0_outputs(1665));
    layer1_outputs(145) <= '1';
    layer1_outputs(146) <= not((layer0_outputs(6618)) and (layer0_outputs(5985)));
    layer1_outputs(147) <= not(layer0_outputs(4984)) or (layer0_outputs(6959));
    layer1_outputs(148) <= '0';
    layer1_outputs(149) <= not((layer0_outputs(2126)) and (layer0_outputs(7327)));
    layer1_outputs(150) <= not(layer0_outputs(958));
    layer1_outputs(151) <= (layer0_outputs(5603)) and not (layer0_outputs(812));
    layer1_outputs(152) <= '1';
    layer1_outputs(153) <= '1';
    layer1_outputs(154) <= layer0_outputs(4273);
    layer1_outputs(155) <= (layer0_outputs(500)) and not (layer0_outputs(7192));
    layer1_outputs(156) <= (layer0_outputs(2065)) and (layer0_outputs(395));
    layer1_outputs(157) <= '1';
    layer1_outputs(158) <= layer0_outputs(5551);
    layer1_outputs(159) <= not(layer0_outputs(3494));
    layer1_outputs(160) <= not((layer0_outputs(111)) or (layer0_outputs(4349)));
    layer1_outputs(161) <= layer0_outputs(5899);
    layer1_outputs(162) <= not((layer0_outputs(4168)) or (layer0_outputs(6531)));
    layer1_outputs(163) <= not(layer0_outputs(5541));
    layer1_outputs(164) <= (layer0_outputs(489)) or (layer0_outputs(6650));
    layer1_outputs(165) <= (layer0_outputs(2540)) and not (layer0_outputs(2916));
    layer1_outputs(166) <= '1';
    layer1_outputs(167) <= (layer0_outputs(3824)) and not (layer0_outputs(6713));
    layer1_outputs(168) <= layer0_outputs(7602);
    layer1_outputs(169) <= not(layer0_outputs(5574)) or (layer0_outputs(6689));
    layer1_outputs(170) <= not(layer0_outputs(6345)) or (layer0_outputs(5572));
    layer1_outputs(171) <= (layer0_outputs(3715)) and not (layer0_outputs(7096));
    layer1_outputs(172) <= (layer0_outputs(444)) or (layer0_outputs(6446));
    layer1_outputs(173) <= (layer0_outputs(2009)) and (layer0_outputs(6250));
    layer1_outputs(174) <= not((layer0_outputs(418)) or (layer0_outputs(5718)));
    layer1_outputs(175) <= layer0_outputs(4518);
    layer1_outputs(176) <= not(layer0_outputs(6111)) or (layer0_outputs(1242));
    layer1_outputs(177) <= not(layer0_outputs(2673));
    layer1_outputs(178) <= not(layer0_outputs(1364));
    layer1_outputs(179) <= (layer0_outputs(578)) and (layer0_outputs(3866));
    layer1_outputs(180) <= not(layer0_outputs(3426));
    layer1_outputs(181) <= not(layer0_outputs(2813));
    layer1_outputs(182) <= layer0_outputs(6851);
    layer1_outputs(183) <= not((layer0_outputs(2152)) and (layer0_outputs(2208)));
    layer1_outputs(184) <= (layer0_outputs(2222)) and not (layer0_outputs(2733));
    layer1_outputs(185) <= layer0_outputs(5115);
    layer1_outputs(186) <= not(layer0_outputs(2709));
    layer1_outputs(187) <= (layer0_outputs(1482)) and not (layer0_outputs(1538));
    layer1_outputs(188) <= not(layer0_outputs(1891)) or (layer0_outputs(132));
    layer1_outputs(189) <= '1';
    layer1_outputs(190) <= not((layer0_outputs(600)) and (layer0_outputs(3590)));
    layer1_outputs(191) <= '0';
    layer1_outputs(192) <= layer0_outputs(7371);
    layer1_outputs(193) <= not((layer0_outputs(1201)) or (layer0_outputs(7280)));
    layer1_outputs(194) <= not((layer0_outputs(2784)) and (layer0_outputs(1393)));
    layer1_outputs(195) <= not(layer0_outputs(981)) or (layer0_outputs(1341));
    layer1_outputs(196) <= layer0_outputs(3013);
    layer1_outputs(197) <= not(layer0_outputs(3982));
    layer1_outputs(198) <= layer0_outputs(5453);
    layer1_outputs(199) <= not(layer0_outputs(3038));
    layer1_outputs(200) <= (layer0_outputs(763)) and (layer0_outputs(1755));
    layer1_outputs(201) <= '0';
    layer1_outputs(202) <= not(layer0_outputs(4096));
    layer1_outputs(203) <= not((layer0_outputs(840)) or (layer0_outputs(1574)));
    layer1_outputs(204) <= not((layer0_outputs(1415)) and (layer0_outputs(1566)));
    layer1_outputs(205) <= (layer0_outputs(944)) and not (layer0_outputs(5354));
    layer1_outputs(206) <= '0';
    layer1_outputs(207) <= not(layer0_outputs(6270));
    layer1_outputs(208) <= (layer0_outputs(4247)) and not (layer0_outputs(7628));
    layer1_outputs(209) <= not(layer0_outputs(6972));
    layer1_outputs(210) <= (layer0_outputs(5029)) xor (layer0_outputs(3057));
    layer1_outputs(211) <= not(layer0_outputs(6892)) or (layer0_outputs(2800));
    layer1_outputs(212) <= '1';
    layer1_outputs(213) <= not(layer0_outputs(7501));
    layer1_outputs(214) <= '0';
    layer1_outputs(215) <= layer0_outputs(7104);
    layer1_outputs(216) <= not(layer0_outputs(6205));
    layer1_outputs(217) <= not(layer0_outputs(5676));
    layer1_outputs(218) <= '0';
    layer1_outputs(219) <= not((layer0_outputs(6246)) or (layer0_outputs(2036)));
    layer1_outputs(220) <= '0';
    layer1_outputs(221) <= not((layer0_outputs(2516)) or (layer0_outputs(4788)));
    layer1_outputs(222) <= not(layer0_outputs(6285));
    layer1_outputs(223) <= (layer0_outputs(5074)) or (layer0_outputs(1487));
    layer1_outputs(224) <= not((layer0_outputs(1634)) and (layer0_outputs(6179)));
    layer1_outputs(225) <= (layer0_outputs(2095)) or (layer0_outputs(3576));
    layer1_outputs(226) <= '1';
    layer1_outputs(227) <= layer0_outputs(70);
    layer1_outputs(228) <= not(layer0_outputs(4894)) or (layer0_outputs(5504));
    layer1_outputs(229) <= '0';
    layer1_outputs(230) <= not(layer0_outputs(6206));
    layer1_outputs(231) <= not(layer0_outputs(1595)) or (layer0_outputs(5212));
    layer1_outputs(232) <= not((layer0_outputs(3642)) and (layer0_outputs(396)));
    layer1_outputs(233) <= (layer0_outputs(2522)) and not (layer0_outputs(3550));
    layer1_outputs(234) <= layer0_outputs(7591);
    layer1_outputs(235) <= (layer0_outputs(4663)) and (layer0_outputs(7614));
    layer1_outputs(236) <= '0';
    layer1_outputs(237) <= (layer0_outputs(4097)) and not (layer0_outputs(3953));
    layer1_outputs(238) <= '0';
    layer1_outputs(239) <= '0';
    layer1_outputs(240) <= not((layer0_outputs(3408)) xor (layer0_outputs(4727)));
    layer1_outputs(241) <= not((layer0_outputs(4573)) or (layer0_outputs(5584)));
    layer1_outputs(242) <= not(layer0_outputs(2509));
    layer1_outputs(243) <= (layer0_outputs(6168)) or (layer0_outputs(5636));
    layer1_outputs(244) <= not((layer0_outputs(5755)) and (layer0_outputs(1730)));
    layer1_outputs(245) <= (layer0_outputs(7431)) or (layer0_outputs(1576));
    layer1_outputs(246) <= '0';
    layer1_outputs(247) <= layer0_outputs(1007);
    layer1_outputs(248) <= not(layer0_outputs(7181)) or (layer0_outputs(4754));
    layer1_outputs(249) <= layer0_outputs(6542);
    layer1_outputs(250) <= not(layer0_outputs(4655));
    layer1_outputs(251) <= '1';
    layer1_outputs(252) <= (layer0_outputs(4738)) and not (layer0_outputs(4651));
    layer1_outputs(253) <= (layer0_outputs(1886)) and (layer0_outputs(6720));
    layer1_outputs(254) <= not((layer0_outputs(228)) or (layer0_outputs(7362)));
    layer1_outputs(255) <= not((layer0_outputs(4304)) or (layer0_outputs(6608)));
    layer1_outputs(256) <= '1';
    layer1_outputs(257) <= (layer0_outputs(6818)) or (layer0_outputs(31));
    layer1_outputs(258) <= not((layer0_outputs(6534)) or (layer0_outputs(2106)));
    layer1_outputs(259) <= (layer0_outputs(5577)) and not (layer0_outputs(7245));
    layer1_outputs(260) <= not(layer0_outputs(2964));
    layer1_outputs(261) <= (layer0_outputs(3538)) or (layer0_outputs(6003));
    layer1_outputs(262) <= not(layer0_outputs(1528));
    layer1_outputs(263) <= (layer0_outputs(6613)) and not (layer0_outputs(1726));
    layer1_outputs(264) <= (layer0_outputs(2547)) and not (layer0_outputs(3606));
    layer1_outputs(265) <= layer0_outputs(3923);
    layer1_outputs(266) <= not(layer0_outputs(6762));
    layer1_outputs(267) <= layer0_outputs(2240);
    layer1_outputs(268) <= (layer0_outputs(6856)) or (layer0_outputs(4195));
    layer1_outputs(269) <= not((layer0_outputs(5970)) and (layer0_outputs(984)));
    layer1_outputs(270) <= not((layer0_outputs(6203)) and (layer0_outputs(5356)));
    layer1_outputs(271) <= not(layer0_outputs(3733));
    layer1_outputs(272) <= not(layer0_outputs(3148));
    layer1_outputs(273) <= not((layer0_outputs(2483)) or (layer0_outputs(3145)));
    layer1_outputs(274) <= (layer0_outputs(1639)) and not (layer0_outputs(1246));
    layer1_outputs(275) <= layer0_outputs(991);
    layer1_outputs(276) <= '0';
    layer1_outputs(277) <= not((layer0_outputs(6743)) and (layer0_outputs(1392)));
    layer1_outputs(278) <= not((layer0_outputs(4412)) or (layer0_outputs(3182)));
    layer1_outputs(279) <= not(layer0_outputs(7114)) or (layer0_outputs(7514));
    layer1_outputs(280) <= not(layer0_outputs(4009));
    layer1_outputs(281) <= layer0_outputs(7293);
    layer1_outputs(282) <= (layer0_outputs(1323)) and not (layer0_outputs(595));
    layer1_outputs(283) <= not((layer0_outputs(4514)) xor (layer0_outputs(3285)));
    layer1_outputs(284) <= '1';
    layer1_outputs(285) <= (layer0_outputs(6440)) and not (layer0_outputs(2581));
    layer1_outputs(286) <= not(layer0_outputs(6277));
    layer1_outputs(287) <= not((layer0_outputs(3344)) and (layer0_outputs(7533)));
    layer1_outputs(288) <= (layer0_outputs(1298)) or (layer0_outputs(5911));
    layer1_outputs(289) <= (layer0_outputs(4521)) and not (layer0_outputs(1999));
    layer1_outputs(290) <= (layer0_outputs(2181)) and not (layer0_outputs(4301));
    layer1_outputs(291) <= (layer0_outputs(5374)) and not (layer0_outputs(293));
    layer1_outputs(292) <= not(layer0_outputs(1995)) or (layer0_outputs(2475));
    layer1_outputs(293) <= not(layer0_outputs(3089));
    layer1_outputs(294) <= not(layer0_outputs(3646)) or (layer0_outputs(3004));
    layer1_outputs(295) <= not(layer0_outputs(6522)) or (layer0_outputs(2334));
    layer1_outputs(296) <= not(layer0_outputs(2999));
    layer1_outputs(297) <= (layer0_outputs(1061)) or (layer0_outputs(1583));
    layer1_outputs(298) <= (layer0_outputs(3624)) and (layer0_outputs(1343));
    layer1_outputs(299) <= (layer0_outputs(1784)) or (layer0_outputs(4732));
    layer1_outputs(300) <= (layer0_outputs(5656)) and not (layer0_outputs(1715));
    layer1_outputs(301) <= (layer0_outputs(2563)) and (layer0_outputs(3855));
    layer1_outputs(302) <= (layer0_outputs(5835)) and (layer0_outputs(7544));
    layer1_outputs(303) <= not(layer0_outputs(1007));
    layer1_outputs(304) <= '0';
    layer1_outputs(305) <= not((layer0_outputs(6049)) or (layer0_outputs(3209)));
    layer1_outputs(306) <= not(layer0_outputs(7564));
    layer1_outputs(307) <= (layer0_outputs(6631)) and not (layer0_outputs(1728));
    layer1_outputs(308) <= not((layer0_outputs(2086)) and (layer0_outputs(3994)));
    layer1_outputs(309) <= layer0_outputs(6978);
    layer1_outputs(310) <= layer0_outputs(7315);
    layer1_outputs(311) <= (layer0_outputs(4577)) and (layer0_outputs(2267));
    layer1_outputs(312) <= not((layer0_outputs(3959)) or (layer0_outputs(6497)));
    layer1_outputs(313) <= (layer0_outputs(4706)) or (layer0_outputs(6065));
    layer1_outputs(314) <= (layer0_outputs(146)) or (layer0_outputs(358));
    layer1_outputs(315) <= layer0_outputs(1183);
    layer1_outputs(316) <= (layer0_outputs(6590)) or (layer0_outputs(915));
    layer1_outputs(317) <= (layer0_outputs(7248)) and not (layer0_outputs(2370));
    layer1_outputs(318) <= (layer0_outputs(4024)) and not (layer0_outputs(3385));
    layer1_outputs(319) <= layer0_outputs(1699);
    layer1_outputs(320) <= not(layer0_outputs(3861));
    layer1_outputs(321) <= '0';
    layer1_outputs(322) <= (layer0_outputs(3784)) and (layer0_outputs(3919));
    layer1_outputs(323) <= not(layer0_outputs(6922)) or (layer0_outputs(4468));
    layer1_outputs(324) <= (layer0_outputs(6863)) and not (layer0_outputs(6363));
    layer1_outputs(325) <= layer0_outputs(5907);
    layer1_outputs(326) <= not(layer0_outputs(1059)) or (layer0_outputs(5926));
    layer1_outputs(327) <= not(layer0_outputs(4924)) or (layer0_outputs(5443));
    layer1_outputs(328) <= '0';
    layer1_outputs(329) <= '1';
    layer1_outputs(330) <= (layer0_outputs(87)) or (layer0_outputs(6820));
    layer1_outputs(331) <= '0';
    layer1_outputs(332) <= not(layer0_outputs(3024)) or (layer0_outputs(2434));
    layer1_outputs(333) <= not((layer0_outputs(5392)) xor (layer0_outputs(2134)));
    layer1_outputs(334) <= not(layer0_outputs(544)) or (layer0_outputs(1622));
    layer1_outputs(335) <= layer0_outputs(5222);
    layer1_outputs(336) <= not(layer0_outputs(5259));
    layer1_outputs(337) <= (layer0_outputs(180)) and not (layer0_outputs(6198));
    layer1_outputs(338) <= not(layer0_outputs(4280));
    layer1_outputs(339) <= '1';
    layer1_outputs(340) <= layer0_outputs(4951);
    layer1_outputs(341) <= (layer0_outputs(3771)) and not (layer0_outputs(7558));
    layer1_outputs(342) <= not(layer0_outputs(2071));
    layer1_outputs(343) <= (layer0_outputs(6896)) or (layer0_outputs(2514));
    layer1_outputs(344) <= not(layer0_outputs(3681)) or (layer0_outputs(1799));
    layer1_outputs(345) <= not(layer0_outputs(2549)) or (layer0_outputs(564));
    layer1_outputs(346) <= not(layer0_outputs(1219)) or (layer0_outputs(2222));
    layer1_outputs(347) <= not((layer0_outputs(3880)) or (layer0_outputs(5823)));
    layer1_outputs(348) <= (layer0_outputs(742)) and not (layer0_outputs(5295));
    layer1_outputs(349) <= '1';
    layer1_outputs(350) <= '0';
    layer1_outputs(351) <= not(layer0_outputs(7110));
    layer1_outputs(352) <= not((layer0_outputs(1956)) or (layer0_outputs(4534)));
    layer1_outputs(353) <= '1';
    layer1_outputs(354) <= (layer0_outputs(6513)) and (layer0_outputs(2101));
    layer1_outputs(355) <= not(layer0_outputs(6815));
    layer1_outputs(356) <= not(layer0_outputs(3173)) or (layer0_outputs(7010));
    layer1_outputs(357) <= not((layer0_outputs(5882)) and (layer0_outputs(3097)));
    layer1_outputs(358) <= not(layer0_outputs(3940)) or (layer0_outputs(4303));
    layer1_outputs(359) <= not(layer0_outputs(852)) or (layer0_outputs(7350));
    layer1_outputs(360) <= '1';
    layer1_outputs(361) <= (layer0_outputs(7471)) xor (layer0_outputs(2671));
    layer1_outputs(362) <= not(layer0_outputs(6112)) or (layer0_outputs(3498));
    layer1_outputs(363) <= not((layer0_outputs(931)) and (layer0_outputs(6068)));
    layer1_outputs(364) <= not(layer0_outputs(3059));
    layer1_outputs(365) <= not(layer0_outputs(3571));
    layer1_outputs(366) <= not(layer0_outputs(3306));
    layer1_outputs(367) <= '0';
    layer1_outputs(368) <= '0';
    layer1_outputs(369) <= not(layer0_outputs(5565)) or (layer0_outputs(2843));
    layer1_outputs(370) <= not(layer0_outputs(6421));
    layer1_outputs(371) <= not(layer0_outputs(5663)) or (layer0_outputs(7226));
    layer1_outputs(372) <= (layer0_outputs(1680)) and not (layer0_outputs(939));
    layer1_outputs(373) <= '1';
    layer1_outputs(374) <= not(layer0_outputs(1565)) or (layer0_outputs(3339));
    layer1_outputs(375) <= '1';
    layer1_outputs(376) <= '1';
    layer1_outputs(377) <= not(layer0_outputs(2079));
    layer1_outputs(378) <= (layer0_outputs(5713)) and not (layer0_outputs(3932));
    layer1_outputs(379) <= not((layer0_outputs(4140)) and (layer0_outputs(834)));
    layer1_outputs(380) <= layer0_outputs(5056);
    layer1_outputs(381) <= not(layer0_outputs(4975));
    layer1_outputs(382) <= layer0_outputs(5734);
    layer1_outputs(383) <= (layer0_outputs(6147)) and (layer0_outputs(3875));
    layer1_outputs(384) <= not((layer0_outputs(1126)) and (layer0_outputs(676)));
    layer1_outputs(385) <= (layer0_outputs(7321)) and not (layer0_outputs(2588));
    layer1_outputs(386) <= not(layer0_outputs(323));
    layer1_outputs(387) <= not(layer0_outputs(3155));
    layer1_outputs(388) <= not((layer0_outputs(2100)) and (layer0_outputs(2072)));
    layer1_outputs(389) <= not(layer0_outputs(6361));
    layer1_outputs(390) <= not((layer0_outputs(6312)) and (layer0_outputs(5873)));
    layer1_outputs(391) <= (layer0_outputs(1672)) and not (layer0_outputs(3353));
    layer1_outputs(392) <= (layer0_outputs(5501)) and not (layer0_outputs(1807));
    layer1_outputs(393) <= not((layer0_outputs(754)) xor (layer0_outputs(7370)));
    layer1_outputs(394) <= layer0_outputs(2304);
    layer1_outputs(395) <= (layer0_outputs(2074)) and (layer0_outputs(5717));
    layer1_outputs(396) <= layer0_outputs(2603);
    layer1_outputs(397) <= not(layer0_outputs(6050));
    layer1_outputs(398) <= (layer0_outputs(60)) or (layer0_outputs(1483));
    layer1_outputs(399) <= not(layer0_outputs(6960)) or (layer0_outputs(4127));
    layer1_outputs(400) <= not(layer0_outputs(712));
    layer1_outputs(401) <= not(layer0_outputs(1707));
    layer1_outputs(402) <= not(layer0_outputs(1127)) or (layer0_outputs(3096));
    layer1_outputs(403) <= (layer0_outputs(6169)) and not (layer0_outputs(4066));
    layer1_outputs(404) <= layer0_outputs(7551);
    layer1_outputs(405) <= '0';
    layer1_outputs(406) <= (layer0_outputs(2096)) or (layer0_outputs(4387));
    layer1_outputs(407) <= '0';
    layer1_outputs(408) <= not(layer0_outputs(6437));
    layer1_outputs(409) <= not(layer0_outputs(2243));
    layer1_outputs(410) <= '0';
    layer1_outputs(411) <= not(layer0_outputs(858)) or (layer0_outputs(1811));
    layer1_outputs(412) <= not(layer0_outputs(6553)) or (layer0_outputs(501));
    layer1_outputs(413) <= layer0_outputs(4167);
    layer1_outputs(414) <= (layer0_outputs(6534)) and not (layer0_outputs(3816));
    layer1_outputs(415) <= not(layer0_outputs(3390)) or (layer0_outputs(208));
    layer1_outputs(416) <= '1';
    layer1_outputs(417) <= not(layer0_outputs(2898));
    layer1_outputs(418) <= not(layer0_outputs(777));
    layer1_outputs(419) <= layer0_outputs(5964);
    layer1_outputs(420) <= not(layer0_outputs(7337));
    layer1_outputs(421) <= (layer0_outputs(7013)) and (layer0_outputs(621));
    layer1_outputs(422) <= not(layer0_outputs(5798)) or (layer0_outputs(5199));
    layer1_outputs(423) <= not(layer0_outputs(440)) or (layer0_outputs(4617));
    layer1_outputs(424) <= (layer0_outputs(3065)) and (layer0_outputs(2376));
    layer1_outputs(425) <= (layer0_outputs(3283)) and (layer0_outputs(3392));
    layer1_outputs(426) <= not(layer0_outputs(3844)) or (layer0_outputs(2061));
    layer1_outputs(427) <= not((layer0_outputs(2840)) and (layer0_outputs(1535)));
    layer1_outputs(428) <= not(layer0_outputs(1118));
    layer1_outputs(429) <= '0';
    layer1_outputs(430) <= (layer0_outputs(6590)) and not (layer0_outputs(5425));
    layer1_outputs(431) <= (layer0_outputs(3907)) xor (layer0_outputs(3910));
    layer1_outputs(432) <= layer0_outputs(5227);
    layer1_outputs(433) <= '1';
    layer1_outputs(434) <= (layer0_outputs(4814)) and not (layer0_outputs(6414));
    layer1_outputs(435) <= (layer0_outputs(1516)) and (layer0_outputs(333));
    layer1_outputs(436) <= not(layer0_outputs(3548));
    layer1_outputs(437) <= not((layer0_outputs(4520)) or (layer0_outputs(3089)));
    layer1_outputs(438) <= not((layer0_outputs(4911)) or (layer0_outputs(4512)));
    layer1_outputs(439) <= not(layer0_outputs(4446));
    layer1_outputs(440) <= not(layer0_outputs(456));
    layer1_outputs(441) <= '1';
    layer1_outputs(442) <= layer0_outputs(2184);
    layer1_outputs(443) <= not((layer0_outputs(1890)) or (layer0_outputs(367)));
    layer1_outputs(444) <= '0';
    layer1_outputs(445) <= not(layer0_outputs(4851));
    layer1_outputs(446) <= not((layer0_outputs(3472)) or (layer0_outputs(4506)));
    layer1_outputs(447) <= layer0_outputs(233);
    layer1_outputs(448) <= (layer0_outputs(183)) and not (layer0_outputs(6509));
    layer1_outputs(449) <= (layer0_outputs(2846)) and not (layer0_outputs(2646));
    layer1_outputs(450) <= not(layer0_outputs(2938)) or (layer0_outputs(7366));
    layer1_outputs(451) <= '1';
    layer1_outputs(452) <= '0';
    layer1_outputs(453) <= not(layer0_outputs(5076));
    layer1_outputs(454) <= layer0_outputs(4248);
    layer1_outputs(455) <= not(layer0_outputs(202));
    layer1_outputs(456) <= not(layer0_outputs(3417));
    layer1_outputs(457) <= layer0_outputs(1812);
    layer1_outputs(458) <= (layer0_outputs(7098)) and (layer0_outputs(952));
    layer1_outputs(459) <= not(layer0_outputs(1814));
    layer1_outputs(460) <= '0';
    layer1_outputs(461) <= not(layer0_outputs(4393));
    layer1_outputs(462) <= (layer0_outputs(7112)) and (layer0_outputs(6650));
    layer1_outputs(463) <= layer0_outputs(2708);
    layer1_outputs(464) <= not(layer0_outputs(3968));
    layer1_outputs(465) <= not((layer0_outputs(5393)) or (layer0_outputs(5339)));
    layer1_outputs(466) <= not(layer0_outputs(2090)) or (layer0_outputs(837));
    layer1_outputs(467) <= '1';
    layer1_outputs(468) <= not((layer0_outputs(4563)) or (layer0_outputs(6582)));
    layer1_outputs(469) <= not((layer0_outputs(5860)) and (layer0_outputs(2406)));
    layer1_outputs(470) <= layer0_outputs(2741);
    layer1_outputs(471) <= '1';
    layer1_outputs(472) <= (layer0_outputs(3262)) and not (layer0_outputs(5608));
    layer1_outputs(473) <= '1';
    layer1_outputs(474) <= not(layer0_outputs(7339));
    layer1_outputs(475) <= layer0_outputs(6835);
    layer1_outputs(476) <= not((layer0_outputs(1475)) xor (layer0_outputs(7256)));
    layer1_outputs(477) <= (layer0_outputs(2961)) and not (layer0_outputs(5527));
    layer1_outputs(478) <= '0';
    layer1_outputs(479) <= (layer0_outputs(3260)) and not (layer0_outputs(1069));
    layer1_outputs(480) <= (layer0_outputs(6570)) or (layer0_outputs(128));
    layer1_outputs(481) <= '1';
    layer1_outputs(482) <= (layer0_outputs(6760)) or (layer0_outputs(7531));
    layer1_outputs(483) <= not(layer0_outputs(6779)) or (layer0_outputs(406));
    layer1_outputs(484) <= (layer0_outputs(6579)) and not (layer0_outputs(889));
    layer1_outputs(485) <= not(layer0_outputs(3916));
    layer1_outputs(486) <= '1';
    layer1_outputs(487) <= not((layer0_outputs(6975)) or (layer0_outputs(3415)));
    layer1_outputs(488) <= (layer0_outputs(4162)) and (layer0_outputs(4002));
    layer1_outputs(489) <= not(layer0_outputs(62));
    layer1_outputs(490) <= not(layer0_outputs(1258)) or (layer0_outputs(3097));
    layer1_outputs(491) <= not((layer0_outputs(4599)) or (layer0_outputs(5899)));
    layer1_outputs(492) <= not(layer0_outputs(2905)) or (layer0_outputs(2260));
    layer1_outputs(493) <= (layer0_outputs(2443)) or (layer0_outputs(7358));
    layer1_outputs(494) <= layer0_outputs(2492);
    layer1_outputs(495) <= not(layer0_outputs(1652)) or (layer0_outputs(6387));
    layer1_outputs(496) <= '0';
    layer1_outputs(497) <= (layer0_outputs(5320)) and not (layer0_outputs(4763));
    layer1_outputs(498) <= (layer0_outputs(5519)) or (layer0_outputs(5034));
    layer1_outputs(499) <= (layer0_outputs(1925)) and not (layer0_outputs(1354));
    layer1_outputs(500) <= not(layer0_outputs(1178)) or (layer0_outputs(4937));
    layer1_outputs(501) <= (layer0_outputs(1845)) and not (layer0_outputs(152));
    layer1_outputs(502) <= not((layer0_outputs(972)) and (layer0_outputs(271)));
    layer1_outputs(503) <= not(layer0_outputs(2034)) or (layer0_outputs(7334));
    layer1_outputs(504) <= (layer0_outputs(2289)) and not (layer0_outputs(5813));
    layer1_outputs(505) <= '0';
    layer1_outputs(506) <= '1';
    layer1_outputs(507) <= (layer0_outputs(4479)) and (layer0_outputs(5277));
    layer1_outputs(508) <= (layer0_outputs(4587)) or (layer0_outputs(1607));
    layer1_outputs(509) <= '0';
    layer1_outputs(510) <= not(layer0_outputs(1407));
    layer1_outputs(511) <= not(layer0_outputs(2300));
    layer1_outputs(512) <= (layer0_outputs(741)) and not (layer0_outputs(961));
    layer1_outputs(513) <= not((layer0_outputs(4132)) and (layer0_outputs(4637)));
    layer1_outputs(514) <= (layer0_outputs(2946)) or (layer0_outputs(6800));
    layer1_outputs(515) <= (layer0_outputs(851)) and not (layer0_outputs(3031));
    layer1_outputs(516) <= '1';
    layer1_outputs(517) <= not(layer0_outputs(2607));
    layer1_outputs(518) <= not(layer0_outputs(3045)) or (layer0_outputs(2845));
    layer1_outputs(519) <= (layer0_outputs(804)) and (layer0_outputs(4790));
    layer1_outputs(520) <= not(layer0_outputs(4428)) or (layer0_outputs(6948));
    layer1_outputs(521) <= not((layer0_outputs(33)) and (layer0_outputs(3378)));
    layer1_outputs(522) <= not(layer0_outputs(2986));
    layer1_outputs(523) <= not((layer0_outputs(1496)) or (layer0_outputs(246)));
    layer1_outputs(524) <= not((layer0_outputs(3041)) or (layer0_outputs(4585)));
    layer1_outputs(525) <= (layer0_outputs(7263)) and not (layer0_outputs(1967));
    layer1_outputs(526) <= (layer0_outputs(7140)) and not (layer0_outputs(5259));
    layer1_outputs(527) <= not(layer0_outputs(3578)) or (layer0_outputs(344));
    layer1_outputs(528) <= not(layer0_outputs(3718));
    layer1_outputs(529) <= not(layer0_outputs(4797)) or (layer0_outputs(1397));
    layer1_outputs(530) <= not(layer0_outputs(4502)) or (layer0_outputs(6568));
    layer1_outputs(531) <= (layer0_outputs(6846)) and not (layer0_outputs(4416));
    layer1_outputs(532) <= not(layer0_outputs(3413));
    layer1_outputs(533) <= '0';
    layer1_outputs(534) <= (layer0_outputs(7048)) xor (layer0_outputs(2812));
    layer1_outputs(535) <= not(layer0_outputs(1611));
    layer1_outputs(536) <= '0';
    layer1_outputs(537) <= not(layer0_outputs(1692));
    layer1_outputs(538) <= (layer0_outputs(6116)) or (layer0_outputs(5994));
    layer1_outputs(539) <= layer0_outputs(279);
    layer1_outputs(540) <= (layer0_outputs(1820)) or (layer0_outputs(5294));
    layer1_outputs(541) <= layer0_outputs(5043);
    layer1_outputs(542) <= not(layer0_outputs(1464));
    layer1_outputs(543) <= '1';
    layer1_outputs(544) <= not(layer0_outputs(2492));
    layer1_outputs(545) <= not(layer0_outputs(3410));
    layer1_outputs(546) <= (layer0_outputs(2117)) xor (layer0_outputs(2715));
    layer1_outputs(547) <= not(layer0_outputs(5262)) or (layer0_outputs(5474));
    layer1_outputs(548) <= layer0_outputs(4462);
    layer1_outputs(549) <= not((layer0_outputs(7517)) and (layer0_outputs(2534)));
    layer1_outputs(550) <= '0';
    layer1_outputs(551) <= layer0_outputs(1347);
    layer1_outputs(552) <= not((layer0_outputs(690)) or (layer0_outputs(659)));
    layer1_outputs(553) <= '0';
    layer1_outputs(554) <= layer0_outputs(5670);
    layer1_outputs(555) <= not((layer0_outputs(5109)) or (layer0_outputs(3874)));
    layer1_outputs(556) <= (layer0_outputs(657)) and not (layer0_outputs(7406));
    layer1_outputs(557) <= not(layer0_outputs(142)) or (layer0_outputs(5762));
    layer1_outputs(558) <= not(layer0_outputs(2946));
    layer1_outputs(559) <= not((layer0_outputs(417)) or (layer0_outputs(4970)));
    layer1_outputs(560) <= layer0_outputs(3922);
    layer1_outputs(561) <= not(layer0_outputs(7332)) or (layer0_outputs(3768));
    layer1_outputs(562) <= not(layer0_outputs(131));
    layer1_outputs(563) <= (layer0_outputs(5558)) or (layer0_outputs(3832));
    layer1_outputs(564) <= (layer0_outputs(5613)) or (layer0_outputs(4650));
    layer1_outputs(565) <= not(layer0_outputs(1915));
    layer1_outputs(566) <= (layer0_outputs(6936)) and not (layer0_outputs(4730));
    layer1_outputs(567) <= (layer0_outputs(2121)) and not (layer0_outputs(4858));
    layer1_outputs(568) <= not(layer0_outputs(40));
    layer1_outputs(569) <= (layer0_outputs(523)) and (layer0_outputs(3124));
    layer1_outputs(570) <= '1';
    layer1_outputs(571) <= (layer0_outputs(2491)) xor (layer0_outputs(5405));
    layer1_outputs(572) <= not(layer0_outputs(5644));
    layer1_outputs(573) <= '0';
    layer1_outputs(574) <= (layer0_outputs(7321)) or (layer0_outputs(7150));
    layer1_outputs(575) <= layer0_outputs(647);
    layer1_outputs(576) <= layer0_outputs(7117);
    layer1_outputs(577) <= not(layer0_outputs(2860)) or (layer0_outputs(4967));
    layer1_outputs(578) <= not((layer0_outputs(7604)) xor (layer0_outputs(5283)));
    layer1_outputs(579) <= not((layer0_outputs(1312)) and (layer0_outputs(7524)));
    layer1_outputs(580) <= not(layer0_outputs(6634));
    layer1_outputs(581) <= not(layer0_outputs(2593)) or (layer0_outputs(2629));
    layer1_outputs(582) <= (layer0_outputs(4036)) and not (layer0_outputs(5393));
    layer1_outputs(583) <= not(layer0_outputs(5984));
    layer1_outputs(584) <= '0';
    layer1_outputs(585) <= (layer0_outputs(6925)) or (layer0_outputs(6773));
    layer1_outputs(586) <= not(layer0_outputs(421)) or (layer0_outputs(3725));
    layer1_outputs(587) <= (layer0_outputs(5277)) or (layer0_outputs(1256));
    layer1_outputs(588) <= layer0_outputs(3218);
    layer1_outputs(589) <= '0';
    layer1_outputs(590) <= (layer0_outputs(4687)) xor (layer0_outputs(5644));
    layer1_outputs(591) <= (layer0_outputs(7584)) or (layer0_outputs(3943));
    layer1_outputs(592) <= not((layer0_outputs(1121)) xor (layer0_outputs(1153)));
    layer1_outputs(593) <= not((layer0_outputs(6920)) xor (layer0_outputs(5764)));
    layer1_outputs(594) <= layer0_outputs(6982);
    layer1_outputs(595) <= (layer0_outputs(2416)) and not (layer0_outputs(5507));
    layer1_outputs(596) <= not((layer0_outputs(6520)) and (layer0_outputs(79)));
    layer1_outputs(597) <= '1';
    layer1_outputs(598) <= not(layer0_outputs(7633));
    layer1_outputs(599) <= not((layer0_outputs(4328)) or (layer0_outputs(796)));
    layer1_outputs(600) <= not(layer0_outputs(3063));
    layer1_outputs(601) <= not(layer0_outputs(290)) or (layer0_outputs(7599));
    layer1_outputs(602) <= '0';
    layer1_outputs(603) <= layer0_outputs(6251);
    layer1_outputs(604) <= layer0_outputs(6978);
    layer1_outputs(605) <= not(layer0_outputs(7317));
    layer1_outputs(606) <= not(layer0_outputs(1011)) or (layer0_outputs(1767));
    layer1_outputs(607) <= '1';
    layer1_outputs(608) <= not(layer0_outputs(5872)) or (layer0_outputs(5727));
    layer1_outputs(609) <= not(layer0_outputs(4629));
    layer1_outputs(610) <= layer0_outputs(3507);
    layer1_outputs(611) <= (layer0_outputs(7378)) and not (layer0_outputs(3941));
    layer1_outputs(612) <= not(layer0_outputs(1194));
    layer1_outputs(613) <= not(layer0_outputs(3583));
    layer1_outputs(614) <= layer0_outputs(6421);
    layer1_outputs(615) <= (layer0_outputs(1699)) xor (layer0_outputs(505));
    layer1_outputs(616) <= not((layer0_outputs(7354)) and (layer0_outputs(7194)));
    layer1_outputs(617) <= layer0_outputs(1764);
    layer1_outputs(618) <= layer0_outputs(3101);
    layer1_outputs(619) <= (layer0_outputs(4796)) and not (layer0_outputs(6488));
    layer1_outputs(620) <= not((layer0_outputs(6564)) and (layer0_outputs(3888)));
    layer1_outputs(621) <= not(layer0_outputs(7256)) or (layer0_outputs(5242));
    layer1_outputs(622) <= (layer0_outputs(6825)) and (layer0_outputs(7068));
    layer1_outputs(623) <= not((layer0_outputs(2027)) or (layer0_outputs(4835)));
    layer1_outputs(624) <= '0';
    layer1_outputs(625) <= (layer0_outputs(245)) and not (layer0_outputs(6242));
    layer1_outputs(626) <= '1';
    layer1_outputs(627) <= layer0_outputs(2035);
    layer1_outputs(628) <= '0';
    layer1_outputs(629) <= (layer0_outputs(5471)) and not (layer0_outputs(4166));
    layer1_outputs(630) <= layer0_outputs(1683);
    layer1_outputs(631) <= not(layer0_outputs(5606)) or (layer0_outputs(1146));
    layer1_outputs(632) <= not((layer0_outputs(1853)) or (layer0_outputs(6386)));
    layer1_outputs(633) <= not(layer0_outputs(5743));
    layer1_outputs(634) <= '1';
    layer1_outputs(635) <= '1';
    layer1_outputs(636) <= layer0_outputs(5543);
    layer1_outputs(637) <= (layer0_outputs(1134)) and not (layer0_outputs(5040));
    layer1_outputs(638) <= not(layer0_outputs(2982)) or (layer0_outputs(384));
    layer1_outputs(639) <= (layer0_outputs(1242)) and not (layer0_outputs(990));
    layer1_outputs(640) <= not((layer0_outputs(7579)) xor (layer0_outputs(2198)));
    layer1_outputs(641) <= (layer0_outputs(5360)) and (layer0_outputs(4617));
    layer1_outputs(642) <= '0';
    layer1_outputs(643) <= not((layer0_outputs(933)) xor (layer0_outputs(7348)));
    layer1_outputs(644) <= (layer0_outputs(3506)) and not (layer0_outputs(4783));
    layer1_outputs(645) <= not((layer0_outputs(195)) and (layer0_outputs(2391)));
    layer1_outputs(646) <= not(layer0_outputs(7564));
    layer1_outputs(647) <= not(layer0_outputs(7193)) or (layer0_outputs(7509));
    layer1_outputs(648) <= not(layer0_outputs(2853));
    layer1_outputs(649) <= '0';
    layer1_outputs(650) <= not((layer0_outputs(6833)) or (layer0_outputs(3431)));
    layer1_outputs(651) <= '0';
    layer1_outputs(652) <= not(layer0_outputs(1854));
    layer1_outputs(653) <= not(layer0_outputs(3429)) or (layer0_outputs(872));
    layer1_outputs(654) <= layer0_outputs(6271);
    layer1_outputs(655) <= not((layer0_outputs(6113)) and (layer0_outputs(4608)));
    layer1_outputs(656) <= not((layer0_outputs(4601)) or (layer0_outputs(2537)));
    layer1_outputs(657) <= (layer0_outputs(2144)) and (layer0_outputs(2525));
    layer1_outputs(658) <= layer0_outputs(6157);
    layer1_outputs(659) <= (layer0_outputs(1104)) and not (layer0_outputs(2808));
    layer1_outputs(660) <= '1';
    layer1_outputs(661) <= not(layer0_outputs(6369));
    layer1_outputs(662) <= not(layer0_outputs(5427)) or (layer0_outputs(2048));
    layer1_outputs(663) <= not((layer0_outputs(6326)) and (layer0_outputs(6556)));
    layer1_outputs(664) <= (layer0_outputs(3818)) and (layer0_outputs(3786));
    layer1_outputs(665) <= layer0_outputs(6511);
    layer1_outputs(666) <= not((layer0_outputs(1010)) or (layer0_outputs(1948)));
    layer1_outputs(667) <= layer0_outputs(5476);
    layer1_outputs(668) <= not((layer0_outputs(7084)) or (layer0_outputs(4442)));
    layer1_outputs(669) <= (layer0_outputs(4781)) and not (layer0_outputs(299));
    layer1_outputs(670) <= layer0_outputs(1753);
    layer1_outputs(671) <= not(layer0_outputs(1990));
    layer1_outputs(672) <= (layer0_outputs(2287)) and not (layer0_outputs(4644));
    layer1_outputs(673) <= (layer0_outputs(4789)) and not (layer0_outputs(7159));
    layer1_outputs(674) <= '1';
    layer1_outputs(675) <= layer0_outputs(5723);
    layer1_outputs(676) <= not(layer0_outputs(2854));
    layer1_outputs(677) <= (layer0_outputs(4717)) and not (layer0_outputs(6020));
    layer1_outputs(678) <= (layer0_outputs(4483)) and not (layer0_outputs(1646));
    layer1_outputs(679) <= '1';
    layer1_outputs(680) <= layer0_outputs(1014);
    layer1_outputs(681) <= (layer0_outputs(6791)) and not (layer0_outputs(1675));
    layer1_outputs(682) <= not(layer0_outputs(429)) or (layer0_outputs(3698));
    layer1_outputs(683) <= '1';
    layer1_outputs(684) <= not(layer0_outputs(3332));
    layer1_outputs(685) <= (layer0_outputs(6746)) or (layer0_outputs(3644));
    layer1_outputs(686) <= not(layer0_outputs(4448));
    layer1_outputs(687) <= layer0_outputs(1453);
    layer1_outputs(688) <= (layer0_outputs(4278)) and not (layer0_outputs(5032));
    layer1_outputs(689) <= (layer0_outputs(2211)) and (layer0_outputs(4809));
    layer1_outputs(690) <= not((layer0_outputs(7031)) and (layer0_outputs(4408)));
    layer1_outputs(691) <= not(layer0_outputs(6454)) or (layer0_outputs(2223));
    layer1_outputs(692) <= layer0_outputs(3313);
    layer1_outputs(693) <= (layer0_outputs(3573)) and not (layer0_outputs(7184));
    layer1_outputs(694) <= '1';
    layer1_outputs(695) <= not(layer0_outputs(5747)) or (layer0_outputs(4450));
    layer1_outputs(696) <= not(layer0_outputs(6094));
    layer1_outputs(697) <= not((layer0_outputs(4911)) and (layer0_outputs(6160)));
    layer1_outputs(698) <= layer0_outputs(970);
    layer1_outputs(699) <= not((layer0_outputs(4234)) and (layer0_outputs(2012)));
    layer1_outputs(700) <= not(layer0_outputs(3537)) or (layer0_outputs(7168));
    layer1_outputs(701) <= not(layer0_outputs(5483));
    layer1_outputs(702) <= layer0_outputs(7);
    layer1_outputs(703) <= not((layer0_outputs(635)) and (layer0_outputs(1616)));
    layer1_outputs(704) <= (layer0_outputs(4826)) and not (layer0_outputs(6046));
    layer1_outputs(705) <= not(layer0_outputs(6471));
    layer1_outputs(706) <= (layer0_outputs(4705)) xor (layer0_outputs(1572));
    layer1_outputs(707) <= not(layer0_outputs(3350));
    layer1_outputs(708) <= not(layer0_outputs(5368));
    layer1_outputs(709) <= (layer0_outputs(4513)) and (layer0_outputs(459));
    layer1_outputs(710) <= layer0_outputs(630);
    layer1_outputs(711) <= '1';
    layer1_outputs(712) <= not(layer0_outputs(3259));
    layer1_outputs(713) <= not(layer0_outputs(1289)) or (layer0_outputs(3523));
    layer1_outputs(714) <= layer0_outputs(2536);
    layer1_outputs(715) <= '0';
    layer1_outputs(716) <= not(layer0_outputs(3804));
    layer1_outputs(717) <= '1';
    layer1_outputs(718) <= '0';
    layer1_outputs(719) <= not(layer0_outputs(6008)) or (layer0_outputs(2697));
    layer1_outputs(720) <= (layer0_outputs(1465)) and (layer0_outputs(2019));
    layer1_outputs(721) <= (layer0_outputs(3312)) and not (layer0_outputs(7673));
    layer1_outputs(722) <= not(layer0_outputs(2642)) or (layer0_outputs(5704));
    layer1_outputs(723) <= (layer0_outputs(6631)) and not (layer0_outputs(5384));
    layer1_outputs(724) <= (layer0_outputs(3074)) or (layer0_outputs(5754));
    layer1_outputs(725) <= (layer0_outputs(3241)) or (layer0_outputs(7546));
    layer1_outputs(726) <= (layer0_outputs(5460)) and not (layer0_outputs(3763));
    layer1_outputs(727) <= '1';
    layer1_outputs(728) <= layer0_outputs(3288);
    layer1_outputs(729) <= layer0_outputs(1727);
    layer1_outputs(730) <= not((layer0_outputs(6302)) or (layer0_outputs(1686)));
    layer1_outputs(731) <= not(layer0_outputs(2191)) or (layer0_outputs(3054));
    layer1_outputs(732) <= (layer0_outputs(1875)) and not (layer0_outputs(6572));
    layer1_outputs(733) <= not(layer0_outputs(2415));
    layer1_outputs(734) <= not((layer0_outputs(2900)) and (layer0_outputs(5537)));
    layer1_outputs(735) <= (layer0_outputs(4081)) and (layer0_outputs(2556));
    layer1_outputs(736) <= (layer0_outputs(108)) or (layer0_outputs(7021));
    layer1_outputs(737) <= layer0_outputs(1677);
    layer1_outputs(738) <= '0';
    layer1_outputs(739) <= layer0_outputs(2599);
    layer1_outputs(740) <= not(layer0_outputs(6811));
    layer1_outputs(741) <= (layer0_outputs(1975)) and not (layer0_outputs(726));
    layer1_outputs(742) <= not((layer0_outputs(5830)) or (layer0_outputs(2005)));
    layer1_outputs(743) <= layer0_outputs(4944);
    layer1_outputs(744) <= not((layer0_outputs(7333)) or (layer0_outputs(3609)));
    layer1_outputs(745) <= not(layer0_outputs(5004)) or (layer0_outputs(7276));
    layer1_outputs(746) <= (layer0_outputs(6745)) and not (layer0_outputs(2102));
    layer1_outputs(747) <= not(layer0_outputs(7038));
    layer1_outputs(748) <= (layer0_outputs(7177)) and not (layer0_outputs(6722));
    layer1_outputs(749) <= (layer0_outputs(6566)) and not (layer0_outputs(4807));
    layer1_outputs(750) <= not((layer0_outputs(7334)) and (layer0_outputs(1508)));
    layer1_outputs(751) <= not(layer0_outputs(5505)) or (layer0_outputs(5806));
    layer1_outputs(752) <= not(layer0_outputs(3379)) or (layer0_outputs(3271));
    layer1_outputs(753) <= (layer0_outputs(857)) and not (layer0_outputs(7461));
    layer1_outputs(754) <= not(layer0_outputs(6301)) or (layer0_outputs(5529));
    layer1_outputs(755) <= layer0_outputs(3855);
    layer1_outputs(756) <= (layer0_outputs(2138)) and not (layer0_outputs(1761));
    layer1_outputs(757) <= (layer0_outputs(3906)) xor (layer0_outputs(3683));
    layer1_outputs(758) <= layer0_outputs(1773);
    layer1_outputs(759) <= layer0_outputs(1295);
    layer1_outputs(760) <= '0';
    layer1_outputs(761) <= not((layer0_outputs(5976)) and (layer0_outputs(7522)));
    layer1_outputs(762) <= (layer0_outputs(4675)) and (layer0_outputs(4872));
    layer1_outputs(763) <= not((layer0_outputs(3679)) or (layer0_outputs(1386)));
    layer1_outputs(764) <= not(layer0_outputs(2760)) or (layer0_outputs(305));
    layer1_outputs(765) <= '0';
    layer1_outputs(766) <= not(layer0_outputs(6265));
    layer1_outputs(767) <= layer0_outputs(4147);
    layer1_outputs(768) <= (layer0_outputs(883)) and not (layer0_outputs(7022));
    layer1_outputs(769) <= not(layer0_outputs(1892));
    layer1_outputs(770) <= not(layer0_outputs(5079)) or (layer0_outputs(4712));
    layer1_outputs(771) <= not(layer0_outputs(3977));
    layer1_outputs(772) <= '1';
    layer1_outputs(773) <= not(layer0_outputs(3945));
    layer1_outputs(774) <= not(layer0_outputs(879)) or (layer0_outputs(6601));
    layer1_outputs(775) <= (layer0_outputs(1958)) and not (layer0_outputs(4508));
    layer1_outputs(776) <= not(layer0_outputs(770));
    layer1_outputs(777) <= not((layer0_outputs(5454)) or (layer0_outputs(5736)));
    layer1_outputs(778) <= not(layer0_outputs(7361));
    layer1_outputs(779) <= not(layer0_outputs(5645));
    layer1_outputs(780) <= layer0_outputs(4010);
    layer1_outputs(781) <= not(layer0_outputs(6264));
    layer1_outputs(782) <= '0';
    layer1_outputs(783) <= '1';
    layer1_outputs(784) <= layer0_outputs(7527);
    layer1_outputs(785) <= not(layer0_outputs(1158));
    layer1_outputs(786) <= not(layer0_outputs(19));
    layer1_outputs(787) <= not(layer0_outputs(4589));
    layer1_outputs(788) <= not(layer0_outputs(5096));
    layer1_outputs(789) <= not(layer0_outputs(5338));
    layer1_outputs(790) <= (layer0_outputs(7241)) and not (layer0_outputs(7336));
    layer1_outputs(791) <= not(layer0_outputs(6757)) or (layer0_outputs(3738));
    layer1_outputs(792) <= (layer0_outputs(7584)) and (layer0_outputs(2998));
    layer1_outputs(793) <= (layer0_outputs(4549)) and not (layer0_outputs(4492));
    layer1_outputs(794) <= (layer0_outputs(2616)) and (layer0_outputs(3883));
    layer1_outputs(795) <= (layer0_outputs(5303)) and not (layer0_outputs(5395));
    layer1_outputs(796) <= '1';
    layer1_outputs(797) <= not(layer0_outputs(464));
    layer1_outputs(798) <= (layer0_outputs(11)) and not (layer0_outputs(3719));
    layer1_outputs(799) <= (layer0_outputs(3632)) and not (layer0_outputs(3562));
    layer1_outputs(800) <= (layer0_outputs(901)) and (layer0_outputs(5617));
    layer1_outputs(801) <= layer0_outputs(4104);
    layer1_outputs(802) <= (layer0_outputs(4794)) or (layer0_outputs(2051));
    layer1_outputs(803) <= '0';
    layer1_outputs(804) <= (layer0_outputs(320)) and not (layer0_outputs(6965));
    layer1_outputs(805) <= (layer0_outputs(6714)) and (layer0_outputs(1885));
    layer1_outputs(806) <= (layer0_outputs(5605)) or (layer0_outputs(4495));
    layer1_outputs(807) <= not((layer0_outputs(6596)) or (layer0_outputs(966)));
    layer1_outputs(808) <= (layer0_outputs(3701)) and (layer0_outputs(4185));
    layer1_outputs(809) <= '0';
    layer1_outputs(810) <= '1';
    layer1_outputs(811) <= not((layer0_outputs(5318)) or (layer0_outputs(2975)));
    layer1_outputs(812) <= not(layer0_outputs(1002));
    layer1_outputs(813) <= not(layer0_outputs(4458)) or (layer0_outputs(7641));
    layer1_outputs(814) <= not(layer0_outputs(3172));
    layer1_outputs(815) <= not(layer0_outputs(2929)) or (layer0_outputs(6560));
    layer1_outputs(816) <= layer0_outputs(2655);
    layer1_outputs(817) <= not(layer0_outputs(5071));
    layer1_outputs(818) <= (layer0_outputs(5030)) and not (layer0_outputs(2738));
    layer1_outputs(819) <= not(layer0_outputs(5813));
    layer1_outputs(820) <= not(layer0_outputs(5736)) or (layer0_outputs(497));
    layer1_outputs(821) <= not(layer0_outputs(5291));
    layer1_outputs(822) <= (layer0_outputs(2298)) or (layer0_outputs(490));
    layer1_outputs(823) <= '0';
    layer1_outputs(824) <= '0';
    layer1_outputs(825) <= not(layer0_outputs(1505));
    layer1_outputs(826) <= not((layer0_outputs(6171)) or (layer0_outputs(6652)));
    layer1_outputs(827) <= layer0_outputs(1594);
    layer1_outputs(828) <= layer0_outputs(5349);
    layer1_outputs(829) <= not(layer0_outputs(3484));
    layer1_outputs(830) <= not((layer0_outputs(3806)) or (layer0_outputs(5331)));
    layer1_outputs(831) <= '0';
    layer1_outputs(832) <= not(layer0_outputs(3345));
    layer1_outputs(833) <= (layer0_outputs(2145)) or (layer0_outputs(2413));
    layer1_outputs(834) <= not((layer0_outputs(2248)) and (layer0_outputs(4558)));
    layer1_outputs(835) <= '0';
    layer1_outputs(836) <= not(layer0_outputs(4547)) or (layer0_outputs(4887));
    layer1_outputs(837) <= layer0_outputs(4417);
    layer1_outputs(838) <= not((layer0_outputs(6293)) and (layer0_outputs(3336)));
    layer1_outputs(839) <= '1';
    layer1_outputs(840) <= (layer0_outputs(4852)) or (layer0_outputs(2487));
    layer1_outputs(841) <= '1';
    layer1_outputs(842) <= layer0_outputs(5978);
    layer1_outputs(843) <= (layer0_outputs(3395)) or (layer0_outputs(2630));
    layer1_outputs(844) <= not(layer0_outputs(5097)) or (layer0_outputs(6997));
    layer1_outputs(845) <= not(layer0_outputs(4153));
    layer1_outputs(846) <= (layer0_outputs(3222)) xor (layer0_outputs(4099));
    layer1_outputs(847) <= layer0_outputs(2992);
    layer1_outputs(848) <= '0';
    layer1_outputs(849) <= not(layer0_outputs(284));
    layer1_outputs(850) <= (layer0_outputs(5160)) and (layer0_outputs(6087));
    layer1_outputs(851) <= not(layer0_outputs(1358)) or (layer0_outputs(2689));
    layer1_outputs(852) <= (layer0_outputs(5304)) or (layer0_outputs(321));
    layer1_outputs(853) <= '1';
    layer1_outputs(854) <= '1';
    layer1_outputs(855) <= not(layer0_outputs(7361)) or (layer0_outputs(4666));
    layer1_outputs(856) <= layer0_outputs(1497);
    layer1_outputs(857) <= layer0_outputs(3763);
    layer1_outputs(858) <= '1';
    layer1_outputs(859) <= '0';
    layer1_outputs(860) <= not(layer0_outputs(4929));
    layer1_outputs(861) <= layer0_outputs(10);
    layer1_outputs(862) <= not(layer0_outputs(34));
    layer1_outputs(863) <= layer0_outputs(298);
    layer1_outputs(864) <= (layer0_outputs(5441)) and not (layer0_outputs(7547));
    layer1_outputs(865) <= not(layer0_outputs(2578));
    layer1_outputs(866) <= layer0_outputs(3731);
    layer1_outputs(867) <= (layer0_outputs(1597)) or (layer0_outputs(5859));
    layer1_outputs(868) <= not((layer0_outputs(1614)) and (layer0_outputs(2358)));
    layer1_outputs(869) <= not(layer0_outputs(2542)) or (layer0_outputs(1203));
    layer1_outputs(870) <= not((layer0_outputs(6172)) or (layer0_outputs(2392)));
    layer1_outputs(871) <= (layer0_outputs(200)) and not (layer0_outputs(6081));
    layer1_outputs(872) <= (layer0_outputs(7185)) or (layer0_outputs(1534));
    layer1_outputs(873) <= (layer0_outputs(4936)) and not (layer0_outputs(3059));
    layer1_outputs(874) <= '1';
    layer1_outputs(875) <= (layer0_outputs(839)) and not (layer0_outputs(1653));
    layer1_outputs(876) <= not(layer0_outputs(1555)) or (layer0_outputs(3751));
    layer1_outputs(877) <= (layer0_outputs(7421)) xor (layer0_outputs(1902));
    layer1_outputs(878) <= (layer0_outputs(4510)) and not (layer0_outputs(1996));
    layer1_outputs(879) <= '0';
    layer1_outputs(880) <= not((layer0_outputs(3568)) and (layer0_outputs(6848)));
    layer1_outputs(881) <= layer0_outputs(6890);
    layer1_outputs(882) <= layer0_outputs(2993);
    layer1_outputs(883) <= layer0_outputs(7116);
    layer1_outputs(884) <= not(layer0_outputs(6263));
    layer1_outputs(885) <= not((layer0_outputs(5912)) or (layer0_outputs(451)));
    layer1_outputs(886) <= layer0_outputs(1934);
    layer1_outputs(887) <= (layer0_outputs(373)) and not (layer0_outputs(2777));
    layer1_outputs(888) <= not((layer0_outputs(859)) or (layer0_outputs(2725)));
    layer1_outputs(889) <= not(layer0_outputs(2571));
    layer1_outputs(890) <= '0';
    layer1_outputs(891) <= not(layer0_outputs(1925)) or (layer0_outputs(7398));
    layer1_outputs(892) <= layer0_outputs(4691);
    layer1_outputs(893) <= (layer0_outputs(7363)) or (layer0_outputs(3197));
    layer1_outputs(894) <= not(layer0_outputs(2309)) or (layer0_outputs(5450));
    layer1_outputs(895) <= not(layer0_outputs(95));
    layer1_outputs(896) <= '1';
    layer1_outputs(897) <= not((layer0_outputs(4953)) xor (layer0_outputs(1897)));
    layer1_outputs(898) <= not((layer0_outputs(7597)) and (layer0_outputs(3362)));
    layer1_outputs(899) <= not(layer0_outputs(7574)) or (layer0_outputs(4769));
    layer1_outputs(900) <= (layer0_outputs(5217)) or (layer0_outputs(2690));
    layer1_outputs(901) <= not((layer0_outputs(2688)) or (layer0_outputs(1383)));
    layer1_outputs(902) <= not(layer0_outputs(6690)) or (layer0_outputs(6551));
    layer1_outputs(903) <= not(layer0_outputs(1293));
    layer1_outputs(904) <= (layer0_outputs(2120)) and not (layer0_outputs(5933));
    layer1_outputs(905) <= not((layer0_outputs(1486)) or (layer0_outputs(6210)));
    layer1_outputs(906) <= not(layer0_outputs(4029));
    layer1_outputs(907) <= (layer0_outputs(2925)) and not (layer0_outputs(3809));
    layer1_outputs(908) <= (layer0_outputs(4146)) and not (layer0_outputs(4169));
    layer1_outputs(909) <= '0';
    layer1_outputs(910) <= not((layer0_outputs(7562)) and (layer0_outputs(4991)));
    layer1_outputs(911) <= (layer0_outputs(7477)) or (layer0_outputs(4143));
    layer1_outputs(912) <= not(layer0_outputs(2948));
    layer1_outputs(913) <= not(layer0_outputs(6050)) or (layer0_outputs(2160));
    layer1_outputs(914) <= not((layer0_outputs(580)) and (layer0_outputs(5047)));
    layer1_outputs(915) <= '0';
    layer1_outputs(916) <= (layer0_outputs(3746)) and (layer0_outputs(1818));
    layer1_outputs(917) <= (layer0_outputs(5258)) and not (layer0_outputs(1629));
    layer1_outputs(918) <= not((layer0_outputs(1885)) or (layer0_outputs(6876)));
    layer1_outputs(919) <= not(layer0_outputs(6933));
    layer1_outputs(920) <= (layer0_outputs(1578)) or (layer0_outputs(5384));
    layer1_outputs(921) <= layer0_outputs(3894);
    layer1_outputs(922) <= '0';
    layer1_outputs(923) <= not(layer0_outputs(2626)) or (layer0_outputs(6573));
    layer1_outputs(924) <= not(layer0_outputs(3517));
    layer1_outputs(925) <= (layer0_outputs(4807)) and not (layer0_outputs(2770));
    layer1_outputs(926) <= '1';
    layer1_outputs(927) <= not(layer0_outputs(3538));
    layer1_outputs(928) <= layer0_outputs(1503);
    layer1_outputs(929) <= layer0_outputs(1536);
    layer1_outputs(930) <= not((layer0_outputs(6871)) or (layer0_outputs(3810)));
    layer1_outputs(931) <= layer0_outputs(3133);
    layer1_outputs(932) <= not(layer0_outputs(3597));
    layer1_outputs(933) <= layer0_outputs(2851);
    layer1_outputs(934) <= layer0_outputs(6191);
    layer1_outputs(935) <= not(layer0_outputs(3051));
    layer1_outputs(936) <= layer0_outputs(3595);
    layer1_outputs(937) <= (layer0_outputs(2096)) or (layer0_outputs(1600));
    layer1_outputs(938) <= not((layer0_outputs(3068)) and (layer0_outputs(900)));
    layer1_outputs(939) <= (layer0_outputs(658)) and not (layer0_outputs(332));
    layer1_outputs(940) <= not(layer0_outputs(1682)) or (layer0_outputs(6355));
    layer1_outputs(941) <= not(layer0_outputs(4144));
    layer1_outputs(942) <= not((layer0_outputs(5270)) xor (layer0_outputs(4549)));
    layer1_outputs(943) <= (layer0_outputs(1363)) or (layer0_outputs(1451));
    layer1_outputs(944) <= not((layer0_outputs(3028)) and (layer0_outputs(3375)));
    layer1_outputs(945) <= not(layer0_outputs(6063));
    layer1_outputs(946) <= not((layer0_outputs(5751)) and (layer0_outputs(80)));
    layer1_outputs(947) <= not(layer0_outputs(1624));
    layer1_outputs(948) <= not((layer0_outputs(7368)) xor (layer0_outputs(6683)));
    layer1_outputs(949) <= '1';
    layer1_outputs(950) <= not(layer0_outputs(3189));
    layer1_outputs(951) <= not((layer0_outputs(6714)) or (layer0_outputs(3619)));
    layer1_outputs(952) <= not(layer0_outputs(6950)) or (layer0_outputs(6554));
    layer1_outputs(953) <= '0';
    layer1_outputs(954) <= not(layer0_outputs(6496));
    layer1_outputs(955) <= not(layer0_outputs(6681)) or (layer0_outputs(1228));
    layer1_outputs(956) <= (layer0_outputs(317)) and not (layer0_outputs(1953));
    layer1_outputs(957) <= (layer0_outputs(114)) and not (layer0_outputs(6434));
    layer1_outputs(958) <= not(layer0_outputs(6786));
    layer1_outputs(959) <= (layer0_outputs(4823)) xor (layer0_outputs(7324));
    layer1_outputs(960) <= (layer0_outputs(4538)) and not (layer0_outputs(4262));
    layer1_outputs(961) <= '1';
    layer1_outputs(962) <= '1';
    layer1_outputs(963) <= not((layer0_outputs(6167)) and (layer0_outputs(3512)));
    layer1_outputs(964) <= (layer0_outputs(2810)) and not (layer0_outputs(7561));
    layer1_outputs(965) <= (layer0_outputs(926)) and (layer0_outputs(7391));
    layer1_outputs(966) <= (layer0_outputs(3966)) and not (layer0_outputs(1805));
    layer1_outputs(967) <= layer0_outputs(3582);
    layer1_outputs(968) <= layer0_outputs(3265);
    layer1_outputs(969) <= not(layer0_outputs(6271)) or (layer0_outputs(5256));
    layer1_outputs(970) <= layer0_outputs(1169);
    layer1_outputs(971) <= (layer0_outputs(1615)) or (layer0_outputs(3075));
    layer1_outputs(972) <= (layer0_outputs(329)) and not (layer0_outputs(5766));
    layer1_outputs(973) <= not(layer0_outputs(4007)) or (layer0_outputs(5521));
    layer1_outputs(974) <= not(layer0_outputs(206)) or (layer0_outputs(4637));
    layer1_outputs(975) <= not((layer0_outputs(5449)) and (layer0_outputs(7385)));
    layer1_outputs(976) <= not(layer0_outputs(954));
    layer1_outputs(977) <= not(layer0_outputs(5627)) or (layer0_outputs(678));
    layer1_outputs(978) <= '0';
    layer1_outputs(979) <= '1';
    layer1_outputs(980) <= not(layer0_outputs(5446));
    layer1_outputs(981) <= not(layer0_outputs(26)) or (layer0_outputs(6918));
    layer1_outputs(982) <= (layer0_outputs(6579)) and (layer0_outputs(7561));
    layer1_outputs(983) <= not(layer0_outputs(6079));
    layer1_outputs(984) <= not(layer0_outputs(1338)) or (layer0_outputs(3231));
    layer1_outputs(985) <= not(layer0_outputs(6721));
    layer1_outputs(986) <= layer0_outputs(4467);
    layer1_outputs(987) <= (layer0_outputs(275)) and not (layer0_outputs(3229));
    layer1_outputs(988) <= (layer0_outputs(5540)) and not (layer0_outputs(2219));
    layer1_outputs(989) <= (layer0_outputs(916)) and not (layer0_outputs(1823));
    layer1_outputs(990) <= layer0_outputs(4370);
    layer1_outputs(991) <= '0';
    layer1_outputs(992) <= (layer0_outputs(6476)) and not (layer0_outputs(7339));
    layer1_outputs(993) <= not((layer0_outputs(6867)) or (layer0_outputs(5282)));
    layer1_outputs(994) <= (layer0_outputs(2802)) and not (layer0_outputs(1143));
    layer1_outputs(995) <= '1';
    layer1_outputs(996) <= (layer0_outputs(7449)) and (layer0_outputs(2318));
    layer1_outputs(997) <= (layer0_outputs(318)) and (layer0_outputs(1781));
    layer1_outputs(998) <= (layer0_outputs(576)) and (layer0_outputs(2519));
    layer1_outputs(999) <= not(layer0_outputs(195));
    layer1_outputs(1000) <= not(layer0_outputs(1374)) or (layer0_outputs(1357));
    layer1_outputs(1001) <= (layer0_outputs(6078)) and not (layer0_outputs(2706));
    layer1_outputs(1002) <= not(layer0_outputs(7082)) or (layer0_outputs(6638));
    layer1_outputs(1003) <= not(layer0_outputs(7544)) or (layer0_outputs(4226));
    layer1_outputs(1004) <= (layer0_outputs(3421)) and not (layer0_outputs(3187));
    layer1_outputs(1005) <= (layer0_outputs(5118)) and (layer0_outputs(6298));
    layer1_outputs(1006) <= not(layer0_outputs(5637)) or (layer0_outputs(2621));
    layer1_outputs(1007) <= (layer0_outputs(3317)) or (layer0_outputs(1911));
    layer1_outputs(1008) <= not(layer0_outputs(1003)) or (layer0_outputs(3214));
    layer1_outputs(1009) <= (layer0_outputs(4642)) and (layer0_outputs(3343));
    layer1_outputs(1010) <= not(layer0_outputs(809)) or (layer0_outputs(1958));
    layer1_outputs(1011) <= not(layer0_outputs(7303)) or (layer0_outputs(7543));
    layer1_outputs(1012) <= '0';
    layer1_outputs(1013) <= layer0_outputs(1243);
    layer1_outputs(1014) <= (layer0_outputs(5280)) and not (layer0_outputs(3072));
    layer1_outputs(1015) <= (layer0_outputs(6151)) and not (layer0_outputs(4451));
    layer1_outputs(1016) <= not((layer0_outputs(3223)) xor (layer0_outputs(6402)));
    layer1_outputs(1017) <= (layer0_outputs(6637)) and not (layer0_outputs(7431));
    layer1_outputs(1018) <= (layer0_outputs(5809)) and not (layer0_outputs(1195));
    layer1_outputs(1019) <= not((layer0_outputs(4470)) and (layer0_outputs(2400)));
    layer1_outputs(1020) <= not((layer0_outputs(4821)) or (layer0_outputs(4616)));
    layer1_outputs(1021) <= not(layer0_outputs(1469));
    layer1_outputs(1022) <= layer0_outputs(2317);
    layer1_outputs(1023) <= (layer0_outputs(96)) and not (layer0_outputs(472));
    layer1_outputs(1024) <= '0';
    layer1_outputs(1025) <= '0';
    layer1_outputs(1026) <= '0';
    layer1_outputs(1027) <= not((layer0_outputs(4)) and (layer0_outputs(4120)));
    layer1_outputs(1028) <= (layer0_outputs(5990)) and (layer0_outputs(1330));
    layer1_outputs(1029) <= not((layer0_outputs(7373)) or (layer0_outputs(7422)));
    layer1_outputs(1030) <= not(layer0_outputs(1645)) or (layer0_outputs(4696));
    layer1_outputs(1031) <= layer0_outputs(3662);
    layer1_outputs(1032) <= not((layer0_outputs(7191)) and (layer0_outputs(1353)));
    layer1_outputs(1033) <= '0';
    layer1_outputs(1034) <= not((layer0_outputs(5417)) and (layer0_outputs(881)));
    layer1_outputs(1035) <= (layer0_outputs(4476)) xor (layer0_outputs(655));
    layer1_outputs(1036) <= not(layer0_outputs(4757)) or (layer0_outputs(5015));
    layer1_outputs(1037) <= layer0_outputs(7306);
    layer1_outputs(1038) <= not(layer0_outputs(6099)) or (layer0_outputs(6479));
    layer1_outputs(1039) <= '0';
    layer1_outputs(1040) <= '1';
    layer1_outputs(1041) <= '1';
    layer1_outputs(1042) <= not(layer0_outputs(1424));
    layer1_outputs(1043) <= (layer0_outputs(3449)) xor (layer0_outputs(3545));
    layer1_outputs(1044) <= (layer0_outputs(5598)) or (layer0_outputs(6558));
    layer1_outputs(1045) <= not((layer0_outputs(232)) or (layer0_outputs(4324)));
    layer1_outputs(1046) <= (layer0_outputs(2125)) and (layer0_outputs(3577));
    layer1_outputs(1047) <= layer0_outputs(1869);
    layer1_outputs(1048) <= not((layer0_outputs(4886)) and (layer0_outputs(612)));
    layer1_outputs(1049) <= (layer0_outputs(4360)) and not (layer0_outputs(450));
    layer1_outputs(1050) <= (layer0_outputs(341)) and not (layer0_outputs(4710));
    layer1_outputs(1051) <= not((layer0_outputs(5025)) or (layer0_outputs(2780)));
    layer1_outputs(1052) <= not(layer0_outputs(2517));
    layer1_outputs(1053) <= not(layer0_outputs(5865));
    layer1_outputs(1054) <= not(layer0_outputs(2613));
    layer1_outputs(1055) <= (layer0_outputs(3046)) and (layer0_outputs(7529));
    layer1_outputs(1056) <= '0';
    layer1_outputs(1057) <= layer0_outputs(1193);
    layer1_outputs(1058) <= layer0_outputs(6529);
    layer1_outputs(1059) <= layer0_outputs(3856);
    layer1_outputs(1060) <= '0';
    layer1_outputs(1061) <= (layer0_outputs(3387)) and not (layer0_outputs(6450));
    layer1_outputs(1062) <= not(layer0_outputs(7580));
    layer1_outputs(1063) <= (layer0_outputs(5116)) and (layer0_outputs(5700));
    layer1_outputs(1064) <= '0';
    layer1_outputs(1065) <= not((layer0_outputs(5127)) xor (layer0_outputs(1151)));
    layer1_outputs(1066) <= (layer0_outputs(1128)) or (layer0_outputs(1056));
    layer1_outputs(1067) <= '1';
    layer1_outputs(1068) <= not(layer0_outputs(3902));
    layer1_outputs(1069) <= layer0_outputs(562);
    layer1_outputs(1070) <= (layer0_outputs(4)) or (layer0_outputs(2405));
    layer1_outputs(1071) <= layer0_outputs(892);
    layer1_outputs(1072) <= (layer0_outputs(154)) xor (layer0_outputs(2637));
    layer1_outputs(1073) <= layer0_outputs(6345);
    layer1_outputs(1074) <= '1';
    layer1_outputs(1075) <= '1';
    layer1_outputs(1076) <= (layer0_outputs(5145)) and (layer0_outputs(6527));
    layer1_outputs(1077) <= not((layer0_outputs(3529)) and (layer0_outputs(7464)));
    layer1_outputs(1078) <= layer0_outputs(1908);
    layer1_outputs(1079) <= not(layer0_outputs(7451));
    layer1_outputs(1080) <= not(layer0_outputs(5245));
    layer1_outputs(1081) <= '1';
    layer1_outputs(1082) <= not((layer0_outputs(5524)) or (layer0_outputs(4568)));
    layer1_outputs(1083) <= layer0_outputs(3651);
    layer1_outputs(1084) <= not((layer0_outputs(5962)) and (layer0_outputs(5870)));
    layer1_outputs(1085) <= layer0_outputs(6715);
    layer1_outputs(1086) <= '1';
    layer1_outputs(1087) <= layer0_outputs(4213);
    layer1_outputs(1088) <= not(layer0_outputs(1966));
    layer1_outputs(1089) <= '1';
    layer1_outputs(1090) <= '0';
    layer1_outputs(1091) <= not((layer0_outputs(6158)) or (layer0_outputs(7243)));
    layer1_outputs(1092) <= not(layer0_outputs(7067));
    layer1_outputs(1093) <= layer0_outputs(1309);
    layer1_outputs(1094) <= (layer0_outputs(1399)) xor (layer0_outputs(4071));
    layer1_outputs(1095) <= not(layer0_outputs(5569)) or (layer0_outputs(1144));
    layer1_outputs(1096) <= (layer0_outputs(805)) and (layer0_outputs(7559));
    layer1_outputs(1097) <= not(layer0_outputs(6841));
    layer1_outputs(1098) <= '0';
    layer1_outputs(1099) <= '1';
    layer1_outputs(1100) <= not(layer0_outputs(3182));
    layer1_outputs(1101) <= not(layer0_outputs(7053));
    layer1_outputs(1102) <= layer0_outputs(3823);
    layer1_outputs(1103) <= layer0_outputs(5371);
    layer1_outputs(1104) <= layer0_outputs(4871);
    layer1_outputs(1105) <= (layer0_outputs(849)) and (layer0_outputs(4173));
    layer1_outputs(1106) <= (layer0_outputs(1756)) or (layer0_outputs(1716));
    layer1_outputs(1107) <= not((layer0_outputs(5455)) and (layer0_outputs(4713)));
    layer1_outputs(1108) <= not(layer0_outputs(2555)) or (layer0_outputs(5297));
    layer1_outputs(1109) <= not(layer0_outputs(1504));
    layer1_outputs(1110) <= (layer0_outputs(3405)) and not (layer0_outputs(1660));
    layer1_outputs(1111) <= (layer0_outputs(7676)) and not (layer0_outputs(3703));
    layer1_outputs(1112) <= '0';
    layer1_outputs(1113) <= not((layer0_outputs(4018)) or (layer0_outputs(4928)));
    layer1_outputs(1114) <= not((layer0_outputs(2410)) and (layer0_outputs(7294)));
    layer1_outputs(1115) <= not(layer0_outputs(5030)) or (layer0_outputs(5611));
    layer1_outputs(1116) <= not((layer0_outputs(4323)) or (layer0_outputs(4934)));
    layer1_outputs(1117) <= not(layer0_outputs(5874)) or (layer0_outputs(5280));
    layer1_outputs(1118) <= '0';
    layer1_outputs(1119) <= (layer0_outputs(7359)) or (layer0_outputs(1778));
    layer1_outputs(1120) <= layer0_outputs(2154);
    layer1_outputs(1121) <= not(layer0_outputs(3688)) or (layer0_outputs(3424));
    layer1_outputs(1122) <= not(layer0_outputs(2912));
    layer1_outputs(1123) <= not((layer0_outputs(4057)) xor (layer0_outputs(1672)));
    layer1_outputs(1124) <= (layer0_outputs(4680)) and not (layer0_outputs(5061));
    layer1_outputs(1125) <= (layer0_outputs(3019)) and not (layer0_outputs(1033));
    layer1_outputs(1126) <= (layer0_outputs(1808)) and not (layer0_outputs(6212));
    layer1_outputs(1127) <= layer0_outputs(2408);
    layer1_outputs(1128) <= '1';
    layer1_outputs(1129) <= not((layer0_outputs(1457)) and (layer0_outputs(5596)));
    layer1_outputs(1130) <= not(layer0_outputs(3924));
    layer1_outputs(1131) <= (layer0_outputs(6584)) and not (layer0_outputs(5113));
    layer1_outputs(1132) <= not(layer0_outputs(4623)) or (layer0_outputs(5838));
    layer1_outputs(1133) <= (layer0_outputs(6510)) and not (layer0_outputs(4956));
    layer1_outputs(1134) <= not(layer0_outputs(5634)) or (layer0_outputs(3826));
    layer1_outputs(1135) <= not((layer0_outputs(3698)) or (layer0_outputs(584)));
    layer1_outputs(1136) <= not(layer0_outputs(4037));
    layer1_outputs(1137) <= not((layer0_outputs(3520)) or (layer0_outputs(6366)));
    layer1_outputs(1138) <= (layer0_outputs(2285)) or (layer0_outputs(151));
    layer1_outputs(1139) <= not(layer0_outputs(7119)) or (layer0_outputs(5778));
    layer1_outputs(1140) <= (layer0_outputs(4045)) or (layer0_outputs(6443));
    layer1_outputs(1141) <= (layer0_outputs(7579)) and not (layer0_outputs(5000));
    layer1_outputs(1142) <= not(layer0_outputs(3414)) or (layer0_outputs(6014));
    layer1_outputs(1143) <= (layer0_outputs(4533)) or (layer0_outputs(5616));
    layer1_outputs(1144) <= not(layer0_outputs(1429));
    layer1_outputs(1145) <= not((layer0_outputs(6883)) xor (layer0_outputs(5652)));
    layer1_outputs(1146) <= layer0_outputs(5041);
    layer1_outputs(1147) <= not((layer0_outputs(3130)) or (layer0_outputs(6145)));
    layer1_outputs(1148) <= not(layer0_outputs(6578));
    layer1_outputs(1149) <= not(layer0_outputs(2559)) or (layer0_outputs(2062));
    layer1_outputs(1150) <= (layer0_outputs(1659)) and not (layer0_outputs(246));
    layer1_outputs(1151) <= (layer0_outputs(7480)) and not (layer0_outputs(6683));
    layer1_outputs(1152) <= layer0_outputs(4282);
    layer1_outputs(1153) <= not(layer0_outputs(5744)) or (layer0_outputs(4531));
    layer1_outputs(1154) <= '0';
    layer1_outputs(1155) <= (layer0_outputs(5553)) and not (layer0_outputs(4397));
    layer1_outputs(1156) <= '1';
    layer1_outputs(1157) <= (layer0_outputs(7089)) and not (layer0_outputs(603));
    layer1_outputs(1158) <= (layer0_outputs(5744)) and (layer0_outputs(1205));
    layer1_outputs(1159) <= layer0_outputs(6810);
    layer1_outputs(1160) <= not(layer0_outputs(2085)) or (layer0_outputs(1791));
    layer1_outputs(1161) <= '0';
    layer1_outputs(1162) <= layer0_outputs(718);
    layer1_outputs(1163) <= (layer0_outputs(4622)) and not (layer0_outputs(704));
    layer1_outputs(1164) <= not((layer0_outputs(4724)) and (layer0_outputs(5917)));
    layer1_outputs(1165) <= '1';
    layer1_outputs(1166) <= layer0_outputs(2296);
    layer1_outputs(1167) <= (layer0_outputs(7519)) xor (layer0_outputs(3150));
    layer1_outputs(1168) <= layer0_outputs(4277);
    layer1_outputs(1169) <= layer0_outputs(1191);
    layer1_outputs(1170) <= not((layer0_outputs(6148)) or (layer0_outputs(1152)));
    layer1_outputs(1171) <= not((layer0_outputs(5884)) xor (layer0_outputs(1589)));
    layer1_outputs(1172) <= '0';
    layer1_outputs(1173) <= not(layer0_outputs(4274)) or (layer0_outputs(4661));
    layer1_outputs(1174) <= '1';
    layer1_outputs(1175) <= not(layer0_outputs(5780)) or (layer0_outputs(1055));
    layer1_outputs(1176) <= not(layer0_outputs(7566)) or (layer0_outputs(5772));
    layer1_outputs(1177) <= not(layer0_outputs(4384)) or (layer0_outputs(5424));
    layer1_outputs(1178) <= not((layer0_outputs(5478)) or (layer0_outputs(339)));
    layer1_outputs(1179) <= '1';
    layer1_outputs(1180) <= not(layer0_outputs(6153));
    layer1_outputs(1181) <= (layer0_outputs(2736)) and not (layer0_outputs(2037));
    layer1_outputs(1182) <= layer0_outputs(6168);
    layer1_outputs(1183) <= not((layer0_outputs(6178)) or (layer0_outputs(6173)));
    layer1_outputs(1184) <= '1';
    layer1_outputs(1185) <= (layer0_outputs(6973)) or (layer0_outputs(1023));
    layer1_outputs(1186) <= (layer0_outputs(81)) and not (layer0_outputs(5954));
    layer1_outputs(1187) <= (layer0_outputs(7611)) and (layer0_outputs(3066));
    layer1_outputs(1188) <= layer0_outputs(4193);
    layer1_outputs(1189) <= not(layer0_outputs(4569));
    layer1_outputs(1190) <= not(layer0_outputs(7507)) or (layer0_outputs(6313));
    layer1_outputs(1191) <= layer0_outputs(2700);
    layer1_outputs(1192) <= (layer0_outputs(6391)) or (layer0_outputs(198));
    layer1_outputs(1193) <= '0';
    layer1_outputs(1194) <= '0';
    layer1_outputs(1195) <= not((layer0_outputs(1852)) and (layer0_outputs(7619)));
    layer1_outputs(1196) <= (layer0_outputs(1545)) and (layer0_outputs(2792));
    layer1_outputs(1197) <= (layer0_outputs(5582)) xor (layer0_outputs(1053));
    layer1_outputs(1198) <= (layer0_outputs(3533)) or (layer0_outputs(4495));
    layer1_outputs(1199) <= (layer0_outputs(179)) and not (layer0_outputs(1712));
    layer1_outputs(1200) <= (layer0_outputs(3151)) or (layer0_outputs(3711));
    layer1_outputs(1201) <= (layer0_outputs(619)) or (layer0_outputs(4311));
    layer1_outputs(1202) <= layer0_outputs(3172);
    layer1_outputs(1203) <= not((layer0_outputs(4231)) or (layer0_outputs(2903)));
    layer1_outputs(1204) <= (layer0_outputs(1904)) and (layer0_outputs(7643));
    layer1_outputs(1205) <= not((layer0_outputs(4839)) or (layer0_outputs(816)));
    layer1_outputs(1206) <= (layer0_outputs(5236)) and not (layer0_outputs(7308));
    layer1_outputs(1207) <= not(layer0_outputs(1373));
    layer1_outputs(1208) <= not(layer0_outputs(3661));
    layer1_outputs(1209) <= (layer0_outputs(5117)) and (layer0_outputs(1515));
    layer1_outputs(1210) <= (layer0_outputs(2943)) and (layer0_outputs(1628));
    layer1_outputs(1211) <= not((layer0_outputs(3514)) or (layer0_outputs(5918)));
    layer1_outputs(1212) <= layer0_outputs(4837);
    layer1_outputs(1213) <= not(layer0_outputs(263));
    layer1_outputs(1214) <= not(layer0_outputs(4023)) or (layer0_outputs(6666));
    layer1_outputs(1215) <= not(layer0_outputs(15)) or (layer0_outputs(4052));
    layer1_outputs(1216) <= not(layer0_outputs(3507));
    layer1_outputs(1217) <= not(layer0_outputs(5378));
    layer1_outputs(1218) <= (layer0_outputs(1405)) and not (layer0_outputs(3359));
    layer1_outputs(1219) <= '0';
    layer1_outputs(1220) <= '1';
    layer1_outputs(1221) <= '0';
    layer1_outputs(1222) <= not((layer0_outputs(3078)) and (layer0_outputs(1436)));
    layer1_outputs(1223) <= not(layer0_outputs(2880));
    layer1_outputs(1224) <= (layer0_outputs(4470)) and (layer0_outputs(6823));
    layer1_outputs(1225) <= '0';
    layer1_outputs(1226) <= not((layer0_outputs(274)) xor (layer0_outputs(1076)));
    layer1_outputs(1227) <= (layer0_outputs(1248)) and not (layer0_outputs(2322));
    layer1_outputs(1228) <= layer0_outputs(5139);
    layer1_outputs(1229) <= '1';
    layer1_outputs(1230) <= not(layer0_outputs(2331));
    layer1_outputs(1231) <= layer0_outputs(2817);
    layer1_outputs(1232) <= not(layer0_outputs(3044));
    layer1_outputs(1233) <= not(layer0_outputs(7308));
    layer1_outputs(1234) <= not((layer0_outputs(4275)) and (layer0_outputs(1931)));
    layer1_outputs(1235) <= not(layer0_outputs(618));
    layer1_outputs(1236) <= '1';
    layer1_outputs(1237) <= not(layer0_outputs(5999)) or (layer0_outputs(4503));
    layer1_outputs(1238) <= (layer0_outputs(5311)) and not (layer0_outputs(1069));
    layer1_outputs(1239) <= layer0_outputs(7152);
    layer1_outputs(1240) <= '0';
    layer1_outputs(1241) <= (layer0_outputs(6592)) or (layer0_outputs(5947));
    layer1_outputs(1242) <= layer0_outputs(1860);
    layer1_outputs(1243) <= layer0_outputs(1962);
    layer1_outputs(1244) <= not(layer0_outputs(238)) or (layer0_outputs(722));
    layer1_outputs(1245) <= layer0_outputs(46);
    layer1_outputs(1246) <= not(layer0_outputs(4636)) or (layer0_outputs(3208));
    layer1_outputs(1247) <= not(layer0_outputs(2163));
    layer1_outputs(1248) <= '1';
    layer1_outputs(1249) <= not((layer0_outputs(3293)) and (layer0_outputs(7080)));
    layer1_outputs(1250) <= layer0_outputs(1887);
    layer1_outputs(1251) <= (layer0_outputs(2960)) xor (layer0_outputs(6810));
    layer1_outputs(1252) <= (layer0_outputs(4032)) and not (layer0_outputs(166));
    layer1_outputs(1253) <= (layer0_outputs(1564)) or (layer0_outputs(3777));
    layer1_outputs(1254) <= (layer0_outputs(5972)) and not (layer0_outputs(6197));
    layer1_outputs(1255) <= not(layer0_outputs(3585));
    layer1_outputs(1256) <= not((layer0_outputs(6506)) or (layer0_outputs(2748)));
    layer1_outputs(1257) <= not(layer0_outputs(3870));
    layer1_outputs(1258) <= '1';
    layer1_outputs(1259) <= '0';
    layer1_outputs(1260) <= '1';
    layer1_outputs(1261) <= layer0_outputs(1285);
    layer1_outputs(1262) <= not(layer0_outputs(4188));
    layer1_outputs(1263) <= layer0_outputs(3612);
    layer1_outputs(1264) <= (layer0_outputs(7009)) and (layer0_outputs(5797));
    layer1_outputs(1265) <= not(layer0_outputs(3684)) or (layer0_outputs(671));
    layer1_outputs(1266) <= layer0_outputs(813);
    layer1_outputs(1267) <= not((layer0_outputs(7444)) and (layer0_outputs(2688)));
    layer1_outputs(1268) <= (layer0_outputs(1648)) and not (layer0_outputs(2417));
    layer1_outputs(1269) <= layer0_outputs(3115);
    layer1_outputs(1270) <= (layer0_outputs(3805)) and not (layer0_outputs(433));
    layer1_outputs(1271) <= not(layer0_outputs(5062)) or (layer0_outputs(7138));
    layer1_outputs(1272) <= not(layer0_outputs(1082)) or (layer0_outputs(6911));
    layer1_outputs(1273) <= layer0_outputs(3048);
    layer1_outputs(1274) <= not(layer0_outputs(7588)) or (layer0_outputs(1375));
    layer1_outputs(1275) <= '0';
    layer1_outputs(1276) <= (layer0_outputs(4387)) and not (layer0_outputs(1664));
    layer1_outputs(1277) <= (layer0_outputs(7669)) and not (layer0_outputs(1502));
    layer1_outputs(1278) <= (layer0_outputs(6272)) and not (layer0_outputs(7178));
    layer1_outputs(1279) <= '1';
    layer1_outputs(1280) <= not(layer0_outputs(980)) or (layer0_outputs(1244));
    layer1_outputs(1281) <= not(layer0_outputs(1805)) or (layer0_outputs(7203));
    layer1_outputs(1282) <= not((layer0_outputs(4355)) and (layer0_outputs(7198)));
    layer1_outputs(1283) <= layer0_outputs(7498);
    layer1_outputs(1284) <= not(layer0_outputs(4190));
    layer1_outputs(1285) <= not(layer0_outputs(6138));
    layer1_outputs(1286) <= not(layer0_outputs(3865));
    layer1_outputs(1287) <= (layer0_outputs(5035)) and not (layer0_outputs(7215));
    layer1_outputs(1288) <= not((layer0_outputs(47)) xor (layer0_outputs(4391)));
    layer1_outputs(1289) <= not((layer0_outputs(772)) and (layer0_outputs(3691)));
    layer1_outputs(1290) <= (layer0_outputs(7142)) and not (layer0_outputs(5268));
    layer1_outputs(1291) <= (layer0_outputs(4821)) and not (layer0_outputs(5297));
    layer1_outputs(1292) <= not(layer0_outputs(3779)) or (layer0_outputs(2330));
    layer1_outputs(1293) <= '1';
    layer1_outputs(1294) <= not(layer0_outputs(6455));
    layer1_outputs(1295) <= (layer0_outputs(7213)) and (layer0_outputs(2781));
    layer1_outputs(1296) <= layer0_outputs(2083);
    layer1_outputs(1297) <= (layer0_outputs(5551)) and not (layer0_outputs(1065));
    layer1_outputs(1298) <= (layer0_outputs(1108)) and (layer0_outputs(3248));
    layer1_outputs(1299) <= layer0_outputs(6356);
    layer1_outputs(1300) <= (layer0_outputs(2669)) and not (layer0_outputs(3064));
    layer1_outputs(1301) <= (layer0_outputs(2328)) and not (layer0_outputs(6444));
    layer1_outputs(1302) <= not(layer0_outputs(521));
    layer1_outputs(1303) <= (layer0_outputs(6607)) and not (layer0_outputs(2131));
    layer1_outputs(1304) <= layer0_outputs(6920);
    layer1_outputs(1305) <= not(layer0_outputs(4833));
    layer1_outputs(1306) <= not(layer0_outputs(5263)) or (layer0_outputs(4274));
    layer1_outputs(1307) <= not(layer0_outputs(4461));
    layer1_outputs(1308) <= '1';
    layer1_outputs(1309) <= (layer0_outputs(3371)) or (layer0_outputs(1914));
    layer1_outputs(1310) <= layer0_outputs(3066);
    layer1_outputs(1311) <= not((layer0_outputs(6129)) or (layer0_outputs(2732)));
    layer1_outputs(1312) <= '1';
    layer1_outputs(1313) <= (layer0_outputs(5368)) or (layer0_outputs(4853));
    layer1_outputs(1314) <= not(layer0_outputs(409));
    layer1_outputs(1315) <= '1';
    layer1_outputs(1316) <= layer0_outputs(3485);
    layer1_outputs(1317) <= '0';
    layer1_outputs(1318) <= not(layer0_outputs(7064)) or (layer0_outputs(7069));
    layer1_outputs(1319) <= not(layer0_outputs(6074));
    layer1_outputs(1320) <= '1';
    layer1_outputs(1321) <= (layer0_outputs(4944)) and not (layer0_outputs(1104));
    layer1_outputs(1322) <= not(layer0_outputs(4018));
    layer1_outputs(1323) <= not(layer0_outputs(7292)) or (layer0_outputs(4112));
    layer1_outputs(1324) <= '1';
    layer1_outputs(1325) <= layer0_outputs(3134);
    layer1_outputs(1326) <= layer0_outputs(4473);
    layer1_outputs(1327) <= layer0_outputs(2835);
    layer1_outputs(1328) <= not(layer0_outputs(623)) or (layer0_outputs(2870));
    layer1_outputs(1329) <= '0';
    layer1_outputs(1330) <= not(layer0_outputs(5155)) or (layer0_outputs(3821));
    layer1_outputs(1331) <= not((layer0_outputs(5371)) and (layer0_outputs(5141)));
    layer1_outputs(1332) <= '1';
    layer1_outputs(1333) <= not(layer0_outputs(6075)) or (layer0_outputs(566));
    layer1_outputs(1334) <= '1';
    layer1_outputs(1335) <= layer0_outputs(56);
    layer1_outputs(1336) <= '0';
    layer1_outputs(1337) <= not((layer0_outputs(1220)) or (layer0_outputs(5620)));
    layer1_outputs(1338) <= not((layer0_outputs(5124)) or (layer0_outputs(270)));
    layer1_outputs(1339) <= layer0_outputs(622);
    layer1_outputs(1340) <= not(layer0_outputs(5784));
    layer1_outputs(1341) <= not((layer0_outputs(1291)) or (layer0_outputs(5706)));
    layer1_outputs(1342) <= not((layer0_outputs(4421)) xor (layer0_outputs(6846)));
    layer1_outputs(1343) <= layer0_outputs(1534);
    layer1_outputs(1344) <= (layer0_outputs(3936)) or (layer0_outputs(4597));
    layer1_outputs(1345) <= not((layer0_outputs(7542)) and (layer0_outputs(4347)));
    layer1_outputs(1346) <= layer0_outputs(4242);
    layer1_outputs(1347) <= (layer0_outputs(6411)) and not (layer0_outputs(4552));
    layer1_outputs(1348) <= not((layer0_outputs(2343)) or (layer0_outputs(3748)));
    layer1_outputs(1349) <= (layer0_outputs(4432)) or (layer0_outputs(6020));
    layer1_outputs(1350) <= '1';
    layer1_outputs(1351) <= not(layer0_outputs(4632));
    layer1_outputs(1352) <= not((layer0_outputs(3395)) or (layer0_outputs(1282)));
    layer1_outputs(1353) <= not((layer0_outputs(5692)) or (layer0_outputs(6750)));
    layer1_outputs(1354) <= not((layer0_outputs(4159)) and (layer0_outputs(6391)));
    layer1_outputs(1355) <= not(layer0_outputs(1395));
    layer1_outputs(1356) <= layer0_outputs(4592);
    layer1_outputs(1357) <= not(layer0_outputs(3479));
    layer1_outputs(1358) <= not(layer0_outputs(872)) or (layer0_outputs(6651));
    layer1_outputs(1359) <= not((layer0_outputs(5078)) or (layer0_outputs(2089)));
    layer1_outputs(1360) <= '0';
    layer1_outputs(1361) <= '0';
    layer1_outputs(1362) <= not(layer0_outputs(387)) or (layer0_outputs(2684));
    layer1_outputs(1363) <= not((layer0_outputs(2825)) and (layer0_outputs(6745)));
    layer1_outputs(1364) <= (layer0_outputs(6258)) and not (layer0_outputs(6874));
    layer1_outputs(1365) <= not((layer0_outputs(6544)) or (layer0_outputs(3983)));
    layer1_outputs(1366) <= not((layer0_outputs(7049)) or (layer0_outputs(1853)));
    layer1_outputs(1367) <= not((layer0_outputs(5335)) and (layer0_outputs(7078)));
    layer1_outputs(1368) <= (layer0_outputs(507)) and (layer0_outputs(3592));
    layer1_outputs(1369) <= '1';
    layer1_outputs(1370) <= '0';
    layer1_outputs(1371) <= '1';
    layer1_outputs(1372) <= (layer0_outputs(517)) and (layer0_outputs(5099));
    layer1_outputs(1373) <= (layer0_outputs(6616)) and not (layer0_outputs(5068));
    layer1_outputs(1374) <= (layer0_outputs(2272)) and (layer0_outputs(3368));
    layer1_outputs(1375) <= not(layer0_outputs(35));
    layer1_outputs(1376) <= layer0_outputs(2039);
    layer1_outputs(1377) <= (layer0_outputs(7485)) or (layer0_outputs(2507));
    layer1_outputs(1378) <= not(layer0_outputs(4565));
    layer1_outputs(1379) <= (layer0_outputs(5385)) and (layer0_outputs(2951));
    layer1_outputs(1380) <= not(layer0_outputs(137));
    layer1_outputs(1381) <= (layer0_outputs(1212)) and not (layer0_outputs(3853));
    layer1_outputs(1382) <= (layer0_outputs(5939)) xor (layer0_outputs(6034));
    layer1_outputs(1383) <= layer0_outputs(1445);
    layer1_outputs(1384) <= layer0_outputs(4067);
    layer1_outputs(1385) <= not((layer0_outputs(6116)) and (layer0_outputs(2883)));
    layer1_outputs(1386) <= (layer0_outputs(63)) or (layer0_outputs(3454));
    layer1_outputs(1387) <= not((layer0_outputs(1981)) or (layer0_outputs(720)));
    layer1_outputs(1388) <= not(layer0_outputs(4389));
    layer1_outputs(1389) <= not(layer0_outputs(3674)) or (layer0_outputs(2731));
    layer1_outputs(1390) <= not(layer0_outputs(3807));
    layer1_outputs(1391) <= (layer0_outputs(1054)) and not (layer0_outputs(6208));
    layer1_outputs(1392) <= '1';
    layer1_outputs(1393) <= not(layer0_outputs(4554)) or (layer0_outputs(493));
    layer1_outputs(1394) <= (layer0_outputs(7237)) xor (layer0_outputs(2532));
    layer1_outputs(1395) <= not(layer0_outputs(560)) or (layer0_outputs(3596));
    layer1_outputs(1396) <= (layer0_outputs(4421)) or (layer0_outputs(4881));
    layer1_outputs(1397) <= not(layer0_outputs(2137)) or (layer0_outputs(6647));
    layer1_outputs(1398) <= layer0_outputs(936);
    layer1_outputs(1399) <= layer0_outputs(3216);
    layer1_outputs(1400) <= (layer0_outputs(4186)) or (layer0_outputs(5513));
    layer1_outputs(1401) <= '0';
    layer1_outputs(1402) <= '0';
    layer1_outputs(1403) <= not(layer0_outputs(6798));
    layer1_outputs(1404) <= layer0_outputs(4630);
    layer1_outputs(1405) <= not(layer0_outputs(5828)) or (layer0_outputs(106));
    layer1_outputs(1406) <= not(layer0_outputs(5693)) or (layer0_outputs(1752));
    layer1_outputs(1407) <= not((layer0_outputs(6999)) or (layer0_outputs(4920)));
    layer1_outputs(1408) <= (layer0_outputs(4630)) and not (layer0_outputs(7673));
    layer1_outputs(1409) <= not((layer0_outputs(7109)) or (layer0_outputs(3113)));
    layer1_outputs(1410) <= '0';
    layer1_outputs(1411) <= not(layer0_outputs(613)) or (layer0_outputs(5470));
    layer1_outputs(1412) <= not((layer0_outputs(3080)) or (layer0_outputs(1355)));
    layer1_outputs(1413) <= (layer0_outputs(5498)) and (layer0_outputs(5876));
    layer1_outputs(1414) <= '0';
    layer1_outputs(1415) <= not(layer0_outputs(4761));
    layer1_outputs(1416) <= not(layer0_outputs(3435));
    layer1_outputs(1417) <= layer0_outputs(597);
    layer1_outputs(1418) <= (layer0_outputs(5658)) or (layer0_outputs(1035));
    layer1_outputs(1419) <= (layer0_outputs(934)) xor (layer0_outputs(5593));
    layer1_outputs(1420) <= (layer0_outputs(6100)) and (layer0_outputs(576));
    layer1_outputs(1421) <= layer0_outputs(7488);
    layer1_outputs(1422) <= not(layer0_outputs(4053)) or (layer0_outputs(2552));
    layer1_outputs(1423) <= '0';
    layer1_outputs(1424) <= not(layer0_outputs(7134)) or (layer0_outputs(4114));
    layer1_outputs(1425) <= layer0_outputs(3211);
    layer1_outputs(1426) <= layer0_outputs(507);
    layer1_outputs(1427) <= '0';
    layer1_outputs(1428) <= layer0_outputs(173);
    layer1_outputs(1429) <= layer0_outputs(287);
    layer1_outputs(1430) <= not(layer0_outputs(1118));
    layer1_outputs(1431) <= not(layer0_outputs(4647));
    layer1_outputs(1432) <= '0';
    layer1_outputs(1433) <= (layer0_outputs(7404)) and not (layer0_outputs(3534));
    layer1_outputs(1434) <= (layer0_outputs(3518)) or (layer0_outputs(3915));
    layer1_outputs(1435) <= not(layer0_outputs(6788)) or (layer0_outputs(274));
    layer1_outputs(1436) <= not(layer0_outputs(211));
    layer1_outputs(1437) <= not((layer0_outputs(929)) or (layer0_outputs(5557)));
    layer1_outputs(1438) <= layer0_outputs(843);
    layer1_outputs(1439) <= not(layer0_outputs(5811));
    layer1_outputs(1440) <= '0';
    layer1_outputs(1441) <= not(layer0_outputs(1903)) or (layer0_outputs(3445));
    layer1_outputs(1442) <= not(layer0_outputs(2892));
    layer1_outputs(1443) <= not(layer0_outputs(5114));
    layer1_outputs(1444) <= not(layer0_outputs(396));
    layer1_outputs(1445) <= (layer0_outputs(1511)) xor (layer0_outputs(4735));
    layer1_outputs(1446) <= layer0_outputs(1512);
    layer1_outputs(1447) <= layer0_outputs(2325);
    layer1_outputs(1448) <= not(layer0_outputs(4882));
    layer1_outputs(1449) <= '0';
    layer1_outputs(1450) <= (layer0_outputs(329)) and not (layer0_outputs(2454));
    layer1_outputs(1451) <= not(layer0_outputs(3808)) or (layer0_outputs(2800));
    layer1_outputs(1452) <= '0';
    layer1_outputs(1453) <= (layer0_outputs(555)) and not (layer0_outputs(5054));
    layer1_outputs(1454) <= not(layer0_outputs(69));
    layer1_outputs(1455) <= not((layer0_outputs(3602)) or (layer0_outputs(4980)));
    layer1_outputs(1456) <= '0';
    layer1_outputs(1457) <= '1';
    layer1_outputs(1458) <= '0';
    layer1_outputs(1459) <= (layer0_outputs(5428)) and not (layer0_outputs(2292));
    layer1_outputs(1460) <= layer0_outputs(7490);
    layer1_outputs(1461) <= (layer0_outputs(7360)) and (layer0_outputs(2779));
    layer1_outputs(1462) <= not((layer0_outputs(916)) and (layer0_outputs(2696)));
    layer1_outputs(1463) <= (layer0_outputs(1010)) and not (layer0_outputs(4472));
    layer1_outputs(1464) <= not(layer0_outputs(3393));
    layer1_outputs(1465) <= not((layer0_outputs(620)) or (layer0_outputs(5459)));
    layer1_outputs(1466) <= (layer0_outputs(6108)) and (layer0_outputs(4638));
    layer1_outputs(1467) <= not(layer0_outputs(6938)) or (layer0_outputs(2753));
    layer1_outputs(1468) <= not((layer0_outputs(7002)) and (layer0_outputs(1000)));
    layer1_outputs(1469) <= layer0_outputs(7375);
    layer1_outputs(1470) <= not(layer0_outputs(2718));
    layer1_outputs(1471) <= not(layer0_outputs(2081));
    layer1_outputs(1472) <= not(layer0_outputs(6921));
    layer1_outputs(1473) <= layer0_outputs(1098);
    layer1_outputs(1474) <= '1';
    layer1_outputs(1475) <= (layer0_outputs(5523)) or (layer0_outputs(162));
    layer1_outputs(1476) <= (layer0_outputs(5373)) and not (layer0_outputs(1));
    layer1_outputs(1477) <= not(layer0_outputs(7450));
    layer1_outputs(1478) <= not(layer0_outputs(7620)) or (layer0_outputs(944));
    layer1_outputs(1479) <= not(layer0_outputs(6092)) or (layer0_outputs(4814));
    layer1_outputs(1480) <= (layer0_outputs(7186)) or (layer0_outputs(1319));
    layer1_outputs(1481) <= not(layer0_outputs(4000)) or (layer0_outputs(2472));
    layer1_outputs(1482) <= not(layer0_outputs(4619));
    layer1_outputs(1483) <= not((layer0_outputs(5306)) and (layer0_outputs(5131)));
    layer1_outputs(1484) <= (layer0_outputs(976)) and not (layer0_outputs(6358));
    layer1_outputs(1485) <= not(layer0_outputs(2512));
    layer1_outputs(1486) <= not(layer0_outputs(7388));
    layer1_outputs(1487) <= not((layer0_outputs(5658)) and (layer0_outputs(5413)));
    layer1_outputs(1488) <= not((layer0_outputs(2240)) or (layer0_outputs(157)));
    layer1_outputs(1489) <= not((layer0_outputs(4468)) and (layer0_outputs(415)));
    layer1_outputs(1490) <= (layer0_outputs(6789)) or (layer0_outputs(5943));
    layer1_outputs(1491) <= (layer0_outputs(3887)) and not (layer0_outputs(2932));
    layer1_outputs(1492) <= (layer0_outputs(5688)) and (layer0_outputs(4191));
    layer1_outputs(1493) <= layer0_outputs(4628);
    layer1_outputs(1494) <= layer0_outputs(986);
    layer1_outputs(1495) <= not(layer0_outputs(7551));
    layer1_outputs(1496) <= not((layer0_outputs(1679)) and (layer0_outputs(7227)));
    layer1_outputs(1497) <= '0';
    layer1_outputs(1498) <= not(layer0_outputs(4335)) or (layer0_outputs(1433));
    layer1_outputs(1499) <= (layer0_outputs(6975)) or (layer0_outputs(521));
    layer1_outputs(1500) <= '0';
    layer1_outputs(1501) <= not(layer0_outputs(2818));
    layer1_outputs(1502) <= '1';
    layer1_outputs(1503) <= (layer0_outputs(4532)) and not (layer0_outputs(972));
    layer1_outputs(1504) <= not(layer0_outputs(7540));
    layer1_outputs(1505) <= not((layer0_outputs(716)) and (layer0_outputs(656)));
    layer1_outputs(1506) <= not(layer0_outputs(7586)) or (layer0_outputs(5756));
    layer1_outputs(1507) <= (layer0_outputs(2249)) or (layer0_outputs(7301));
    layer1_outputs(1508) <= not((layer0_outputs(5729)) and (layer0_outputs(7502)));
    layer1_outputs(1509) <= '1';
    layer1_outputs(1510) <= (layer0_outputs(3199)) and not (layer0_outputs(2515));
    layer1_outputs(1511) <= not((layer0_outputs(7119)) and (layer0_outputs(4022)));
    layer1_outputs(1512) <= not((layer0_outputs(6443)) or (layer0_outputs(7524)));
    layer1_outputs(1513) <= not(layer0_outputs(687)) or (layer0_outputs(6541));
    layer1_outputs(1514) <= '0';
    layer1_outputs(1515) <= layer0_outputs(7621);
    layer1_outputs(1516) <= not(layer0_outputs(5080));
    layer1_outputs(1517) <= not(layer0_outputs(3843)) or (layer0_outputs(298));
    layer1_outputs(1518) <= '0';
    layer1_outputs(1519) <= (layer0_outputs(3137)) and (layer0_outputs(1216));
    layer1_outputs(1520) <= not(layer0_outputs(1231));
    layer1_outputs(1521) <= not(layer0_outputs(6948));
    layer1_outputs(1522) <= '0';
    layer1_outputs(1523) <= (layer0_outputs(3980)) and not (layer0_outputs(3863));
    layer1_outputs(1524) <= layer0_outputs(1236);
    layer1_outputs(1525) <= (layer0_outputs(4927)) and not (layer0_outputs(6423));
    layer1_outputs(1526) <= (layer0_outputs(3755)) and not (layer0_outputs(3866));
    layer1_outputs(1527) <= not((layer0_outputs(2364)) or (layer0_outputs(6778)));
    layer1_outputs(1528) <= not(layer0_outputs(1278)) or (layer0_outputs(889));
    layer1_outputs(1529) <= layer0_outputs(5746);
    layer1_outputs(1530) <= not((layer0_outputs(1612)) and (layer0_outputs(2226)));
    layer1_outputs(1531) <= not((layer0_outputs(3900)) and (layer0_outputs(6440)));
    layer1_outputs(1532) <= not(layer0_outputs(6245));
    layer1_outputs(1533) <= not(layer0_outputs(5158));
    layer1_outputs(1534) <= not(layer0_outputs(7077));
    layer1_outputs(1535) <= (layer0_outputs(1691)) xor (layer0_outputs(3333));
    layer1_outputs(1536) <= not(layer0_outputs(5728)) or (layer0_outputs(1938));
    layer1_outputs(1537) <= '1';
    layer1_outputs(1538) <= not((layer0_outputs(1880)) xor (layer0_outputs(494)));
    layer1_outputs(1539) <= not(layer0_outputs(6565));
    layer1_outputs(1540) <= layer0_outputs(1186);
    layer1_outputs(1541) <= not((layer0_outputs(5831)) and (layer0_outputs(1785)));
    layer1_outputs(1542) <= not(layer0_outputs(5012));
    layer1_outputs(1543) <= not((layer0_outputs(4355)) xor (layer0_outputs(7223)));
    layer1_outputs(1544) <= not((layer0_outputs(649)) or (layer0_outputs(3693)));
    layer1_outputs(1545) <= '1';
    layer1_outputs(1546) <= layer0_outputs(5812);
    layer1_outputs(1547) <= (layer0_outputs(7573)) and not (layer0_outputs(1783));
    layer1_outputs(1548) <= not(layer0_outputs(3116));
    layer1_outputs(1549) <= (layer0_outputs(3157)) and not (layer0_outputs(3491));
    layer1_outputs(1550) <= (layer0_outputs(7404)) or (layer0_outputs(4912));
    layer1_outputs(1551) <= (layer0_outputs(3818)) and not (layer0_outputs(2316));
    layer1_outputs(1552) <= layer0_outputs(7611);
    layer1_outputs(1553) <= '1';
    layer1_outputs(1554) <= not(layer0_outputs(3156));
    layer1_outputs(1555) <= not(layer0_outputs(154));
    layer1_outputs(1556) <= not(layer0_outputs(1893));
    layer1_outputs(1557) <= not((layer0_outputs(7199)) and (layer0_outputs(7355)));
    layer1_outputs(1558) <= (layer0_outputs(4981)) or (layer0_outputs(6216));
    layer1_outputs(1559) <= not(layer0_outputs(3458));
    layer1_outputs(1560) <= (layer0_outputs(1115)) and not (layer0_outputs(1065));
    layer1_outputs(1561) <= not(layer0_outputs(72)) or (layer0_outputs(7056));
    layer1_outputs(1562) <= not((layer0_outputs(3906)) and (layer0_outputs(3332)));
    layer1_outputs(1563) <= (layer0_outputs(5475)) and (layer0_outputs(4516));
    layer1_outputs(1564) <= not(layer0_outputs(727)) or (layer0_outputs(4536));
    layer1_outputs(1565) <= not(layer0_outputs(1227));
    layer1_outputs(1566) <= (layer0_outputs(2176)) or (layer0_outputs(7525));
    layer1_outputs(1567) <= not((layer0_outputs(4327)) or (layer0_outputs(265)));
    layer1_outputs(1568) <= not(layer0_outputs(4769)) or (layer0_outputs(5110));
    layer1_outputs(1569) <= not(layer0_outputs(391));
    layer1_outputs(1570) <= (layer0_outputs(5106)) and not (layer0_outputs(1577));
    layer1_outputs(1571) <= layer0_outputs(2055);
    layer1_outputs(1572) <= (layer0_outputs(7619)) and not (layer0_outputs(5481));
    layer1_outputs(1573) <= not(layer0_outputs(4012));
    layer1_outputs(1574) <= '1';
    layer1_outputs(1575) <= (layer0_outputs(6052)) and not (layer0_outputs(2377));
    layer1_outputs(1576) <= '1';
    layer1_outputs(1577) <= (layer0_outputs(3501)) and not (layer0_outputs(6834));
    layer1_outputs(1578) <= '1';
    layer1_outputs(1579) <= not(layer0_outputs(2721)) or (layer0_outputs(4886));
    layer1_outputs(1580) <= not((layer0_outputs(5621)) and (layer0_outputs(2544)));
    layer1_outputs(1581) <= (layer0_outputs(222)) or (layer0_outputs(3587));
    layer1_outputs(1582) <= (layer0_outputs(2036)) or (layer0_outputs(2579));
    layer1_outputs(1583) <= not((layer0_outputs(3901)) or (layer0_outputs(1898)));
    layer1_outputs(1584) <= layer0_outputs(6306);
    layer1_outputs(1585) <= not(layer0_outputs(3389)) or (layer0_outputs(2399));
    layer1_outputs(1586) <= (layer0_outputs(6365)) and not (layer0_outputs(5724));
    layer1_outputs(1587) <= '0';
    layer1_outputs(1588) <= not(layer0_outputs(2575));
    layer1_outputs(1589) <= (layer0_outputs(3053)) xor (layer0_outputs(4995));
    layer1_outputs(1590) <= layer0_outputs(3967);
    layer1_outputs(1591) <= '0';
    layer1_outputs(1592) <= (layer0_outputs(7346)) and (layer0_outputs(2520));
    layer1_outputs(1593) <= layer0_outputs(4218);
    layer1_outputs(1594) <= not(layer0_outputs(7130)) or (layer0_outputs(811));
    layer1_outputs(1595) <= layer0_outputs(7123);
    layer1_outputs(1596) <= '0';
    layer1_outputs(1597) <= not((layer0_outputs(2471)) and (layer0_outputs(2154)));
    layer1_outputs(1598) <= '0';
    layer1_outputs(1599) <= not((layer0_outputs(1551)) or (layer0_outputs(4720)));
    layer1_outputs(1600) <= not(layer0_outputs(6272));
    layer1_outputs(1601) <= not((layer0_outputs(1310)) and (layer0_outputs(1706)));
    layer1_outputs(1602) <= (layer0_outputs(982)) or (layer0_outputs(1643));
    layer1_outputs(1603) <= (layer0_outputs(1850)) and not (layer0_outputs(117));
    layer1_outputs(1604) <= not((layer0_outputs(3084)) xor (layer0_outputs(5754)));
    layer1_outputs(1605) <= not(layer0_outputs(7608));
    layer1_outputs(1606) <= layer0_outputs(1503);
    layer1_outputs(1607) <= layer0_outputs(1525);
    layer1_outputs(1608) <= layer0_outputs(5159);
    layer1_outputs(1609) <= not((layer0_outputs(5966)) and (layer0_outputs(404)));
    layer1_outputs(1610) <= not(layer0_outputs(3369));
    layer1_outputs(1611) <= '1';
    layer1_outputs(1612) <= not(layer0_outputs(6686)) or (layer0_outputs(7473));
    layer1_outputs(1613) <= not(layer0_outputs(3161)) or (layer0_outputs(4993));
    layer1_outputs(1614) <= (layer0_outputs(1712)) or (layer0_outputs(6710));
    layer1_outputs(1615) <= not((layer0_outputs(4773)) or (layer0_outputs(2706)));
    layer1_outputs(1616) <= not((layer0_outputs(13)) or (layer0_outputs(3352)));
    layer1_outputs(1617) <= (layer0_outputs(3443)) and not (layer0_outputs(2675));
    layer1_outputs(1618) <= (layer0_outputs(741)) or (layer0_outputs(6517));
    layer1_outputs(1619) <= (layer0_outputs(2213)) and not (layer0_outputs(6030));
    layer1_outputs(1620) <= not(layer0_outputs(4357)) or (layer0_outputs(864));
    layer1_outputs(1621) <= not(layer0_outputs(3758)) or (layer0_outputs(2115));
    layer1_outputs(1622) <= not(layer0_outputs(3564)) or (layer0_outputs(2042));
    layer1_outputs(1623) <= (layer0_outputs(1237)) and (layer0_outputs(5714));
    layer1_outputs(1624) <= (layer0_outputs(2546)) and (layer0_outputs(3166));
    layer1_outputs(1625) <= not(layer0_outputs(4511)) or (layer0_outputs(4485));
    layer1_outputs(1626) <= not((layer0_outputs(2028)) or (layer0_outputs(2828)));
    layer1_outputs(1627) <= not(layer0_outputs(1941));
    layer1_outputs(1628) <= not(layer0_outputs(932));
    layer1_outputs(1629) <= layer0_outputs(2088);
    layer1_outputs(1630) <= not(layer0_outputs(5465)) or (layer0_outputs(5295));
    layer1_outputs(1631) <= (layer0_outputs(5072)) xor (layer0_outputs(3657));
    layer1_outputs(1632) <= layer0_outputs(6431);
    layer1_outputs(1633) <= (layer0_outputs(214)) or (layer0_outputs(3401));
    layer1_outputs(1634) <= '1';
    layer1_outputs(1635) <= not(layer0_outputs(6852));
    layer1_outputs(1636) <= not((layer0_outputs(1778)) or (layer0_outputs(6897)));
    layer1_outputs(1637) <= not((layer0_outputs(6010)) or (layer0_outputs(1733)));
    layer1_outputs(1638) <= not((layer0_outputs(7383)) or (layer0_outputs(3979)));
    layer1_outputs(1639) <= not(layer0_outputs(7277));
    layer1_outputs(1640) <= not(layer0_outputs(882));
    layer1_outputs(1641) <= '1';
    layer1_outputs(1642) <= '0';
    layer1_outputs(1643) <= not(layer0_outputs(7478));
    layer1_outputs(1644) <= '0';
    layer1_outputs(1645) <= (layer0_outputs(3420)) or (layer0_outputs(6716));
    layer1_outputs(1646) <= not(layer0_outputs(7313)) or (layer0_outputs(1417));
    layer1_outputs(1647) <= (layer0_outputs(2135)) and not (layer0_outputs(474));
    layer1_outputs(1648) <= (layer0_outputs(1128)) and (layer0_outputs(6615));
    layer1_outputs(1649) <= not((layer0_outputs(2021)) or (layer0_outputs(3532)));
    layer1_outputs(1650) <= not(layer0_outputs(1550));
    layer1_outputs(1651) <= not(layer0_outputs(4208));
    layer1_outputs(1652) <= (layer0_outputs(1047)) and (layer0_outputs(5399));
    layer1_outputs(1653) <= '0';
    layer1_outputs(1654) <= layer0_outputs(7254);
    layer1_outputs(1655) <= (layer0_outputs(1348)) and (layer0_outputs(251));
    layer1_outputs(1656) <= (layer0_outputs(6826)) and not (layer0_outputs(1404));
    layer1_outputs(1657) <= '0';
    layer1_outputs(1658) <= not(layer0_outputs(483));
    layer1_outputs(1659) <= not(layer0_outputs(3470));
    layer1_outputs(1660) <= not(layer0_outputs(5051)) or (layer0_outputs(4176));
    layer1_outputs(1661) <= (layer0_outputs(395)) xor (layer0_outputs(99));
    layer1_outputs(1662) <= not((layer0_outputs(4531)) or (layer0_outputs(3312)));
    layer1_outputs(1663) <= layer0_outputs(1947);
    layer1_outputs(1664) <= layer0_outputs(6660);
    layer1_outputs(1665) <= not(layer0_outputs(709)) or (layer0_outputs(4095));
    layer1_outputs(1666) <= (layer0_outputs(4611)) and not (layer0_outputs(4076));
    layer1_outputs(1667) <= '0';
    layer1_outputs(1668) <= not(layer0_outputs(370));
    layer1_outputs(1669) <= (layer0_outputs(20)) and not (layer0_outputs(6646));
    layer1_outputs(1670) <= not((layer0_outputs(538)) and (layer0_outputs(7471)));
    layer1_outputs(1671) <= '0';
    layer1_outputs(1672) <= '1';
    layer1_outputs(1673) <= not(layer0_outputs(77)) or (layer0_outputs(6636));
    layer1_outputs(1674) <= not((layer0_outputs(5690)) or (layer0_outputs(5195)));
    layer1_outputs(1675) <= layer0_outputs(1309);
    layer1_outputs(1676) <= layer0_outputs(7424);
    layer1_outputs(1677) <= (layer0_outputs(6827)) and (layer0_outputs(6057));
    layer1_outputs(1678) <= not(layer0_outputs(6492));
    layer1_outputs(1679) <= not((layer0_outputs(7356)) and (layer0_outputs(5965)));
    layer1_outputs(1680) <= (layer0_outputs(942)) and (layer0_outputs(6521));
    layer1_outputs(1681) <= (layer0_outputs(5530)) and not (layer0_outputs(3258));
    layer1_outputs(1682) <= not(layer0_outputs(4802)) or (layer0_outputs(7287));
    layer1_outputs(1683) <= not((layer0_outputs(2791)) and (layer0_outputs(5193)));
    layer1_outputs(1684) <= not(layer0_outputs(1337));
    layer1_outputs(1685) <= not((layer0_outputs(2541)) or (layer0_outputs(6727)));
    layer1_outputs(1686) <= '0';
    layer1_outputs(1687) <= not(layer0_outputs(6004));
    layer1_outputs(1688) <= '0';
    layer1_outputs(1689) <= (layer0_outputs(3603)) or (layer0_outputs(5832));
    layer1_outputs(1690) <= not(layer0_outputs(2889)) or (layer0_outputs(3334));
    layer1_outputs(1691) <= not((layer0_outputs(4616)) or (layer0_outputs(352)));
    layer1_outputs(1692) <= (layer0_outputs(4673)) and not (layer0_outputs(5423));
    layer1_outputs(1693) <= (layer0_outputs(4546)) and (layer0_outputs(7195));
    layer1_outputs(1694) <= (layer0_outputs(5254)) and (layer0_outputs(2157));
    layer1_outputs(1695) <= not(layer0_outputs(2675));
    layer1_outputs(1696) <= layer0_outputs(2911);
    layer1_outputs(1697) <= (layer0_outputs(390)) and not (layer0_outputs(337));
    layer1_outputs(1698) <= layer0_outputs(1456);
    layer1_outputs(1699) <= (layer0_outputs(6555)) or (layer0_outputs(1418));
    layer1_outputs(1700) <= (layer0_outputs(5857)) and not (layer0_outputs(723));
    layer1_outputs(1701) <= '0';
    layer1_outputs(1702) <= (layer0_outputs(5989)) xor (layer0_outputs(4039));
    layer1_outputs(1703) <= '0';
    layer1_outputs(1704) <= not(layer0_outputs(3875));
    layer1_outputs(1705) <= not(layer0_outputs(3442)) or (layer0_outputs(7265));
    layer1_outputs(1706) <= '0';
    layer1_outputs(1707) <= (layer0_outputs(3557)) and not (layer0_outputs(6733));
    layer1_outputs(1708) <= not((layer0_outputs(2997)) or (layer0_outputs(5093)));
    layer1_outputs(1709) <= '0';
    layer1_outputs(1710) <= (layer0_outputs(3502)) and (layer0_outputs(4023));
    layer1_outputs(1711) <= (layer0_outputs(6330)) or (layer0_outputs(7063));
    layer1_outputs(1712) <= not(layer0_outputs(499)) or (layer0_outputs(6760));
    layer1_outputs(1713) <= not((layer0_outputs(4412)) xor (layer0_outputs(5544)));
    layer1_outputs(1714) <= layer0_outputs(1028);
    layer1_outputs(1715) <= (layer0_outputs(5149)) and (layer0_outputs(1247));
    layer1_outputs(1716) <= layer0_outputs(1135);
    layer1_outputs(1717) <= not(layer0_outputs(5346)) or (layer0_outputs(746));
    layer1_outputs(1718) <= (layer0_outputs(2739)) and not (layer0_outputs(2433));
    layer1_outputs(1719) <= not(layer0_outputs(4553));
    layer1_outputs(1720) <= not((layer0_outputs(1049)) or (layer0_outputs(7176)));
    layer1_outputs(1721) <= '1';
    layer1_outputs(1722) <= layer0_outputs(4329);
    layer1_outputs(1723) <= not((layer0_outputs(5187)) or (layer0_outputs(7568)));
    layer1_outputs(1724) <= not((layer0_outputs(6666)) or (layer0_outputs(3728)));
    layer1_outputs(1725) <= '1';
    layer1_outputs(1726) <= not((layer0_outputs(5304)) and (layer0_outputs(3043)));
    layer1_outputs(1727) <= not(layer0_outputs(2469));
    layer1_outputs(1728) <= not(layer0_outputs(1737)) or (layer0_outputs(5916));
    layer1_outputs(1729) <= (layer0_outputs(6643)) and (layer0_outputs(5520));
    layer1_outputs(1730) <= (layer0_outputs(275)) and not (layer0_outputs(6015));
    layer1_outputs(1731) <= not(layer0_outputs(2239));
    layer1_outputs(1732) <= '1';
    layer1_outputs(1733) <= (layer0_outputs(3877)) and (layer0_outputs(3404));
    layer1_outputs(1734) <= not(layer0_outputs(627)) or (layer0_outputs(4729));
    layer1_outputs(1735) <= '0';
    layer1_outputs(1736) <= not((layer0_outputs(3261)) or (layer0_outputs(5342)));
    layer1_outputs(1737) <= '1';
    layer1_outputs(1738) <= layer0_outputs(1346);
    layer1_outputs(1739) <= not((layer0_outputs(4926)) and (layer0_outputs(978)));
    layer1_outputs(1740) <= (layer0_outputs(723)) and not (layer0_outputs(3092));
    layer1_outputs(1741) <= not((layer0_outputs(6053)) or (layer0_outputs(1480)));
    layer1_outputs(1742) <= not(layer0_outputs(1574));
    layer1_outputs(1743) <= (layer0_outputs(3437)) and not (layer0_outputs(6227));
    layer1_outputs(1744) <= '0';
    layer1_outputs(1745) <= '0';
    layer1_outputs(1746) <= not((layer0_outputs(2004)) or (layer0_outputs(6730)));
    layer1_outputs(1747) <= (layer0_outputs(1340)) and (layer0_outputs(3316));
    layer1_outputs(1748) <= layer0_outputs(1588);
    layer1_outputs(1749) <= layer0_outputs(2199);
    layer1_outputs(1750) <= not(layer0_outputs(2875)) or (layer0_outputs(2122));
    layer1_outputs(1751) <= layer0_outputs(5150);
    layer1_outputs(1752) <= layer0_outputs(4284);
    layer1_outputs(1753) <= layer0_outputs(6645);
    layer1_outputs(1754) <= '1';
    layer1_outputs(1755) <= not((layer0_outputs(2136)) and (layer0_outputs(3825)));
    layer1_outputs(1756) <= '0';
    layer1_outputs(1757) <= '1';
    layer1_outputs(1758) <= '1';
    layer1_outputs(1759) <= '0';
    layer1_outputs(1760) <= (layer0_outputs(4791)) and not (layer0_outputs(5511));
    layer1_outputs(1761) <= (layer0_outputs(5850)) and not (layer0_outputs(7057));
    layer1_outputs(1762) <= not(layer0_outputs(6842));
    layer1_outputs(1763) <= '0';
    layer1_outputs(1764) <= (layer0_outputs(6330)) and not (layer0_outputs(1946));
    layer1_outputs(1765) <= (layer0_outputs(1792)) and (layer0_outputs(3372));
    layer1_outputs(1766) <= not((layer0_outputs(2374)) or (layer0_outputs(3722)));
    layer1_outputs(1767) <= (layer0_outputs(4034)) and not (layer0_outputs(7654));
    layer1_outputs(1768) <= not((layer0_outputs(3330)) or (layer0_outputs(2070)));
    layer1_outputs(1769) <= '0';
    layer1_outputs(1770) <= layer0_outputs(3458);
    layer1_outputs(1771) <= not(layer0_outputs(5028));
    layer1_outputs(1772) <= '0';
    layer1_outputs(1773) <= (layer0_outputs(3436)) and not (layer0_outputs(2664));
    layer1_outputs(1774) <= (layer0_outputs(7088)) or (layer0_outputs(5816));
    layer1_outputs(1775) <= (layer0_outputs(2439)) and not (layer0_outputs(3034));
    layer1_outputs(1776) <= not(layer0_outputs(1021)) or (layer0_outputs(4031));
    layer1_outputs(1777) <= '0';
    layer1_outputs(1778) <= layer0_outputs(4041);
    layer1_outputs(1779) <= '1';
    layer1_outputs(1780) <= (layer0_outputs(6114)) and not (layer0_outputs(3712));
    layer1_outputs(1781) <= '0';
    layer1_outputs(1782) <= '1';
    layer1_outputs(1783) <= not((layer0_outputs(6989)) xor (layer0_outputs(3901)));
    layer1_outputs(1784) <= (layer0_outputs(5884)) and (layer0_outputs(5410));
    layer1_outputs(1785) <= '1';
    layer1_outputs(1786) <= '1';
    layer1_outputs(1787) <= (layer0_outputs(2538)) or (layer0_outputs(2891));
    layer1_outputs(1788) <= '1';
    layer1_outputs(1789) <= not(layer0_outputs(1416)) or (layer0_outputs(6886));
    layer1_outputs(1790) <= '0';
    layer1_outputs(1791) <= (layer0_outputs(2237)) and not (layer0_outputs(388));
    layer1_outputs(1792) <= (layer0_outputs(5639)) and not (layer0_outputs(1326));
    layer1_outputs(1793) <= not((layer0_outputs(3970)) and (layer0_outputs(7609)));
    layer1_outputs(1794) <= not(layer0_outputs(1630));
    layer1_outputs(1795) <= not(layer0_outputs(5228));
    layer1_outputs(1796) <= (layer0_outputs(5321)) and not (layer0_outputs(2456));
    layer1_outputs(1797) <= layer0_outputs(116);
    layer1_outputs(1798) <= '1';
    layer1_outputs(1799) <= layer0_outputs(2760);
    layer1_outputs(1800) <= (layer0_outputs(2100)) and not (layer0_outputs(5152));
    layer1_outputs(1801) <= not(layer0_outputs(4474));
    layer1_outputs(1802) <= not(layer0_outputs(2931)) or (layer0_outputs(1109));
    layer1_outputs(1803) <= layer0_outputs(6341);
    layer1_outputs(1804) <= not((layer0_outputs(6562)) xor (layer0_outputs(7055)));
    layer1_outputs(1805) <= not(layer0_outputs(6236)) or (layer0_outputs(3792));
    layer1_outputs(1806) <= not((layer0_outputs(7541)) and (layer0_outputs(6115)));
    layer1_outputs(1807) <= not(layer0_outputs(6813));
    layer1_outputs(1808) <= not(layer0_outputs(5273)) or (layer0_outputs(5451));
    layer1_outputs(1809) <= (layer0_outputs(6839)) or (layer0_outputs(3162));
    layer1_outputs(1810) <= (layer0_outputs(1384)) and (layer0_outputs(1531));
    layer1_outputs(1811) <= layer0_outputs(3310);
    layer1_outputs(1812) <= (layer0_outputs(605)) and (layer0_outputs(147));
    layer1_outputs(1813) <= (layer0_outputs(3473)) and (layer0_outputs(524));
    layer1_outputs(1814) <= (layer0_outputs(2119)) or (layer0_outputs(672));
    layer1_outputs(1815) <= not(layer0_outputs(423));
    layer1_outputs(1816) <= (layer0_outputs(4070)) and not (layer0_outputs(2052));
    layer1_outputs(1817) <= '0';
    layer1_outputs(1818) <= layer0_outputs(4918);
    layer1_outputs(1819) <= (layer0_outputs(5538)) and (layer0_outputs(4060));
    layer1_outputs(1820) <= '0';
    layer1_outputs(1821) <= not(layer0_outputs(6456));
    layer1_outputs(1822) <= (layer0_outputs(700)) and not (layer0_outputs(7571));
    layer1_outputs(1823) <= (layer0_outputs(4124)) and (layer0_outputs(2709));
    layer1_outputs(1824) <= not(layer0_outputs(6572));
    layer1_outputs(1825) <= layer0_outputs(193);
    layer1_outputs(1826) <= not((layer0_outputs(182)) and (layer0_outputs(3584)));
    layer1_outputs(1827) <= not(layer0_outputs(3405)) or (layer0_outputs(178));
    layer1_outputs(1828) <= layer0_outputs(1452);
    layer1_outputs(1829) <= (layer0_outputs(5702)) and not (layer0_outputs(3645));
    layer1_outputs(1830) <= not((layer0_outputs(4820)) or (layer0_outputs(41)));
    layer1_outputs(1831) <= layer0_outputs(1443);
    layer1_outputs(1832) <= not((layer0_outputs(5225)) and (layer0_outputs(7552)));
    layer1_outputs(1833) <= not((layer0_outputs(5796)) and (layer0_outputs(5548)));
    layer1_outputs(1834) <= layer0_outputs(2341);
    layer1_outputs(1835) <= not(layer0_outputs(7067));
    layer1_outputs(1836) <= not(layer0_outputs(2313));
    layer1_outputs(1837) <= (layer0_outputs(7416)) and (layer0_outputs(3861));
    layer1_outputs(1838) <= (layer0_outputs(2539)) and (layer0_outputs(6785));
    layer1_outputs(1839) <= not(layer0_outputs(2756)) or (layer0_outputs(2607));
    layer1_outputs(1840) <= not((layer0_outputs(5923)) and (layer0_outputs(283)));
    layer1_outputs(1841) <= not(layer0_outputs(4996));
    layer1_outputs(1842) <= not(layer0_outputs(5698));
    layer1_outputs(1843) <= not(layer0_outputs(6156));
    layer1_outputs(1844) <= not((layer0_outputs(1005)) or (layer0_outputs(6305)));
    layer1_outputs(1845) <= layer0_outputs(2290);
    layer1_outputs(1846) <= (layer0_outputs(5046)) xor (layer0_outputs(338));
    layer1_outputs(1847) <= '0';
    layer1_outputs(1848) <= (layer0_outputs(6553)) and not (layer0_outputs(6695));
    layer1_outputs(1849) <= not(layer0_outputs(7669));
    layer1_outputs(1850) <= not(layer0_outputs(4972));
    layer1_outputs(1851) <= layer0_outputs(6343);
    layer1_outputs(1852) <= (layer0_outputs(3)) or (layer0_outputs(5081));
    layer1_outputs(1853) <= layer0_outputs(2693);
    layer1_outputs(1854) <= not(layer0_outputs(968)) or (layer0_outputs(7387));
    layer1_outputs(1855) <= not((layer0_outputs(4475)) and (layer0_outputs(167)));
    layer1_outputs(1856) <= layer0_outputs(3257);
    layer1_outputs(1857) <= (layer0_outputs(7242)) or (layer0_outputs(7180));
    layer1_outputs(1858) <= not((layer0_outputs(4697)) and (layer0_outputs(1734)));
    layer1_outputs(1859) <= '0';
    layer1_outputs(1860) <= '1';
    layer1_outputs(1861) <= (layer0_outputs(3743)) or (layer0_outputs(547));
    layer1_outputs(1862) <= not(layer0_outputs(6266)) or (layer0_outputs(5731));
    layer1_outputs(1863) <= not(layer0_outputs(260));
    layer1_outputs(1864) <= not(layer0_outputs(233));
    layer1_outputs(1865) <= '1';
    layer1_outputs(1866) <= not((layer0_outputs(5503)) or (layer0_outputs(1798)));
    layer1_outputs(1867) <= (layer0_outputs(832)) and not (layer0_outputs(3665));
    layer1_outputs(1868) <= '1';
    layer1_outputs(1869) <= layer0_outputs(912);
    layer1_outputs(1870) <= '1';
    layer1_outputs(1871) <= '0';
    layer1_outputs(1872) <= layer0_outputs(2112);
    layer1_outputs(1873) <= not(layer0_outputs(4165)) or (layer0_outputs(1554));
    layer1_outputs(1874) <= '1';
    layer1_outputs(1875) <= layer0_outputs(776);
    layer1_outputs(1876) <= (layer0_outputs(91)) and not (layer0_outputs(685));
    layer1_outputs(1877) <= (layer0_outputs(4962)) and not (layer0_outputs(3727));
    layer1_outputs(1878) <= (layer0_outputs(6468)) and not (layer0_outputs(6668));
    layer1_outputs(1879) <= layer0_outputs(1757);
    layer1_outputs(1880) <= layer0_outputs(2069);
    layer1_outputs(1881) <= layer0_outputs(5516);
    layer1_outputs(1882) <= not(layer0_outputs(1750));
    layer1_outputs(1883) <= not(layer0_outputs(1987));
    layer1_outputs(1884) <= (layer0_outputs(447)) xor (layer0_outputs(5915));
    layer1_outputs(1885) <= (layer0_outputs(4744)) and not (layer0_outputs(6125));
    layer1_outputs(1886) <= layer0_outputs(4033);
    layer1_outputs(1887) <= '0';
    layer1_outputs(1888) <= (layer0_outputs(6157)) and not (layer0_outputs(4404));
    layer1_outputs(1889) <= layer0_outputs(4647);
    layer1_outputs(1890) <= not(layer0_outputs(7167)) or (layer0_outputs(5942));
    layer1_outputs(1891) <= not((layer0_outputs(4222)) or (layer0_outputs(6267)));
    layer1_outputs(1892) <= (layer0_outputs(3690)) and not (layer0_outputs(6735));
    layer1_outputs(1893) <= not(layer0_outputs(541));
    layer1_outputs(1894) <= '1';
    layer1_outputs(1895) <= '0';
    layer1_outputs(1896) <= layer0_outputs(2118);
    layer1_outputs(1897) <= layer0_outputs(2692);
    layer1_outputs(1898) <= '0';
    layer1_outputs(1899) <= (layer0_outputs(3744)) or (layer0_outputs(2962));
    layer1_outputs(1900) <= not(layer0_outputs(7679));
    layer1_outputs(1901) <= not((layer0_outputs(5085)) xor (layer0_outputs(4238)));
    layer1_outputs(1902) <= not(layer0_outputs(4556));
    layer1_outputs(1903) <= (layer0_outputs(3418)) and not (layer0_outputs(3596));
    layer1_outputs(1904) <= '0';
    layer1_outputs(1905) <= layer0_outputs(855);
    layer1_outputs(1906) <= '1';
    layer1_outputs(1907) <= '0';
    layer1_outputs(1908) <= not((layer0_outputs(2164)) xor (layer0_outputs(446)));
    layer1_outputs(1909) <= not(layer0_outputs(4870));
    layer1_outputs(1910) <= not((layer0_outputs(4526)) or (layer0_outputs(675)));
    layer1_outputs(1911) <= layer0_outputs(2185);
    layer1_outputs(1912) <= layer0_outputs(7180);
    layer1_outputs(1913) <= (layer0_outputs(6024)) and not (layer0_outputs(3383));
    layer1_outputs(1914) <= (layer0_outputs(6275)) and (layer0_outputs(3767));
    layer1_outputs(1915) <= (layer0_outputs(4735)) and (layer0_outputs(1619));
    layer1_outputs(1916) <= not((layer0_outputs(703)) and (layer0_outputs(2259)));
    layer1_outputs(1917) <= not(layer0_outputs(6463));
    layer1_outputs(1918) <= not((layer0_outputs(1457)) and (layer0_outputs(7120)));
    layer1_outputs(1919) <= (layer0_outputs(6697)) and (layer0_outputs(2570));
    layer1_outputs(1920) <= '1';
    layer1_outputs(1921) <= '0';
    layer1_outputs(1922) <= not(layer0_outputs(3444)) or (layer0_outputs(2357));
    layer1_outputs(1923) <= '0';
    layer1_outputs(1924) <= '0';
    layer1_outputs(1925) <= (layer0_outputs(920)) and (layer0_outputs(5645));
    layer1_outputs(1926) <= (layer0_outputs(4423)) and not (layer0_outputs(4921));
    layer1_outputs(1927) <= (layer0_outputs(6070)) or (layer0_outputs(1036));
    layer1_outputs(1928) <= layer0_outputs(4183);
    layer1_outputs(1929) <= not(layer0_outputs(2847));
    layer1_outputs(1930) <= (layer0_outputs(2798)) and not (layer0_outputs(3072));
    layer1_outputs(1931) <= not(layer0_outputs(4390)) or (layer0_outputs(2893));
    layer1_outputs(1932) <= (layer0_outputs(5207)) and not (layer0_outputs(2557));
    layer1_outputs(1933) <= '1';
    layer1_outputs(1934) <= layer0_outputs(390);
    layer1_outputs(1935) <= (layer0_outputs(3775)) xor (layer0_outputs(2281));
    layer1_outputs(1936) <= layer0_outputs(1292);
    layer1_outputs(1937) <= not((layer0_outputs(3321)) or (layer0_outputs(6061)));
    layer1_outputs(1938) <= '1';
    layer1_outputs(1939) <= not((layer0_outputs(7434)) xor (layer0_outputs(6195)));
    layer1_outputs(1940) <= not(layer0_outputs(1253));
    layer1_outputs(1941) <= not(layer0_outputs(5426));
    layer1_outputs(1942) <= not(layer0_outputs(7603)) or (layer0_outputs(5018));
    layer1_outputs(1943) <= (layer0_outputs(6259)) or (layer0_outputs(4645));
    layer1_outputs(1944) <= '1';
    layer1_outputs(1945) <= (layer0_outputs(6151)) and not (layer0_outputs(7563));
    layer1_outputs(1946) <= not((layer0_outputs(6939)) or (layer0_outputs(1013)));
    layer1_outputs(1947) <= not(layer0_outputs(2750)) or (layer0_outputs(5563));
    layer1_outputs(1948) <= layer0_outputs(6713);
    layer1_outputs(1949) <= '1';
    layer1_outputs(1950) <= not(layer0_outputs(4119));
    layer1_outputs(1951) <= (layer0_outputs(3475)) and not (layer0_outputs(5486));
    layer1_outputs(1952) <= (layer0_outputs(6826)) and not (layer0_outputs(7018));
    layer1_outputs(1953) <= layer0_outputs(2188);
    layer1_outputs(1954) <= not(layer0_outputs(1859)) or (layer0_outputs(4416));
    layer1_outputs(1955) <= not((layer0_outputs(2883)) or (layer0_outputs(6322)));
    layer1_outputs(1956) <= not(layer0_outputs(5502));
    layer1_outputs(1957) <= not((layer0_outputs(7129)) or (layer0_outputs(2822)));
    layer1_outputs(1958) <= '0';
    layer1_outputs(1959) <= not(layer0_outputs(3893)) or (layer0_outputs(6559));
    layer1_outputs(1960) <= '0';
    layer1_outputs(1961) <= (layer0_outputs(3234)) or (layer0_outputs(5953));
    layer1_outputs(1962) <= '0';
    layer1_outputs(1963) <= not(layer0_outputs(2793)) or (layer0_outputs(5776));
    layer1_outputs(1964) <= not(layer0_outputs(2187));
    layer1_outputs(1965) <= not(layer0_outputs(4849));
    layer1_outputs(1966) <= layer0_outputs(2427);
    layer1_outputs(1967) <= (layer0_outputs(1250)) and (layer0_outputs(4219));
    layer1_outputs(1968) <= not(layer0_outputs(2450)) or (layer0_outputs(2052));
    layer1_outputs(1969) <= layer0_outputs(5490);
    layer1_outputs(1970) <= not(layer0_outputs(543));
    layer1_outputs(1971) <= (layer0_outputs(3202)) or (layer0_outputs(2210));
    layer1_outputs(1972) <= layer0_outputs(2114);
    layer1_outputs(1973) <= '1';
    layer1_outputs(1974) <= (layer0_outputs(4200)) and not (layer0_outputs(3994));
    layer1_outputs(1975) <= '0';
    layer1_outputs(1976) <= '0';
    layer1_outputs(1977) <= '0';
    layer1_outputs(1978) <= layer0_outputs(6367);
    layer1_outputs(1979) <= (layer0_outputs(4794)) and not (layer0_outputs(2810));
    layer1_outputs(1980) <= not(layer0_outputs(5978)) or (layer0_outputs(7228));
    layer1_outputs(1981) <= layer0_outputs(7033);
    layer1_outputs(1982) <= not(layer0_outputs(1029)) or (layer0_outputs(4753));
    layer1_outputs(1983) <= (layer0_outputs(985)) or (layer0_outputs(2310));
    layer1_outputs(1984) <= '1';
    layer1_outputs(1985) <= '1';
    layer1_outputs(1986) <= '0';
    layer1_outputs(1987) <= layer0_outputs(3753);
    layer1_outputs(1988) <= not(layer0_outputs(7251)) or (layer0_outputs(5670));
    layer1_outputs(1989) <= (layer0_outputs(4245)) or (layer0_outputs(7073));
    layer1_outputs(1990) <= '0';
    layer1_outputs(1991) <= (layer0_outputs(4233)) and (layer0_outputs(2892));
    layer1_outputs(1992) <= layer0_outputs(1163);
    layer1_outputs(1993) <= not(layer0_outputs(5985));
    layer1_outputs(1994) <= (layer0_outputs(4853)) and not (layer0_outputs(1618));
    layer1_outputs(1995) <= not(layer0_outputs(1208));
    layer1_outputs(1996) <= not(layer0_outputs(5019));
    layer1_outputs(1997) <= not(layer0_outputs(3988));
    layer1_outputs(1998) <= not(layer0_outputs(3966)) or (layer0_outputs(1441));
    layer1_outputs(1999) <= not(layer0_outputs(105));
    layer1_outputs(2000) <= not(layer0_outputs(6824)) or (layer0_outputs(3544));
    layer1_outputs(2001) <= not((layer0_outputs(124)) and (layer0_outputs(5651)));
    layer1_outputs(2002) <= (layer0_outputs(2747)) xor (layer0_outputs(7202));
    layer1_outputs(2003) <= '0';
    layer1_outputs(2004) <= not(layer0_outputs(2137)) or (layer0_outputs(6883));
    layer1_outputs(2005) <= '1';
    layer1_outputs(2006) <= (layer0_outputs(6955)) or (layer0_outputs(3325));
    layer1_outputs(2007) <= not((layer0_outputs(4793)) or (layer0_outputs(2120)));
    layer1_outputs(2008) <= (layer0_outputs(1225)) and (layer0_outputs(5996));
    layer1_outputs(2009) <= not((layer0_outputs(4145)) and (layer0_outputs(733)));
    layer1_outputs(2010) <= not((layer0_outputs(4957)) or (layer0_outputs(4114)));
    layer1_outputs(2011) <= not(layer0_outputs(4879)) or (layer0_outputs(234));
    layer1_outputs(2012) <= (layer0_outputs(7583)) and (layer0_outputs(1493));
    layer1_outputs(2013) <= not(layer0_outputs(1189));
    layer1_outputs(2014) <= layer0_outputs(4319);
    layer1_outputs(2015) <= not(layer0_outputs(2378)) or (layer0_outputs(2201));
    layer1_outputs(2016) <= '1';
    layer1_outputs(2017) <= layer0_outputs(4915);
    layer1_outputs(2018) <= (layer0_outputs(7176)) and not (layer0_outputs(5560));
    layer1_outputs(2019) <= layer0_outputs(634);
    layer1_outputs(2020) <= layer0_outputs(4176);
    layer1_outputs(2021) <= not(layer0_outputs(2163));
    layer1_outputs(2022) <= (layer0_outputs(48)) and not (layer0_outputs(790));
    layer1_outputs(2023) <= not(layer0_outputs(4687)) or (layer0_outputs(3598));
    layer1_outputs(2024) <= (layer0_outputs(4635)) or (layer0_outputs(4251));
    layer1_outputs(2025) <= (layer0_outputs(3635)) or (layer0_outputs(4138));
    layer1_outputs(2026) <= not(layer0_outputs(4033)) or (layer0_outputs(7218));
    layer1_outputs(2027) <= not(layer0_outputs(1657));
    layer1_outputs(2028) <= '1';
    layer1_outputs(2029) <= not(layer0_outputs(5276));
    layer1_outputs(2030) <= '0';
    layer1_outputs(2031) <= (layer0_outputs(5049)) or (layer0_outputs(6221));
    layer1_outputs(2032) <= not(layer0_outputs(694)) or (layer0_outputs(1957));
    layer1_outputs(2033) <= '1';
    layer1_outputs(2034) <= '0';
    layer1_outputs(2035) <= not(layer0_outputs(7419));
    layer1_outputs(2036) <= '1';
    layer1_outputs(2037) <= not(layer0_outputs(7652));
    layer1_outputs(2038) <= '1';
    layer1_outputs(2039) <= '0';
    layer1_outputs(2040) <= layer0_outputs(4424);
    layer1_outputs(2041) <= (layer0_outputs(4959)) and (layer0_outputs(184));
    layer1_outputs(2042) <= '0';
    layer1_outputs(2043) <= layer0_outputs(5178);
    layer1_outputs(2044) <= (layer0_outputs(5422)) xor (layer0_outputs(4225));
    layer1_outputs(2045) <= (layer0_outputs(3567)) and not (layer0_outputs(198));
    layer1_outputs(2046) <= not((layer0_outputs(4480)) and (layer0_outputs(7652)));
    layer1_outputs(2047) <= (layer0_outputs(6233)) and not (layer0_outputs(5887));
    layer1_outputs(2048) <= not(layer0_outputs(1012));
    layer1_outputs(2049) <= not((layer0_outputs(6950)) and (layer0_outputs(1440)));
    layer1_outputs(2050) <= not((layer0_outputs(6832)) or (layer0_outputs(2683)));
    layer1_outputs(2051) <= not(layer0_outputs(3095)) or (layer0_outputs(7046));
    layer1_outputs(2052) <= not(layer0_outputs(7401));
    layer1_outputs(2053) <= (layer0_outputs(4514)) or (layer0_outputs(2245));
    layer1_outputs(2054) <= not(layer0_outputs(5313));
    layer1_outputs(2055) <= not(layer0_outputs(475));
    layer1_outputs(2056) <= '1';
    layer1_outputs(2057) <= not((layer0_outputs(5421)) and (layer0_outputs(4553)));
    layer1_outputs(2058) <= (layer0_outputs(1245)) and not (layer0_outputs(6863));
    layer1_outputs(2059) <= (layer0_outputs(4857)) or (layer0_outputs(2579));
    layer1_outputs(2060) <= layer0_outputs(3476);
    layer1_outputs(2061) <= not((layer0_outputs(6587)) and (layer0_outputs(7662)));
    layer1_outputs(2062) <= (layer0_outputs(7086)) or (layer0_outputs(3400));
    layer1_outputs(2063) <= layer0_outputs(7442);
    layer1_outputs(2064) <= not((layer0_outputs(532)) and (layer0_outputs(2758)));
    layer1_outputs(2065) <= not(layer0_outputs(2414));
    layer1_outputs(2066) <= not(layer0_outputs(2375)) or (layer0_outputs(6362));
    layer1_outputs(2067) <= not(layer0_outputs(3991));
    layer1_outputs(2068) <= (layer0_outputs(4978)) and (layer0_outputs(5883));
    layer1_outputs(2069) <= not(layer0_outputs(6188)) or (layer0_outputs(5833));
    layer1_outputs(2070) <= '0';
    layer1_outputs(2071) <= not(layer0_outputs(2365));
    layer1_outputs(2072) <= (layer0_outputs(1203)) or (layer0_outputs(6629));
    layer1_outputs(2073) <= '0';
    layer1_outputs(2074) <= not((layer0_outputs(3221)) or (layer0_outputs(1046)));
    layer1_outputs(2075) <= not((layer0_outputs(2151)) and (layer0_outputs(2002)));
    layer1_outputs(2076) <= (layer0_outputs(1789)) or (layer0_outputs(6801));
    layer1_outputs(2077) <= not((layer0_outputs(7634)) or (layer0_outputs(420)));
    layer1_outputs(2078) <= (layer0_outputs(4762)) and not (layer0_outputs(3103));
    layer1_outputs(2079) <= not(layer0_outputs(1747));
    layer1_outputs(2080) <= not(layer0_outputs(4567));
    layer1_outputs(2081) <= not(layer0_outputs(6033));
    layer1_outputs(2082) <= '0';
    layer1_outputs(2083) <= (layer0_outputs(4666)) and (layer0_outputs(3033));
    layer1_outputs(2084) <= not(layer0_outputs(6737));
    layer1_outputs(2085) <= not(layer0_outputs(2344));
    layer1_outputs(2086) <= (layer0_outputs(4179)) xor (layer0_outputs(168));
    layer1_outputs(2087) <= layer0_outputs(7106);
    layer1_outputs(2088) <= '1';
    layer1_outputs(2089) <= not(layer0_outputs(1261));
    layer1_outputs(2090) <= not((layer0_outputs(1061)) or (layer0_outputs(4539)));
    layer1_outputs(2091) <= not(layer0_outputs(3574));
    layer1_outputs(2092) <= not(layer0_outputs(3486)) or (layer0_outputs(4456));
    layer1_outputs(2093) <= (layer0_outputs(6577)) xor (layer0_outputs(2324));
    layer1_outputs(2094) <= not(layer0_outputs(3811));
    layer1_outputs(2095) <= (layer0_outputs(1196)) and (layer0_outputs(10));
    layer1_outputs(2096) <= layer0_outputs(6587);
    layer1_outputs(2097) <= not(layer0_outputs(3535));
    layer1_outputs(2098) <= not(layer0_outputs(5116)) or (layer0_outputs(4334));
    layer1_outputs(2099) <= not((layer0_outputs(454)) xor (layer0_outputs(121)));
    layer1_outputs(2100) <= not((layer0_outputs(4913)) and (layer0_outputs(3731)));
    layer1_outputs(2101) <= (layer0_outputs(5695)) and (layer0_outputs(1800));
    layer1_outputs(2102) <= not(layer0_outputs(2685));
    layer1_outputs(2103) <= not((layer0_outputs(3665)) and (layer0_outputs(6231)));
    layer1_outputs(2104) <= '1';
    layer1_outputs(2105) <= not((layer0_outputs(7570)) or (layer0_outputs(6096)));
    layer1_outputs(2106) <= layer0_outputs(6262);
    layer1_outputs(2107) <= (layer0_outputs(7509)) and (layer0_outputs(5707));
    layer1_outputs(2108) <= not(layer0_outputs(500));
    layer1_outputs(2109) <= layer0_outputs(5655);
    layer1_outputs(2110) <= (layer0_outputs(4181)) and not (layer0_outputs(1206));
    layer1_outputs(2111) <= (layer0_outputs(2411)) and not (layer0_outputs(5526));
    layer1_outputs(2112) <= '1';
    layer1_outputs(2113) <= (layer0_outputs(3477)) and (layer0_outputs(3076));
    layer1_outputs(2114) <= '0';
    layer1_outputs(2115) <= '1';
    layer1_outputs(2116) <= not((layer0_outputs(2495)) and (layer0_outputs(4287)));
    layer1_outputs(2117) <= (layer0_outputs(2335)) and (layer0_outputs(891));
    layer1_outputs(2118) <= not(layer0_outputs(6254));
    layer1_outputs(2119) <= layer0_outputs(6648);
    layer1_outputs(2120) <= layer0_outputs(2677);
    layer1_outputs(2121) <= not(layer0_outputs(7667)) or (layer0_outputs(1045));
    layer1_outputs(2122) <= not(layer0_outputs(3942)) or (layer0_outputs(4236));
    layer1_outputs(2123) <= (layer0_outputs(4665)) and (layer0_outputs(6334));
    layer1_outputs(2124) <= (layer0_outputs(2759)) and not (layer0_outputs(4334));
    layer1_outputs(2125) <= not(layer0_outputs(1439)) or (layer0_outputs(3895));
    layer1_outputs(2126) <= (layer0_outputs(6122)) and not (layer0_outputs(7442));
    layer1_outputs(2127) <= not(layer0_outputs(6687));
    layer1_outputs(2128) <= not(layer0_outputs(7300)) or (layer0_outputs(3333));
    layer1_outputs(2129) <= (layer0_outputs(6047)) and not (layer0_outputs(201));
    layer1_outputs(2130) <= not((layer0_outputs(1544)) and (layer0_outputs(4613)));
    layer1_outputs(2131) <= not(layer0_outputs(3799)) or (layer0_outputs(7059));
    layer1_outputs(2132) <= (layer0_outputs(1817)) and not (layer0_outputs(6389));
    layer1_outputs(2133) <= (layer0_outputs(7396)) or (layer0_outputs(1468));
    layer1_outputs(2134) <= layer0_outputs(5164);
    layer1_outputs(2135) <= '0';
    layer1_outputs(2136) <= not(layer0_outputs(6500));
    layer1_outputs(2137) <= not(layer0_outputs(487)) or (layer0_outputs(4396));
    layer1_outputs(2138) <= '0';
    layer1_outputs(2139) <= (layer0_outputs(4523)) and not (layer0_outputs(6453));
    layer1_outputs(2140) <= not(layer0_outputs(4084)) or (layer0_outputs(4795));
    layer1_outputs(2141) <= not((layer0_outputs(4139)) or (layer0_outputs(6783)));
    layer1_outputs(2142) <= (layer0_outputs(5027)) and (layer0_outputs(6012));
    layer1_outputs(2143) <= layer0_outputs(1902);
    layer1_outputs(2144) <= not((layer0_outputs(2944)) and (layer0_outputs(3230)));
    layer1_outputs(2145) <= not(layer0_outputs(3188)) or (layer0_outputs(2108));
    layer1_outputs(2146) <= not((layer0_outputs(1899)) or (layer0_outputs(838)));
    layer1_outputs(2147) <= (layer0_outputs(3847)) and (layer0_outputs(5196));
    layer1_outputs(2148) <= layer0_outputs(4780);
    layer1_outputs(2149) <= layer0_outputs(134);
    layer1_outputs(2150) <= (layer0_outputs(6923)) and not (layer0_outputs(98));
    layer1_outputs(2151) <= not(layer0_outputs(3925)) or (layer0_outputs(2727));
    layer1_outputs(2152) <= (layer0_outputs(343)) or (layer0_outputs(3559));
    layer1_outputs(2153) <= (layer0_outputs(4427)) or (layer0_outputs(5781));
    layer1_outputs(2154) <= '1';
    layer1_outputs(2155) <= not((layer0_outputs(2698)) or (layer0_outputs(251)));
    layer1_outputs(2156) <= not((layer0_outputs(4378)) and (layer0_outputs(4571)));
    layer1_outputs(2157) <= not(layer0_outputs(2077));
    layer1_outputs(2158) <= not(layer0_outputs(7250));
    layer1_outputs(2159) <= '1';
    layer1_outputs(2160) <= not(layer0_outputs(49));
    layer1_outputs(2161) <= not(layer0_outputs(1197));
    layer1_outputs(2162) <= (layer0_outputs(6528)) and not (layer0_outputs(296));
    layer1_outputs(2163) <= (layer0_outputs(2416)) or (layer0_outputs(5910));
    layer1_outputs(2164) <= not(layer0_outputs(2341)) or (layer0_outputs(2272));
    layer1_outputs(2165) <= '0';
    layer1_outputs(2166) <= not(layer0_outputs(4001)) or (layer0_outputs(4192));
    layer1_outputs(2167) <= not((layer0_outputs(4178)) and (layer0_outputs(1651)));
    layer1_outputs(2168) <= layer0_outputs(1268);
    layer1_outputs(2169) <= not(layer0_outputs(1742));
    layer1_outputs(2170) <= layer0_outputs(2204);
    layer1_outputs(2171) <= not((layer0_outputs(3920)) and (layer0_outputs(838)));
    layer1_outputs(2172) <= not(layer0_outputs(6582));
    layer1_outputs(2173) <= '0';
    layer1_outputs(2174) <= not((layer0_outputs(3534)) and (layer0_outputs(1205)));
    layer1_outputs(2175) <= not((layer0_outputs(5204)) or (layer0_outputs(1346)));
    layer1_outputs(2176) <= (layer0_outputs(5145)) and not (layer0_outputs(783));
    layer1_outputs(2177) <= not(layer0_outputs(311));
    layer1_outputs(2178) <= layer0_outputs(277);
    layer1_outputs(2179) <= not(layer0_outputs(5039)) or (layer0_outputs(12));
    layer1_outputs(2180) <= not(layer0_outputs(4227)) or (layer0_outputs(3457));
    layer1_outputs(2181) <= not(layer0_outputs(6734)) or (layer0_outputs(2740));
    layer1_outputs(2182) <= (layer0_outputs(2922)) xor (layer0_outputs(1253));
    layer1_outputs(2183) <= layer0_outputs(1422);
    layer1_outputs(2184) <= not((layer0_outputs(5792)) and (layer0_outputs(2311)));
    layer1_outputs(2185) <= not((layer0_outputs(3537)) and (layer0_outputs(3188)));
    layer1_outputs(2186) <= not(layer0_outputs(3429));
    layer1_outputs(2187) <= layer0_outputs(451);
    layer1_outputs(2188) <= (layer0_outputs(5016)) and (layer0_outputs(5758));
    layer1_outputs(2189) <= (layer0_outputs(766)) and (layer0_outputs(3867));
    layer1_outputs(2190) <= (layer0_outputs(1168)) and not (layer0_outputs(6543));
    layer1_outputs(2191) <= not(layer0_outputs(3198)) or (layer0_outputs(1172));
    layer1_outputs(2192) <= '0';
    layer1_outputs(2193) <= not(layer0_outputs(3956));
    layer1_outputs(2194) <= (layer0_outputs(571)) and (layer0_outputs(4855));
    layer1_outputs(2195) <= '0';
    layer1_outputs(2196) <= not((layer0_outputs(1453)) and (layer0_outputs(4391)));
    layer1_outputs(2197) <= not((layer0_outputs(4088)) and (layer0_outputs(2371)));
    layer1_outputs(2198) <= (layer0_outputs(2487)) or (layer0_outputs(5248));
    layer1_outputs(2199) <= not(layer0_outputs(5905));
    layer1_outputs(2200) <= not(layer0_outputs(6629)) or (layer0_outputs(3254));
    layer1_outputs(2201) <= (layer0_outputs(4458)) xor (layer0_outputs(258));
    layer1_outputs(2202) <= not(layer0_outputs(210)) or (layer0_outputs(1718));
    layer1_outputs(2203) <= '1';
    layer1_outputs(2204) <= not((layer0_outputs(2253)) and (layer0_outputs(3439)));
    layer1_outputs(2205) <= layer0_outputs(6887);
    layer1_outputs(2206) <= (layer0_outputs(5336)) and not (layer0_outputs(3010));
    layer1_outputs(2207) <= layer0_outputs(1508);
    layer1_outputs(2208) <= not(layer0_outputs(5984));
    layer1_outputs(2209) <= (layer0_outputs(2939)) and not (layer0_outputs(1315));
    layer1_outputs(2210) <= not(layer0_outputs(5433));
    layer1_outputs(2211) <= (layer0_outputs(6051)) or (layer0_outputs(6558));
    layer1_outputs(2212) <= layer0_outputs(5279);
    layer1_outputs(2213) <= not((layer0_outputs(4435)) and (layer0_outputs(1372)));
    layer1_outputs(2214) <= not(layer0_outputs(1604)) or (layer0_outputs(1667));
    layer1_outputs(2215) <= (layer0_outputs(7008)) and not (layer0_outputs(7661));
    layer1_outputs(2216) <= layer0_outputs(560);
    layer1_outputs(2217) <= layer0_outputs(1581);
    layer1_outputs(2218) <= '1';
    layer1_outputs(2219) <= not((layer0_outputs(7262)) and (layer0_outputs(780)));
    layer1_outputs(2220) <= not(layer0_outputs(2432));
    layer1_outputs(2221) <= '1';
    layer1_outputs(2222) <= (layer0_outputs(2713)) or (layer0_outputs(7507));
    layer1_outputs(2223) <= not(layer0_outputs(2979));
    layer1_outputs(2224) <= '0';
    layer1_outputs(2225) <= not((layer0_outputs(690)) or (layer0_outputs(829)));
    layer1_outputs(2226) <= (layer0_outputs(1939)) or (layer0_outputs(4008));
    layer1_outputs(2227) <= (layer0_outputs(678)) and not (layer0_outputs(6269));
    layer1_outputs(2228) <= not(layer0_outputs(5093));
    layer1_outputs(2229) <= '1';
    layer1_outputs(2230) <= '0';
    layer1_outputs(2231) <= not(layer0_outputs(4771));
    layer1_outputs(2232) <= not(layer0_outputs(4013)) or (layer0_outputs(523));
    layer1_outputs(2233) <= not((layer0_outputs(2110)) or (layer0_outputs(2687)));
    layer1_outputs(2234) <= layer0_outputs(1563);
    layer1_outputs(2235) <= not(layer0_outputs(527)) or (layer0_outputs(516));
    layer1_outputs(2236) <= not(layer0_outputs(6969));
    layer1_outputs(2237) <= layer0_outputs(5057);
    layer1_outputs(2238) <= layer0_outputs(1860);
    layer1_outputs(2239) <= not(layer0_outputs(7039)) or (layer0_outputs(6422));
    layer1_outputs(2240) <= not(layer0_outputs(1032)) or (layer0_outputs(6695));
    layer1_outputs(2241) <= not(layer0_outputs(7370)) or (layer0_outputs(6213));
    layer1_outputs(2242) <= '0';
    layer1_outputs(2243) <= (layer0_outputs(1863)) and not (layer0_outputs(4778));
    layer1_outputs(2244) <= layer0_outputs(7382);
    layer1_outputs(2245) <= (layer0_outputs(1633)) and not (layer0_outputs(644));
    layer1_outputs(2246) <= layer0_outputs(5436);
    layer1_outputs(2247) <= not(layer0_outputs(5687));
    layer1_outputs(2248) <= layer0_outputs(6277);
    layer1_outputs(2249) <= not((layer0_outputs(1647)) and (layer0_outputs(2155)));
    layer1_outputs(2250) <= not((layer0_outputs(7539)) and (layer0_outputs(100)));
    layer1_outputs(2251) <= '0';
    layer1_outputs(2252) <= '1';
    layer1_outputs(2253) <= not((layer0_outputs(1077)) or (layer0_outputs(2930)));
    layer1_outputs(2254) <= not(layer0_outputs(5096)) or (layer0_outputs(1331));
    layer1_outputs(2255) <= (layer0_outputs(1323)) or (layer0_outputs(1073));
    layer1_outputs(2256) <= layer0_outputs(1331);
    layer1_outputs(2257) <= '1';
    layer1_outputs(2258) <= layer0_outputs(4265);
    layer1_outputs(2259) <= not(layer0_outputs(4903));
    layer1_outputs(2260) <= layer0_outputs(2208);
    layer1_outputs(2261) <= not((layer0_outputs(3599)) xor (layer0_outputs(3660)));
    layer1_outputs(2262) <= layer0_outputs(4721);
    layer1_outputs(2263) <= '1';
    layer1_outputs(2264) <= not(layer0_outputs(4302));
    layer1_outputs(2265) <= (layer0_outputs(4908)) and (layer0_outputs(5630));
    layer1_outputs(2266) <= (layer0_outputs(5668)) and not (layer0_outputs(1398));
    layer1_outputs(2267) <= layer0_outputs(5244);
    layer1_outputs(2268) <= layer0_outputs(1460);
    layer1_outputs(2269) <= layer0_outputs(7106);
    layer1_outputs(2270) <= (layer0_outputs(98)) and (layer0_outputs(6704));
    layer1_outputs(2271) <= not((layer0_outputs(4730)) and (layer0_outputs(7129)));
    layer1_outputs(2272) <= (layer0_outputs(5679)) and not (layer0_outputs(6867));
    layer1_outputs(2273) <= not(layer0_outputs(7320));
    layer1_outputs(2274) <= (layer0_outputs(498)) and not (layer0_outputs(2357));
    layer1_outputs(2275) <= (layer0_outputs(2615)) and not (layer0_outputs(2711));
    layer1_outputs(2276) <= not(layer0_outputs(3828));
    layer1_outputs(2277) <= not((layer0_outputs(522)) xor (layer0_outputs(3500)));
    layer1_outputs(2278) <= '1';
    layer1_outputs(2279) <= '0';
    layer1_outputs(2280) <= '0';
    layer1_outputs(2281) <= not((layer0_outputs(2153)) and (layer0_outputs(3031)));
    layer1_outputs(2282) <= (layer0_outputs(2806)) and (layer0_outputs(2373));
    layer1_outputs(2283) <= (layer0_outputs(430)) and not (layer0_outputs(3407));
    layer1_outputs(2284) <= '0';
    layer1_outputs(2285) <= not((layer0_outputs(666)) or (layer0_outputs(4850)));
    layer1_outputs(2286) <= not((layer0_outputs(5947)) or (layer0_outputs(4682)));
    layer1_outputs(2287) <= '1';
    layer1_outputs(2288) <= (layer0_outputs(4525)) and not (layer0_outputs(6707));
    layer1_outputs(2289) <= '1';
    layer1_outputs(2290) <= (layer0_outputs(4260)) or (layer0_outputs(2877));
    layer1_outputs(2291) <= not((layer0_outputs(7122)) or (layer0_outputs(1159)));
    layer1_outputs(2292) <= not(layer0_outputs(1265));
    layer1_outputs(2293) <= (layer0_outputs(6597)) and not (layer0_outputs(2858));
    layer1_outputs(2294) <= '0';
    layer1_outputs(2295) <= not((layer0_outputs(1937)) or (layer0_outputs(6324)));
    layer1_outputs(2296) <= (layer0_outputs(332)) or (layer0_outputs(6960));
    layer1_outputs(2297) <= not(layer0_outputs(3216));
    layer1_outputs(2298) <= not(layer0_outputs(1590));
    layer1_outputs(2299) <= not(layer0_outputs(5214));
    layer1_outputs(2300) <= not(layer0_outputs(6805));
    layer1_outputs(2301) <= not(layer0_outputs(4828)) or (layer0_outputs(5495));
    layer1_outputs(2302) <= (layer0_outputs(3999)) and (layer0_outputs(3340));
    layer1_outputs(2303) <= not((layer0_outputs(2162)) and (layer0_outputs(857)));
    layer1_outputs(2304) <= layer0_outputs(3181);
    layer1_outputs(2305) <= not((layer0_outputs(4626)) or (layer0_outputs(453)));
    layer1_outputs(2306) <= not(layer0_outputs(1111));
    layer1_outputs(2307) <= '1';
    layer1_outputs(2308) <= (layer0_outputs(3381)) and (layer0_outputs(2837));
    layer1_outputs(2309) <= (layer0_outputs(408)) and not (layer0_outputs(4343));
    layer1_outputs(2310) <= not(layer0_outputs(1312));
    layer1_outputs(2311) <= (layer0_outputs(2797)) and not (layer0_outputs(3981));
    layer1_outputs(2312) <= not((layer0_outputs(171)) or (layer0_outputs(845)));
    layer1_outputs(2313) <= '1';
    layer1_outputs(2314) <= (layer0_outputs(4375)) or (layer0_outputs(5510));
    layer1_outputs(2315) <= '0';
    layer1_outputs(2316) <= layer0_outputs(6765);
    layer1_outputs(2317) <= '1';
    layer1_outputs(2318) <= not(layer0_outputs(5150));
    layer1_outputs(2319) <= not((layer0_outputs(2381)) and (layer0_outputs(662)));
    layer1_outputs(2320) <= '1';
    layer1_outputs(2321) <= not(layer0_outputs(4645)) or (layer0_outputs(5827));
    layer1_outputs(2322) <= layer0_outputs(6478);
    layer1_outputs(2323) <= (layer0_outputs(3421)) and not (layer0_outputs(3277));
    layer1_outputs(2324) <= not(layer0_outputs(7458));
    layer1_outputs(2325) <= (layer0_outputs(1169)) or (layer0_outputs(924));
    layer1_outputs(2326) <= (layer0_outputs(2805)) and not (layer0_outputs(7101));
    layer1_outputs(2327) <= (layer0_outputs(2360)) and (layer0_outputs(2774));
    layer1_outputs(2328) <= (layer0_outputs(6732)) and not (layer0_outputs(3765));
    layer1_outputs(2329) <= layer0_outputs(266);
    layer1_outputs(2330) <= layer0_outputs(4385);
    layer1_outputs(2331) <= (layer0_outputs(6075)) or (layer0_outputs(6530));
    layer1_outputs(2332) <= '1';
    layer1_outputs(2333) <= '0';
    layer1_outputs(2334) <= not((layer0_outputs(5457)) or (layer0_outputs(48)));
    layer1_outputs(2335) <= '0';
    layer1_outputs(2336) <= (layer0_outputs(5439)) and not (layer0_outputs(3466));
    layer1_outputs(2337) <= not((layer0_outputs(3876)) or (layer0_outputs(6940)));
    layer1_outputs(2338) <= (layer0_outputs(4102)) and (layer0_outputs(1671));
    layer1_outputs(2339) <= layer0_outputs(4659);
    layer1_outputs(2340) <= not(layer0_outputs(5453));
    layer1_outputs(2341) <= not(layer0_outputs(1744)) or (layer0_outputs(5684));
    layer1_outputs(2342) <= '1';
    layer1_outputs(2343) <= (layer0_outputs(163)) and not (layer0_outputs(6170));
    layer1_outputs(2344) <= (layer0_outputs(190)) and not (layer0_outputs(1522));
    layer1_outputs(2345) <= not(layer0_outputs(6934));
    layer1_outputs(2346) <= not((layer0_outputs(3980)) and (layer0_outputs(3392)));
    layer1_outputs(2347) <= not(layer0_outputs(7298)) or (layer0_outputs(5932));
    layer1_outputs(2348) <= not(layer0_outputs(1273));
    layer1_outputs(2349) <= not((layer0_outputs(2682)) or (layer0_outputs(5643)));
    layer1_outputs(2350) <= '1';
    layer1_outputs(2351) <= not((layer0_outputs(7042)) or (layer0_outputs(6451)));
    layer1_outputs(2352) <= layer0_outputs(1269);
    layer1_outputs(2353) <= (layer0_outputs(3610)) and (layer0_outputs(7569));
    layer1_outputs(2354) <= (layer0_outputs(6321)) or (layer0_outputs(6519));
    layer1_outputs(2355) <= (layer0_outputs(2628)) and not (layer0_outputs(1180));
    layer1_outputs(2356) <= not(layer0_outputs(4897)) or (layer0_outputs(5271));
    layer1_outputs(2357) <= not((layer0_outputs(616)) or (layer0_outputs(3476)));
    layer1_outputs(2358) <= layer0_outputs(197);
    layer1_outputs(2359) <= '0';
    layer1_outputs(2360) <= not(layer0_outputs(6692));
    layer1_outputs(2361) <= '1';
    layer1_outputs(2362) <= '1';
    layer1_outputs(2363) <= not(layer0_outputs(4863));
    layer1_outputs(2364) <= layer0_outputs(7072);
    layer1_outputs(2365) <= not(layer0_outputs(5188)) or (layer0_outputs(5989));
    layer1_outputs(2366) <= not(layer0_outputs(7672));
    layer1_outputs(2367) <= not(layer0_outputs(5314));
    layer1_outputs(2368) <= not((layer0_outputs(2644)) or (layer0_outputs(2338)));
    layer1_outputs(2369) <= (layer0_outputs(2046)) and not (layer0_outputs(2907));
    layer1_outputs(2370) <= '0';
    layer1_outputs(2371) <= layer0_outputs(7324);
    layer1_outputs(2372) <= not(layer0_outputs(2448)) or (layer0_outputs(5845));
    layer1_outputs(2373) <= (layer0_outputs(3760)) xor (layer0_outputs(6816));
    layer1_outputs(2374) <= not(layer0_outputs(5702)) or (layer0_outputs(2975));
    layer1_outputs(2375) <= '1';
    layer1_outputs(2376) <= (layer0_outputs(4441)) or (layer0_outputs(307));
    layer1_outputs(2377) <= not((layer0_outputs(1944)) and (layer0_outputs(2647)));
    layer1_outputs(2378) <= not((layer0_outputs(2174)) or (layer0_outputs(7254)));
    layer1_outputs(2379) <= not(layer0_outputs(4981));
    layer1_outputs(2380) <= not(layer0_outputs(3710));
    layer1_outputs(2381) <= not(layer0_outputs(6979));
    layer1_outputs(2382) <= '0';
    layer1_outputs(2383) <= not(layer0_outputs(749));
    layer1_outputs(2384) <= '0';
    layer1_outputs(2385) <= not((layer0_outputs(3590)) or (layer0_outputs(3467)));
    layer1_outputs(2386) <= layer0_outputs(6131);
    layer1_outputs(2387) <= '1';
    layer1_outputs(2388) <= not(layer0_outputs(2848)) or (layer0_outputs(96));
    layer1_outputs(2389) <= (layer0_outputs(4110)) and not (layer0_outputs(2827));
    layer1_outputs(2390) <= '0';
    layer1_outputs(2391) <= layer0_outputs(2828);
    layer1_outputs(2392) <= (layer0_outputs(1410)) xor (layer0_outputs(2740));
    layer1_outputs(2393) <= not((layer0_outputs(1824)) or (layer0_outputs(6827)));
    layer1_outputs(2394) <= (layer0_outputs(1387)) or (layer0_outputs(6988));
    layer1_outputs(2395) <= layer0_outputs(2243);
    layer1_outputs(2396) <= not(layer0_outputs(7216));
    layer1_outputs(2397) <= (layer0_outputs(5664)) or (layer0_outputs(2626));
    layer1_outputs(2398) <= '1';
    layer1_outputs(2399) <= not(layer0_outputs(6848)) or (layer0_outputs(4882));
    layer1_outputs(2400) <= layer0_outputs(5119);
    layer1_outputs(2401) <= not(layer0_outputs(819));
    layer1_outputs(2402) <= not(layer0_outputs(4576)) or (layer0_outputs(413));
    layer1_outputs(2403) <= not(layer0_outputs(4889)) or (layer0_outputs(4899));
    layer1_outputs(2404) <= (layer0_outputs(5333)) and not (layer0_outputs(4422));
    layer1_outputs(2405) <= (layer0_outputs(7556)) and not (layer0_outputs(2598));
    layer1_outputs(2406) <= layer0_outputs(2302);
    layer1_outputs(2407) <= '0';
    layer1_outputs(2408) <= (layer0_outputs(5728)) and not (layer0_outputs(3868));
    layer1_outputs(2409) <= layer0_outputs(2469);
    layer1_outputs(2410) <= (layer0_outputs(2482)) or (layer0_outputs(2130));
    layer1_outputs(2411) <= not((layer0_outputs(2417)) and (layer0_outputs(1883)));
    layer1_outputs(2412) <= not(layer0_outputs(7215)) or (layer0_outputs(3233));
    layer1_outputs(2413) <= not(layer0_outputs(7607));
    layer1_outputs(2414) <= '1';
    layer1_outputs(2415) <= (layer0_outputs(2424)) and not (layer0_outputs(5335));
    layer1_outputs(2416) <= (layer0_outputs(7025)) xor (layer0_outputs(6412));
    layer1_outputs(2417) <= '0';
    layer1_outputs(2418) <= layer0_outputs(5600);
    layer1_outputs(2419) <= not((layer0_outputs(4615)) or (layer0_outputs(4733)));
    layer1_outputs(2420) <= layer0_outputs(1277);
    layer1_outputs(2421) <= '0';
    layer1_outputs(2422) <= not((layer0_outputs(82)) and (layer0_outputs(3902)));
    layer1_outputs(2423) <= not(layer0_outputs(1347)) or (layer0_outputs(268));
    layer1_outputs(2424) <= layer0_outputs(3635);
    layer1_outputs(2425) <= (layer0_outputs(3219)) and not (layer0_outputs(2764));
    layer1_outputs(2426) <= layer0_outputs(3294);
    layer1_outputs(2427) <= not((layer0_outputs(141)) and (layer0_outputs(4409)));
    layer1_outputs(2428) <= '1';
    layer1_outputs(2429) <= (layer0_outputs(4430)) and not (layer0_outputs(3961));
    layer1_outputs(2430) <= not(layer0_outputs(1576)) or (layer0_outputs(1908));
    layer1_outputs(2431) <= '0';
    layer1_outputs(2432) <= not(layer0_outputs(3198)) or (layer0_outputs(1910));
    layer1_outputs(2433) <= not((layer0_outputs(7515)) or (layer0_outputs(912)));
    layer1_outputs(2434) <= (layer0_outputs(653)) and not (layer0_outputs(2015));
    layer1_outputs(2435) <= not((layer0_outputs(4182)) or (layer0_outputs(7003)));
    layer1_outputs(2436) <= not(layer0_outputs(2517)) or (layer0_outputs(1142));
    layer1_outputs(2437) <= not(layer0_outputs(2071));
    layer1_outputs(2438) <= '1';
    layer1_outputs(2439) <= '0';
    layer1_outputs(2440) <= not((layer0_outputs(3394)) and (layer0_outputs(5778)));
    layer1_outputs(2441) <= not(layer0_outputs(5083)) or (layer0_outputs(16));
    layer1_outputs(2442) <= layer0_outputs(4533);
    layer1_outputs(2443) <= layer0_outputs(519);
    layer1_outputs(2444) <= (layer0_outputs(5930)) and (layer0_outputs(6005));
    layer1_outputs(2445) <= layer0_outputs(6574);
    layer1_outputs(2446) <= (layer0_outputs(4633)) xor (layer0_outputs(2561));
    layer1_outputs(2447) <= layer0_outputs(7583);
    layer1_outputs(2448) <= not(layer0_outputs(1385)) or (layer0_outputs(3907));
    layer1_outputs(2449) <= '1';
    layer1_outputs(2450) <= layer0_outputs(4201);
    layer1_outputs(2451) <= layer0_outputs(4354);
    layer1_outputs(2452) <= (layer0_outputs(7626)) and not (layer0_outputs(4535));
    layer1_outputs(2453) <= (layer0_outputs(7310)) and not (layer0_outputs(6881));
    layer1_outputs(2454) <= '0';
    layer1_outputs(2455) <= not(layer0_outputs(905));
    layer1_outputs(2456) <= '1';
    layer1_outputs(2457) <= '1';
    layer1_outputs(2458) <= '0';
    layer1_outputs(2459) <= layer0_outputs(2231);
    layer1_outputs(2460) <= '0';
    layer1_outputs(2461) <= layer0_outputs(6074);
    layer1_outputs(2462) <= not((layer0_outputs(6178)) and (layer0_outputs(2989)));
    layer1_outputs(2463) <= (layer0_outputs(729)) and not (layer0_outputs(3209));
    layer1_outputs(2464) <= not(layer0_outputs(6946));
    layer1_outputs(2465) <= not(layer0_outputs(2167));
    layer1_outputs(2466) <= not(layer0_outputs(409)) or (layer0_outputs(7325));
    layer1_outputs(2467) <= layer0_outputs(480);
    layer1_outputs(2468) <= '1';
    layer1_outputs(2469) <= not(layer0_outputs(6095));
    layer1_outputs(2470) <= '1';
    layer1_outputs(2471) <= (layer0_outputs(6977)) or (layer0_outputs(360));
    layer1_outputs(2472) <= not(layer0_outputs(7265));
    layer1_outputs(2473) <= layer0_outputs(36);
    layer1_outputs(2474) <= (layer0_outputs(947)) and not (layer0_outputs(7648));
    layer1_outputs(2475) <= (layer0_outputs(3033)) and (layer0_outputs(5805));
    layer1_outputs(2476) <= (layer0_outputs(491)) and not (layer0_outputs(6117));
    layer1_outputs(2477) <= '1';
    layer1_outputs(2478) <= (layer0_outputs(7546)) and not (layer0_outputs(3153));
    layer1_outputs(2479) <= not((layer0_outputs(6673)) or (layer0_outputs(6420)));
    layer1_outputs(2480) <= not((layer0_outputs(3443)) or (layer0_outputs(3141)));
    layer1_outputs(2481) <= layer0_outputs(6628);
    layer1_outputs(2482) <= '1';
    layer1_outputs(2483) <= layer0_outputs(5680);
    layer1_outputs(2484) <= '1';
    layer1_outputs(2485) <= '1';
    layer1_outputs(2486) <= (layer0_outputs(2498)) or (layer0_outputs(6044));
    layer1_outputs(2487) <= not(layer0_outputs(5649));
    layer1_outputs(2488) <= not((layer0_outputs(4501)) or (layer0_outputs(847)));
    layer1_outputs(2489) <= (layer0_outputs(3331)) and not (layer0_outputs(1481));
    layer1_outputs(2490) <= (layer0_outputs(3781)) xor (layer0_outputs(4148));
    layer1_outputs(2491) <= '1';
    layer1_outputs(2492) <= not(layer0_outputs(6424)) or (layer0_outputs(467));
    layer1_outputs(2493) <= layer0_outputs(4524);
    layer1_outputs(2494) <= not((layer0_outputs(6071)) or (layer0_outputs(1099)));
    layer1_outputs(2495) <= not((layer0_outputs(1703)) or (layer0_outputs(159)));
    layer1_outputs(2496) <= not(layer0_outputs(6677)) or (layer0_outputs(5436));
    layer1_outputs(2497) <= (layer0_outputs(6240)) and not (layer0_outputs(2038));
    layer1_outputs(2498) <= (layer0_outputs(1869)) and not (layer0_outputs(6208));
    layer1_outputs(2499) <= layer0_outputs(975);
    layer1_outputs(2500) <= layer0_outputs(5194);
    layer1_outputs(2501) <= layer0_outputs(5703);
    layer1_outputs(2502) <= not(layer0_outputs(1945));
    layer1_outputs(2503) <= not(layer0_outputs(4747));
    layer1_outputs(2504) <= (layer0_outputs(4560)) and not (layer0_outputs(2165));
    layer1_outputs(2505) <= '0';
    layer1_outputs(2506) <= (layer0_outputs(4383)) and (layer0_outputs(1535));
    layer1_outputs(2507) <= (layer0_outputs(4990)) and not (layer0_outputs(540));
    layer1_outputs(2508) <= (layer0_outputs(4233)) xor (layer0_outputs(2873));
    layer1_outputs(2509) <= (layer0_outputs(6233)) and (layer0_outputs(5650));
    layer1_outputs(2510) <= not(layer0_outputs(1124)) or (layer0_outputs(221));
    layer1_outputs(2511) <= (layer0_outputs(6747)) and not (layer0_outputs(237));
    layer1_outputs(2512) <= not(layer0_outputs(5836));
    layer1_outputs(2513) <= (layer0_outputs(6940)) and not (layer0_outputs(6447));
    layer1_outputs(2514) <= not((layer0_outputs(5373)) xor (layer0_outputs(6737)));
    layer1_outputs(2515) <= not(layer0_outputs(5575));
    layer1_outputs(2516) <= (layer0_outputs(965)) and not (layer0_outputs(5147));
    layer1_outputs(2517) <= layer0_outputs(2057);
    layer1_outputs(2518) <= (layer0_outputs(7126)) or (layer0_outputs(3592));
    layer1_outputs(2519) <= '0';
    layer1_outputs(2520) <= not(layer0_outputs(4958)) or (layer0_outputs(5991));
    layer1_outputs(2521) <= '1';
    layer1_outputs(2522) <= (layer0_outputs(4462)) and (layer0_outputs(6598));
    layer1_outputs(2523) <= '1';
    layer1_outputs(2524) <= '0';
    layer1_outputs(2525) <= not(layer0_outputs(7387)) or (layer0_outputs(3038));
    layer1_outputs(2526) <= not((layer0_outputs(3087)) and (layer0_outputs(6403)));
    layer1_outputs(2527) <= not((layer0_outputs(7455)) xor (layer0_outputs(55)));
    layer1_outputs(2528) <= not(layer0_outputs(426)) or (layer0_outputs(2346));
    layer1_outputs(2529) <= not(layer0_outputs(5875)) or (layer0_outputs(2539));
    layer1_outputs(2530) <= (layer0_outputs(3821)) and (layer0_outputs(6457));
    layer1_outputs(2531) <= not(layer0_outputs(3155)) or (layer0_outputs(3359));
    layer1_outputs(2532) <= not(layer0_outputs(7007)) or (layer0_outputs(91));
    layer1_outputs(2533) <= not((layer0_outputs(2037)) xor (layer0_outputs(5386)));
    layer1_outputs(2534) <= not(layer0_outputs(4847));
    layer1_outputs(2535) <= (layer0_outputs(682)) and not (layer0_outputs(3683));
    layer1_outputs(2536) <= layer0_outputs(6705);
    layer1_outputs(2537) <= layer0_outputs(3156);
    layer1_outputs(2538) <= '0';
    layer1_outputs(2539) <= '1';
    layer1_outputs(2540) <= '0';
    layer1_outputs(2541) <= (layer0_outputs(487)) or (layer0_outputs(2));
    layer1_outputs(2542) <= not((layer0_outputs(186)) and (layer0_outputs(220)));
    layer1_outputs(2543) <= layer0_outputs(2682);
    layer1_outputs(2544) <= not(layer0_outputs(3636)) or (layer0_outputs(6705));
    layer1_outputs(2545) <= layer0_outputs(1413);
    layer1_outputs(2546) <= not(layer0_outputs(2549));
    layer1_outputs(2547) <= layer0_outputs(1063);
    layer1_outputs(2548) <= (layer0_outputs(4946)) and not (layer0_outputs(6945));
    layer1_outputs(2549) <= (layer0_outputs(1700)) or (layer0_outputs(4287));
    layer1_outputs(2550) <= '1';
    layer1_outputs(2551) <= (layer0_outputs(5183)) and not (layer0_outputs(6730));
    layer1_outputs(2552) <= layer0_outputs(6299);
    layer1_outputs(2553) <= not((layer0_outputs(4899)) and (layer0_outputs(1940)));
    layer1_outputs(2554) <= not(layer0_outputs(5667)) or (layer0_outputs(342));
    layer1_outputs(2555) <= layer0_outputs(4268);
    layer1_outputs(2556) <= '1';
    layer1_outputs(2557) <= (layer0_outputs(2401)) and not (layer0_outputs(7591));
    layer1_outputs(2558) <= not(layer0_outputs(7329));
    layer1_outputs(2559) <= not(layer0_outputs(534));
    layer1_outputs(2560) <= not(layer0_outputs(641)) or (layer0_outputs(324));
    layer1_outputs(2561) <= not((layer0_outputs(2156)) or (layer0_outputs(6139)));
    layer1_outputs(2562) <= layer0_outputs(4710);
    layer1_outputs(2563) <= not(layer0_outputs(2991));
    layer1_outputs(2564) <= not(layer0_outputs(885));
    layer1_outputs(2565) <= (layer0_outputs(5282)) or (layer0_outputs(3713));
    layer1_outputs(2566) <= not(layer0_outputs(2385));
    layer1_outputs(2567) <= layer0_outputs(542);
    layer1_outputs(2568) <= not(layer0_outputs(5312)) or (layer0_outputs(4614));
    layer1_outputs(2569) <= not(layer0_outputs(7475)) or (layer0_outputs(4437));
    layer1_outputs(2570) <= not((layer0_outputs(437)) or (layer0_outputs(1001)));
    layer1_outputs(2571) <= layer0_outputs(3918);
    layer1_outputs(2572) <= not((layer0_outputs(2523)) or (layer0_outputs(3670)));
    layer1_outputs(2573) <= not(layer0_outputs(6541)) or (layer0_outputs(328));
    layer1_outputs(2574) <= not((layer0_outputs(1761)) and (layer0_outputs(369)));
    layer1_outputs(2575) <= '1';
    layer1_outputs(2576) <= '0';
    layer1_outputs(2577) <= layer0_outputs(2801);
    layer1_outputs(2578) <= not((layer0_outputs(1594)) or (layer0_outputs(2783)));
    layer1_outputs(2579) <= (layer0_outputs(456)) or (layer0_outputs(6575));
    layer1_outputs(2580) <= (layer0_outputs(1893)) or (layer0_outputs(2809));
    layer1_outputs(2581) <= layer0_outputs(6297);
    layer1_outputs(2582) <= '0';
    layer1_outputs(2583) <= not((layer0_outputs(1670)) and (layer0_outputs(4755)));
    layer1_outputs(2584) <= layer0_outputs(1927);
    layer1_outputs(2585) <= not((layer0_outputs(4001)) and (layer0_outputs(7342)));
    layer1_outputs(2586) <= layer0_outputs(3510);
    layer1_outputs(2587) <= not((layer0_outputs(4113)) and (layer0_outputs(6218)));
    layer1_outputs(2588) <= not((layer0_outputs(2221)) and (layer0_outputs(1649)));
    layer1_outputs(2589) <= (layer0_outputs(4711)) and not (layer0_outputs(6128));
    layer1_outputs(2590) <= not(layer0_outputs(6703)) or (layer0_outputs(7500));
    layer1_outputs(2591) <= (layer0_outputs(5487)) and (layer0_outputs(1494));
    layer1_outputs(2592) <= not(layer0_outputs(1819)) or (layer0_outputs(5273));
    layer1_outputs(2593) <= '1';
    layer1_outputs(2594) <= not((layer0_outputs(6012)) and (layer0_outputs(3355)));
    layer1_outputs(2595) <= layer0_outputs(4726);
    layer1_outputs(2596) <= not(layer0_outputs(234)) or (layer0_outputs(1664));
    layer1_outputs(2597) <= layer0_outputs(4581);
    layer1_outputs(2598) <= not(layer0_outputs(2297)) or (layer0_outputs(54));
    layer1_outputs(2599) <= (layer0_outputs(5855)) and not (layer0_outputs(1240));
    layer1_outputs(2600) <= not(layer0_outputs(4062));
    layer1_outputs(2601) <= not((layer0_outputs(6449)) or (layer0_outputs(4996)));
    layer1_outputs(2602) <= '0';
    layer1_outputs(2603) <= (layer0_outputs(5363)) and not (layer0_outputs(6539));
    layer1_outputs(2604) <= not(layer0_outputs(4194));
    layer1_outputs(2605) <= not(layer0_outputs(7253));
    layer1_outputs(2606) <= not((layer0_outputs(6189)) and (layer0_outputs(5008)));
    layer1_outputs(2607) <= '0';
    layer1_outputs(2608) <= '1';
    layer1_outputs(2609) <= not((layer0_outputs(4266)) and (layer0_outputs(5535)));
    layer1_outputs(2610) <= (layer0_outputs(1652)) and not (layer0_outputs(1770));
    layer1_outputs(2611) <= (layer0_outputs(2528)) and not (layer0_outputs(6812));
    layer1_outputs(2612) <= '1';
    layer1_outputs(2613) <= (layer0_outputs(637)) and (layer0_outputs(6663));
    layer1_outputs(2614) <= not(layer0_outputs(886));
    layer1_outputs(2615) <= not(layer0_outputs(7637)) or (layer0_outputs(3012));
    layer1_outputs(2616) <= not(layer0_outputs(1836));
    layer1_outputs(2617) <= layer0_outputs(4405);
    layer1_outputs(2618) <= not(layer0_outputs(791));
    layer1_outputs(2619) <= not(layer0_outputs(5911)) or (layer0_outputs(2870));
    layer1_outputs(2620) <= '1';
    layer1_outputs(2621) <= not(layer0_outputs(7318));
    layer1_outputs(2622) <= (layer0_outputs(7312)) and (layer0_outputs(3505));
    layer1_outputs(2623) <= layer0_outputs(2408);
    layer1_outputs(2624) <= not(layer0_outputs(6102));
    layer1_outputs(2625) <= not((layer0_outputs(5581)) or (layer0_outputs(5768)));
    layer1_outputs(2626) <= not((layer0_outputs(5916)) or (layer0_outputs(4818)));
    layer1_outputs(2627) <= (layer0_outputs(2099)) or (layer0_outputs(2397));
    layer1_outputs(2628) <= not((layer0_outputs(1871)) and (layer0_outputs(7554)));
    layer1_outputs(2629) <= not(layer0_outputs(3830));
    layer1_outputs(2630) <= not(layer0_outputs(350));
    layer1_outputs(2631) <= '0';
    layer1_outputs(2632) <= not((layer0_outputs(389)) or (layer0_outputs(5179)));
    layer1_outputs(2633) <= not((layer0_outputs(5208)) and (layer0_outputs(5581)));
    layer1_outputs(2634) <= layer0_outputs(5952);
    layer1_outputs(2635) <= not(layer0_outputs(1927)) or (layer0_outputs(7136));
    layer1_outputs(2636) <= layer0_outputs(4708);
    layer1_outputs(2637) <= not(layer0_outputs(2270));
    layer1_outputs(2638) <= (layer0_outputs(2699)) and (layer0_outputs(3937));
    layer1_outputs(2639) <= not(layer0_outputs(5084)) or (layer0_outputs(1745));
    layer1_outputs(2640) <= (layer0_outputs(654)) and not (layer0_outputs(3807));
    layer1_outputs(2641) <= not((layer0_outputs(2888)) and (layer0_outputs(2241)));
    layer1_outputs(2642) <= (layer0_outputs(2842)) and (layer0_outputs(1606));
    layer1_outputs(2643) <= not(layer0_outputs(6589));
    layer1_outputs(2644) <= not((layer0_outputs(3338)) or (layer0_outputs(2728)));
    layer1_outputs(2645) <= '0';
    layer1_outputs(2646) <= not(layer0_outputs(1728));
    layer1_outputs(2647) <= not(layer0_outputs(2907)) or (layer0_outputs(7435));
    layer1_outputs(2648) <= not(layer0_outputs(4859)) or (layer0_outputs(5198));
    layer1_outputs(2649) <= (layer0_outputs(7027)) and not (layer0_outputs(2904));
    layer1_outputs(2650) <= layer0_outputs(4895);
    layer1_outputs(2651) <= not(layer0_outputs(4658));
    layer1_outputs(2652) <= (layer0_outputs(1585)) and not (layer0_outputs(4641));
    layer1_outputs(2653) <= layer0_outputs(4624);
    layer1_outputs(2654) <= not(layer0_outputs(4689)) or (layer0_outputs(6376));
    layer1_outputs(2655) <= '1';
    layer1_outputs(2656) <= (layer0_outputs(1038)) or (layer0_outputs(5667));
    layer1_outputs(2657) <= (layer0_outputs(1839)) or (layer0_outputs(4820));
    layer1_outputs(2658) <= not(layer0_outputs(6146)) or (layer0_outputs(2826));
    layer1_outputs(2659) <= (layer0_outputs(6718)) and (layer0_outputs(1828));
    layer1_outputs(2660) <= (layer0_outputs(3543)) and not (layer0_outputs(4988));
    layer1_outputs(2661) <= layer0_outputs(6753);
    layer1_outputs(2662) <= (layer0_outputs(4303)) or (layer0_outputs(5459));
    layer1_outputs(2663) <= '0';
    layer1_outputs(2664) <= layer0_outputs(4143);
    layer1_outputs(2665) <= '1';
    layer1_outputs(2666) <= (layer0_outputs(1735)) and not (layer0_outputs(4993));
    layer1_outputs(2667) <= (layer0_outputs(2386)) or (layer0_outputs(3711));
    layer1_outputs(2668) <= not((layer0_outputs(270)) or (layer0_outputs(7153)));
    layer1_outputs(2669) <= '0';
    layer1_outputs(2670) <= layer0_outputs(4377);
    layer1_outputs(2671) <= layer0_outputs(1324);
    layer1_outputs(2672) <= '1';
    layer1_outputs(2673) <= not(layer0_outputs(5721));
    layer1_outputs(2674) <= not((layer0_outputs(5189)) xor (layer0_outputs(6424)));
    layer1_outputs(2675) <= (layer0_outputs(7590)) or (layer0_outputs(2045));
    layer1_outputs(2676) <= '0';
    layer1_outputs(2677) <= '1';
    layer1_outputs(2678) <= (layer0_outputs(6380)) or (layer0_outputs(929));
    layer1_outputs(2679) <= '1';
    layer1_outputs(2680) <= not((layer0_outputs(7545)) or (layer0_outputs(2396)));
    layer1_outputs(2681) <= '1';
    layer1_outputs(2682) <= (layer0_outputs(126)) and not (layer0_outputs(3682));
    layer1_outputs(2683) <= not((layer0_outputs(615)) or (layer0_outputs(2714)));
    layer1_outputs(2684) <= (layer0_outputs(3798)) or (layer0_outputs(1627));
    layer1_outputs(2685) <= '0';
    layer1_outputs(2686) <= not((layer0_outputs(6061)) and (layer0_outputs(7092)));
    layer1_outputs(2687) <= not(layer0_outputs(1123));
    layer1_outputs(2688) <= not(layer0_outputs(7083)) or (layer0_outputs(2589));
    layer1_outputs(2689) <= '0';
    layer1_outputs(2690) <= (layer0_outputs(2217)) and not (layer0_outputs(4217));
    layer1_outputs(2691) <= not(layer0_outputs(4262));
    layer1_outputs(2692) <= not((layer0_outputs(6551)) xor (layer0_outputs(2383)));
    layer1_outputs(2693) <= (layer0_outputs(380)) and not (layer0_outputs(7058));
    layer1_outputs(2694) <= not(layer0_outputs(2251));
    layer1_outputs(2695) <= not((layer0_outputs(5461)) or (layer0_outputs(5330)));
    layer1_outputs(2696) <= not(layer0_outputs(5798));
    layer1_outputs(2697) <= layer0_outputs(4115);
    layer1_outputs(2698) <= (layer0_outputs(2712)) and not (layer0_outputs(304));
    layer1_outputs(2699) <= (layer0_outputs(1843)) and not (layer0_outputs(1643));
    layer1_outputs(2700) <= not((layer0_outputs(5497)) and (layer0_outputs(3393)));
    layer1_outputs(2701) <= (layer0_outputs(4003)) and not (layer0_outputs(3829));
    layer1_outputs(2702) <= '0';
    layer1_outputs(2703) <= not(layer0_outputs(4301));
    layer1_outputs(2704) <= '1';
    layer1_outputs(2705) <= (layer0_outputs(5264)) and not (layer0_outputs(3007));
    layer1_outputs(2706) <= '0';
    layer1_outputs(2707) <= layer0_outputs(2980);
    layer1_outputs(2708) <= (layer0_outputs(230)) and not (layer0_outputs(6495));
    layer1_outputs(2709) <= (layer0_outputs(3553)) and (layer0_outputs(3397));
    layer1_outputs(2710) <= not((layer0_outputs(1152)) and (layer0_outputs(1404)));
    layer1_outputs(2711) <= (layer0_outputs(4253)) and not (layer0_outputs(3699));
    layer1_outputs(2712) <= not(layer0_outputs(1790));
    layer1_outputs(2713) <= not(layer0_outputs(1740)) or (layer0_outputs(280));
    layer1_outputs(2714) <= '1';
    layer1_outputs(2715) <= '0';
    layer1_outputs(2716) <= '0';
    layer1_outputs(2717) <= not(layer0_outputs(3847));
    layer1_outputs(2718) <= not(layer0_outputs(7621));
    layer1_outputs(2719) <= not(layer0_outputs(3163)) or (layer0_outputs(938));
    layer1_outputs(2720) <= layer0_outputs(5010);
    layer1_outputs(2721) <= (layer0_outputs(6642)) or (layer0_outputs(7182));
    layer1_outputs(2722) <= not((layer0_outputs(1921)) and (layer0_outputs(7651)));
    layer1_outputs(2723) <= (layer0_outputs(5156)) and not (layer0_outputs(4499));
    layer1_outputs(2724) <= (layer0_outputs(3675)) and (layer0_outputs(5348));
    layer1_outputs(2725) <= not(layer0_outputs(2574)) or (layer0_outputs(7521));
    layer1_outputs(2726) <= not(layer0_outputs(2054));
    layer1_outputs(2727) <= (layer0_outputs(2214)) and (layer0_outputs(5316));
    layer1_outputs(2728) <= (layer0_outputs(2326)) or (layer0_outputs(2380));
    layer1_outputs(2729) <= (layer0_outputs(6459)) and not (layer0_outputs(7536));
    layer1_outputs(2730) <= '0';
    layer1_outputs(2731) <= not(layer0_outputs(2640)) or (layer0_outputs(4113));
    layer1_outputs(2732) <= layer0_outputs(6127);
    layer1_outputs(2733) <= not((layer0_outputs(1393)) and (layer0_outputs(5343)));
    layer1_outputs(2734) <= not(layer0_outputs(820)) or (layer0_outputs(591));
    layer1_outputs(2735) <= layer0_outputs(5108);
    layer1_outputs(2736) <= (layer0_outputs(5732)) and not (layer0_outputs(3838));
    layer1_outputs(2737) <= not(layer0_outputs(3183));
    layer1_outputs(2738) <= (layer0_outputs(5980)) and not (layer0_outputs(1516));
    layer1_outputs(2739) <= not(layer0_outputs(1173));
    layer1_outputs(2740) <= not((layer0_outputs(2982)) and (layer0_outputs(2310)));
    layer1_outputs(2741) <= not(layer0_outputs(1714));
    layer1_outputs(2742) <= '0';
    layer1_outputs(2743) <= '1';
    layer1_outputs(2744) <= (layer0_outputs(5365)) or (layer0_outputs(5869));
    layer1_outputs(2745) <= not((layer0_outputs(2274)) and (layer0_outputs(6334)));
    layer1_outputs(2746) <= not(layer0_outputs(4440));
    layer1_outputs(2747) <= not(layer0_outputs(5501)) or (layer0_outputs(751));
    layer1_outputs(2748) <= (layer0_outputs(1132)) or (layer0_outputs(6772));
    layer1_outputs(2749) <= not((layer0_outputs(2210)) and (layer0_outputs(6832)));
    layer1_outputs(2750) <= not(layer0_outputs(3947));
    layer1_outputs(2751) <= (layer0_outputs(6601)) and not (layer0_outputs(7653));
    layer1_outputs(2752) <= not((layer0_outputs(6228)) or (layer0_outputs(2575)));
    layer1_outputs(2753) <= (layer0_outputs(739)) xor (layer0_outputs(4965));
    layer1_outputs(2754) <= '1';
    layer1_outputs(2755) <= (layer0_outputs(1631)) and (layer0_outputs(2171));
    layer1_outputs(2756) <= (layer0_outputs(1828)) or (layer0_outputs(3977));
    layer1_outputs(2757) <= layer0_outputs(7569);
    layer1_outputs(2758) <= not((layer0_outputs(2097)) or (layer0_outputs(957)));
    layer1_outputs(2759) <= (layer0_outputs(2632)) xor (layer0_outputs(7550));
    layer1_outputs(2760) <= not(layer0_outputs(4880));
    layer1_outputs(2761) <= layer0_outputs(7371);
    layer1_outputs(2762) <= '0';
    layer1_outputs(2763) <= (layer0_outputs(4245)) and (layer0_outputs(4073));
    layer1_outputs(2764) <= not(layer0_outputs(4619)) or (layer0_outputs(7197));
    layer1_outputs(2765) <= '0';
    layer1_outputs(2766) <= layer0_outputs(7330);
    layer1_outputs(2767) <= layer0_outputs(7233);
    layer1_outputs(2768) <= (layer0_outputs(2622)) and not (layer0_outputs(6365));
    layer1_outputs(2769) <= layer0_outputs(4082);
    layer1_outputs(2770) <= (layer0_outputs(717)) and not (layer0_outputs(6963));
    layer1_outputs(2771) <= not(layer0_outputs(285)) or (layer0_outputs(6870));
    layer1_outputs(2772) <= not(layer0_outputs(2148));
    layer1_outputs(2773) <= not(layer0_outputs(2540));
    layer1_outputs(2774) <= (layer0_outputs(7347)) and not (layer0_outputs(2880));
    layer1_outputs(2775) <= (layer0_outputs(2325)) and not (layer0_outputs(2586));
    layer1_outputs(2776) <= not(layer0_outputs(5879)) or (layer0_outputs(5473));
    layer1_outputs(2777) <= (layer0_outputs(4277)) or (layer0_outputs(4025));
    layer1_outputs(2778) <= not(layer0_outputs(5587)) or (layer0_outputs(2277));
    layer1_outputs(2779) <= not(layer0_outputs(3073));
    layer1_outputs(2780) <= layer0_outputs(90);
    layer1_outputs(2781) <= '1';
    layer1_outputs(2782) <= layer0_outputs(5683);
    layer1_outputs(2783) <= layer0_outputs(2582);
    layer1_outputs(2784) <= layer0_outputs(7454);
    layer1_outputs(2785) <= not(layer0_outputs(6016));
    layer1_outputs(2786) <= (layer0_outputs(5394)) and not (layer0_outputs(3741));
    layer1_outputs(2787) <= not(layer0_outputs(3884)) or (layer0_outputs(6436));
    layer1_outputs(2788) <= layer0_outputs(3002);
    layer1_outputs(2789) <= '1';
    layer1_outputs(2790) <= not(layer0_outputs(2141)) or (layer0_outputs(1954));
    layer1_outputs(2791) <= (layer0_outputs(2146)) or (layer0_outputs(6159));
    layer1_outputs(2792) <= (layer0_outputs(47)) and (layer0_outputs(6322));
    layer1_outputs(2793) <= (layer0_outputs(568)) xor (layer0_outputs(767));
    layer1_outputs(2794) <= not(layer0_outputs(4594)) or (layer0_outputs(6097));
    layer1_outputs(2795) <= (layer0_outputs(6010)) and (layer0_outputs(6268));
    layer1_outputs(2796) <= (layer0_outputs(3490)) or (layer0_outputs(799));
    layer1_outputs(2797) <= not((layer0_outputs(6044)) and (layer0_outputs(4429)));
    layer1_outputs(2798) <= (layer0_outputs(3788)) or (layer0_outputs(4577));
    layer1_outputs(2799) <= (layer0_outputs(4598)) and not (layer0_outputs(2660));
    layer1_outputs(2800) <= not(layer0_outputs(984));
    layer1_outputs(2801) <= not((layer0_outputs(1443)) or (layer0_outputs(2865)));
    layer1_outputs(2802) <= not(layer0_outputs(2441));
    layer1_outputs(2803) <= layer0_outputs(506);
    layer1_outputs(2804) <= layer0_outputs(4683);
    layer1_outputs(2805) <= (layer0_outputs(2876)) and not (layer0_outputs(5871));
    layer1_outputs(2806) <= layer0_outputs(3277);
    layer1_outputs(2807) <= not(layer0_outputs(1016)) or (layer0_outputs(3814));
    layer1_outputs(2808) <= '1';
    layer1_outputs(2809) <= '1';
    layer1_outputs(2810) <= (layer0_outputs(698)) and not (layer0_outputs(3782));
    layer1_outputs(2811) <= not((layer0_outputs(1901)) xor (layer0_outputs(3904)));
    layer1_outputs(2812) <= not(layer0_outputs(2191));
    layer1_outputs(2813) <= not(layer0_outputs(4158)) or (layer0_outputs(4483));
    layer1_outputs(2814) <= not(layer0_outputs(2654));
    layer1_outputs(2815) <= not(layer0_outputs(1013)) or (layer0_outputs(4501));
    layer1_outputs(2816) <= layer0_outputs(4718);
    layer1_outputs(2817) <= (layer0_outputs(4169)) or (layer0_outputs(4775));
    layer1_outputs(2818) <= (layer0_outputs(5353)) and not (layer0_outputs(108));
    layer1_outputs(2819) <= (layer0_outputs(7247)) and not (layer0_outputs(2224));
    layer1_outputs(2820) <= not(layer0_outputs(2278)) or (layer0_outputs(3270));
    layer1_outputs(2821) <= (layer0_outputs(4078)) and not (layer0_outputs(2295));
    layer1_outputs(2822) <= '0';
    layer1_outputs(2823) <= (layer0_outputs(6182)) and (layer0_outputs(3631));
    layer1_outputs(2824) <= layer0_outputs(4051);
    layer1_outputs(2825) <= not((layer0_outputs(2837)) or (layer0_outputs(11)));
    layer1_outputs(2826) <= '0';
    layer1_outputs(2827) <= (layer0_outputs(7436)) and not (layer0_outputs(958));
    layer1_outputs(2828) <= layer0_outputs(6396);
    layer1_outputs(2829) <= not(layer0_outputs(2821));
    layer1_outputs(2830) <= layer0_outputs(1276);
    layer1_outputs(2831) <= '1';
    layer1_outputs(2832) <= not(layer0_outputs(4126)) or (layer0_outputs(4125));
    layer1_outputs(2833) <= (layer0_outputs(4211)) or (layer0_outputs(2497));
    layer1_outputs(2834) <= '1';
    layer1_outputs(2835) <= (layer0_outputs(2044)) or (layer0_outputs(7565));
    layer1_outputs(2836) <= '1';
    layer1_outputs(2837) <= '1';
    layer1_outputs(2838) <= not((layer0_outputs(7222)) and (layer0_outputs(7213)));
    layer1_outputs(2839) <= '0';
    layer1_outputs(2840) <= '0';
    layer1_outputs(2841) <= (layer0_outputs(5224)) and not (layer0_outputs(6485));
    layer1_outputs(2842) <= not((layer0_outputs(563)) or (layer0_outputs(3870)));
    layer1_outputs(2843) <= '1';
    layer1_outputs(2844) <= not(layer0_outputs(2855)) or (layer0_outputs(6550));
    layer1_outputs(2845) <= (layer0_outputs(1779)) or (layer0_outputs(1051));
    layer1_outputs(2846) <= '0';
    layer1_outputs(2847) <= (layer0_outputs(7132)) and (layer0_outputs(6068));
    layer1_outputs(2848) <= not((layer0_outputs(5358)) xor (layer0_outputs(6244)));
    layer1_outputs(2849) <= layer0_outputs(4203);
    layer1_outputs(2850) <= '0';
    layer1_outputs(2851) <= not((layer0_outputs(2388)) or (layer0_outputs(4172)));
    layer1_outputs(2852) <= not((layer0_outputs(5852)) or (layer0_outputs(3139)));
    layer1_outputs(2853) <= (layer0_outputs(1501)) and not (layer0_outputs(2293));
    layer1_outputs(2854) <= not(layer0_outputs(4116));
    layer1_outputs(2855) <= not(layer0_outputs(2395));
    layer1_outputs(2856) <= (layer0_outputs(6446)) and not (layer0_outputs(697));
    layer1_outputs(2857) <= (layer0_outputs(3820)) and not (layer0_outputs(4479));
    layer1_outputs(2858) <= not((layer0_outputs(6885)) xor (layer0_outputs(5207)));
    layer1_outputs(2859) <= (layer0_outputs(4063)) and not (layer0_outputs(2033));
    layer1_outputs(2860) <= '0';
    layer1_outputs(2861) <= not(layer0_outputs(5477)) or (layer0_outputs(3213));
    layer1_outputs(2862) <= not(layer0_outputs(7212)) or (layer0_outputs(5714));
    layer1_outputs(2863) <= not((layer0_outputs(141)) or (layer0_outputs(4767)));
    layer1_outputs(2864) <= layer0_outputs(164);
    layer1_outputs(2865) <= (layer0_outputs(1630)) and not (layer0_outputs(5351));
    layer1_outputs(2866) <= (layer0_outputs(594)) xor (layer0_outputs(2576));
    layer1_outputs(2867) <= not(layer0_outputs(3020));
    layer1_outputs(2868) <= (layer0_outputs(5130)) and (layer0_outputs(3122));
    layer1_outputs(2869) <= not((layer0_outputs(2227)) and (layer0_outputs(5130)));
    layer1_outputs(2870) <= not(layer0_outputs(1636));
    layer1_outputs(2871) <= '0';
    layer1_outputs(2872) <= not(layer0_outputs(7096)) or (layer0_outputs(7616));
    layer1_outputs(2873) <= (layer0_outputs(983)) and not (layer0_outputs(4691));
    layer1_outputs(2874) <= not(layer0_outputs(7649));
    layer1_outputs(2875) <= (layer0_outputs(7153)) and not (layer0_outputs(6837));
    layer1_outputs(2876) <= not(layer0_outputs(7466)) or (layer0_outputs(5187));
    layer1_outputs(2877) <= not(layer0_outputs(5438)) or (layer0_outputs(1093));
    layer1_outputs(2878) <= '1';
    layer1_outputs(2879) <= (layer0_outputs(215)) xor (layer0_outputs(5308));
    layer1_outputs(2880) <= (layer0_outputs(2591)) or (layer0_outputs(6315));
    layer1_outputs(2881) <= '0';
    layer1_outputs(2882) <= not(layer0_outputs(3206));
    layer1_outputs(2883) <= not(layer0_outputs(2401));
    layer1_outputs(2884) <= not((layer0_outputs(952)) and (layer0_outputs(6211)));
    layer1_outputs(2885) <= layer0_outputs(1009);
    layer1_outputs(2886) <= '1';
    layer1_outputs(2887) <= not((layer0_outputs(3909)) and (layer0_outputs(757)));
    layer1_outputs(2888) <= '0';
    layer1_outputs(2889) <= (layer0_outputs(3820)) or (layer0_outputs(3775));
    layer1_outputs(2890) <= not(layer0_outputs(6489)) or (layer0_outputs(1546));
    layer1_outputs(2891) <= (layer0_outputs(4077)) and not (layer0_outputs(3036));
    layer1_outputs(2892) <= not(layer0_outputs(1753)) or (layer0_outputs(3877));
    layer1_outputs(2893) <= not(layer0_outputs(404));
    layer1_outputs(2894) <= '1';
    layer1_outputs(2895) <= not((layer0_outputs(4383)) or (layer0_outputs(3325)));
    layer1_outputs(2896) <= '1';
    layer1_outputs(2897) <= not((layer0_outputs(1776)) and (layer0_outputs(3408)));
    layer1_outputs(2898) <= '1';
    layer1_outputs(2899) <= not(layer0_outputs(744));
    layer1_outputs(2900) <= (layer0_outputs(4297)) xor (layer0_outputs(169));
    layer1_outputs(2901) <= (layer0_outputs(5745)) or (layer0_outputs(3499));
    layer1_outputs(2902) <= layer0_outputs(2221);
    layer1_outputs(2903) <= layer0_outputs(6930);
    layer1_outputs(2904) <= '1';
    layer1_outputs(2905) <= not(layer0_outputs(5885)) or (layer0_outputs(4026));
    layer1_outputs(2906) <= layer0_outputs(977);
    layer1_outputs(2907) <= (layer0_outputs(5802)) and (layer0_outputs(4685));
    layer1_outputs(2908) <= not((layer0_outputs(163)) or (layer0_outputs(4604)));
    layer1_outputs(2909) <= '1';
    layer1_outputs(2910) <= (layer0_outputs(7116)) and not (layer0_outputs(3104));
    layer1_outputs(2911) <= layer0_outputs(4826);
    layer1_outputs(2912) <= not(layer0_outputs(1532)) or (layer0_outputs(6776));
    layer1_outputs(2913) <= layer0_outputs(4681);
    layer1_outputs(2914) <= '1';
    layer1_outputs(2915) <= '0';
    layer1_outputs(2916) <= layer0_outputs(2627);
    layer1_outputs(2917) <= '0';
    layer1_outputs(2918) <= '0';
    layer1_outputs(2919) <= not(layer0_outputs(3398)) or (layer0_outputs(3689));
    layer1_outputs(2920) <= layer0_outputs(1591);
    layer1_outputs(2921) <= '1';
    layer1_outputs(2922) <= not(layer0_outputs(6141));
    layer1_outputs(2923) <= not((layer0_outputs(3830)) and (layer0_outputs(5786)));
    layer1_outputs(2924) <= not(layer0_outputs(844)) or (layer0_outputs(6926));
    layer1_outputs(2925) <= layer0_outputs(3948);
    layer1_outputs(2926) <= not(layer0_outputs(1063));
    layer1_outputs(2927) <= '1';
    layer1_outputs(2928) <= '0';
    layer1_outputs(2929) <= layer0_outputs(639);
    layer1_outputs(2930) <= not(layer0_outputs(1378)) or (layer0_outputs(1674));
    layer1_outputs(2931) <= (layer0_outputs(875)) or (layer0_outputs(1187));
    layer1_outputs(2932) <= layer0_outputs(3944);
    layer1_outputs(2933) <= (layer0_outputs(7323)) and not (layer0_outputs(2553));
    layer1_outputs(2934) <= (layer0_outputs(6700)) and (layer0_outputs(1587));
    layer1_outputs(2935) <= (layer0_outputs(4711)) and (layer0_outputs(6964));
    layer1_outputs(2936) <= not(layer0_outputs(6860)) or (layer0_outputs(6474));
    layer1_outputs(2937) <= (layer0_outputs(4094)) and not (layer0_outputs(2879));
    layer1_outputs(2938) <= (layer0_outputs(2996)) and not (layer0_outputs(7146));
    layer1_outputs(2939) <= layer0_outputs(2665);
    layer1_outputs(2940) <= not((layer0_outputs(5991)) or (layer0_outputs(6025)));
    layer1_outputs(2941) <= not((layer0_outputs(5729)) or (layer0_outputs(2535)));
    layer1_outputs(2942) <= not(layer0_outputs(5182));
    layer1_outputs(2943) <= '1';
    layer1_outputs(2944) <= layer0_outputs(3761);
    layer1_outputs(2945) <= not(layer0_outputs(5298));
    layer1_outputs(2946) <= '1';
    layer1_outputs(2947) <= '1';
    layer1_outputs(2948) <= (layer0_outputs(3854)) and not (layer0_outputs(143));
    layer1_outputs(2949) <= not((layer0_outputs(1094)) and (layer0_outputs(3207)));
    layer1_outputs(2950) <= layer0_outputs(6660);
    layer1_outputs(2951) <= not(layer0_outputs(239)) or (layer0_outputs(2011));
    layer1_outputs(2952) <= not(layer0_outputs(3655)) or (layer0_outputs(2537));
    layer1_outputs(2953) <= '1';
    layer1_outputs(2954) <= '1';
    layer1_outputs(2955) <= '0';
    layer1_outputs(2956) <= layer0_outputs(123);
    layer1_outputs(2957) <= not(layer0_outputs(5867)) or (layer0_outputs(7445));
    layer1_outputs(2958) <= '1';
    layer1_outputs(2959) <= not(layer0_outputs(6862));
    layer1_outputs(2960) <= not(layer0_outputs(7247));
    layer1_outputs(2961) <= (layer0_outputs(1563)) and not (layer0_outputs(3435));
    layer1_outputs(2962) <= '1';
    layer1_outputs(2963) <= (layer0_outputs(5192)) and (layer0_outputs(1605));
    layer1_outputs(2964) <= '1';
    layer1_outputs(2965) <= (layer0_outputs(4743)) and (layer0_outputs(4559));
    layer1_outputs(2966) <= '1';
    layer1_outputs(2967) <= '0';
    layer1_outputs(2968) <= (layer0_outputs(4139)) xor (layer0_outputs(1667));
    layer1_outputs(2969) <= not((layer0_outputs(5935)) or (layer0_outputs(3658)));
    layer1_outputs(2970) <= layer0_outputs(2179);
    layer1_outputs(2971) <= not(layer0_outputs(3023));
    layer1_outputs(2972) <= not(layer0_outputs(2382)) or (layer0_outputs(1198));
    layer1_outputs(2973) <= not(layer0_outputs(1654)) or (layer0_outputs(6808));
    layer1_outputs(2974) <= not((layer0_outputs(509)) xor (layer0_outputs(5941)));
    layer1_outputs(2975) <= layer0_outputs(7655);
    layer1_outputs(2976) <= (layer0_outputs(539)) and not (layer0_outputs(446));
    layer1_outputs(2977) <= not(layer0_outputs(3671));
    layer1_outputs(2978) <= '1';
    layer1_outputs(2979) <= not(layer0_outputs(6082));
    layer1_outputs(2980) <= '0';
    layer1_outputs(2981) <= layer0_outputs(2266);
    layer1_outputs(2982) <= not(layer0_outputs(2769)) or (layer0_outputs(4541));
    layer1_outputs(2983) <= '1';
    layer1_outputs(2984) <= not(layer0_outputs(6507)) or (layer0_outputs(3611));
    layer1_outputs(2985) <= (layer0_outputs(302)) xor (layer0_outputs(1948));
    layer1_outputs(2986) <= not(layer0_outputs(6483)) or (layer0_outputs(6448));
    layer1_outputs(2987) <= not(layer0_outputs(3545)) or (layer0_outputs(142));
    layer1_outputs(2988) <= (layer0_outputs(554)) and (layer0_outputs(3250));
    layer1_outputs(2989) <= not(layer0_outputs(3561));
    layer1_outputs(2990) <= not((layer0_outputs(824)) or (layer0_outputs(537)));
    layer1_outputs(2991) <= (layer0_outputs(5820)) and not (layer0_outputs(2898));
    layer1_outputs(2992) <= not(layer0_outputs(3481)) or (layer0_outputs(3026));
    layer1_outputs(2993) <= (layer0_outputs(3598)) or (layer0_outputs(4365));
    layer1_outputs(2994) <= '1';
    layer1_outputs(2995) <= not((layer0_outputs(6041)) or (layer0_outputs(5913)));
    layer1_outputs(2996) <= not((layer0_outputs(1409)) xor (layer0_outputs(6258)));
    layer1_outputs(2997) <= not(layer0_outputs(4403));
    layer1_outputs(2998) <= '1';
    layer1_outputs(2999) <= not(layer0_outputs(2670));
    layer1_outputs(3000) <= not((layer0_outputs(3428)) or (layer0_outputs(6132)));
    layer1_outputs(3001) <= '0';
    layer1_outputs(3002) <= '0';
    layer1_outputs(3003) <= (layer0_outputs(5237)) or (layer0_outputs(5168));
    layer1_outputs(3004) <= not(layer0_outputs(5783));
    layer1_outputs(3005) <= layer0_outputs(4000);
    layer1_outputs(3006) <= not(layer0_outputs(4135)) or (layer0_outputs(326));
    layer1_outputs(3007) <= '0';
    layer1_outputs(3008) <= (layer0_outputs(960)) and not (layer0_outputs(7629));
    layer1_outputs(3009) <= '1';
    layer1_outputs(3010) <= layer0_outputs(3423);
    layer1_outputs(3011) <= layer0_outputs(4805);
    layer1_outputs(3012) <= not(layer0_outputs(7671)) or (layer0_outputs(1802));
    layer1_outputs(3013) <= layer0_outputs(35);
    layer1_outputs(3014) <= not((layer0_outputs(491)) or (layer0_outputs(479)));
    layer1_outputs(3015) <= not(layer0_outputs(3101));
    layer1_outputs(3016) <= not(layer0_outputs(6840)) or (layer0_outputs(4606));
    layer1_outputs(3017) <= (layer0_outputs(1175)) or (layer0_outputs(2743));
    layer1_outputs(3018) <= layer0_outputs(7617);
    layer1_outputs(3019) <= (layer0_outputs(2695)) and not (layer0_outputs(226));
    layer1_outputs(3020) <= (layer0_outputs(7625)) or (layer0_outputs(2177));
    layer1_outputs(3021) <= '0';
    layer1_outputs(3022) <= layer0_outputs(7535);
    layer1_outputs(3023) <= layer0_outputs(1337);
    layer1_outputs(3024) <= layer0_outputs(2584);
    layer1_outputs(3025) <= '0';
    layer1_outputs(3026) <= (layer0_outputs(6688)) and (layer0_outputs(1980));
    layer1_outputs(3027) <= not((layer0_outputs(5906)) or (layer0_outputs(2481)));
    layer1_outputs(3028) <= '1';
    layer1_outputs(3029) <= '1';
    layer1_outputs(3030) <= not((layer0_outputs(1578)) and (layer0_outputs(3008)));
    layer1_outputs(3031) <= (layer0_outputs(4381)) and not (layer0_outputs(2882));
    layer1_outputs(3032) <= layer0_outputs(3629);
    layer1_outputs(3033) <= '1';
    layer1_outputs(3034) <= layer0_outputs(7428);
    layer1_outputs(3035) <= '0';
    layer1_outputs(3036) <= not((layer0_outputs(7391)) or (layer0_outputs(2965)));
    layer1_outputs(3037) <= '0';
    layer1_outputs(3038) <= not(layer0_outputs(1638)) or (layer0_outputs(4582));
    layer1_outputs(3039) <= layer0_outputs(4705);
    layer1_outputs(3040) <= not(layer0_outputs(6991));
    layer1_outputs(3041) <= not((layer0_outputs(4230)) or (layer0_outputs(36)));
    layer1_outputs(3042) <= layer0_outputs(717);
    layer1_outputs(3043) <= not(layer0_outputs(245));
    layer1_outputs(3044) <= layer0_outputs(1129);
    layer1_outputs(3045) <= '0';
    layer1_outputs(3046) <= '1';
    layer1_outputs(3047) <= not(layer0_outputs(6532)) or (layer0_outputs(5414));
    layer1_outputs(3048) <= not(layer0_outputs(4481));
    layer1_outputs(3049) <= not(layer0_outputs(6927)) or (layer0_outputs(5375));
    layer1_outputs(3050) <= layer0_outputs(7638);
    layer1_outputs(3051) <= '0';
    layer1_outputs(3052) <= not((layer0_outputs(2483)) or (layer0_outputs(7296)));
    layer1_outputs(3053) <= (layer0_outputs(3149)) and not (layer0_outputs(617));
    layer1_outputs(3054) <= not(layer0_outputs(5292)) or (layer0_outputs(6616));
    layer1_outputs(3055) <= (layer0_outputs(3293)) and not (layer0_outputs(4929));
    layer1_outputs(3056) <= not(layer0_outputs(4042));
    layer1_outputs(3057) <= not(layer0_outputs(6575)) or (layer0_outputs(3493));
    layer1_outputs(3058) <= layer0_outputs(5766);
    layer1_outputs(3059) <= '0';
    layer1_outputs(3060) <= (layer0_outputs(1394)) and not (layer0_outputs(6339));
    layer1_outputs(3061) <= not(layer0_outputs(5839));
    layer1_outputs(3062) <= not((layer0_outputs(1904)) xor (layer0_outputs(363)));
    layer1_outputs(3063) <= not(layer0_outputs(4512)) or (layer0_outputs(7543));
    layer1_outputs(3064) <= (layer0_outputs(1091)) and not (layer0_outputs(5959));
    layer1_outputs(3065) <= not(layer0_outputs(5194)) or (layer0_outputs(2612));
    layer1_outputs(3066) <= not((layer0_outputs(5747)) and (layer0_outputs(1961)));
    layer1_outputs(3067) <= not((layer0_outputs(3279)) or (layer0_outputs(4530)));
    layer1_outputs(3068) <= (layer0_outputs(3451)) or (layer0_outputs(5895));
    layer1_outputs(3069) <= '0';
    layer1_outputs(3070) <= layer0_outputs(106);
    layer1_outputs(3071) <= '0';
    layer1_outputs(3072) <= layer0_outputs(2885);
    layer1_outputs(3073) <= layer0_outputs(525);
    layer1_outputs(3074) <= '1';
    layer1_outputs(3075) <= not(layer0_outputs(663));
    layer1_outputs(3076) <= (layer0_outputs(3672)) and not (layer0_outputs(5322));
    layer1_outputs(3077) <= (layer0_outputs(1088)) and not (layer0_outputs(810));
    layer1_outputs(3078) <= not(layer0_outputs(7318)) or (layer0_outputs(7174));
    layer1_outputs(3079) <= not(layer0_outputs(4321)) or (layer0_outputs(7376));
    layer1_outputs(3080) <= not(layer0_outputs(6604)) or (layer0_outputs(7640));
    layer1_outputs(3081) <= layer0_outputs(2433);
    layer1_outputs(3082) <= layer0_outputs(4783);
    layer1_outputs(3083) <= not(layer0_outputs(590)) or (layer0_outputs(1741));
    layer1_outputs(3084) <= layer0_outputs(67);
    layer1_outputs(3085) <= not(layer0_outputs(3430));
    layer1_outputs(3086) <= not(layer0_outputs(4068));
    layer1_outputs(3087) <= not((layer0_outputs(216)) or (layer0_outputs(2081)));
    layer1_outputs(3088) <= not(layer0_outputs(3569)) or (layer0_outputs(2393));
    layer1_outputs(3089) <= not((layer0_outputs(207)) xor (layer0_outputs(5710)));
    layer1_outputs(3090) <= (layer0_outputs(7115)) and not (layer0_outputs(583));
    layer1_outputs(3091) <= not(layer0_outputs(6958)) or (layer0_outputs(3186));
    layer1_outputs(3092) <= not((layer0_outputs(5555)) and (layer0_outputs(12)));
    layer1_outputs(3093) <= (layer0_outputs(810)) and (layer0_outputs(5582));
    layer1_outputs(3094) <= not(layer0_outputs(7476));
    layer1_outputs(3095) <= (layer0_outputs(105)) and not (layer0_outputs(2623));
    layer1_outputs(3096) <= not(layer0_outputs(7299));
    layer1_outputs(3097) <= (layer0_outputs(5799)) and (layer0_outputs(4057));
    layer1_outputs(3098) <= '1';
    layer1_outputs(3099) <= '1';
    layer1_outputs(3100) <= layer0_outputs(6435);
    layer1_outputs(3101) <= layer0_outputs(2234);
    layer1_outputs(3102) <= (layer0_outputs(4500)) and not (layer0_outputs(4748));
    layer1_outputs(3103) <= layer0_outputs(4198);
    layer1_outputs(3104) <= '0';
    layer1_outputs(3105) <= '1';
    layer1_outputs(3106) <= not((layer0_outputs(3254)) and (layer0_outputs(506)));
    layer1_outputs(3107) <= (layer0_outputs(1864)) and (layer0_outputs(3795));
    layer1_outputs(3108) <= (layer0_outputs(7100)) and not (layer0_outputs(5566));
    layer1_outputs(3109) <= '1';
    layer1_outputs(3110) <= not((layer0_outputs(878)) and (layer0_outputs(880)));
    layer1_outputs(3111) <= not((layer0_outputs(6342)) and (layer0_outputs(5699)));
    layer1_outputs(3112) <= (layer0_outputs(5557)) and not (layer0_outputs(4471));
    layer1_outputs(3113) <= layer0_outputs(6630);
    layer1_outputs(3114) <= not(layer0_outputs(7220));
    layer1_outputs(3115) <= '0';
    layer1_outputs(3116) <= layer0_outputs(4477);
    layer1_outputs(3117) <= layer0_outputs(794);
    layer1_outputs(3118) <= not((layer0_outputs(1478)) or (layer0_outputs(5912)));
    layer1_outputs(3119) <= (layer0_outputs(5035)) and (layer0_outputs(4216));
    layer1_outputs(3120) <= '1';
    layer1_outputs(3121) <= (layer0_outputs(3287)) and not (layer0_outputs(6787));
    layer1_outputs(3122) <= (layer0_outputs(4186)) and not (layer0_outputs(3026));
    layer1_outputs(3123) <= not((layer0_outputs(1431)) or (layer0_outputs(3976)));
    layer1_outputs(3124) <= not(layer0_outputs(3770)) or (layer0_outputs(2232));
    layer1_outputs(3125) <= not((layer0_outputs(5230)) or (layer0_outputs(6678)));
    layer1_outputs(3126) <= (layer0_outputs(6048)) and (layer0_outputs(1543));
    layer1_outputs(3127) <= not((layer0_outputs(4947)) and (layer0_outputs(1612)));
    layer1_outputs(3128) <= '0';
    layer1_outputs(3129) <= layer0_outputs(7513);
    layer1_outputs(3130) <= not((layer0_outputs(4588)) and (layer0_outputs(1382)));
    layer1_outputs(3131) <= '0';
    layer1_outputs(3132) <= not((layer0_outputs(6031)) and (layer0_outputs(2478)));
    layer1_outputs(3133) <= layer0_outputs(2550);
    layer1_outputs(3134) <= not((layer0_outputs(3309)) or (layer0_outputs(5801)));
    layer1_outputs(3135) <= layer0_outputs(4804);
    layer1_outputs(3136) <= (layer0_outputs(2957)) and not (layer0_outputs(1975));
    layer1_outputs(3137) <= not(layer0_outputs(650)) or (layer0_outputs(3496));
    layer1_outputs(3138) <= '1';
    layer1_outputs(3139) <= (layer0_outputs(5748)) and (layer0_outputs(955));
    layer1_outputs(3140) <= (layer0_outputs(6306)) and not (layer0_outputs(2582));
    layer1_outputs(3141) <= not((layer0_outputs(1313)) and (layer0_outputs(4618)));
    layer1_outputs(3142) <= not(layer0_outputs(4197)) or (layer0_outputs(5817));
    layer1_outputs(3143) <= (layer0_outputs(3554)) or (layer0_outputs(3803));
    layer1_outputs(3144) <= (layer0_outputs(253)) or (layer0_outputs(6034));
    layer1_outputs(3145) <= not((layer0_outputs(3125)) xor (layer0_outputs(6018)));
    layer1_outputs(3146) <= (layer0_outputs(1200)) or (layer0_outputs(2233));
    layer1_outputs(3147) <= '0';
    layer1_outputs(3148) <= layer0_outputs(316);
    layer1_outputs(3149) <= not(layer0_outputs(559));
    layer1_outputs(3150) <= (layer0_outputs(4100)) and not (layer0_outputs(3588));
    layer1_outputs(3151) <= not(layer0_outputs(7131)) or (layer0_outputs(967));
    layer1_outputs(3152) <= (layer0_outputs(5531)) and not (layer0_outputs(518));
    layer1_outputs(3153) <= (layer0_outputs(4182)) xor (layer0_outputs(2007));
    layer1_outputs(3154) <= not((layer0_outputs(7152)) and (layer0_outputs(4633)));
    layer1_outputs(3155) <= '1';
    layer1_outputs(3156) <= (layer0_outputs(3657)) or (layer0_outputs(3671));
    layer1_outputs(3157) <= not(layer0_outputs(7429)) or (layer0_outputs(6685));
    layer1_outputs(3158) <= layer0_outputs(6003);
    layer1_outputs(3159) <= '1';
    layer1_outputs(3160) <= layer0_outputs(6205);
    layer1_outputs(3161) <= layer0_outputs(1750);
    layer1_outputs(3162) <= layer0_outputs(5849);
    layer1_outputs(3163) <= '0';
    layer1_outputs(3164) <= not(layer0_outputs(424)) or (layer0_outputs(1296));
    layer1_outputs(3165) <= '1';
    layer1_outputs(3166) <= '0';
    layer1_outputs(3167) <= not((layer0_outputs(3454)) or (layer0_outputs(6661)));
    layer1_outputs(3168) <= (layer0_outputs(5973)) or (layer0_outputs(2981));
    layer1_outputs(3169) <= not(layer0_outputs(4745)) or (layer0_outputs(442));
    layer1_outputs(3170) <= '1';
    layer1_outputs(3171) <= layer0_outputs(7050);
    layer1_outputs(3172) <= '1';
    layer1_outputs(3173) <= layer0_outputs(2094);
    layer1_outputs(3174) <= layer0_outputs(2500);
    layer1_outputs(3175) <= layer0_outputs(2372);
    layer1_outputs(3176) <= (layer0_outputs(6853)) and not (layer0_outputs(694));
    layer1_outputs(3177) <= layer0_outputs(406);
    layer1_outputs(3178) <= not((layer0_outputs(333)) and (layer0_outputs(546)));
    layer1_outputs(3179) <= '0';
    layer1_outputs(3180) <= '1';
    layer1_outputs(3181) <= (layer0_outputs(1353)) or (layer0_outputs(3273));
    layer1_outputs(3182) <= not(layer0_outputs(41)) or (layer0_outputs(7267));
    layer1_outputs(3183) <= '0';
    layer1_outputs(3184) <= not(layer0_outputs(1085)) or (layer0_outputs(4680));
    layer1_outputs(3185) <= not(layer0_outputs(3748));
    layer1_outputs(3186) <= (layer0_outputs(6790)) or (layer0_outputs(1722));
    layer1_outputs(3187) <= not(layer0_outputs(821)) or (layer0_outputs(583));
    layer1_outputs(3188) <= '0';
    layer1_outputs(3189) <= '0';
    layer1_outputs(3190) <= not(layer0_outputs(39));
    layer1_outputs(3191) <= (layer0_outputs(6706)) and not (layer0_outputs(3468));
    layer1_outputs(3192) <= '0';
    layer1_outputs(3193) <= not(layer0_outputs(6649)) or (layer0_outputs(4648));
    layer1_outputs(3194) <= layer0_outputs(5888);
    layer1_outputs(3195) <= (layer0_outputs(975)) and not (layer0_outputs(4056));
    layer1_outputs(3196) <= '1';
    layer1_outputs(3197) <= (layer0_outputs(4636)) and not (layer0_outputs(4028));
    layer1_outputs(3198) <= layer0_outputs(604);
    layer1_outputs(3199) <= '0';
    layer1_outputs(3200) <= not(layer0_outputs(6996)) or (layer0_outputs(480));
    layer1_outputs(3201) <= '1';
    layer1_outputs(3202) <= '0';
    layer1_outputs(3203) <= '0';
    layer1_outputs(3204) <= not(layer0_outputs(4856));
    layer1_outputs(3205) <= '0';
    layer1_outputs(3206) <= layer0_outputs(1155);
    layer1_outputs(3207) <= (layer0_outputs(6164)) xor (layer0_outputs(1461));
    layer1_outputs(3208) <= '0';
    layer1_outputs(3209) <= not(layer0_outputs(4655)) or (layer0_outputs(2406));
    layer1_outputs(3210) <= '1';
    layer1_outputs(3211) <= '1';
    layer1_outputs(3212) <= '0';
    layer1_outputs(3213) <= not(layer0_outputs(1498));
    layer1_outputs(3214) <= '0';
    layer1_outputs(3215) <= '1';
    layer1_outputs(3216) <= not(layer0_outputs(1398));
    layer1_outputs(3217) <= '1';
    layer1_outputs(3218) <= not((layer0_outputs(5370)) and (layer0_outputs(5706)));
    layer1_outputs(3219) <= not(layer0_outputs(3138));
    layer1_outputs(3220) <= (layer0_outputs(477)) and (layer0_outputs(3021));
    layer1_outputs(3221) <= (layer0_outputs(1214)) or (layer0_outputs(3171));
    layer1_outputs(3222) <= '1';
    layer1_outputs(3223) <= layer0_outputs(2235);
    layer1_outputs(3224) <= not(layer0_outputs(7036));
    layer1_outputs(3225) <= layer0_outputs(4668);
    layer1_outputs(3226) <= layer0_outputs(6190);
    layer1_outputs(3227) <= not((layer0_outputs(6194)) or (layer0_outputs(520)));
    layer1_outputs(3228) <= not((layer0_outputs(4408)) and (layer0_outputs(6076)));
    layer1_outputs(3229) <= '1';
    layer1_outputs(3230) <= '0';
    layer1_outputs(3231) <= not(layer0_outputs(6280)) or (layer0_outputs(7363));
    layer1_outputs(3232) <= '0';
    layer1_outputs(3233) <= (layer0_outputs(850)) or (layer0_outputs(1765));
    layer1_outputs(3234) <= (layer0_outputs(1500)) and (layer0_outputs(1212));
    layer1_outputs(3235) <= layer0_outputs(3938);
    layer1_outputs(3236) <= not(layer0_outputs(987));
    layer1_outputs(3237) <= (layer0_outputs(5988)) xor (layer0_outputs(4598));
    layer1_outputs(3238) <= (layer0_outputs(3364)) or (layer0_outputs(2003));
    layer1_outputs(3239) <= not((layer0_outputs(1429)) or (layer0_outputs(898)));
    layer1_outputs(3240) <= not((layer0_outputs(953)) or (layer0_outputs(4336)));
    layer1_outputs(3241) <= (layer0_outputs(1271)) or (layer0_outputs(2266));
    layer1_outputs(3242) <= not(layer0_outputs(2140)) or (layer0_outputs(1895));
    layer1_outputs(3243) <= layer0_outputs(136);
    layer1_outputs(3244) <= not(layer0_outputs(2079)) or (layer0_outputs(1631));
    layer1_outputs(3245) <= '0';
    layer1_outputs(3246) <= (layer0_outputs(7183)) or (layer0_outputs(956));
    layer1_outputs(3247) <= not(layer0_outputs(4923)) or (layer0_outputs(1714));
    layer1_outputs(3248) <= layer0_outputs(7125);
    layer1_outputs(3249) <= '1';
    layer1_outputs(3250) <= not(layer0_outputs(5416));
    layer1_outputs(3251) <= layer0_outputs(609);
    layer1_outputs(3252) <= (layer0_outputs(5411)) xor (layer0_outputs(2319));
    layer1_outputs(3253) <= '1';
    layer1_outputs(3254) <= '1';
    layer1_outputs(3255) <= (layer0_outputs(1470)) and not (layer0_outputs(152));
    layer1_outputs(3256) <= (layer0_outputs(1430)) and (layer0_outputs(1855));
    layer1_outputs(3257) <= not(layer0_outputs(801));
    layer1_outputs(3258) <= (layer0_outputs(2461)) and not (layer0_outputs(2101));
    layer1_outputs(3259) <= '0';
    layer1_outputs(3260) <= not(layer0_outputs(3717));
    layer1_outputs(3261) <= not(layer0_outputs(1234)) or (layer0_outputs(7557));
    layer1_outputs(3262) <= '0';
    layer1_outputs(3263) <= (layer0_outputs(2001)) and (layer0_outputs(4732));
    layer1_outputs(3264) <= not(layer0_outputs(7316)) or (layer0_outputs(1762));
    layer1_outputs(3265) <= layer0_outputs(6122);
    layer1_outputs(3266) <= not(layer0_outputs(4252));
    layer1_outputs(3267) <= not(layer0_outputs(937)) or (layer0_outputs(3379));
    layer1_outputs(3268) <= not((layer0_outputs(7065)) or (layer0_outputs(68)));
    layer1_outputs(3269) <= not((layer0_outputs(28)) and (layer0_outputs(4731)));
    layer1_outputs(3270) <= not(layer0_outputs(7231)) or (layer0_outputs(7290));
    layer1_outputs(3271) <= '0';
    layer1_outputs(3272) <= layer0_outputs(5946);
    layer1_outputs(3273) <= '1';
    layer1_outputs(3274) <= not(layer0_outputs(5220));
    layer1_outputs(3275) <= not(layer0_outputs(7224)) or (layer0_outputs(6709));
    layer1_outputs(3276) <= layer0_outputs(5804);
    layer1_outputs(3277) <= '0';
    layer1_outputs(3278) <= not(layer0_outputs(365));
    layer1_outputs(3279) <= '0';
    layer1_outputs(3280) <= (layer0_outputs(4347)) and not (layer0_outputs(3304));
    layer1_outputs(3281) <= (layer0_outputs(4718)) or (layer0_outputs(1820));
    layer1_outputs(3282) <= not(layer0_outputs(3500)) or (layer0_outputs(1789));
    layer1_outputs(3283) <= (layer0_outputs(7035)) and (layer0_outputs(2595));
    layer1_outputs(3284) <= not(layer0_outputs(3174)) or (layer0_outputs(5573));
    layer1_outputs(3285) <= not(layer0_outputs(3397));
    layer1_outputs(3286) <= '0';
    layer1_outputs(3287) <= layer0_outputs(3183);
    layer1_outputs(3288) <= '0';
    layer1_outputs(3289) <= '0';
    layer1_outputs(3290) <= not(layer0_outputs(1234));
    layer1_outputs(3291) <= '1';
    layer1_outputs(3292) <= (layer0_outputs(1501)) and (layer0_outputs(7582));
    layer1_outputs(3293) <= (layer0_outputs(225)) or (layer0_outputs(1850));
    layer1_outputs(3294) <= not((layer0_outputs(706)) and (layer0_outputs(187)));
    layer1_outputs(3295) <= not(layer0_outputs(740));
    layer1_outputs(3296) <= not((layer0_outputs(3300)) and (layer0_outputs(4964)));
    layer1_outputs(3297) <= not((layer0_outputs(5550)) or (layer0_outputs(2485)));
    layer1_outputs(3298) <= not(layer0_outputs(3670)) or (layer0_outputs(3692));
    layer1_outputs(3299) <= '0';
    layer1_outputs(3300) <= (layer0_outputs(657)) and not (layer0_outputs(7626));
    layer1_outputs(3301) <= not((layer0_outputs(1200)) or (layer0_outputs(3415)));
    layer1_outputs(3302) <= not(layer0_outputs(761));
    layer1_outputs(3303) <= (layer0_outputs(3879)) or (layer0_outputs(4817));
    layer1_outputs(3304) <= not(layer0_outputs(2343));
    layer1_outputs(3305) <= layer0_outputs(6946);
    layer1_outputs(3306) <= not(layer0_outputs(1870)) or (layer0_outputs(2387));
    layer1_outputs(3307) <= not(layer0_outputs(6039)) or (layer0_outputs(42));
    layer1_outputs(3308) <= not(layer0_outputs(2609)) or (layer0_outputs(2495));
    layer1_outputs(3309) <= not(layer0_outputs(6100)) or (layer0_outputs(584));
    layer1_outputs(3310) <= not((layer0_outputs(1633)) or (layer0_outputs(6876)));
    layer1_outputs(3311) <= layer0_outputs(1254);
    layer1_outputs(3312) <= '1';
    layer1_outputs(3313) <= not(layer0_outputs(4588)) or (layer0_outputs(6999));
    layer1_outputs(3314) <= (layer0_outputs(6563)) and (layer0_outputs(1006));
    layer1_outputs(3315) <= layer0_outputs(1795);
    layer1_outputs(3316) <= '0';
    layer1_outputs(3317) <= not(layer0_outputs(1174));
    layer1_outputs(3318) <= '1';
    layer1_outputs(3319) <= layer0_outputs(903);
    layer1_outputs(3320) <= '0';
    layer1_outputs(3321) <= not(layer0_outputs(6606));
    layer1_outputs(3322) <= not(layer0_outputs(821)) or (layer0_outputs(5598));
    layer1_outputs(3323) <= '1';
    layer1_outputs(3324) <= not((layer0_outputs(6893)) or (layer0_outputs(3859)));
    layer1_outputs(3325) <= not(layer0_outputs(2129)) or (layer0_outputs(2411));
    layer1_outputs(3326) <= not(layer0_outputs(493)) or (layer0_outputs(7367));
    layer1_outputs(3327) <= (layer0_outputs(1427)) and (layer0_outputs(6177));
    layer1_outputs(3328) <= '0';
    layer1_outputs(3329) <= (layer0_outputs(528)) and (layer0_outputs(9));
    layer1_outputs(3330) <= '0';
    layer1_outputs(3331) <= (layer0_outputs(673)) and not (layer0_outputs(3843));
    layer1_outputs(3332) <= (layer0_outputs(3260)) or (layer0_outputs(4505));
    layer1_outputs(3333) <= not((layer0_outputs(4381)) xor (layer0_outputs(7351)));
    layer1_outputs(3334) <= '0';
    layer1_outputs(3335) <= '0';
    layer1_outputs(3336) <= (layer0_outputs(1219)) and not (layer0_outputs(7408));
    layer1_outputs(3337) <= not(layer0_outputs(950)) or (layer0_outputs(3149));
    layer1_outputs(3338) <= '0';
    layer1_outputs(3339) <= not(layer0_outputs(1198));
    layer1_outputs(3340) <= not((layer0_outputs(1070)) xor (layer0_outputs(5732)));
    layer1_outputs(3341) <= '1';
    layer1_outputs(3342) <= not(layer0_outputs(3728)) or (layer0_outputs(1552));
    layer1_outputs(3343) <= not(layer0_outputs(6090)) or (layer0_outputs(3542));
    layer1_outputs(3344) <= not(layer0_outputs(1080)) or (layer0_outputs(4433));
    layer1_outputs(3345) <= '0';
    layer1_outputs(3346) <= layer0_outputs(1540);
    layer1_outputs(3347) <= not(layer0_outputs(996));
    layer1_outputs(3348) <= layer0_outputs(5044);
    layer1_outputs(3349) <= not((layer0_outputs(4774)) and (layer0_outputs(710)));
    layer1_outputs(3350) <= '1';
    layer1_outputs(3351) <= not((layer0_outputs(5017)) or (layer0_outputs(1441)));
    layer1_outputs(3352) <= not((layer0_outputs(3351)) and (layer0_outputs(7512)));
    layer1_outputs(3353) <= '1';
    layer1_outputs(3354) <= (layer0_outputs(3447)) or (layer0_outputs(5840));
    layer1_outputs(3355) <= not(layer0_outputs(4415));
    layer1_outputs(3356) <= layer0_outputs(4312);
    layer1_outputs(3357) <= (layer0_outputs(4806)) xor (layer0_outputs(2987));
    layer1_outputs(3358) <= layer0_outputs(5359);
    layer1_outputs(3359) <= not(layer0_outputs(6972)) or (layer0_outputs(5180));
    layer1_outputs(3360) <= not((layer0_outputs(6879)) and (layer0_outputs(5704)));
    layer1_outputs(3361) <= layer0_outputs(1471);
    layer1_outputs(3362) <= not((layer0_outputs(2491)) or (layer0_outputs(4843)));
    layer1_outputs(3363) <= (layer0_outputs(4659)) or (layer0_outputs(3955));
    layer1_outputs(3364) <= not(layer0_outputs(5765));
    layer1_outputs(3365) <= not(layer0_outputs(4593));
    layer1_outputs(3366) <= not(layer0_outputs(905));
    layer1_outputs(3367) <= (layer0_outputs(3362)) or (layer0_outputs(5055));
    layer1_outputs(3368) <= not(layer0_outputs(2786));
    layer1_outputs(3369) <= '0';
    layer1_outputs(3370) <= (layer0_outputs(7281)) and not (layer0_outputs(5185));
    layer1_outputs(3371) <= (layer0_outputs(7241)) and not (layer0_outputs(2766));
    layer1_outputs(3372) <= '1';
    layer1_outputs(3373) <= layer0_outputs(357);
    layer1_outputs(3374) <= not(layer0_outputs(2116));
    layer1_outputs(3375) <= layer0_outputs(2442);
    layer1_outputs(3376) <= not(layer0_outputs(3857));
    layer1_outputs(3377) <= not(layer0_outputs(5418));
    layer1_outputs(3378) <= not((layer0_outputs(1685)) xor (layer0_outputs(5027)));
    layer1_outputs(3379) <= not(layer0_outputs(2641));
    layer1_outputs(3380) <= not((layer0_outputs(5077)) or (layer0_outputs(2992)));
    layer1_outputs(3381) <= not(layer0_outputs(6817)) or (layer0_outputs(4338));
    layer1_outputs(3382) <= (layer0_outputs(732)) and not (layer0_outputs(4746));
    layer1_outputs(3383) <= (layer0_outputs(6779)) and not (layer0_outputs(3858));
    layer1_outputs(3384) <= '0';
    layer1_outputs(3385) <= not(layer0_outputs(6229)) or (layer0_outputs(1479));
    layer1_outputs(3386) <= '0';
    layer1_outputs(3387) <= '0';
    layer1_outputs(3388) <= not(layer0_outputs(3124)) or (layer0_outputs(3527));
    layer1_outputs(3389) <= not(layer0_outputs(1058));
    layer1_outputs(3390) <= layer0_outputs(1507);
    layer1_outputs(3391) <= not(layer0_outputs(1086)) or (layer0_outputs(2797));
    layer1_outputs(3392) <= layer0_outputs(2660);
    layer1_outputs(3393) <= not(layer0_outputs(5383));
    layer1_outputs(3394) <= not(layer0_outputs(4610)) or (layer0_outputs(22));
    layer1_outputs(3395) <= not(layer0_outputs(6612)) or (layer0_outputs(485));
    layer1_outputs(3396) <= not(layer0_outputs(5946)) or (layer0_outputs(6699));
    layer1_outputs(3397) <= '1';
    layer1_outputs(3398) <= layer0_outputs(559);
    layer1_outputs(3399) <= not((layer0_outputs(5678)) and (layer0_outputs(7210)));
    layer1_outputs(3400) <= not((layer0_outputs(2215)) or (layer0_outputs(2278)));
    layer1_outputs(3401) <= (layer0_outputs(867)) and not (layer0_outputs(2397));
    layer1_outputs(3402) <= '0';
    layer1_outputs(3403) <= not(layer0_outputs(7645)) or (layer0_outputs(7635));
    layer1_outputs(3404) <= '1';
    layer1_outputs(3405) <= not((layer0_outputs(7668)) or (layer0_outputs(994)));
    layer1_outputs(3406) <= (layer0_outputs(2942)) or (layer0_outputs(3006));
    layer1_outputs(3407) <= not(layer0_outputs(3999)) or (layer0_outputs(1233));
    layer1_outputs(3408) <= '0';
    layer1_outputs(3409) <= (layer0_outputs(58)) or (layer0_outputs(374));
    layer1_outputs(3410) <= (layer0_outputs(6368)) and not (layer0_outputs(6214));
    layer1_outputs(3411) <= not(layer0_outputs(4931)) or (layer0_outputs(4785));
    layer1_outputs(3412) <= '0';
    layer1_outputs(3413) <= (layer0_outputs(4177)) and not (layer0_outputs(637));
    layer1_outputs(3414) <= (layer0_outputs(3940)) xor (layer0_outputs(6016));
    layer1_outputs(3415) <= (layer0_outputs(7210)) and not (layer0_outputs(5988));
    layer1_outputs(3416) <= not((layer0_outputs(5609)) xor (layer0_outputs(5779)));
    layer1_outputs(3417) <= '1';
    layer1_outputs(3418) <= (layer0_outputs(643)) and not (layer0_outputs(5112));
    layer1_outputs(3419) <= '0';
    layer1_outputs(3420) <= (layer0_outputs(280)) xor (layer0_outputs(1626));
    layer1_outputs(3421) <= (layer0_outputs(6120)) and (layer0_outputs(394));
    layer1_outputs(3422) <= not(layer0_outputs(2156)) or (layer0_outputs(7592));
    layer1_outputs(3423) <= not(layer0_outputs(3412)) or (layer0_outputs(5098));
    layer1_outputs(3424) <= layer0_outputs(1548);
    layer1_outputs(3425) <= not((layer0_outputs(1852)) and (layer0_outputs(3154)));
    layer1_outputs(3426) <= '0';
    layer1_outputs(3427) <= (layer0_outputs(1800)) and not (layer0_outputs(3386));
    layer1_outputs(3428) <= not(layer0_outputs(3091)) or (layer0_outputs(356));
    layer1_outputs(3429) <= (layer0_outputs(1543)) or (layer0_outputs(4072));
    layer1_outputs(3430) <= (layer0_outputs(5028)) xor (layer0_outputs(7201));
    layer1_outputs(3431) <= '0';
    layer1_outputs(3432) <= (layer0_outputs(6502)) and not (layer0_outputs(1391));
    layer1_outputs(3433) <= not((layer0_outputs(5936)) and (layer0_outputs(1876)));
    layer1_outputs(3434) <= layer0_outputs(6658);
    layer1_outputs(3435) <= (layer0_outputs(4082)) and (layer0_outputs(5549));
    layer1_outputs(3436) <= not(layer0_outputs(6105));
    layer1_outputs(3437) <= (layer0_outputs(4406)) or (layer0_outputs(7355));
    layer1_outputs(3438) <= not(layer0_outputs(6943));
    layer1_outputs(3439) <= not(layer0_outputs(4858)) or (layer0_outputs(2384));
    layer1_outputs(3440) <= layer0_outputs(6226);
    layer1_outputs(3441) <= (layer0_outputs(1933)) and (layer0_outputs(5224));
    layer1_outputs(3442) <= not(layer0_outputs(1166));
    layer1_outputs(3443) <= (layer0_outputs(3764)) xor (layer0_outputs(468));
    layer1_outputs(3444) <= '1';
    layer1_outputs(3445) <= (layer0_outputs(5808)) or (layer0_outputs(6223));
    layer1_outputs(3446) <= not(layer0_outputs(5163));
    layer1_outputs(3447) <= not(layer0_outputs(3074)) or (layer0_outputs(5463));
    layer1_outputs(3448) <= not((layer0_outputs(6966)) and (layer0_outputs(2793)));
    layer1_outputs(3449) <= not(layer0_outputs(6283)) or (layer0_outputs(7174));
    layer1_outputs(3450) <= not((layer0_outputs(4097)) or (layer0_outputs(4877)));
    layer1_outputs(3451) <= '0';
    layer1_outputs(3452) <= '0';
    layer1_outputs(3453) <= '1';
    layer1_outputs(3454) <= layer0_outputs(5377);
    layer1_outputs(3455) <= layer0_outputs(4949);
    layer1_outputs(3456) <= (layer0_outputs(4096)) and not (layer0_outputs(4587));
    layer1_outputs(3457) <= (layer0_outputs(6530)) and not (layer0_outputs(2455));
    layer1_outputs(3458) <= '1';
    layer1_outputs(3459) <= layer0_outputs(599);
    layer1_outputs(3460) <= not(layer0_outputs(1448)) or (layer0_outputs(1320));
    layer1_outputs(3461) <= (layer0_outputs(513)) and (layer0_outputs(7248));
    layer1_outputs(3462) <= not((layer0_outputs(2332)) xor (layer0_outputs(1992)));
    layer1_outputs(3463) <= (layer0_outputs(1644)) or (layer0_outputs(4751));
    layer1_outputs(3464) <= '0';
    layer1_outputs(3465) <= not((layer0_outputs(1944)) and (layer0_outputs(6720)));
    layer1_outputs(3466) <= layer0_outputs(1702);
    layer1_outputs(3467) <= '0';
    layer1_outputs(3468) <= (layer0_outputs(5753)) and not (layer0_outputs(7332));
    layer1_outputs(3469) <= not(layer0_outputs(6143));
    layer1_outputs(3470) <= layer0_outputs(880);
    layer1_outputs(3471) <= layer0_outputs(3621);
    layer1_outputs(3472) <= not(layer0_outputs(4693)) or (layer0_outputs(4360));
    layer1_outputs(3473) <= '0';
    layer1_outputs(3474) <= not(layer0_outputs(4854));
    layer1_outputs(3475) <= layer0_outputs(460);
    layer1_outputs(3476) <= (layer0_outputs(4199)) and not (layer0_outputs(6307));
    layer1_outputs(3477) <= (layer0_outputs(798)) or (layer0_outputs(6547));
    layer1_outputs(3478) <= layer0_outputs(7510);
    layer1_outputs(3479) <= '0';
    layer1_outputs(3480) <= not(layer0_outputs(5011));
    layer1_outputs(3481) <= layer0_outputs(4784);
    layer1_outputs(3482) <= not(layer0_outputs(4130));
    layer1_outputs(3483) <= '0';
    layer1_outputs(3484) <= not((layer0_outputs(4579)) or (layer0_outputs(2230)));
    layer1_outputs(3485) <= layer0_outputs(890);
    layer1_outputs(3486) <= not(layer0_outputs(937)) or (layer0_outputs(5662));
    layer1_outputs(3487) <= layer0_outputs(6725);
    layer1_outputs(3488) <= (layer0_outputs(5891)) and (layer0_outputs(3487));
    layer1_outputs(3489) <= (layer0_outputs(5949)) and (layer0_outputs(222));
    layer1_outputs(3490) <= not((layer0_outputs(5036)) or (layer0_outputs(997)));
    layer1_outputs(3491) <= '1';
    layer1_outputs(3492) <= not((layer0_outputs(5104)) or (layer0_outputs(2990)));
    layer1_outputs(3493) <= '0';
    layer1_outputs(3494) <= '0';
    layer1_outputs(3495) <= (layer0_outputs(6397)) or (layer0_outputs(3646));
    layer1_outputs(3496) <= not(layer0_outputs(5666));
    layer1_outputs(3497) <= not(layer0_outputs(5605));
    layer1_outputs(3498) <= (layer0_outputs(2974)) and not (layer0_outputs(2212));
    layer1_outputs(3499) <= layer0_outputs(7165);
    layer1_outputs(3500) <= '0';
    layer1_outputs(3501) <= not(layer0_outputs(7439));
    layer1_outputs(3502) <= layer0_outputs(1499);
    layer1_outputs(3503) <= (layer0_outputs(4884)) and (layer0_outputs(4878));
    layer1_outputs(3504) <= '0';
    layer1_outputs(3505) <= (layer0_outputs(5554)) or (layer0_outputs(6721));
    layer1_outputs(3506) <= not((layer0_outputs(6675)) xor (layer0_outputs(3196)));
    layer1_outputs(3507) <= (layer0_outputs(2000)) and not (layer0_outputs(735));
    layer1_outputs(3508) <= (layer0_outputs(1797)) or (layer0_outputs(2955));
    layer1_outputs(3509) <= not(layer0_outputs(5066));
    layer1_outputs(3510) <= '0';
    layer1_outputs(3511) <= (layer0_outputs(6633)) and not (layer0_outputs(7374));
    layer1_outputs(3512) <= not(layer0_outputs(2290)) or (layer0_outputs(6836));
    layer1_outputs(3513) <= (layer0_outputs(509)) or (layer0_outputs(7430));
    layer1_outputs(3514) <= (layer0_outputs(7230)) or (layer0_outputs(6087));
    layer1_outputs(3515) <= not(layer0_outputs(6066)) or (layer0_outputs(803));
    layer1_outputs(3516) <= not(layer0_outputs(788)) or (layer0_outputs(969));
    layer1_outputs(3517) <= (layer0_outputs(6)) and not (layer0_outputs(1410));
    layer1_outputs(3518) <= '0';
    layer1_outputs(3519) <= not((layer0_outputs(6000)) and (layer0_outputs(5070)));
    layer1_outputs(3520) <= (layer0_outputs(3579)) and not (layer0_outputs(2334));
    layer1_outputs(3521) <= layer0_outputs(6911);
    layer1_outputs(3522) <= '1';
    layer1_outputs(3523) <= '0';
    layer1_outputs(3524) <= not((layer0_outputs(2808)) and (layer0_outputs(5379)));
    layer1_outputs(3525) <= not(layer0_outputs(3969));
    layer1_outputs(3526) <= (layer0_outputs(4640)) or (layer0_outputs(3381));
    layer1_outputs(3527) <= (layer0_outputs(326)) and not (layer0_outputs(1172));
    layer1_outputs(3528) <= (layer0_outputs(4341)) or (layer0_outputs(2977));
    layer1_outputs(3529) <= not(layer0_outputs(5960));
    layer1_outputs(3530) <= (layer0_outputs(7494)) or (layer0_outputs(5708));
    layer1_outputs(3531) <= layer0_outputs(4815);
    layer1_outputs(3532) <= layer0_outputs(3912);
    layer1_outputs(3533) <= (layer0_outputs(4255)) and (layer0_outputs(5084));
    layer1_outputs(3534) <= not((layer0_outputs(1083)) or (layer0_outputs(4586)));
    layer1_outputs(3535) <= not(layer0_outputs(424)) or (layer0_outputs(2413));
    layer1_outputs(3536) <= (layer0_outputs(7577)) and not (layer0_outputs(4444));
    layer1_outputs(3537) <= not(layer0_outputs(3560)) or (layer0_outputs(1089));
    layer1_outputs(3538) <= not((layer0_outputs(6655)) and (layer0_outputs(1459)));
    layer1_outputs(3539) <= not((layer0_outputs(2904)) or (layer0_outputs(3844)));
    layer1_outputs(3540) <= not(layer0_outputs(6581)) or (layer0_outputs(2897));
    layer1_outputs(3541) <= not(layer0_outputs(577));
    layer1_outputs(3542) <= layer0_outputs(1523);
    layer1_outputs(3543) <= not((layer0_outputs(6931)) and (layer0_outputs(6499)));
    layer1_outputs(3544) <= (layer0_outputs(3262)) or (layer0_outputs(2561));
    layer1_outputs(3545) <= not(layer0_outputs(2421));
    layer1_outputs(3546) <= (layer0_outputs(1989)) and (layer0_outputs(4683));
    layer1_outputs(3547) <= not((layer0_outputs(610)) or (layer0_outputs(5131)));
    layer1_outputs(3548) <= (layer0_outputs(4102)) or (layer0_outputs(7512));
    layer1_outputs(3549) <= '0';
    layer1_outputs(3550) <= not((layer0_outputs(1758)) or (layer0_outputs(2121)));
    layer1_outputs(3551) <= layer0_outputs(3100);
    layer1_outputs(3552) <= not(layer0_outputs(6684)) or (layer0_outputs(7150));
    layer1_outputs(3553) <= not(layer0_outputs(5716)) or (layer0_outputs(1201));
    layer1_outputs(3554) <= not(layer0_outputs(313)) or (layer0_outputs(2521));
    layer1_outputs(3555) <= not(layer0_outputs(7490));
    layer1_outputs(3556) <= not(layer0_outputs(6357));
    layer1_outputs(3557) <= not(layer0_outputs(3102)) or (layer0_outputs(4865));
    layer1_outputs(3558) <= not(layer0_outputs(7070));
    layer1_outputs(3559) <= layer0_outputs(4703);
    layer1_outputs(3560) <= (layer0_outputs(2460)) or (layer0_outputs(3441));
    layer1_outputs(3561) <= layer0_outputs(4992);
    layer1_outputs(3562) <= (layer0_outputs(5737)) and not (layer0_outputs(6458));
    layer1_outputs(3563) <= not((layer0_outputs(17)) and (layer0_outputs(6001)));
    layer1_outputs(3564) <= layer0_outputs(4519);
    layer1_outputs(3565) <= '1';
    layer1_outputs(3566) <= '1';
    layer1_outputs(3567) <= not((layer0_outputs(7330)) or (layer0_outputs(1210)));
    layer1_outputs(3568) <= layer0_outputs(4399);
    layer1_outputs(3569) <= not(layer0_outputs(6922)) or (layer0_outputs(2638));
    layer1_outputs(3570) <= layer0_outputs(6465);
    layer1_outputs(3571) <= not(layer0_outputs(3133));
    layer1_outputs(3572) <= (layer0_outputs(1434)) and not (layer0_outputs(315));
    layer1_outputs(3573) <= not(layer0_outputs(6207)) or (layer0_outputs(7020));
    layer1_outputs(3574) <= not((layer0_outputs(2915)) or (layer0_outputs(2029)));
    layer1_outputs(3575) <= (layer0_outputs(3290)) or (layer0_outputs(4940));
    layer1_outputs(3576) <= layer0_outputs(3896);
    layer1_outputs(3577) <= not(layer0_outputs(2322));
    layer1_outputs(3578) <= layer0_outputs(2304);
    layer1_outputs(3579) <= '1';
    layer1_outputs(3580) <= (layer0_outputs(5927)) and (layer0_outputs(7660));
    layer1_outputs(3581) <= not(layer0_outputs(102));
    layer1_outputs(3582) <= layer0_outputs(753);
    layer1_outputs(3583) <= (layer0_outputs(2614)) and not (layer0_outputs(43));
    layer1_outputs(3584) <= not((layer0_outputs(4011)) and (layer0_outputs(1986)));
    layer1_outputs(3585) <= not((layer0_outputs(1978)) xor (layer0_outputs(5024)));
    layer1_outputs(3586) <= layer0_outputs(667);
    layer1_outputs(3587) <= (layer0_outputs(272)) and (layer0_outputs(4618));
    layer1_outputs(3588) <= not(layer0_outputs(1580));
    layer1_outputs(3589) <= not(layer0_outputs(5618));
    layer1_outputs(3590) <= '1';
    layer1_outputs(3591) <= (layer0_outputs(893)) and not (layer0_outputs(6962));
    layer1_outputs(3592) <= layer0_outputs(4326);
    layer1_outputs(3593) <= not((layer0_outputs(4332)) and (layer0_outputs(7130)));
    layer1_outputs(3594) <= not(layer0_outputs(5484)) or (layer0_outputs(3170));
    layer1_outputs(3595) <= '0';
    layer1_outputs(3596) <= not((layer0_outputs(7320)) or (layer0_outputs(7179)));
    layer1_outputs(3597) <= not(layer0_outputs(3733));
    layer1_outputs(3598) <= '1';
    layer1_outputs(3599) <= not(layer0_outputs(7245));
    layer1_outputs(3600) <= layer0_outputs(4941);
    layer1_outputs(3601) <= '1';
    layer1_outputs(3602) <= not(layer0_outputs(6505)) or (layer0_outputs(5973));
    layer1_outputs(3603) <= layer0_outputs(4991);
    layer1_outputs(3604) <= '0';
    layer1_outputs(3605) <= (layer0_outputs(6529)) and (layer0_outputs(5400));
    layer1_outputs(3606) <= layer0_outputs(6591);
    layer1_outputs(3607) <= not((layer0_outputs(5767)) and (layer0_outputs(6203)));
    layer1_outputs(3608) <= '1';
    layer1_outputs(3609) <= (layer0_outputs(6264)) or (layer0_outputs(1806));
    layer1_outputs(3610) <= not(layer0_outputs(5937));
    layer1_outputs(3611) <= not(layer0_outputs(2606));
    layer1_outputs(3612) <= not(layer0_outputs(5800)) or (layer0_outputs(6702));
    layer1_outputs(3613) <= '1';
    layer1_outputs(3614) <= not(layer0_outputs(3914));
    layer1_outputs(3615) <= (layer0_outputs(3105)) and not (layer0_outputs(32));
    layer1_outputs(3616) <= not(layer0_outputs(4366)) or (layer0_outputs(1492));
    layer1_outputs(3617) <= not(layer0_outputs(4979));
    layer1_outputs(3618) <= not((layer0_outputs(5775)) or (layer0_outputs(6900)));
    layer1_outputs(3619) <= layer0_outputs(6212);
    layer1_outputs(3620) <= not((layer0_outputs(7566)) or (layer0_outputs(6568)));
    layer1_outputs(3621) <= '0';
    layer1_outputs(3622) <= not(layer0_outputs(4677));
    layer1_outputs(3623) <= not(layer0_outputs(7403)) or (layer0_outputs(3756));
    layer1_outputs(3624) <= (layer0_outputs(6086)) and not (layer0_outputs(1450));
    layer1_outputs(3625) <= not((layer0_outputs(6995)) and (layer0_outputs(7429)));
    layer1_outputs(3626) <= not((layer0_outputs(1919)) or (layer0_outputs(1533)));
    layer1_outputs(3627) <= layer0_outputs(5158);
    layer1_outputs(3628) <= (layer0_outputs(7043)) or (layer0_outputs(230));
    layer1_outputs(3629) <= not((layer0_outputs(5981)) and (layer0_outputs(1689)));
    layer1_outputs(3630) <= '1';
    layer1_outputs(3631) <= layer0_outputs(2199);
    layer1_outputs(3632) <= layer0_outputs(6260);
    layer1_outputs(3633) <= (layer0_outputs(3184)) or (layer0_outputs(7316));
    layer1_outputs(3634) <= not((layer0_outputs(3315)) and (layer0_outputs(6887)));
    layer1_outputs(3635) <= not((layer0_outputs(709)) and (layer0_outputs(2927)));
    layer1_outputs(3636) <= '1';
    layer1_outputs(3637) <= (layer0_outputs(3688)) and not (layer0_outputs(683));
    layer1_outputs(3638) <= layer0_outputs(781);
    layer1_outputs(3639) <= not(layer0_outputs(2288));
    layer1_outputs(3640) <= not(layer0_outputs(4507)) or (layer0_outputs(1110));
    layer1_outputs(3641) <= not(layer0_outputs(5222));
    layer1_outputs(3642) <= (layer0_outputs(3191)) and (layer0_outputs(7638));
    layer1_outputs(3643) <= not(layer0_outputs(4134));
    layer1_outputs(3644) <= '1';
    layer1_outputs(3645) <= (layer0_outputs(85)) and (layer0_outputs(7567));
    layer1_outputs(3646) <= not(layer0_outputs(4013));
    layer1_outputs(3647) <= not(layer0_outputs(219));
    layer1_outputs(3648) <= (layer0_outputs(4420)) and not (layer0_outputs(3269));
    layer1_outputs(3649) <= not((layer0_outputs(5934)) and (layer0_outputs(3986)));
    layer1_outputs(3650) <= not(layer0_outputs(3570)) or (layer0_outputs(1961));
    layer1_outputs(3651) <= not((layer0_outputs(6225)) and (layer0_outputs(1)));
    layer1_outputs(3652) <= (layer0_outputs(1810)) or (layer0_outputs(3166));
    layer1_outputs(3653) <= (layer0_outputs(3354)) or (layer0_outputs(75));
    layer1_outputs(3654) <= not((layer0_outputs(3451)) and (layer0_outputs(6006)));
    layer1_outputs(3655) <= layer0_outputs(5758);
    layer1_outputs(3656) <= (layer0_outputs(693)) and not (layer0_outputs(5486));
    layer1_outputs(3657) <= not(layer0_outputs(4282)) or (layer0_outputs(4869));
    layer1_outputs(3658) <= layer0_outputs(3930);
    layer1_outputs(3659) <= layer0_outputs(6498);
    layer1_outputs(3660) <= not(layer0_outputs(655));
    layer1_outputs(3661) <= not(layer0_outputs(3060));
    layer1_outputs(3662) <= (layer0_outputs(7571)) and not (layer0_outputs(6926));
    layer1_outputs(3663) <= not((layer0_outputs(484)) and (layer0_outputs(4927)));
    layer1_outputs(3664) <= (layer0_outputs(7411)) and (layer0_outputs(6753));
    layer1_outputs(3665) <= (layer0_outputs(5715)) and not (layer0_outputs(3259));
    layer1_outputs(3666) <= not(layer0_outputs(1455)) or (layer0_outputs(2568));
    layer1_outputs(3667) <= not((layer0_outputs(4367)) or (layer0_outputs(1704)));
    layer1_outputs(3668) <= '1';
    layer1_outputs(3669) <= not(layer0_outputs(2335)) or (layer0_outputs(1584));
    layer1_outputs(3670) <= layer0_outputs(6678);
    layer1_outputs(3671) <= '1';
    layer1_outputs(3672) <= not(layer0_outputs(1920));
    layer1_outputs(3673) <= '0';
    layer1_outputs(3674) <= '1';
    layer1_outputs(3675) <= layer0_outputs(3261);
    layer1_outputs(3676) <= (layer0_outputs(5305)) and (layer0_outputs(4595));
    layer1_outputs(3677) <= not((layer0_outputs(3752)) or (layer0_outputs(4900)));
    layer1_outputs(3678) <= (layer0_outputs(7657)) and not (layer0_outputs(930));
    layer1_outputs(3679) <= not(layer0_outputs(806)) or (layer0_outputs(1162));
    layer1_outputs(3680) <= not(layer0_outputs(7263)) or (layer0_outputs(3811));
    layer1_outputs(3681) <= (layer0_outputs(7612)) and (layer0_outputs(7016));
    layer1_outputs(3682) <= layer0_outputs(5713);
    layer1_outputs(3683) <= '1';
    layer1_outputs(3684) <= not(layer0_outputs(3778)) or (layer0_outputs(3021));
    layer1_outputs(3685) <= not(layer0_outputs(6665));
    layer1_outputs(3686) <= '0';
    layer1_outputs(3687) <= '1';
    layer1_outputs(3688) <= (layer0_outputs(4299)) and (layer0_outputs(4448));
    layer1_outputs(3689) <= layer0_outputs(1990);
    layer1_outputs(3690) <= not(layer0_outputs(7647));
    layer1_outputs(3691) <= layer0_outputs(1527);
    layer1_outputs(3692) <= layer0_outputs(5226);
    layer1_outputs(3693) <= (layer0_outputs(6970)) and not (layer0_outputs(4985));
    layer1_outputs(3694) <= not(layer0_outputs(1019)) or (layer0_outputs(2238));
    layer1_outputs(3695) <= '0';
    layer1_outputs(3696) <= not((layer0_outputs(7646)) xor (layer0_outputs(2694)));
    layer1_outputs(3697) <= not(layer0_outputs(7436));
    layer1_outputs(3698) <= '1';
    layer1_outputs(3699) <= layer0_outputs(4600);
    layer1_outputs(3700) <= (layer0_outputs(5055)) or (layer0_outputs(3690));
    layer1_outputs(3701) <= (layer0_outputs(5726)) and not (layer0_outputs(3356));
    layer1_outputs(3702) <= layer0_outputs(4390);
    layer1_outputs(3703) <= (layer0_outputs(7014)) and (layer0_outputs(499));
    layer1_outputs(3704) <= not((layer0_outputs(1919)) or (layer0_outputs(5575)));
    layer1_outputs(3705) <= not(layer0_outputs(6815)) or (layer0_outputs(4829));
    layer1_outputs(3706) <= not((layer0_outputs(6185)) and (layer0_outputs(4819)));
    layer1_outputs(3707) <= (layer0_outputs(1097)) or (layer0_outputs(4392));
    layer1_outputs(3708) <= layer0_outputs(5537);
    layer1_outputs(3709) <= layer0_outputs(4707);
    layer1_outputs(3710) <= '0';
    layer1_outputs(3711) <= '1';
    layer1_outputs(3712) <= not(layer0_outputs(3295));
    layer1_outputs(3713) <= layer0_outputs(397);
    layer1_outputs(3714) <= (layer0_outputs(2484)) and not (layer0_outputs(4207));
    layer1_outputs(3715) <= not(layer0_outputs(7671)) or (layer0_outputs(5773));
    layer1_outputs(3716) <= not((layer0_outputs(3933)) and (layer0_outputs(700)));
    layer1_outputs(3717) <= not(layer0_outputs(299)) or (layer0_outputs(5324));
    layer1_outputs(3718) <= (layer0_outputs(4559)) and (layer0_outputs(6057));
    layer1_outputs(3719) <= not(layer0_outputs(5162)) or (layer0_outputs(6144));
    layer1_outputs(3720) <= (layer0_outputs(3253)) and not (layer0_outputs(2287));
    layer1_outputs(3721) <= not(layer0_outputs(917)) or (layer0_outputs(5675));
    layer1_outputs(3722) <= (layer0_outputs(946)) and not (layer0_outputs(5576));
    layer1_outputs(3723) <= (layer0_outputs(1060)) and not (layer0_outputs(3608));
    layer1_outputs(3724) <= (layer0_outputs(6467)) and not (layer0_outputs(822));
    layer1_outputs(3725) <= '0';
    layer1_outputs(3726) <= '1';
    layer1_outputs(3727) <= not((layer0_outputs(1311)) xor (layer0_outputs(2894)));
    layer1_outputs(3728) <= not(layer0_outputs(1843)) or (layer0_outputs(4047));
    layer1_outputs(3729) <= not(layer0_outputs(6802)) or (layer0_outputs(890));
    layer1_outputs(3730) <= not(layer0_outputs(309)) or (layer0_outputs(4660));
    layer1_outputs(3731) <= layer0_outputs(5125);
    layer1_outputs(3732) <= layer0_outputs(5353);
    layer1_outputs(3733) <= layer0_outputs(1176);
    layer1_outputs(3734) <= layer0_outputs(1292);
    layer1_outputs(3735) <= '0';
    layer1_outputs(3736) <= (layer0_outputs(2398)) and (layer0_outputs(3623));
    layer1_outputs(3737) <= (layer0_outputs(1345)) and not (layer0_outputs(2503));
    layer1_outputs(3738) <= not(layer0_outputs(6146)) or (layer0_outputs(750));
    layer1_outputs(3739) <= not(layer0_outputs(1283)) or (layer0_outputs(3447));
    layer1_outputs(3740) <= (layer0_outputs(5497)) xor (layer0_outputs(5040));
    layer1_outputs(3741) <= '0';
    layer1_outputs(3742) <= (layer0_outputs(3611)) xor (layer0_outputs(95));
    layer1_outputs(3743) <= (layer0_outputs(5787)) and not (layer0_outputs(5971));
    layer1_outputs(3744) <= (layer0_outputs(3323)) and not (layer0_outputs(2459));
    layer1_outputs(3745) <= layer0_outputs(4259);
    layer1_outputs(3746) <= layer0_outputs(6509);
    layer1_outputs(3747) <= (layer0_outputs(2463)) and not (layer0_outputs(2211));
    layer1_outputs(3748) <= not(layer0_outputs(2886));
    layer1_outputs(3749) <= not(layer0_outputs(1623));
    layer1_outputs(3750) <= '1';
    layer1_outputs(3751) <= (layer0_outputs(2723)) and (layer0_outputs(5243));
    layer1_outputs(3752) <= not((layer0_outputs(4855)) and (layer0_outputs(5066)));
    layer1_outputs(3753) <= not((layer0_outputs(5715)) and (layer0_outputs(1981)));
    layer1_outputs(3754) <= not(layer0_outputs(1081)) or (layer0_outputs(7304));
    layer1_outputs(3755) <= not((layer0_outputs(6204)) and (layer0_outputs(7462)));
    layer1_outputs(3756) <= (layer0_outputs(7251)) or (layer0_outputs(1168));
    layer1_outputs(3757) <= layer0_outputs(2649);
    layer1_outputs(3758) <= layer0_outputs(5083);
    layer1_outputs(3759) <= not((layer0_outputs(72)) and (layer0_outputs(3191)));
    layer1_outputs(3760) <= layer0_outputs(5191);
    layer1_outputs(3761) <= not(layer0_outputs(4829));
    layer1_outputs(3762) <= '1';
    layer1_outputs(3763) <= layer0_outputs(6459);
    layer1_outputs(3764) <= layer0_outputs(3767);
    layer1_outputs(3765) <= '0';
    layer1_outputs(3766) <= not((layer0_outputs(3301)) and (layer0_outputs(5649)));
    layer1_outputs(3767) <= layer0_outputs(2952);
    layer1_outputs(3768) <= '1';
    layer1_outputs(3769) <= not(layer0_outputs(257));
    layer1_outputs(3770) <= not(layer0_outputs(5347));
    layer1_outputs(3771) <= '0';
    layer1_outputs(3772) <= '1';
    layer1_outputs(3773) <= not((layer0_outputs(642)) and (layer0_outputs(3765)));
    layer1_outputs(3774) <= (layer0_outputs(66)) and not (layer0_outputs(3361));
    layer1_outputs(3775) <= layer0_outputs(5672);
    layer1_outputs(3776) <= layer0_outputs(5843);
    layer1_outputs(3777) <= layer0_outputs(4488);
    layer1_outputs(3778) <= (layer0_outputs(4704)) and not (layer0_outputs(6226));
    layer1_outputs(3779) <= (layer0_outputs(1617)) or (layer0_outputs(1983));
    layer1_outputs(3780) <= not((layer0_outputs(6595)) and (layer0_outputs(5366)));
    layer1_outputs(3781) <= '1';
    layer1_outputs(3782) <= layer0_outputs(169);
    layer1_outputs(3783) <= not((layer0_outputs(7537)) or (layer0_outputs(2643)));
    layer1_outputs(3784) <= (layer0_outputs(4336)) or (layer0_outputs(3643));
    layer1_outputs(3785) <= '0';
    layer1_outputs(3786) <= (layer0_outputs(4087)) and not (layer0_outputs(7326));
    layer1_outputs(3787) <= '1';
    layer1_outputs(3788) <= not(layer0_outputs(4016));
    layer1_outputs(3789) <= not(layer0_outputs(5140));
    layer1_outputs(3790) <= (layer0_outputs(703)) or (layer0_outputs(5739));
    layer1_outputs(3791) <= not(layer0_outputs(662)) or (layer0_outputs(2570));
    layer1_outputs(3792) <= not(layer0_outputs(624));
    layer1_outputs(3793) <= (layer0_outputs(7259)) and not (layer0_outputs(3003));
    layer1_outputs(3794) <= '0';
    layer1_outputs(3795) <= not(layer0_outputs(1795)) or (layer0_outputs(5126));
    layer1_outputs(3796) <= (layer0_outputs(5473)) and (layer0_outputs(2505));
    layer1_outputs(3797) <= not(layer0_outputs(421)) or (layer0_outputs(3506));
    layer1_outputs(3798) <= (layer0_outputs(4606)) and not (layer0_outputs(2894));
    layer1_outputs(3799) <= (layer0_outputs(5949)) and not (layer0_outputs(959));
    layer1_outputs(3800) <= '0';
    layer1_outputs(3801) <= not((layer0_outputs(648)) xor (layer0_outputs(2806)));
    layer1_outputs(3802) <= not((layer0_outputs(4308)) or (layer0_outputs(46)));
    layer1_outputs(3803) <= '0';
    layer1_outputs(3804) <= not((layer0_outputs(1888)) and (layer0_outputs(4045)));
    layer1_outputs(3805) <= not(layer0_outputs(868)) or (layer0_outputs(1038));
    layer1_outputs(3806) <= not((layer0_outputs(5232)) and (layer0_outputs(6676)));
    layer1_outputs(3807) <= not(layer0_outputs(6691)) or (layer0_outputs(6812));
    layer1_outputs(3808) <= not(layer0_outputs(3299));
    layer1_outputs(3809) <= (layer0_outputs(257)) or (layer0_outputs(3950));
    layer1_outputs(3810) <= '0';
    layer1_outputs(3811) <= (layer0_outputs(4450)) and not (layer0_outputs(833));
    layer1_outputs(3812) <= (layer0_outputs(1782)) and not (layer0_outputs(6043));
    layer1_outputs(3813) <= layer0_outputs(795);
    layer1_outputs(3814) <= (layer0_outputs(749)) and not (layer0_outputs(4594));
    layer1_outputs(3815) <= (layer0_outputs(1976)) and (layer0_outputs(6393));
    layer1_outputs(3816) <= not(layer0_outputs(6902));
    layer1_outputs(3817) <= (layer0_outputs(4742)) or (layer0_outputs(4466));
    layer1_outputs(3818) <= '0';
    layer1_outputs(3819) <= (layer0_outputs(6109)) and not (layer0_outputs(549));
    layer1_outputs(3820) <= layer0_outputs(5037);
    layer1_outputs(3821) <= layer0_outputs(4798);
    layer1_outputs(3822) <= '0';
    layer1_outputs(3823) <= not(layer0_outputs(3594)) or (layer0_outputs(5794));
    layer1_outputs(3824) <= (layer0_outputs(3664)) or (layer0_outputs(7360));
    layer1_outputs(3825) <= (layer0_outputs(873)) and not (layer0_outputs(674));
    layer1_outputs(3826) <= (layer0_outputs(579)) and not (layer0_outputs(4917));
    layer1_outputs(3827) <= not(layer0_outputs(2477));
    layer1_outputs(3828) <= '1';
    layer1_outputs(3829) <= not(layer0_outputs(6379));
    layer1_outputs(3830) <= layer0_outputs(4175);
    layer1_outputs(3831) <= layer0_outputs(3784);
    layer1_outputs(3832) <= '1';
    layer1_outputs(3833) <= (layer0_outputs(1074)) and not (layer0_outputs(7418));
    layer1_outputs(3834) <= (layer0_outputs(4372)) and not (layer0_outputs(4356));
    layer1_outputs(3835) <= (layer0_outputs(2345)) and not (layer0_outputs(2911));
    layer1_outputs(3836) <= not((layer0_outputs(3801)) xor (layer0_outputs(2073)));
    layer1_outputs(3837) <= not((layer0_outputs(4895)) or (layer0_outputs(6383)));
    layer1_outputs(3838) <= not((layer0_outputs(3714)) or (layer0_outputs(1718)));
    layer1_outputs(3839) <= (layer0_outputs(1686)) and (layer0_outputs(4924));
    layer1_outputs(3840) <= '1';
    layer1_outputs(3841) <= '0';
    layer1_outputs(3842) <= not(layer0_outputs(7522)) or (layer0_outputs(3770));
    layer1_outputs(3843) <= not(layer0_outputs(7384));
    layer1_outputs(3844) <= not(layer0_outputs(4397));
    layer1_outputs(3845) <= not(layer0_outputs(5205)) or (layer0_outputs(342));
    layer1_outputs(3846) <= layer0_outputs(5755);
    layer1_outputs(3847) <= layer0_outputs(296);
    layer1_outputs(3848) <= '1';
    layer1_outputs(3849) <= (layer0_outputs(2672)) xor (layer0_outputs(6701));
    layer1_outputs(3850) <= layer0_outputs(4564);
    layer1_outputs(3851) <= '0';
    layer1_outputs(3852) <= not((layer0_outputs(3515)) and (layer0_outputs(7102)));
    layer1_outputs(3853) <= '0';
    layer1_outputs(3854) <= layer0_outputs(4561);
    layer1_outputs(3855) <= not(layer0_outputs(459));
    layer1_outputs(3856) <= not(layer0_outputs(4151));
    layer1_outputs(3857) <= (layer0_outputs(7257)) and (layer0_outputs(5097));
    layer1_outputs(3858) <= not((layer0_outputs(5796)) or (layer0_outputs(6611)));
    layer1_outputs(3859) <= not(layer0_outputs(7663)) or (layer0_outputs(5340));
    layer1_outputs(3860) <= '1';
    layer1_outputs(3861) <= layer0_outputs(7135);
    layer1_outputs(3862) <= (layer0_outputs(4284)) and not (layer0_outputs(1250));
    layer1_outputs(3863) <= (layer0_outputs(5149)) and not (layer0_outputs(6909));
    layer1_outputs(3864) <= layer0_outputs(6537);
    layer1_outputs(3865) <= not((layer0_outputs(4453)) xor (layer0_outputs(4094)));
    layer1_outputs(3866) <= not((layer0_outputs(2420)) or (layer0_outputs(4913)));
    layer1_outputs(3867) <= not(layer0_outputs(4438));
    layer1_outputs(3868) <= not((layer0_outputs(5995)) or (layer0_outputs(1336)));
    layer1_outputs(3869) <= not(layer0_outputs(6932));
    layer1_outputs(3870) <= (layer0_outputs(6101)) and not (layer0_outputs(6857));
    layer1_outputs(3871) <= not((layer0_outputs(5584)) or (layer0_outputs(4688)));
    layer1_outputs(3872) <= not(layer0_outputs(5294));
    layer1_outputs(3873) <= (layer0_outputs(6496)) and (layer0_outputs(6577));
    layer1_outputs(3874) <= layer0_outputs(6404);
    layer1_outputs(3875) <= layer0_outputs(4955);
    layer1_outputs(3876) <= '0';
    layer1_outputs(3877) <= '1';
    layer1_outputs(3878) <= not(layer0_outputs(5588));
    layer1_outputs(3879) <= layer0_outputs(5731);
    layer1_outputs(3880) <= not(layer0_outputs(6349));
    layer1_outputs(3881) <= not(layer0_outputs(7331));
    layer1_outputs(3882) <= (layer0_outputs(4698)) and not (layer0_outputs(1075));
    layer1_outputs(3883) <= '1';
    layer1_outputs(3884) <= not(layer0_outputs(3251));
    layer1_outputs(3885) <= not(layer0_outputs(3504));
    layer1_outputs(3886) <= '1';
    layer1_outputs(3887) <= not((layer0_outputs(1537)) xor (layer0_outputs(2639)));
    layer1_outputs(3888) <= layer0_outputs(1726);
    layer1_outputs(3889) <= (layer0_outputs(5319)) or (layer0_outputs(2612));
    layer1_outputs(3890) <= not(layer0_outputs(5773));
    layer1_outputs(3891) <= not((layer0_outputs(3373)) or (layer0_outputs(6269)));
    layer1_outputs(3892) <= '0';
    layer1_outputs(3893) <= not(layer0_outputs(7618)) or (layer0_outputs(4844));
    layer1_outputs(3894) <= (layer0_outputs(42)) and not (layer0_outputs(1979));
    layer1_outputs(3895) <= not(layer0_outputs(4860)) or (layer0_outputs(5629));
    layer1_outputs(3896) <= not(layer0_outputs(825));
    layer1_outputs(3897) <= '1';
    layer1_outputs(3898) <= '0';
    layer1_outputs(3899) <= layer0_outputs(6232);
    layer1_outputs(3900) <= layer0_outputs(7038);
    layer1_outputs(3901) <= (layer0_outputs(3391)) and not (layer0_outputs(2078));
    layer1_outputs(3902) <= '0';
    layer1_outputs(3903) <= not(layer0_outputs(1684)) or (layer0_outputs(4902));
    layer1_outputs(3904) <= layer0_outputs(6944);
    layer1_outputs(3905) <= not(layer0_outputs(7079));
    layer1_outputs(3906) <= not(layer0_outputs(1580)) or (layer0_outputs(888));
    layer1_outputs(3907) <= (layer0_outputs(5048)) or (layer0_outputs(754));
    layer1_outputs(3908) <= '0';
    layer1_outputs(3909) <= '0';
    layer1_outputs(3910) <= not(layer0_outputs(3079));
    layer1_outputs(3911) <= (layer0_outputs(1032)) and not (layer0_outputs(3750));
    layer1_outputs(3912) <= '1';
    layer1_outputs(3913) <= not(layer0_outputs(4294));
    layer1_outputs(3914) <= (layer0_outputs(1916)) xor (layer0_outputs(2730));
    layer1_outputs(3915) <= (layer0_outputs(7290)) and (layer0_outputs(4526));
    layer1_outputs(3916) <= (layer0_outputs(1388)) and not (layer0_outputs(6526));
    layer1_outputs(3917) <= not(layer0_outputs(1923)) or (layer0_outputs(3853));
    layer1_outputs(3918) <= layer0_outputs(4132);
    layer1_outputs(3919) <= layer0_outputs(4740);
    layer1_outputs(3920) <= not(layer0_outputs(1287));
    layer1_outputs(3921) <= not(layer0_outputs(6410)) or (layer0_outputs(1715));
    layer1_outputs(3922) <= (layer0_outputs(2227)) xor (layer0_outputs(1964));
    layer1_outputs(3923) <= (layer0_outputs(6861)) and not (layer0_outputs(2184));
    layer1_outputs(3924) <= not(layer0_outputs(2024)) or (layer0_outputs(4880));
    layer1_outputs(3925) <= (layer0_outputs(3673)) and not (layer0_outputs(2565));
    layer1_outputs(3926) <= (layer0_outputs(5230)) and (layer0_outputs(1164));
    layer1_outputs(3927) <= '0';
    layer1_outputs(3928) <= not((layer0_outputs(1267)) or (layer0_outputs(2025)));
    layer1_outputs(3929) <= layer0_outputs(4411);
    layer1_outputs(3930) <= not((layer0_outputs(5703)) and (layer0_outputs(911)));
    layer1_outputs(3931) <= not(layer0_outputs(7502));
    layer1_outputs(3932) <= not(layer0_outputs(7453));
    layer1_outputs(3933) <= not((layer0_outputs(4300)) or (layer0_outputs(1471)));
    layer1_outputs(3934) <= not(layer0_outputs(1772)) or (layer0_outputs(3159));
    layer1_outputs(3935) <= not(layer0_outputs(182)) or (layer0_outputs(1977));
    layer1_outputs(3936) <= not((layer0_outputs(782)) and (layer0_outputs(4157)));
    layer1_outputs(3937) <= '1';
    layer1_outputs(3938) <= '0';
    layer1_outputs(3939) <= not((layer0_outputs(668)) and (layer0_outputs(585)));
    layer1_outputs(3940) <= (layer0_outputs(6758)) or (layer0_outputs(789));
    layer1_outputs(3941) <= '1';
    layer1_outputs(3942) <= not((layer0_outputs(217)) xor (layer0_outputs(1235)));
    layer1_outputs(3943) <= not((layer0_outputs(2558)) xor (layer0_outputs(4494)));
    layer1_outputs(3944) <= '0';
    layer1_outputs(3945) <= '1';
    layer1_outputs(3946) <= not((layer0_outputs(1157)) xor (layer0_outputs(6894)));
    layer1_outputs(3947) <= not((layer0_outputs(5462)) and (layer0_outputs(6984)));
    layer1_outputs(3948) <= not(layer0_outputs(7589)) or (layer0_outputs(5429));
    layer1_outputs(3949) <= not((layer0_outputs(4919)) and (layer0_outputs(351)));
    layer1_outputs(3950) <= not(layer0_outputs(2160)) or (layer0_outputs(2348));
    layer1_outputs(3951) <= (layer0_outputs(2776)) and (layer0_outputs(5098));
    layer1_outputs(3952) <= '1';
    layer1_outputs(3953) <= not(layer0_outputs(5997)) or (layer0_outputs(7413));
    layer1_outputs(3954) <= not((layer0_outputs(7045)) or (layer0_outputs(771)));
    layer1_outputs(3955) <= (layer0_outputs(6838)) and (layer0_outputs(2166));
    layer1_outputs(3956) <= layer0_outputs(2748);
    layer1_outputs(3957) <= (layer0_outputs(240)) and not (layer0_outputs(3251));
    layer1_outputs(3958) <= (layer0_outputs(897)) and (layer0_outputs(4485));
    layer1_outputs(3959) <= not((layer0_outputs(1518)) or (layer0_outputs(3485)));
    layer1_outputs(3960) <= not((layer0_outputs(2047)) xor (layer0_outputs(5179)));
    layer1_outputs(3961) <= (layer0_outputs(627)) and not (layer0_outputs(5571));
    layer1_outputs(3962) <= not(layer0_outputs(4007));
    layer1_outputs(3963) <= (layer0_outputs(1367)) and not (layer0_outputs(879));
    layer1_outputs(3964) <= '1';
    layer1_outputs(3965) <= layer0_outputs(68);
    layer1_outputs(3966) <= '0';
    layer1_outputs(3967) <= layer0_outputs(7175);
    layer1_outputs(3968) <= not((layer0_outputs(6333)) and (layer0_outputs(3558)));
    layer1_outputs(3969) <= not((layer0_outputs(6854)) and (layer0_outputs(2422)));
    layer1_outputs(3970) <= (layer0_outputs(6540)) and not (layer0_outputs(849));
    layer1_outputs(3971) <= not((layer0_outputs(2726)) or (layer0_outputs(2857)));
    layer1_outputs(3972) <= '1';
    layer1_outputs(3973) <= (layer0_outputs(5394)) or (layer0_outputs(5186));
    layer1_outputs(3974) <= not(layer0_outputs(6180)) or (layer0_outputs(2566));
    layer1_outputs(3975) <= (layer0_outputs(84)) or (layer0_outputs(7217));
    layer1_outputs(3976) <= not(layer0_outputs(378));
    layer1_outputs(3977) <= layer0_outputs(172);
    layer1_outputs(3978) <= (layer0_outputs(6672)) and (layer0_outputs(3152));
    layer1_outputs(3979) <= not((layer0_outputs(5867)) and (layer0_outputs(5205)));
    layer1_outputs(3980) <= (layer0_outputs(2764)) and not (layer0_outputs(7485));
    layer1_outputs(3981) <= layer0_outputs(14);
    layer1_outputs(3982) <= not(layer0_outputs(5920));
    layer1_outputs(3983) <= (layer0_outputs(5299)) and not (layer0_outputs(6143));
    layer1_outputs(3984) <= not(layer0_outputs(5549)) or (layer0_outputs(547));
    layer1_outputs(3985) <= not((layer0_outputs(6630)) or (layer0_outputs(6418)));
    layer1_outputs(3986) <= not(layer0_outputs(6085));
    layer1_outputs(3987) <= '0';
    layer1_outputs(3988) <= not(layer0_outputs(570)) or (layer0_outputs(4298));
    layer1_outputs(3989) <= '1';
    layer1_outputs(3990) <= layer0_outputs(5660);
    layer1_outputs(3991) <= not(layer0_outputs(3090)) or (layer0_outputs(4596));
    layer1_outputs(3992) <= not((layer0_outputs(403)) or (layer0_outputs(279)));
    layer1_outputs(3993) <= '1';
    layer1_outputs(3994) <= '1';
    layer1_outputs(3995) <= '1';
    layer1_outputs(3996) <= (layer0_outputs(4939)) and (layer0_outputs(3214));
    layer1_outputs(3997) <= not((layer0_outputs(1668)) and (layer0_outputs(322)));
    layer1_outputs(3998) <= not(layer0_outputs(2529)) or (layer0_outputs(761));
    layer1_outputs(3999) <= '1';
    layer1_outputs(4000) <= '1';
    layer1_outputs(4001) <= '0';
    layer1_outputs(4002) <= not(layer0_outputs(3055)) or (layer0_outputs(5776));
    layer1_outputs(4003) <= '1';
    layer1_outputs(4004) <= '1';
    layer1_outputs(4005) <= not(layer0_outputs(1245));
    layer1_outputs(4006) <= not((layer0_outputs(5924)) or (layer0_outputs(7482)));
    layer1_outputs(4007) <= '0';
    layer1_outputs(4008) <= not(layer0_outputs(6191));
    layer1_outputs(4009) <= not((layer0_outputs(5542)) or (layer0_outputs(2203)));
    layer1_outputs(4010) <= not(layer0_outputs(7048));
    layer1_outputs(4011) <= not((layer0_outputs(1029)) xor (layer0_outputs(3666)));
    layer1_outputs(4012) <= not((layer0_outputs(7118)) and (layer0_outputs(6344)));
    layer1_outputs(4013) <= (layer0_outputs(5413)) and not (layer0_outputs(7610));
    layer1_outputs(4014) <= not(layer0_outputs(6919));
    layer1_outputs(4015) <= not((layer0_outputs(2035)) and (layer0_outputs(4051)));
    layer1_outputs(4016) <= '0';
    layer1_outputs(4017) <= (layer0_outputs(124)) or (layer0_outputs(2432));
    layer1_outputs(4018) <= layer0_outputs(374);
    layer1_outputs(4019) <= (layer0_outputs(4269)) and not (layer0_outputs(5314));
    layer1_outputs(4020) <= not((layer0_outputs(5283)) or (layer0_outputs(955)));
    layer1_outputs(4021) <= not(layer0_outputs(2957)) or (layer0_outputs(779));
    layer1_outputs(4022) <= not((layer0_outputs(964)) and (layer0_outputs(1364)));
    layer1_outputs(4023) <= not(layer0_outputs(5140)) or (layer0_outputs(5235));
    layer1_outputs(4024) <= not(layer0_outputs(1529));
    layer1_outputs(4025) <= not((layer0_outputs(811)) or (layer0_outputs(5897)));
    layer1_outputs(4026) <= (layer0_outputs(2991)) and (layer0_outputs(4620));
    layer1_outputs(4027) <= not(layer0_outputs(2919));
    layer1_outputs(4028) <= not((layer0_outputs(1162)) xor (layer0_outputs(7473)));
    layer1_outputs(4029) <= layer0_outputs(4014);
    layer1_outputs(4030) <= not(layer0_outputs(5261));
    layer1_outputs(4031) <= (layer0_outputs(3835)) or (layer0_outputs(7028));
    layer1_outputs(4032) <= not((layer0_outputs(1230)) or (layer0_outputs(23)));
    layer1_outputs(4033) <= not(layer0_outputs(5892));
    layer1_outputs(4034) <= not((layer0_outputs(1786)) or (layer0_outputs(3136)));
    layer1_outputs(4035) <= (layer0_outputs(2794)) and not (layer0_outputs(1062));
    layer1_outputs(4036) <= not(layer0_outputs(5386));
    layer1_outputs(4037) <= (layer0_outputs(1064)) or (layer0_outputs(4311));
    layer1_outputs(4038) <= not(layer0_outputs(5880));
    layer1_outputs(4039) <= (layer0_outputs(742)) and (layer0_outputs(6076));
    layer1_outputs(4040) <= layer0_outputs(4363);
    layer1_outputs(4041) <= (layer0_outputs(6533)) and not (layer0_outputs(13));
    layer1_outputs(4042) <= (layer0_outputs(210)) or (layer0_outputs(4438));
    layer1_outputs(4043) <= '1';
    layer1_outputs(4044) <= not((layer0_outputs(2849)) or (layer0_outputs(6355)));
    layer1_outputs(4045) <= (layer0_outputs(2059)) and not (layer0_outputs(7060));
    layer1_outputs(4046) <= not(layer0_outputs(6239)) or (layer0_outputs(7430));
    layer1_outputs(4047) <= not(layer0_outputs(3252)) or (layer0_outputs(6517));
    layer1_outputs(4048) <= (layer0_outputs(2172)) or (layer0_outputs(1374));
    layer1_outputs(4049) <= not(layer0_outputs(4988)) or (layer0_outputs(5412));
    layer1_outputs(4050) <= not((layer0_outputs(6831)) or (layer0_outputs(6199)));
    layer1_outputs(4051) <= not((layer0_outputs(3239)) or (layer0_outputs(7205)));
    layer1_outputs(4052) <= (layer0_outputs(5517)) and not (layer0_outputs(2861));
    layer1_outputs(4053) <= (layer0_outputs(5683)) or (layer0_outputs(3008));
    layer1_outputs(4054) <= (layer0_outputs(3658)) and not (layer0_outputs(3693));
    layer1_outputs(4055) <= not(layer0_outputs(5272));
    layer1_outputs(4056) <= (layer0_outputs(7007)) and not (layer0_outputs(6011));
    layer1_outputs(4057) <= (layer0_outputs(2967)) or (layer0_outputs(1609));
    layer1_outputs(4058) <= not(layer0_outputs(1513));
    layer1_outputs(4059) <= not(layer0_outputs(5515));
    layer1_outputs(4060) <= not(layer0_outputs(6439)) or (layer0_outputs(1510));
    layer1_outputs(4061) <= '1';
    layer1_outputs(4062) <= layer0_outputs(6125);
    layer1_outputs(4063) <= layer0_outputs(7146);
    layer1_outputs(4064) <= not(layer0_outputs(436)) or (layer0_outputs(6580));
    layer1_outputs(4065) <= layer0_outputs(3085);
    layer1_outputs(4066) <= not(layer0_outputs(6399));
    layer1_outputs(4067) <= '0';
    layer1_outputs(4068) <= layer0_outputs(3511);
    layer1_outputs(4069) <= not((layer0_outputs(7344)) and (layer0_outputs(3802)));
    layer1_outputs(4070) <= (layer0_outputs(6712)) and not (layer0_outputs(7205));
    layer1_outputs(4071) <= (layer0_outputs(6749)) and not (layer0_outputs(5538));
    layer1_outputs(4072) <= not(layer0_outputs(7172));
    layer1_outputs(4073) <= '0';
    layer1_outputs(4074) <= layer0_outputs(45);
    layer1_outputs(4075) <= (layer0_outputs(4915)) and not (layer0_outputs(5877));
    layer1_outputs(4076) <= (layer0_outputs(4831)) and not (layer0_outputs(37));
    layer1_outputs(4077) <= not((layer0_outputs(6619)) or (layer0_outputs(1489)));
    layer1_outputs(4078) <= (layer0_outputs(1936)) and (layer0_outputs(6186));
    layer1_outputs(4079) <= not(layer0_outputs(2048)) or (layer0_outputs(1147));
    layer1_outputs(4080) <= not((layer0_outputs(4126)) and (layer0_outputs(3663)));
    layer1_outputs(4081) <= '1';
    layer1_outputs(4082) <= not(layer0_outputs(4798));
    layer1_outputs(4083) <= (layer0_outputs(3497)) and not (layer0_outputs(294));
    layer1_outputs(4084) <= not((layer0_outputs(5233)) or (layer0_outputs(2451)));
    layer1_outputs(4085) <= layer0_outputs(1204);
    layer1_outputs(4086) <= (layer0_outputs(3112)) or (layer0_outputs(6706));
    layer1_outputs(4087) <= not(layer0_outputs(2524)) or (layer0_outputs(5251));
    layer1_outputs(4088) <= not(layer0_outputs(6620)) or (layer0_outputs(5056));
    layer1_outputs(4089) <= (layer0_outputs(7166)) and not (layer0_outputs(7440));
    layer1_outputs(4090) <= not(layer0_outputs(7298));
    layer1_outputs(4091) <= not(layer0_outputs(4312));
    layer1_outputs(4092) <= not(layer0_outputs(2691));
    layer1_outputs(4093) <= '1';
    layer1_outputs(4094) <= not((layer0_outputs(7666)) and (layer0_outputs(1607)));
    layer1_outputs(4095) <= not(layer0_outputs(7258)) or (layer0_outputs(5410));
    layer1_outputs(4096) <= '0';
    layer1_outputs(4097) <= layer0_outputs(3067);
    layer1_outputs(4098) <= (layer0_outputs(248)) and (layer0_outputs(2410));
    layer1_outputs(4099) <= not(layer0_outputs(5476));
    layer1_outputs(4100) <= (layer0_outputs(6785)) xor (layer0_outputs(2929));
    layer1_outputs(4101) <= '0';
    layer1_outputs(4102) <= '0';
    layer1_outputs(4103) <= '0';
    layer1_outputs(4104) <= not((layer0_outputs(572)) xor (layer0_outputs(2790)));
    layer1_outputs(4105) <= not((layer0_outputs(2161)) and (layer0_outputs(6009)));
    layer1_outputs(4106) <= (layer0_outputs(4856)) and not (layer0_outputs(4716));
    layer1_outputs(4107) <= (layer0_outputs(587)) and (layer0_outputs(5111));
    layer1_outputs(4108) <= not(layer0_outputs(5868));
    layer1_outputs(4109) <= not(layer0_outputs(7197));
    layer1_outputs(4110) <= (layer0_outputs(6017)) and not (layer0_outputs(3813));
    layer1_outputs(4111) <= '0';
    layer1_outputs(4112) <= (layer0_outputs(5659)) or (layer0_outputs(3800));
    layer1_outputs(4113) <= not(layer0_outputs(1568));
    layer1_outputs(4114) <= '1';
    layer1_outputs(4115) <= '0';
    layer1_outputs(4116) <= (layer0_outputs(5330)) and not (layer0_outputs(2110));
    layer1_outputs(4117) <= not(layer0_outputs(241));
    layer1_outputs(4118) <= '0';
    layer1_outputs(4119) <= not(layer0_outputs(7636));
    layer1_outputs(4120) <= (layer0_outputs(6416)) and not (layer0_outputs(413));
    layer1_outputs(4121) <= (layer0_outputs(335)) or (layer0_outputs(2822));
    layer1_outputs(4122) <= not(layer0_outputs(5154));
    layer1_outputs(4123) <= not(layer0_outputs(2744)) or (layer0_outputs(4426));
    layer1_outputs(4124) <= not(layer0_outputs(7157));
    layer1_outputs(4125) <= layer0_outputs(4477);
    layer1_outputs(4126) <= not(layer0_outputs(3114));
    layer1_outputs(4127) <= (layer0_outputs(4612)) or (layer0_outputs(5060));
    layer1_outputs(4128) <= not(layer0_outputs(5025)) or (layer0_outputs(773));
    layer1_outputs(4129) <= layer0_outputs(3081);
    layer1_outputs(4130) <= not((layer0_outputs(5552)) and (layer0_outputs(4174)));
    layer1_outputs(4131) <= (layer0_outputs(6627)) and not (layer0_outputs(3637));
    layer1_outputs(4132) <= '1';
    layer1_outputs(4133) <= (layer0_outputs(2159)) and not (layer0_outputs(1732));
    layer1_outputs(4134) <= '1';
    layer1_outputs(4135) <= not((layer0_outputs(5344)) xor (layer0_outputs(802)));
    layer1_outputs(4136) <= not((layer0_outputs(2206)) and (layer0_outputs(1763)));
    layer1_outputs(4137) <= '1';
    layer1_outputs(4138) <= not(layer0_outputs(4229)) or (layer0_outputs(5752));
    layer1_outputs(4139) <= not(layer0_outputs(439));
    layer1_outputs(4140) <= not(layer0_outputs(4590));
    layer1_outputs(4141) <= not((layer0_outputs(745)) or (layer0_outputs(249)));
    layer1_outputs(4142) <= (layer0_outputs(139)) and (layer0_outputs(2385));
    layer1_outputs(4143) <= (layer0_outputs(4779)) and not (layer0_outputs(6550));
    layer1_outputs(4144) <= '1';
    layer1_outputs(4145) <= '0';
    layer1_outputs(4146) <= not(layer0_outputs(6308)) or (layer0_outputs(2306));
    layer1_outputs(4147) <= (layer0_outputs(3118)) and not (layer0_outputs(765));
    layer1_outputs(4148) <= (layer0_outputs(6021)) and (layer0_outputs(2686));
    layer1_outputs(4149) <= '1';
    layer1_outputs(4150) <= not(layer0_outputs(2821));
    layer1_outputs(4151) <= layer0_outputs(410);
    layer1_outputs(4152) <= (layer0_outputs(2470)) and not (layer0_outputs(3712));
    layer1_outputs(4153) <= not((layer0_outputs(3931)) and (layer0_outputs(7647)));
    layer1_outputs(4154) <= not(layer0_outputs(5817));
    layer1_outputs(4155) <= (layer0_outputs(2452)) and not (layer0_outputs(5738));
    layer1_outputs(4156) <= not(layer0_outputs(3547)) or (layer0_outputs(2796));
    layer1_outputs(4157) <= (layer0_outputs(4152)) and not (layer0_outputs(1428));
    layer1_outputs(4158) <= '1';
    layer1_outputs(4159) <= '1';
    layer1_outputs(4160) <= '1';
    layer1_outputs(4161) <= '0';
    layer1_outputs(4162) <= (layer0_outputs(3610)) or (layer0_outputs(3616));
    layer1_outputs(4163) <= not(layer0_outputs(665));
    layer1_outputs(4164) <= not(layer0_outputs(2016)) or (layer0_outputs(5347));
    layer1_outputs(4165) <= not(layer0_outputs(3996)) or (layer0_outputs(1849));
    layer1_outputs(4166) <= not(layer0_outputs(2630));
    layer1_outputs(4167) <= not(layer0_outputs(5561));
    layer1_outputs(4168) <= not((layer0_outputs(3464)) and (layer0_outputs(5154)));
    layer1_outputs(4169) <= layer0_outputs(5401);
    layer1_outputs(4170) <= not(layer0_outputs(5514));
    layer1_outputs(4171) <= layer0_outputs(2437);
    layer1_outputs(4172) <= (layer0_outputs(3533)) and not (layer0_outputs(715));
    layer1_outputs(4173) <= '1';
    layer1_outputs(4174) <= (layer0_outputs(5936)) and not (layer0_outputs(1208));
    layer1_outputs(4175) <= layer0_outputs(5266);
    layer1_outputs(4176) <= layer0_outputs(3836);
    layer1_outputs(4177) <= not(layer0_outputs(3744));
    layer1_outputs(4178) <= (layer0_outputs(3826)) and not (layer0_outputs(3406));
    layer1_outputs(4179) <= '1';
    layer1_outputs(4180) <= '0';
    layer1_outputs(4181) <= not(layer0_outputs(5201));
    layer1_outputs(4182) <= '1';
    layer1_outputs(4183) <= not(layer0_outputs(2951));
    layer1_outputs(4184) <= not(layer0_outputs(1271));
    layer1_outputs(4185) <= not(layer0_outputs(4310));
    layer1_outputs(4186) <= layer0_outputs(677);
    layer1_outputs(4187) <= (layer0_outputs(6766)) and not (layer0_outputs(4136));
    layer1_outputs(4188) <= '1';
    layer1_outputs(4189) <= layer0_outputs(966);
    layer1_outputs(4190) <= (layer0_outputs(6693)) or (layer0_outputs(5572));
    layer1_outputs(4191) <= not(layer0_outputs(138));
    layer1_outputs(4192) <= '1';
    layer1_outputs(4193) <= not(layer0_outputs(3453)) or (layer0_outputs(3885));
    layer1_outputs(4194) <= not(layer0_outputs(4135)) or (layer0_outputs(4058));
    layer1_outputs(4195) <= '1';
    layer1_outputs(4196) <= not(layer0_outputs(4914)) or (layer0_outputs(5979));
    layer1_outputs(4197) <= not((layer0_outputs(5815)) or (layer0_outputs(3200)));
    layer1_outputs(4198) <= '0';
    layer1_outputs(4199) <= '0';
    layer1_outputs(4200) <= (layer0_outputs(4206)) and not (layer0_outputs(2658));
    layer1_outputs(4201) <= not((layer0_outputs(5266)) or (layer0_outputs(1875)));
    layer1_outputs(4202) <= layer0_outputs(2550);
    layer1_outputs(4203) <= (layer0_outputs(6598)) or (layer0_outputs(4481));
    layer1_outputs(4204) <= not(layer0_outputs(1804));
    layer1_outputs(4205) <= not(layer0_outputs(823)) or (layer0_outputs(552));
    layer1_outputs(4206) <= layer0_outputs(6871);
    layer1_outputs(4207) <= '1';
    layer1_outputs(4208) <= '0';
    layer1_outputs(4209) <= '1';
    layer1_outputs(4210) <= (layer0_outputs(2500)) and not (layer0_outputs(3355));
    layer1_outputs(4211) <= '0';
    layer1_outputs(4212) <= not((layer0_outputs(4572)) and (layer0_outputs(6350)));
    layer1_outputs(4213) <= not(layer0_outputs(2664));
    layer1_outputs(4214) <= (layer0_outputs(2988)) and not (layer0_outputs(5445));
    layer1_outputs(4215) <= layer0_outputs(3859);
    layer1_outputs(4216) <= '0';
    layer1_outputs(4217) <= (layer0_outputs(4178)) and (layer0_outputs(7649));
    layer1_outputs(4218) <= not(layer0_outputs(5343)) or (layer0_outputs(2093));
    layer1_outputs(4219) <= not((layer0_outputs(1115)) and (layer0_outputs(6637)));
    layer1_outputs(4220) <= '1';
    layer1_outputs(4221) <= not(layer0_outputs(7459));
    layer1_outputs(4222) <= '0';
    layer1_outputs(4223) <= (layer0_outputs(4241)) and not (layer0_outputs(2765));
    layer1_outputs(4224) <= layer0_outputs(3846);
    layer1_outputs(4225) <= (layer0_outputs(6612)) and not (layer0_outputs(5075));
    layer1_outputs(4226) <= not((layer0_outputs(7433)) or (layer0_outputs(2186)));
    layer1_outputs(4227) <= (layer0_outputs(6894)) and not (layer0_outputs(4052));
    layer1_outputs(4228) <= layer0_outputs(1514);
    layer1_outputs(4229) <= not(layer0_outputs(5333));
    layer1_outputs(4230) <= (layer0_outputs(7542)) and (layer0_outputs(4504));
    layer1_outputs(4231) <= not(layer0_outputs(5213)) or (layer0_outputs(2535));
    layer1_outputs(4232) <= (layer0_outputs(2645)) and (layer0_outputs(213));
    layer1_outputs(4233) <= (layer0_outputs(702)) and (layer0_outputs(4432));
    layer1_outputs(4234) <= layer0_outputs(243);
    layer1_outputs(4235) <= (layer0_outputs(7392)) and (layer0_outputs(2562));
    layer1_outputs(4236) <= '0';
    layer1_outputs(4237) <= not(layer0_outputs(7508));
    layer1_outputs(4238) <= layer0_outputs(2073);
    layer1_outputs(4239) <= layer0_outputs(883);
    layer1_outputs(4240) <= (layer0_outputs(1932)) and not (layer0_outputs(5725));
    layer1_outputs(4241) <= '1';
    layer1_outputs(4242) <= layer0_outputs(6311);
    layer1_outputs(4243) <= (layer0_outputs(1888)) and not (layer0_outputs(1161));
    layer1_outputs(4244) <= '1';
    layer1_outputs(4245) <= layer0_outputs(7239);
    layer1_outputs(4246) <= (layer0_outputs(7639)) or (layer0_outputs(5547));
    layer1_outputs(4247) <= '1';
    layer1_outputs(4248) <= not(layer0_outputs(196));
    layer1_outputs(4249) <= not(layer0_outputs(704)) or (layer0_outputs(4777));
    layer1_outputs(4250) <= '1';
    layer1_outputs(4251) <= not((layer0_outputs(457)) and (layer0_outputs(751)));
    layer1_outputs(4252) <= '0';
    layer1_outputs(4253) <= (layer0_outputs(1455)) xor (layer0_outputs(6085));
    layer1_outputs(4254) <= not(layer0_outputs(3893));
    layer1_outputs(4255) <= not((layer0_outputs(3030)) or (layer0_outputs(2920)));
    layer1_outputs(4256) <= not((layer0_outputs(3306)) or (layer0_outputs(2885)));
    layer1_outputs(4257) <= layer0_outputs(1324);
    layer1_outputs(4258) <= layer0_outputs(5440);
    layer1_outputs(4259) <= not((layer0_outputs(1933)) or (layer0_outputs(6585)));
    layer1_outputs(4260) <= (layer0_outputs(4720)) and (layer0_outputs(2510));
    layer1_outputs(4261) <= (layer0_outputs(488)) and (layer0_outputs(4792));
    layer1_outputs(4262) <= '1';
    layer1_outputs(4263) <= (layer0_outputs(2544)) and not (layer0_outputs(1390));
    layer1_outputs(4264) <= (layer0_outputs(6951)) and not (layer0_outputs(5555));
    layer1_outputs(4265) <= (layer0_outputs(6253)) and not (layer0_outputs(7409));
    layer1_outputs(4266) <= (layer0_outputs(7392)) or (layer0_outputs(4400));
    layer1_outputs(4267) <= layer0_outputs(5184);
    layer1_outputs(4268) <= not(layer0_outputs(4465));
    layer1_outputs(4269) <= (layer0_outputs(3127)) and not (layer0_outputs(2710));
    layer1_outputs(4270) <= not(layer0_outputs(1829));
    layer1_outputs(4271) <= not(layer0_outputs(3328)) or (layer0_outputs(7423));
    layer1_outputs(4272) <= not(layer0_outputs(6583)) or (layer0_outputs(360));
    layer1_outputs(4273) <= not(layer0_outputs(1666));
    layer1_outputs(4274) <= (layer0_outputs(6298)) xor (layer0_outputs(2355));
    layer1_outputs(4275) <= not(layer0_outputs(3764)) or (layer0_outputs(7537));
    layer1_outputs(4276) <= (layer0_outputs(4215)) and (layer0_outputs(7092));
    layer1_outputs(4277) <= (layer0_outputs(2104)) and (layer0_outputs(1956));
    layer1_outputs(4278) <= layer0_outputs(6882);
    layer1_outputs(4279) <= (layer0_outputs(1442)) and not (layer0_outputs(2662));
    layer1_outputs(4280) <= layer0_outputs(6377);
    layer1_outputs(4281) <= not((layer0_outputs(1650)) and (layer0_outputs(6430)));
    layer1_outputs(4282) <= '1';
    layer1_outputs(4283) <= layer0_outputs(3394);
    layer1_outputs(4284) <= layer0_outputs(5787);
    layer1_outputs(4285) <= layer0_outputs(4084);
    layer1_outputs(4286) <= not(layer0_outputs(3090));
    layer1_outputs(4287) <= (layer0_outputs(3469)) and (layer0_outputs(2496));
    layer1_outputs(4288) <= (layer0_outputs(4469)) and not (layer0_outputs(4566));
    layer1_outputs(4289) <= not(layer0_outputs(2751));
    layer1_outputs(4290) <= layer0_outputs(2236);
    layer1_outputs(4291) <= not(layer0_outputs(4721)) or (layer0_outputs(4025));
    layer1_outputs(4292) <= not(layer0_outputs(4537));
    layer1_outputs(4293) <= (layer0_outputs(1596)) and not (layer0_outputs(716));
    layer1_outputs(4294) <= not(layer0_outputs(3557)) or (layer0_outputs(3094));
    layer1_outputs(4295) <= not((layer0_outputs(3997)) and (layer0_outputs(4185)));
    layer1_outputs(4296) <= not(layer0_outputs(4482)) or (layer0_outputs(1766));
    layer1_outputs(4297) <= layer0_outputs(7576);
    layer1_outputs(4298) <= not((layer0_outputs(3619)) or (layer0_outputs(639)));
    layer1_outputs(4299) <= not(layer0_outputs(1521));
    layer1_outputs(4300) <= not((layer0_outputs(1469)) or (layer0_outputs(6079)));
    layer1_outputs(4301) <= not(layer0_outputs(940));
    layer1_outputs(4302) <= not(layer0_outputs(2711));
    layer1_outputs(4303) <= not((layer0_outputs(3138)) and (layer0_outputs(831)));
    layer1_outputs(4304) <= (layer0_outputs(5415)) and (layer0_outputs(170));
    layer1_outputs(4305) <= layer0_outputs(4041);
    layer1_outputs(4306) <= not((layer0_outputs(5944)) and (layer0_outputs(3647)));
    layer1_outputs(4307) <= not((layer0_outputs(6504)) and (layer0_outputs(317)));
    layer1_outputs(4308) <= not((layer0_outputs(4551)) or (layer0_outputs(6133)));
    layer1_outputs(4309) <= '0';
    layer1_outputs(4310) <= not((layer0_outputs(2873)) or (layer0_outputs(5833)));
    layer1_outputs(4311) <= (layer0_outputs(7109)) and not (layer0_outputs(591));
    layer1_outputs(4312) <= not((layer0_outputs(4105)) and (layer0_outputs(1475)));
    layer1_outputs(4313) <= '0';
    layer1_outputs(4314) <= '0';
    layer1_outputs(4315) <= '0';
    layer1_outputs(4316) <= '1';
    layer1_outputs(4317) <= '0';
    layer1_outputs(4318) <= (layer0_outputs(5261)) and not (layer0_outputs(5920));
    layer1_outputs(4319) <= '0';
    layer1_outputs(4320) <= not(layer0_outputs(6734));
    layer1_outputs(4321) <= not((layer0_outputs(7326)) or (layer0_outputs(5789)));
    layer1_outputs(4322) <= (layer0_outputs(7171)) and (layer0_outputs(4307));
    layer1_outputs(4323) <= (layer0_outputs(3927)) and not (layer0_outputs(442));
    layer1_outputs(4324) <= not(layer0_outputs(4276)) or (layer0_outputs(5527));
    layer1_outputs(4325) <= '0';
    layer1_outputs(4326) <= '1';
    layer1_outputs(4327) <= (layer0_outputs(1467)) and not (layer0_outputs(2781));
    layer1_outputs(4328) <= (layer0_outputs(3472)) or (layer0_outputs(7643));
    layer1_outputs(4329) <= (layer0_outputs(2224)) and not (layer0_outputs(7305));
    layer1_outputs(4330) <= not(layer0_outputs(4584));
    layer1_outputs(4331) <= (layer0_outputs(3771)) and not (layer0_outputs(4812));
    layer1_outputs(4332) <= (layer0_outputs(118)) and not (layer0_outputs(5434));
    layer1_outputs(4333) <= not(layer0_outputs(6136));
    layer1_outputs(4334) <= (layer0_outputs(2526)) and (layer0_outputs(1238));
    layer1_outputs(4335) <= (layer0_outputs(3882)) and (layer0_outputs(5290));
    layer1_outputs(4336) <= '0';
    layer1_outputs(4337) <= (layer0_outputs(3587)) and (layer0_outputs(510));
    layer1_outputs(4338) <= (layer0_outputs(7103)) and (layer0_outputs(5738));
    layer1_outputs(4339) <= (layer0_outputs(2351)) and not (layer0_outputs(294));
    layer1_outputs(4340) <= (layer0_outputs(1239)) and not (layer0_outputs(7668));
    layer1_outputs(4341) <= (layer0_outputs(2547)) and not (layer0_outputs(1197));
    layer1_outputs(4342) <= '1';
    layer1_outputs(4343) <= (layer0_outputs(1496)) and (layer0_outputs(4065));
    layer1_outputs(4344) <= '0';
    layer1_outputs(4345) <= (layer0_outputs(6814)) and (layer0_outputs(1803));
    layer1_outputs(4346) <= '0';
    layer1_outputs(4347) <= layer0_outputs(943);
    layer1_outputs(4348) <= (layer0_outputs(110)) xor (layer0_outputs(5073));
    layer1_outputs(4349) <= '0';
    layer1_outputs(4350) <= (layer0_outputs(3065)) xor (layer0_outputs(6386));
    layer1_outputs(4351) <= not(layer0_outputs(2988));
    layer1_outputs(4352) <= layer0_outputs(3626);
    layer1_outputs(4353) <= layer0_outputs(1422);
    layer1_outputs(4354) <= '0';
    layer1_outputs(4355) <= not((layer0_outputs(7357)) or (layer0_outputs(6820)));
    layer1_outputs(4356) <= (layer0_outputs(2107)) xor (layer0_outputs(6945));
    layer1_outputs(4357) <= layer0_outputs(6392);
    layer1_outputs(4358) <= not(layer0_outputs(875));
    layer1_outputs(4359) <= '1';
    layer1_outputs(4360) <= '0';
    layer1_outputs(4361) <= (layer0_outputs(7188)) or (layer0_outputs(2872));
    layer1_outputs(4362) <= (layer0_outputs(2155)) and not (layer0_outputs(1139));
    layer1_outputs(4363) <= not(layer0_outputs(681));
    layer1_outputs(4364) <= not(layer0_outputs(4315));
    layer1_outputs(4365) <= not((layer0_outputs(5597)) and (layer0_outputs(5188)));
    layer1_outputs(4366) <= '0';
    layer1_outputs(4367) <= not(layer0_outputs(5471));
    layer1_outputs(4368) <= not((layer0_outputs(2745)) and (layer0_outputs(4717)));
    layer1_outputs(4369) <= not(layer0_outputs(2093));
    layer1_outputs(4370) <= not(layer0_outputs(7225));
    layer1_outputs(4371) <= '0';
    layer1_outputs(4372) <= (layer0_outputs(2180)) and (layer0_outputs(6248));
    layer1_outputs(4373) <= '1';
    layer1_outputs(4374) <= not(layer0_outputs(1068)) or (layer0_outputs(1967));
    layer1_outputs(4375) <= not(layer0_outputs(6299));
    layer1_outputs(4376) <= not(layer0_outputs(4985)) or (layer0_outputs(6921));
    layer1_outputs(4377) <= not(layer0_outputs(6752));
    layer1_outputs(4378) <= layer0_outputs(6724);
    layer1_outputs(4379) <= '0';
    layer1_outputs(4380) <= '0';
    layer1_outputs(4381) <= layer0_outputs(6909);
    layer1_outputs(4382) <= not(layer0_outputs(3357));
    layer1_outputs(4383) <= '0';
    layer1_outputs(4384) <= not(layer0_outputs(7095));
    layer1_outputs(4385) <= not(layer0_outputs(2332)) or (layer0_outputs(3414));
    layer1_outputs(4386) <= not(layer0_outputs(2845)) or (layer0_outputs(7229));
    layer1_outputs(4387) <= not(layer0_outputs(4973));
    layer1_outputs(4388) <= not(layer0_outputs(4768));
    layer1_outputs(4389) <= layer0_outputs(5128);
    layer1_outputs(4390) <= layer0_outputs(1769);
    layer1_outputs(4391) <= (layer0_outputs(1521)) and not (layer0_outputs(2486));
    layer1_outputs(4392) <= (layer0_outputs(1174)) and (layer0_outputs(2174));
    layer1_outputs(4393) <= not(layer0_outputs(1240)) or (layer0_outputs(1491));
    layer1_outputs(4394) <= not(layer0_outputs(6300)) or (layer0_outputs(5337));
    layer1_outputs(4395) <= (layer0_outputs(7623)) and not (layer0_outputs(3998));
    layer1_outputs(4396) <= layer0_outputs(3947);
    layer1_outputs(4397) <= not((layer0_outputs(1668)) or (layer0_outputs(5709)));
    layer1_outputs(4398) <= layer0_outputs(3889);
    layer1_outputs(4399) <= '1';
    layer1_outputs(4400) <= not(layer0_outputs(6450));
    layer1_outputs(4401) <= not(layer0_outputs(5481));
    layer1_outputs(4402) <= (layer0_outputs(2704)) and (layer0_outputs(4011));
    layer1_outputs(4403) <= not(layer0_outputs(2956)) or (layer0_outputs(1097));
    layer1_outputs(4404) <= (layer0_outputs(7578)) and (layer0_outputs(1722));
    layer1_outputs(4405) <= (layer0_outputs(4464)) and not (layer0_outputs(2423));
    layer1_outputs(4406) <= not((layer0_outputs(6840)) and (layer0_outputs(5274)));
    layer1_outputs(4407) <= not(layer0_outputs(165)) or (layer0_outputs(2176));
    layer1_outputs(4408) <= not(layer0_outputs(1655));
    layer1_outputs(4409) <= layer0_outputs(800);
    layer1_outputs(4410) <= not(layer0_outputs(6763));
    layer1_outputs(4411) <= (layer0_outputs(6276)) and not (layer0_outputs(5255));
    layer1_outputs(4412) <= (layer0_outputs(6406)) and (layer0_outputs(4678));
    layer1_outputs(4413) <= not(layer0_outputs(64)) or (layer0_outputs(15));
    layer1_outputs(4414) <= not(layer0_outputs(3126)) or (layer0_outputs(3718));
    layer1_outputs(4415) <= not(layer0_outputs(2708)) or (layer0_outputs(6538));
    layer1_outputs(4416) <= layer0_outputs(5763);
    layer1_outputs(4417) <= '0';
    layer1_outputs(4418) <= (layer0_outputs(3279)) and not (layer0_outputs(5633));
    layer1_outputs(4419) <= layer0_outputs(529);
    layer1_outputs(4420) <= not((layer0_outputs(7076)) and (layer0_outputs(4403)));
    layer1_outputs(4421) <= '0';
    layer1_outputs(4422) <= not(layer0_outputs(734));
    layer1_outputs(4423) <= not(layer0_outputs(3742)) or (layer0_outputs(3704));
    layer1_outputs(4424) <= (layer0_outputs(120)) and not (layer0_outputs(200));
    layer1_outputs(4425) <= not(layer0_outputs(1248));
    layer1_outputs(4426) <= not((layer0_outputs(684)) or (layer0_outputs(2313)));
    layer1_outputs(4427) <= (layer0_outputs(5516)) and (layer0_outputs(2819));
    layer1_outputs(4428) <= not(layer0_outputs(6194)) or (layer0_outputs(1504));
    layer1_outputs(4429) <= '1';
    layer1_outputs(4430) <= not(layer0_outputs(7594));
    layer1_outputs(4431) <= '0';
    layer1_outputs(4432) <= '0';
    layer1_outputs(4433) <= not((layer0_outputs(2488)) or (layer0_outputs(1577)));
    layer1_outputs(4434) <= '1';
    layer1_outputs(4435) <= (layer0_outputs(3178)) or (layer0_outputs(1539));
    layer1_outputs(4436) <= (layer0_outputs(1340)) and not (layer0_outputs(1564));
    layer1_outputs(4437) <= layer0_outputs(5232);
    layer1_outputs(4438) <= '0';
    layer1_outputs(4439) <= not((layer0_outputs(6374)) and (layer0_outputs(5031)));
    layer1_outputs(4440) <= not(layer0_outputs(5546));
    layer1_outputs(4441) <= not(layer0_outputs(3351)) or (layer0_outputs(7417));
    layer1_outputs(4442) <= '1';
    layer1_outputs(4443) <= layer0_outputs(2473);
    layer1_outputs(4444) <= '1';
    layer1_outputs(4445) <= not((layer0_outputs(4528)) or (layer0_outputs(5906)));
    layer1_outputs(4446) <= (layer0_outputs(4639)) and not (layer0_outputs(5448));
    layer1_outputs(4447) <= not((layer0_outputs(6954)) and (layer0_outputs(3171)));
    layer1_outputs(4448) <= '1';
    layer1_outputs(4449) <= layer0_outputs(6865);
    layer1_outputs(4450) <= layer0_outputs(1100);
    layer1_outputs(4451) <= '0';
    layer1_outputs(4452) <= '1';
    layer1_outputs(4453) <= (layer0_outputs(5494)) and not (layer0_outputs(974));
    layer1_outputs(4454) <= layer0_outputs(2778);
    layer1_outputs(4455) <= (layer0_outputs(5590)) and (layer0_outputs(3504));
    layer1_outputs(4456) <= not(layer0_outputs(5901)) or (layer0_outputs(1054));
    layer1_outputs(4457) <= (layer0_outputs(7121)) or (layer0_outputs(5254));
    layer1_outputs(4458) <= '0';
    layer1_outputs(4459) <= not(layer0_outputs(876));
    layer1_outputs(4460) <= '1';
    layer1_outputs(4461) <= not(layer0_outputs(531)) or (layer0_outputs(1338));
    layer1_outputs(4462) <= not((layer0_outputs(6428)) and (layer0_outputs(2250)));
    layer1_outputs(4463) <= (layer0_outputs(6501)) and not (layer0_outputs(2514));
    layer1_outputs(4464) <= not(layer0_outputs(2109));
    layer1_outputs(4465) <= (layer0_outputs(125)) or (layer0_outputs(4758));
    layer1_outputs(4466) <= (layer0_outputs(3464)) and (layer0_outputs(6327));
    layer1_outputs(4467) <= not((layer0_outputs(4841)) or (layer0_outputs(3709)));
    layer1_outputs(4468) <= not(layer0_outputs(7145)) or (layer0_outputs(4715));
    layer1_outputs(4469) <= not((layer0_outputs(3287)) or (layer0_outputs(903)));
    layer1_outputs(4470) <= (layer0_outputs(6461)) and not (layer0_outputs(3541));
    layer1_outputs(4471) <= not((layer0_outputs(6470)) or (layer0_outputs(4948)));
    layer1_outputs(4472) <= not(layer0_outputs(363)) or (layer0_outputs(3083));
    layer1_outputs(4473) <= layer0_outputs(310);
    layer1_outputs(4474) <= (layer0_outputs(6538)) and (layer0_outputs(784));
    layer1_outputs(4475) <= not((layer0_outputs(563)) and (layer0_outputs(7032)));
    layer1_outputs(4476) <= not(layer0_outputs(5069)) or (layer0_outputs(1808));
    layer1_outputs(4477) <= not((layer0_outputs(4581)) or (layer0_outputs(3432)));
    layer1_outputs(4478) <= (layer0_outputs(2692)) or (layer0_outputs(1123));
    layer1_outputs(4479) <= '1';
    layer1_outputs(4480) <= (layer0_outputs(4983)) and not (layer0_outputs(3806));
    layer1_outputs(4481) <= not(layer0_outputs(1479)) or (layer0_outputs(5225));
    layer1_outputs(4482) <= (layer0_outputs(236)) and (layer0_outputs(2678));
    layer1_outputs(4483) <= layer0_outputs(1000);
    layer1_outputs(4484) <= '0';
    layer1_outputs(4485) <= '1';
    layer1_outputs(4486) <= not(layer0_outputs(6803));
    layer1_outputs(4487) <= (layer0_outputs(5390)) or (layer0_outputs(4567));
    layer1_outputs(4488) <= (layer0_outputs(3839)) or (layer0_outputs(1190));
    layer1_outputs(4489) <= '1';
    layer1_outputs(4490) <= not((layer0_outputs(6957)) and (layer0_outputs(1473)));
    layer1_outputs(4491) <= not((layer0_outputs(6115)) or (layer0_outputs(2790)));
    layer1_outputs(4492) <= '0';
    layer1_outputs(4493) <= not(layer0_outputs(6230));
    layer1_outputs(4494) <= (layer0_outputs(1283)) and not (layer0_outputs(7136));
    layer1_outputs(4495) <= (layer0_outputs(6696)) and (layer0_outputs(2055));
    layer1_outputs(4496) <= (layer0_outputs(6132)) and not (layer0_outputs(5088));
    layer1_outputs(4497) <= (layer0_outputs(3367)) and not (layer0_outputs(1765));
    layer1_outputs(4498) <= '0';
    layer1_outputs(4499) <= '0';
    layer1_outputs(4500) <= not((layer0_outputs(4816)) xor (layer0_outputs(1444)));
    layer1_outputs(4501) <= '1';
    layer1_outputs(4502) <= not((layer0_outputs(4540)) and (layer0_outputs(5325)));
    layer1_outputs(4503) <= '0';
    layer1_outputs(4504) <= not((layer0_outputs(2680)) xor (layer0_outputs(1966)));
    layer1_outputs(4505) <= (layer0_outputs(5250)) and (layer0_outputs(6736));
    layer1_outputs(4506) <= not(layer0_outputs(1657)) or (layer0_outputs(3833));
    layer1_outputs(4507) <= layer0_outputs(4382);
    layer1_outputs(4508) <= (layer0_outputs(795)) or (layer0_outputs(2910));
    layer1_outputs(4509) <= (layer0_outputs(373)) and not (layer0_outputs(592));
    layer1_outputs(4510) <= (layer0_outputs(7012)) and not (layer0_outputs(4938));
    layer1_outputs(4511) <= not((layer0_outputs(3897)) and (layer0_outputs(5123)));
    layer1_outputs(4512) <= not(layer0_outputs(7493)) or (layer0_outputs(6470));
    layer1_outputs(4513) <= layer0_outputs(3815);
    layer1_outputs(4514) <= not((layer0_outputs(6285)) and (layer0_outputs(3725)));
    layer1_outputs(4515) <= not(layer0_outputs(6464));
    layer1_outputs(4516) <= not(layer0_outputs(6223));
    layer1_outputs(4517) <= (layer0_outputs(7425)) and not (layer0_outputs(656));
    layer1_outputs(4518) <= not(layer0_outputs(2407));
    layer1_outputs(4519) <= not(layer0_outputs(3058)) or (layer0_outputs(2197));
    layer1_outputs(4520) <= (layer0_outputs(1955)) and not (layer0_outputs(4130));
    layer1_outputs(4521) <= '1';
    layer1_outputs(4522) <= '1';
    layer1_outputs(4523) <= not((layer0_outputs(4255)) or (layer0_outputs(3215)));
    layer1_outputs(4524) <= not(layer0_outputs(1199)) or (layer0_outputs(5493));
    layer1_outputs(4525) <= not(layer0_outputs(4395)) or (layer0_outputs(1189));
    layer1_outputs(4526) <= layer0_outputs(6427);
    layer1_outputs(4527) <= not((layer0_outputs(1096)) and (layer0_outputs(7556)));
    layer1_outputs(4528) <= not(layer0_outputs(7105)) or (layer0_outputs(204));
    layer1_outputs(4529) <= '1';
    layer1_outputs(4530) <= '1';
    layer1_outputs(4531) <= (layer0_outputs(2789)) and not (layer0_outputs(3301));
    layer1_outputs(4532) <= not((layer0_outputs(7666)) and (layer0_outputs(6460)));
    layer1_outputs(4533) <= layer0_outputs(5176);
    layer1_outputs(4534) <= (layer0_outputs(2888)) xor (layer0_outputs(6072));
    layer1_outputs(4535) <= not((layer0_outputs(4498)) or (layer0_outputs(7160)));
    layer1_outputs(4536) <= not((layer0_outputs(2662)) or (layer0_outputs(552)));
    layer1_outputs(4537) <= not(layer0_outputs(4240)) or (layer0_outputs(3607));
    layer1_outputs(4538) <= (layer0_outputs(6319)) and not (layer0_outputs(7056));
    layer1_outputs(4539) <= layer0_outputs(1024);
    layer1_outputs(4540) <= layer0_outputs(6694);
    layer1_outputs(4541) <= '1';
    layer1_outputs(4542) <= '1';
    layer1_outputs(4543) <= layer0_outputs(3434);
    layer1_outputs(4544) <= (layer0_outputs(139)) and not (layer0_outputs(7628));
    layer1_outputs(4545) <= not(layer0_outputs(1057));
    layer1_outputs(4546) <= layer0_outputs(696);
    layer1_outputs(4547) <= not((layer0_outputs(5826)) or (layer0_outputs(1304)));
    layer1_outputs(4548) <= not((layer0_outputs(7462)) or (layer0_outputs(5689)));
    layer1_outputs(4549) <= not((layer0_outputs(352)) and (layer0_outputs(1117)));
    layer1_outputs(4550) <= not(layer0_outputs(4737)) or (layer0_outputs(6970));
    layer1_outputs(4551) <= '0';
    layer1_outputs(4552) <= '0';
    layer1_outputs(4553) <= (layer0_outputs(2773)) and not (layer0_outputs(6405));
    layer1_outputs(4554) <= layer0_outputs(2807);
    layer1_outputs(4555) <= (layer0_outputs(2796)) and not (layer0_outputs(2922));
    layer1_outputs(4556) <= layer0_outputs(2751);
    layer1_outputs(4557) <= not((layer0_outputs(2523)) xor (layer0_outputs(3388)));
    layer1_outputs(4558) <= not(layer0_outputs(6798)) or (layer0_outputs(5982));
    layer1_outputs(4559) <= layer0_outputs(2839);
    layer1_outputs(4560) <= (layer0_outputs(2686)) and (layer0_outputs(6570));
    layer1_outputs(4561) <= '0';
    layer1_outputs(4562) <= (layer0_outputs(2934)) and not (layer0_outputs(3232));
    layer1_outputs(4563) <= layer0_outputs(2703);
    layer1_outputs(4564) <= '0';
    layer1_outputs(4565) <= '0';
    layer1_outputs(4566) <= not(layer0_outputs(3103));
    layer1_outputs(4567) <= not(layer0_outputs(5982)) or (layer0_outputs(2479));
    layer1_outputs(4568) <= '0';
    layer1_outputs(4569) <= not(layer0_outputs(6755));
    layer1_outputs(4570) <= '1';
    layer1_outputs(4571) <= '0';
    layer1_outputs(4572) <= '0';
    layer1_outputs(4573) <= layer0_outputs(2139);
    layer1_outputs(4574) <= '1';
    layer1_outputs(4575) <= layer0_outputs(231);
    layer1_outputs(4576) <= not((layer0_outputs(4157)) and (layer0_outputs(2505)));
    layer1_outputs(4577) <= layer0_outputs(4812);
    layer1_outputs(4578) <= layer0_outputs(6571);
    layer1_outputs(4579) <= not(layer0_outputs(6403));
    layer1_outputs(4580) <= not(layer0_outputs(4650)) or (layer0_outputs(930));
    layer1_outputs(4581) <= (layer0_outputs(1090)) and (layer0_outputs(5739));
    layer1_outputs(4582) <= not((layer0_outputs(6898)) or (layer0_outputs(3889)));
    layer1_outputs(4583) <= not(layer0_outputs(7641)) or (layer0_outputs(1341));
    layer1_outputs(4584) <= layer0_outputs(5135);
    layer1_outputs(4585) <= not((layer0_outputs(5937)) and (layer0_outputs(1522)));
    layer1_outputs(4586) <= (layer0_outputs(4376)) or (layer0_outputs(5651));
    layer1_outputs(4587) <= (layer0_outputs(307)) or (layer0_outputs(2225));
    layer1_outputs(4588) <= layer0_outputs(4951);
    layer1_outputs(4589) <= (layer0_outputs(6819)) and (layer0_outputs(6875));
    layer1_outputs(4590) <= (layer0_outputs(7675)) and (layer0_outputs(792));
    layer1_outputs(4591) <= not(layer0_outputs(1911));
    layer1_outputs(4592) <= not(layer0_outputs(6979));
    layer1_outputs(4593) <= layer0_outputs(6098);
    layer1_outputs(4594) <= layer0_outputs(144);
    layer1_outputs(4595) <= (layer0_outputs(6981)) and (layer0_outputs(6907));
    layer1_outputs(4596) <= layer0_outputs(5022);
    layer1_outputs(4597) <= '0';
    layer1_outputs(4598) <= not(layer0_outputs(4314)) or (layer0_outputs(1874));
    layer1_outputs(4599) <= layer0_outputs(886);
    layer1_outputs(4600) <= layer0_outputs(855);
    layer1_outputs(4601) <= not(layer0_outputs(3990)) or (layer0_outputs(3335));
    layer1_outputs(4602) <= not(layer0_outputs(5352));
    layer1_outputs(4603) <= layer0_outputs(5247);
    layer1_outputs(4604) <= '0';
    layer1_outputs(4605) <= (layer0_outputs(5594)) or (layer0_outputs(2465));
    layer1_outputs(4606) <= not(layer0_outputs(6219)) or (layer0_outputs(6329));
    layer1_outputs(4607) <= (layer0_outputs(713)) and not (layer0_outputs(143));
    layer1_outputs(4608) <= not(layer0_outputs(3417));
    layer1_outputs(4609) <= layer0_outputs(4115);
    layer1_outputs(4610) <= (layer0_outputs(3617)) or (layer0_outputs(899));
    layer1_outputs(4611) <= (layer0_outputs(5665)) xor (layer0_outputs(5721));
    layer1_outputs(4612) <= not(layer0_outputs(1811)) or (layer0_outputs(4202));
    layer1_outputs(4613) <= layer0_outputs(1555);
    layer1_outputs(4614) <= (layer0_outputs(6988)) and (layer0_outputs(3474));
    layer1_outputs(4615) <= '0';
    layer1_outputs(4616) <= not(layer0_outputs(244)) or (layer0_outputs(2129));
    layer1_outputs(4617) <= (layer0_outputs(759)) and (layer0_outputs(2269));
    layer1_outputs(4618) <= not(layer0_outputs(6626));
    layer1_outputs(4619) <= layer0_outputs(7349);
    layer1_outputs(4620) <= not((layer0_outputs(2135)) and (layer0_outputs(7017)));
    layer1_outputs(4621) <= (layer0_outputs(3467)) and not (layer0_outputs(3874));
    layer1_outputs(4622) <= '1';
    layer1_outputs(4623) <= not(layer0_outputs(4840));
    layer1_outputs(4624) <= (layer0_outputs(3281)) and not (layer0_outputs(5336));
    layer1_outputs(4625) <= not(layer0_outputs(1241));
    layer1_outputs(4626) <= not((layer0_outputs(74)) xor (layer0_outputs(4797)));
    layer1_outputs(4627) <= layer0_outputs(7120);
    layer1_outputs(4628) <= (layer0_outputs(6898)) xor (layer0_outputs(5253));
    layer1_outputs(4629) <= (layer0_outputs(4345)) or (layer0_outputs(5740));
    layer1_outputs(4630) <= not((layer0_outputs(2259)) or (layer0_outputs(3195)));
    layer1_outputs(4631) <= (layer0_outputs(837)) and (layer0_outputs(5599));
    layer1_outputs(4632) <= layer0_outputs(3088);
    layer1_outputs(4633) <= '1';
    layer1_outputs(4634) <= layer0_outputs(4298);
    layer1_outputs(4635) <= (layer0_outputs(1355)) or (layer0_outputs(3482));
    layer1_outputs(4636) <= (layer0_outputs(636)) and not (layer0_outputs(5461));
    layer1_outputs(4637) <= not((layer0_outputs(3242)) and (layer0_outputs(7294)));
    layer1_outputs(4638) <= not(layer0_outputs(2882));
    layer1_outputs(4639) <= (layer0_outputs(3959)) and (layer0_outputs(3719));
    layer1_outputs(4640) <= (layer0_outputs(4925)) and not (layer0_outputs(179));
    layer1_outputs(4641) <= not(layer0_outputs(6707));
    layer1_outputs(4642) <= (layer0_outputs(6858)) and (layer0_outputs(3035));
    layer1_outputs(4643) <= not((layer0_outputs(7327)) or (layer0_outputs(264)));
    layer1_outputs(4644) <= not(layer0_outputs(6041)) or (layer0_outputs(4714));
    layer1_outputs(4645) <= not(layer0_outputs(2995)) or (layer0_outputs(798));
    layer1_outputs(4646) <= layer0_outputs(5810);
    layer1_outputs(4647) <= (layer0_outputs(387)) or (layer0_outputs(5201));
    layer1_outputs(4648) <= layer0_outputs(5388);
    layer1_outputs(4649) <= layer0_outputs(2175);
    layer1_outputs(4650) <= '0';
    layer1_outputs(4651) <= not(layer0_outputs(4350)) or (layer0_outputs(5975));
    layer1_outputs(4652) <= (layer0_outputs(193)) and (layer0_outputs(3793));
    layer1_outputs(4653) <= not(layer0_outputs(5614)) or (layer0_outputs(1696));
    layer1_outputs(4654) <= not(layer0_outputs(7266));
    layer1_outputs(4655) <= layer0_outputs(724);
    layer1_outputs(4656) <= not(layer0_outputs(5356));
    layer1_outputs(4657) <= '0';
    layer1_outputs(4658) <= layer0_outputs(4467);
    layer1_outputs(4659) <= layer0_outputs(3617);
    layer1_outputs(4660) <= '1';
    layer1_outputs(4661) <= (layer0_outputs(4542)) and (layer0_outputs(1621));
    layer1_outputs(4662) <= not(layer0_outputs(4974));
    layer1_outputs(4663) <= '1';
    layer1_outputs(4664) <= (layer0_outputs(4605)) and not (layer0_outputs(2354));
    layer1_outputs(4665) <= layer0_outputs(191);
    layer1_outputs(4666) <= not(layer0_outputs(2683));
    layer1_outputs(4667) <= (layer0_outputs(7273)) or (layer0_outputs(4380));
    layer1_outputs(4668) <= layer0_outputs(4086);
    layer1_outputs(4669) <= not(layer0_outputs(628)) or (layer0_outputs(3550));
    layer1_outputs(4670) <= '1';
    layer1_outputs(4671) <= (layer0_outputs(2600)) or (layer0_outputs(3120));
    layer1_outputs(4672) <= not((layer0_outputs(1352)) or (layer0_outputs(86)));
    layer1_outputs(4673) <= not(layer0_outputs(2639)) or (layer0_outputs(7534));
    layer1_outputs(4674) <= '1';
    layer1_outputs(4675) <= not(layer0_outputs(4313)) or (layer0_outputs(2801));
    layer1_outputs(4676) <= (layer0_outputs(6947)) or (layer0_outputs(2761));
    layer1_outputs(4677) <= '0';
    layer1_outputs(4678) <= layer0_outputs(6796);
    layer1_outputs(4679) <= (layer0_outputs(6351)) and (layer0_outputs(5256));
    layer1_outputs(4680) <= not(layer0_outputs(941));
    layer1_outputs(4681) <= not((layer0_outputs(4874)) xor (layer0_outputs(6187)));
    layer1_outputs(4682) <= layer0_outputs(1736);
    layer1_outputs(4683) <= '1';
    layer1_outputs(4684) <= '0';
    layer1_outputs(4685) <= '0';
    layer1_outputs(4686) <= layer0_outputs(4604);
    layer1_outputs(4687) <= (layer0_outputs(3749)) or (layer0_outputs(2458));
    layer1_outputs(4688) <= (layer0_outputs(4474)) xor (layer0_outputs(5685));
    layer1_outputs(4689) <= (layer0_outputs(2819)) and not (layer0_outputs(1796));
    layer1_outputs(4690) <= (layer0_outputs(7342)) and not (layer0_outputs(1992));
    layer1_outputs(4691) <= '0';
    layer1_outputs(4692) <= (layer0_outputs(1866)) or (layer0_outputs(3676));
    layer1_outputs(4693) <= not(layer0_outputs(4031));
    layer1_outputs(4694) <= '1';
    layer1_outputs(4695) <= not((layer0_outputs(3076)) and (layer0_outputs(4170)));
    layer1_outputs(4696) <= (layer0_outputs(5890)) or (layer0_outputs(1868));
    layer1_outputs(4697) <= not((layer0_outputs(114)) or (layer0_outputs(415)));
    layer1_outputs(4698) <= layer0_outputs(7235);
    layer1_outputs(4699) <= not(layer0_outputs(4125));
    layer1_outputs(4700) <= '0';
    layer1_outputs(4701) <= (layer0_outputs(7538)) and not (layer0_outputs(4909));
    layer1_outputs(4702) <= layer0_outputs(5182);
    layer1_outputs(4703) <= not(layer0_outputs(112)) or (layer0_outputs(3850));
    layer1_outputs(4704) <= not((layer0_outputs(3012)) or (layer0_outputs(1857)));
    layer1_outputs(4705) <= layer0_outputs(6026);
    layer1_outputs(4706) <= (layer0_outputs(6314)) and not (layer0_outputs(6958));
    layer1_outputs(4707) <= layer0_outputs(7665);
    layer1_outputs(4708) <= layer0_outputs(4089);
    layer1_outputs(4709) <= (layer0_outputs(2604)) and (layer0_outputs(4259));
    layer1_outputs(4710) <= layer0_outputs(2864);
    layer1_outputs(4711) <= layer0_outputs(5229);
    layer1_outputs(4712) <= not(layer0_outputs(4997));
    layer1_outputs(4713) <= not((layer0_outputs(618)) or (layer0_outputs(7402)));
    layer1_outputs(4714) <= (layer0_outputs(1825)) and (layer0_outputs(6742));
    layer1_outputs(4715) <= not(layer0_outputs(3679));
    layer1_outputs(4716) <= '1';
    layer1_outputs(4717) <= not(layer0_outputs(3758)) or (layer0_outputs(7336));
    layer1_outputs(4718) <= layer0_outputs(2734);
    layer1_outputs(4719) <= (layer0_outputs(21)) and not (layer0_outputs(454));
    layer1_outputs(4720) <= not(layer0_outputs(5641));
    layer1_outputs(4721) <= (layer0_outputs(113)) xor (layer0_outputs(7575));
    layer1_outputs(4722) <= (layer0_outputs(6224)) or (layer0_outputs(1223));
    layer1_outputs(4723) <= not(layer0_outputs(297));
    layer1_outputs(4724) <= (layer0_outputs(5387)) and (layer0_outputs(3697));
    layer1_outputs(4725) <= layer0_outputs(6728);
    layer1_outputs(4726) <= not(layer0_outputs(2945));
    layer1_outputs(4727) <= not((layer0_outputs(5086)) and (layer0_outputs(6712)));
    layer1_outputs(4728) <= layer0_outputs(1068);
    layer1_outputs(4729) <= layer0_outputs(6985);
    layer1_outputs(4730) <= not(layer0_outputs(5722));
    layer1_outputs(4731) <= '1';
    layer1_outputs(4732) <= (layer0_outputs(2274)) and not (layer0_outputs(137));
    layer1_outputs(4733) <= not(layer0_outputs(599));
    layer1_outputs(4734) <= layer0_outputs(1963);
    layer1_outputs(4735) <= not(layer0_outputs(971));
    layer1_outputs(4736) <= layer0_outputs(4799);
    layer1_outputs(4737) <= '1';
    layer1_outputs(4738) <= not(layer0_outputs(4773));
    layer1_outputs(4739) <= '1';
    layer1_outputs(4740) <= not(layer0_outputs(127));
    layer1_outputs(4741) <= not(layer0_outputs(4522)) or (layer0_outputs(4092));
    layer1_outputs(4742) <= '1';
    layer1_outputs(4743) <= not((layer0_outputs(6220)) and (layer0_outputs(5612)));
    layer1_outputs(4744) <= (layer0_outputs(3724)) or (layer0_outputs(2938));
    layer1_outputs(4745) <= '1';
    layer1_outputs(4746) <= layer0_outputs(3772);
    layer1_outputs(4747) <= not((layer0_outputs(2762)) and (layer0_outputs(6409)));
    layer1_outputs(4748) <= '1';
    layer1_outputs(4749) <= not((layer0_outputs(1033)) or (layer0_outputs(7124)));
    layer1_outputs(4750) <= not(layer0_outputs(6181)) or (layer0_outputs(539));
    layer1_outputs(4751) <= (layer0_outputs(3680)) or (layer0_outputs(5502));
    layer1_outputs(4752) <= not((layer0_outputs(4603)) or (layer0_outputs(6150)));
    layer1_outputs(4753) <= not((layer0_outputs(2841)) and (layer0_outputs(5474)));
    layer1_outputs(4754) <= '0';
    layer1_outputs(4755) <= '0';
    layer1_outputs(4756) <= (layer0_outputs(5088)) or (layer0_outputs(7131));
    layer1_outputs(4757) <= layer0_outputs(5783);
    layer1_outputs(4758) <= '1';
    layer1_outputs(4759) <= (layer0_outputs(7286)) and not (layer0_outputs(6290));
    layer1_outputs(4760) <= not(layer0_outputs(6718)) or (layer0_outputs(1727));
    layer1_outputs(4761) <= not(layer0_outputs(203)) or (layer0_outputs(2914));
    layer1_outputs(4762) <= not(layer0_outputs(1387)) or (layer0_outputs(4459));
    layer1_outputs(4763) <= '0';
    layer1_outputs(4764) <= (layer0_outputs(5444)) and not (layer0_outputs(2144));
    layer1_outputs(4765) <= '0';
    layer1_outputs(4766) <= not(layer0_outputs(2280));
    layer1_outputs(4767) <= (layer0_outputs(2082)) xor (layer0_outputs(962));
    layer1_outputs(4768) <= (layer0_outputs(3668)) and not (layer0_outputs(2635));
    layer1_outputs(4769) <= not(layer0_outputs(3952)) or (layer0_outputs(1290));
    layer1_outputs(4770) <= layer0_outputs(1787);
    layer1_outputs(4771) <= '1';
    layer1_outputs(4772) <= layer0_outputs(2887);
    layer1_outputs(4773) <= not(layer0_outputs(1129)) or (layer0_outputs(5452));
    layer1_outputs(4774) <= not((layer0_outputs(3716)) and (layer0_outputs(5069)));
    layer1_outputs(4775) <= not(layer0_outputs(1402));
    layer1_outputs(4776) <= not(layer0_outputs(4318));
    layer1_outputs(4777) <= layer0_outputs(5057);
    layer1_outputs(4778) <= '0';
    layer1_outputs(4779) <= not((layer0_outputs(622)) and (layer0_outputs(1167)));
    layer1_outputs(4780) <= not((layer0_outputs(6942)) xor (layer0_outputs(7042)));
    layer1_outputs(4781) <= (layer0_outputs(3949)) and not (layer0_outputs(3210));
    layer1_outputs(4782) <= (layer0_outputs(4595)) and (layer0_outputs(2836));
    layer1_outputs(4783) <= (layer0_outputs(4722)) or (layer0_outputs(1662));
    layer1_outputs(4784) <= '0';
    layer1_outputs(4785) <= not((layer0_outputs(4419)) and (layer0_outputs(5046)));
    layer1_outputs(4786) <= (layer0_outputs(6234)) and not (layer0_outputs(7486));
    layer1_outputs(4787) <= not((layer0_outputs(3634)) and (layer0_outputs(2699)));
    layer1_outputs(4788) <= not((layer0_outputs(1812)) or (layer0_outputs(3975)));
    layer1_outputs(4789) <= layer0_outputs(1257);
    layer1_outputs(4790) <= not((layer0_outputs(7353)) and (layer0_outputs(400)));
    layer1_outputs(4791) <= not(layer0_outputs(4002));
    layer1_outputs(4792) <= not(layer0_outputs(932));
    layer1_outputs(4793) <= layer0_outputs(5020);
    layer1_outputs(4794) <= (layer0_outputs(3556)) or (layer0_outputs(2218));
    layer1_outputs(4795) <= not((layer0_outputs(3890)) xor (layer0_outputs(5623)));
    layer1_outputs(4796) <= not((layer0_outputs(4508)) xor (layer0_outputs(7409)));
    layer1_outputs(4797) <= (layer0_outputs(1020)) and not (layer0_outputs(7511));
    layer1_outputs(4798) <= layer0_outputs(291);
    layer1_outputs(4799) <= (layer0_outputs(1418)) or (layer0_outputs(5919));
    layer1_outputs(4800) <= not(layer0_outputs(5675)) or (layer0_outputs(5272));
    layer1_outputs(4801) <= not((layer0_outputs(2588)) and (layer0_outputs(1748)));
    layer1_outputs(4802) <= (layer0_outputs(4945)) and not (layer0_outputs(5871));
    layer1_outputs(4803) <= (layer0_outputs(1448)) and not (layer0_outputs(6262));
    layer1_outputs(4804) <= '0';
    layer1_outputs(4805) <= not((layer0_outputs(2598)) and (layer0_outputs(925)));
    layer1_outputs(4806) <= not(layer0_outputs(7291));
    layer1_outputs(4807) <= '1';
    layer1_outputs(4808) <= (layer0_outputs(5111)) and (layer0_outputs(384));
    layer1_outputs(4809) <= '0';
    layer1_outputs(4810) <= (layer0_outputs(5634)) and not (layer0_outputs(4779));
    layer1_outputs(4811) <= not((layer0_outputs(6943)) xor (layer0_outputs(2611)));
    layer1_outputs(4812) <= (layer0_outputs(362)) or (layer0_outputs(957));
    layer1_outputs(4813) <= layer0_outputs(244);
    layer1_outputs(4814) <= '1';
    layer1_outputs(4815) <= (layer0_outputs(1763)) xor (layer0_outputs(2124));
    layer1_outputs(4816) <= (layer0_outputs(4624)) or (layer0_outputs(2853));
    layer1_outputs(4817) <= not(layer0_outputs(3668));
    layer1_outputs(4818) <= (layer0_outputs(1896)) and not (layer0_outputs(4258));
    layer1_outputs(4819) <= (layer0_outputs(3972)) or (layer0_outputs(398));
    layer1_outputs(4820) <= not((layer0_outputs(2279)) or (layer0_outputs(548)));
    layer1_outputs(4821) <= '1';
    layer1_outputs(4822) <= not(layer0_outputs(2862)) or (layer0_outputs(2668));
    layer1_outputs(4823) <= not((layer0_outputs(6390)) xor (layer0_outputs(5561)));
    layer1_outputs(4824) <= (layer0_outputs(7402)) and not (layer0_outputs(5601));
    layer1_outputs(4825) <= not((layer0_outputs(4788)) and (layer0_outputs(4443)));
    layer1_outputs(4826) <= (layer0_outputs(524)) and not (layer0_outputs(7108));
    layer1_outputs(4827) <= not((layer0_outputs(5081)) or (layer0_outputs(5615)));
    layer1_outputs(4828) <= (layer0_outputs(6957)) and not (layer0_outputs(6532));
    layer1_outputs(4829) <= not(layer0_outputs(5709));
    layer1_outputs(4830) <= (layer0_outputs(850)) or (layer0_outputs(4916));
    layer1_outputs(4831) <= not(layer0_outputs(2476)) or (layer0_outputs(2881));
    layer1_outputs(4832) <= not(layer0_outputs(1112));
    layer1_outputs(4833) <= '1';
    layer1_outputs(4834) <= '0';
    layer1_outputs(4835) <= not(layer0_outputs(4431));
    layer1_outputs(4836) <= (layer0_outputs(3948)) and (layer0_outputs(2657));
    layer1_outputs(4837) <= '0';
    layer1_outputs(4838) <= '1';
    layer1_outputs(4839) <= (layer0_outputs(596)) and not (layer0_outputs(6685));
    layer1_outputs(4840) <= (layer0_outputs(3152)) and (layer0_outputs(4306));
    layer1_outputs(4841) <= layer0_outputs(6167);
    layer1_outputs(4842) <= '0';
    layer1_outputs(4843) <= '0';
    layer1_outputs(4844) <= not(layer0_outputs(18));
    layer1_outputs(4845) <= not((layer0_outputs(7079)) and (layer0_outputs(4806)));
    layer1_outputs(4846) <= (layer0_outputs(6084)) and not (layer0_outputs(2340));
    layer1_outputs(4847) <= not((layer0_outputs(807)) and (layer0_outputs(947)));
    layer1_outputs(4848) <= (layer0_outputs(4510)) or (layer0_outputs(2618));
    layer1_outputs(4849) <= not((layer0_outputs(1050)) and (layer0_outputs(3286)));
    layer1_outputs(4850) <= not(layer0_outputs(7479)) or (layer0_outputs(3548));
    layer1_outputs(4851) <= '1';
    layer1_outputs(4852) <= layer0_outputs(2294);
    layer1_outputs(4853) <= (layer0_outputs(6908)) and not (layer0_outputs(3663));
    layer1_outputs(4854) <= not(layer0_outputs(4231)) or (layer0_outputs(4206));
    layer1_outputs(4855) <= layer0_outputs(4833);
    layer1_outputs(4856) <= layer0_outputs(6592);
    layer1_outputs(4857) <= '1';
    layer1_outputs(4858) <= not(layer0_outputs(4802));
    layer1_outputs(4859) <= not(layer0_outputs(7631)) or (layer0_outputs(5814));
    layer1_outputs(4860) <= not((layer0_outputs(6430)) and (layer0_outputs(2521)));
    layer1_outputs(4861) <= not(layer0_outputs(6062)) or (layer0_outputs(6080));
    layer1_outputs(4862) <= not((layer0_outputs(1383)) or (layer0_outputs(4957)));
    layer1_outputs(4863) <= layer0_outputs(6317);
    layer1_outputs(4864) <= not(layer0_outputs(6378)) or (layer0_outputs(6040));
    layer1_outputs(4865) <= not(layer0_outputs(4961)) or (layer0_outputs(4357));
    layer1_outputs(4866) <= '1';
    layer1_outputs(4867) <= layer0_outputs(677);
    layer1_outputs(4868) <= '0';
    layer1_outputs(4869) <= not((layer0_outputs(5293)) and (layer0_outputs(6412)));
    layer1_outputs(4870) <= not(layer0_outputs(2021));
    layer1_outputs(4871) <= (layer0_outputs(4762)) and not (layer0_outputs(553));
    layer1_outputs(4872) <= not(layer0_outputs(5038)) or (layer0_outputs(3562));
    layer1_outputs(4873) <= not(layer0_outputs(5562)) or (layer0_outputs(5653));
    layer1_outputs(4874) <= (layer0_outputs(441)) and (layer0_outputs(7199));
    layer1_outputs(4875) <= layer0_outputs(1361);
    layer1_outputs(4876) <= not(layer0_outputs(6983));
    layer1_outputs(4877) <= layer0_outputs(1573);
    layer1_outputs(4878) <= layer0_outputs(2455);
    layer1_outputs(4879) <= layer0_outputs(4254);
    layer1_outputs(4880) <= (layer0_outputs(3975)) and not (layer0_outputs(7244));
    layer1_outputs(4881) <= not((layer0_outputs(2192)) and (layer0_outputs(6469)));
    layer1_outputs(4882) <= not(layer0_outputs(3810)) or (layer0_outputs(6489));
    layer1_outputs(4883) <= not(layer0_outputs(2902));
    layer1_outputs(4884) <= (layer0_outputs(458)) or (layer0_outputs(7422));
    layer1_outputs(4885) <= '0';
    layer1_outputs(4886) <= (layer0_outputs(74)) and not (layer0_outputs(5829));
    layer1_outputs(4887) <= not(layer0_outputs(7249));
    layer1_outputs(4888) <= (layer0_outputs(6414)) and (layer0_outputs(3885));
    layer1_outputs(4889) <= not(layer0_outputs(6031));
    layer1_outputs(4890) <= (layer0_outputs(3270)) and not (layer0_outputs(3249));
    layer1_outputs(4891) <= (layer0_outputs(281)) and (layer0_outputs(2206));
    layer1_outputs(4892) <= (layer0_outputs(2765)) and not (layer0_outputs(1928));
    layer1_outputs(4893) <= '0';
    layer1_outputs(4894) <= (layer0_outputs(2147)) and not (layer0_outputs(5430));
    layer1_outputs(4895) <= not((layer0_outputs(4106)) or (layer0_outputs(3574)));
    layer1_outputs(4896) <= layer0_outputs(4679);
    layer1_outputs(4897) <= layer0_outputs(6681);
    layer1_outputs(4898) <= layer0_outputs(1658);
    layer1_outputs(4899) <= not(layer0_outputs(2655)) or (layer0_outputs(1909));
    layer1_outputs(4900) <= (layer0_outputs(6206)) and not (layer0_outputs(3104));
    layer1_outputs(4901) <= (layer0_outputs(5016)) and not (layer0_outputs(4204));
    layer1_outputs(4902) <= (layer0_outputs(1416)) or (layer0_outputs(410));
    layer1_outputs(4903) <= not(layer0_outputs(5819));
    layer1_outputs(4904) <= not((layer0_outputs(5858)) and (layer0_outputs(1775)));
    layer1_outputs(4905) <= layer0_outputs(1519);
    layer1_outputs(4906) <= not((layer0_outputs(318)) and (layer0_outputs(6913)));
    layer1_outputs(4907) <= '1';
    layer1_outputs(4908) <= not((layer0_outputs(5635)) or (layer0_outputs(5464)));
    layer1_outputs(4909) <= '0';
    layer1_outputs(4910) <= not(layer0_outputs(6089)) or (layer0_outputs(4552));
    layer1_outputs(4911) <= not(layer0_outputs(1454));
    layer1_outputs(4912) <= (layer0_outputs(3409)) and (layer0_outputs(5718));
    layer1_outputs(4913) <= not(layer0_outputs(2987)) or (layer0_outputs(4823));
    layer1_outputs(4914) <= (layer0_outputs(5609)) and not (layer0_outputs(5048));
    layer1_outputs(4915) <= (layer0_outputs(558)) and not (layer0_outputs(7585));
    layer1_outputs(4916) <= (layer0_outputs(4257)) and not (layer0_outputs(1573));
    layer1_outputs(4917) <= (layer0_outputs(5977)) and (layer0_outputs(6919));
    layer1_outputs(4918) <= '1';
    layer1_outputs(4919) <= not((layer0_outputs(3852)) or (layer0_outputs(854)));
    layer1_outputs(4920) <= not(layer0_outputs(3851));
    layer1_outputs(4921) <= not(layer0_outputs(4076));
    layer1_outputs(4922) <= not(layer0_outputs(1974));
    layer1_outputs(4923) <= '0';
    layer1_outputs(4924) <= not((layer0_outputs(3952)) and (layer0_outputs(5597)));
    layer1_outputs(4925) <= not(layer0_outputs(6094));
    layer1_outputs(4926) <= '0';
    layer1_outputs(4927) <= not(layer0_outputs(2973));
    layer1_outputs(4928) <= layer0_outputs(2656);
    layer1_outputs(4929) <= (layer0_outputs(4449)) and not (layer0_outputs(931));
    layer1_outputs(4930) <= not(layer0_outputs(2183));
    layer1_outputs(4931) <= layer0_outputs(4838);
    layer1_outputs(4932) <= not(layer0_outputs(6744)) or (layer0_outputs(3993));
    layer1_outputs(4933) <= '1';
    layer1_outputs(4934) <= not((layer0_outputs(3908)) or (layer0_outputs(2082)));
    layer1_outputs(4935) <= not(layer0_outputs(5966)) or (layer0_outputs(1663));
    layer1_outputs(4936) <= '1';
    layer1_outputs(4937) <= (layer0_outputs(1137)) xor (layer0_outputs(5626));
    layer1_outputs(4938) <= layer0_outputs(5323);
    layer1_outputs(4939) <= layer0_outputs(5443);
    layer1_outputs(4940) <= not(layer0_outputs(4288));
    layer1_outputs(4941) <= '0';
    layer1_outputs(4942) <= '0';
    layer1_outputs(4943) <= (layer0_outputs(3389)) and not (layer0_outputs(2799));
    layer1_outputs(4944) <= not((layer0_outputs(1230)) or (layer0_outputs(5281)));
    layer1_outputs(4945) <= not(layer0_outputs(3913)) or (layer0_outputs(6657));
    layer1_outputs(4946) <= not(layer0_outputs(4305));
    layer1_outputs(4947) <= not(layer0_outputs(6184)) or (layer0_outputs(4021));
    layer1_outputs(4948) <= not(layer0_outputs(6522)) or (layer0_outputs(4669));
    layer1_outputs(4949) <= not((layer0_outputs(6632)) or (layer0_outputs(2463)));
    layer1_outputs(4950) <= not(layer0_outputs(1713));
    layer1_outputs(4951) <= not(layer0_outputs(3051));
    layer1_outputs(4952) <= not(layer0_outputs(695)) or (layer0_outputs(3258));
    layer1_outputs(4953) <= '0';
    layer1_outputs(4954) <= layer0_outputs(511);
    layer1_outputs(4955) <= (layer0_outputs(6821)) or (layer0_outputs(1098));
    layer1_outputs(4956) <= (layer0_outputs(2815)) and (layer0_outputs(345));
    layer1_outputs(4957) <= not(layer0_outputs(1072)) or (layer0_outputs(5545));
    layer1_outputs(4958) <= (layer0_outputs(84)) and not (layer0_outputs(1697));
    layer1_outputs(4959) <= not(layer0_outputs(3180));
    layer1_outputs(4960) <= layer0_outputs(3519);
    layer1_outputs(4961) <= not(layer0_outputs(2440));
    layer1_outputs(4962) <= not(layer0_outputs(4642));
    layer1_outputs(4963) <= (layer0_outputs(5835)) or (layer0_outputs(815));
    layer1_outputs(4964) <= not((layer0_outputs(608)) or (layer0_outputs(425)));
    layer1_outputs(4965) <= (layer0_outputs(3539)) xor (layer0_outputs(6325));
    layer1_outputs(4966) <= not((layer0_outputs(1369)) and (layer0_outputs(3710)));
    layer1_outputs(4967) <= not(layer0_outputs(397));
    layer1_outputs(4968) <= '0';
    layer1_outputs(4969) <= '1';
    layer1_outputs(4970) <= not(layer0_outputs(1182));
    layer1_outputs(4971) <= (layer0_outputs(5913)) and not (layer0_outputs(1903));
    layer1_outputs(4972) <= not((layer0_outputs(1571)) or (layer0_outputs(113)));
    layer1_outputs(4973) <= '1';
    layer1_outputs(4974) <= '0';
    layer1_outputs(4975) <= layer0_outputs(6799);
    layer1_outputs(4976) <= not(layer0_outputs(5101));
    layer1_outputs(4977) <= layer0_outputs(2125);
    layer1_outputs(4978) <= not((layer0_outputs(4092)) or (layer0_outputs(6091)));
    layer1_outputs(4979) <= '0';
    layer1_outputs(4980) <= (layer0_outputs(5994)) or (layer0_outputs(4061));
    layer1_outputs(4981) <= layer0_outputs(2580);
    layer1_outputs(4982) <= (layer0_outputs(1484)) or (layer0_outputs(7134));
    layer1_outputs(4983) <= not((layer0_outputs(1833)) or (layer0_outputs(6354)));
    layer1_outputs(4984) <= '1';
    layer1_outputs(4985) <= layer0_outputs(2700);
    layer1_outputs(4986) <= not(layer0_outputs(4596));
    layer1_outputs(4987) <= '0';
    layer1_outputs(4988) <= (layer0_outputs(5070)) or (layer0_outputs(6431));
    layer1_outputs(4989) <= '1';
    layer1_outputs(4990) <= (layer0_outputs(3618)) and (layer0_outputs(2344));
    layer1_outputs(4991) <= layer0_outputs(7015);
    layer1_outputs(4992) <= layer0_outputs(303);
    layer1_outputs(4993) <= layer0_outputs(2327);
    layer1_outputs(4994) <= '1';
    layer1_outputs(4995) <= not((layer0_outputs(1494)) and (layer0_outputs(7302)));
    layer1_outputs(4996) <= '1';
    layer1_outputs(4997) <= (layer0_outputs(178)) and not (layer0_outputs(3735));
    layer1_outputs(4998) <= not(layer0_outputs(4734)) or (layer0_outputs(1868));
    layer1_outputs(4999) <= not(layer0_outputs(6193)) or (layer0_outputs(1671));
    layer1_outputs(5000) <= not(layer0_outputs(5903)) or (layer0_outputs(708));
    layer1_outputs(5001) <= not((layer0_outputs(956)) xor (layer0_outputs(5512)));
    layer1_outputs(5002) <= '0';
    layer1_outputs(5003) <= not(layer0_outputs(1262)) or (layer0_outputs(4813));
    layer1_outputs(5004) <= not((layer0_outputs(267)) and (layer0_outputs(5890)));
    layer1_outputs(5005) <= layer0_outputs(865);
    layer1_outputs(5006) <= not(layer0_outputs(6928));
    layer1_outputs(5007) <= '0';
    layer1_outputs(5008) <= layer0_outputs(5196);
    layer1_outputs(5009) <= not(layer0_outputs(3010)) or (layer0_outputs(2064));
    layer1_outputs(5010) <= not((layer0_outputs(2234)) and (layer0_outputs(194)));
    layer1_outputs(5011) <= '0';
    layer1_outputs(5012) <= (layer0_outputs(5928)) and not (layer0_outputs(3412));
    layer1_outputs(5013) <= not((layer0_outputs(6822)) or (layer0_outputs(1333)));
    layer1_outputs(5014) <= not(layer0_outputs(4044)) or (layer0_outputs(5379));
    layer1_outputs(5015) <= not(layer0_outputs(1998));
    layer1_outputs(5016) <= '1';
    layer1_outputs(5017) <= layer0_outputs(3227);
    layer1_outputs(5018) <= (layer0_outputs(7288)) or (layer0_outputs(2823));
    layer1_outputs(5019) <= (layer0_outputs(5956)) and not (layer0_outputs(502));
    layer1_outputs(5020) <= '1';
    layer1_outputs(5021) <= not(layer0_outputs(5375));
    layer1_outputs(5022) <= layer0_outputs(611);
    layer1_outputs(5023) <= not(layer0_outputs(5242)) or (layer0_outputs(928));
    layer1_outputs(5024) <= not(layer0_outputs(3919)) or (layer0_outputs(1905));
    layer1_outputs(5025) <= layer0_outputs(1087);
    layer1_outputs(5026) <= '1';
    layer1_outputs(5027) <= layer0_outputs(2893);
    layer1_outputs(5028) <= not(layer0_outputs(3054));
    layer1_outputs(5029) <= '1';
    layer1_outputs(5030) <= not(layer0_outputs(2903)) or (layer0_outputs(7344));
    layer1_outputs(5031) <= not(layer0_outputs(3436)) or (layer0_outputs(1379));
    layer1_outputs(5032) <= (layer0_outputs(3850)) and (layer0_outputs(6477));
    layer1_outputs(5033) <= (layer0_outputs(1368)) and not (layer0_outputs(4517));
    layer1_outputs(5034) <= not(layer0_outputs(2829)) or (layer0_outputs(5485));
    layer1_outputs(5035) <= (layer0_outputs(836)) and not (layer0_outputs(7505));
    layer1_outputs(5036) <= (layer0_outputs(5492)) and not (layer0_outputs(2377));
    layer1_outputs(5037) <= (layer0_outputs(83)) and not (layer0_outputs(2909));
    layer1_outputs(5038) <= (layer0_outputs(3677)) or (layer0_outputs(52));
    layer1_outputs(5039) <= (layer0_outputs(118)) and not (layer0_outputs(814));
    layer1_outputs(5040) <= '1';
    layer1_outputs(5041) <= (layer0_outputs(2336)) and not (layer0_outputs(1681));
    layer1_outputs(5042) <= (layer0_outputs(6869)) or (layer0_outputs(1746));
    layer1_outputs(5043) <= not(layer0_outputs(4269));
    layer1_outputs(5044) <= '1';
    layer1_outputs(5045) <= (layer0_outputs(5948)) and (layer0_outputs(6617));
    layer1_outputs(5046) <= (layer0_outputs(2314)) or (layer0_outputs(2974));
    layer1_outputs(5047) <= '0';
    layer1_outputs(5048) <= not((layer0_outputs(2890)) and (layer0_outputs(3380)));
    layer1_outputs(5049) <= (layer0_outputs(153)) and not (layer0_outputs(682));
    layer1_outputs(5050) <= not(layer0_outputs(732)) or (layer0_outputs(721));
    layer1_outputs(5051) <= not(layer0_outputs(1557)) or (layer0_outputs(1184));
    layer1_outputs(5052) <= not(layer0_outputs(7011));
    layer1_outputs(5053) <= (layer0_outputs(4515)) and (layer0_outputs(2117));
    layer1_outputs(5054) <= (layer0_outputs(1423)) and not (layer0_outputs(5252));
    layer1_outputs(5055) <= (layer0_outputs(1682)) and not (layer0_outputs(5720));
    layer1_outputs(5056) <= layer0_outputs(6536);
    layer1_outputs(5057) <= '1';
    layer1_outputs(5058) <= '0';
    layer1_outputs(5059) <= layer0_outputs(5488);
    layer1_outputs(5060) <= (layer0_outputs(4966)) and not (layer0_outputs(7147));
    layer1_outputs(5061) <= layer0_outputs(4543);
    layer1_outputs(5062) <= not(layer0_outputs(4332));
    layer1_outputs(5063) <= not(layer0_outputs(774)) or (layer0_outputs(4071));
    layer1_outputs(5064) <= (layer0_outputs(5307)) and not (layer0_outputs(7577));
    layer1_outputs(5065) <= (layer0_outputs(1090)) and not (layer0_outputs(2403));
    layer1_outputs(5066) <= not((layer0_outputs(3078)) or (layer0_outputs(2264)));
    layer1_outputs(5067) <= not(layer0_outputs(7123)) or (layer0_outputs(1738));
    layer1_outputs(5068) <= not(layer0_outputs(6461)) or (layer0_outputs(3460));
    layer1_outputs(5069) <= (layer0_outputs(2941)) and (layer0_outputs(6398));
    layer1_outputs(5070) <= (layer0_outputs(259)) and not (layer0_outputs(6809));
    layer1_outputs(5071) <= '0';
    layer1_outputs(5072) <= layer0_outputs(4267);
    layer1_outputs(5073) <= not(layer0_outputs(3348)) or (layer0_outputs(7499));
    layer1_outputs(5074) <= '0';
    layer1_outputs(5075) <= (layer0_outputs(3413)) and not (layer0_outputs(5958));
    layer1_outputs(5076) <= not(layer0_outputs(7228)) or (layer0_outputs(7162));
    layer1_outputs(5077) <= (layer0_outputs(3984)) and not (layer0_outputs(7437));
    layer1_outputs(5078) <= layer0_outputs(7184);
    layer1_outputs(5079) <= '0';
    layer1_outputs(5080) <= (layer0_outputs(2167)) and not (layer0_outputs(3819));
    layer1_outputs(5081) <= layer0_outputs(4877);
    layer1_outputs(5082) <= (layer0_outputs(7165)) and not (layer0_outputs(6915));
    layer1_outputs(5083) <= not(layer0_outputs(7214));
    layer1_outputs(5084) <= layer0_outputs(301);
    layer1_outputs(5085) <= layer0_outputs(4948);
    layer1_outputs(5086) <= not(layer0_outputs(2745)) or (layer0_outputs(3382));
    layer1_outputs(5087) <= layer0_outputs(306);
    layer1_outputs(5088) <= not((layer0_outputs(109)) xor (layer0_outputs(2816)));
    layer1_outputs(5089) <= '1';
    layer1_outputs(5090) <= not(layer0_outputs(3660));
    layer1_outputs(5091) <= layer0_outputs(5100);
    layer1_outputs(5092) <= '1';
    layer1_outputs(5093) <= (layer0_outputs(6093)) and (layer0_outputs(3577));
    layer1_outputs(5094) <= layer0_outputs(4213);
    layer1_outputs(5095) <= layer0_outputs(504);
    layer1_outputs(5096) <= '1';
    layer1_outputs(5097) <= not(layer0_outputs(2530));
    layer1_outputs(5098) <= not(layer0_outputs(2077));
    layer1_outputs(5099) <= '0';
    layer1_outputs(5100) <= '0';
    layer1_outputs(5101) <= '0';
    layer1_outputs(5102) <= not(layer0_outputs(6065)) or (layer0_outputs(1294));
    layer1_outputs(5103) <= (layer0_outputs(2522)) and (layer0_outputs(7665));
    layer1_outputs(5104) <= layer0_outputs(1747);
    layer1_outputs(5105) <= not(layer0_outputs(5153));
    layer1_outputs(5106) <= (layer0_outputs(2451)) and not (layer0_outputs(6413));
    layer1_outputs(5107) <= (layer0_outputs(37)) and (layer0_outputs(4433));
    layer1_outputs(5108) <= '1';
    layer1_outputs(5109) <= not((layer0_outputs(134)) or (layer0_outputs(758)));
    layer1_outputs(5110) <= not((layer0_outputs(4152)) and (layer0_outputs(4578)));
    layer1_outputs(5111) <= '1';
    layer1_outputs(5112) <= layer0_outputs(2474);
    layer1_outputs(5113) <= not(layer0_outputs(5880)) or (layer0_outputs(5814));
    layer1_outputs(5114) <= layer0_outputs(4945);
    layer1_outputs(5115) <= '1';
    layer1_outputs(5116) <= not(layer0_outputs(4572));
    layer1_outputs(5117) <= layer0_outputs(5124);
    layer1_outputs(5118) <= not(layer0_outputs(5595));
    layer1_outputs(5119) <= '1';
    layer1_outputs(5120) <= not(layer0_outputs(110));
    layer1_outputs(5121) <= layer0_outputs(4491);
    layer1_outputs(5122) <= '0';
    layer1_outputs(5123) <= layer0_outputs(6360);
    layer1_outputs(5124) <= layer0_outputs(2354);
    layer1_outputs(5125) <= not(layer0_outputs(6597)) or (layer0_outputs(3440));
    layer1_outputs(5126) <= not(layer0_outputs(6002));
    layer1_outputs(5127) <= (layer0_outputs(6663)) and (layer0_outputs(827));
    layer1_outputs(5128) <= (layer0_outputs(3348)) and not (layer0_outputs(5918));
    layer1_outputs(5129) <= not((layer0_outputs(2006)) and (layer0_outputs(1759)));
    layer1_outputs(5130) <= not(layer0_outputs(314));
    layer1_outputs(5131) <= layer0_outputs(6934);
    layer1_outputs(5132) <= '0';
    layer1_outputs(5133) <= not((layer0_outputs(2020)) or (layer0_outputs(4497)));
    layer1_outputs(5134) <= layer0_outputs(4947);
    layer1_outputs(5135) <= (layer0_outputs(775)) and not (layer0_outputs(4195));
    layer1_outputs(5136) <= not((layer0_outputs(6751)) or (layer0_outputs(2484)));
    layer1_outputs(5137) <= not((layer0_outputs(2730)) xor (layer0_outputs(1177)));
    layer1_outputs(5138) <= layer0_outputs(4652);
    layer1_outputs(5139) <= '1';
    layer1_outputs(5140) <= layer0_outputs(1261);
    layer1_outputs(5141) <= layer0_outputs(2426);
    layer1_outputs(5142) <= layer0_outputs(5957);
    layer1_outputs(5143) <= (layer0_outputs(3734)) and not (layer0_outputs(4290));
    layer1_outputs(5144) <= layer0_outputs(3991);
    layer1_outputs(5145) <= (layer0_outputs(1052)) xor (layer0_outputs(3963));
    layer1_outputs(5146) <= layer0_outputs(1430);
    layer1_outputs(5147) <= not(layer0_outputs(3144));
    layer1_outputs(5148) <= not(layer0_outputs(83));
    layer1_outputs(5149) <= not((layer0_outputs(5157)) xor (layer0_outputs(6033)));
    layer1_outputs(5150) <= (layer0_outputs(6091)) and (layer0_outputs(425));
    layer1_outputs(5151) <= (layer0_outputs(92)) xor (layer0_outputs(3377));
    layer1_outputs(5152) <= (layer0_outputs(6523)) and not (layer0_outputs(171));
    layer1_outputs(5153) <= layer0_outputs(1254);
    layer1_outputs(5154) <= not(layer0_outputs(7041));
    layer1_outputs(5155) <= layer0_outputs(385);
    layer1_outputs(5156) <= (layer0_outputs(3311)) and not (layer0_outputs(6047));
    layer1_outputs(5157) <= not(layer0_outputs(5211));
    layer1_outputs(5158) <= (layer0_outputs(2337)) and not (layer0_outputs(3511));
    layer1_outputs(5159) <= (layer0_outputs(5252)) xor (layer0_outputs(2320));
    layer1_outputs(5160) <= (layer0_outputs(4078)) and not (layer0_outputs(3530));
    layer1_outputs(5161) <= (layer0_outputs(5052)) and (layer0_outputs(5089));
    layer1_outputs(5162) <= not(layer0_outputs(4490)) or (layer0_outputs(3549));
    layer1_outputs(5163) <= not(layer0_outputs(7033)) or (layer0_outputs(1392));
    layer1_outputs(5164) <= '1';
    layer1_outputs(5165) <= not((layer0_outputs(7472)) and (layer0_outputs(2098)));
    layer1_outputs(5166) <= not(layer0_outputs(3483));
    layer1_outputs(5167) <= not(layer0_outputs(5806)) or (layer0_outputs(6058));
    layer1_outputs(5168) <= not((layer0_outputs(5791)) xor (layer0_outputs(3848)));
    layer1_outputs(5169) <= '1';
    layer1_outputs(5170) <= not(layer0_outputs(6968)) or (layer0_outputs(3625));
    layer1_outputs(5171) <= layer0_outputs(738);
    layer1_outputs(5172) <= not((layer0_outputs(7632)) or (layer0_outputs(527)));
    layer1_outputs(5173) <= not((layer0_outputs(2258)) and (layer0_outputs(1914)));
    layer1_outputs(5174) <= '1';
    layer1_outputs(5175) <= (layer0_outputs(6777)) and not (layer0_outputs(7196));
    layer1_outputs(5176) <= not(layer0_outputs(755));
    layer1_outputs(5177) <= (layer0_outputs(2394)) or (layer0_outputs(1400));
    layer1_outputs(5178) <= layer0_outputs(1806);
    layer1_outputs(5179) <= not(layer0_outputs(2886));
    layer1_outputs(5180) <= layer0_outputs(6778);
    layer1_outputs(5181) <= not(layer0_outputs(3374));
    layer1_outputs(5182) <= layer0_outputs(2264);
    layer1_outputs(5183) <= layer0_outputs(1229);
    layer1_outputs(5184) <= layer0_outputs(5631);
    layer1_outputs(5185) <= not(layer0_outputs(6953));
    layer1_outputs(5186) <= layer0_outputs(4712);
    layer1_outputs(5187) <= not(layer0_outputs(4954));
    layer1_outputs(5188) <= (layer0_outputs(4410)) or (layer0_outputs(5457));
    layer1_outputs(5189) <= layer0_outputs(6038);
    layer1_outputs(5190) <= not(layer0_outputs(7547)) or (layer0_outputs(5897));
    layer1_outputs(5191) <= '0';
    layer1_outputs(5192) <= not(layer0_outputs(1343));
    layer1_outputs(5193) <= not((layer0_outputs(1549)) or (layer0_outputs(2583)));
    layer1_outputs(5194) <= layer0_outputs(4413);
    layer1_outputs(5195) <= not((layer0_outputs(5698)) or (layer0_outputs(1491)));
    layer1_outputs(5196) <= '0';
    layer1_outputs(5197) <= not(layer0_outputs(2714));
    layer1_outputs(5198) <= layer0_outputs(6310);
    layer1_outputs(5199) <= layer0_outputs(6557);
    layer1_outputs(5200) <= not(layer0_outputs(218)) or (layer0_outputs(6373));
    layer1_outputs(5201) <= '1';
    layer1_outputs(5202) <= layer0_outputs(235);
    layer1_outputs(5203) <= not(layer0_outputs(2809));
    layer1_outputs(5204) <= '1';
    layer1_outputs(5205) <= not((layer0_outputs(5854)) or (layer0_outputs(7341)));
    layer1_outputs(5206) <= (layer0_outputs(455)) and (layer0_outputs(6818));
    layer1_outputs(5207) <= layer0_outputs(2731);
    layer1_outputs(5208) <= not(layer0_outputs(508));
    layer1_outputs(5209) <= not(layer0_outputs(327));
    layer1_outputs(5210) <= layer0_outputs(3680);
    layer1_outputs(5211) <= '1';
    layer1_outputs(5212) <= not(layer0_outputs(5677)) or (layer0_outputs(6381));
    layer1_outputs(5213) <= not((layer0_outputs(7606)) or (layer0_outputs(1709)));
    layer1_outputs(5214) <= not(layer0_outputs(7375));
    layer1_outputs(5215) <= not((layer0_outputs(3659)) or (layer0_outputs(808)));
    layer1_outputs(5216) <= not((layer0_outputs(885)) or (layer0_outputs(386)));
    layer1_outputs(5217) <= '0';
    layer1_outputs(5218) <= layer0_outputs(3540);
    layer1_outputs(5219) <= (layer0_outputs(7493)) and not (layer0_outputs(5107));
    layer1_outputs(5220) <= not((layer0_outputs(4891)) and (layer0_outputs(3461)));
    layer1_outputs(5221) <= (layer0_outputs(2478)) or (layer0_outputs(1931));
    layer1_outputs(5222) <= not(layer0_outputs(6727)) or (layer0_outputs(2895));
    layer1_outputs(5223) <= '1';
    layer1_outputs(5224) <= '0';
    layer1_outputs(5225) <= '0';
    layer1_outputs(5226) <= layer0_outputs(6565);
    layer1_outputs(5227) <= '1';
    layer1_outputs(5228) <= '0';
    layer1_outputs(5229) <= layer0_outputs(2139);
    layer1_outputs(5230) <= not(layer0_outputs(7167));
    layer1_outputs(5231) <= '0';
    layer1_outputs(5232) <= '1';
    layer1_outputs(5233) <= (layer0_outputs(1160)) xor (layer0_outputs(714));
    layer1_outputs(5234) <= not(layer0_outputs(6824)) or (layer0_outputs(5445));
    layer1_outputs(5235) <= '0';
    layer1_outputs(5236) <= '0';
    layer1_outputs(5237) <= '0';
    layer1_outputs(5238) <= layer0_outputs(3666);
    layer1_outputs(5239) <= '1';
    layer1_outputs(5240) <= not(layer0_outputs(5580)) or (layer0_outputs(4702));
    layer1_outputs(5241) <= not(layer0_outputs(4407));
    layer1_outputs(5242) <= not(layer0_outputs(1084)) or (layer0_outputs(7460));
    layer1_outputs(5243) <= '0';
    layer1_outputs(5244) <= not(layer0_outputs(7244));
    layer1_outputs(5245) <= not(layer0_outputs(334)) or (layer0_outputs(2792));
    layer1_outputs(5246) <= layer0_outputs(1119);
    layer1_outputs(5247) <= (layer0_outputs(3003)) or (layer0_outputs(7500));
    layer1_outputs(5248) <= (layer0_outputs(4545)) and not (layer0_outputs(6181));
    layer1_outputs(5249) <= not(layer0_outputs(4752)) or (layer0_outputs(3457));
    layer1_outputs(5250) <= not(layer0_outputs(6813));
    layer1_outputs(5251) <= not(layer0_outputs(2679));
    layer1_outputs(5252) <= layer0_outputs(7061);
    layer1_outputs(5253) <= not(layer0_outputs(3802)) or (layer0_outputs(1281));
    layer1_outputs(5254) <= layer0_outputs(140);
    layer1_outputs(5255) <= '0';
    layer1_outputs(5256) <= not(layer0_outputs(5358));
    layer1_outputs(5257) <= layer0_outputs(7044);
    layer1_outputs(5258) <= not((layer0_outputs(3974)) or (layer0_outputs(1365)));
    layer1_outputs(5259) <= not((layer0_outputs(3951)) or (layer0_outputs(4237)));
    layer1_outputs(5260) <= not(layer0_outputs(1481));
    layer1_outputs(5261) <= '1';
    layer1_outputs(5262) <= not((layer0_outputs(6974)) or (layer0_outputs(1444)));
    layer1_outputs(5263) <= (layer0_outputs(3578)) and not (layer0_outputs(5203));
    layer1_outputs(5264) <= not(layer0_outputs(7031)) or (layer0_outputs(2753));
    layer1_outputs(5265) <= layer0_outputs(1266);
    layer1_outputs(5266) <= not(layer0_outputs(1001));
    layer1_outputs(5267) <= not(layer0_outputs(7156)) or (layer0_outputs(1141));
    layer1_outputs(5268) <= not(layer0_outputs(463)) or (layer0_outputs(6523));
    layer1_outputs(5269) <= not(layer0_outputs(4384));
    layer1_outputs(5270) <= '1';
    layer1_outputs(5271) <= (layer0_outputs(3186)) and not (layer0_outputs(5284));
    layer1_outputs(5272) <= not((layer0_outputs(1059)) or (layer0_outputs(5017)));
    layer1_outputs(5273) <= (layer0_outputs(4372)) and (layer0_outputs(1161));
    layer1_outputs(5274) <= layer0_outputs(2670);
    layer1_outputs(5275) <= (layer0_outputs(5769)) or (layer0_outputs(5064));
    layer1_outputs(5276) <= not(layer0_outputs(5749));
    layer1_outputs(5277) <= (layer0_outputs(4643)) or (layer0_outputs(519));
    layer1_outputs(5278) <= (layer0_outputs(203)) or (layer0_outputs(3267));
    layer1_outputs(5279) <= not((layer0_outputs(7034)) or (layer0_outputs(1505)));
    layer1_outputs(5280) <= not(layer0_outputs(5976));
    layer1_outputs(5281) <= '0';
    layer1_outputs(5282) <= '1';
    layer1_outputs(5283) <= (layer0_outputs(4122)) and (layer0_outputs(6752));
    layer1_outputs(5284) <= layer0_outputs(1279);
    layer1_outputs(5285) <= '0';
    layer1_outputs(5286) <= (layer0_outputs(3388)) and not (layer0_outputs(7437));
    layer1_outputs(5287) <= (layer0_outputs(2083)) and (layer0_outputs(1817));
    layer1_outputs(5288) <= layer0_outputs(308);
    layer1_outputs(5289) <= layer0_outputs(2049);
    layer1_outputs(5290) <= not(layer0_outputs(2312));
    layer1_outputs(5291) <= (layer0_outputs(5019)) and not (layer0_outputs(654));
    layer1_outputs(5292) <= not((layer0_outputs(6797)) xor (layer0_outputs(3402)));
    layer1_outputs(5293) <= not(layer0_outputs(4215));
    layer1_outputs(5294) <= not((layer0_outputs(3285)) and (layer0_outputs(7072)));
    layer1_outputs(5295) <= not((layer0_outputs(736)) and (layer0_outputs(7297)));
    layer1_outputs(5296) <= not(layer0_outputs(3475));
    layer1_outputs(5297) <= not(layer0_outputs(3687));
    layer1_outputs(5298) <= not(layer0_outputs(2908));
    layer1_outputs(5299) <= not(layer0_outputs(1698)) or (layer0_outputs(1116));
    layer1_outputs(5300) <= layer0_outputs(6634);
    layer1_outputs(5301) <= '0';
    layer1_outputs(5302) <= '0';
    layer1_outputs(5303) <= (layer0_outputs(3247)) and not (layer0_outputs(5385));
    layer1_outputs(5304) <= layer0_outputs(2532);
    layer1_outputs(5305) <= not((layer0_outputs(4261)) and (layer0_outputs(1618)));
    layer1_outputs(5306) <= not((layer0_outputs(2701)) or (layer0_outputs(6936)));
    layer1_outputs(5307) <= not(layer0_outputs(5065)) or (layer0_outputs(4439));
    layer1_outputs(5308) <= (layer0_outputs(3695)) and (layer0_outputs(1264));
    layer1_outputs(5309) <= not(layer0_outputs(3278));
    layer1_outputs(5310) <= not((layer0_outputs(6361)) and (layer0_outputs(3109)));
    layer1_outputs(5311) <= layer0_outputs(4353);
    layer1_outputs(5312) <= layer0_outputs(7661);
    layer1_outputs(5313) <= not(layer0_outputs(549)) or (layer0_outputs(2615));
    layer1_outputs(5314) <= not((layer0_outputs(375)) and (layer0_outputs(2733)));
    layer1_outputs(5315) <= not((layer0_outputs(4369)) and (layer0_outputs(2669)));
    layer1_outputs(5316) <= (layer0_outputs(5586)) and not (layer0_outputs(6545));
    layer1_outputs(5317) <= not((layer0_outputs(7080)) or (layer0_outputs(6783)));
    layer1_outputs(5318) <= not((layer0_outputs(1827)) and (layer0_outputs(4140)));
    layer1_outputs(5319) <= (layer0_outputs(602)) and not (layer0_outputs(135));
    layer1_outputs(5320) <= not(layer0_outputs(436)) or (layer0_outputs(399));
    layer1_outputs(5321) <= (layer0_outputs(1985)) and (layer0_outputs(5257));
    layer1_outputs(5322) <= '0';
    layer1_outputs(5323) <= not(layer0_outputs(3961)) or (layer0_outputs(3366));
    layer1_outputs(5324) <= (layer0_outputs(2836)) and (layer0_outputs(3696));
    layer1_outputs(5325) <= layer0_outputs(1044);
    layer1_outputs(5326) <= not(layer0_outputs(1846));
    layer1_outputs(5327) <= not(layer0_outputs(5716)) or (layer0_outputs(1772));
    layer1_outputs(5328) <= not((layer0_outputs(6022)) or (layer0_outputs(2362)));
    layer1_outputs(5329) <= (layer0_outputs(7030)) and (layer0_outputs(5842));
    layer1_outputs(5330) <= '0';
    layer1_outputs(5331) <= not((layer0_outputs(2370)) and (layer0_outputs(4980)));
    layer1_outputs(5332) <= not(layer0_outputs(4393));
    layer1_outputs(5333) <= layer0_outputs(1637);
    layer1_outputs(5334) <= not((layer0_outputs(7528)) and (layer0_outputs(1111)));
    layer1_outputs(5335) <= '1';
    layer1_outputs(5336) <= layer0_outputs(3565);
    layer1_outputs(5337) <= not(layer0_outputs(2518)) or (layer0_outputs(5078));
    layer1_outputs(5338) <= '1';
    layer1_outputs(5339) <= (layer0_outputs(7314)) and not (layer0_outputs(2890));
    layer1_outputs(5340) <= (layer0_outputs(7345)) or (layer0_outputs(5114));
    layer1_outputs(5341) <= layer0_outputs(3184);
    layer1_outputs(5342) <= not((layer0_outputs(3988)) xor (layer0_outputs(4161)));
    layer1_outputs(5343) <= not(layer0_outputs(4905)) or (layer0_outputs(2802));
    layer1_outputs(5344) <= (layer0_outputs(3989)) or (layer0_outputs(305));
    layer1_outputs(5345) <= layer0_outputs(4161);
    layer1_outputs(5346) <= '1';
    layer1_outputs(5347) <= not(layer0_outputs(6588));
    layer1_outputs(5348) <= '1';
    layer1_outputs(5349) <= not(layer0_outputs(1971));
    layer1_outputs(5350) <= (layer0_outputs(5902)) or (layer0_outputs(1196));
    layer1_outputs(5351) <= (layer0_outputs(6136)) or (layer0_outputs(4189));
    layer1_outputs(5352) <= layer0_outputs(5289);
    layer1_outputs(5353) <= layer0_outputs(393);
    layer1_outputs(5354) <= layer0_outputs(4817);
    layer1_outputs(5355) <= (layer0_outputs(5993)) and (layer0_outputs(3022));
    layer1_outputs(5356) <= layer0_outputs(358);
    layer1_outputs(5357) <= not(layer0_outputs(2869));
    layer1_outputs(5358) <= not(layer0_outputs(1559));
    layer1_outputs(5359) <= (layer0_outputs(4098)) or (layer0_outputs(440));
    layer1_outputs(5360) <= '1';
    layer1_outputs(5361) <= not(layer0_outputs(4043)) or (layer0_outputs(2876));
    layer1_outputs(5362) <= layer0_outputs(6130);
    layer1_outputs(5363) <= (layer0_outputs(5522)) xor (layer0_outputs(6821));
    layer1_outputs(5364) <= not(layer0_outputs(1717));
    layer1_outputs(5365) <= not(layer0_outputs(3176)) or (layer0_outputs(3284));
    layer1_outputs(5366) <= not(layer0_outputs(6088)) or (layer0_outputs(1640));
    layer1_outputs(5367) <= not((layer0_outputs(6710)) xor (layer0_outputs(2489)));
    layer1_outputs(5368) <= not(layer0_outputs(6843));
    layer1_outputs(5369) <= not(layer0_outputs(346));
    layer1_outputs(5370) <= not(layer0_outputs(1550));
    layer1_outputs(5371) <= layer0_outputs(3315);
    layer1_outputs(5372) <= not((layer0_outputs(2439)) xor (layer0_outputs(2668)));
    layer1_outputs(5373) <= '0';
    layer1_outputs(5374) <= not(layer0_outputs(7227)) or (layer0_outputs(2027));
    layer1_outputs(5375) <= not((layer0_outputs(7085)) and (layer0_outputs(319)));
    layer1_outputs(5376) <= not(layer0_outputs(428)) or (layer0_outputs(1830));
    layer1_outputs(5377) <= not((layer0_outputs(4348)) or (layer0_outputs(1344)));
    layer1_outputs(5378) <= layer0_outputs(7560);
    layer1_outputs(5379) <= not(layer0_outputs(227)) or (layer0_outputs(5799));
    layer1_outputs(5380) <= not(layer0_outputs(6797)) or (layer0_outputs(3275));
    layer1_outputs(5381) <= not(layer0_outputs(4296));
    layer1_outputs(5382) <= not(layer0_outputs(4405)) or (layer0_outputs(3694));
    layer1_outputs(5383) <= '0';
    layer1_outputs(5384) <= (layer0_outputs(6749)) and not (layer0_outputs(913));
    layer1_outputs(5385) <= layer0_outputs(7319);
    layer1_outputs(5386) <= not(layer0_outputs(6661));
    layer1_outputs(5387) <= not(layer0_outputs(4079));
    layer1_outputs(5388) <= (layer0_outputs(7117)) or (layer0_outputs(4079));
    layer1_outputs(5389) <= '1';
    layer1_outputs(5390) <= not(layer0_outputs(1154)) or (layer0_outputs(6781));
    layer1_outputs(5391) <= '1';
    layer1_outputs(5392) <= layer0_outputs(3203);
    layer1_outputs(5393) <= (layer0_outputs(6895)) or (layer0_outputs(3217));
    layer1_outputs(5394) <= (layer0_outputs(1255)) and not (layer0_outputs(6472));
    layer1_outputs(5395) <= (layer0_outputs(2738)) or (layer0_outputs(3623));
    layer1_outputs(5396) <= layer0_outputs(6884);
    layer1_outputs(5397) <= '0';
    layer1_outputs(5398) <= layer0_outputs(2667);
    layer1_outputs(5399) <= (layer0_outputs(802)) and (layer0_outputs(5209));
    layer1_outputs(5400) <= not(layer0_outputs(1530)) or (layer0_outputs(5983));
    layer1_outputs(5401) <= '0';
    layer1_outputs(5402) <= '1';
    layer1_outputs(5403) <= '0';
    layer1_outputs(5404) <= (layer0_outputs(4575)) and not (layer0_outputs(6114));
    layer1_outputs(5405) <= (layer0_outputs(5195)) and not (layer0_outputs(5119));
    layer1_outputs(5406) <= (layer0_outputs(1229)) and (layer0_outputs(2931));
    layer1_outputs(5407) <= (layer0_outputs(3824)) or (layer0_outputs(5001));
    layer1_outputs(5408) <= (layer0_outputs(2307)) and not (layer0_outputs(3695));
    layer1_outputs(5409) <= '1';
    layer1_outputs(5410) <= '0';
    layer1_outputs(5411) <= '0';
    layer1_outputs(5412) <= '0';
    layer1_outputs(5413) <= not(layer0_outputs(6481)) or (layer0_outputs(6273));
    layer1_outputs(5414) <= not(layer0_outputs(211)) or (layer0_outputs(1419));
    layer1_outputs(5415) <= not((layer0_outputs(3334)) or (layer0_outputs(2207)));
    layer1_outputs(5416) <= not(layer0_outputs(6761));
    layer1_outputs(5417) <= (layer0_outputs(2600)) and not (layer0_outputs(629));
    layer1_outputs(5418) <= layer0_outputs(6098);
    layer1_outputs(5419) <= not((layer0_outputs(6164)) or (layer0_outputs(401)));
    layer1_outputs(5420) <= (layer0_outputs(3120)) and not (layer0_outputs(1953));
    layer1_outputs(5421) <= not(layer0_outputs(7376)) or (layer0_outputs(4420));
    layer1_outputs(5422) <= layer0_outputs(5635);
    layer1_outputs(5423) <= layer0_outputs(5771);
    layer1_outputs(5424) <= '1';
    layer1_outputs(5425) <= (layer0_outputs(5638)) and not (layer0_outputs(2918));
    layer1_outputs(5426) <= (layer0_outputs(6147)) and not (layer0_outputs(7305));
    layer1_outputs(5427) <= (layer0_outputs(2457)) and not (layer0_outputs(2319));
    layer1_outputs(5428) <= not(layer0_outputs(4614));
    layer1_outputs(5429) <= layer0_outputs(6359);
    layer1_outputs(5430) <= '0';
    layer1_outputs(5431) <= '1';
    layer1_outputs(5432) <= not(layer0_outputs(660));
    layer1_outputs(5433) <= not(layer0_outputs(291));
    layer1_outputs(5434) <= not(layer0_outputs(1222)) or (layer0_outputs(1997));
    layer1_outputs(5435) <= '1';
    layer1_outputs(5436) <= (layer0_outputs(4003)) and not (layer0_outputs(4499));
    layer1_outputs(5437) <= (layer0_outputs(101)) and not (layer0_outputs(3518));
    layer1_outputs(5438) <= layer0_outputs(4811);
    layer1_outputs(5439) <= layer0_outputs(4463);
    layer1_outputs(5440) <= not((layer0_outputs(1583)) and (layer0_outputs(7679)));
    layer1_outputs(5441) <= layer0_outputs(3110);
    layer1_outputs(5442) <= layer0_outputs(961);
    layer1_outputs(5443) <= not(layer0_outputs(726));
    layer1_outputs(5444) <= not(layer0_outputs(6332));
    layer1_outputs(5445) <= (layer0_outputs(3380)) and not (layer0_outputs(4513));
    layer1_outputs(5446) <= (layer0_outputs(7674)) and not (layer0_outputs(7481));
    layer1_outputs(5447) <= layer0_outputs(7291);
    layer1_outputs(5448) <= (layer0_outputs(30)) and (layer0_outputs(1500));
    layer1_outputs(5449) <= not(layer0_outputs(2011)) or (layer0_outputs(1335));
    layer1_outputs(5450) <= not((layer0_outputs(6356)) and (layer0_outputs(6698)));
    layer1_outputs(5451) <= not(layer0_outputs(7640));
    layer1_outputs(5452) <= '0';
    layer1_outputs(5453) <= (layer0_outputs(7127)) or (layer0_outputs(4243));
    layer1_outputs(5454) <= (layer0_outputs(7139)) or (layer0_outputs(1178));
    layer1_outputs(5455) <= '1';
    layer1_outputs(5456) <= layer0_outputs(3809);
    layer1_outputs(5457) <= not(layer0_outputs(2002));
    layer1_outputs(5458) <= not(layer0_outputs(6754));
    layer1_outputs(5459) <= layer0_outputs(4943);
    layer1_outputs(5460) <= layer0_outputs(2059);
    layer1_outputs(5461) <= not((layer0_outputs(2248)) and (layer0_outputs(4778)));
    layer1_outputs(5462) <= (layer0_outputs(319)) or (layer0_outputs(4689));
    layer1_outputs(5463) <= (layer0_outputs(3630)) xor (layer0_outputs(2742));
    layer1_outputs(5464) <= (layer0_outputs(6113)) and not (layer0_outputs(3933));
    layer1_outputs(5465) <= not(layer0_outputs(5271));
    layer1_outputs(5466) <= layer0_outputs(6382);
    layer1_outputs(5467) <= not((layer0_outputs(478)) or (layer0_outputs(876)));
    layer1_outputs(5468) <= (layer0_outputs(923)) or (layer0_outputs(6275));
    layer1_outputs(5469) <= (layer0_outputs(7377)) and not (layer0_outputs(420));
    layer1_outputs(5470) <= layer0_outputs(2347);
    layer1_outputs(5471) <= not((layer0_outputs(7124)) or (layer0_outputs(4766)));
    layer1_outputs(5472) <= not(layer0_outputs(5240));
    layer1_outputs(5473) <= not((layer0_outputs(2294)) or (layer0_outputs(6180)));
    layer1_outputs(5474) <= (layer0_outputs(5367)) and not (layer0_outputs(359));
    layer1_outputs(5475) <= not(layer0_outputs(2066));
    layer1_outputs(5476) <= (layer0_outputs(1924)) and not (layer0_outputs(4527));
    layer1_outputs(5477) <= (layer0_outputs(7434)) xor (layer0_outputs(3176));
    layer1_outputs(5478) <= layer0_outputs(2990);
    layer1_outputs(5479) <= '1';
    layer1_outputs(5480) <= not((layer0_outputs(6239)) or (layer0_outputs(6834)));
    layer1_outputs(5481) <= not(layer0_outputs(2317));
    layer1_outputs(5482) <= (layer0_outputs(1263)) and not (layer0_outputs(1680));
    layer1_outputs(5483) <= layer0_outputs(7206);
    layer1_outputs(5484) <= '1';
    layer1_outputs(5485) <= layer0_outputs(5811);
    layer1_outputs(5486) <= not(layer0_outputs(4443));
    layer1_outputs(5487) <= not(layer0_outputs(7175)) or (layer0_outputs(3897));
    layer1_outputs(5488) <= '0';
    layer1_outputs(5489) <= (layer0_outputs(7271)) and (layer0_outputs(3308));
    layer1_outputs(5490) <= not(layer0_outputs(3102));
    layer1_outputs(5491) <= layer0_outputs(3422);
    layer1_outputs(5492) <= layer0_outputs(4356);
    layer1_outputs(5493) <= (layer0_outputs(2364)) and not (layer0_outputs(4385));
    layer1_outputs(5494) <= (layer0_outputs(460)) or (layer0_outputs(2091));
    layer1_outputs(5495) <= not((layer0_outputs(5442)) and (layer0_outputs(5382)));
    layer1_outputs(5496) <= not(layer0_outputs(398)) or (layer0_outputs(4054));
    layer1_outputs(5497) <= (layer0_outputs(641)) and not (layer0_outputs(5903));
    layer1_outputs(5498) <= not(layer0_outputs(2383)) or (layer0_outputs(1432));
    layer1_outputs(5499) <= not(layer0_outputs(7515));
    layer1_outputs(5500) <= '1';
    layer1_outputs(5501) <= (layer0_outputs(6526)) and not (layer0_outputs(2249));
    layer1_outputs(5502) <= not(layer0_outputs(6761)) or (layer0_outputs(3917));
    layer1_outputs(5503) <= '0';
    layer1_outputs(5504) <= '0';
    layer1_outputs(5505) <= '1';
    layer1_outputs(5506) <= (layer0_outputs(5428)) and not (layer0_outputs(2565));
    layer1_outputs(5507) <= '1';
    layer1_outputs(5508) <= layer0_outputs(3446);
    layer1_outputs(5509) <= not(layer0_outputs(3211)) or (layer0_outputs(2559));
    layer1_outputs(5510) <= (layer0_outputs(6719)) and (layer0_outputs(4374));
    layer1_outputs(5511) <= not((layer0_outputs(5637)) xor (layer0_outputs(3524)));
    layer1_outputs(5512) <= (layer0_outputs(5544)) and (layer0_outputs(7107));
    layer1_outputs(5513) <= not((layer0_outputs(3782)) or (layer0_outputs(7147)));
    layer1_outputs(5514) <= layer0_outputs(6243);
    layer1_outputs(5515) <= layer0_outputs(1400);
    layer1_outputs(5516) <= '1';
    layer1_outputs(5517) <= not(layer0_outputs(633));
    layer1_outputs(5518) <= not(layer0_outputs(5243)) or (layer0_outputs(1336));
    layer1_outputs(5519) <= not((layer0_outputs(24)) or (layer0_outputs(5147)));
    layer1_outputs(5520) <= (layer0_outputs(6885)) and not (layer0_outputs(4584));
    layer1_outputs(5521) <= not(layer0_outputs(4665));
    layer1_outputs(5522) <= '1';
    layer1_outputs(5523) <= not(layer0_outputs(199));
    layer1_outputs(5524) <= (layer0_outputs(794)) and (layer0_outputs(1730));
    layer1_outputs(5525) <= not(layer0_outputs(6139));
    layer1_outputs(5526) <= (layer0_outputs(7356)) and not (layer0_outputs(6341));
    layer1_outputs(5527) <= layer0_outputs(992);
    layer1_outputs(5528) <= not(layer0_outputs(6927)) or (layer0_outputs(758));
    layer1_outputs(5529) <= not(layer0_outputs(4698));
    layer1_outputs(5530) <= not((layer0_outputs(432)) xor (layer0_outputs(189)));
    layer1_outputs(5531) <= not((layer0_outputs(7476)) and (layer0_outputs(963)));
    layer1_outputs(5532) <= (layer0_outputs(5839)) and (layer0_outputs(5296));
    layer1_outputs(5533) <= (layer0_outputs(4615)) or (layer0_outputs(4767));
    layer1_outputs(5534) <= '1';
    layer1_outputs(5535) <= not(layer0_outputs(5533));
    layer1_outputs(5536) <= layer0_outputs(2618);
    layer1_outputs(5537) <= layer0_outputs(2107);
    layer1_outputs(5538) <= not(layer0_outputs(3542));
    layer1_outputs(5539) <= '1';
    layer1_outputs(5540) <= layer0_outputs(5170);
    layer1_outputs(5541) <= layer0_outputs(3422);
    layer1_outputs(5542) <= layer0_outputs(5770);
    layer1_outputs(5543) <= not((layer0_outputs(6482)) and (layer0_outputs(2013)));
    layer1_outputs(5544) <= (layer0_outputs(5003)) and not (layer0_outputs(7095));
    layer1_outputs(5545) <= not(layer0_outputs(7530)) or (layer0_outputs(4289));
    layer1_outputs(5546) <= (layer0_outputs(7488)) and not (layer0_outputs(3762));
    layer1_outputs(5547) <= (layer0_outputs(2031)) xor (layer0_outputs(6160));
    layer1_outputs(5548) <= (layer0_outputs(2355)) or (layer0_outputs(2229));
    layer1_outputs(5549) <= not(layer0_outputs(866));
    layer1_outputs(5550) <= not(layer0_outputs(4288));
    layer1_outputs(5551) <= not(layer0_outputs(1086)) or (layer0_outputs(7271));
    layer1_outputs(5552) <= not((layer0_outputs(6814)) and (layer0_outputs(117)));
    layer1_outputs(5553) <= not((layer0_outputs(2930)) xor (layer0_outputs(2548)));
    layer1_outputs(5554) <= layer0_outputs(5407);
    layer1_outputs(5555) <= (layer0_outputs(5168)) and (layer0_outputs(1227));
    layer1_outputs(5556) <= layer0_outputs(6739);
    layer1_outputs(5557) <= not(layer0_outputs(2431));
    layer1_outputs(5558) <= not(layer0_outputs(2283)) or (layer0_outputs(3846));
    layer1_outputs(5559) <= not((layer0_outputs(4525)) or (layer0_outputs(982)));
    layer1_outputs(5560) <= not(layer0_outputs(4878)) or (layer0_outputs(578));
    layer1_outputs(5561) <= not(layer0_outputs(4260));
    layer1_outputs(5562) <= not(layer0_outputs(3625));
    layer1_outputs(5563) <= not(layer0_outputs(4219)) or (layer0_outputs(7456));
    layer1_outputs(5564) <= not(layer0_outputs(5851)) or (layer0_outputs(514));
    layer1_outputs(5565) <= '1';
    layer1_outputs(5566) <= (layer0_outputs(5808)) and (layer0_outputs(4609));
    layer1_outputs(5567) <= not(layer0_outputs(4699)) or (layer0_outputs(5762));
    layer1_outputs(5568) <= (layer0_outputs(438)) and not (layer0_outputs(5212));
    layer1_outputs(5569) <= layer0_outputs(7506);
    layer1_outputs(5570) <= (layer0_outputs(6331)) and not (layer0_outputs(5887));
    layer1_outputs(5571) <= (layer0_outputs(2702)) and not (layer0_outputs(1517));
    layer1_outputs(5572) <= '1';
    layer1_outputs(5573) <= (layer0_outputs(2850)) and not (layer0_outputs(6595));
    layer1_outputs(5574) <= layer0_outputs(6775);
    layer1_outputs(5575) <= not(layer0_outputs(1170)) or (layer0_outputs(5215));
    layer1_outputs(5576) <= not(layer0_outputs(582));
    layer1_outputs(5577) <= not(layer0_outputs(3720)) or (layer0_outputs(1798));
    layer1_outputs(5578) <= '0';
    layer1_outputs(5579) <= not(layer0_outputs(4916)) or (layer0_outputs(756));
    layer1_outputs(5580) <= not((layer0_outputs(4211)) or (layer0_outputs(4149)));
    layer1_outputs(5581) <= (layer0_outputs(4522)) and (layer0_outputs(4065));
    layer1_outputs(5582) <= not((layer0_outputs(5535)) and (layer0_outputs(4862)));
    layer1_outputs(5583) <= '0';
    layer1_outputs(5584) <= not(layer0_outputs(4764)) or (layer0_outputs(2296));
    layer1_outputs(5585) <= not(layer0_outputs(6769));
    layer1_outputs(5586) <= not(layer0_outputs(1822));
    layer1_outputs(5587) <= '0';
    layer1_outputs(5588) <= layer0_outputs(5642);
    layer1_outputs(5589) <= (layer0_outputs(630)) or (layer0_outputs(1946));
    layer1_outputs(5590) <= (layer0_outputs(510)) and not (layer0_outputs(7663));
    layer1_outputs(5591) <= not(layer0_outputs(1438));
    layer1_outputs(5592) <= not((layer0_outputs(6599)) or (layer0_outputs(5206)));
    layer1_outputs(5593) <= not(layer0_outputs(160));
    layer1_outputs(5594) <= '0';
    layer1_outputs(5595) <= not(layer0_outputs(4612));
    layer1_outputs(5596) <= (layer0_outputs(1371)) or (layer0_outputs(1055));
    layer1_outputs(5597) <= not(layer0_outputs(5819));
    layer1_outputs(5598) <= (layer0_outputs(5014)) and not (layer0_outputs(6502));
    layer1_outputs(5599) <= not(layer0_outputs(6404));
    layer1_outputs(5600) <= '1';
    layer1_outputs(5601) <= (layer0_outputs(3686)) or (layer0_outputs(3218));
    layer1_outputs(5602) <= not((layer0_outputs(7518)) xor (layer0_outputs(2459)));
    layer1_outputs(5603) <= not(layer0_outputs(797)) or (layer0_outputs(3608));
    layer1_outputs(5604) <= '0';
    layer1_outputs(5605) <= '1';
    layer1_outputs(5606) <= (layer0_outputs(5136)) and (layer0_outputs(2900));
    layer1_outputs(5607) <= not(layer0_outputs(3050)) or (layer0_outputs(575));
    layer1_outputs(5608) <= (layer0_outputs(2281)) and not (layer0_outputs(1856));
    layer1_outputs(5609) <= '0';
    layer1_outputs(5610) <= layer0_outputs(187);
    layer1_outputs(5611) <= not(layer0_outputs(6856)) or (layer0_outputs(943));
    layer1_outputs(5612) <= (layer0_outputs(1839)) or (layer0_outputs(6961));
    layer1_outputs(5613) <= layer0_outputs(7269);
    layer1_outputs(5614) <= layer0_outputs(7317);
    layer1_outputs(5615) <= layer0_outputs(6200);
    layer1_outputs(5616) <= not(layer0_outputs(1781));
    layer1_outputs(5617) <= (layer0_outputs(573)) and not (layer0_outputs(5968));
    layer1_outputs(5618) <= (layer0_outputs(5112)) or (layer0_outputs(7399));
    layer1_outputs(5619) <= '1';
    layer1_outputs(5620) <= not(layer0_outputs(6452));
    layer1_outputs(5621) <= layer0_outputs(2954);
    layer1_outputs(5622) <= '0';
    layer1_outputs(5623) <= (layer0_outputs(684)) or (layer0_outputs(5688));
    layer1_outputs(5624) <= not(layer0_outputs(2162)) or (layer0_outputs(973));
    layer1_outputs(5625) <= not(layer0_outputs(5532)) or (layer0_outputs(1480));
    layer1_outputs(5626) <= (layer0_outputs(2476)) and not (layer0_outputs(843));
    layer1_outputs(5627) <= not(layer0_outputs(2078)) or (layer0_outputs(3684));
    layer1_outputs(5628) <= not(layer0_outputs(2663)) or (layer0_outputs(5148));
    layer1_outputs(5629) <= not((layer0_outputs(3410)) or (layer0_outputs(2638)));
    layer1_outputs(5630) <= not(layer0_outputs(5694));
    layer1_outputs(5631) <= not((layer0_outputs(2705)) or (layer0_outputs(6514)));
    layer1_outputs(5632) <= layer0_outputs(6369);
    layer1_outputs(5633) <= (layer0_outputs(5307)) or (layer0_outputs(4627));
    layer1_outputs(5634) <= not(layer0_outputs(6153));
    layer1_outputs(5635) <= '0';
    layer1_outputs(5636) <= '0';
    layer1_outputs(5637) <= not(layer0_outputs(155));
    layer1_outputs(5638) <= '1';
    layer1_outputs(5639) <= not((layer0_outputs(6990)) or (layer0_outputs(4304)));
    layer1_outputs(5640) <= (layer0_outputs(5464)) and (layer0_outputs(5624));
    layer1_outputs(5641) <= (layer0_outputs(724)) and not (layer0_outputs(4106));
    layer1_outputs(5642) <= (layer0_outputs(6525)) and not (layer0_outputs(242));
    layer1_outputs(5643) <= not((layer0_outputs(6806)) and (layer0_outputs(1399)));
    layer1_outputs(5644) <= not(layer0_outputs(3034));
    layer1_outputs(5645) <= not((layer0_outputs(5466)) or (layer0_outputs(1818)));
    layer1_outputs(5646) <= not((layer0_outputs(5864)) and (layer0_outputs(4469)));
    layer1_outputs(5647) <= (layer0_outputs(6407)) and not (layer0_outputs(5104));
    layer1_outputs(5648) <= layer0_outputs(4351);
    layer1_outputs(5649) <= not(layer0_outputs(5959)) or (layer0_outputs(3585));
    layer1_outputs(5650) <= not(layer0_outputs(4337)) or (layer0_outputs(2044));
    layer1_outputs(5651) <= (layer0_outputs(6209)) and (layer0_outputs(452));
    layer1_outputs(5652) <= not((layer0_outputs(3898)) or (layer0_outputs(5724)));
    layer1_outputs(5653) <= not(layer0_outputs(650)) or (layer0_outputs(4827));
    layer1_outputs(5654) <= not(layer0_outputs(2339)) or (layer0_outputs(6415));
    layer1_outputs(5655) <= layer0_outputs(5466);
    layer1_outputs(5656) <= '1';
    layer1_outputs(5657) <= (layer0_outputs(2409)) and not (layer0_outputs(2619));
    layer1_outputs(5658) <= not(layer0_outputs(2978)) or (layer0_outputs(3563));
    layer1_outputs(5659) <= layer0_outputs(3984);
    layer1_outputs(5660) <= '1';
    layer1_outputs(5661) <= layer0_outputs(4222);
    layer1_outputs(5662) <= not(layer0_outputs(2707));
    layer1_outputs(5663) <= (layer0_outputs(819)) xor (layer0_outputs(5053));
    layer1_outputs(5664) <= not(layer0_outputs(2878)) or (layer0_outputs(1182));
    layer1_outputs(5665) <= '1';
    layer1_outputs(5666) <= '1';
    layer1_outputs(5667) <= layer0_outputs(1700);
    layer1_outputs(5668) <= (layer0_outputs(1558)) and not (layer0_outputs(1316));
    layer1_outputs(5669) <= '0';
    layer1_outputs(5670) <= not(layer0_outputs(4326));
    layer1_outputs(5671) <= layer0_outputs(6449);
    layer1_outputs(5672) <= not(layer0_outputs(6621));
    layer1_outputs(5673) <= '1';
    layer1_outputs(5674) <= not(layer0_outputs(3478));
    layer1_outputs(5675) <= not(layer0_outputs(2551));
    layer1_outputs(5676) <= layer0_outputs(4977);
    layer1_outputs(5677) <= not(layer0_outputs(2158)) or (layer0_outputs(2318));
    layer1_outputs(5678) <= (layer0_outputs(311)) and not (layer0_outputs(2362));
    layer1_outputs(5679) <= (layer0_outputs(5504)) and not (layer0_outputs(4564));
    layer1_outputs(5680) <= not(layer0_outputs(6187)) or (layer0_outputs(223));
    layer1_outputs(5681) <= (layer0_outputs(4883)) and not (layer0_outputs(2352));
    layer1_outputs(5682) <= layer0_outputs(2490);
    layer1_outputs(5683) <= not(layer0_outputs(913));
    layer1_outputs(5684) <= '1';
    layer1_outputs(5685) <= '0';
    layer1_outputs(5686) <= not(layer0_outputs(5950));
    layer1_outputs(5687) <= layer0_outputs(3199);
    layer1_outputs(5688) <= '0';
    layer1_outputs(5689) <= (layer0_outputs(1297)) and not (layer0_outputs(1982));
    layer1_outputs(5690) <= (layer0_outputs(884)) and not (layer0_outputs(4674));
    layer1_outputs(5691) <= layer0_outputs(2916);
    layer1_outputs(5692) <= not(layer0_outputs(1978)) or (layer0_outputs(6535));
    layer1_outputs(5693) <= (layer0_outputs(1830)) and not (layer0_outputs(1965));
    layer1_outputs(5694) <= '1';
    layer1_outputs(5695) <= (layer0_outputs(1678)) and (layer0_outputs(2901));
    layer1_outputs(5696) <= not(layer0_outputs(645)) or (layer0_outputs(1891));
    layer1_outputs(5697) <= layer0_outputs(7482);
    layer1_outputs(5698) <= '0';
    layer1_outputs(5699) <= not(layer0_outputs(4307)) or (layer0_outputs(6674));
    layer1_outputs(5700) <= (layer0_outputs(7610)) and not (layer0_outputs(6425));
    layer1_outputs(5701) <= not(layer0_outputs(2601));
    layer1_outputs(5702) <= (layer0_outputs(4077)) xor (layer0_outputs(377));
    layer1_outputs(5703) <= not(layer0_outputs(818));
    layer1_outputs(5704) <= '0';
    layer1_outputs(5705) <= '0';
    layer1_outputs(5706) <= layer0_outputs(5404);
    layer1_outputs(5707) <= (layer0_outputs(7657)) and not (layer0_outputs(3492));
    layer1_outputs(5708) <= '0';
    layer1_outputs(5709) <= (layer0_outputs(5079)) and not (layer0_outputs(7535));
    layer1_outputs(5710) <= (layer0_outputs(5697)) and not (layer0_outputs(6486));
    layer1_outputs(5711) <= not(layer0_outputs(2017));
    layer1_outputs(5712) <= not(layer0_outputs(3349));
    layer1_outputs(5713) <= '1';
    layer1_outputs(5714) <= not((layer0_outputs(1316)) or (layer0_outputs(5345)));
    layer1_outputs(5715) <= (layer0_outputs(7026)) or (layer0_outputs(2145));
    layer1_outputs(5716) <= not(layer0_outputs(6807)) or (layer0_outputs(6790));
    layer1_outputs(5717) <= '1';
    layer1_outputs(5718) <= not((layer0_outputs(638)) xor (layer0_outputs(6460)));
    layer1_outputs(5719) <= (layer0_outputs(7651)) and (layer0_outputs(5559));
    layer1_outputs(5720) <= '1';
    layer1_outputs(5721) <= (layer0_outputs(1388)) and not (layer0_outputs(2757));
    layer1_outputs(5722) <= not(layer0_outputs(6284)) or (layer0_outputs(295));
    layer1_outputs(5723) <= layer0_outputs(7568);
    layer1_outputs(5724) <= (layer0_outputs(7382)) and not (layer0_outputs(3002));
    layer1_outputs(5725) <= '0';
    layer1_outputs(5726) <= (layer0_outputs(3144)) and not (layer0_outputs(5146));
    layer1_outputs(5727) <= layer0_outputs(5388);
    layer1_outputs(5728) <= (layer0_outputs(5797)) or (layer0_outputs(7309));
    layer1_outputs(5729) <= not((layer0_outputs(3827)) xor (layer0_outputs(6830)));
    layer1_outputs(5730) <= not(layer0_outputs(3345)) or (layer0_outputs(6135));
    layer1_outputs(5731) <= not(layer0_outputs(1528)) or (layer0_outputs(6199));
    layer1_outputs(5732) <= (layer0_outputs(6413)) and not (layer0_outputs(7155));
    layer1_outputs(5733) <= layer0_outputs(2431);
    layer1_outputs(5734) <= layer0_outputs(1880);
    layer1_outputs(5735) <= not(layer0_outputs(2803)) or (layer0_outputs(4209));
    layer1_outputs(5736) <= layer0_outputs(3730);
    layer1_outputs(5737) <= not(layer0_outputs(6279));
    layer1_outputs(5738) <= (layer0_outputs(2348)) and not (layer0_outputs(6748));
    layer1_outputs(5739) <= not((layer0_outputs(4398)) or (layer0_outputs(7054)));
    layer1_outputs(5740) <= layer0_outputs(5915);
    layer1_outputs(5741) <= layer0_outputs(5881);
    layer1_outputs(5742) <= not((layer0_outputs(2449)) or (layer0_outputs(5617)));
    layer1_outputs(5743) <= layer0_outputs(7395);
    layer1_outputs(5744) <= not(layer0_outputs(1960));
    layer1_outputs(5745) <= (layer0_outputs(6881)) and not (layer0_outputs(535));
    layer1_outputs(5746) <= not((layer0_outputs(4455)) or (layer0_outputs(3627)));
    layer1_outputs(5747) <= not(layer0_outputs(313));
    layer1_outputs(5748) <= (layer0_outputs(3742)) and (layer0_outputs(2256));
    layer1_outputs(5749) <= (layer0_outputs(7670)) or (layer0_outputs(174));
    layer1_outputs(5750) <= layer0_outputs(6769);
    layer1_outputs(5751) <= (layer0_outputs(44)) and (layer0_outputs(3238));
    layer1_outputs(5752) <= '0';
    layer1_outputs(5753) <= (layer0_outputs(2566)) or (layer0_outputs(938));
    layer1_outputs(5754) <= (layer0_outputs(3335)) and not (layer0_outputs(775));
    layer1_outputs(5755) <= layer0_outputs(7450);
    layer1_outputs(5756) <= '1';
    layer1_outputs(5757) <= '0';
    layer1_outputs(5758) <= (layer0_outputs(4987)) and not (layer0_outputs(2851));
    layer1_outputs(5759) <= '1';
    layer1_outputs(5760) <= (layer0_outputs(4611)) and (layer0_outputs(6234));
    layer1_outputs(5761) <= (layer0_outputs(6755)) or (layer0_outputs(5350));
    layer1_outputs(5762) <= layer0_outputs(6931);
    layer1_outputs(5763) <= not(layer0_outputs(7349));
    layer1_outputs(5764) <= '1';
    layer1_outputs(5765) <= (layer0_outputs(6495)) and not (layer0_outputs(6624));
    layer1_outputs(5766) <= (layer0_outputs(7178)) or (layer0_outputs(5633));
    layer1_outputs(5767) <= (layer0_outputs(310)) and not (layer0_outputs(6930));
    layer1_outputs(5768) <= '0';
    layer1_outputs(5769) <= '0';
    layer1_outputs(5770) <= layer0_outputs(7166);
    layer1_outputs(5771) <= not(layer0_outputs(6627)) or (layer0_outputs(3425));
    layer1_outputs(5772) <= not(layer0_outputs(4999)) or (layer0_outputs(5489));
    layer1_outputs(5773) <= layer0_outputs(7284);
    layer1_outputs(5774) <= (layer0_outputs(5050)) or (layer0_outputs(2087));
    layer1_outputs(5775) <= not(layer0_outputs(6609)) or (layer0_outputs(3560));
    layer1_outputs(5776) <= layer0_outputs(1486);
    layer1_outputs(5777) <= not(layer0_outputs(3111));
    layer1_outputs(5778) <= (layer0_outputs(4008)) and (layer0_outputs(6255));
    layer1_outputs(5779) <= not(layer0_outputs(4607)) or (layer0_outputs(129));
    layer1_outputs(5780) <= (layer0_outputs(2534)) and not (layer0_outputs(5921));
    layer1_outputs(5781) <= '1';
    layer1_outputs(5782) <= '0';
    layer1_outputs(5783) <= not((layer0_outputs(3878)) and (layer0_outputs(7393)));
    layer1_outputs(5784) <= not((layer0_outputs(3799)) or (layer0_outputs(383)));
    layer1_outputs(5785) <= not(layer0_outputs(5002)) or (layer0_outputs(2447));
    layer1_outputs(5786) <= layer0_outputs(6547);
    layer1_outputs(5787) <= '0';
    layer1_outputs(5788) <= layer0_outputs(453);
    layer1_outputs(5789) <= not((layer0_outputs(2599)) or (layer0_outputs(2284)));
    layer1_outputs(5790) <= layer0_outputs(5087);
    layer1_outputs(5791) <= (layer0_outputs(6102)) and not (layer0_outputs(6328));
    layer1_outputs(5792) <= layer0_outputs(160);
    layer1_outputs(5793) <= (layer0_outputs(2326)) and not (layer0_outputs(5106));
    layer1_outputs(5794) <= '0';
    layer1_outputs(5795) <= not((layer0_outputs(6062)) and (layer0_outputs(3374)));
    layer1_outputs(5796) <= layer0_outputs(5904);
    layer1_outputs(5797) <= (layer0_outputs(686)) or (layer0_outputs(4565));
    layer1_outputs(5798) <= not((layer0_outputs(4042)) and (layer0_outputs(4394)));
    layer1_outputs(5799) <= not((layer0_outputs(2729)) or (layer0_outputs(401)));
    layer1_outputs(5800) <= not((layer0_outputs(3700)) or (layer0_outputs(231)));
    layer1_outputs(5801) <= not((layer0_outputs(4723)) xor (layer0_outputs(6172)));
    layer1_outputs(5802) <= not(layer0_outputs(6490)) or (layer0_outputs(1711));
    layer1_outputs(5803) <= not(layer0_outputs(4085));
    layer1_outputs(5804) <= not((layer0_outputs(1073)) or (layer0_outputs(1867)));
    layer1_outputs(5805) <= not(layer0_outputs(4093)) or (layer0_outputs(1658));
    layer1_outputs(5806) <= '0';
    layer1_outputs(5807) <= not((layer0_outputs(334)) or (layer0_outputs(6054)));
    layer1_outputs(5808) <= layer0_outputs(5508);
    layer1_outputs(5809) <= '1';
    layer1_outputs(5810) <= not(layer0_outputs(7012)) or (layer0_outputs(5285));
    layer1_outputs(5811) <= not(layer0_outputs(4221)) or (layer0_outputs(7664));
    layer1_outputs(5812) <= not((layer0_outputs(5125)) and (layer0_outputs(4860)));
    layer1_outputs(5813) <= not((layer0_outputs(644)) or (layer0_outputs(429)));
    layer1_outputs(5814) <= (layer0_outputs(7190)) and not (layer0_outputs(5650));
    layer1_outputs(5815) <= '1';
    layer1_outputs(5816) <= not(layer0_outputs(6302)) or (layer0_outputs(4488));
    layer1_outputs(5817) <= not(layer0_outputs(2040));
    layer1_outputs(5818) <= (layer0_outputs(5213)) and not (layer0_outputs(4935));
    layer1_outputs(5819) <= not(layer0_outputs(928));
    layer1_outputs(5820) <= layer0_outputs(4272);
    layer1_outputs(5821) <= not(layer0_outputs(3954));
    layer1_outputs(5822) <= layer0_outputs(940);
    layer1_outputs(5823) <= '0';
    layer1_outputs(5824) <= not(layer0_outputs(6118));
    layer1_outputs(5825) <= '1';
    layer1_outputs(5826) <= (layer0_outputs(3347)) or (layer0_outputs(3935));
    layer1_outputs(5827) <= (layer0_outputs(2415)) or (layer0_outputs(4746));
    layer1_outputs(5828) <= '1';
    layer1_outputs(5829) <= layer0_outputs(2926);
    layer1_outputs(5830) <= layer0_outputs(6715);
    layer1_outputs(5831) <= not((layer0_outputs(4700)) or (layer0_outputs(2986)));
    layer1_outputs(5832) <= '0';
    layer1_outputs(5833) <= '0';
    layer1_outputs(5834) <= layer0_outputs(4748);
    layer1_outputs(5835) <= '0';
    layer1_outputs(5836) <= not((layer0_outputs(1792)) and (layer0_outputs(2298)));
    layer1_outputs(5837) <= '1';
    layer1_outputs(5838) <= layer0_outputs(2033);
    layer1_outputs(5839) <= layer0_outputs(3276);
    layer1_outputs(5840) <= not((layer0_outputs(5828)) and (layer0_outputs(2181)));
    layer1_outputs(5841) <= not((layer0_outputs(3056)) and (layer0_outputs(5938)));
    layer1_outputs(5842) <= not((layer0_outputs(6366)) xor (layer0_outputs(473)));
    layer1_outputs(5843) <= not(layer0_outputs(965)) or (layer0_outputs(2395));
    layer1_outputs(5844) <= layer0_outputs(768);
    layer1_outputs(5845) <= not((layer0_outputs(5843)) or (layer0_outputs(2674)));
    layer1_outputs(5846) <= '1';
    layer1_outputs(5847) <= (layer0_outputs(5847)) and not (layer0_outputs(1202));
    layer1_outputs(5848) <= not((layer0_outputs(2970)) or (layer0_outputs(3271)));
    layer1_outputs(5849) <= (layer0_outputs(1148)) and not (layer0_outputs(3201));
    layer1_outputs(5850) <= (layer0_outputs(5181)) and not (layer0_outputs(4116));
    layer1_outputs(5851) <= not(layer0_outputs(3894));
    layer1_outputs(5852) <= '0';
    layer1_outputs(5853) <= '1';
    layer1_outputs(5854) <= not(layer0_outputs(7644));
    layer1_outputs(5855) <= (layer0_outputs(3363)) and (layer0_outputs(598));
    layer1_outputs(5856) <= not(layer0_outputs(1053));
    layer1_outputs(5857) <= '1';
    layer1_outputs(5858) <= (layer0_outputs(598)) and not (layer0_outputs(6462));
    layer1_outputs(5859) <= '1';
    layer1_outputs(5860) <= (layer0_outputs(7364)) and (layer0_outputs(6176));
    layer1_outputs(5861) <= layer0_outputs(919);
    layer1_outputs(5862) <= layer0_outputs(558);
    layer1_outputs(5863) <= '0';
    layer1_outputs(5864) <= (layer0_outputs(4971)) and (layer0_outputs(7405));
    layer1_outputs(5865) <= layer0_outputs(5268);
    layer1_outputs(5866) <= '1';
    layer1_outputs(5867) <= not(layer0_outputs(6067));
    layer1_outputs(5868) <= layer0_outputs(5933);
    layer1_outputs(5869) <= not(layer0_outputs(1724)) or (layer0_outputs(6473));
    layer1_outputs(5870) <= not(layer0_outputs(1950));
    layer1_outputs(5871) <= not(layer0_outputs(7041));
    layer1_outputs(5872) <= not((layer0_outputs(4493)) or (layer0_outputs(5352)));
    layer1_outputs(5873) <= '0';
    layer1_outputs(5874) <= (layer0_outputs(6914)) and not (layer0_outputs(7347));
    layer1_outputs(5875) <= layer0_outputs(17);
    layer1_outputs(5876) <= layer0_outputs(7632);
    layer1_outputs(5877) <= not((layer0_outputs(822)) xor (layer0_outputs(3041)));
    layer1_outputs(5878) <= '1';
    layer1_outputs(5879) <= not((layer0_outputs(7353)) or (layer0_outputs(2533)));
    layer1_outputs(5880) <= not(layer0_outputs(799)) or (layer0_outputs(1291));
    layer1_outputs(5881) <= (layer0_outputs(2983)) and (layer0_outputs(3720));
    layer1_outputs(5882) <= (layer0_outputs(6855)) and not (layer0_outputs(496));
    layer1_outputs(5883) <= '0';
    layer1_outputs(5884) <= not((layer0_outputs(3115)) or (layer0_outputs(2014)));
    layer1_outputs(5885) <= not(layer0_outputs(4946)) or (layer0_outputs(4952));
    layer1_outputs(5886) <= (layer0_outputs(2623)) and not (layer0_outputs(6673));
    layer1_outputs(5887) <= (layer0_outputs(6949)) or (layer0_outputs(7580));
    layer1_outputs(5888) <= layer0_outputs(5659);
    layer1_outputs(5889) <= (layer0_outputs(6870)) xor (layer0_outputs(1559));
    layer1_outputs(5890) <= (layer0_outputs(6767)) and not (layer0_outputs(5923));
    layer1_outputs(5891) <= '1';
    layer1_outputs(5892) <= (layer0_outputs(3378)) or (layer0_outputs(5622));
    layer1_outputs(5893) <= (layer0_outputs(1912)) and (layer0_outputs(1572));
    layer1_outputs(5894) <= '1';
    layer1_outputs(5895) <= '1';
    layer1_outputs(5896) <= not(layer0_outputs(2356)) or (layer0_outputs(4149));
    layer1_outputs(5897) <= not(layer0_outputs(4112));
    layer1_outputs(5898) <= not(layer0_outputs(4460));
    layer1_outputs(5899) <= '1';
    layer1_outputs(5900) <= not((layer0_outputs(87)) or (layer0_outputs(4072)));
    layer1_outputs(5901) <= not((layer0_outputs(3953)) or (layer0_outputs(2252)));
    layer1_outputs(5902) <= not(layer0_outputs(2513)) or (layer0_outputs(1370));
    layer1_outputs(5903) <= (layer0_outputs(7397)) and not (layer0_outputs(5267));
    layer1_outputs(5904) <= layer0_outputs(529);
    layer1_outputs(5905) <= '0';
    layer1_outputs(5906) <= not((layer0_outputs(7377)) and (layer0_outputs(7053)));
    layer1_outputs(5907) <= (layer0_outputs(6780)) and not (layer0_outputs(1608));
    layer1_outputs(5908) <= not(layer0_outputs(3606)) or (layer0_outputs(6401));
    layer1_outputs(5909) <= (layer0_outputs(1403)) and not (layer0_outputs(612));
    layer1_outputs(5910) <= (layer0_outputs(4638)) and (layer0_outputs(6735));
    layer1_outputs(5911) <= layer0_outputs(5021);
    layer1_outputs(5912) <= not(layer0_outputs(7341));
    layer1_outputs(5913) <= (layer0_outputs(1663)) and (layer0_outputs(594));
    layer1_outputs(5914) <= not(layer0_outputs(7441));
    layer1_outputs(5915) <= not((layer0_outputs(7189)) or (layer0_outputs(752)));
    layer1_outputs(5916) <= not(layer0_outputs(5372));
    layer1_outputs(5917) <= '1';
    layer1_outputs(5918) <= not(layer0_outputs(261)) or (layer0_outputs(2147));
    layer1_outputs(5919) <= '1';
    layer1_outputs(5920) <= (layer0_outputs(4523)) xor (layer0_outputs(5306));
    layer1_outputs(5921) <= not((layer0_outputs(4109)) or (layer0_outputs(2770)));
    layer1_outputs(5922) <= '0';
    layer1_outputs(5923) <= (layer0_outputs(2170)) and not (layer0_outputs(1460));
    layer1_outputs(5924) <= '1';
    layer1_outputs(5925) <= not(layer0_outputs(1621));
    layer1_outputs(5926) <= not(layer0_outputs(1912));
    layer1_outputs(5927) <= (layer0_outputs(2252)) and not (layer0_outputs(5726));
    layer1_outputs(5928) <= (layer0_outputs(4350)) and not (layer0_outputs(534));
    layer1_outputs(5929) <= not(layer0_outputs(3286)) or (layer0_outputs(7468));
    layer1_outputs(5930) <= not((layer0_outputs(5113)) and (layer0_outputs(725)));
    layer1_outputs(5931) <= (layer0_outputs(2889)) or (layer0_outputs(1640));
    layer1_outputs(5932) <= not(layer0_outputs(7574));
    layer1_outputs(5933) <= '0';
    layer1_outputs(5934) <= '1';
    layer1_outputs(5935) <= not(layer0_outputs(4414));
    layer1_outputs(5936) <= (layer0_outputs(2180)) and not (layer0_outputs(7520));
    layer1_outputs(5937) <= (layer0_outputs(971)) and not (layer0_outputs(6569));
    layer1_outputs(5938) <= '1';
    layer1_outputs(5939) <= layer0_outputs(4621);
    layer1_outputs(5940) <= not((layer0_outputs(2860)) and (layer0_outputs(1836)));
    layer1_outputs(5941) <= not((layer0_outputs(236)) and (layer0_outputs(4319)));
    layer1_outputs(5942) <= not(layer0_outputs(1634)) or (layer0_outputs(6021));
    layer1_outputs(5943) <= layer0_outputs(7202);
    layer1_outputs(5944) <= (layer0_outputs(6709)) and not (layer0_outputs(7274));
    layer1_outputs(5945) <= (layer0_outputs(6280)) or (layer0_outputs(6890));
    layer1_outputs(5946) <= layer0_outputs(6408);
    layer1_outputs(5947) <= not((layer0_outputs(3621)) or (layer0_outputs(680)));
    layer1_outputs(5948) <= '1';
    layer1_outputs(5949) <= not(layer0_outputs(6574));
    layer1_outputs(5950) <= not(layer0_outputs(7398));
    layer1_outputs(5951) <= not((layer0_outputs(1884)) or (layer0_outputs(5346)));
    layer1_outputs(5952) <= (layer0_outputs(3512)) and (layer0_outputs(6320));
    layer1_outputs(5953) <= not(layer0_outputs(6904)) or (layer0_outputs(2361));
    layer1_outputs(5954) <= layer0_outputs(719);
    layer1_outputs(5955) <= (layer0_outputs(670)) and not (layer0_outputs(2444));
    layer1_outputs(5956) <= (layer0_outputs(2123)) and not (layer0_outputs(482));
    layer1_outputs(5957) <= (layer0_outputs(50)) and (layer0_outputs(3117));
    layer1_outputs(5958) <= '1';
    layer1_outputs(5959) <= layer0_outputs(3583);
    layer1_outputs(5960) <= not((layer0_outputs(2190)) and (layer0_outputs(2247)));
    layer1_outputs(5961) <= not(layer0_outputs(5841)) or (layer0_outputs(2657));
    layer1_outputs(5962) <= not(layer0_outputs(3759)) or (layer0_outputs(7658));
    layer1_outputs(5963) <= not(layer0_outputs(3)) or (layer0_outputs(4089));
    layer1_outputs(5964) <= not(layer0_outputs(636)) or (layer0_outputs(5092));
    layer1_outputs(5965) <= (layer0_outputs(7622)) or (layer0_outputs(2920));
    layer1_outputs(5966) <= not((layer0_outputs(3797)) or (layer0_outputs(776)));
    layer1_outputs(5967) <= not(layer0_outputs(5128)) or (layer0_outputs(2130));
    layer1_outputs(5968) <= (layer0_outputs(900)) and (layer0_outputs(490));
    layer1_outputs(5969) <= not(layer0_outputs(830));
    layer1_outputs(5970) <= not((layer0_outputs(5033)) and (layer0_outputs(3581)));
    layer1_outputs(5971) <= not(layer0_outputs(2361));
    layer1_outputs(5972) <= (layer0_outputs(2112)) or (layer0_outputs(3491));
    layer1_outputs(5973) <= layer0_outputs(2910);
    layer1_outputs(5974) <= (layer0_outputs(1411)) or (layer0_outputs(1036));
    layer1_outputs(5975) <= not((layer0_outputs(2515)) and (layer0_outputs(2681)));
    layer1_outputs(5976) <= not(layer0_outputs(1922));
    layer1_outputs(5977) <= (layer0_outputs(3303)) and (layer0_outputs(2057));
    layer1_outputs(5978) <= not(layer0_outputs(7573)) or (layer0_outputs(2610));
    layer1_outputs(5979) <= not(layer0_outputs(1788)) or (layer0_outputs(4851));
    layer1_outputs(5980) <= (layer0_outputs(6177)) and not (layer0_outputs(750));
    layer1_outputs(5981) <= (layer0_outputs(7266)) and not (layer0_outputs(1930));
    layer1_outputs(5982) <= layer0_outputs(4589);
    layer1_outputs(5983) <= (layer0_outputs(2367)) xor (layer0_outputs(1190));
    layer1_outputs(5984) <= '0';
    layer1_outputs(5985) <= not(layer0_outputs(4960));
    layer1_outputs(5986) <= layer0_outputs(6442);
    layer1_outputs(5987) <= '0';
    layer1_outputs(5988) <= layer0_outputs(728);
    layer1_outputs(5989) <= '1';
    layer1_outputs(5990) <= not(layer0_outputs(3781));
    layer1_outputs(5991) <= not((layer0_outputs(1080)) and (layer0_outputs(3291)));
    layer1_outputs(5992) <= layer0_outputs(4108);
    layer1_outputs(5993) <= not(layer0_outputs(1674));
    layer1_outputs(5994) <= layer0_outputs(5760);
    layer1_outputs(5995) <= layer0_outputs(295);
    layer1_outputs(5996) <= not((layer0_outputs(4237)) or (layer0_outputs(1570)));
    layer1_outputs(5997) <= '1';
    layer1_outputs(5998) <= layer0_outputs(3070);
    layer1_outputs(5999) <= not(layer0_outputs(6731));
    layer1_outputs(6000) <= not((layer0_outputs(1026)) and (layer0_outputs(4281)));
    layer1_outputs(6001) <= '1';
    layer1_outputs(6002) <= not(layer0_outputs(2538)) or (layer0_outputs(3738));
    layer1_outputs(6003) <= not((layer0_outputs(2321)) and (layer0_outputs(3375)));
    layer1_outputs(6004) <= '0';
    layer1_outputs(6005) <= (layer0_outputs(569)) and not (layer0_outputs(3018));
    layer1_outputs(6006) <= not(layer0_outputs(6288)) or (layer0_outputs(63));
    layer1_outputs(6007) <= not(layer0_outputs(4142)) or (layer0_outputs(1382));
    layer1_outputs(6008) <= not(layer0_outputs(4302));
    layer1_outputs(6009) <= (layer0_outputs(3356)) and not (layer0_outputs(5970));
    layer1_outputs(6010) <= '1';
    layer1_outputs(6011) <= not((layer0_outputs(2394)) and (layer0_outputs(5067)));
    layer1_outputs(6012) <= not(layer0_outputs(3477));
    layer1_outputs(6013) <= not(layer0_outputs(3593)) or (layer0_outputs(1344));
    layer1_outputs(6014) <= layer0_outputs(6135);
    layer1_outputs(6015) <= (layer0_outputs(5642)) and not (layer0_outputs(6624));
    layer1_outputs(6016) <= (layer0_outputs(7616)) and not (layer0_outputs(592));
    layer1_outputs(6017) <= (layer0_outputs(1877)) xor (layer0_outputs(4375));
    layer1_outputs(6018) <= (layer0_outputs(1588)) and not (layer0_outputs(5041));
    layer1_outputs(6019) <= (layer0_outputs(5556)) or (layer0_outputs(1299));
    layer1_outputs(6020) <= not((layer0_outputs(4100)) and (layer0_outputs(93)));
    layer1_outputs(6021) <= (layer0_outputs(1952)) and (layer0_outputs(6439));
    layer1_outputs(6022) <= (layer0_outputs(2807)) xor (layer0_outputs(2421));
    layer1_outputs(6023) <= '1';
    layer1_outputs(6024) <= layer0_outputs(4296);
    layer1_outputs(6025) <= not(layer0_outputs(2932));
    layer1_outputs(6026) <= not(layer0_outputs(1262));
    layer1_outputs(6027) <= not(layer0_outputs(1959)) or (layer0_outputs(5611));
    layer1_outputs(6028) <= '0';
    layer1_outputs(6029) <= (layer0_outputs(4695)) and not (layer0_outputs(5869));
    layer1_outputs(6030) <= not((layer0_outputs(1556)) or (layer0_outputs(7011)));
    layer1_outputs(6031) <= (layer0_outputs(3352)) and not (layer0_outputs(1221));
    layer1_outputs(6032) <= not((layer0_outputs(904)) or (layer0_outputs(6111)));
    layer1_outputs(6033) <= layer0_outputs(262);
    layer1_outputs(6034) <= '1';
    layer1_outputs(6035) <= '0';
    layer1_outputs(6036) <= layer0_outputs(7309);
    layer1_outputs(6037) <= (layer0_outputs(3584)) or (layer0_outputs(6506));
    layer1_outputs(6038) <= layer0_outputs(6780);
    layer1_outputs(6039) <= layer0_outputs(6273);
    layer1_outputs(6040) <= (layer0_outputs(5432)) xor (layer0_outputs(2043));
    layer1_outputs(6041) <= (layer0_outputs(3299)) and not (layer0_outputs(3812));
    layer1_outputs(6042) <= (layer0_outputs(5927)) and not (layer0_outputs(2720));
    layer1_outputs(6043) <= layer0_outputs(5824);
    layer1_outputs(6044) <= (layer0_outputs(4489)) and (layer0_outputs(6237));
    layer1_outputs(6045) <= (layer0_outputs(2269)) and not (layer0_outputs(3420));
    layer1_outputs(6046) <= not(layer0_outputs(999));
    layer1_outputs(6047) <= layer0_outputs(6703);
    layer1_outputs(6048) <= (layer0_outputs(554)) and (layer0_outputs(793));
    layer1_outputs(6049) <= layer0_outputs(151);
    layer1_outputs(6050) <= (layer0_outputs(2653)) and (layer0_outputs(1490));
    layer1_outputs(6051) <= not(layer0_outputs(1224)) or (layer0_outputs(7405));
    layer1_outputs(6052) <= (layer0_outputs(2029)) and not (layer0_outputs(3455));
    layer1_outputs(6053) <= '1';
    layer1_outputs(6054) <= not(layer0_outputs(5120));
    layer1_outputs(6055) <= not(layer0_outputs(7030));
    layer1_outputs(6056) <= layer0_outputs(6515);
    layer1_outputs(6057) <= not((layer0_outputs(5197)) and (layer0_outputs(7113)));
    layer1_outputs(6058) <= (layer0_outputs(5391)) or (layer0_outputs(3817));
    layer1_outputs(6059) <= layer0_outputs(205);
    layer1_outputs(6060) <= not(layer0_outputs(4621));
    layer1_outputs(6061) <= (layer0_outputs(1269)) and not (layer0_outputs(2677));
    layer1_outputs(6062) <= not((layer0_outputs(7455)) or (layer0_outputs(7219)));
    layer1_outputs(6063) <= '1';
    layer1_outputs(6064) <= '0';
    layer1_outputs(6065) <= (layer0_outputs(4131)) and (layer0_outputs(3525));
    layer1_outputs(6066) <= not(layer0_outputs(381));
    layer1_outputs(6067) <= (layer0_outputs(3700)) and not (layer0_outputs(7303));
    layer1_outputs(6068) <= not(layer0_outputs(4146));
    layer1_outputs(6069) <= not(layer0_outputs(5720)) or (layer0_outputs(2286));
    layer1_outputs(6070) <= '1';
    layer1_outputs(6071) <= layer0_outputs(2393);
    layer1_outputs(6072) <= (layer0_outputs(3052)) and (layer0_outputs(2871));
    layer1_outputs(6073) <= (layer0_outputs(4201)) and not (layer0_outputs(253));
    layer1_outputs(6074) <= not((layer0_outputs(897)) or (layer0_outputs(7203)));
    layer1_outputs(6075) <= layer0_outputs(7283);
    layer1_outputs(6076) <= '1';
    layer1_outputs(6077) <= not((layer0_outputs(3923)) or (layer0_outputs(800)));
    layer1_outputs(6078) <= '1';
    layer1_outputs(6079) <= not(layer0_outputs(4685));
    layer1_outputs(6080) <= not(layer0_outputs(2358)) or (layer0_outputs(2017));
    layer1_outputs(6081) <= '0';
    layer1_outputs(6082) <= '1';
    layer1_outputs(6083) <= '1';
    layer1_outputs(6084) <= not(layer0_outputs(2299));
    layer1_outputs(6085) <= layer0_outputs(5026);
    layer1_outputs(6086) <= not(layer0_outputs(4090)) or (layer0_outputs(5033));
    layer1_outputs(6087) <= '1';
    layer1_outputs(6088) <= (layer0_outputs(3148)) or (layer0_outputs(7055));
    layer1_outputs(6089) <= (layer0_outputs(6183)) and not (layer0_outputs(7390));
    layer1_outputs(6090) <= not(layer0_outputs(5275));
    layer1_outputs(6091) <= (layer0_outputs(5791)) and (layer0_outputs(5958));
    layer1_outputs(6092) <= not(layer0_outputs(2275)) or (layer0_outputs(7463));
    layer1_outputs(6093) <= layer0_outputs(3264);
    layer1_outputs(6094) <= (layer0_outputs(1593)) and not (layer0_outputs(5935));
    layer1_outputs(6095) <= (layer0_outputs(3478)) and not (layer0_outputs(7204));
    layer1_outputs(6096) <= not(layer0_outputs(7002));
    layer1_outputs(6097) <= not(layer0_outputs(5922));
    layer1_outputs(6098) <= '0';
    layer1_outputs(6099) <= not(layer0_outputs(3778));
    layer1_outputs(6100) <= layer0_outputs(6029);
    layer1_outputs(6101) <= not(layer0_outputs(3918));
    layer1_outputs(6102) <= '0';
    layer1_outputs(6103) <= '0';
    layer1_outputs(6104) <= not((layer0_outputs(3001)) or (layer0_outputs(2024)));
    layer1_outputs(6105) <= '0';
    layer1_outputs(6106) <= not(layer0_outputs(2232)) or (layer0_outputs(4327));
    layer1_outputs(6107) <= (layer0_outputs(3686)) and not (layer0_outputs(1099));
    layer1_outputs(6108) <= not(layer0_outputs(7236));
    layer1_outputs(6109) <= layer0_outputs(1570);
    layer1_outputs(6110) <= not(layer0_outputs(4868)) or (layer0_outputs(3655));
    layer1_outputs(6111) <= '1';
    layer1_outputs(6112) <= (layer0_outputs(3628)) or (layer0_outputs(1209));
    layer1_outputs(6113) <= not(layer0_outputs(1734)) or (layer0_outputs(7137));
    layer1_outputs(6114) <= not((layer0_outputs(2265)) or (layer0_outputs(1375)));
    layer1_outputs(6115) <= (layer0_outputs(3450)) xor (layer0_outputs(5360));
    layer1_outputs(6116) <= (layer0_outputs(3957)) and (layer0_outputs(660));
    layer1_outputs(6117) <= not((layer0_outputs(3028)) or (layer0_outputs(468)));
    layer1_outputs(6118) <= not(layer0_outputs(5723));
    layer1_outputs(6119) <= '0';
    layer1_outputs(6120) <= not((layer0_outputs(1988)) and (layer0_outputs(4673)));
    layer1_outputs(6121) <= layer0_outputs(5792);
    layer1_outputs(6122) <= layer0_outputs(1272);
    layer1_outputs(6123) <= not(layer0_outputs(5370));
    layer1_outputs(6124) <= not(layer0_outputs(5932));
    layer1_outputs(6125) <= (layer0_outputs(3455)) and not (layer0_outputs(403));
    layer1_outputs(6126) <= not((layer0_outputs(7432)) or (layer0_outputs(7307)));
    layer1_outputs(6127) <= layer0_outputs(5181);
    layer1_outputs(6128) <= layer0_outputs(2603);
    layer1_outputs(6129) <= '0';
    layer1_outputs(6130) <= '0';
    layer1_outputs(6131) <= not(layer0_outputs(993)) or (layer0_outputs(5875));
    layer1_outputs(6132) <= not(layer0_outputs(4362));
    layer1_outputs(6133) <= layer0_outputs(5507);
    layer1_outputs(6134) <= not((layer0_outputs(2666)) or (layer0_outputs(6653)));
    layer1_outputs(6135) <= (layer0_outputs(6316)) or (layer0_outputs(3062));
    layer1_outputs(6136) <= not(layer0_outputs(4805)) or (layer0_outputs(676));
    layer1_outputs(6137) <= not(layer0_outputs(6202));
    layer1_outputs(6138) <= not(layer0_outputs(2636)) or (layer0_outputs(3753));
    layer1_outputs(6139) <= not(layer0_outputs(3463));
    layer1_outputs(6140) <= not((layer0_outputs(6432)) or (layer0_outputs(2229)));
    layer1_outputs(6141) <= layer0_outputs(6248);
    layer1_outputs(6142) <= (layer0_outputs(934)) or (layer0_outputs(2755));
    layer1_outputs(6143) <= not(layer0_outputs(4370)) or (layer0_outputs(5803));
    layer1_outputs(6144) <= not((layer0_outputs(1052)) or (layer0_outputs(2480)));
    layer1_outputs(6145) <= not((layer0_outputs(2964)) xor (layer0_outputs(1527)));
    layer1_outputs(6146) <= '0';
    layer1_outputs(6147) <= not((layer0_outputs(6214)) or (layer0_outputs(736)));
    layer1_outputs(6148) <= (layer0_outputs(476)) and not (layer0_outputs(1434));
    layer1_outputs(6149) <= '0';
    layer1_outputs(6150) <= '0';
    layer1_outputs(6151) <= '1';
    layer1_outputs(6152) <= not(layer0_outputs(4297)) or (layer0_outputs(1318));
    layer1_outputs(6153) <= not((layer0_outputs(1377)) or (layer0_outputs(6138)));
    layer1_outputs(6154) <= (layer0_outputs(620)) or (layer0_outputs(3194));
    layer1_outputs(6155) <= layer0_outputs(626);
    layer1_outputs(6156) <= not(layer0_outputs(4273));
    layer1_outputs(6157) <= (layer0_outputs(2525)) or (layer0_outputs(5191));
    layer1_outputs(6158) <= not((layer0_outputs(7217)) or (layer0_outputs(5866)));
    layer1_outputs(6159) <= not(layer0_outputs(4926)) or (layer0_outputs(6117));
    layer1_outputs(6160) <= (layer0_outputs(7268)) and (layer0_outputs(4959));
    layer1_outputs(6161) <= not(layer0_outputs(1462)) or (layer0_outputs(5840));
    layer1_outputs(6162) <= not(layer0_outputs(2567)) or (layer0_outputs(65));
    layer1_outputs(6163) <= (layer0_outputs(5969)) or (layer0_outputs(2075));
    layer1_outputs(6164) <= not(layer0_outputs(3595)) or (layer0_outputs(3676));
    layer1_outputs(6165) <= (layer0_outputs(3480)) and not (layer0_outputs(346));
    layer1_outputs(6166) <= (layer0_outputs(7499)) and not (layer0_outputs(7503));
    layer1_outputs(6167) <= layer0_outputs(1590);
    layer1_outputs(6168) <= layer0_outputs(7065);
    layer1_outputs(6169) <= layer0_outputs(4729);
    layer1_outputs(6170) <= not((layer0_outputs(3924)) and (layer0_outputs(5364)));
    layer1_outputs(6171) <= not((layer0_outputs(1445)) xor (layer0_outputs(1126)));
    layer1_outputs(6172) <= (layer0_outputs(212)) xor (layer0_outputs(6474));
    layer1_outputs(6173) <= layer0_outputs(3350);
    layer1_outputs(6174) <= not((layer0_outputs(1484)) and (layer0_outputs(4845)));
    layer1_outputs(6175) <= (layer0_outputs(1597)) and not (layer0_outputs(1644));
    layer1_outputs(6176) <= (layer0_outputs(2835)) or (layer0_outputs(3836));
    layer1_outputs(6177) <= not(layer0_outputs(5021));
    layer1_outputs(6178) <= not(layer0_outputs(653));
    layer1_outputs(6179) <= (layer0_outputs(3841)) or (layer0_outputs(3290));
    layer1_outputs(6180) <= not((layer0_outputs(6368)) or (layer0_outputs(2261)));
    layer1_outputs(6181) <= not(layer0_outputs(5001)) or (layer0_outputs(4331));
    layer1_outputs(6182) <= layer0_outputs(6548);
    layer1_outputs(6183) <= not(layer0_outputs(3365));
    layer1_outputs(6184) <= (layer0_outputs(6238)) and (layer0_outputs(265));
    layer1_outputs(6185) <= '1';
    layer1_outputs(6186) <= (layer0_outputs(7589)) and (layer0_outputs(4471));
    layer1_outputs(6187) <= (layer0_outputs(5893)) or (layer0_outputs(2787));
    layer1_outputs(6188) <= '0';
    layer1_outputs(6189) <= (layer0_outputs(7612)) and not (layer0_outputs(3400));
    layer1_outputs(6190) <= not(layer0_outputs(2996)) or (layer0_outputs(2656));
    layer1_outputs(6191) <= (layer0_outputs(540)) and (layer0_outputs(3708));
    layer1_outputs(6192) <= not(layer0_outputs(1370));
    layer1_outputs(6193) <= not((layer0_outputs(86)) and (layer0_outputs(895)));
    layer1_outputs(6194) <= (layer0_outputs(1222)) and not (layer0_outputs(4098));
    layer1_outputs(6195) <= (layer0_outputs(2151)) and not (layer0_outputs(5415));
    layer1_outputs(6196) <= (layer0_outputs(6576)) and not (layer0_outputs(6822));
    layer1_outputs(6197) <= not((layer0_outputs(1878)) or (layer0_outputs(951)));
    layer1_outputs(6198) <= not((layer0_outputs(5861)) or (layer0_outputs(4354)));
    layer1_outputs(6199) <= not((layer0_outputs(1624)) or (layer0_outputs(1691)));
    layer1_outputs(6200) <= (layer0_outputs(4367)) or (layer0_outputs(829));
    layer1_outputs(6201) <= '1';
    layer1_outputs(6202) <= '0';
    layer1_outputs(6203) <= not(layer0_outputs(6725)) or (layer0_outputs(2563));
    layer1_outputs(6204) <= not((layer0_outputs(969)) and (layer0_outputs(1882)));
    layer1_outputs(6205) <= (layer0_outputs(1669)) and (layer0_outputs(4517));
    layer1_outputs(6206) <= not(layer0_outputs(1994));
    layer1_outputs(6207) <= '1';
    layer1_outputs(6208) <= (layer0_outputs(7045)) or (layer0_outputs(4530));
    layer1_outputs(6209) <= '0';
    layer1_outputs(6210) <= layer0_outputs(2868);
    layer1_outputs(6211) <= not(layer0_outputs(368)) or (layer0_outputs(5608));
    layer1_outputs(6212) <= not(layer0_outputs(7598)) or (layer0_outputs(3739));
    layer1_outputs(6213) <= layer0_outputs(7650);
    layer1_outputs(6214) <= not(layer0_outputs(3136));
    layer1_outputs(6215) <= '1';
    layer1_outputs(6216) <= (layer0_outputs(7218)) and not (layer0_outputs(3122));
    layer1_outputs(6217) <= '0';
    layer1_outputs(6218) <= not(layer0_outputs(3740));
    layer1_outputs(6219) <= layer0_outputs(3709);
    layer1_outputs(6220) <= layer0_outputs(1871);
    layer1_outputs(6221) <= '0';
    layer1_outputs(6222) <= '1';
    layer1_outputs(6223) <= not(layer0_outputs(5433)) or (layer0_outputs(6983));
    layer1_outputs(6224) <= not(layer0_outputs(3510));
    layer1_outputs(6225) <= not(layer0_outputs(6986)) or (layer0_outputs(4170));
    layer1_outputs(6226) <= not(layer0_outputs(1823)) or (layer0_outputs(4667));
    layer1_outputs(6227) <= not((layer0_outputs(4406)) and (layer0_outputs(3373)));
    layer1_outputs(6228) <= not((layer0_outputs(6358)) or (layer0_outputs(1973)));
    layer1_outputs(6229) <= not(layer0_outputs(3058));
    layer1_outputs(6230) <= (layer0_outputs(375)) and (layer0_outputs(2554));
    layer1_outputs(6231) <= layer0_outputs(632);
    layer1_outputs(6232) <= not(layer0_outputs(861));
    layer1_outputs(6233) <= (layer0_outputs(3000)) and not (layer0_outputs(6070));
    layer1_outputs(6234) <= not((layer0_outputs(2510)) or (layer0_outputs(5589)));
    layer1_outputs(6235) <= not((layer0_outputs(6962)) and (layer0_outputs(7418)));
    layer1_outputs(6236) <= not(layer0_outputs(2193));
    layer1_outputs(6237) <= (layer0_outputs(2315)) or (layer0_outputs(5945));
    layer1_outputs(6238) <= '1';
    layer1_outputs(6239) <= not((layer0_outputs(3272)) and (layer0_outputs(1017)));
    layer1_outputs(6240) <= layer0_outputs(4825);
    layer1_outputs(6241) <= not(layer0_outputs(2933));
    layer1_outputs(6242) <= not((layer0_outputs(2276)) or (layer0_outputs(2529)));
    layer1_outputs(6243) <= layer0_outputs(7082);
    layer1_outputs(6244) <= not((layer0_outputs(4834)) or (layer0_outputs(3456)));
    layer1_outputs(6245) <= '0';
    layer1_outputs(6246) <= layer0_outputs(3840);
    layer1_outputs(6247) <= (layer0_outputs(4542)) and not (layer0_outputs(4609));
    layer1_outputs(6248) <= '0';
    layer1_outputs(6249) <= not(layer0_outputs(351)) or (layer0_outputs(248));
    layer1_outputs(6250) <= (layer0_outputs(7427)) and (layer0_outputs(3653));
    layer1_outputs(6251) <= not(layer0_outputs(4628));
    layer1_outputs(6252) <= '0';
    layer1_outputs(6253) <= not((layer0_outputs(4205)) or (layer0_outputs(1993)));
    layer1_outputs(6254) <= layer0_outputs(1614);
    layer1_outputs(6255) <= (layer0_outputs(5579)) or (layer0_outputs(50));
    layer1_outputs(6256) <= '1';
    layer1_outputs(6257) <= layer0_outputs(2202);
    layer1_outputs(6258) <= not(layer0_outputs(6247));
    layer1_outputs(6259) <= '0';
    layer1_outputs(6260) <= (layer0_outputs(518)) or (layer0_outputs(5180));
    layer1_outputs(6261) <= not(layer0_outputs(1669)) or (layer0_outputs(145));
    layer1_outputs(6262) <= (layer0_outputs(2149)) or (layer0_outputs(6739));
    layer1_outputs(6263) <= (layer0_outputs(1122)) and not (layer0_outputs(6872));
    layer1_outputs(6264) <= layer0_outputs(2746);
    layer1_outputs(6265) <= layer0_outputs(6052);
    layer1_outputs(6266) <= not((layer0_outputs(7523)) and (layer0_outputs(3565)));
    layer1_outputs(6267) <= not(layer0_outputs(1342));
    layer1_outputs(6268) <= (layer0_outputs(4239)) or (layer0_outputs(4164));
    layer1_outputs(6269) <= (layer0_outputs(1156)) or (layer0_outputs(1713));
    layer1_outputs(6270) <= not(layer0_outputs(6390));
    layer1_outputs(6271) <= not(layer0_outputs(5441));
    layer1_outputs(6272) <= not(layer0_outputs(3852));
    layer1_outputs(6273) <= not(layer0_outputs(5822));
    layer1_outputs(6274) <= '1';
    layer1_outputs(6275) <= not(layer0_outputs(3235)) or (layer0_outputs(6380));
    layer1_outputs(6276) <= not((layer0_outputs(7195)) or (layer0_outputs(817)));
    layer1_outputs(6277) <= not(layer0_outputs(6300)) or (layer0_outputs(6144));
    layer1_outputs(6278) <= not((layer0_outputs(316)) or (layer0_outputs(4046)));
    layer1_outputs(6279) <= '1';
    layer1_outputs(6280) <= not((layer0_outputs(3292)) and (layer0_outputs(4197)));
    layer1_outputs(6281) <= (layer0_outputs(5750)) and not (layer0_outputs(6649));
    layer1_outputs(6282) <= layer0_outputs(845);
    layer1_outputs(6283) <= not(layer0_outputs(1165));
    layer1_outputs(6284) <= '1';
    layer1_outputs(6285) <= layer0_outputs(2896);
    layer1_outputs(6286) <= not(layer0_outputs(71));
    layer1_outputs(6287) <= not(layer0_outputs(3019)) or (layer0_outputs(3426));
    layer1_outputs(6288) <= layer0_outputs(6540);
    layer1_outputs(6289) <= not((layer0_outputs(1506)) and (layer0_outputs(5815)));
    layer1_outputs(6290) <= (layer0_outputs(5077)) or (layer0_outputs(5469));
    layer1_outputs(6291) <= not(layer0_outputs(737));
    layer1_outputs(6292) <= '1';
    layer1_outputs(6293) <= '0';
    layer1_outputs(6294) <= layer0_outputs(3638);
    layer1_outputs(6295) <= (layer0_outputs(3783)) xor (layer0_outputs(1319));
    layer1_outputs(6296) <= not(layer0_outputs(4901));
    layer1_outputs(6297) <= not(layer0_outputs(4969)) or (layer0_outputs(4749));
    layer1_outputs(6298) <= '1';
    layer1_outputs(6299) <= '1';
    layer1_outputs(6300) <= not(layer0_outputs(5249));
    layer1_outputs(6301) <= '1';
    layer1_outputs(6302) <= not(layer0_outputs(6543)) or (layer0_outputs(1366));
    layer1_outputs(6303) <= '1';
    layer1_outputs(6304) <= '0';
    layer1_outputs(6305) <= layer0_outputs(9);
    layer1_outputs(6306) <= (layer0_outputs(1495)) xor (layer0_outputs(858));
    layer1_outputs(6307) <= not(layer0_outputs(1970)) or (layer0_outputs(7559));
    layer1_outputs(6308) <= (layer0_outputs(6974)) and not (layer0_outputs(731));
    layer1_outputs(6309) <= not(layer0_outputs(5571));
    layer1_outputs(6310) <= not(layer0_outputs(6189));
    layer1_outputs(6311) <= '1';
    layer1_outputs(6312) <= not((layer0_outputs(5202)) and (layer0_outputs(6654)));
    layer1_outputs(6313) <= not(layer0_outputs(1649)) or (layer0_outputs(6000));
    layer1_outputs(6314) <= (layer0_outputs(936)) and not (layer0_outputs(2396));
    layer1_outputs(6315) <= layer0_outputs(2007);
    layer1_outputs(6316) <= (layer0_outputs(960)) or (layer0_outputs(1524));
    layer1_outputs(6317) <= not(layer0_outputs(4972)) or (layer0_outputs(5381));
    layer1_outputs(6318) <= (layer0_outputs(4744)) and (layer0_outputs(4047));
    layer1_outputs(6319) <= not((layer0_outputs(3495)) and (layer0_outputs(3884)));
    layer1_outputs(6320) <= (layer0_outputs(3958)) and not (layer0_outputs(3882));
    layer1_outputs(6321) <= not(layer0_outputs(29));
    layer1_outputs(6322) <= '0';
    layer1_outputs(6323) <= not(layer0_outputs(7162)) or (layer0_outputs(1381));
    layer1_outputs(6324) <= '0';
    layer1_outputs(6325) <= '1';
    layer1_outputs(6326) <= '0';
    layer1_outputs(6327) <= (layer0_outputs(3269)) or (layer0_outputs(7555));
    layer1_outputs(6328) <= not(layer0_outputs(115));
    layer1_outputs(6329) <= not((layer0_outputs(2097)) and (layer0_outputs(3489)));
    layer1_outputs(6330) <= not((layer0_outputs(5925)) and (layer0_outputs(5624)));
    layer1_outputs(6331) <= not(layer0_outputs(3438));
    layer1_outputs(6332) <= not(layer0_outputs(2689)) or (layer0_outputs(6488));
    layer1_outputs(6333) <= (layer0_outputs(6433)) and not (layer0_outputs(2614));
    layer1_outputs(6334) <= not((layer0_outputs(5309)) and (layer0_outputs(1066)));
    layer1_outputs(6335) <= not(layer0_outputs(3157)) or (layer0_outputs(2050));
    layer1_outputs(6336) <= not(layer0_outputs(1423));
    layer1_outputs(6337) <= '0';
    layer1_outputs(6338) <= (layer0_outputs(1255)) and (layer0_outputs(4279));
    layer1_outputs(6339) <= not(layer0_outputs(4171));
    layer1_outputs(6340) <= '1';
    layer1_outputs(6341) <= (layer0_outputs(4623)) and not (layer0_outputs(5109));
    layer1_outputs(6342) <= (layer0_outputs(4437)) and not (layer0_outputs(167));
    layer1_outputs(6343) <= not(layer0_outputs(1586)) or (layer0_outputs(4866));
    layer1_outputs(6344) <= '0';
    layer1_outputs(6345) <= not(layer0_outputs(2178)) or (layer0_outputs(606));
    layer1_outputs(6346) <= not(layer0_outputs(1988)) or (layer0_outputs(5342));
    layer1_outputs(6347) <= '1';
    layer1_outputs(6348) <= (layer0_outputs(2263)) and not (layer0_outputs(1752));
    layer1_outputs(6349) <= '1';
    layer1_outputs(6350) <= (layer0_outputs(664)) and not (layer0_outputs(581));
    layer1_outputs(6351) <= not(layer0_outputs(7061));
    layer1_outputs(6352) <= layer0_outputs(1030);
    layer1_outputs(6353) <= not(layer0_outputs(337)) or (layer0_outputs(1263));
    layer1_outputs(6354) <= layer0_outputs(6968);
    layer1_outputs(6355) <= not((layer0_outputs(3930)) or (layer0_outputs(4852)));
    layer1_outputs(6356) <= (layer0_outputs(3825)) and not (layer0_outputs(6152));
    layer1_outputs(6357) <= not(layer0_outputs(348)) or (layer0_outputs(1561));
    layer1_outputs(6358) <= layer0_outputs(4349);
    layer1_outputs(6359) <= (layer0_outputs(727)) and not (layer0_outputs(1440));
    layer1_outputs(6360) <= layer0_outputs(4601);
    layer1_outputs(6361) <= (layer0_outputs(5219)) and (layer0_outputs(5874));
    layer1_outputs(6362) <= (layer0_outputs(5316)) and not (layer0_outputs(6693));
    layer1_outputs(6363) <= (layer0_outputs(6351)) or (layer0_outputs(6740));
    layer1_outputs(6364) <= not((layer0_outputs(4163)) or (layer0_outputs(6215)));
    layer1_outputs(6365) <= (layer0_outputs(5508)) and not (layer0_outputs(7457));
    layer1_outputs(6366) <= (layer0_outputs(2424)) xor (layer0_outputs(3524));
    layer1_outputs(6367) <= (layer0_outputs(364)) and not (layer0_outputs(2613));
    layer1_outputs(6368) <= not(layer0_outputs(4602)) or (layer0_outputs(5380));
    layer1_outputs(6369) <= not(layer0_outputs(327)) or (layer0_outputs(3323));
    layer1_outputs(6370) <= layer0_outputs(2937);
    layer1_outputs(6371) <= layer0_outputs(5412);
    layer1_outputs(6372) <= '0';
    layer1_outputs(6373) <= '1';
    layer1_outputs(6374) <= (layer0_outputs(2118)) and not (layer0_outputs(1121));
    layer1_outputs(6375) <= layer0_outputs(5169);
    layer1_outputs(6376) <= '0';
    layer1_outputs(6377) <= not(layer0_outputs(1723)) or (layer0_outputs(2074));
    layer1_outputs(6378) <= layer0_outputs(4445);
    layer1_outputs(6379) <= not(layer0_outputs(665));
    layer1_outputs(6380) <= (layer0_outputs(5364)) and not (layer0_outputs(5010));
    layer1_outputs(6381) <= '0';
    layer1_outputs(6382) <= not((layer0_outputs(1710)) and (layer0_outputs(1897)));
    layer1_outputs(6383) <= not(layer0_outputs(297)) or (layer0_outputs(1082));
    layer1_outputs(6384) <= (layer0_outputs(6795)) and not (layer0_outputs(1005));
    layer1_outputs(6385) <= (layer0_outputs(2282)) and (layer0_outputs(467));
    layer1_outputs(6386) <= (layer0_outputs(1265)) and not (layer0_outputs(7289));
    layer1_outputs(6387) <= not(layer0_outputs(1288));
    layer1_outputs(6388) <= layer0_outputs(4848);
    layer1_outputs(6389) <= not(layer0_outputs(2905));
    layer1_outputs(6390) <= not(layer0_outputs(783));
    layer1_outputs(6391) <= not(layer0_outputs(4239));
    layer1_outputs(6392) <= (layer0_outputs(4166)) and not (layer0_outputs(3943));
    layer1_outputs(6393) <= '1';
    layer1_outputs(6394) <= not(layer0_outputs(4268));
    layer1_outputs(6395) <= not(layer0_outputs(128)) or (layer0_outputs(5498));
    layer1_outputs(6396) <= '0';
    layer1_outputs(6397) <= (layer0_outputs(2430)) and not (layer0_outputs(7656));
    layer1_outputs(6398) <= layer0_outputs(5784);
    layer1_outputs(6399) <= (layer0_outputs(5664)) or (layer0_outputs(209));
    layer1_outputs(6400) <= (layer0_outputs(851)) or (layer0_outputs(2442));
    layer1_outputs(6401) <= (layer0_outputs(6908)) and (layer0_outputs(1821));
    layer1_outputs(6402) <= not(layer0_outputs(5059));
    layer1_outputs(6403) <= '1';
    layer1_outputs(6404) <= (layer0_outputs(2195)) or (layer0_outputs(7598));
    layer1_outputs(6405) <= layer0_outputs(6384);
    layer1_outputs(6406) <= '0';
    layer1_outputs(6407) <= '1';
    layer1_outputs(6408) <= layer0_outputs(6141);
    layer1_outputs(6409) <= layer0_outputs(512);
    layer1_outputs(6410) <= layer0_outputs(812);
    layer1_outputs(6411) <= (layer0_outputs(5332)) and not (layer0_outputs(740));
    layer1_outputs(6412) <= not(layer0_outputs(1968)) or (layer0_outputs(2602));
    layer1_outputs(6413) <= (layer0_outputs(6019)) and not (layer0_outputs(5369));
    layer1_outputs(6414) <= layer0_outputs(1835);
    layer1_outputs(6415) <= '0';
    layer1_outputs(6416) <= not((layer0_outputs(6623)) or (layer0_outputs(3177)));
    layer1_outputs(6417) <= '0';
    layer1_outputs(6418) <= (layer0_outputs(3737)) or (layer0_outputs(2462));
    layer1_outputs(6419) <= not(layer0_outputs(2782));
    layer1_outputs(6420) <= not(layer0_outputs(4388));
    layer1_outputs(6421) <= not((layer0_outputs(3052)) or (layer0_outputs(730)));
    layer1_outputs(6422) <= '0';
    layer1_outputs(6423) <= layer0_outputs(7246);
    layer1_outputs(6424) <= (layer0_outputs(640)) and (layer0_outputs(4774));
    layer1_outputs(6425) <= (layer0_outputs(2454)) and (layer0_outputs(5816));
    layer1_outputs(6426) <= (layer0_outputs(2404)) and (layer0_outputs(3244));
    layer1_outputs(6427) <= not((layer0_outputs(7252)) or (layer0_outputs(5838)));
    layer1_outputs(6428) <= '1';
    layer1_outputs(6429) <= layer0_outputs(2091);
    layer1_outputs(6430) <= (layer0_outputs(6762)) and (layer0_outputs(5032));
    layer1_outputs(6431) <= '0';
    layer1_outputs(6432) <= '0';
    layer1_outputs(6433) <= not(layer0_outputs(5696)) or (layer0_outputs(3023));
    layer1_outputs(6434) <= not(layer0_outputs(53)) or (layer0_outputs(1804));
    layer1_outputs(6435) <= (layer0_outputs(382)) and (layer0_outputs(7572));
    layer1_outputs(6436) <= not(layer0_outputs(4024));
    layer1_outputs(6437) <= layer0_outputs(648);
    layer1_outputs(6438) <= '0';
    layer1_outputs(6439) <= (layer0_outputs(4961)) and not (layer0_outputs(5037));
    layer1_outputs(6440) <= (layer0_outputs(1185)) or (layer0_outputs(5493));
    layer1_outputs(6441) <= not(layer0_outputs(377));
    layer1_outputs(6442) <= not(layer0_outputs(696));
    layer1_outputs(6443) <= not(layer0_outputs(7128)) or (layer0_outputs(4365));
    layer1_outputs(6444) <= (layer0_outputs(4101)) and (layer0_outputs(5631));
    layer1_outputs(6445) <= (layer0_outputs(1571)) and not (layer0_outputs(6162));
    layer1_outputs(6446) <= not(layer0_outputs(1089)) or (layer0_outputs(7204));
    layer1_outputs(6447) <= layer0_outputs(4646);
    layer1_outputs(6448) <= '1';
    layer1_outputs(6449) <= '1';
    layer1_outputs(6450) <= not(layer0_outputs(4286)) or (layer0_outputs(7590));
    layer1_outputs(6451) <= (layer0_outputs(7090)) or (layer0_outputs(5929));
    layer1_outputs(6452) <= not((layer0_outputs(6610)) or (layer0_outputs(550)));
    layer1_outputs(6453) <= layer0_outputs(1300);
    layer1_outputs(6454) <= layer0_outputs(5757);
    layer1_outputs(6455) <= layer0_outputs(923);
    layer1_outputs(6456) <= not((layer0_outputs(1824)) and (layer0_outputs(1017)));
    layer1_outputs(6457) <= not((layer0_outputs(5662)) or (layer0_outputs(5834)));
    layer1_outputs(6458) <= '0';
    layer1_outputs(6459) <= '0';
    layer1_outputs(6460) <= not((layer0_outputs(7261)) and (layer0_outputs(5403)));
    layer1_outputs(6461) <= not(layer0_outputs(5821));
    layer1_outputs(6462) <= (layer0_outputs(1159)) and not (layer0_outputs(4127));
    layer1_outputs(6463) <= not(layer0_outputs(5263));
    layer1_outputs(6464) <= not((layer0_outputs(5825)) or (layer0_outputs(3193)));
    layer1_outputs(6465) <= not(layer0_outputs(3004));
    layer1_outputs(6466) <= not(layer0_outputs(6656)) or (layer0_outputs(1846));
    layer1_outputs(6467) <= (layer0_outputs(1693)) or (layer0_outputs(2960));
    layer1_outputs(6468) <= '1';
    layer1_outputs(6469) <= (layer0_outputs(7519)) and not (layer0_outputs(3822));
    layer1_outputs(6470) <= '1';
    layer1_outputs(6471) <= not((layer0_outputs(1729)) or (layer0_outputs(7675)));
    layer1_outputs(6472) <= (layer0_outputs(3314)) or (layer0_outputs(1139));
    layer1_outputs(6473) <= layer0_outputs(6278);
    layer1_outputs(6474) <= layer0_outputs(1130);
    layer1_outputs(6475) <= not(layer0_outputs(6740));
    layer1_outputs(6476) <= not(layer0_outputs(2400)) or (layer0_outputs(6476));
    layer1_outputs(6477) <= (layer0_outputs(3282)) and not (layer0_outputs(4484));
    layer1_outputs(6478) <= layer0_outputs(680);
    layer1_outputs(6479) <= not(layer0_outputs(7603)) or (layer0_outputs(3605));
    layer1_outputs(6480) <= not(layer0_outputs(4341)) or (layer0_outputs(2969));
    layer1_outputs(6481) <= not(layer0_outputs(7505));
    layer1_outputs(6482) <= not(layer0_outputs(2371)) or (layer0_outputs(6959));
    layer1_outputs(6483) <= '1';
    layer1_outputs(6484) <= layer0_outputs(4569);
    layer1_outputs(6485) <= layer0_outputs(4874);
    layer1_outputs(6486) <= (layer0_outputs(4240)) and (layer0_outputs(3582));
    layer1_outputs(6487) <= (layer0_outputs(3473)) or (layer0_outputs(6702));
    layer1_outputs(6488) <= (layer0_outputs(7613)) and not (layer0_outputs(3095));
    layer1_outputs(6489) <= (layer0_outputs(3401)) and not (layer0_outputs(1302));
    layer1_outputs(6490) <= not((layer0_outputs(315)) or (layer0_outputs(3761)));
    layer1_outputs(6491) <= '1';
    layer1_outputs(6492) <= layer0_outputs(1952);
    layer1_outputs(6493) <= '1';
    layer1_outputs(6494) <= '0';
    layer1_outputs(6495) <= not(layer0_outputs(1259)) or (layer0_outputs(2088));
    layer1_outputs(6496) <= not(layer0_outputs(7270));
    layer1_outputs(6497) <= (layer0_outputs(3499)) and (layer0_outputs(3022));
    layer1_outputs(6498) <= (layer0_outputs(3791)) and not (layer0_outputs(5751));
    layer1_outputs(6499) <= not((layer0_outputs(5406)) and (layer0_outputs(6503)));
    layer1_outputs(6500) <= (layer0_outputs(3164)) or (layer0_outputs(5968));
    layer1_outputs(6501) <= (layer0_outputs(3343)) and not (layer0_outputs(3559));
    layer1_outputs(6502) <= not(layer0_outputs(2921)) or (layer0_outputs(4174));
    layer1_outputs(6503) <= layer0_outputs(5515);
    layer1_outputs(6504) <= '0';
    layer1_outputs(6505) <= '1';
    layer1_outputs(6506) <= (layer0_outputs(1547)) or (layer0_outputs(2597));
    layer1_outputs(6507) <= '1';
    layer1_outputs(6508) <= (layer0_outputs(2217)) and (layer0_outputs(4064));
    layer1_outputs(6509) <= '0';
    layer1_outputs(6510) <= not(layer0_outputs(3227));
    layer1_outputs(6511) <= not((layer0_outputs(261)) and (layer0_outputs(4930)));
    layer1_outputs(6512) <= (layer0_outputs(4344)) or (layer0_outputs(3780));
    layer1_outputs(6513) <= (layer0_outputs(2084)) or (layer0_outputs(5129));
    layer1_outputs(6514) <= layer0_outputs(6215);
    layer1_outputs(6515) <= '0';
    layer1_outputs(6516) <= not((layer0_outputs(3330)) or (layer0_outputs(6625)));
    layer1_outputs(6517) <= (layer0_outputs(2583)) and not (layer0_outputs(1760));
    layer1_outputs(6518) <= (layer0_outputs(767)) and not (layer0_outputs(1704));
    layer1_outputs(6519) <= (layer0_outputs(7470)) or (layer0_outputs(895));
    layer1_outputs(6520) <= (layer0_outputs(349)) and (layer0_outputs(4250));
    layer1_outputs(6521) <= not((layer0_outputs(4413)) and (layer0_outputs(3233)));
    layer1_outputs(6522) <= (layer0_outputs(6554)) xor (layer0_outputs(1611));
    layer1_outputs(6523) <= not((layer0_outputs(4846)) and (layer0_outputs(7667)));
    layer1_outputs(6524) <= layer0_outputs(2787);
    layer1_outputs(6525) <= (layer0_outputs(1829)) and not (layer0_outputs(5733));
    layer1_outputs(6526) <= not((layer0_outputs(3195)) or (layer0_outputs(869)));
    layer1_outputs(6527) <= not(layer0_outputs(1315)) or (layer0_outputs(7242));
    layer1_outputs(6528) <= (layer0_outputs(3496)) and (layer0_outputs(2466));
    layer1_outputs(6529) <= layer0_outputs(2374);
    layer1_outputs(6530) <= not((layer0_outputs(2531)) and (layer0_outputs(78)));
    layer1_outputs(6531) <= layer0_outputs(781);
    layer1_outputs(6532) <= '0';
    layer1_outputs(6533) <= '0';
    layer1_outputs(6534) <= (layer0_outputs(2715)) and not (layer0_outputs(1774));
    layer1_outputs(6535) <= not((layer0_outputs(1915)) and (layer0_outputs(6025)));
    layer1_outputs(6536) <= '1';
    layer1_outputs(6537) <= (layer0_outputs(4271)) and (layer0_outputs(1140));
    layer1_outputs(6538) <= layer0_outputs(3801);
    layer1_outputs(6539) <= not(layer0_outputs(5092)) or (layer0_outputs(6119));
    layer1_outputs(6540) <= layer0_outputs(5872);
    layer1_outputs(6541) <= not(layer0_outputs(4997));
    layer1_outputs(6542) <= not((layer0_outputs(3609)) and (layer0_outputs(2314)));
    layer1_outputs(6543) <= not((layer0_outputs(1582)) and (layer0_outputs(5311)));
    layer1_outputs(6544) <= (layer0_outputs(5786)) and not (layer0_outputs(3319));
    layer1_outputs(6545) <= layer0_outputs(6891);
    layer1_outputs(6546) <= not(layer0_outputs(5162)) or (layer0_outputs(6252));
    layer1_outputs(6547) <= not(layer0_outputs(5065)) or (layer0_outputs(1096));
    layer1_outputs(6548) <= not(layer0_outputs(5963));
    layer1_outputs(6549) <= not((layer0_outputs(5142)) or (layer0_outputs(7097)));
    layer1_outputs(6550) <= not((layer0_outputs(6726)) and (layer0_outputs(7364)));
    layer1_outputs(6551) <= '1';
    layer1_outputs(6552) <= not(layer0_outputs(3656)) or (layer0_outputs(3200));
    layer1_outputs(6553) <= not(layer0_outputs(1542));
    layer1_outputs(6554) <= not((layer0_outputs(5216)) and (layer0_outputs(1929)));
    layer1_outputs(6555) <= not(layer0_outputs(239));
    layer1_outputs(6556) <= (layer0_outputs(97)) and not (layer0_outputs(6664));
    layer1_outputs(6557) <= (layer0_outputs(3441)) and not (layer0_outputs(3581));
    layer1_outputs(6558) <= not(layer0_outputs(5319)) or (layer0_outputs(6875));
    layer1_outputs(6559) <= layer0_outputs(4465);
    layer1_outputs(6560) <= '0';
    layer1_outputs(6561) <= layer0_outputs(7549);
    layer1_outputs(6562) <= not(layer0_outputs(1707));
    layer1_outputs(6563) <= not((layer0_outputs(1687)) or (layer0_outputs(6042)));
    layer1_outputs(6564) <= not(layer0_outputs(5818)) or (layer0_outputs(669));
    layer1_outputs(6565) <= (layer0_outputs(5239)) and not (layer0_outputs(4742));
    layer1_outputs(6566) <= '0';
    layer1_outputs(6567) <= not((layer0_outputs(434)) and (layer0_outputs(5567)));
    layer1_outputs(6568) <= not(layer0_outputs(601));
    layer1_outputs(6569) <= '1';
    layer1_outputs(6570) <= not(layer0_outputs(4333));
    layer1_outputs(6571) <= (layer0_outputs(2075)) and not (layer0_outputs(78));
    layer1_outputs(6572) <= '1';
    layer1_outputs(6573) <= layer0_outputs(336);
    layer1_outputs(6574) <= (layer0_outputs(2652)) and (layer0_outputs(6626));
    layer1_outputs(6575) <= layer0_outputs(4395);
    layer1_outputs(6576) <= '0';
    layer1_outputs(6577) <= '0';
    layer1_outputs(6578) <= layer0_outputs(5943);
    layer1_outputs(6579) <= layer0_outputs(5853);
    layer1_outputs(6580) <= '1';
    layer1_outputs(6581) <= layer0_outputs(4709);
    layer1_outputs(6582) <= layer0_outputs(4295);
    layer1_outputs(6583) <= not(layer0_outputs(4306)) or (layer0_outputs(543));
    layer1_outputs(6584) <= '0';
    layer1_outputs(6585) <= not(layer0_outputs(4837));
    layer1_outputs(6586) <= '0';
    layer1_outputs(6587) <= layer0_outputs(3193);
    layer1_outputs(6588) <= not(layer0_outputs(1156)) or (layer0_outputs(2833));
    layer1_outputs(6589) <= (layer0_outputs(476)) and (layer0_outputs(5770));
    layer1_outputs(6590) <= '0';
    layer1_outputs(6591) <= '1';
    layer1_outputs(6592) <= layer0_outputs(827);
    layer1_outputs(6593) <= layer0_outputs(7278);
    layer1_outputs(6594) <= '1';
    layer1_outputs(6595) <= layer0_outputs(2775);
    layer1_outputs(6596) <= '1';
    layer1_outputs(6597) <= (layer0_outputs(2543)) and (layer0_outputs(3808));
    layer1_outputs(6598) <= '0';
    layer1_outputs(6599) <= not(layer0_outputs(3737));
    layer1_outputs(6600) <= layer0_outputs(7655);
    layer1_outputs(6601) <= '1';
    layer1_outputs(6602) <= '0';
    layer1_outputs(6603) <= (layer0_outputs(6842)) and not (layer0_outputs(2132));
    layer1_outputs(6604) <= not((layer0_outputs(3488)) and (layer0_outputs(4267)));
    layer1_outputs(6605) <= '0';
    layer1_outputs(6606) <= not(layer0_outputs(4221));
    layer1_outputs(6607) <= not(layer0_outputs(4547)) or (layer0_outputs(7415));
    layer1_outputs(6608) <= not(layer0_outputs(5278)) or (layer0_outputs(7044));
    layer1_outputs(6609) <= layer0_outputs(2462);
    layer1_outputs(6610) <= not((layer0_outputs(4919)) and (layer0_outputs(6998)));
    layer1_outputs(6611) <= (layer0_outputs(2569)) or (layer0_outputs(3281));
    layer1_outputs(6612) <= not(layer0_outputs(2771));
    layer1_outputs(6613) <= (layer0_outputs(4568)) and (layer0_outputs(3278));
    layer1_outputs(6614) <= layer0_outputs(1733);
    layer1_outputs(6615) <= (layer0_outputs(6104)) or (layer0_outputs(3632));
    layer1_outputs(6616) <= '1';
    layer1_outputs(6617) <= not(layer0_outputs(354));
    layer1_outputs(6618) <= not(layer0_outputs(2844));
    layer1_outputs(6619) <= '0';
    layer1_outputs(6620) <= (layer0_outputs(3049)) and not (layer0_outputs(1211));
    layer1_outputs(6621) <= (layer0_outputs(6494)) and not (layer0_outputs(4279));
    layer1_outputs(6622) <= layer0_outputs(6282);
    layer1_outputs(6623) <= layer0_outputs(4765);
    layer1_outputs(6624) <= not(layer0_outputs(57));
    layer1_outputs(6625) <= not(layer0_outputs(4242));
    layer1_outputs(6626) <= '1';
    layer1_outputs(6627) <= not(layer0_outputs(3677)) or (layer0_outputs(2058));
    layer1_outputs(6628) <= (layer0_outputs(7286)) and (layer0_outputs(1171));
    layer1_outputs(6629) <= (layer0_outputs(2474)) or (layer0_outputs(2004));
    layer1_outputs(6630) <= layer0_outputs(5492);
    layer1_outputs(6631) <= not((layer0_outputs(1359)) and (layer0_outputs(4235)));
    layer1_outputs(6632) <= (layer0_outputs(2756)) and not (layer0_outputs(5876));
    layer1_outputs(6633) <= (layer0_outputs(6238)) and (layer0_outputs(6844));
    layer1_outputs(6634) <= (layer0_outputs(1509)) and not (layer0_outputs(6987));
    layer1_outputs(6635) <= not((layer0_outputs(393)) or (layer0_outputs(379)));
    layer1_outputs(6636) <= not(layer0_outputs(3025)) or (layer0_outputs(841));
    layer1_outputs(6637) <= not(layer0_outputs(2141));
    layer1_outputs(6638) <= not(layer0_outputs(4893));
    layer1_outputs(6639) <= (layer0_outputs(6028)) and not (layer0_outputs(4989));
    layer1_outputs(6640) <= not(layer0_outputs(34)) or (layer0_outputs(6078));
    layer1_outputs(6641) <= layer0_outputs(6751);
    layer1_outputs(6642) <= '1';
    layer1_outputs(6643) <= (layer0_outputs(6644)) xor (layer0_outputs(5227));
    layer1_outputs(6644) <= not(layer0_outputs(418)) or (layer0_outputs(4210));
    layer1_outputs(6645) <= (layer0_outputs(2878)) and (layer0_outputs(1176));
    layer1_outputs(6646) <= not(layer0_outputs(5777)) or (layer0_outputs(6844));
    layer1_outputs(6647) <= not((layer0_outputs(6723)) or (layer0_outputs(4006)));
    layer1_outputs(6648) <= (layer0_outputs(4466)) or (layer0_outputs(2569));
    layer1_outputs(6649) <= not(layer0_outputs(2868));
    layer1_outputs(6650) <= not((layer0_outputs(6338)) and (layer0_outputs(2242)));
    layer1_outputs(6651) <= not(layer0_outputs(2752));
    layer1_outputs(6652) <= '1';
    layer1_outputs(6653) <= '0';
    layer1_outputs(6654) <= layer0_outputs(1862);
    layer1_outputs(6655) <= (layer0_outputs(7426)) or (layer0_outputs(5173));
    layer1_outputs(6656) <= (layer0_outputs(2271)) and not (layer0_outputs(3776));
    layer1_outputs(6657) <= (layer0_outputs(2651)) or (layer0_outputs(1043));
    layer1_outputs(6658) <= not(layer0_outputs(2948));
    layer1_outputs(6659) <= not((layer0_outputs(2389)) and (layer0_outputs(5218)));
    layer1_outputs(6660) <= not((layer0_outputs(2257)) or (layer0_outputs(2685)));
    layer1_outputs(6661) <= not(layer0_outputs(6291));
    layer1_outputs(6662) <= '1';
    layer1_outputs(6663) <= not(layer0_outputs(3327)) or (layer0_outputs(602));
    layer1_outputs(6664) <= not(layer0_outputs(2976));
    layer1_outputs(6665) <= (layer0_outputs(6584)) and not (layer0_outputs(2959));
    layer1_outputs(6666) <= (layer0_outputs(3082)) or (layer0_outputs(4968));
    layer1_outputs(6667) <= '1';
    layer1_outputs(6668) <= not(layer0_outputs(6864)) or (layer0_outputs(1435));
    layer1_outputs(6669) <= '0';
    layer1_outputs(6670) <= (layer0_outputs(6614)) or (layer0_outputs(3867));
    layer1_outputs(6671) <= not(layer0_outputs(6196));
    layer1_outputs(6672) <= layer0_outputs(4896);
    layer1_outputs(6673) <= layer0_outputs(3081);
    layer1_outputs(6674) <= layer0_outputs(4407);
    layer1_outputs(6675) <= (layer0_outputs(1708)) and not (layer0_outputs(262));
    layer1_outputs(6676) <= not((layer0_outputs(668)) xor (layer0_outputs(4032)));
    layer1_outputs(6677) <= not(layer0_outputs(6499));
    layer1_outputs(6678) <= (layer0_outputs(1959)) and not (layer0_outputs(1367));
    layer1_outputs(6679) <= '1';
    layer1_outputs(6680) <= (layer0_outputs(5630)) and not (layer0_outputs(1863));
    layer1_outputs(6681) <= not(layer0_outputs(3093));
    layer1_outputs(6682) <= not((layer0_outputs(2572)) and (layer0_outputs(907)));
    layer1_outputs(6683) <= '1';
    layer1_outputs(6684) <= (layer0_outputs(7469)) and (layer0_outputs(1238));
    layer1_outputs(6685) <= not(layer0_outputs(6708)) or (layer0_outputs(367));
    layer1_outputs(6686) <= (layer0_outputs(5847)) and (layer0_outputs(2485));
    layer1_outputs(6687) <= (layer0_outputs(6371)) and not (layer0_outputs(1825));
    layer1_outputs(6688) <= (layer0_outputs(7141)) and not (layer0_outputs(1526));
    layer1_outputs(6689) <= '0';
    layer1_outputs(6690) <= not(layer0_outputs(5756)) or (layer0_outputs(2824));
    layer1_outputs(6691) <= (layer0_outputs(3284)) or (layer0_outputs(1101));
    layer1_outputs(6692) <= (layer0_outputs(6323)) and (layer0_outputs(6804));
    layer1_outputs(6693) <= not(layer0_outputs(5361)) or (layer0_outputs(5341));
    layer1_outputs(6694) <= not(layer0_outputs(2729));
    layer1_outputs(6695) <= not((layer0_outputs(3142)) or (layer0_outputs(7446)));
    layer1_outputs(6696) <= '0';
    layer1_outputs(6697) <= not(layer0_outputs(3942));
    layer1_outputs(6698) <= (layer0_outputs(4133)) or (layer0_outputs(925));
    layer1_outputs(6699) <= not(layer0_outputs(180)) or (layer0_outputs(856));
    layer1_outputs(6700) <= (layer0_outputs(3554)) or (layer0_outputs(260));
    layer1_outputs(6701) <= layer0_outputs(7281);
    layer1_outputs(6702) <= not(layer0_outputs(7243)) or (layer0_outputs(5788));
    layer1_outputs(6703) <= '0';
    layer1_outputs(6704) <= (layer0_outputs(2527)) and not (layer0_outputs(970));
    layer1_outputs(6705) <= (layer0_outputs(1220)) or (layer0_outputs(7050));
    layer1_outputs(6706) <= '0';
    layer1_outputs(6707) <= layer0_outputs(6222);
    layer1_outputs(6708) <= (layer0_outputs(3238)) and not (layer0_outputs(2486));
    layer1_outputs(6709) <= (layer0_outputs(7004)) and not (layer0_outputs(3067));
    layer1_outputs(6710) <= layer0_outputs(3871);
    layer1_outputs(6711) <= '1';
    layer1_outputs(6712) <= not(layer0_outputs(6973));
    layer1_outputs(6713) <= not(layer0_outputs(1892));
    layer1_outputs(6714) <= (layer0_outputs(4763)) or (layer0_outputs(3530));
    layer1_outputs(6715) <= not((layer0_outputs(7220)) or (layer0_outputs(2586)));
    layer1_outputs(6716) <= (layer0_outputs(7063)) and not (layer0_outputs(5302));
    layer1_outputs(6717) <= not((layer0_outputs(2342)) and (layer0_outputs(3519)));
    layer1_outputs(6718) <= (layer0_outputs(4080)) and not (layer0_outputs(3735));
    layer1_outputs(6719) <= not(layer0_outputs(4891)) or (layer0_outputs(2418));
    layer1_outputs(6720) <= (layer0_outputs(4305)) and not (layer0_outputs(6254));
    layer1_outputs(6721) <= '0';
    layer1_outputs(6722) <= '0';
    layer1_outputs(6723) <= (layer0_outputs(7514)) and not (layer0_outputs(6594));
    layer1_outputs(6724) <= (layer0_outputs(5463)) and not (layer0_outputs(4857));
    layer1_outputs(6725) <= (layer0_outputs(1313)) xor (layer0_outputs(6432));
    layer1_outputs(6726) <= (layer0_outputs(6605)) or (layer0_outputs(2839));
    layer1_outputs(6727) <= (layer0_outputs(4749)) and not (layer0_outputs(7489));
    layer1_outputs(6728) <= '1';
    layer1_outputs(6729) <= layer0_outputs(6559);
    layer1_outputs(6730) <= not(layer0_outputs(5964)) or (layer0_outputs(6651));
    layer1_outputs(6731) <= (layer0_outputs(666)) or (layer0_outputs(4632));
    layer1_outputs(6732) <= not(layer0_outputs(2791)) or (layer0_outputs(3403));
    layer1_outputs(6733) <= '1';
    layer1_outputs(6734) <= '1';
    layer1_outputs(6735) <= '0';
    layer1_outputs(6736) <= (layer0_outputs(6337)) and (layer0_outputs(3514));
    layer1_outputs(6737) <= layer0_outputs(1322);
    layer1_outputs(6738) <= layer0_outputs(324);
    layer1_outputs(6739) <= (layer0_outputs(1695)) or (layer0_outputs(1426));
    layer1_outputs(6740) <= not(layer0_outputs(4028));
    layer1_outputs(6741) <= not(layer0_outputs(51));
    layer1_outputs(6742) <= not((layer0_outputs(3291)) or (layer0_outputs(2691)));
    layer1_outputs(6743) <= '1';
    layer1_outputs(6744) <= not(layer0_outputs(3153));
    layer1_outputs(6745) <= not((layer0_outputs(7331)) or (layer0_outputs(6291)));
    layer1_outputs(6746) <= not((layer0_outputs(5437)) and (layer0_outputs(613)));
    layer1_outputs(6747) <= not(layer0_outputs(6711));
    layer1_outputs(6748) <= not(layer0_outputs(5699)) or (layer0_outputs(1424));
    layer1_outputs(6749) <= not((layer0_outputs(3204)) or (layer0_outputs(3015)));
    layer1_outputs(6750) <= (layer0_outputs(870)) and (layer0_outputs(3437));
    layer1_outputs(6751) <= not(layer0_outputs(1979));
    layer1_outputs(6752) <= (layer0_outputs(365)) and not (layer0_outputs(6901));
    layer1_outputs(6753) <= not((layer0_outputs(1223)) and (layer0_outputs(7567)));
    layer1_outputs(6754) <= not((layer0_outputs(3543)) and (layer0_outputs(4168)));
    layer1_outputs(6755) <= layer0_outputs(4953);
    layer1_outputs(6756) <= not(layer0_outputs(6454));
    layer1_outputs(6757) <= not((layer0_outputs(2188)) and (layer0_outputs(3131)));
    layer1_outputs(6758) <= not(layer0_outputs(6539));
    layer1_outputs(6759) <= layer0_outputs(722);
    layer1_outputs(6760) <= not((layer0_outputs(6401)) or (layer0_outputs(2177)));
    layer1_outputs(6761) <= (layer0_outputs(2056)) and (layer0_outputs(156));
    layer1_outputs(6762) <= not(layer0_outputs(4658));
    layer1_outputs(6763) <= (layer0_outputs(5063)) and not (layer0_outputs(6742));
    layer1_outputs(6764) <= '0';
    layer1_outputs(6765) <= not(layer0_outputs(7013));
    layer1_outputs(6766) <= (layer0_outputs(4590)) and (layer0_outputs(3862));
    layer1_outputs(6767) <= not(layer0_outputs(3268));
    layer1_outputs(6768) <= '1';
    layer1_outputs(6769) <= not(layer0_outputs(603));
    layer1_outputs(6770) <= '0';
    layer1_outputs(6771) <= '1';
    layer1_outputs(6772) <= not(layer0_outputs(1277));
    layer1_outputs(6773) <= not(layer0_outputs(5450));
    layer1_outputs(6774) <= (layer0_outputs(438)) and not (layer0_outputs(4055));
    layer1_outputs(6775) <= (layer0_outputs(4842)) and not (layer0_outputs(5846));
    layer1_outputs(6776) <= layer0_outputs(1145);
    layer1_outputs(6777) <= layer0_outputs(3857);
    layer1_outputs(6778) <= not((layer0_outputs(1816)) or (layer0_outputs(1989)));
    layer1_outputs(6779) <= layer0_outputs(4786);
    layer1_outputs(6780) <= layer0_outputs(574);
    layer1_outputs(6781) <= '1';
    layer1_outputs(6782) <= not(layer0_outputs(32)) or (layer0_outputs(174));
    layer1_outputs(6783) <= layer0_outputs(6393);
    layer1_outputs(6784) <= '1';
    layer1_outputs(6785) <= not(layer0_outputs(43));
    layer1_outputs(6786) <= not(layer0_outputs(2831)) or (layer0_outputs(2513));
    layer1_outputs(6787) <= not(layer0_outputs(1947));
    layer1_outputs(6788) <= (layer0_outputs(4339)) and (layer0_outputs(2149));
    layer1_outputs(6789) <= not((layer0_outputs(4133)) and (layer0_outputs(5359)));
    layer1_outputs(6790) <= (layer0_outputs(1103)) and (layer0_outputs(2237));
    layer1_outputs(6791) <= not((layer0_outputs(2736)) or (layer0_outputs(2165)));
    layer1_outputs(6792) <= (layer0_outputs(5948)) and (layer0_outputs(5221));
    layer1_outputs(6793) <= (layer0_outputs(4053)) or (layer0_outputs(6699));
    layer1_outputs(6794) <= '0';
    layer1_outputs(6795) <= '0';
    layer1_outputs(6796) <= not(layer0_outputs(1791));
    layer1_outputs(6797) <= '1';
    layer1_outputs(6798) <= not(layer0_outputs(1122));
    layer1_outputs(6799) <= not(layer0_outputs(1548)) or (layer0_outputs(1226));
    layer1_outputs(6800) <= (layer0_outputs(6600)) and not (layer0_outputs(431));
    layer1_outputs(6801) <= (layer0_outputs(2884)) and (layer0_outputs(3069));
    layer1_outputs(6802) <= layer0_outputs(4686);
    layer1_outputs(6803) <= '0';
    layer1_outputs(6804) <= (layer0_outputs(1257)) and not (layer0_outputs(6684));
    layer1_outputs(6805) <= (layer0_outputs(312)) or (layer0_outputs(5705));
    layer1_outputs(6806) <= not((layer0_outputs(4941)) xor (layer0_outputs(833)));
    layer1_outputs(6807) <= not((layer0_outputs(7477)) and (layer0_outputs(7279)));
    layer1_outputs(6808) <= '1';
    layer1_outputs(6809) <= '1';
    layer1_outputs(6810) <= (layer0_outputs(1074)) and not (layer0_outputs(5253));
    layer1_outputs(6811) <= not(layer0_outputs(4271)) or (layer0_outputs(814));
    layer1_outputs(6812) <= '0';
    layer1_outputs(6813) <= not(layer0_outputs(5426));
    layer1_outputs(6814) <= layer0_outputs(4599);
    layer1_outputs(6815) <= '1';
    layer1_outputs(6816) <= not(layer0_outputs(589));
    layer1_outputs(6817) <= (layer0_outputs(4699)) and not (layer0_outputs(6980));
    layer1_outputs(6818) <= layer0_outputs(301);
    layer1_outputs(6819) <= (layer0_outputs(4183)) and (layer0_outputs(7088));
    layer1_outputs(6820) <= (layer0_outputs(4141)) and not (layer0_outputs(2245));
    layer1_outputs(6821) <= not((layer0_outputs(2339)) or (layer0_outputs(1678)));
    layer1_outputs(6822) <= not(layer0_outputs(5197)) or (layer0_outputs(3210));
    layer1_outputs(6823) <= (layer0_outputs(1939)) or (layer0_outputs(3572));
    layer1_outputs(6824) <= not(layer0_outputs(5618));
    layer1_outputs(6825) <= (layer0_outputs(1275)) and (layer0_outputs(2351));
    layer1_outputs(6826) <= not(layer0_outputs(5673));
    layer1_outputs(6827) <= '0';
    layer1_outputs(6828) <= not(layer0_outputs(5652)) or (layer0_outputs(6015));
    layer1_outputs(6829) <= not(layer0_outputs(6241)) or (layer0_outputs(2127));
    layer1_outputs(6830) <= '0';
    layer1_outputs(6831) <= not(layer0_outputs(3696));
    layer1_outputs(6832) <= (layer0_outputs(7214)) and (layer0_outputs(2228));
    layer1_outputs(6833) <= not(layer0_outputs(7581));
    layer1_outputs(6834) <= layer0_outputs(5434);
    layer1_outputs(6835) <= (layer0_outputs(2464)) and not (layer0_outputs(2705));
    layer1_outputs(6836) <= '1';
    layer1_outputs(6837) <= '0';
    layer1_outputs(6838) <= not(layer0_outputs(1166));
    layer1_outputs(6839) <= not(layer0_outputs(4249));
    layer1_outputs(6840) <= (layer0_outputs(2291)) and not (layer0_outputs(5785));
    layer1_outputs(6841) <= '1';
    layer1_outputs(6842) <= not((layer0_outputs(4811)) and (layer0_outputs(5646)));
    layer1_outputs(6843) <= not(layer0_outputs(6889));
    layer1_outputs(6844) <= layer0_outputs(6004);
    layer1_outputs(6845) <= not(layer0_outputs(252));
    layer1_outputs(6846) <= not(layer0_outputs(7115));
    layer1_outputs(6847) <= (layer0_outputs(2778)) and not (layer0_outputs(5287));
    layer1_outputs(6848) <= not(layer0_outputs(5006)) or (layer0_outputs(2303));
    layer1_outputs(6849) <= layer0_outputs(5689);
    layer1_outputs(6850) <= (layer0_outputs(229)) and not (layer0_outputs(3769));
    layer1_outputs(6851) <= layer0_outputs(6726);
    layer1_outputs(6852) <= layer0_outputs(6303);
    layer1_outputs(6853) <= not(layer0_outputs(2969)) or (layer0_outputs(61));
    layer1_outputs(6854) <= '0';
    layer1_outputs(6855) <= layer0_outputs(743);
    layer1_outputs(6856) <= not(layer0_outputs(4005)) or (layer0_outputs(5058));
    layer1_outputs(6857) <= not(layer0_outputs(5018)) or (layer0_outputs(5592));
    layer1_outputs(6858) <= layer0_outputs(1191);
    layer1_outputs(6859) <= (layer0_outputs(7536)) xor (layer0_outputs(7383));
    layer1_outputs(6860) <= layer0_outputs(5292);
    layer1_outputs(6861) <= (layer0_outputs(2774)) and not (layer0_outputs(3053));
    layer1_outputs(6862) <= not((layer0_outputs(5300)) and (layer0_outputs(1002)));
    layer1_outputs(6863) <= not(layer0_outputs(2443));
    layer1_outputs(6864) <= '1';
    layer1_outputs(6865) <= layer0_outputs(2390);
    layer1_outputs(6866) <= not(layer0_outputs(3694));
    layer1_outputs(6867) <= not((layer0_outputs(232)) or (layer0_outputs(5886)));
    layer1_outputs(6868) <= not(layer0_outputs(1127));
    layer1_outputs(6869) <= not(layer0_outputs(3552)) or (layer0_outputs(7631));
    layer1_outputs(6870) <= layer0_outputs(1102);
    layer1_outputs(6871) <= not((layer0_outputs(2713)) or (layer0_outputs(4200)));
    layer1_outputs(6872) <= not(layer0_outputs(4865)) or (layer0_outputs(3055));
    layer1_outputs(6873) <= (layer0_outputs(2927)) and not (layer0_outputs(196));
    layer1_outputs(6874) <= not(layer0_outputs(4238));
    layer1_outputs(6875) <= not(layer0_outputs(5603));
    layer1_outputs(6876) <= '1';
    layer1_outputs(6877) <= (layer0_outputs(3634)) and not (layer0_outputs(1417));
    layer1_outputs(6878) <= layer0_outputs(3179);
    layer1_outputs(6879) <= not((layer0_outputs(2446)) xor (layer0_outputs(97)));
    layer1_outputs(6880) <= '0';
    layer1_outputs(6881) <= not(layer0_outputs(6294));
    layer1_outputs(6882) <= not(layer0_outputs(6508)) or (layer0_outputs(2419));
    layer1_outputs(6883) <= '1';
    layer1_outputs(6884) <= layer0_outputs(3888);
    layer1_outputs(6885) <= not(layer0_outputs(3881));
    layer1_outputs(6886) <= '0';
    layer1_outputs(6887) <= '1';
    layer1_outputs(6888) <= (layer0_outputs(6850)) and not (layer0_outputs(7));
    layer1_outputs(6889) <= (layer0_outputs(5419)) and not (layer0_outputs(5625));
    layer1_outputs(6890) <= layer0_outputs(6981);
    layer1_outputs(6891) <= (layer0_outputs(224)) and not (layer0_outputs(6976));
    layer1_outputs(6892) <= not((layer0_outputs(1509)) or (layer0_outputs(6059)));
    layer1_outputs(6893) <= not(layer0_outputs(2329)) or (layer0_outputs(1581));
    layer1_outputs(6894) <= layer0_outputs(3605);
    layer1_outputs(6895) <= '1';
    layer1_outputs(6896) <= (layer0_outputs(4425)) and not (layer0_outputs(6320));
    layer1_outputs(6897) <= not(layer0_outputs(492)) or (layer0_outputs(7678));
    layer1_outputs(6898) <= not((layer0_outputs(4402)) or (layer0_outputs(6385)));
    layer1_outputs(6899) <= not((layer0_outputs(3642)) or (layer0_outputs(4706)));
    layer1_outputs(6900) <= not(layer0_outputs(5680));
    layer1_outputs(6901) <= (layer0_outputs(2235)) and (layer0_outputs(5613));
    layer1_outputs(6902) <= (layer0_outputs(4134)) and (layer0_outputs(2966));
    layer1_outputs(6903) <= '0';
    layer1_outputs(6904) <= (layer0_outputs(1213)) and (layer0_outputs(5910));
    layer1_outputs(6905) <= layer0_outputs(5759);
    layer1_outputs(6906) <= '0';
    layer1_outputs(6907) <= (layer0_outputs(5286)) and not (layer0_outputs(3173));
    layer1_outputs(6908) <= '1';
    layer1_outputs(6909) <= '1';
    layer1_outputs(6910) <= '0';
    layer1_outputs(6911) <= '1';
    layer1_outputs(6912) <= '1';
    layer1_outputs(6913) <= not(layer0_outputs(1900));
    layer1_outputs(6914) <= '0';
    layer1_outputs(6915) <= layer0_outputs(5740);
    layer1_outputs(6916) <= (layer0_outputs(5694)) and not (layer0_outputs(4054));
    layer1_outputs(6917) <= (layer0_outputs(2830)) or (layer0_outputs(4885));
    layer1_outputs(6918) <= '0';
    layer1_outputs(6919) <= not((layer0_outputs(5138)) or (layer0_outputs(6546)));
    layer1_outputs(6920) <= layer0_outputs(5482);
    layer1_outputs(6921) <= not((layer0_outputs(5656)) and (layer0_outputs(5325)));
    layer1_outputs(6922) <= (layer0_outputs(5317)) and (layer0_outputs(3564));
    layer1_outputs(6923) <= layer0_outputs(2681);
    layer1_outputs(6924) <= (layer0_outputs(5629)) or (layer0_outputs(5374));
    layer1_outputs(6925) <= (layer0_outputs(4017)) or (layer0_outputs(5563));
    layer1_outputs(6926) <= layer0_outputs(6768);
    layer1_outputs(6927) <= '0';
    layer1_outputs(6928) <= layer0_outputs(7314);
    layer1_outputs(6929) <= not(layer0_outputs(1641)) or (layer0_outputs(3316));
    layer1_outputs(6930) <= (layer0_outputs(6123)) and not (layer0_outputs(256));
    layer1_outputs(6931) <= layer0_outputs(7440);
    layer1_outputs(6932) <= layer0_outputs(7143);
    layer1_outputs(6933) <= '1';
    layer1_outputs(6934) <= not(layer0_outputs(5004));
    layer1_outputs(6935) <= not((layer0_outputs(5790)) or (layer0_outputs(4602)));
    layer1_outputs(6936) <= '1';
    layer1_outputs(6937) <= not(layer0_outputs(2742));
    layer1_outputs(6938) <= layer0_outputs(6578);
    layer1_outputs(6939) <= not(layer0_outputs(3876)) or (layer0_outputs(7272));
    layer1_outputs(6940) <= layer0_outputs(3007);
    layer1_outputs(6941) <= (layer0_outputs(1179)) and (layer0_outputs(5750));
    layer1_outputs(6942) <= not((layer0_outputs(5809)) and (layer0_outputs(3759)));
    layer1_outputs(6943) <= (layer0_outputs(6873)) or (layer0_outputs(4968));
    layer1_outputs(6944) <= not(layer0_outputs(2133));
    layer1_outputs(6945) <= not((layer0_outputs(5354)) or (layer0_outputs(4059)));
    layer1_outputs(6946) <= layer0_outputs(3546);
    layer1_outputs(6947) <= '1';
    layer1_outputs(6948) <= not((layer0_outputs(1756)) or (layer0_outputs(1955)));
    layer1_outputs(6949) <= (layer0_outputs(4570)) and not (layer0_outputs(2168));
    layer1_outputs(6950) <= layer0_outputs(5039);
    layer1_outputs(6951) <= not(layer0_outputs(6086)) or (layer0_outputs(309));
    layer1_outputs(6952) <= (layer0_outputs(3835)) or (layer0_outputs(2788));
    layer1_outputs(6953) <= '1';
    layer1_outputs(6954) <= '0';
    layer1_outputs(6955) <= layer0_outputs(7424);
    layer1_outputs(6956) <= '1';
    layer1_outputs(6957) <= layer0_outputs(4330);
    layer1_outputs(6958) <= '0';
    layer1_outputs(6959) <= not((layer0_outputs(2161)) or (layer0_outputs(6006)));
    layer1_outputs(6960) <= not(layer0_outputs(3230)) or (layer0_outputs(4803));
    layer1_outputs(6961) <= not(layer0_outputs(5834));
    layer1_outputs(6962) <= not(layer0_outputs(4266));
    layer1_outputs(6963) <= layer0_outputs(7425);
    layer1_outputs(6964) <= not(layer0_outputs(1627)) or (layer0_outputs(3631));
    layer1_outputs(6965) <= not(layer0_outputs(7678)) or (layer0_outputs(1408));
    layer1_outputs(6966) <= (layer0_outputs(2291)) or (layer0_outputs(4225));
    layer1_outputs(6967) <= not(layer0_outputs(1167)) or (layer0_outputs(7615));
    layer1_outputs(6968) <= layer0_outputs(2812);
    layer1_outputs(6969) <= layer0_outputs(2545);
    layer1_outputs(6970) <= not((layer0_outputs(2798)) or (layer0_outputs(6888)));
    layer1_outputs(6971) <= not(layer0_outputs(6103));
    layer1_outputs(6972) <= layer0_outputs(1040);
    layer1_outputs(6973) <= not(layer0_outputs(2906)) or (layer0_outputs(4667));
    layer1_outputs(6974) <= not(layer0_outputs(1286)) or (layer0_outputs(3800));
    layer1_outputs(6975) <= not((layer0_outputs(4364)) and (layer0_outputs(7575)));
    layer1_outputs(6976) <= not((layer0_outputs(2153)) or (layer0_outputs(2250)));
    layer1_outputs(6977) <= (layer0_outputs(5355)) and (layer0_outputs(1603));
    layer1_outputs(6978) <= not((layer0_outputs(1813)) and (layer0_outputs(2201)));
    layer1_outputs(6979) <= (layer0_outputs(6417)) or (layer0_outputs(119));
    layer1_outputs(6980) <= (layer0_outputs(2436)) or (layer0_outputs(1363));
    layer1_outputs(6981) <= not(layer0_outputs(5559));
    layer1_outputs(6982) <= layer0_outputs(5382);
    layer1_outputs(6983) <= '1';
    layer1_outputs(6984) <= (layer0_outputs(2402)) and (layer0_outputs(6851));
    layer1_outputs(6985) <= layer0_outputs(103);
    layer1_outputs(6986) <= (layer0_outputs(3603)) and not (layer0_outputs(3868));
    layer1_outputs(6987) <= (layer0_outputs(40)) and (layer0_outputs(4758));
    layer1_outputs(6988) <= (layer0_outputs(369)) or (layer0_outputs(2659));
    layer1_outputs(6989) <= not((layer0_outputs(1710)) or (layer0_outputs(6776)));
    layer1_outputs(6990) <= not(layer0_outputs(729)) or (layer0_outputs(3858));
    layer1_outputs(6991) <= not(layer0_outputs(2053));
    layer1_outputs(6992) <= (layer0_outputs(7014)) and not (layer0_outputs(967));
    layer1_outputs(6993) <= layer0_outputs(5133);
    layer1_outputs(6994) <= not((layer0_outputs(4789)) and (layer0_outputs(4671)));
    layer1_outputs(6995) <= (layer0_outputs(2954)) and not (layer0_outputs(2785));
    layer1_outputs(6996) <= (layer0_outputs(73)) or (layer0_outputs(3204));
    layer1_outputs(6997) <= (layer0_outputs(530)) and not (layer0_outputs(6419));
    layer1_outputs(6998) <= '1';
    layer1_outputs(6999) <= '0';
    layer1_outputs(7000) <= not(layer0_outputs(1826));
    layer1_outputs(7001) <= '0';
    layer1_outputs(7002) <= (layer0_outputs(906)) and not (layer0_outputs(4657));
    layer1_outputs(7003) <= (layer0_outputs(2124)) and (layer0_outputs(2923));
    layer1_outputs(7004) <= not((layer0_outputs(5891)) or (layer0_outputs(2019)));
    layer1_outputs(7005) <= not(layer0_outputs(1458)) or (layer0_outputs(6441));
    layer1_outputs(7006) <= not(layer0_outputs(3167)) or (layer0_outputs(1838));
    layer1_outputs(7007) <= layer0_outputs(5332);
    layer1_outputs(7008) <= not(layer0_outputs(4550)) or (layer0_outputs(1306));
    layer1_outputs(7009) <= (layer0_outputs(5547)) and not (layer0_outputs(7648));
    layer1_outputs(7010) <= not(layer0_outputs(541)) or (layer0_outputs(5986));
    layer1_outputs(7011) <= layer0_outputs(1366);
    layer1_outputs(7012) <= not(layer0_outputs(3236)) or (layer0_outputs(3790));
    layer1_outputs(7013) <= not(layer0_outputs(2094));
    layer1_outputs(7014) <= (layer0_outputs(6987)) and not (layer0_outputs(6917));
    layer1_outputs(7015) <= '1';
    layer1_outputs(7016) <= not(layer0_outputs(6791));
    layer1_outputs(7017) <= '1';
    layer1_outputs(7018) <= (layer0_outputs(6354)) and not (layer0_outputs(1027));
    layer1_outputs(7019) <= not(layer0_outputs(4772));
    layer1_outputs(7020) <= not(layer0_outputs(1406)) or (layer0_outputs(6563));
    layer1_outputs(7021) <= '1';
    layer1_outputs(7022) <= not(layer0_outputs(6486));
    layer1_outputs(7023) <= (layer0_outputs(7496)) or (layer0_outputs(4863));
    layer1_outputs(7024) <= layer0_outputs(3842);
    layer1_outputs(7025) <= '1';
    layer1_outputs(7026) <= '1';
    layer1_outputs(7027) <= not(layer0_outputs(3448));
    layer1_outputs(7028) <= not(layer0_outputs(1802));
    layer1_outputs(7029) <= not(layer0_outputs(1766));
    layer1_outputs(7030) <= not((layer0_outputs(1796)) or (layer0_outputs(7333)));
    layer1_outputs(7031) <= '1';
    layer1_outputs(7032) <= not(layer0_outputs(3079)) or (layer0_outputs(6123));
    layer1_outputs(7033) <= not(layer0_outputs(4330));
    layer1_outputs(7034) <= not(layer0_outputs(828));
    layer1_outputs(7035) <= '0';
    layer1_outputs(7036) <= layer0_outputs(3368);
    layer1_outputs(7037) <= not((layer0_outputs(276)) xor (layer0_outputs(5166)));
    layer1_outputs(7038) <= layer0_outputs(3314);
    layer1_outputs(7039) <= '0';
    layer1_outputs(7040) <= (layer0_outputs(7200)) and not (layer0_outputs(4210));
    layer1_outputs(7041) <= not(layer0_outputs(748));
    layer1_outputs(7042) <= '1';
    layer1_outputs(7043) <= (layer0_outputs(1610)) and (layer0_outputs(3747));
    layer1_outputs(7044) <= '0';
    layer1_outputs(7045) <= (layer0_outputs(273)) or (layer0_outputs(4351));
    layer1_outputs(7046) <= (layer0_outputs(1381)) and not (layer0_outputs(734));
    layer1_outputs(7047) <= not((layer0_outputs(6991)) or (layer0_outputs(5103)));
    layer1_outputs(7048) <= (layer0_outputs(6567)) and (layer0_outputs(4918));
    layer1_outputs(7049) <= (layer0_outputs(2945)) or (layer0_outputs(6327));
    layer1_outputs(7050) <= (layer0_outputs(4482)) and not (layer0_outputs(3849));
    layer1_outputs(7051) <= layer0_outputs(2205);
    layer1_outputs(7052) <= not((layer0_outputs(4309)) xor (layer0_outputs(3745)));
    layer1_outputs(7053) <= layer0_outputs(5686);
    layer1_outputs(7054) <= layer0_outputs(941);
    layer1_outputs(7055) <= '0';
    layer1_outputs(7056) <= (layer0_outputs(209)) and not (layer0_outputs(3891));
    layer1_outputs(7057) <= (layer0_outputs(1294)) or (layer0_outputs(2070));
    layer1_outputs(7058) <= '1';
    layer1_outputs(7059) <= not(layer0_outputs(4004));
    layer1_outputs(7060) <= layer0_outputs(1926);
    layer1_outputs(7061) <= not((layer0_outputs(5788)) or (layer0_outputs(3128)));
    layer1_outputs(7062) <= (layer0_outputs(465)) or (layer0_outputs(3450));
    layer1_outputs(7063) <= '1';
    layer1_outputs(7064) <= not(layer0_outputs(7084)) or (layer0_outputs(481));
    layer1_outputs(7065) <= '1';
    layer1_outputs(7066) <= (layer0_outputs(6118)) and not (layer0_outputs(2702));
    layer1_outputs(7067) <= not(layer0_outputs(3165)) or (layer0_outputs(1030));
    layer1_outputs(7068) <= layer0_outputs(2777);
    layer1_outputs(7069) <= not(layer0_outputs(4922));
    layer1_outputs(7070) <= layer0_outputs(2546);
    layer1_outputs(7071) <= (layer0_outputs(1180)) xor (layer0_outputs(7441));
    layer1_outputs(7072) <= not((layer0_outputs(472)) and (layer0_outputs(1022)));
    layer1_outputs(7073) <= not((layer0_outputs(6897)) and (layer0_outputs(264)));
    layer1_outputs(7074) <= not(layer0_outputs(3483));
    layer1_outputs(7075) <= '0';
    layer1_outputs(7076) <= (layer0_outputs(640)) and not (layer0_outputs(6295));
    layer1_outputs(7077) <= not((layer0_outputs(1016)) and (layer0_outputs(188)));
    layer1_outputs(7078) <= (layer0_outputs(3734)) or (layer0_outputs(5327));
    layer1_outputs(7079) <= (layer0_outputs(6217)) or (layer0_outputs(1186));
    layer1_outputs(7080) <= (layer0_outputs(3892)) or (layer0_outputs(2592));
    layer1_outputs(7081) <= not((layer0_outputs(0)) and (layer0_outputs(6829)));
    layer1_outputs(7082) <= not((layer0_outputs(1762)) or (layer0_outputs(2445)));
    layer1_outputs(7083) <= not(layer0_outputs(866)) or (layer0_outputs(4338));
    layer1_outputs(7084) <= (layer0_outputs(412)) and not (layer0_outputs(4212));
    layer1_outputs(7085) <= not(layer0_outputs(752));
    layer1_outputs(7086) <= not((layer0_outputs(864)) or (layer0_outputs(3586)));
    layer1_outputs(7087) <= not(layer0_outputs(4591));
    layer1_outputs(7088) <= not(layer0_outputs(4249));
    layer1_outputs(7089) <= not(layer0_outputs(6801));
    layer1_outputs(7090) <= not(layer0_outputs(671)) or (layer0_outputs(6689));
    layer1_outputs(7091) <= '0';
    layer1_outputs(7092) <= not(layer0_outputs(237));
    layer1_outputs(7093) <= '1';
    layer1_outputs(7094) <= (layer0_outputs(7635)) and not (layer0_outputs(2717));
    layer1_outputs(7095) <= not((layer0_outputs(7121)) and (layer0_outputs(58)));
    layer1_outputs(7096) <= layer0_outputs(5596);
    layer1_outputs(7097) <= (layer0_outputs(5539)) and not (layer0_outputs(5855));
    layer1_outputs(7098) <= not(layer0_outputs(3851));
    layer1_outputs(7099) <= (layer0_outputs(7068)) and not (layer0_outputs(5175));
    layer1_outputs(7100) <= '1';
    layer1_outputs(7101) <= not((layer0_outputs(3049)) or (layer0_outputs(3865)));
    layer1_outputs(7102) <= '0';
    layer1_outputs(7103) <= (layer0_outputs(7348)) and not (layer0_outputs(6374));
    layer1_outputs(7104) <= layer0_outputs(2143);
    layer1_outputs(7105) <= (layer0_outputs(5639)) and (layer0_outputs(7491));
    layer1_outputs(7106) <= (layer0_outputs(1003)) and not (layer0_outputs(3944));
    layer1_outputs(7107) <= not((layer0_outputs(1148)) and (layer0_outputs(6490)));
    layer1_outputs(7108) <= not((layer0_outputs(6555)) or (layer0_outputs(7097)));
    layer1_outputs(7109) <= '0';
    layer1_outputs(7110) <= '0';
    layer1_outputs(7111) <= '0';
    layer1_outputs(7112) <= layer0_outputs(1144);
    layer1_outputs(7113) <= (layer0_outputs(3970)) and (layer0_outputs(6561));
    layer1_outputs(7114) <= not((layer0_outputs(1241)) and (layer0_outputs(219)));
    layer1_outputs(7115) <= (layer0_outputs(6493)) and (layer0_outputs(7601));
    layer1_outputs(7116) <= not((layer0_outputs(2667)) or (layer0_outputs(1769)));
    layer1_outputs(7117) <= not((layer0_outputs(4750)) or (layer0_outputs(3832)));
    layer1_outputs(7118) <= (layer0_outputs(5565)) and (layer0_outputs(3337));
    layer1_outputs(7119) <= layer0_outputs(7207);
    layer1_outputs(7120) <= layer0_outputs(130);
    layer1_outputs(7121) <= not((layer0_outputs(3140)) and (layer0_outputs(224)));
    layer1_outputs(7122) <= (layer0_outputs(831)) and not (layer0_outputs(204));
    layer1_outputs(7123) <= layer0_outputs(7074);
    layer1_outputs(7124) <= (layer0_outputs(7642)) and (layer0_outputs(6874));
    layer1_outputs(7125) <= layer0_outputs(1673);
    layer1_outputs(7126) <= not(layer0_outputs(6503));
    layer1_outputs(7127) <= not((layer0_outputs(5542)) and (layer0_outputs(2216)));
    layer1_outputs(7128) <= not(layer0_outputs(7645));
    layer1_outputs(7129) <= not((layer0_outputs(4081)) and (layer0_outputs(2268)));
    layer1_outputs(7130) <= not(layer0_outputs(6665));
    layer1_outputs(7131) <= layer0_outputs(5329);
    layer1_outputs(7132) <= not(layer0_outputs(3630)) or (layer0_outputs(104));
    layer1_outputs(7133) <= (layer0_outputs(6024)) or (layer0_outputs(5340));
    layer1_outputs(7134) <= (layer0_outputs(2589)) and not (layer0_outputs(6186));
    layer1_outputs(7135) <= '1';
    layer1_outputs(7136) <= not(layer0_outputs(2254)) or (layer0_outputs(3936));
    layer1_outputs(7137) <= layer0_outputs(4737);
    layer1_outputs(7138) <= (layer0_outputs(1431)) and (layer0_outputs(2560));
    layer1_outputs(7139) <= not(layer0_outputs(3062));
    layer1_outputs(7140) <= not(layer0_outputs(4020)) or (layer0_outputs(3967));
    layer1_outputs(7141) <= not(layer0_outputs(4904)) or (layer0_outputs(7194));
    layer1_outputs(7142) <= '1';
    layer1_outputs(7143) <= (layer0_outputs(5577)) and not (layer0_outputs(4690));
    layer1_outputs(7144) <= not(layer0_outputs(3221));
    layer1_outputs(7145) <= '0';
    layer1_outputs(7146) <= layer0_outputs(1599);
    layer1_outputs(7147) <= layer0_outputs(5200);
    layer1_outputs(7148) <= '1';
    layer1_outputs(7149) <= not(layer0_outputs(3746));
    layer1_outputs(7150) <= (layer0_outputs(3614)) and not (layer0_outputs(1695));
    layer1_outputs(7151) <= layer0_outputs(3340);
    layer1_outputs(7152) <= (layer0_outputs(784)) and not (layer0_outputs(787));
    layer1_outputs(7153) <= not(layer0_outputs(7299)) or (layer0_outputs(5532));
    layer1_outputs(7154) <= not((layer0_outputs(4050)) xor (layer0_outputs(1413)));
    layer1_outputs(7155) <= layer0_outputs(4923);
    layer1_outputs(7156) <= not(layer0_outputs(2606));
    layer1_outputs(7157) <= not(layer0_outputs(5511));
    layer1_outputs(7158) <= (layer0_outputs(7051)) and not (layer0_outputs(609));
    layer1_outputs(7159) <= not(layer0_outputs(94));
    layer1_outputs(7160) <= (layer0_outputs(4272)) and (layer0_outputs(5719));
    layer1_outputs(7161) <= layer0_outputs(1719);
    layer1_outputs(7162) <= '1';
    layer1_outputs(7163) <= layer0_outputs(5955);
    layer1_outputs(7164) <= (layer0_outputs(3996)) and (layer0_outputs(6207));
    layer1_outputs(7165) <= not((layer0_outputs(853)) and (layer0_outputs(7511)));
    layer1_outputs(7166) <= '0';
    layer1_outputs(7167) <= not(layer0_outputs(5595)) or (layer0_outputs(7528));
    layer1_outputs(7168) <= (layer0_outputs(3951)) and not (layer0_outputs(3502));
    layer1_outputs(7169) <= not(layer0_outputs(31));
    layer1_outputs(7170) <= (layer0_outputs(3177)) or (layer0_outputs(1622));
    layer1_outputs(7171) <= not(layer0_outputs(6335)) or (layer0_outputs(3001));
    layer1_outputs(7172) <= (layer0_outputs(2674)) or (layer0_outputs(1211));
    layer1_outputs(7173) <= not(layer0_outputs(6343));
    layer1_outputs(7174) <= not(layer0_outputs(443)) or (layer0_outputs(3084));
    layer1_outputs(7175) <= '0';
    layer1_outputs(7176) <= layer0_outputs(2697);
    layer1_outputs(7177) <= layer0_outputs(4768);
    layer1_outputs(7178) <= layer0_outputs(1862);
    layer1_outputs(7179) <= layer0_outputs(698);
    layer1_outputs(7180) <= layer0_outputs(7622);
    layer1_outputs(7181) <= layer0_outputs(1035);
    layer1_outputs(7182) <= '0';
    layer1_outputs(7183) <= (layer0_outputs(979)) or (layer0_outputs(2826));
    layer1_outputs(7184) <= '0';
    layer1_outputs(7185) <= (layer0_outputs(289)) xor (layer0_outputs(5172));
    layer1_outputs(7186) <= not(layer0_outputs(4316));
    layer1_outputs(7187) <= layer0_outputs(3070);
    layer1_outputs(7188) <= not(layer0_outputs(2703));
    layer1_outputs(7189) <= (layer0_outputs(6378)) and not (layer0_outputs(1651));
    layer1_outputs(7190) <= (layer0_outputs(7443)) and not (layer0_outputs(7410));
    layer1_outputs(7191) <= not(layer0_outputs(3201));
    layer1_outputs(7192) <= layer0_outputs(871);
    layer1_outputs(7193) <= (layer0_outputs(2723)) xor (layer0_outputs(1493));
    layer1_outputs(7194) <= not(layer0_outputs(7234)) or (layer0_outputs(1923));
    layer1_outputs(7195) <= (layer0_outputs(5992)) or (layer0_outputs(2864));
    layer1_outputs(7196) <= (layer0_outputs(756)) and not (layer0_outputs(7452));
    layer1_outputs(7197) <= not(layer0_outputs(719)) or (layer0_outputs(1373));
    layer1_outputs(7198) <= not((layer0_outputs(3777)) xor (layer0_outputs(7557)));
    layer1_outputs(7199) <= '1';
    layer1_outputs(7200) <= layer0_outputs(1905);
    layer1_outputs(7201) <= not(layer0_outputs(2213)) or (layer0_outputs(4627));
    layer1_outputs(7202) <= (layer0_outputs(6236)) or (layer0_outputs(7289));
    layer1_outputs(7203) <= (layer0_outputs(5931)) and not (layer0_outputs(4196));
    layer1_outputs(7204) <= not((layer0_outputs(6838)) and (layer0_outputs(6387)));
    layer1_outputs(7205) <= layer0_outputs(842);
    layer1_outputs(7206) <= not(layer0_outputs(557));
    layer1_outputs(7207) <= not((layer0_outputs(1078)) or (layer0_outputs(896)));
    layer1_outputs(7208) <= not(layer0_outputs(1602));
    layer1_outputs(7209) <= layer0_outputs(6400);
    layer1_outputs(7210) <= not((layer0_outputs(5735)) and (layer0_outputs(5020)));
    layer1_outputs(7211) <= not(layer0_outputs(6505)) or (layer0_outputs(5064));
    layer1_outputs(7212) <= not((layer0_outputs(7311)) or (layer0_outputs(4107)));
    layer1_outputs(7213) <= not(layer0_outputs(871));
    layer1_outputs(7214) <= not((layer0_outputs(4660)) or (layer0_outputs(1785)));
    layer1_outputs(7215) <= (layer0_outputs(2010)) or (layer0_outputs(3371));
    layer1_outputs(7216) <= not(layer0_outputs(1896));
    layer1_outputs(7217) <= not(layer0_outputs(5824)) or (layer0_outputs(407));
    layer1_outputs(7218) <= not((layer0_outputs(6410)) or (layer0_outputs(3057)));
    layer1_outputs(7219) <= '0';
    layer1_outputs(7220) <= not(layer0_outputs(6619));
    layer1_outputs(7221) <= (layer0_outputs(6218)) and (layer0_outputs(1917));
    layer1_outputs(7222) <= not((layer0_outputs(1195)) and (layer0_outputs(4664)));
    layer1_outputs(7223) <= '1';
    layer1_outputs(7224) <= not(layer0_outputs(2301)) or (layer0_outputs(235));
    layer1_outputs(7225) <= (layer0_outputs(7234)) and not (layer0_outputs(7311));
    layer1_outputs(7226) <= (layer0_outputs(3833)) or (layer0_outputs(5907));
    layer1_outputs(7227) <= not(layer0_outputs(5315));
    layer1_outputs(7228) <= (layer0_outputs(494)) xor (layer0_outputs(2511));
    layer1_outputs(7229) <= '0';
    layer1_outputs(7230) <= not(layer0_outputs(149));
    layer1_outputs(7231) <= layer0_outputs(4844);
    layer1_outputs(7232) <= '1';
    layer1_outputs(7233) <= not((layer0_outputs(3135)) xor (layer0_outputs(4451)));
    layer1_outputs(7234) <= '1';
    layer1_outputs(7235) <= not(layer0_outputs(5123));
    layer1_outputs(7236) <= not(layer0_outputs(5730));
    layer1_outputs(7237) <= '0';
    layer1_outputs(7238) <= not((layer0_outputs(3569)) or (layer0_outputs(6064)));
    layer1_outputs(7239) <= (layer0_outputs(6845)) and not (layer0_outputs(6759));
    layer1_outputs(7240) <= (layer0_outputs(7472)) and (layer0_outputs(5240));
    layer1_outputs(7241) <= not((layer0_outputs(1913)) or (layer0_outputs(2039)));
    layer1_outputs(7242) <= layer0_outputs(3099);
    layer1_outputs(7243) <= (layer0_outputs(7479)) xor (layer0_outputs(6437));
    layer1_outputs(7244) <= '0';
    layer1_outputs(7245) <= layer0_outputs(7187);
    layer1_outputs(7246) <= not(layer0_outputs(434)) or (layer0_outputs(5961));
    layer1_outputs(7247) <= not(layer0_outputs(5496)) or (layer0_outputs(463));
    layer1_outputs(7248) <= not((layer0_outputs(2122)) or (layer0_outputs(1474)));
    layer1_outputs(7249) <= layer0_outputs(1407);
    layer1_outputs(7250) <= '0';
    layer1_outputs(7251) <= not(layer0_outputs(3137));
    layer1_outputs(7252) <= (layer0_outputs(1389)) and not (layer0_outputs(1842));
    layer1_outputs(7253) <= not(layer0_outputs(6089));
    layer1_outputs(7254) <= layer0_outputs(4253);
    layer1_outputs(7255) <= (layer0_outputs(1217)) and (layer0_outputs(5745));
    layer1_outputs(7256) <= not(layer0_outputs(7177)) or (layer0_outputs(5697));
    layer1_outputs(7257) <= (layer0_outputs(366)) and not (layer0_outputs(5807));
    layer1_outputs(7258) <= '1';
    layer1_outputs(7259) <= '1';
    layer1_outputs(7260) <= not(layer0_outputs(5134)) or (layer0_outputs(2972));
    layer1_outputs(7261) <= not(layer0_outputs(6434));
    layer1_outputs(7262) <= (layer0_outputs(2080)) and not (layer0_outputs(5660));
    layer1_outputs(7263) <= '0';
    layer1_outputs(7264) <= (layer0_outputs(4414)) or (layer0_outputs(402));
    layer1_outputs(7265) <= (layer0_outputs(7075)) and not (layer0_outputs(93));
    layer1_outputs(7266) <= (layer0_outputs(1377)) or (layer0_outputs(5681));
    layer1_outputs(7267) <= (layer0_outputs(4753)) and not (layer0_outputs(6969));
    layer1_outputs(7268) <= layer0_outputs(4528);
    layer1_outputs(7269) <= (layer0_outputs(7420)) or (layer0_outputs(4739));
    layer1_outputs(7270) <= not(layer0_outputs(4731)) or (layer0_outputs(6596));
    layer1_outputs(7271) <= layer0_outputs(5878);
    layer1_outputs(7272) <= (layer0_outputs(6982)) and not (layer0_outputs(2895));
    layer1_outputs(7273) <= not(layer0_outputs(6381)) or (layer0_outputs(6789));
    layer1_outputs(7274) <= (layer0_outputs(6516)) and not (layer0_outputs(1094));
    layer1_outputs(7275) <= not((layer0_outputs(4932)) or (layer0_outputs(3347)));
    layer1_outputs(7276) <= not((layer0_outputs(6878)) and (layer0_outputs(4546)));
    layer1_outputs(7277) <= (layer0_outputs(121)) or (layer0_outputs(7085));
    layer1_outputs(7278) <= (layer0_outputs(2721)) and not (layer0_outputs(3346));
    layer1_outputs(7279) <= (layer0_outputs(5734)) and not (layer0_outputs(5377));
    layer1_outputs(7280) <= not((layer0_outputs(5757)) or (layer0_outputs(30)));
    layer1_outputs(7281) <= '0';
    layer1_outputs(7282) <= (layer0_outputs(1360)) and not (layer0_outputs(6484));
    layer1_outputs(7283) <= '1';
    layer1_outputs(7284) <= (layer0_outputs(7144)) and not (layer0_outputs(445));
    layer1_outputs(7285) <= not(layer0_outputs(4676)) or (layer0_outputs(5211));
    layer1_outputs(7286) <= (layer0_outputs(1380)) and (layer0_outputs(3675));
    layer1_outputs(7287) <= not((layer0_outputs(853)) or (layer0_outputs(4910)));
    layer1_outputs(7288) <= '1';
    layer1_outputs(7289) <= not(layer0_outputs(813)) or (layer0_outputs(3243));
    layer1_outputs(7290) <= (layer0_outputs(5725)) and not (layer0_outputs(7000));
    layer1_outputs(7291) <= not((layer0_outputs(2771)) and (layer0_outputs(760)));
    layer1_outputs(7292) <= '1';
    layer1_outputs(7293) <= not(layer0_outputs(120));
    layer1_outputs(7294) <= (layer0_outputs(4770)) and not (layer0_outputs(5967));
    layer1_outputs(7295) <= (layer0_outputs(2901)) and not (layer0_outputs(564));
    layer1_outputs(7296) <= not((layer0_outputs(6353)) xor (layer0_outputs(4010)));
    layer1_outputs(7297) <= '1';
    layer1_outputs(7298) <= not((layer0_outputs(5296)) and (layer0_outputs(790)));
    layer1_outputs(7299) <= (layer0_outputs(7435)) or (layer0_outputs(2635));
    layer1_outputs(7300) <= not(layer0_outputs(921));
    layer1_outputs(7301) <= layer0_outputs(7219);
    layer1_outputs(7302) <= layer0_outputs(6379);
    layer1_outputs(7303) <= not(layer0_outputs(2560));
    layer1_outputs(7304) <= not(layer0_outputs(6763));
    layer1_outputs(7305) <= not(layer0_outputs(6904));
    layer1_outputs(7306) <= '1';
    layer1_outputs(7307) <= (layer0_outputs(5470)) and (layer0_outputs(7025));
    layer1_outputs(7308) <= (layer0_outputs(6453)) and (layer0_outputs(5270));
    layer1_outputs(7309) <= not(layer0_outputs(6884)) or (layer0_outputs(1993));
    layer1_outputs(7310) <= (layer0_outputs(586)) and (layer0_outputs(4867));
    layer1_outputs(7311) <= (layer0_outputs(5954)) and not (layer0_outputs(3903));
    layer1_outputs(7312) <= not((layer0_outputs(1070)) and (layer0_outputs(112)));
    layer1_outputs(7313) <= not(layer0_outputs(6185)) or (layer0_outputs(6880));
    layer1_outputs(7314) <= (layer0_outputs(7138)) and not (layer0_outputs(985));
    layer1_outputs(7315) <= not(layer0_outputs(5023)) or (layer0_outputs(1506));
    layer1_outputs(7316) <= '1';
    layer1_outputs(7317) <= not(layer0_outputs(4500)) or (layer0_outputs(3232));
    layer1_outputs(7318) <= layer0_outputs(4681);
    layer1_outputs(7319) <= (layer0_outputs(3118)) and not (layer0_outputs(1532));
    layer1_outputs(7320) <= not(layer0_outputs(3732));
    layer1_outputs(7321) <= not((layer0_outputs(4447)) and (layer0_outputs(6843)));
    layer1_outputs(7322) <= (layer0_outputs(1477)) or (layer0_outputs(3297));
    layer1_outputs(7323) <= not((layer0_outputs(1301)) or (layer0_outputs(4866)));
    layer1_outputs(7324) <= not((layer0_outputs(5700)) or (layer0_outputs(6809)));
    layer1_outputs(7325) <= not(layer0_outputs(4373)) or (layer0_outputs(1995));
    layer1_outputs(7326) <= '0';
    layer1_outputs(7327) <= '1';
    layer1_outputs(7328) <= '0';
    layer1_outputs(7329) <= not(layer0_outputs(1043));
    layer1_outputs(7330) <= (layer0_outputs(1702)) and not (layer0_outputs(6265));
    layer1_outputs(7331) <= '0';
    layer1_outputs(7332) <= (layer0_outputs(7335)) and (layer0_outputs(5851));
    layer1_outputs(7333) <= not(layer0_outputs(271)) or (layer0_outputs(1547));
    layer1_outputs(7334) <= (layer0_outputs(3973)) and not (layer0_outputs(1589));
    layer1_outputs(7335) <= not(layer0_outputs(6865));
    layer1_outputs(7336) <= not((layer0_outputs(3762)) or (layer0_outputs(4747)));
    layer1_outputs(7337) <= '0';
    layer1_outputs(7338) <= not(layer0_outputs(1844));
    layer1_outputs(7339) <= not((layer0_outputs(4597)) or (layer0_outputs(4908)));
    layer1_outputs(7340) <= not(layer0_outputs(6331));
    layer1_outputs(7341) <= (layer0_outputs(5202)) or (layer0_outputs(3409));
    layer1_outputs(7342) <= (layer0_outputs(2407)) and (layer0_outputs(6030));
    layer1_outputs(7343) <= (layer0_outputs(2899)) or (layer0_outputs(5400));
    layer1_outputs(7344) <= (layer0_outputs(3231)) and (layer0_outputs(4994));
    layer1_outputs(7345) <= not(layer0_outputs(2388)) or (layer0_outputs(3129));
    layer1_outputs(7346) <= not(layer0_outputs(5793)) or (layer0_outputs(502));
    layer1_outputs(7347) <= (layer0_outputs(6729)) and not (layer0_outputs(2874));
    layer1_outputs(7348) <= (layer0_outputs(185)) and not (layer0_outputs(223));
    layer1_outputs(7349) <= not(layer0_outputs(371)) or (layer0_outputs(1683));
    layer1_outputs(7350) <= (layer0_outputs(2258)) and (layer0_outputs(533));
    layer1_outputs(7351) <= '1';
    layer1_outputs(7352) <= '1';
    layer1_outputs(7353) <= (layer0_outputs(5586)) and not (layer0_outputs(4246));
    layer1_outputs(7354) <= not((layer0_outputs(1273)) or (layer0_outputs(917)));
    layer1_outputs(7355) <= layer0_outputs(6158);
    layer1_outputs(7356) <= layer0_outputs(7098);
    layer1_outputs(7357) <= not(layer0_outputs(4439)) or (layer0_outputs(570));
    layer1_outputs(7358) <= (layer0_outputs(6670)) and not (layer0_outputs(7073));
    layer1_outputs(7359) <= (layer0_outputs(4545)) and not (layer0_outputs(5856));
    layer1_outputs(7360) <= (layer0_outputs(7386)) and (layer0_outputs(6155));
    layer1_outputs(7361) <= '0';
    layer1_outputs(7362) <= not(layer0_outputs(3346));
    layer1_outputs(7363) <= '1';
    layer1_outputs(7364) <= (layer0_outputs(4261)) and (layer0_outputs(1314));
    layer1_outputs(7365) <= not(layer0_outputs(4285));
    layer1_outputs(7366) <= not(layer0_outputs(7040));
    layer1_outputs(7367) <= not(layer0_outputs(4520));
    layer1_outputs(7368) <= not(layer0_outputs(6512)) or (layer0_outputs(7439));
    layer1_outputs(7369) <= '0';
    layer1_outputs(7370) <= '0';
    layer1_outputs(7371) <= layer0_outputs(3295);
    layer1_outputs(7372) <= '1';
    layer1_outputs(7373) <= not((layer0_outputs(4230)) or (layer0_outputs(4491)));
    layer1_outputs(7374) <= not(layer0_outputs(5174)) or (layer0_outputs(1027));
    layer1_outputs(7375) <= not(layer0_outputs(1088));
    layer1_outputs(7376) <= (layer0_outputs(1401)) and not (layer0_outputs(4724));
    layer1_outputs(7377) <= not(layer0_outputs(2320));
    layer1_outputs(7378) <= (layer0_outputs(2651)) or (layer0_outputs(2726));
    layer1_outputs(7379) <= (layer0_outputs(6399)) and not (layer0_outputs(3521));
    layer1_outputs(7380) <= not(layer0_outputs(212)) or (layer0_outputs(3185));
    layer1_outputs(7381) <= (layer0_outputs(1075)) or (layer0_outputs(3659));
    layer1_outputs(7382) <= not(layer0_outputs(1748)) or (layer0_outputs(1476));
    layer1_outputs(7383) <= not(layer0_outputs(548));
    layer1_outputs(7384) <= not(layer0_outputs(4223)) or (layer0_outputs(2942));
    layer1_outputs(7385) <= not(layer0_outputs(4435)) or (layer0_outputs(7187));
    layer1_outputs(7386) <= not((layer0_outputs(7412)) xor (layer0_outputs(4668)));
    layer1_outputs(7387) <= '1';
    layer1_outputs(7388) <= '0';
    layer1_outputs(7389) <= (layer0_outputs(1339)) or (layer0_outputs(3721));
    layer1_outputs(7390) <= not(layer0_outputs(1847)) or (layer0_outputs(5767));
    layer1_outputs(7391) <= (layer0_outputs(881)) and not (layer0_outputs(2435));
    layer1_outputs(7392) <= (layer0_outputs(1218)) or (layer0_outputs(6770));
    layer1_outputs(7393) <= (layer0_outputs(3879)) and (layer0_outputs(2725));
    layer1_outputs(7394) <= not(layer0_outputs(1270));
    layer1_outputs(7395) <= not(layer0_outputs(3637));
    layer1_outputs(7396) <= '0';
    layer1_outputs(7397) <= not((layer0_outputs(2634)) and (layer0_outputs(2212)));
    layer1_outputs(7398) <= not((layer0_outputs(3522)) or (layer0_outputs(1595)));
    layer1_outputs(7399) <= not(layer0_outputs(479)) or (layer0_outputs(4790));
    layer1_outputs(7400) <= (layer0_outputs(580)) and not (layer0_outputs(888));
    layer1_outputs(7401) <= layer0_outputs(6823);
    layer1_outputs(7402) <= '0';
    layer1_outputs(7403) <= not(layer0_outputs(5337));
    layer1_outputs(7404) <= (layer0_outputs(5467)) xor (layer0_outputs(4022));
    layer1_outputs(7405) <= not(layer0_outputs(7368));
    layer1_outputs(7406) <= not((layer0_outputs(6893)) or (layer0_outputs(1184)));
    layer1_outputs(7407) <= layer0_outputs(5287);
    layer1_outputs(7408) <= layer0_outputs(288);
    layer1_outputs(7409) <= not(layer0_outputs(3572));
    layer1_outputs(7410) <= (layer0_outputs(7654)) and not (layer0_outputs(256));
    layer1_outputs(7411) <= layer0_outputs(6348);
    layer1_outputs(7412) <= not(layer0_outputs(4524));
    layer1_outputs(7413) <= not((layer0_outputs(6018)) and (layer0_outputs(6618)));
    layer1_outputs(7414) <= layer0_outputs(1721);
    layer1_outputs(7415) <= (layer0_outputs(4180)) and not (layer0_outputs(5072));
    layer1_outputs(7416) <= layer0_outputs(2671);
    layer1_outputs(7417) <= '0';
    layer1_outputs(7418) <= (layer0_outputs(782)) and not (layer0_outputs(5793));
    layer1_outputs(7419) <= (layer0_outputs(1642)) and (layer0_outputs(1670));
    layer1_outputs(7420) <= layer0_outputs(3566);
    layer1_outputs(7421) <= not((layer0_outputs(4325)) or (layer0_outputs(2622)));
    layer1_outputs(7422) <= not((layer0_outputs(1553)) or (layer0_outputs(914)));
    layer1_outputs(7423) <= (layer0_outputs(5210)) and (layer0_outputs(267));
    layer1_outputs(7424) <= (layer0_outputs(6013)) or (layer0_outputs(7190));
    layer1_outputs(7425) <= not(layer0_outputs(1239)) or (layer0_outputs(3442));
    layer1_outputs(7426) <= '0';
    layer1_outputs(7427) <= '0';
    layer1_outputs(7428) <= not(layer0_outputs(6535));
    layer1_outputs(7429) <= (layer0_outputs(6326)) or (layer0_outputs(3252));
    layer1_outputs(7430) <= not((layer0_outputs(667)) and (layer0_outputs(1072)));
    layer1_outputs(7431) <= (layer0_outputs(1042)) and (layer0_outputs(998));
    layer1_outputs(7432) <= layer0_outputs(1551);
    layer1_outputs(7433) <= not(layer0_outputs(1199));
    layer1_outputs(7434) <= (layer0_outputs(3341)) and (layer0_outputs(3922));
    layer1_outputs(7435) <= '1';
    layer1_outputs(7436) <= '0';
    layer1_outputs(7437) <= '0';
    layer1_outputs(7438) <= '0';
    layer1_outputs(7439) <= not((layer0_outputs(4310)) or (layer0_outputs(6008)));
    layer1_outputs(7440) <= (layer0_outputs(4118)) or (layer0_outputs(6289));
    layer1_outputs(7441) <= '1';
    layer1_outputs(7442) <= (layer0_outputs(2573)) and not (layer0_outputs(419));
    layer1_outputs(7443) <= layer0_outputs(6175);
    layer1_outputs(7444) <= '0';
    layer1_outputs(7445) <= not(layer0_outputs(1362)) or (layer0_outputs(350));
    layer1_outputs(7446) <= (layer0_outputs(3689)) and not (layer0_outputs(705));
    layer1_outputs(7447) <= layer0_outputs(6108);
    layer1_outputs(7448) <= layer0_outputs(6646);
    layer1_outputs(7449) <= (layer0_outputs(6081)) and not (layer0_outputs(2412));
    layer1_outputs(7450) <= not(layer0_outputs(4027));
    layer1_outputs(7451) <= '0';
    layer1_outputs(7452) <= (layer0_outputs(634)) and (layer0_outputs(1438));
    layer1_outputs(7453) <= (layer0_outputs(3535)) and (layer0_outputs(2584));
    layer1_outputs(7454) <= (layer0_outputs(614)) xor (layer0_outputs(1842));
    layer1_outputs(7455) <= not((layer0_outputs(626)) xor (layer0_outputs(461)));
    layer1_outputs(7456) <= not(layer0_outputs(765)) or (layer0_outputs(730));
    layer1_outputs(7457) <= '1';
    layer1_outputs(7458) <= layer0_outputs(5159);
    layer1_outputs(7459) <= not((layer0_outputs(3257)) or (layer0_outputs(161)));
    layer1_outputs(7460) <= not((layer0_outputs(572)) and (layer0_outputs(1529)));
    layer1_outputs(7461) <= '1';
    layer1_outputs(7462) <= layer0_outputs(6303);
    layer1_outputs(7463) <= not(layer0_outputs(6829));
    layer1_outputs(7464) <= (layer0_outputs(7279)) and (layer0_outputs(6965));
    layer1_outputs(7465) <= (layer0_outputs(7403)) and not (layer0_outputs(3228));
    layer1_outputs(7466) <= not(layer0_outputs(918)) or (layer0_outputs(7037));
    layer1_outputs(7467) <= layer0_outputs(4548);
    layer1_outputs(7468) <= layer0_outputs(303);
    layer1_outputs(7469) <= (layer0_outputs(1822)) and not (layer0_outputs(2710));
    layer1_outputs(7470) <= layer0_outputs(3439);
    layer1_outputs(7471) <= layer0_outputs(3386);
    layer1_outputs(7472) <= '1';
    layer1_outputs(7473) <= (layer0_outputs(3489)) and (layer0_outputs(780));
    layer1_outputs(7474) <= (layer0_outputs(51)) and not (layer0_outputs(4040));
    layer1_outputs(7475) <= layer0_outputs(4352);
    layer1_outputs(7476) <= not(layer0_outputs(6438)) or (layer0_outputs(2246));
    layer1_outputs(7477) <= layer0_outputs(1232);
    layer1_outputs(7478) <= (layer0_outputs(6119)) and not (layer0_outputs(5765));
    layer1_outputs(7479) <= layer0_outputs(79);
    layer1_outputs(7480) <= not(layer0_outputs(2282));
    layer1_outputs(7481) <= not(layer0_outputs(861));
    layer1_outputs(7482) <= '1';
    layer1_outputs(7483) <= (layer0_outputs(6985)) xor (layer0_outputs(3048));
    layer1_outputs(7484) <= '0';
    layer1_outputs(7485) <= '0';
    layer1_outputs(7486) <= layer0_outputs(7555);
    layer1_outputs(7487) <= '0';
    layer1_outputs(7488) <= (layer0_outputs(2518)) and (layer0_outputs(5045));
    layer1_outputs(7489) <= not(layer0_outputs(4515));
    layer1_outputs(7490) <= layer0_outputs(6567);
    layer1_outputs(7491) <= (layer0_outputs(5341)) and not (layer0_outputs(6521));
    layer1_outputs(7492) <= not(layer0_outputs(1066)) or (layer0_outputs(1095));
    layer1_outputs(7493) <= '0';
    layer1_outputs(7494) <= not(layer0_outputs(7432)) or (layer0_outputs(4480));
    layer1_outputs(7495) <= layer0_outputs(5523);
    layer1_outputs(7496) <= layer0_outputs(7310);
    layer1_outputs(7497) <= (layer0_outputs(689)) or (layer0_outputs(1133));
    layer1_outputs(7498) <= '1';
    layer1_outputs(7499) <= '0';
    layer1_outputs(7500) <= (layer0_outputs(7260)) or (layer0_outputs(7539));
    layer1_outputs(7501) <= (layer0_outputs(964)) and (layer0_outputs(3964));
    layer1_outputs(7502) <= not(layer0_outputs(3774));
    layer1_outputs(7503) <= layer0_outputs(1034);
    layer1_outputs(7504) <= (layer0_outputs(3146)) and (layer0_outputs(3042));
    layer1_outputs(7505) <= not(layer0_outputs(5310));
    layer1_outputs(7506) <= not(layer0_outputs(225));
    layer1_outputs(7507) <= not((layer0_outputs(3513)) xor (layer0_outputs(215)));
    layer1_outputs(7508) <= '1';
    layer1_outputs(7509) <= layer0_outputs(3416);
    layer1_outputs(7510) <= (layer0_outputs(6027)) and not (layer0_outputs(5914));
    layer1_outputs(7511) <= layer0_outputs(5241);
    layer1_outputs(7512) <= not(layer0_outputs(7394));
    layer1_outputs(7513) <= (layer0_outputs(910)) xor (layer0_outputs(3063));
    layer1_outputs(7514) <= not(layer0_outputs(2843));
    layer1_outputs(7515) <= not((layer0_outputs(5626)) or (layer0_outputs(4073)));
    layer1_outputs(7516) <= '1';
    layer1_outputs(7517) <= '1';
    layer1_outputs(7518) <= not((layer0_outputs(73)) xor (layer0_outputs(4452)));
    layer1_outputs(7519) <= layer0_outputs(3294);
    layer1_outputs(7520) <= '1';
    layer1_outputs(7521) <= not(layer0_outputs(1746));
    layer1_outputs(7522) <= '0';
    layer1_outputs(7523) <= not(layer0_outputs(2138));
    layer1_outputs(7524) <= (layer0_outputs(948)) and not (layer0_outputs(1694));
    layer1_outputs(7525) <= (layer0_outputs(2436)) and (layer0_outputs(7586));
    layer1_outputs(7526) <= not(layer0_outputs(6880));
    layer1_outputs(7527) <= not((layer0_outputs(5925)) and (layer0_outputs(4103)));
    layer1_outputs(7528) <= not(layer0_outputs(2977)) or (layer0_outputs(4832));
    layer1_outputs(7529) <= not(layer0_outputs(6696));
    layer1_outputs(7530) <= (layer0_outputs(777)) or (layer0_outputs(2896));
    layer1_outputs(7531) <= not(layer0_outputs(1867));
    layer1_outputs(7532) <= (layer0_outputs(3732)) and (layer0_outputs(3222));
    layer1_outputs(7533) <= (layer0_outputs(628)) or (layer0_outputs(863));
    layer1_outputs(7534) <= (layer0_outputs(2621)) and not (layer0_outputs(208));
    layer1_outputs(7535) <= (layer0_outputs(435)) and not (layer0_outputs(6445));
    layer1_outputs(7536) <= '1';
    layer1_outputs(7537) <= not((layer0_outputs(6611)) and (layer0_outputs(6915)));
    layer1_outputs(7538) <= layer0_outputs(1739);
    layer1_outputs(7539) <= (layer0_outputs(1023)) xor (layer0_outputs(4639));
    layer1_outputs(7540) <= layer0_outputs(3168);
    layer1_outputs(7541) <= '0';
    layer1_outputs(7542) <= '0';
    layer1_outputs(7543) <= layer0_outputs(6066);
    layer1_outputs(7544) <= (layer0_outputs(6825)) and not (layer0_outputs(1390));
    layer1_outputs(7545) <= not((layer0_outputs(1468)) or (layer0_outputs(1428)));
    layer1_outputs(7546) <= not(layer0_outputs(5477));
    layer1_outputs(7547) <= not(layer0_outputs(2414)) or (layer0_outputs(5752));
    layer1_outputs(7548) <= layer0_outputs(4111);
    layer1_outputs(7549) <= not(layer0_outputs(2242)) or (layer0_outputs(1719));
    layer1_outputs(7550) <= (layer0_outputs(6905)) and (layer0_outputs(6537));
    layer1_outputs(7551) <= not(layer0_outputs(5638)) or (layer0_outputs(2608));
    layer1_outputs(7552) <= layer0_outputs(7032);
    layer1_outputs(7553) <= '0';
    layer1_outputs(7554) <= (layer0_outputs(6498)) or (layer0_outputs(3544));
    layer1_outputs(7555) <= not(layer0_outputs(7296)) or (layer0_outputs(1754));
    layer1_outputs(7556) <= (layer0_outputs(1485)) or (layer0_outputs(3575));
    layer1_outputs(7557) <= '0';
    layer1_outputs(7558) <= (layer0_outputs(6966)) and not (layer0_outputs(283));
    layer1_outputs(7559) <= (layer0_outputs(2342)) and not (layer0_outputs(7001));
    layer1_outputs(7560) <= (layer0_outputs(1109)) and not (layer0_outputs(4316));
    layer1_outputs(7561) <= not(layer0_outputs(3179));
    layer1_outputs(7562) <= not(layer0_outputs(1907));
    layer1_outputs(7563) <= '0';
    layer1_outputs(7564) <= '0';
    layer1_outputs(7565) <= '1';
    layer1_outputs(7566) <= '0';
    layer1_outputs(7567) <= not(layer0_outputs(4281)) or (layer0_outputs(6766));
    layer1_outputs(7568) <= layer0_outputs(5185);
    layer1_outputs(7569) <= (layer0_outputs(7633)) and not (layer0_outputs(177));
    layer1_outputs(7570) <= not(layer0_outputs(3842));
    layer1_outputs(7571) <= not(layer0_outputs(2333));
    layer1_outputs(7572) <= (layer0_outputs(7624)) and not (layer0_outputs(6882));
    layer1_outputs(7573) <= (layer0_outputs(4226)) xor (layer0_outputs(447));
    layer1_outputs(7574) <= layer0_outputs(1163);
    layer1_outputs(7575) <= not(layer0_outputs(5529)) or (layer0_outputs(5053));
    layer1_outputs(7576) <= (layer0_outputs(5472)) or (layer0_outputs(6643));
    layer1_outputs(7577) <= not((layer0_outputs(3237)) or (layer0_outputs(3273)));
    layer1_outputs(7578) <= not(layer0_outputs(5908));
    layer1_outputs(7579) <= layer0_outputs(4537);
    layer1_outputs(7580) <= not(layer0_outputs(1744));
    layer1_outputs(7581) <= layer0_outputs(2752);
    layer1_outputs(7582) <= not((layer0_outputs(129)) or (layer0_outputs(5237)));
    layer1_outputs(7583) <= not((layer0_outputs(7142)) and (layer0_outputs(1758)));
    layer1_outputs(7584) <= not(layer0_outputs(2472)) or (layer0_outputs(7340));
    layer1_outputs(7585) <= not(layer0_outputs(5144));
    layer1_outputs(7586) <= not(layer0_outputs(2834)) or (layer0_outputs(914));
    layer1_outputs(7587) <= layer0_outputs(4232);
    layer1_outputs(7588) <= (layer0_outputs(6953)) or (layer0_outputs(7617));
    layer1_outputs(7589) <= '1';
    layer1_outputs(7590) <= (layer0_outputs(5061)) and not (layer0_outputs(3463));
    layer1_outputs(7591) <= (layer0_outputs(7600)) and not (layer0_outputs(2032));
    layer1_outputs(7592) <= (layer0_outputs(4228)) xor (layer0_outputs(7233));
    layer1_outputs(7593) <= '0';
    layer1_outputs(7594) <= not(layer0_outputs(911));
    layer1_outputs(7595) <= not(layer0_outputs(1881)) or (layer0_outputs(7103));
    layer1_outputs(7596) <= not(layer0_outputs(3431));
    layer1_outputs(7597) <= (layer0_outputs(3016)) and not (layer0_outputs(6463));
    layer1_outputs(7598) <= not((layer0_outputs(4027)) and (layer0_outputs(2971)));
    layer1_outputs(7599) <= layer0_outputs(6828);
    layer1_outputs(7600) <= '1';
    layer1_outputs(7601) <= not(layer0_outputs(808));
    layer1_outputs(7602) <= (layer0_outputs(2627)) and not (layer0_outputs(902));
    layer1_outputs(7603) <= not(layer0_outputs(6690));
    layer1_outputs(7604) <= not(layer0_outputs(5171));
    layer1_outputs(7605) <= not(layer0_outputs(5312));
    layer1_outputs(7606) <= layer0_outputs(2288);
    layer1_outputs(7607) <= layer0_outputs(6110);
    layer1_outputs(7608) <= (layer0_outputs(4293)) and (layer0_outputs(1692));
    layer1_outputs(7609) <= not(layer0_outputs(632));
    layer1_outputs(7610) <= '1';
    layer1_outputs(7611) <= not(layer0_outputs(4034)) or (layer0_outputs(5067));
    layer1_outputs(7612) <= layer0_outputs(4670);
    layer1_outputs(7613) <= (layer0_outputs(6411)) and not (layer0_outputs(2113));
    layer1_outputs(7614) <= '0';
    layer1_outputs(7615) <= layer0_outputs(1213);
    layer1_outputs(7616) <= (layer0_outputs(1380)) and not (layer0_outputs(6750));
    layer1_outputs(7617) <= not((layer0_outputs(1308)) or (layer0_outputs(2754)));
    layer1_outputs(7618) <= '1';
    layer1_outputs(7619) <= not(layer0_outputs(1112));
    layer1_outputs(7620) <= not(layer0_outputs(2620));
    layer1_outputs(7621) <= not(layer0_outputs(6787));
    layer1_outputs(7622) <= not(layer0_outputs(2331));
    layer1_outputs(7623) <= not(layer0_outputs(4760));
    layer1_outputs(7624) <= not(layer0_outputs(4177)) or (layer0_outputs(5983));
    layer1_outputs(7625) <= not((layer0_outputs(5344)) or (layer0_outputs(2831)));
    layer1_outputs(7626) <= not((layer0_outputs(2967)) or (layer0_outputs(4492)));
    layer1_outputs(7627) <= not(layer0_outputs(1901)) or (layer0_outputs(328));
    layer1_outputs(7628) <= not((layer0_outputs(7182)) or (layer0_outputs(2152)));
    layer1_outputs(7629) <= (layer0_outputs(2936)) and (layer0_outputs(4344));
    layer1_outputs(7630) <= not((layer0_outputs(3905)) and (layer0_outputs(201)));
    layer1_outputs(7631) <= (layer0_outputs(1260)) and not (layer0_outputs(3460));
    layer1_outputs(7632) <= not(layer0_outputs(4992));
    layer1_outputs(7633) <= '1';
    layer1_outputs(7634) <= not(layer0_outputs(569));
    layer1_outputs(7635) <= '1';
    layer1_outputs(7636) <= (layer0_outputs(3729)) and not (layer0_outputs(6442));
    layer1_outputs(7637) <= (layer0_outputs(3098)) and not (layer0_outputs(1472));
    layer1_outputs(7638) <= not(layer0_outputs(1962));
    layer1_outputs(7639) <= '0';
    layer1_outputs(7640) <= (layer0_outputs(7111)) xor (layer0_outputs(5326));
    layer1_outputs(7641) <= '1';
    layer1_outputs(7642) <= not((layer0_outputs(600)) or (layer0_outputs(4199)));
    layer1_outputs(7643) <= not(layer0_outputs(4876)) or (layer0_outputs(7016));
    layer1_outputs(7644) <= '0';
    layer1_outputs(7645) <= not(layer0_outputs(5570)) or (layer0_outputs(1832));
    layer1_outputs(7646) <= (layer0_outputs(1084)) and not (layer0_outputs(6935));
    layer1_outputs(7647) <= (layer0_outputs(3246)) and (layer0_outputs(7268));
    layer1_outputs(7648) <= layer0_outputs(4760);
    layer1_outputs(7649) <= layer0_outputs(1135);
    layer1_outputs(7650) <= (layer0_outputs(3649)) and not (layer0_outputs(3727));
    layer1_outputs(7651) <= '1';
    layer1_outputs(7652) <= (layer0_outputs(5286)) or (layer0_outputs(2785));
    layer1_outputs(7653) <= (layer0_outputs(1217)) and not (layer0_outputs(5167));
    layer1_outputs(7654) <= (layer0_outputs(5587)) and not (layer0_outputs(3501));
    layer1_outputs(7655) <= layer0_outputs(1041);
    layer1_outputs(7656) <= layer0_outputs(5671);
    layer1_outputs(7657) <= not((layer0_outputs(3280)) and (layer0_outputs(6093)));
    layer1_outputs(7658) <= not((layer0_outputs(3224)) and (layer0_outputs(6465)));
    layer1_outputs(7659) <= '0';
    layer1_outputs(7660) <= (layer0_outputs(2794)) and (layer0_outputs(6406));
    layer1_outputs(7661) <= layer0_outputs(3636);
    layer1_outputs(7662) <= '1';
    layer1_outputs(7663) <= not((layer0_outputs(6841)) and (layer0_outputs(2116)));
    layer1_outputs(7664) <= layer0_outputs(536);
    layer1_outputs(7665) <= not(layer0_outputs(672));
    layer1_outputs(7666) <= layer0_outputs(7380);
    layer1_outputs(7667) <= '1';
    layer1_outputs(7668) <= (layer0_outputs(778)) and not (layer0_outputs(3829));
    layer1_outputs(7669) <= (layer0_outputs(6288)) or (layer0_outputs(6617));
    layer1_outputs(7670) <= not(layer0_outputs(5524));
    layer1_outputs(7671) <= not((layer0_outputs(6228)) and (layer0_outputs(927)));
    layer1_outputs(7672) <= not((layer0_outputs(3310)) and (layer0_outputs(1307)));
    layer1_outputs(7673) <= not(layer0_outputs(2297));
    layer1_outputs(7674) <= (layer0_outputs(4795)) or (layer0_outputs(5448));
    layer1_outputs(7675) <= not((layer0_outputs(4862)) and (layer0_outputs(2214)));
    layer1_outputs(7676) <= (layer0_outputs(1107)) and not (layer0_outputs(6071));
    layer1_outputs(7677) <= not(layer0_outputs(2448));
    layer1_outputs(7678) <= '0';
    layer1_outputs(7679) <= layer0_outputs(1790);
    layer2_outputs(0) <= '0';
    layer2_outputs(1) <= layer1_outputs(3162);
    layer2_outputs(2) <= not(layer1_outputs(6972)) or (layer1_outputs(2105));
    layer2_outputs(3) <= layer1_outputs(4106);
    layer2_outputs(4) <= (layer1_outputs(5655)) xor (layer1_outputs(1952));
    layer2_outputs(5) <= layer1_outputs(3186);
    layer2_outputs(6) <= layer1_outputs(3672);
    layer2_outputs(7) <= (layer1_outputs(7445)) and not (layer1_outputs(7657));
    layer2_outputs(8) <= (layer1_outputs(885)) and not (layer1_outputs(6628));
    layer2_outputs(9) <= not(layer1_outputs(1995));
    layer2_outputs(10) <= not((layer1_outputs(2011)) and (layer1_outputs(1036)));
    layer2_outputs(11) <= not(layer1_outputs(6045));
    layer2_outputs(12) <= '1';
    layer2_outputs(13) <= not(layer1_outputs(4016)) or (layer1_outputs(6225));
    layer2_outputs(14) <= layer1_outputs(1669);
    layer2_outputs(15) <= not(layer1_outputs(240)) or (layer1_outputs(6386));
    layer2_outputs(16) <= not(layer1_outputs(6475));
    layer2_outputs(17) <= not((layer1_outputs(7044)) and (layer1_outputs(472)));
    layer2_outputs(18) <= not((layer1_outputs(1965)) or (layer1_outputs(943)));
    layer2_outputs(19) <= not(layer1_outputs(5618));
    layer2_outputs(20) <= not(layer1_outputs(5172));
    layer2_outputs(21) <= not(layer1_outputs(5979));
    layer2_outputs(22) <= not((layer1_outputs(3529)) and (layer1_outputs(2952)));
    layer2_outputs(23) <= not(layer1_outputs(847)) or (layer1_outputs(4917));
    layer2_outputs(24) <= layer1_outputs(4209);
    layer2_outputs(25) <= not(layer1_outputs(1565)) or (layer1_outputs(489));
    layer2_outputs(26) <= not((layer1_outputs(3287)) or (layer1_outputs(2487)));
    layer2_outputs(27) <= layer1_outputs(609);
    layer2_outputs(28) <= (layer1_outputs(7419)) and not (layer1_outputs(5855));
    layer2_outputs(29) <= not((layer1_outputs(6751)) or (layer1_outputs(4160)));
    layer2_outputs(30) <= layer1_outputs(3804);
    layer2_outputs(31) <= '0';
    layer2_outputs(32) <= not(layer1_outputs(7007));
    layer2_outputs(33) <= (layer1_outputs(1102)) and not (layer1_outputs(7150));
    layer2_outputs(34) <= '0';
    layer2_outputs(35) <= not(layer1_outputs(1093));
    layer2_outputs(36) <= not((layer1_outputs(6440)) or (layer1_outputs(5447)));
    layer2_outputs(37) <= '0';
    layer2_outputs(38) <= (layer1_outputs(1384)) or (layer1_outputs(6725));
    layer2_outputs(39) <= '0';
    layer2_outputs(40) <= not(layer1_outputs(1288));
    layer2_outputs(41) <= not(layer1_outputs(4554));
    layer2_outputs(42) <= (layer1_outputs(5167)) or (layer1_outputs(758));
    layer2_outputs(43) <= not(layer1_outputs(4196));
    layer2_outputs(44) <= not(layer1_outputs(5587)) or (layer1_outputs(3879));
    layer2_outputs(45) <= not(layer1_outputs(232)) or (layer1_outputs(4002));
    layer2_outputs(46) <= (layer1_outputs(106)) and (layer1_outputs(2857));
    layer2_outputs(47) <= layer1_outputs(2167);
    layer2_outputs(48) <= not(layer1_outputs(3315)) or (layer1_outputs(3557));
    layer2_outputs(49) <= not(layer1_outputs(3251));
    layer2_outputs(50) <= (layer1_outputs(2969)) or (layer1_outputs(1244));
    layer2_outputs(51) <= (layer1_outputs(423)) or (layer1_outputs(7421));
    layer2_outputs(52) <= layer1_outputs(5855);
    layer2_outputs(53) <= not(layer1_outputs(7333)) or (layer1_outputs(3246));
    layer2_outputs(54) <= '1';
    layer2_outputs(55) <= not(layer1_outputs(5605)) or (layer1_outputs(5899));
    layer2_outputs(56) <= layer1_outputs(999);
    layer2_outputs(57) <= not((layer1_outputs(189)) or (layer1_outputs(5829)));
    layer2_outputs(58) <= not(layer1_outputs(6543));
    layer2_outputs(59) <= not(layer1_outputs(1960)) or (layer1_outputs(1553));
    layer2_outputs(60) <= not(layer1_outputs(6176));
    layer2_outputs(61) <= '0';
    layer2_outputs(62) <= layer1_outputs(6022);
    layer2_outputs(63) <= (layer1_outputs(651)) and not (layer1_outputs(6236));
    layer2_outputs(64) <= (layer1_outputs(998)) and not (layer1_outputs(6544));
    layer2_outputs(65) <= not((layer1_outputs(866)) or (layer1_outputs(214)));
    layer2_outputs(66) <= layer1_outputs(3501);
    layer2_outputs(67) <= layer1_outputs(6670);
    layer2_outputs(68) <= not((layer1_outputs(6970)) or (layer1_outputs(242)));
    layer2_outputs(69) <= (layer1_outputs(4249)) and (layer1_outputs(7021));
    layer2_outputs(70) <= layer1_outputs(7051);
    layer2_outputs(71) <= (layer1_outputs(4967)) and (layer1_outputs(7471));
    layer2_outputs(72) <= (layer1_outputs(3259)) and not (layer1_outputs(1323));
    layer2_outputs(73) <= not(layer1_outputs(5970)) or (layer1_outputs(6551));
    layer2_outputs(74) <= not(layer1_outputs(1368)) or (layer1_outputs(4323));
    layer2_outputs(75) <= not(layer1_outputs(3008));
    layer2_outputs(76) <= not(layer1_outputs(3121)) or (layer1_outputs(3075));
    layer2_outputs(77) <= '0';
    layer2_outputs(78) <= not((layer1_outputs(1398)) and (layer1_outputs(2311)));
    layer2_outputs(79) <= (layer1_outputs(2315)) and not (layer1_outputs(4250));
    layer2_outputs(80) <= not(layer1_outputs(2710)) or (layer1_outputs(3536));
    layer2_outputs(81) <= (layer1_outputs(6554)) and not (layer1_outputs(7027));
    layer2_outputs(82) <= not(layer1_outputs(1143)) or (layer1_outputs(5372));
    layer2_outputs(83) <= '0';
    layer2_outputs(84) <= not((layer1_outputs(3700)) xor (layer1_outputs(1508)));
    layer2_outputs(85) <= (layer1_outputs(5999)) or (layer1_outputs(1988));
    layer2_outputs(86) <= not(layer1_outputs(1049)) or (layer1_outputs(6335));
    layer2_outputs(87) <= (layer1_outputs(3650)) and not (layer1_outputs(4014));
    layer2_outputs(88) <= (layer1_outputs(2843)) and not (layer1_outputs(2097));
    layer2_outputs(89) <= not((layer1_outputs(4913)) or (layer1_outputs(3264)));
    layer2_outputs(90) <= not(layer1_outputs(5039)) or (layer1_outputs(2486));
    layer2_outputs(91) <= not(layer1_outputs(1297)) or (layer1_outputs(807));
    layer2_outputs(92) <= (layer1_outputs(5563)) or (layer1_outputs(2540));
    layer2_outputs(93) <= not(layer1_outputs(2693));
    layer2_outputs(94) <= (layer1_outputs(7424)) and not (layer1_outputs(1840));
    layer2_outputs(95) <= not((layer1_outputs(6894)) and (layer1_outputs(4328)));
    layer2_outputs(96) <= not(layer1_outputs(5946)) or (layer1_outputs(412));
    layer2_outputs(97) <= '0';
    layer2_outputs(98) <= '1';
    layer2_outputs(99) <= not((layer1_outputs(2)) or (layer1_outputs(3858)));
    layer2_outputs(100) <= (layer1_outputs(7259)) or (layer1_outputs(1222));
    layer2_outputs(101) <= (layer1_outputs(2427)) or (layer1_outputs(5290));
    layer2_outputs(102) <= not(layer1_outputs(1205));
    layer2_outputs(103) <= (layer1_outputs(216)) and (layer1_outputs(5746));
    layer2_outputs(104) <= not((layer1_outputs(4679)) and (layer1_outputs(4641)));
    layer2_outputs(105) <= not(layer1_outputs(3692));
    layer2_outputs(106) <= not(layer1_outputs(4546)) or (layer1_outputs(4517));
    layer2_outputs(107) <= (layer1_outputs(5757)) and (layer1_outputs(6270));
    layer2_outputs(108) <= not(layer1_outputs(4175));
    layer2_outputs(109) <= '0';
    layer2_outputs(110) <= not(layer1_outputs(5801));
    layer2_outputs(111) <= not((layer1_outputs(7389)) and (layer1_outputs(5970)));
    layer2_outputs(112) <= not(layer1_outputs(3166)) or (layer1_outputs(7136));
    layer2_outputs(113) <= not(layer1_outputs(5072));
    layer2_outputs(114) <= not(layer1_outputs(1383));
    layer2_outputs(115) <= not((layer1_outputs(2866)) and (layer1_outputs(6318)));
    layer2_outputs(116) <= (layer1_outputs(6864)) and not (layer1_outputs(1685));
    layer2_outputs(117) <= not((layer1_outputs(312)) or (layer1_outputs(764)));
    layer2_outputs(118) <= (layer1_outputs(5266)) and not (layer1_outputs(678));
    layer2_outputs(119) <= not(layer1_outputs(5407));
    layer2_outputs(120) <= not(layer1_outputs(1924));
    layer2_outputs(121) <= layer1_outputs(6450);
    layer2_outputs(122) <= not((layer1_outputs(7064)) or (layer1_outputs(2136)));
    layer2_outputs(123) <= not((layer1_outputs(3993)) and (layer1_outputs(3507)));
    layer2_outputs(124) <= not((layer1_outputs(7066)) and (layer1_outputs(7151)));
    layer2_outputs(125) <= '0';
    layer2_outputs(126) <= layer1_outputs(6995);
    layer2_outputs(127) <= '0';
    layer2_outputs(128) <= (layer1_outputs(4776)) and not (layer1_outputs(4821));
    layer2_outputs(129) <= layer1_outputs(2119);
    layer2_outputs(130) <= not(layer1_outputs(3990)) or (layer1_outputs(6282));
    layer2_outputs(131) <= not(layer1_outputs(244));
    layer2_outputs(132) <= (layer1_outputs(2129)) or (layer1_outputs(3577));
    layer2_outputs(133) <= not(layer1_outputs(6635)) or (layer1_outputs(92));
    layer2_outputs(134) <= layer1_outputs(5640);
    layer2_outputs(135) <= '0';
    layer2_outputs(136) <= layer1_outputs(3893);
    layer2_outputs(137) <= '1';
    layer2_outputs(138) <= not(layer1_outputs(1138));
    layer2_outputs(139) <= '1';
    layer2_outputs(140) <= (layer1_outputs(7056)) or (layer1_outputs(905));
    layer2_outputs(141) <= not(layer1_outputs(1963)) or (layer1_outputs(2522));
    layer2_outputs(142) <= '0';
    layer2_outputs(143) <= layer1_outputs(6742);
    layer2_outputs(144) <= '1';
    layer2_outputs(145) <= not((layer1_outputs(7247)) and (layer1_outputs(6522)));
    layer2_outputs(146) <= not(layer1_outputs(342));
    layer2_outputs(147) <= (layer1_outputs(4105)) and not (layer1_outputs(4376));
    layer2_outputs(148) <= '1';
    layer2_outputs(149) <= (layer1_outputs(4577)) and not (layer1_outputs(6826));
    layer2_outputs(150) <= layer1_outputs(5971);
    layer2_outputs(151) <= (layer1_outputs(2076)) and not (layer1_outputs(5615));
    layer2_outputs(152) <= (layer1_outputs(3899)) or (layer1_outputs(130));
    layer2_outputs(153) <= not(layer1_outputs(1682));
    layer2_outputs(154) <= (layer1_outputs(6190)) or (layer1_outputs(5461));
    layer2_outputs(155) <= layer1_outputs(2660);
    layer2_outputs(156) <= (layer1_outputs(2382)) and (layer1_outputs(7402));
    layer2_outputs(157) <= layer1_outputs(1979);
    layer2_outputs(158) <= not(layer1_outputs(4303));
    layer2_outputs(159) <= (layer1_outputs(5469)) and not (layer1_outputs(2904));
    layer2_outputs(160) <= (layer1_outputs(3364)) xor (layer1_outputs(1328));
    layer2_outputs(161) <= layer1_outputs(4284);
    layer2_outputs(162) <= (layer1_outputs(5396)) or (layer1_outputs(6375));
    layer2_outputs(163) <= not(layer1_outputs(4518)) or (layer1_outputs(7543));
    layer2_outputs(164) <= layer1_outputs(1306);
    layer2_outputs(165) <= layer1_outputs(5999);
    layer2_outputs(166) <= (layer1_outputs(2713)) or (layer1_outputs(3137));
    layer2_outputs(167) <= layer1_outputs(3379);
    layer2_outputs(168) <= layer1_outputs(2434);
    layer2_outputs(169) <= not((layer1_outputs(1097)) or (layer1_outputs(1160)));
    layer2_outputs(170) <= not(layer1_outputs(7207));
    layer2_outputs(171) <= (layer1_outputs(4477)) and not (layer1_outputs(2757));
    layer2_outputs(172) <= '0';
    layer2_outputs(173) <= not(layer1_outputs(1142));
    layer2_outputs(174) <= not((layer1_outputs(7526)) and (layer1_outputs(5328)));
    layer2_outputs(175) <= layer1_outputs(3730);
    layer2_outputs(176) <= '0';
    layer2_outputs(177) <= not((layer1_outputs(492)) and (layer1_outputs(5915)));
    layer2_outputs(178) <= not(layer1_outputs(3615));
    layer2_outputs(179) <= not(layer1_outputs(7103));
    layer2_outputs(180) <= layer1_outputs(576);
    layer2_outputs(181) <= not(layer1_outputs(1733)) or (layer1_outputs(3078));
    layer2_outputs(182) <= (layer1_outputs(6710)) and (layer1_outputs(2296));
    layer2_outputs(183) <= not((layer1_outputs(2039)) and (layer1_outputs(4690)));
    layer2_outputs(184) <= not((layer1_outputs(6460)) and (layer1_outputs(3651)));
    layer2_outputs(185) <= '0';
    layer2_outputs(186) <= layer1_outputs(1266);
    layer2_outputs(187) <= not((layer1_outputs(4590)) xor (layer1_outputs(5167)));
    layer2_outputs(188) <= not((layer1_outputs(1517)) and (layer1_outputs(4360)));
    layer2_outputs(189) <= not(layer1_outputs(1470));
    layer2_outputs(190) <= not(layer1_outputs(4242));
    layer2_outputs(191) <= '1';
    layer2_outputs(192) <= (layer1_outputs(6752)) and not (layer1_outputs(1236));
    layer2_outputs(193) <= not(layer1_outputs(7511));
    layer2_outputs(194) <= not((layer1_outputs(5346)) or (layer1_outputs(3210)));
    layer2_outputs(195) <= (layer1_outputs(4937)) and not (layer1_outputs(6874));
    layer2_outputs(196) <= (layer1_outputs(4667)) and not (layer1_outputs(544));
    layer2_outputs(197) <= not(layer1_outputs(2037));
    layer2_outputs(198) <= layer1_outputs(306);
    layer2_outputs(199) <= not(layer1_outputs(2015));
    layer2_outputs(200) <= '0';
    layer2_outputs(201) <= '0';
    layer2_outputs(202) <= not(layer1_outputs(4190));
    layer2_outputs(203) <= (layer1_outputs(7146)) xor (layer1_outputs(5914));
    layer2_outputs(204) <= (layer1_outputs(2708)) and not (layer1_outputs(3513));
    layer2_outputs(205) <= not((layer1_outputs(4435)) or (layer1_outputs(3978)));
    layer2_outputs(206) <= '1';
    layer2_outputs(207) <= (layer1_outputs(1349)) and (layer1_outputs(219));
    layer2_outputs(208) <= (layer1_outputs(7019)) and (layer1_outputs(6289));
    layer2_outputs(209) <= (layer1_outputs(5202)) xor (layer1_outputs(312));
    layer2_outputs(210) <= not(layer1_outputs(5535)) or (layer1_outputs(6517));
    layer2_outputs(211) <= not(layer1_outputs(2477));
    layer2_outputs(212) <= not((layer1_outputs(2531)) and (layer1_outputs(1283)));
    layer2_outputs(213) <= not(layer1_outputs(5716));
    layer2_outputs(214) <= '0';
    layer2_outputs(215) <= not(layer1_outputs(6766)) or (layer1_outputs(3497));
    layer2_outputs(216) <= not((layer1_outputs(1473)) and (layer1_outputs(462)));
    layer2_outputs(217) <= not((layer1_outputs(1094)) and (layer1_outputs(2630)));
    layer2_outputs(218) <= not(layer1_outputs(7220));
    layer2_outputs(219) <= not(layer1_outputs(5154));
    layer2_outputs(220) <= (layer1_outputs(6352)) and not (layer1_outputs(6556));
    layer2_outputs(221) <= (layer1_outputs(5474)) and (layer1_outputs(1847));
    layer2_outputs(222) <= '0';
    layer2_outputs(223) <= '0';
    layer2_outputs(224) <= not((layer1_outputs(1087)) and (layer1_outputs(3366)));
    layer2_outputs(225) <= layer1_outputs(5764);
    layer2_outputs(226) <= (layer1_outputs(1780)) and not (layer1_outputs(1321));
    layer2_outputs(227) <= (layer1_outputs(5752)) and not (layer1_outputs(1165));
    layer2_outputs(228) <= not(layer1_outputs(2477));
    layer2_outputs(229) <= not((layer1_outputs(4641)) and (layer1_outputs(51)));
    layer2_outputs(230) <= layer1_outputs(2873);
    layer2_outputs(231) <= not(layer1_outputs(5285)) or (layer1_outputs(7439));
    layer2_outputs(232) <= not(layer1_outputs(4887)) or (layer1_outputs(4101));
    layer2_outputs(233) <= not(layer1_outputs(5238)) or (layer1_outputs(3995));
    layer2_outputs(234) <= '0';
    layer2_outputs(235) <= not((layer1_outputs(6368)) or (layer1_outputs(7467)));
    layer2_outputs(236) <= (layer1_outputs(1846)) or (layer1_outputs(3752));
    layer2_outputs(237) <= not(layer1_outputs(3727)) or (layer1_outputs(2886));
    layer2_outputs(238) <= (layer1_outputs(5486)) xor (layer1_outputs(2367));
    layer2_outputs(239) <= not(layer1_outputs(4111)) or (layer1_outputs(1537));
    layer2_outputs(240) <= not(layer1_outputs(5695));
    layer2_outputs(241) <= not(layer1_outputs(737));
    layer2_outputs(242) <= not(layer1_outputs(4940)) or (layer1_outputs(2560));
    layer2_outputs(243) <= not(layer1_outputs(1141)) or (layer1_outputs(1132));
    layer2_outputs(244) <= '0';
    layer2_outputs(245) <= '0';
    layer2_outputs(246) <= not((layer1_outputs(7000)) and (layer1_outputs(3468)));
    layer2_outputs(247) <= (layer1_outputs(5512)) and (layer1_outputs(3741));
    layer2_outputs(248) <= not(layer1_outputs(393));
    layer2_outputs(249) <= not((layer1_outputs(3858)) and (layer1_outputs(5800)));
    layer2_outputs(250) <= '0';
    layer2_outputs(251) <= not(layer1_outputs(1850)) or (layer1_outputs(4896));
    layer2_outputs(252) <= '0';
    layer2_outputs(253) <= not(layer1_outputs(6039));
    layer2_outputs(254) <= not(layer1_outputs(6160));
    layer2_outputs(255) <= layer1_outputs(1967);
    layer2_outputs(256) <= not(layer1_outputs(719));
    layer2_outputs(257) <= '0';
    layer2_outputs(258) <= '0';
    layer2_outputs(259) <= not(layer1_outputs(2605)) or (layer1_outputs(4301));
    layer2_outputs(260) <= (layer1_outputs(1783)) xor (layer1_outputs(4638));
    layer2_outputs(261) <= layer1_outputs(2602);
    layer2_outputs(262) <= layer1_outputs(3617);
    layer2_outputs(263) <= not(layer1_outputs(4320)) or (layer1_outputs(5320));
    layer2_outputs(264) <= not(layer1_outputs(4387));
    layer2_outputs(265) <= not(layer1_outputs(5770));
    layer2_outputs(266) <= (layer1_outputs(6575)) and not (layer1_outputs(1829));
    layer2_outputs(267) <= (layer1_outputs(993)) and not (layer1_outputs(4519));
    layer2_outputs(268) <= (layer1_outputs(6510)) or (layer1_outputs(1182));
    layer2_outputs(269) <= not((layer1_outputs(606)) and (layer1_outputs(4018)));
    layer2_outputs(270) <= not(layer1_outputs(2079));
    layer2_outputs(271) <= '1';
    layer2_outputs(272) <= not(layer1_outputs(7343));
    layer2_outputs(273) <= layer1_outputs(3177);
    layer2_outputs(274) <= (layer1_outputs(7112)) and not (layer1_outputs(2208));
    layer2_outputs(275) <= not((layer1_outputs(2692)) or (layer1_outputs(6372)));
    layer2_outputs(276) <= not(layer1_outputs(6410));
    layer2_outputs(277) <= (layer1_outputs(352)) or (layer1_outputs(5798));
    layer2_outputs(278) <= not((layer1_outputs(4501)) or (layer1_outputs(977)));
    layer2_outputs(279) <= (layer1_outputs(2601)) and not (layer1_outputs(3827));
    layer2_outputs(280) <= layer1_outputs(5054);
    layer2_outputs(281) <= not((layer1_outputs(6690)) and (layer1_outputs(2805)));
    layer2_outputs(282) <= not(layer1_outputs(789)) or (layer1_outputs(4614));
    layer2_outputs(283) <= '0';
    layer2_outputs(284) <= layer1_outputs(2592);
    layer2_outputs(285) <= not(layer1_outputs(2406));
    layer2_outputs(286) <= (layer1_outputs(2418)) and not (layer1_outputs(4203));
    layer2_outputs(287) <= '0';
    layer2_outputs(288) <= layer1_outputs(4595);
    layer2_outputs(289) <= not(layer1_outputs(5714));
    layer2_outputs(290) <= not(layer1_outputs(1065));
    layer2_outputs(291) <= (layer1_outputs(2501)) and not (layer1_outputs(2515));
    layer2_outputs(292) <= not((layer1_outputs(4759)) or (layer1_outputs(2824)));
    layer2_outputs(293) <= not((layer1_outputs(3840)) and (layer1_outputs(7437)));
    layer2_outputs(294) <= '1';
    layer2_outputs(295) <= not(layer1_outputs(4273));
    layer2_outputs(296) <= layer1_outputs(3739);
    layer2_outputs(297) <= layer1_outputs(3663);
    layer2_outputs(298) <= '0';
    layer2_outputs(299) <= not(layer1_outputs(6700)) or (layer1_outputs(3704));
    layer2_outputs(300) <= not((layer1_outputs(5788)) or (layer1_outputs(3671)));
    layer2_outputs(301) <= '0';
    layer2_outputs(302) <= '1';
    layer2_outputs(303) <= '0';
    layer2_outputs(304) <= not(layer1_outputs(286));
    layer2_outputs(305) <= not(layer1_outputs(5822));
    layer2_outputs(306) <= not((layer1_outputs(5233)) and (layer1_outputs(206)));
    layer2_outputs(307) <= '0';
    layer2_outputs(308) <= (layer1_outputs(5010)) and not (layer1_outputs(7648));
    layer2_outputs(309) <= layer1_outputs(846);
    layer2_outputs(310) <= (layer1_outputs(4686)) and (layer1_outputs(3545));
    layer2_outputs(311) <= layer1_outputs(2889);
    layer2_outputs(312) <= not(layer1_outputs(6507)) or (layer1_outputs(2840));
    layer2_outputs(313) <= layer1_outputs(2719);
    layer2_outputs(314) <= layer1_outputs(4356);
    layer2_outputs(315) <= layer1_outputs(76);
    layer2_outputs(316) <= (layer1_outputs(6115)) or (layer1_outputs(5109));
    layer2_outputs(317) <= '0';
    layer2_outputs(318) <= (layer1_outputs(2543)) or (layer1_outputs(1631));
    layer2_outputs(319) <= layer1_outputs(5152);
    layer2_outputs(320) <= layer1_outputs(7459);
    layer2_outputs(321) <= '0';
    layer2_outputs(322) <= not((layer1_outputs(6539)) or (layer1_outputs(1934)));
    layer2_outputs(323) <= '0';
    layer2_outputs(324) <= not((layer1_outputs(4601)) or (layer1_outputs(1124)));
    layer2_outputs(325) <= (layer1_outputs(5110)) and not (layer1_outputs(197));
    layer2_outputs(326) <= layer1_outputs(3474);
    layer2_outputs(327) <= not(layer1_outputs(1915));
    layer2_outputs(328) <= not(layer1_outputs(6153));
    layer2_outputs(329) <= layer1_outputs(1020);
    layer2_outputs(330) <= (layer1_outputs(4133)) or (layer1_outputs(6205));
    layer2_outputs(331) <= (layer1_outputs(5613)) and not (layer1_outputs(3125));
    layer2_outputs(332) <= (layer1_outputs(1270)) and (layer1_outputs(6789));
    layer2_outputs(333) <= layer1_outputs(3471);
    layer2_outputs(334) <= (layer1_outputs(4177)) xor (layer1_outputs(378));
    layer2_outputs(335) <= (layer1_outputs(3971)) and not (layer1_outputs(7223));
    layer2_outputs(336) <= layer1_outputs(1434);
    layer2_outputs(337) <= layer1_outputs(3206);
    layer2_outputs(338) <= not((layer1_outputs(3880)) and (layer1_outputs(2580)));
    layer2_outputs(339) <= (layer1_outputs(6574)) and not (layer1_outputs(3977));
    layer2_outputs(340) <= not(layer1_outputs(5697));
    layer2_outputs(341) <= (layer1_outputs(6256)) or (layer1_outputs(4179));
    layer2_outputs(342) <= not(layer1_outputs(3401));
    layer2_outputs(343) <= '1';
    layer2_outputs(344) <= (layer1_outputs(1090)) xor (layer1_outputs(3626));
    layer2_outputs(345) <= (layer1_outputs(636)) or (layer1_outputs(1030));
    layer2_outputs(346) <= not(layer1_outputs(1793));
    layer2_outputs(347) <= (layer1_outputs(6720)) and (layer1_outputs(3690));
    layer2_outputs(348) <= not((layer1_outputs(5014)) and (layer1_outputs(7178)));
    layer2_outputs(349) <= (layer1_outputs(3789)) and (layer1_outputs(2047));
    layer2_outputs(350) <= '0';
    layer2_outputs(351) <= not(layer1_outputs(266));
    layer2_outputs(352) <= (layer1_outputs(6179)) xor (layer1_outputs(3771));
    layer2_outputs(353) <= '0';
    layer2_outputs(354) <= (layer1_outputs(6779)) and not (layer1_outputs(4553));
    layer2_outputs(355) <= not(layer1_outputs(2877)) or (layer1_outputs(6426));
    layer2_outputs(356) <= not(layer1_outputs(6659));
    layer2_outputs(357) <= layer1_outputs(164);
    layer2_outputs(358) <= not((layer1_outputs(7515)) and (layer1_outputs(7331)));
    layer2_outputs(359) <= not(layer1_outputs(4238)) or (layer1_outputs(6562));
    layer2_outputs(360) <= (layer1_outputs(2712)) xor (layer1_outputs(2438));
    layer2_outputs(361) <= layer1_outputs(469);
    layer2_outputs(362) <= not(layer1_outputs(2132));
    layer2_outputs(363) <= not(layer1_outputs(572)) or (layer1_outputs(4027));
    layer2_outputs(364) <= (layer1_outputs(3928)) and (layer1_outputs(1347));
    layer2_outputs(365) <= (layer1_outputs(5836)) or (layer1_outputs(6300));
    layer2_outputs(366) <= not(layer1_outputs(2134));
    layer2_outputs(367) <= (layer1_outputs(6598)) and (layer1_outputs(4893));
    layer2_outputs(368) <= (layer1_outputs(1091)) and (layer1_outputs(5362));
    layer2_outputs(369) <= not((layer1_outputs(6699)) or (layer1_outputs(5728)));
    layer2_outputs(370) <= not(layer1_outputs(881));
    layer2_outputs(371) <= (layer1_outputs(3633)) and not (layer1_outputs(4764));
    layer2_outputs(372) <= not((layer1_outputs(2089)) or (layer1_outputs(2571)));
    layer2_outputs(373) <= '1';
    layer2_outputs(374) <= layer1_outputs(3489);
    layer2_outputs(375) <= not(layer1_outputs(444)) or (layer1_outputs(6789));
    layer2_outputs(376) <= not((layer1_outputs(1848)) or (layer1_outputs(1241)));
    layer2_outputs(377) <= '0';
    layer2_outputs(378) <= not((layer1_outputs(155)) or (layer1_outputs(619)));
    layer2_outputs(379) <= (layer1_outputs(7493)) and not (layer1_outputs(5614));
    layer2_outputs(380) <= not((layer1_outputs(1181)) or (layer1_outputs(299)));
    layer2_outputs(381) <= not(layer1_outputs(307));
    layer2_outputs(382) <= not(layer1_outputs(2885)) or (layer1_outputs(4835));
    layer2_outputs(383) <= not(layer1_outputs(5288));
    layer2_outputs(384) <= not((layer1_outputs(7230)) or (layer1_outputs(7044)));
    layer2_outputs(385) <= (layer1_outputs(1229)) and (layer1_outputs(1893));
    layer2_outputs(386) <= not(layer1_outputs(2651));
    layer2_outputs(387) <= layer1_outputs(6050);
    layer2_outputs(388) <= layer1_outputs(1399);
    layer2_outputs(389) <= (layer1_outputs(4778)) and not (layer1_outputs(1378));
    layer2_outputs(390) <= (layer1_outputs(5948)) or (layer1_outputs(4774));
    layer2_outputs(391) <= not(layer1_outputs(1229));
    layer2_outputs(392) <= not((layer1_outputs(4267)) or (layer1_outputs(3485)));
    layer2_outputs(393) <= (layer1_outputs(4355)) and not (layer1_outputs(7109));
    layer2_outputs(394) <= '1';
    layer2_outputs(395) <= not(layer1_outputs(2906));
    layer2_outputs(396) <= layer1_outputs(5615);
    layer2_outputs(397) <= '1';
    layer2_outputs(398) <= layer1_outputs(7495);
    layer2_outputs(399) <= not((layer1_outputs(3352)) or (layer1_outputs(4222)));
    layer2_outputs(400) <= not(layer1_outputs(2817));
    layer2_outputs(401) <= not(layer1_outputs(1500));
    layer2_outputs(402) <= layer1_outputs(1140);
    layer2_outputs(403) <= (layer1_outputs(2033)) and not (layer1_outputs(2085));
    layer2_outputs(404) <= not((layer1_outputs(1272)) and (layer1_outputs(4853)));
    layer2_outputs(405) <= not(layer1_outputs(5141));
    layer2_outputs(406) <= (layer1_outputs(3742)) and not (layer1_outputs(2096));
    layer2_outputs(407) <= not((layer1_outputs(4384)) or (layer1_outputs(5091)));
    layer2_outputs(408) <= not(layer1_outputs(6469));
    layer2_outputs(409) <= '0';
    layer2_outputs(410) <= '1';
    layer2_outputs(411) <= '1';
    layer2_outputs(412) <= not((layer1_outputs(250)) and (layer1_outputs(4374)));
    layer2_outputs(413) <= layer1_outputs(7003);
    layer2_outputs(414) <= not(layer1_outputs(6030)) or (layer1_outputs(1909));
    layer2_outputs(415) <= '0';
    layer2_outputs(416) <= (layer1_outputs(3634)) and not (layer1_outputs(6870));
    layer2_outputs(417) <= (layer1_outputs(537)) and not (layer1_outputs(1808));
    layer2_outputs(418) <= not(layer1_outputs(1147)) or (layer1_outputs(3389));
    layer2_outputs(419) <= not((layer1_outputs(2800)) or (layer1_outputs(4064)));
    layer2_outputs(420) <= (layer1_outputs(3442)) and not (layer1_outputs(979));
    layer2_outputs(421) <= (layer1_outputs(676)) or (layer1_outputs(3456));
    layer2_outputs(422) <= layer1_outputs(5561);
    layer2_outputs(423) <= not(layer1_outputs(6761)) or (layer1_outputs(4808));
    layer2_outputs(424) <= layer1_outputs(1322);
    layer2_outputs(425) <= (layer1_outputs(7225)) or (layer1_outputs(2298));
    layer2_outputs(426) <= not(layer1_outputs(7475));
    layer2_outputs(427) <= '1';
    layer2_outputs(428) <= (layer1_outputs(620)) and not (layer1_outputs(7141));
    layer2_outputs(429) <= (layer1_outputs(3844)) and not (layer1_outputs(1749));
    layer2_outputs(430) <= not(layer1_outputs(5904)) or (layer1_outputs(3855));
    layer2_outputs(431) <= (layer1_outputs(2412)) or (layer1_outputs(4766));
    layer2_outputs(432) <= not(layer1_outputs(6046));
    layer2_outputs(433) <= '0';
    layer2_outputs(434) <= not(layer1_outputs(5879)) or (layer1_outputs(2732));
    layer2_outputs(435) <= '0';
    layer2_outputs(436) <= layer1_outputs(3853);
    layer2_outputs(437) <= (layer1_outputs(7448)) and not (layer1_outputs(1561));
    layer2_outputs(438) <= (layer1_outputs(3255)) and not (layer1_outputs(5242));
    layer2_outputs(439) <= layer1_outputs(5251);
    layer2_outputs(440) <= not((layer1_outputs(5180)) and (layer1_outputs(4712)));
    layer2_outputs(441) <= '1';
    layer2_outputs(442) <= (layer1_outputs(3043)) and not (layer1_outputs(194));
    layer2_outputs(443) <= layer1_outputs(5811);
    layer2_outputs(444) <= '1';
    layer2_outputs(445) <= not(layer1_outputs(4547)) or (layer1_outputs(5529));
    layer2_outputs(446) <= (layer1_outputs(1842)) or (layer1_outputs(2474));
    layer2_outputs(447) <= not(layer1_outputs(5416));
    layer2_outputs(448) <= layer1_outputs(6520);
    layer2_outputs(449) <= not(layer1_outputs(6705));
    layer2_outputs(450) <= not((layer1_outputs(6387)) and (layer1_outputs(3866)));
    layer2_outputs(451) <= '1';
    layer2_outputs(452) <= layer1_outputs(3153);
    layer2_outputs(453) <= (layer1_outputs(4524)) and not (layer1_outputs(910));
    layer2_outputs(454) <= not(layer1_outputs(2422));
    layer2_outputs(455) <= not(layer1_outputs(2680));
    layer2_outputs(456) <= layer1_outputs(326);
    layer2_outputs(457) <= (layer1_outputs(3619)) and not (layer1_outputs(6010));
    layer2_outputs(458) <= (layer1_outputs(4017)) and (layer1_outputs(7114));
    layer2_outputs(459) <= not((layer1_outputs(1189)) and (layer1_outputs(2895)));
    layer2_outputs(460) <= '0';
    layer2_outputs(461) <= not((layer1_outputs(542)) or (layer1_outputs(5134)));
    layer2_outputs(462) <= not(layer1_outputs(2262)) or (layer1_outputs(4105));
    layer2_outputs(463) <= '0';
    layer2_outputs(464) <= not((layer1_outputs(5692)) or (layer1_outputs(4420)));
    layer2_outputs(465) <= not((layer1_outputs(6731)) or (layer1_outputs(4655)));
    layer2_outputs(466) <= (layer1_outputs(4648)) and not (layer1_outputs(5021));
    layer2_outputs(467) <= not(layer1_outputs(262));
    layer2_outputs(468) <= not(layer1_outputs(1529));
    layer2_outputs(469) <= (layer1_outputs(978)) xor (layer1_outputs(561));
    layer2_outputs(470) <= (layer1_outputs(94)) or (layer1_outputs(3435));
    layer2_outputs(471) <= (layer1_outputs(3349)) and not (layer1_outputs(5509));
    layer2_outputs(472) <= '1';
    layer2_outputs(473) <= (layer1_outputs(179)) and not (layer1_outputs(7661));
    layer2_outputs(474) <= not(layer1_outputs(4791));
    layer2_outputs(475) <= layer1_outputs(1214);
    layer2_outputs(476) <= not(layer1_outputs(3156));
    layer2_outputs(477) <= '1';
    layer2_outputs(478) <= '0';
    layer2_outputs(479) <= layer1_outputs(3297);
    layer2_outputs(480) <= (layer1_outputs(7404)) and not (layer1_outputs(4080));
    layer2_outputs(481) <= not((layer1_outputs(5444)) and (layer1_outputs(1996)));
    layer2_outputs(482) <= layer1_outputs(2826);
    layer2_outputs(483) <= not((layer1_outputs(7366)) or (layer1_outputs(7648)));
    layer2_outputs(484) <= (layer1_outputs(3351)) or (layer1_outputs(275));
    layer2_outputs(485) <= not((layer1_outputs(646)) and (layer1_outputs(7410)));
    layer2_outputs(486) <= not((layer1_outputs(6571)) and (layer1_outputs(6823)));
    layer2_outputs(487) <= '1';
    layer2_outputs(488) <= (layer1_outputs(5370)) and not (layer1_outputs(2052));
    layer2_outputs(489) <= not(layer1_outputs(2451));
    layer2_outputs(490) <= not(layer1_outputs(4883)) or (layer1_outputs(4077));
    layer2_outputs(491) <= not((layer1_outputs(3381)) or (layer1_outputs(2553)));
    layer2_outputs(492) <= '1';
    layer2_outputs(493) <= not(layer1_outputs(3288)) or (layer1_outputs(2107));
    layer2_outputs(494) <= layer1_outputs(6499);
    layer2_outputs(495) <= not((layer1_outputs(7444)) and (layer1_outputs(2538)));
    layer2_outputs(496) <= (layer1_outputs(5988)) xor (layer1_outputs(181));
    layer2_outputs(497) <= (layer1_outputs(677)) or (layer1_outputs(6686));
    layer2_outputs(498) <= not(layer1_outputs(3281));
    layer2_outputs(499) <= (layer1_outputs(1625)) and not (layer1_outputs(440));
    layer2_outputs(500) <= not((layer1_outputs(1403)) or (layer1_outputs(1454)));
    layer2_outputs(501) <= (layer1_outputs(61)) and not (layer1_outputs(7242));
    layer2_outputs(502) <= layer1_outputs(1246);
    layer2_outputs(503) <= not((layer1_outputs(4704)) xor (layer1_outputs(7595)));
    layer2_outputs(504) <= layer1_outputs(511);
    layer2_outputs(505) <= (layer1_outputs(5724)) and (layer1_outputs(5882));
    layer2_outputs(506) <= layer1_outputs(937);
    layer2_outputs(507) <= layer1_outputs(4591);
    layer2_outputs(508) <= (layer1_outputs(434)) and not (layer1_outputs(3652));
    layer2_outputs(509) <= layer1_outputs(7484);
    layer2_outputs(510) <= (layer1_outputs(5056)) and (layer1_outputs(2647));
    layer2_outputs(511) <= '0';
    layer2_outputs(512) <= '0';
    layer2_outputs(513) <= not(layer1_outputs(4120)) or (layer1_outputs(1748));
    layer2_outputs(514) <= layer1_outputs(4769);
    layer2_outputs(515) <= '0';
    layer2_outputs(516) <= layer1_outputs(4057);
    layer2_outputs(517) <= not(layer1_outputs(2371));
    layer2_outputs(518) <= layer1_outputs(5596);
    layer2_outputs(519) <= layer1_outputs(518);
    layer2_outputs(520) <= layer1_outputs(5863);
    layer2_outputs(521) <= not((layer1_outputs(779)) or (layer1_outputs(1162)));
    layer2_outputs(522) <= (layer1_outputs(3233)) or (layer1_outputs(5979));
    layer2_outputs(523) <= (layer1_outputs(3946)) or (layer1_outputs(4026));
    layer2_outputs(524) <= not(layer1_outputs(4922)) or (layer1_outputs(2283));
    layer2_outputs(525) <= layer1_outputs(3126);
    layer2_outputs(526) <= layer1_outputs(2806);
    layer2_outputs(527) <= '1';
    layer2_outputs(528) <= layer1_outputs(7652);
    layer2_outputs(529) <= (layer1_outputs(3681)) and not (layer1_outputs(4988));
    layer2_outputs(530) <= layer1_outputs(813);
    layer2_outputs(531) <= (layer1_outputs(6494)) and (layer1_outputs(1026));
    layer2_outputs(532) <= layer1_outputs(3543);
    layer2_outputs(533) <= not((layer1_outputs(2488)) and (layer1_outputs(984)));
    layer2_outputs(534) <= (layer1_outputs(5854)) and not (layer1_outputs(5082));
    layer2_outputs(535) <= layer1_outputs(4128);
    layer2_outputs(536) <= (layer1_outputs(913)) and (layer1_outputs(5247));
    layer2_outputs(537) <= not((layer1_outputs(5299)) or (layer1_outputs(6453)));
    layer2_outputs(538) <= not(layer1_outputs(2684));
    layer2_outputs(539) <= '0';
    layer2_outputs(540) <= not(layer1_outputs(7272));
    layer2_outputs(541) <= '0';
    layer2_outputs(542) <= layer1_outputs(4469);
    layer2_outputs(543) <= not(layer1_outputs(2392));
    layer2_outputs(544) <= not(layer1_outputs(945)) or (layer1_outputs(707));
    layer2_outputs(545) <= not((layer1_outputs(6464)) and (layer1_outputs(2009)));
    layer2_outputs(546) <= layer1_outputs(6100);
    layer2_outputs(547) <= not(layer1_outputs(6703));
    layer2_outputs(548) <= (layer1_outputs(3401)) or (layer1_outputs(4856));
    layer2_outputs(549) <= layer1_outputs(1446);
    layer2_outputs(550) <= not((layer1_outputs(4689)) and (layer1_outputs(220)));
    layer2_outputs(551) <= not(layer1_outputs(7561));
    layer2_outputs(552) <= not((layer1_outputs(5553)) xor (layer1_outputs(7595)));
    layer2_outputs(553) <= layer1_outputs(5343);
    layer2_outputs(554) <= layer1_outputs(1554);
    layer2_outputs(555) <= not(layer1_outputs(4564)) or (layer1_outputs(6797));
    layer2_outputs(556) <= not(layer1_outputs(77)) or (layer1_outputs(4814));
    layer2_outputs(557) <= not((layer1_outputs(1728)) or (layer1_outputs(4927)));
    layer2_outputs(558) <= not(layer1_outputs(7673));
    layer2_outputs(559) <= '1';
    layer2_outputs(560) <= not(layer1_outputs(2164));
    layer2_outputs(561) <= (layer1_outputs(4329)) and not (layer1_outputs(1650));
    layer2_outputs(562) <= (layer1_outputs(245)) and not (layer1_outputs(1499));
    layer2_outputs(563) <= not(layer1_outputs(3831)) or (layer1_outputs(2095));
    layer2_outputs(564) <= '0';
    layer2_outputs(565) <= (layer1_outputs(3791)) or (layer1_outputs(7597));
    layer2_outputs(566) <= (layer1_outputs(5991)) or (layer1_outputs(7613));
    layer2_outputs(567) <= (layer1_outputs(1981)) and (layer1_outputs(1544));
    layer2_outputs(568) <= (layer1_outputs(4617)) and not (layer1_outputs(5198));
    layer2_outputs(569) <= not(layer1_outputs(4930));
    layer2_outputs(570) <= layer1_outputs(5531);
    layer2_outputs(571) <= not(layer1_outputs(1233)) or (layer1_outputs(5190));
    layer2_outputs(572) <= not((layer1_outputs(2345)) and (layer1_outputs(2364)));
    layer2_outputs(573) <= (layer1_outputs(5031)) xor (layer1_outputs(4997));
    layer2_outputs(574) <= '1';
    layer2_outputs(575) <= (layer1_outputs(3048)) and not (layer1_outputs(4295));
    layer2_outputs(576) <= (layer1_outputs(5558)) or (layer1_outputs(6612));
    layer2_outputs(577) <= not(layer1_outputs(3163)) or (layer1_outputs(5192));
    layer2_outputs(578) <= (layer1_outputs(2102)) and not (layer1_outputs(5907));
    layer2_outputs(579) <= not(layer1_outputs(7552));
    layer2_outputs(580) <= not((layer1_outputs(5210)) and (layer1_outputs(6185)));
    layer2_outputs(581) <= '0';
    layer2_outputs(582) <= layer1_outputs(2405);
    layer2_outputs(583) <= not(layer1_outputs(5486));
    layer2_outputs(584) <= not(layer1_outputs(4903)) or (layer1_outputs(3358));
    layer2_outputs(585) <= not(layer1_outputs(7315));
    layer2_outputs(586) <= (layer1_outputs(652)) and not (layer1_outputs(1137));
    layer2_outputs(587) <= (layer1_outputs(2127)) and not (layer1_outputs(4757));
    layer2_outputs(588) <= (layer1_outputs(2227)) and not (layer1_outputs(7396));
    layer2_outputs(589) <= not(layer1_outputs(3376)) or (layer1_outputs(3448));
    layer2_outputs(590) <= layer1_outputs(4559);
    layer2_outputs(591) <= '0';
    layer2_outputs(592) <= not(layer1_outputs(5619));
    layer2_outputs(593) <= not(layer1_outputs(3249));
    layer2_outputs(594) <= (layer1_outputs(7411)) and not (layer1_outputs(6475));
    layer2_outputs(595) <= (layer1_outputs(3774)) and not (layer1_outputs(4279));
    layer2_outputs(596) <= layer1_outputs(5128);
    layer2_outputs(597) <= layer1_outputs(3289);
    layer2_outputs(598) <= not((layer1_outputs(4584)) or (layer1_outputs(5638)));
    layer2_outputs(599) <= not(layer1_outputs(1758)) or (layer1_outputs(1850));
    layer2_outputs(600) <= layer1_outputs(4878);
    layer2_outputs(601) <= not(layer1_outputs(1023));
    layer2_outputs(602) <= not((layer1_outputs(2135)) and (layer1_outputs(882)));
    layer2_outputs(603) <= (layer1_outputs(4381)) and (layer1_outputs(3800));
    layer2_outputs(604) <= not(layer1_outputs(5009)) or (layer1_outputs(4579));
    layer2_outputs(605) <= not(layer1_outputs(6189)) or (layer1_outputs(7497));
    layer2_outputs(606) <= not(layer1_outputs(5860)) or (layer1_outputs(3348));
    layer2_outputs(607) <= layer1_outputs(3084);
    layer2_outputs(608) <= '0';
    layer2_outputs(609) <= (layer1_outputs(2820)) and not (layer1_outputs(5932));
    layer2_outputs(610) <= '0';
    layer2_outputs(611) <= '1';
    layer2_outputs(612) <= layer1_outputs(4672);
    layer2_outputs(613) <= (layer1_outputs(5517)) and not (layer1_outputs(137));
    layer2_outputs(614) <= not((layer1_outputs(2126)) and (layer1_outputs(2914)));
    layer2_outputs(615) <= '1';
    layer2_outputs(616) <= (layer1_outputs(2016)) or (layer1_outputs(2482));
    layer2_outputs(617) <= '0';
    layer2_outputs(618) <= layer1_outputs(4270);
    layer2_outputs(619) <= layer1_outputs(6578);
    layer2_outputs(620) <= not((layer1_outputs(842)) and (layer1_outputs(2388)));
    layer2_outputs(621) <= not(layer1_outputs(5780));
    layer2_outputs(622) <= (layer1_outputs(7550)) or (layer1_outputs(793));
    layer2_outputs(623) <= (layer1_outputs(6650)) or (layer1_outputs(3822));
    layer2_outputs(624) <= not(layer1_outputs(2690));
    layer2_outputs(625) <= '1';
    layer2_outputs(626) <= not(layer1_outputs(2335)) or (layer1_outputs(669));
    layer2_outputs(627) <= layer1_outputs(1382);
    layer2_outputs(628) <= '1';
    layer2_outputs(629) <= layer1_outputs(4706);
    layer2_outputs(630) <= not(layer1_outputs(4912));
    layer2_outputs(631) <= (layer1_outputs(943)) and not (layer1_outputs(1170));
    layer2_outputs(632) <= (layer1_outputs(5735)) and not (layer1_outputs(4530));
    layer2_outputs(633) <= (layer1_outputs(2498)) and (layer1_outputs(6525));
    layer2_outputs(634) <= not(layer1_outputs(5374)) or (layer1_outputs(1467));
    layer2_outputs(635) <= not((layer1_outputs(7614)) or (layer1_outputs(7508)));
    layer2_outputs(636) <= not(layer1_outputs(7290));
    layer2_outputs(637) <= '1';
    layer2_outputs(638) <= not(layer1_outputs(198));
    layer2_outputs(639) <= (layer1_outputs(5143)) or (layer1_outputs(1493));
    layer2_outputs(640) <= not(layer1_outputs(4867));
    layer2_outputs(641) <= (layer1_outputs(7081)) and not (layer1_outputs(6900));
    layer2_outputs(642) <= not(layer1_outputs(4998)) or (layer1_outputs(2383));
    layer2_outputs(643) <= (layer1_outputs(5565)) and not (layer1_outputs(4457));
    layer2_outputs(644) <= '1';
    layer2_outputs(645) <= not((layer1_outputs(587)) or (layer1_outputs(7452)));
    layer2_outputs(646) <= not(layer1_outputs(5918));
    layer2_outputs(647) <= '1';
    layer2_outputs(648) <= (layer1_outputs(4380)) and not (layer1_outputs(1));
    layer2_outputs(649) <= not((layer1_outputs(5277)) or (layer1_outputs(5136)));
    layer2_outputs(650) <= not((layer1_outputs(6675)) or (layer1_outputs(3267)));
    layer2_outputs(651) <= not(layer1_outputs(2411)) or (layer1_outputs(5696));
    layer2_outputs(652) <= layer1_outputs(1340);
    layer2_outputs(653) <= not(layer1_outputs(7500)) or (layer1_outputs(7596));
    layer2_outputs(654) <= not(layer1_outputs(2031)) or (layer1_outputs(249));
    layer2_outputs(655) <= (layer1_outputs(2381)) xor (layer1_outputs(7297));
    layer2_outputs(656) <= not((layer1_outputs(2751)) and (layer1_outputs(6129)));
    layer2_outputs(657) <= (layer1_outputs(4098)) and not (layer1_outputs(4202));
    layer2_outputs(658) <= (layer1_outputs(2632)) and not (layer1_outputs(647));
    layer2_outputs(659) <= not(layer1_outputs(7129));
    layer2_outputs(660) <= (layer1_outputs(3275)) and (layer1_outputs(994));
    layer2_outputs(661) <= (layer1_outputs(2671)) or (layer1_outputs(3603));
    layer2_outputs(662) <= layer1_outputs(5422);
    layer2_outputs(663) <= '1';
    layer2_outputs(664) <= '0';
    layer2_outputs(665) <= '1';
    layer2_outputs(666) <= '0';
    layer2_outputs(667) <= '0';
    layer2_outputs(668) <= layer1_outputs(705);
    layer2_outputs(669) <= '0';
    layer2_outputs(670) <= (layer1_outputs(1471)) and not (layer1_outputs(3282));
    layer2_outputs(671) <= '1';
    layer2_outputs(672) <= (layer1_outputs(6977)) and not (layer1_outputs(1722));
    layer2_outputs(673) <= (layer1_outputs(319)) and not (layer1_outputs(6587));
    layer2_outputs(674) <= '0';
    layer2_outputs(675) <= layer1_outputs(5880);
    layer2_outputs(676) <= not(layer1_outputs(109));
    layer2_outputs(677) <= not(layer1_outputs(3620));
    layer2_outputs(678) <= layer1_outputs(3031);
    layer2_outputs(679) <= not(layer1_outputs(310));
    layer2_outputs(680) <= not(layer1_outputs(766));
    layer2_outputs(681) <= not((layer1_outputs(2770)) or (layer1_outputs(2511)));
    layer2_outputs(682) <= (layer1_outputs(3202)) and not (layer1_outputs(3760));
    layer2_outputs(683) <= not(layer1_outputs(4652)) or (layer1_outputs(7360));
    layer2_outputs(684) <= layer1_outputs(933);
    layer2_outputs(685) <= (layer1_outputs(4575)) xor (layer1_outputs(817));
    layer2_outputs(686) <= (layer1_outputs(4511)) and not (layer1_outputs(215));
    layer2_outputs(687) <= (layer1_outputs(6533)) and not (layer1_outputs(1883));
    layer2_outputs(688) <= layer1_outputs(5795);
    layer2_outputs(689) <= not(layer1_outputs(7055)) or (layer1_outputs(4159));
    layer2_outputs(690) <= '0';
    layer2_outputs(691) <= '1';
    layer2_outputs(692) <= layer1_outputs(1532);
    layer2_outputs(693) <= layer1_outputs(2109);
    layer2_outputs(694) <= not(layer1_outputs(6951)) or (layer1_outputs(3459));
    layer2_outputs(695) <= not(layer1_outputs(4265)) or (layer1_outputs(1117));
    layer2_outputs(696) <= (layer1_outputs(7558)) and (layer1_outputs(1141));
    layer2_outputs(697) <= '0';
    layer2_outputs(698) <= '1';
    layer2_outputs(699) <= not((layer1_outputs(4284)) and (layer1_outputs(7642)));
    layer2_outputs(700) <= not(layer1_outputs(6516));
    layer2_outputs(701) <= not((layer1_outputs(384)) or (layer1_outputs(3485)));
    layer2_outputs(702) <= layer1_outputs(4740);
    layer2_outputs(703) <= (layer1_outputs(423)) and (layer1_outputs(773));
    layer2_outputs(704) <= (layer1_outputs(710)) or (layer1_outputs(659));
    layer2_outputs(705) <= layer1_outputs(6265);
    layer2_outputs(706) <= not((layer1_outputs(2845)) and (layer1_outputs(6860)));
    layer2_outputs(707) <= '1';
    layer2_outputs(708) <= '1';
    layer2_outputs(709) <= not(layer1_outputs(1059));
    layer2_outputs(710) <= '1';
    layer2_outputs(711) <= '1';
    layer2_outputs(712) <= (layer1_outputs(2196)) or (layer1_outputs(7474));
    layer2_outputs(713) <= '1';
    layer2_outputs(714) <= (layer1_outputs(6702)) or (layer1_outputs(4995));
    layer2_outputs(715) <= not(layer1_outputs(3659));
    layer2_outputs(716) <= not((layer1_outputs(4911)) or (layer1_outputs(6006)));
    layer2_outputs(717) <= '0';
    layer2_outputs(718) <= layer1_outputs(6776);
    layer2_outputs(719) <= not(layer1_outputs(3857)) or (layer1_outputs(3607));
    layer2_outputs(720) <= layer1_outputs(3278);
    layer2_outputs(721) <= not(layer1_outputs(48));
    layer2_outputs(722) <= layer1_outputs(356);
    layer2_outputs(723) <= (layer1_outputs(1575)) or (layer1_outputs(5351));
    layer2_outputs(724) <= not(layer1_outputs(1105));
    layer2_outputs(725) <= '0';
    layer2_outputs(726) <= layer1_outputs(1697);
    layer2_outputs(727) <= (layer1_outputs(4563)) and not (layer1_outputs(2110));
    layer2_outputs(728) <= layer1_outputs(294);
    layer2_outputs(729) <= layer1_outputs(6229);
    layer2_outputs(730) <= (layer1_outputs(3578)) and not (layer1_outputs(2481));
    layer2_outputs(731) <= layer1_outputs(6519);
    layer2_outputs(732) <= layer1_outputs(5404);
    layer2_outputs(733) <= not(layer1_outputs(3508));
    layer2_outputs(734) <= not(layer1_outputs(439)) or (layer1_outputs(7079));
    layer2_outputs(735) <= '1';
    layer2_outputs(736) <= not(layer1_outputs(295));
    layer2_outputs(737) <= layer1_outputs(775);
    layer2_outputs(738) <= not(layer1_outputs(2223)) or (layer1_outputs(53));
    layer2_outputs(739) <= layer1_outputs(3504);
    layer2_outputs(740) <= layer1_outputs(3847);
    layer2_outputs(741) <= (layer1_outputs(6905)) and not (layer1_outputs(2890));
    layer2_outputs(742) <= (layer1_outputs(1687)) and not (layer1_outputs(3222));
    layer2_outputs(743) <= not(layer1_outputs(4804)) or (layer1_outputs(3668));
    layer2_outputs(744) <= not(layer1_outputs(2299));
    layer2_outputs(745) <= not(layer1_outputs(1078)) or (layer1_outputs(4157));
    layer2_outputs(746) <= '0';
    layer2_outputs(747) <= not(layer1_outputs(5362)) or (layer1_outputs(5278));
    layer2_outputs(748) <= layer1_outputs(2239);
    layer2_outputs(749) <= '0';
    layer2_outputs(750) <= (layer1_outputs(14)) and (layer1_outputs(6026));
    layer2_outputs(751) <= not((layer1_outputs(3000)) or (layer1_outputs(6887)));
    layer2_outputs(752) <= not((layer1_outputs(5216)) and (layer1_outputs(5987)));
    layer2_outputs(753) <= not(layer1_outputs(4782));
    layer2_outputs(754) <= not(layer1_outputs(5475)) or (layer1_outputs(579));
    layer2_outputs(755) <= not((layer1_outputs(45)) or (layer1_outputs(3818)));
    layer2_outputs(756) <= not(layer1_outputs(2763));
    layer2_outputs(757) <= not((layer1_outputs(370)) and (layer1_outputs(2061)));
    layer2_outputs(758) <= not((layer1_outputs(3142)) and (layer1_outputs(4127)));
    layer2_outputs(759) <= '1';
    layer2_outputs(760) <= not((layer1_outputs(2336)) and (layer1_outputs(409)));
    layer2_outputs(761) <= not(layer1_outputs(6235));
    layer2_outputs(762) <= layer1_outputs(883);
    layer2_outputs(763) <= not(layer1_outputs(2733));
    layer2_outputs(764) <= layer1_outputs(849);
    layer2_outputs(765) <= '0';
    layer2_outputs(766) <= (layer1_outputs(2783)) and not (layer1_outputs(6500));
    layer2_outputs(767) <= (layer1_outputs(6669)) and (layer1_outputs(3419));
    layer2_outputs(768) <= layer1_outputs(4790);
    layer2_outputs(769) <= not(layer1_outputs(1429));
    layer2_outputs(770) <= (layer1_outputs(338)) or (layer1_outputs(4079));
    layer2_outputs(771) <= (layer1_outputs(3555)) and not (layer1_outputs(5310));
    layer2_outputs(772) <= not(layer1_outputs(3101));
    layer2_outputs(773) <= not(layer1_outputs(5141)) or (layer1_outputs(3972));
    layer2_outputs(774) <= '1';
    layer2_outputs(775) <= '1';
    layer2_outputs(776) <= not(layer1_outputs(3193)) or (layer1_outputs(2512));
    layer2_outputs(777) <= not(layer1_outputs(5473));
    layer2_outputs(778) <= (layer1_outputs(3788)) xor (layer1_outputs(6943));
    layer2_outputs(779) <= '1';
    layer2_outputs(780) <= (layer1_outputs(927)) and (layer1_outputs(1341));
    layer2_outputs(781) <= layer1_outputs(5921);
    layer2_outputs(782) <= not(layer1_outputs(4272));
    layer2_outputs(783) <= not(layer1_outputs(120));
    layer2_outputs(784) <= not(layer1_outputs(188));
    layer2_outputs(785) <= '0';
    layer2_outputs(786) <= not(layer1_outputs(4936)) or (layer1_outputs(3919));
    layer2_outputs(787) <= layer1_outputs(1338);
    layer2_outputs(788) <= (layer1_outputs(4523)) and not (layer1_outputs(6193));
    layer2_outputs(789) <= '1';
    layer2_outputs(790) <= layer1_outputs(2549);
    layer2_outputs(791) <= not(layer1_outputs(6731));
    layer2_outputs(792) <= not(layer1_outputs(5052)) or (layer1_outputs(4864));
    layer2_outputs(793) <= (layer1_outputs(2346)) and (layer1_outputs(1288));
    layer2_outputs(794) <= not((layer1_outputs(4736)) and (layer1_outputs(5118)));
    layer2_outputs(795) <= not((layer1_outputs(7442)) and (layer1_outputs(6434)));
    layer2_outputs(796) <= (layer1_outputs(5674)) and not (layer1_outputs(1068));
    layer2_outputs(797) <= '1';
    layer2_outputs(798) <= layer1_outputs(7217);
    layer2_outputs(799) <= layer1_outputs(5985);
    layer2_outputs(800) <= not((layer1_outputs(507)) or (layer1_outputs(6853)));
    layer2_outputs(801) <= layer1_outputs(7339);
    layer2_outputs(802) <= '1';
    layer2_outputs(803) <= '0';
    layer2_outputs(804) <= not(layer1_outputs(2146)) or (layer1_outputs(5962));
    layer2_outputs(805) <= '1';
    layer2_outputs(806) <= '1';
    layer2_outputs(807) <= (layer1_outputs(12)) and (layer1_outputs(1514));
    layer2_outputs(808) <= not(layer1_outputs(3055));
    layer2_outputs(809) <= not(layer1_outputs(5673)) or (layer1_outputs(3238));
    layer2_outputs(810) <= not(layer1_outputs(1879)) or (layer1_outputs(7128));
    layer2_outputs(811) <= (layer1_outputs(6508)) and not (layer1_outputs(1332));
    layer2_outputs(812) <= '0';
    layer2_outputs(813) <= not((layer1_outputs(524)) or (layer1_outputs(4056)));
    layer2_outputs(814) <= layer1_outputs(1899);
    layer2_outputs(815) <= (layer1_outputs(4185)) or (layer1_outputs(2900));
    layer2_outputs(816) <= not(layer1_outputs(2755)) or (layer1_outputs(6498));
    layer2_outputs(817) <= not(layer1_outputs(4156));
    layer2_outputs(818) <= layer1_outputs(1331);
    layer2_outputs(819) <= not(layer1_outputs(6304)) or (layer1_outputs(204));
    layer2_outputs(820) <= (layer1_outputs(4568)) and (layer1_outputs(2217));
    layer2_outputs(821) <= not(layer1_outputs(7617));
    layer2_outputs(822) <= not((layer1_outputs(3691)) or (layer1_outputs(525)));
    layer2_outputs(823) <= not((layer1_outputs(196)) and (layer1_outputs(2438)));
    layer2_outputs(824) <= not(layer1_outputs(5790));
    layer2_outputs(825) <= not(layer1_outputs(7147));
    layer2_outputs(826) <= not(layer1_outputs(4534));
    layer2_outputs(827) <= (layer1_outputs(3600)) and (layer1_outputs(4162));
    layer2_outputs(828) <= '1';
    layer2_outputs(829) <= not(layer1_outputs(3749)) or (layer1_outputs(795));
    layer2_outputs(830) <= (layer1_outputs(4509)) and (layer1_outputs(4187));
    layer2_outputs(831) <= '1';
    layer2_outputs(832) <= '0';
    layer2_outputs(833) <= not(layer1_outputs(5633));
    layer2_outputs(834) <= not((layer1_outputs(4083)) and (layer1_outputs(6620)));
    layer2_outputs(835) <= not(layer1_outputs(2169));
    layer2_outputs(836) <= (layer1_outputs(485)) or (layer1_outputs(5438));
    layer2_outputs(837) <= not(layer1_outputs(7091)) or (layer1_outputs(6307));
    layer2_outputs(838) <= layer1_outputs(5524);
    layer2_outputs(839) <= '1';
    layer2_outputs(840) <= not(layer1_outputs(1879)) or (layer1_outputs(2254));
    layer2_outputs(841) <= not(layer1_outputs(2277)) or (layer1_outputs(4723));
    layer2_outputs(842) <= not(layer1_outputs(2513));
    layer2_outputs(843) <= (layer1_outputs(5426)) and not (layer1_outputs(5963));
    layer2_outputs(844) <= layer1_outputs(2217);
    layer2_outputs(845) <= not(layer1_outputs(7094));
    layer2_outputs(846) <= '0';
    layer2_outputs(847) <= not(layer1_outputs(7415));
    layer2_outputs(848) <= (layer1_outputs(2111)) and (layer1_outputs(6125));
    layer2_outputs(849) <= not(layer1_outputs(4481)) or (layer1_outputs(4810));
    layer2_outputs(850) <= not(layer1_outputs(5084));
    layer2_outputs(851) <= not((layer1_outputs(175)) or (layer1_outputs(6471)));
    layer2_outputs(852) <= not(layer1_outputs(2625));
    layer2_outputs(853) <= (layer1_outputs(2152)) and not (layer1_outputs(5299));
    layer2_outputs(854) <= (layer1_outputs(1953)) and not (layer1_outputs(1581));
    layer2_outputs(855) <= layer1_outputs(1577);
    layer2_outputs(856) <= (layer1_outputs(1099)) xor (layer1_outputs(5089));
    layer2_outputs(857) <= not(layer1_outputs(5547)) or (layer1_outputs(5923));
    layer2_outputs(858) <= '0';
    layer2_outputs(859) <= '0';
    layer2_outputs(860) <= (layer1_outputs(1037)) and not (layer1_outputs(2713));
    layer2_outputs(861) <= not(layer1_outputs(3437));
    layer2_outputs(862) <= (layer1_outputs(6442)) and not (layer1_outputs(2304));
    layer2_outputs(863) <= not(layer1_outputs(4521));
    layer2_outputs(864) <= not(layer1_outputs(3011));
    layer2_outputs(865) <= (layer1_outputs(6873)) or (layer1_outputs(592));
    layer2_outputs(866) <= (layer1_outputs(732)) and not (layer1_outputs(7051));
    layer2_outputs(867) <= '0';
    layer2_outputs(868) <= (layer1_outputs(5599)) xor (layer1_outputs(5338));
    layer2_outputs(869) <= not(layer1_outputs(1304));
    layer2_outputs(870) <= not(layer1_outputs(2896));
    layer2_outputs(871) <= '0';
    layer2_outputs(872) <= (layer1_outputs(6366)) and not (layer1_outputs(3187));
    layer2_outputs(873) <= not(layer1_outputs(2288)) or (layer1_outputs(6496));
    layer2_outputs(874) <= not((layer1_outputs(5375)) and (layer1_outputs(7236)));
    layer2_outputs(875) <= layer1_outputs(4539);
    layer2_outputs(876) <= (layer1_outputs(1230)) or (layer1_outputs(27));
    layer2_outputs(877) <= '1';
    layer2_outputs(878) <= layer1_outputs(6328);
    layer2_outputs(879) <= (layer1_outputs(29)) xor (layer1_outputs(5471));
    layer2_outputs(880) <= not(layer1_outputs(7036));
    layer2_outputs(881) <= (layer1_outputs(4371)) and not (layer1_outputs(459));
    layer2_outputs(882) <= not((layer1_outputs(7607)) xor (layer1_outputs(201)));
    layer2_outputs(883) <= not((layer1_outputs(6730)) or (layer1_outputs(1067)));
    layer2_outputs(884) <= layer1_outputs(503);
    layer2_outputs(885) <= not(layer1_outputs(7640));
    layer2_outputs(886) <= not(layer1_outputs(4369)) or (layer1_outputs(354));
    layer2_outputs(887) <= not(layer1_outputs(159));
    layer2_outputs(888) <= not(layer1_outputs(1594));
    layer2_outputs(889) <= layer1_outputs(980);
    layer2_outputs(890) <= (layer1_outputs(3679)) and not (layer1_outputs(4447));
    layer2_outputs(891) <= not((layer1_outputs(7488)) or (layer1_outputs(7036)));
    layer2_outputs(892) <= not(layer1_outputs(1129));
    layer2_outputs(893) <= '1';
    layer2_outputs(894) <= layer1_outputs(6138);
    layer2_outputs(895) <= (layer1_outputs(1057)) and (layer1_outputs(2600));
    layer2_outputs(896) <= not(layer1_outputs(6897));
    layer2_outputs(897) <= not((layer1_outputs(4586)) or (layer1_outputs(6960)));
    layer2_outputs(898) <= (layer1_outputs(2842)) and not (layer1_outputs(4282));
    layer2_outputs(899) <= (layer1_outputs(5349)) and (layer1_outputs(4765));
    layer2_outputs(900) <= not(layer1_outputs(344));
    layer2_outputs(901) <= not(layer1_outputs(6435)) or (layer1_outputs(5784));
    layer2_outputs(902) <= layer1_outputs(768);
    layer2_outputs(903) <= (layer1_outputs(7017)) or (layer1_outputs(5825));
    layer2_outputs(904) <= not(layer1_outputs(2140)) or (layer1_outputs(7289));
    layer2_outputs(905) <= (layer1_outputs(2729)) and (layer1_outputs(257));
    layer2_outputs(906) <= '1';
    layer2_outputs(907) <= (layer1_outputs(2458)) and (layer1_outputs(3383));
    layer2_outputs(908) <= layer1_outputs(3362);
    layer2_outputs(909) <= '1';
    layer2_outputs(910) <= '1';
    layer2_outputs(911) <= '1';
    layer2_outputs(912) <= layer1_outputs(5740);
    layer2_outputs(913) <= not(layer1_outputs(5426)) or (layer1_outputs(2366));
    layer2_outputs(914) <= '1';
    layer2_outputs(915) <= not(layer1_outputs(6943));
    layer2_outputs(916) <= not(layer1_outputs(6854)) or (layer1_outputs(2686));
    layer2_outputs(917) <= layer1_outputs(6976);
    layer2_outputs(918) <= (layer1_outputs(2961)) and (layer1_outputs(7350));
    layer2_outputs(919) <= layer1_outputs(632);
    layer2_outputs(920) <= '0';
    layer2_outputs(921) <= '1';
    layer2_outputs(922) <= (layer1_outputs(7075)) and not (layer1_outputs(2864));
    layer2_outputs(923) <= layer1_outputs(146);
    layer2_outputs(924) <= not((layer1_outputs(1602)) or (layer1_outputs(6899)));
    layer2_outputs(925) <= not(layer1_outputs(3394));
    layer2_outputs(926) <= '0';
    layer2_outputs(927) <= not((layer1_outputs(864)) and (layer1_outputs(2818)));
    layer2_outputs(928) <= '1';
    layer2_outputs(929) <= not(layer1_outputs(6382)) or (layer1_outputs(3808));
    layer2_outputs(930) <= (layer1_outputs(7127)) or (layer1_outputs(4310));
    layer2_outputs(931) <= not(layer1_outputs(6967)) or (layer1_outputs(6256));
    layer2_outputs(932) <= '1';
    layer2_outputs(933) <= layer1_outputs(4930);
    layer2_outputs(934) <= not(layer1_outputs(595)) or (layer1_outputs(5577));
    layer2_outputs(935) <= not(layer1_outputs(2329));
    layer2_outputs(936) <= layer1_outputs(4613);
    layer2_outputs(937) <= not((layer1_outputs(4557)) and (layer1_outputs(2933)));
    layer2_outputs(938) <= (layer1_outputs(7092)) or (layer1_outputs(1905));
    layer2_outputs(939) <= layer1_outputs(1217);
    layer2_outputs(940) <= not(layer1_outputs(5399));
    layer2_outputs(941) <= '1';
    layer2_outputs(942) <= (layer1_outputs(1885)) and (layer1_outputs(4850));
    layer2_outputs(943) <= layer1_outputs(1560);
    layer2_outputs(944) <= not((layer1_outputs(4290)) or (layer1_outputs(2891)));
    layer2_outputs(945) <= (layer1_outputs(5135)) and not (layer1_outputs(7601));
    layer2_outputs(946) <= not(layer1_outputs(5936)) or (layer1_outputs(4777));
    layer2_outputs(947) <= not((layer1_outputs(5747)) and (layer1_outputs(2158)));
    layer2_outputs(948) <= (layer1_outputs(3680)) and (layer1_outputs(3834));
    layer2_outputs(949) <= not(layer1_outputs(5308)) or (layer1_outputs(6611));
    layer2_outputs(950) <= not(layer1_outputs(4446));
    layer2_outputs(951) <= (layer1_outputs(3522)) xor (layer1_outputs(4059));
    layer2_outputs(952) <= (layer1_outputs(5159)) and (layer1_outputs(4212));
    layer2_outputs(953) <= layer1_outputs(4512);
    layer2_outputs(954) <= (layer1_outputs(6052)) and not (layer1_outputs(7015));
    layer2_outputs(955) <= '0';
    layer2_outputs(956) <= '1';
    layer2_outputs(957) <= '0';
    layer2_outputs(958) <= not(layer1_outputs(3071));
    layer2_outputs(959) <= '1';
    layer2_outputs(960) <= (layer1_outputs(4303)) and not (layer1_outputs(5382));
    layer2_outputs(961) <= not((layer1_outputs(3105)) or (layer1_outputs(834)));
    layer2_outputs(962) <= not(layer1_outputs(5644)) or (layer1_outputs(6385));
    layer2_outputs(963) <= not(layer1_outputs(869)) or (layer1_outputs(1156));
    layer2_outputs(964) <= (layer1_outputs(1054)) and not (layer1_outputs(5959));
    layer2_outputs(965) <= not((layer1_outputs(6914)) or (layer1_outputs(1878)));
    layer2_outputs(966) <= not(layer1_outputs(6492));
    layer2_outputs(967) <= (layer1_outputs(6113)) and not (layer1_outputs(7545));
    layer2_outputs(968) <= '0';
    layer2_outputs(969) <= not((layer1_outputs(5452)) and (layer1_outputs(3067)));
    layer2_outputs(970) <= layer1_outputs(18);
    layer2_outputs(971) <= (layer1_outputs(1076)) and (layer1_outputs(1799));
    layer2_outputs(972) <= not((layer1_outputs(631)) or (layer1_outputs(4231)));
    layer2_outputs(973) <= '1';
    layer2_outputs(974) <= not((layer1_outputs(3253)) or (layer1_outputs(6554)));
    layer2_outputs(975) <= not((layer1_outputs(1829)) and (layer1_outputs(1705)));
    layer2_outputs(976) <= not(layer1_outputs(621));
    layer2_outputs(977) <= not(layer1_outputs(7106)) or (layer1_outputs(5169));
    layer2_outputs(978) <= not((layer1_outputs(1057)) or (layer1_outputs(4772)));
    layer2_outputs(979) <= not(layer1_outputs(2059)) or (layer1_outputs(4270));
    layer2_outputs(980) <= (layer1_outputs(5109)) and not (layer1_outputs(1563));
    layer2_outputs(981) <= layer1_outputs(581);
    layer2_outputs(982) <= not(layer1_outputs(6716));
    layer2_outputs(983) <= (layer1_outputs(1548)) and (layer1_outputs(3808));
    layer2_outputs(984) <= (layer1_outputs(6747)) and not (layer1_outputs(4574));
    layer2_outputs(985) <= layer1_outputs(4103);
    layer2_outputs(986) <= '0';
    layer2_outputs(987) <= '0';
    layer2_outputs(988) <= not(layer1_outputs(6276)) or (layer1_outputs(4688));
    layer2_outputs(989) <= '1';
    layer2_outputs(990) <= layer1_outputs(5592);
    layer2_outputs(991) <= not((layer1_outputs(5027)) or (layer1_outputs(6443)));
    layer2_outputs(992) <= not(layer1_outputs(4255)) or (layer1_outputs(6738));
    layer2_outputs(993) <= (layer1_outputs(1040)) or (layer1_outputs(2781));
    layer2_outputs(994) <= layer1_outputs(4122);
    layer2_outputs(995) <= not(layer1_outputs(4263));
    layer2_outputs(996) <= (layer1_outputs(1150)) and (layer1_outputs(4740));
    layer2_outputs(997) <= '0';
    layer2_outputs(998) <= (layer1_outputs(1800)) and not (layer1_outputs(5381));
    layer2_outputs(999) <= not(layer1_outputs(143)) or (layer1_outputs(1027));
    layer2_outputs(1000) <= not(layer1_outputs(2318));
    layer2_outputs(1001) <= layer1_outputs(1162);
    layer2_outputs(1002) <= not(layer1_outputs(7154));
    layer2_outputs(1003) <= not(layer1_outputs(3750));
    layer2_outputs(1004) <= layer1_outputs(6451);
    layer2_outputs(1005) <= layer1_outputs(1025);
    layer2_outputs(1006) <= not(layer1_outputs(3154)) or (layer1_outputs(5646));
    layer2_outputs(1007) <= (layer1_outputs(6913)) and not (layer1_outputs(5171));
    layer2_outputs(1008) <= (layer1_outputs(2637)) and not (layer1_outputs(6585));
    layer2_outputs(1009) <= not(layer1_outputs(5386));
    layer2_outputs(1010) <= '1';
    layer2_outputs(1011) <= (layer1_outputs(3190)) and not (layer1_outputs(105));
    layer2_outputs(1012) <= not(layer1_outputs(3905));
    layer2_outputs(1013) <= not((layer1_outputs(4921)) and (layer1_outputs(5654)));
    layer2_outputs(1014) <= not((layer1_outputs(3501)) or (layer1_outputs(705)));
    layer2_outputs(1015) <= not((layer1_outputs(6438)) and (layer1_outputs(236)));
    layer2_outputs(1016) <= layer1_outputs(1789);
    layer2_outputs(1017) <= layer1_outputs(2662);
    layer2_outputs(1018) <= (layer1_outputs(6802)) and (layer1_outputs(6139));
    layer2_outputs(1019) <= not(layer1_outputs(6305)) or (layer1_outputs(3689));
    layer2_outputs(1020) <= not((layer1_outputs(4397)) and (layer1_outputs(5144)));
    layer2_outputs(1021) <= layer1_outputs(5743);
    layer2_outputs(1022) <= not(layer1_outputs(7371));
    layer2_outputs(1023) <= (layer1_outputs(3660)) and not (layer1_outputs(4713));
    layer2_outputs(1024) <= (layer1_outputs(1842)) and not (layer1_outputs(5621));
    layer2_outputs(1025) <= (layer1_outputs(6326)) or (layer1_outputs(2537));
    layer2_outputs(1026) <= (layer1_outputs(2372)) and (layer1_outputs(4797));
    layer2_outputs(1027) <= not(layer1_outputs(4892)) or (layer1_outputs(946));
    layer2_outputs(1028) <= not(layer1_outputs(2234));
    layer2_outputs(1029) <= (layer1_outputs(5571)) or (layer1_outputs(3763));
    layer2_outputs(1030) <= (layer1_outputs(4504)) or (layer1_outputs(1220));
    layer2_outputs(1031) <= not(layer1_outputs(7181));
    layer2_outputs(1032) <= layer1_outputs(4972);
    layer2_outputs(1033) <= layer1_outputs(7300);
    layer2_outputs(1034) <= '0';
    layer2_outputs(1035) <= layer1_outputs(5041);
    layer2_outputs(1036) <= not(layer1_outputs(7511)) or (layer1_outputs(7531));
    layer2_outputs(1037) <= '0';
    layer2_outputs(1038) <= '1';
    layer2_outputs(1039) <= not(layer1_outputs(3465)) or (layer1_outputs(127));
    layer2_outputs(1040) <= (layer1_outputs(5006)) and (layer1_outputs(6444));
    layer2_outputs(1041) <= layer1_outputs(2060);
    layer2_outputs(1042) <= not((layer1_outputs(5157)) or (layer1_outputs(3041)));
    layer2_outputs(1043) <= '1';
    layer2_outputs(1044) <= not(layer1_outputs(5472));
    layer2_outputs(1045) <= layer1_outputs(4559);
    layer2_outputs(1046) <= '1';
    layer2_outputs(1047) <= (layer1_outputs(6904)) and (layer1_outputs(1115));
    layer2_outputs(1048) <= not(layer1_outputs(3805));
    layer2_outputs(1049) <= (layer1_outputs(3889)) or (layer1_outputs(2581));
    layer2_outputs(1050) <= '1';
    layer2_outputs(1051) <= not(layer1_outputs(4021));
    layer2_outputs(1052) <= (layer1_outputs(1652)) and not (layer1_outputs(1643));
    layer2_outputs(1053) <= not(layer1_outputs(6685)) or (layer1_outputs(497));
    layer2_outputs(1054) <= not(layer1_outputs(5607)) or (layer1_outputs(6332));
    layer2_outputs(1055) <= not(layer1_outputs(1331));
    layer2_outputs(1056) <= (layer1_outputs(1692)) and (layer1_outputs(7376));
    layer2_outputs(1057) <= (layer1_outputs(6991)) and not (layer1_outputs(850));
    layer2_outputs(1058) <= layer1_outputs(4254);
    layer2_outputs(1059) <= not(layer1_outputs(821));
    layer2_outputs(1060) <= not(layer1_outputs(3502));
    layer2_outputs(1061) <= layer1_outputs(6529);
    layer2_outputs(1062) <= not(layer1_outputs(917)) or (layer1_outputs(3624));
    layer2_outputs(1063) <= not(layer1_outputs(5490));
    layer2_outputs(1064) <= (layer1_outputs(1230)) or (layer1_outputs(7671));
    layer2_outputs(1065) <= (layer1_outputs(1077)) and (layer1_outputs(5055));
    layer2_outputs(1066) <= layer1_outputs(1494);
    layer2_outputs(1067) <= not((layer1_outputs(1891)) and (layer1_outputs(4324)));
    layer2_outputs(1068) <= not((layer1_outputs(6424)) or (layer1_outputs(2292)));
    layer2_outputs(1069) <= not(layer1_outputs(3730));
    layer2_outputs(1070) <= '1';
    layer2_outputs(1071) <= '0';
    layer2_outputs(1072) <= (layer1_outputs(4487)) and not (layer1_outputs(1700));
    layer2_outputs(1073) <= layer1_outputs(46);
    layer2_outputs(1074) <= layer1_outputs(2394);
    layer2_outputs(1075) <= '1';
    layer2_outputs(1076) <= not(layer1_outputs(1408));
    layer2_outputs(1077) <= (layer1_outputs(3054)) xor (layer1_outputs(7524));
    layer2_outputs(1078) <= '0';
    layer2_outputs(1079) <= not(layer1_outputs(119));
    layer2_outputs(1080) <= not(layer1_outputs(2687));
    layer2_outputs(1081) <= not(layer1_outputs(7006));
    layer2_outputs(1082) <= layer1_outputs(320);
    layer2_outputs(1083) <= '1';
    layer2_outputs(1084) <= not(layer1_outputs(2484));
    layer2_outputs(1085) <= layer1_outputs(6203);
    layer2_outputs(1086) <= (layer1_outputs(7622)) and (layer1_outputs(1930));
    layer2_outputs(1087) <= layer1_outputs(4599);
    layer2_outputs(1088) <= not(layer1_outputs(3924));
    layer2_outputs(1089) <= not(layer1_outputs(3175)) or (layer1_outputs(5001));
    layer2_outputs(1090) <= not(layer1_outputs(229)) or (layer1_outputs(2796));
    layer2_outputs(1091) <= layer1_outputs(6219);
    layer2_outputs(1092) <= not(layer1_outputs(5413));
    layer2_outputs(1093) <= not(layer1_outputs(4342));
    layer2_outputs(1094) <= layer1_outputs(2257);
    layer2_outputs(1095) <= not((layer1_outputs(4390)) and (layer1_outputs(2254)));
    layer2_outputs(1096) <= '1';
    layer2_outputs(1097) <= '0';
    layer2_outputs(1098) <= (layer1_outputs(4580)) and not (layer1_outputs(4033));
    layer2_outputs(1099) <= '0';
    layer2_outputs(1100) <= '1';
    layer2_outputs(1101) <= (layer1_outputs(6436)) and not (layer1_outputs(1433));
    layer2_outputs(1102) <= '1';
    layer2_outputs(1103) <= (layer1_outputs(3321)) and not (layer1_outputs(5697));
    layer2_outputs(1104) <= (layer1_outputs(4642)) and not (layer1_outputs(470));
    layer2_outputs(1105) <= not(layer1_outputs(6779));
    layer2_outputs(1106) <= (layer1_outputs(5981)) and not (layer1_outputs(4247));
    layer2_outputs(1107) <= layer1_outputs(6197);
    layer2_outputs(1108) <= not((layer1_outputs(5519)) or (layer1_outputs(5207)));
    layer2_outputs(1109) <= not(layer1_outputs(5234));
    layer2_outputs(1110) <= (layer1_outputs(1142)) or (layer1_outputs(5903));
    layer2_outputs(1111) <= (layer1_outputs(6054)) and (layer1_outputs(20));
    layer2_outputs(1112) <= '0';
    layer2_outputs(1113) <= layer1_outputs(5102);
    layer2_outputs(1114) <= not((layer1_outputs(6377)) or (layer1_outputs(1033)));
    layer2_outputs(1115) <= not(layer1_outputs(2655));
    layer2_outputs(1116) <= not(layer1_outputs(1125)) or (layer1_outputs(4004));
    layer2_outputs(1117) <= not(layer1_outputs(1327)) or (layer1_outputs(6743));
    layer2_outputs(1118) <= (layer1_outputs(3942)) and not (layer1_outputs(7393));
    layer2_outputs(1119) <= (layer1_outputs(5279)) and not (layer1_outputs(5650));
    layer2_outputs(1120) <= not(layer1_outputs(823));
    layer2_outputs(1121) <= '1';
    layer2_outputs(1122) <= '1';
    layer2_outputs(1123) <= not((layer1_outputs(7048)) and (layer1_outputs(5909)));
    layer2_outputs(1124) <= layer1_outputs(5511);
    layer2_outputs(1125) <= '1';
    layer2_outputs(1126) <= not(layer1_outputs(5925)) or (layer1_outputs(218));
    layer2_outputs(1127) <= layer1_outputs(4792);
    layer2_outputs(1128) <= '0';
    layer2_outputs(1129) <= not(layer1_outputs(908)) or (layer1_outputs(7212));
    layer2_outputs(1130) <= (layer1_outputs(3005)) or (layer1_outputs(1779));
    layer2_outputs(1131) <= layer1_outputs(3216);
    layer2_outputs(1132) <= not((layer1_outputs(6208)) or (layer1_outputs(398)));
    layer2_outputs(1133) <= '0';
    layer2_outputs(1134) <= layer1_outputs(5398);
    layer2_outputs(1135) <= not((layer1_outputs(5187)) and (layer1_outputs(124)));
    layer2_outputs(1136) <= layer1_outputs(2357);
    layer2_outputs(1137) <= not(layer1_outputs(6000)) or (layer1_outputs(1716));
    layer2_outputs(1138) <= not(layer1_outputs(460)) or (layer1_outputs(3999));
    layer2_outputs(1139) <= not((layer1_outputs(3081)) and (layer1_outputs(2448)));
    layer2_outputs(1140) <= not((layer1_outputs(337)) and (layer1_outputs(4423)));
    layer2_outputs(1141) <= (layer1_outputs(6104)) and (layer1_outputs(4586));
    layer2_outputs(1142) <= '0';
    layer2_outputs(1143) <= not((layer1_outputs(7313)) or (layer1_outputs(1483)));
    layer2_outputs(1144) <= '1';
    layer2_outputs(1145) <= (layer1_outputs(1549)) and not (layer1_outputs(6605));
    layer2_outputs(1146) <= not(layer1_outputs(928));
    layer2_outputs(1147) <= (layer1_outputs(151)) and (layer1_outputs(6298));
    layer2_outputs(1148) <= layer1_outputs(992);
    layer2_outputs(1149) <= not((layer1_outputs(3212)) xor (layer1_outputs(2423)));
    layer2_outputs(1150) <= (layer1_outputs(7084)) and not (layer1_outputs(7594));
    layer2_outputs(1151) <= not(layer1_outputs(6152)) or (layer1_outputs(1388));
    layer2_outputs(1152) <= layer1_outputs(4430);
    layer2_outputs(1153) <= not(layer1_outputs(1947)) or (layer1_outputs(5976));
    layer2_outputs(1154) <= '0';
    layer2_outputs(1155) <= layer1_outputs(4040);
    layer2_outputs(1156) <= not((layer1_outputs(399)) or (layer1_outputs(3823)));
    layer2_outputs(1157) <= (layer1_outputs(2158)) or (layer1_outputs(6267));
    layer2_outputs(1158) <= not(layer1_outputs(7304)) or (layer1_outputs(2381));
    layer2_outputs(1159) <= layer1_outputs(2253);
    layer2_outputs(1160) <= '0';
    layer2_outputs(1161) <= (layer1_outputs(368)) and not (layer1_outputs(4428));
    layer2_outputs(1162) <= not((layer1_outputs(1489)) or (layer1_outputs(2100)));
    layer2_outputs(1163) <= layer1_outputs(181);
    layer2_outputs(1164) <= (layer1_outputs(558)) or (layer1_outputs(6047));
    layer2_outputs(1165) <= not(layer1_outputs(3884));
    layer2_outputs(1166) <= (layer1_outputs(926)) and (layer1_outputs(4092));
    layer2_outputs(1167) <= (layer1_outputs(3568)) and (layer1_outputs(1491));
    layer2_outputs(1168) <= not((layer1_outputs(1519)) or (layer1_outputs(6515)));
    layer2_outputs(1169) <= not((layer1_outputs(6546)) and (layer1_outputs(2948)));
    layer2_outputs(1170) <= (layer1_outputs(2316)) and not (layer1_outputs(6313));
    layer2_outputs(1171) <= layer1_outputs(4341);
    layer2_outputs(1172) <= (layer1_outputs(4067)) xor (layer1_outputs(3541));
    layer2_outputs(1173) <= not(layer1_outputs(173)) or (layer1_outputs(729));
    layer2_outputs(1174) <= (layer1_outputs(7651)) and not (layer1_outputs(1803));
    layer2_outputs(1175) <= layer1_outputs(2951);
    layer2_outputs(1176) <= not(layer1_outputs(4711));
    layer2_outputs(1177) <= not(layer1_outputs(5314)) or (layer1_outputs(4719));
    layer2_outputs(1178) <= not(layer1_outputs(1925)) or (layer1_outputs(7460));
    layer2_outputs(1179) <= not((layer1_outputs(2018)) and (layer1_outputs(7071)));
    layer2_outputs(1180) <= '0';
    layer2_outputs(1181) <= '1';
    layer2_outputs(1182) <= '0';
    layer2_outputs(1183) <= '1';
    layer2_outputs(1184) <= '0';
    layer2_outputs(1185) <= (layer1_outputs(3133)) and not (layer1_outputs(7189));
    layer2_outputs(1186) <= not(layer1_outputs(6985));
    layer2_outputs(1187) <= (layer1_outputs(1019)) and not (layer1_outputs(7554));
    layer2_outputs(1188) <= not(layer1_outputs(426));
    layer2_outputs(1189) <= layer1_outputs(6907);
    layer2_outputs(1190) <= not(layer1_outputs(4243));
    layer2_outputs(1191) <= '1';
    layer2_outputs(1192) <= not(layer1_outputs(669)) or (layer1_outputs(1324));
    layer2_outputs(1193) <= layer1_outputs(6950);
    layer2_outputs(1194) <= '0';
    layer2_outputs(1195) <= (layer1_outputs(5691)) or (layer1_outputs(3130));
    layer2_outputs(1196) <= not((layer1_outputs(2816)) and (layer1_outputs(5058)));
    layer2_outputs(1197) <= not(layer1_outputs(3367));
    layer2_outputs(1198) <= not(layer1_outputs(2661));
    layer2_outputs(1199) <= not(layer1_outputs(4958)) or (layer1_outputs(1961));
    layer2_outputs(1200) <= (layer1_outputs(3044)) or (layer1_outputs(2144));
    layer2_outputs(1201) <= (layer1_outputs(6732)) or (layer1_outputs(6942));
    layer2_outputs(1202) <= not(layer1_outputs(6704));
    layer2_outputs(1203) <= not((layer1_outputs(5590)) or (layer1_outputs(791)));
    layer2_outputs(1204) <= (layer1_outputs(3380)) and not (layer1_outputs(6635));
    layer2_outputs(1205) <= '1';
    layer2_outputs(1206) <= not((layer1_outputs(5953)) or (layer1_outputs(332)));
    layer2_outputs(1207) <= not((layer1_outputs(7616)) or (layer1_outputs(6405)));
    layer2_outputs(1208) <= layer1_outputs(222);
    layer2_outputs(1209) <= not((layer1_outputs(7070)) and (layer1_outputs(4661)));
    layer2_outputs(1210) <= (layer1_outputs(7337)) and (layer1_outputs(5160));
    layer2_outputs(1211) <= (layer1_outputs(2545)) and not (layer1_outputs(1851));
    layer2_outputs(1212) <= layer1_outputs(3069);
    layer2_outputs(1213) <= not(layer1_outputs(5414));
    layer2_outputs(1214) <= layer1_outputs(3838);
    layer2_outputs(1215) <= not((layer1_outputs(3144)) and (layer1_outputs(1518)));
    layer2_outputs(1216) <= '1';
    layer2_outputs(1217) <= (layer1_outputs(3682)) and not (layer1_outputs(3404));
    layer2_outputs(1218) <= not((layer1_outputs(1698)) xor (layer1_outputs(4410)));
    layer2_outputs(1219) <= layer1_outputs(4775);
    layer2_outputs(1220) <= not(layer1_outputs(2391));
    layer2_outputs(1221) <= not((layer1_outputs(6938)) xor (layer1_outputs(7513)));
    layer2_outputs(1222) <= layer1_outputs(6155);
    layer2_outputs(1223) <= not(layer1_outputs(1800));
    layer2_outputs(1224) <= (layer1_outputs(7254)) and (layer1_outputs(5543));
    layer2_outputs(1225) <= (layer1_outputs(3767)) or (layer1_outputs(500));
    layer2_outputs(1226) <= layer1_outputs(363);
    layer2_outputs(1227) <= not(layer1_outputs(3205)) or (layer1_outputs(4282));
    layer2_outputs(1228) <= '1';
    layer2_outputs(1229) <= not(layer1_outputs(4082));
    layer2_outputs(1230) <= not(layer1_outputs(2386));
    layer2_outputs(1231) <= not(layer1_outputs(5777)) or (layer1_outputs(1585));
    layer2_outputs(1232) <= (layer1_outputs(6301)) or (layer1_outputs(2754));
    layer2_outputs(1233) <= (layer1_outputs(2933)) and not (layer1_outputs(156));
    layer2_outputs(1234) <= '1';
    layer2_outputs(1235) <= not(layer1_outputs(4874));
    layer2_outputs(1236) <= (layer1_outputs(1744)) and not (layer1_outputs(1034));
    layer2_outputs(1237) <= (layer1_outputs(3186)) and not (layer1_outputs(1484));
    layer2_outputs(1238) <= (layer1_outputs(4741)) and (layer1_outputs(1190));
    layer2_outputs(1239) <= not((layer1_outputs(2448)) and (layer1_outputs(3364)));
    layer2_outputs(1240) <= not(layer1_outputs(2087));
    layer2_outputs(1241) <= layer1_outputs(3240);
    layer2_outputs(1242) <= '1';
    layer2_outputs(1243) <= (layer1_outputs(7052)) and (layer1_outputs(2401));
    layer2_outputs(1244) <= not(layer1_outputs(532));
    layer2_outputs(1245) <= not((layer1_outputs(5314)) or (layer1_outputs(2771)));
    layer2_outputs(1246) <= not((layer1_outputs(5400)) or (layer1_outputs(6074)));
    layer2_outputs(1247) <= not((layer1_outputs(5594)) or (layer1_outputs(2202)));
    layer2_outputs(1248) <= '1';
    layer2_outputs(1249) <= not(layer1_outputs(6921)) or (layer1_outputs(7029));
    layer2_outputs(1250) <= not((layer1_outputs(5069)) or (layer1_outputs(1543)));
    layer2_outputs(1251) <= not((layer1_outputs(6662)) or (layer1_outputs(4373)));
    layer2_outputs(1252) <= '1';
    layer2_outputs(1253) <= not(layer1_outputs(2562)) or (layer1_outputs(4219));
    layer2_outputs(1254) <= (layer1_outputs(3587)) and not (layer1_outputs(2409));
    layer2_outputs(1255) <= (layer1_outputs(6899)) and not (layer1_outputs(4445));
    layer2_outputs(1256) <= not(layer1_outputs(3963));
    layer2_outputs(1257) <= layer1_outputs(6334);
    layer2_outputs(1258) <= not(layer1_outputs(3910)) or (layer1_outputs(3301));
    layer2_outputs(1259) <= (layer1_outputs(5606)) or (layer1_outputs(7089));
    layer2_outputs(1260) <= not((layer1_outputs(6358)) or (layer1_outputs(2168)));
    layer2_outputs(1261) <= not(layer1_outputs(2069));
    layer2_outputs(1262) <= '0';
    layer2_outputs(1263) <= not(layer1_outputs(4513)) or (layer1_outputs(2067));
    layer2_outputs(1264) <= not((layer1_outputs(7555)) and (layer1_outputs(1648)));
    layer2_outputs(1265) <= (layer1_outputs(1817)) and not (layer1_outputs(1839));
    layer2_outputs(1266) <= (layer1_outputs(6599)) and (layer1_outputs(6187));
    layer2_outputs(1267) <= not(layer1_outputs(5969));
    layer2_outputs(1268) <= '1';
    layer2_outputs(1269) <= not((layer1_outputs(1862)) or (layer1_outputs(1134)));
    layer2_outputs(1270) <= '0';
    layer2_outputs(1271) <= not(layer1_outputs(1824));
    layer2_outputs(1272) <= layer1_outputs(7245);
    layer2_outputs(1273) <= '1';
    layer2_outputs(1274) <= '1';
    layer2_outputs(1275) <= not((layer1_outputs(3878)) or (layer1_outputs(4832)));
    layer2_outputs(1276) <= not(layer1_outputs(4266));
    layer2_outputs(1277) <= not(layer1_outputs(1844)) or (layer1_outputs(717));
    layer2_outputs(1278) <= layer1_outputs(2907);
    layer2_outputs(1279) <= (layer1_outputs(4756)) or (layer1_outputs(405));
    layer2_outputs(1280) <= layer1_outputs(6501);
    layer2_outputs(1281) <= not(layer1_outputs(5744));
    layer2_outputs(1282) <= layer1_outputs(5259);
    layer2_outputs(1283) <= (layer1_outputs(6001)) and (layer1_outputs(4572));
    layer2_outputs(1284) <= not(layer1_outputs(5834)) or (layer1_outputs(1612));
    layer2_outputs(1285) <= layer1_outputs(6463);
    layer2_outputs(1286) <= not(layer1_outputs(5975));
    layer2_outputs(1287) <= (layer1_outputs(7022)) and not (layer1_outputs(2187));
    layer2_outputs(1288) <= '0';
    layer2_outputs(1289) <= layer1_outputs(4398);
    layer2_outputs(1290) <= not((layer1_outputs(4739)) or (layer1_outputs(2009)));
    layer2_outputs(1291) <= '0';
    layer2_outputs(1292) <= not((layer1_outputs(464)) and (layer1_outputs(3983)));
    layer2_outputs(1293) <= not(layer1_outputs(2259)) or (layer1_outputs(472));
    layer2_outputs(1294) <= not((layer1_outputs(104)) or (layer1_outputs(2185)));
    layer2_outputs(1295) <= '1';
    layer2_outputs(1296) <= layer1_outputs(4681);
    layer2_outputs(1297) <= not(layer1_outputs(5980));
    layer2_outputs(1298) <= '1';
    layer2_outputs(1299) <= layer1_outputs(3645);
    layer2_outputs(1300) <= not(layer1_outputs(1168));
    layer2_outputs(1301) <= (layer1_outputs(3263)) and not (layer1_outputs(6719));
    layer2_outputs(1302) <= not(layer1_outputs(6884));
    layer2_outputs(1303) <= not((layer1_outputs(1922)) and (layer1_outputs(235)));
    layer2_outputs(1304) <= not((layer1_outputs(1140)) or (layer1_outputs(5653)));
    layer2_outputs(1305) <= not(layer1_outputs(5683));
    layer2_outputs(1306) <= not((layer1_outputs(7618)) or (layer1_outputs(7077)));
    layer2_outputs(1307) <= layer1_outputs(6360);
    layer2_outputs(1308) <= (layer1_outputs(5225)) and (layer1_outputs(4961));
    layer2_outputs(1309) <= not(layer1_outputs(1299));
    layer2_outputs(1310) <= not(layer1_outputs(6746));
    layer2_outputs(1311) <= (layer1_outputs(4356)) and not (layer1_outputs(5340));
    layer2_outputs(1312) <= (layer1_outputs(7326)) and not (layer1_outputs(3538));
    layer2_outputs(1313) <= (layer1_outputs(4073)) and not (layer1_outputs(5840));
    layer2_outputs(1314) <= (layer1_outputs(2051)) and (layer1_outputs(4468));
    layer2_outputs(1315) <= not(layer1_outputs(1526));
    layer2_outputs(1316) <= layer1_outputs(1059);
    layer2_outputs(1317) <= (layer1_outputs(3862)) or (layer1_outputs(7534));
    layer2_outputs(1318) <= not(layer1_outputs(2259)) or (layer1_outputs(4257));
    layer2_outputs(1319) <= (layer1_outputs(7263)) and not (layer1_outputs(910));
    layer2_outputs(1320) <= (layer1_outputs(5215)) and not (layer1_outputs(4086));
    layer2_outputs(1321) <= '1';
    layer2_outputs(1322) <= '1';
    layer2_outputs(1323) <= (layer1_outputs(7484)) and (layer1_outputs(6760));
    layer2_outputs(1324) <= layer1_outputs(5004);
    layer2_outputs(1325) <= layer1_outputs(2633);
    layer2_outputs(1326) <= '1';
    layer2_outputs(1327) <= not(layer1_outputs(2882)) or (layer1_outputs(3662));
    layer2_outputs(1328) <= layer1_outputs(7632);
    layer2_outputs(1329) <= not(layer1_outputs(4986)) or (layer1_outputs(277));
    layer2_outputs(1330) <= (layer1_outputs(3726)) or (layer1_outputs(7193));
    layer2_outputs(1331) <= not((layer1_outputs(4979)) and (layer1_outputs(835)));
    layer2_outputs(1332) <= (layer1_outputs(7061)) or (layer1_outputs(4052));
    layer2_outputs(1333) <= layer1_outputs(3460);
    layer2_outputs(1334) <= '1';
    layer2_outputs(1335) <= not(layer1_outputs(6854)) or (layer1_outputs(1873));
    layer2_outputs(1336) <= layer1_outputs(347);
    layer2_outputs(1337) <= '1';
    layer2_outputs(1338) <= layer1_outputs(4632);
    layer2_outputs(1339) <= (layer1_outputs(971)) and not (layer1_outputs(4341));
    layer2_outputs(1340) <= not((layer1_outputs(6793)) or (layer1_outputs(2421)));
    layer2_outputs(1341) <= not(layer1_outputs(6012));
    layer2_outputs(1342) <= (layer1_outputs(6077)) and not (layer1_outputs(6187));
    layer2_outputs(1343) <= not(layer1_outputs(3868)) or (layer1_outputs(7436));
    layer2_outputs(1344) <= not(layer1_outputs(5274));
    layer2_outputs(1345) <= not(layer1_outputs(6018)) or (layer1_outputs(279));
    layer2_outputs(1346) <= not((layer1_outputs(4869)) or (layer1_outputs(187)));
    layer2_outputs(1347) <= (layer1_outputs(6959)) or (layer1_outputs(960));
    layer2_outputs(1348) <= layer1_outputs(5406);
    layer2_outputs(1349) <= layer1_outputs(5229);
    layer2_outputs(1350) <= layer1_outputs(5663);
    layer2_outputs(1351) <= (layer1_outputs(2286)) and not (layer1_outputs(4306));
    layer2_outputs(1352) <= not((layer1_outputs(6790)) or (layer1_outputs(1299)));
    layer2_outputs(1353) <= not((layer1_outputs(4521)) or (layer1_outputs(5809)));
    layer2_outputs(1354) <= '0';
    layer2_outputs(1355) <= (layer1_outputs(6745)) or (layer1_outputs(2220));
    layer2_outputs(1356) <= not(layer1_outputs(1961)) or (layer1_outputs(4455));
    layer2_outputs(1357) <= not(layer1_outputs(2182));
    layer2_outputs(1358) <= layer1_outputs(3363);
    layer2_outputs(1359) <= not(layer1_outputs(2737));
    layer2_outputs(1360) <= '0';
    layer2_outputs(1361) <= (layer1_outputs(236)) or (layer1_outputs(7489));
    layer2_outputs(1362) <= not(layer1_outputs(1769)) or (layer1_outputs(6008));
    layer2_outputs(1363) <= not(layer1_outputs(47));
    layer2_outputs(1364) <= not((layer1_outputs(239)) or (layer1_outputs(3876)));
    layer2_outputs(1365) <= not(layer1_outputs(2328)) or (layer1_outputs(1280));
    layer2_outputs(1366) <= layer1_outputs(3220);
    layer2_outputs(1367) <= layer1_outputs(3113);
    layer2_outputs(1368) <= layer1_outputs(6900);
    layer2_outputs(1369) <= not(layer1_outputs(6929));
    layer2_outputs(1370) <= (layer1_outputs(3958)) and not (layer1_outputs(1332));
    layer2_outputs(1371) <= layer1_outputs(1495);
    layer2_outputs(1372) <= not((layer1_outputs(7259)) or (layer1_outputs(872)));
    layer2_outputs(1373) <= layer1_outputs(1727);
    layer2_outputs(1374) <= not((layer1_outputs(2043)) or (layer1_outputs(2178)));
    layer2_outputs(1375) <= not((layer1_outputs(6026)) or (layer1_outputs(3343)));
    layer2_outputs(1376) <= not(layer1_outputs(3325));
    layer2_outputs(1377) <= (layer1_outputs(2064)) or (layer1_outputs(551));
    layer2_outputs(1378) <= (layer1_outputs(5239)) and (layer1_outputs(6218));
    layer2_outputs(1379) <= not(layer1_outputs(6363)) or (layer1_outputs(2625));
    layer2_outputs(1380) <= not(layer1_outputs(5403));
    layer2_outputs(1381) <= '1';
    layer2_outputs(1382) <= (layer1_outputs(5875)) or (layer1_outputs(4552));
    layer2_outputs(1383) <= not((layer1_outputs(2108)) and (layer1_outputs(5580)));
    layer2_outputs(1384) <= not((layer1_outputs(6787)) or (layer1_outputs(6217)));
    layer2_outputs(1385) <= '0';
    layer2_outputs(1386) <= '0';
    layer2_outputs(1387) <= not((layer1_outputs(1825)) or (layer1_outputs(747)));
    layer2_outputs(1388) <= (layer1_outputs(5012)) or (layer1_outputs(2456));
    layer2_outputs(1389) <= (layer1_outputs(1730)) or (layer1_outputs(6574));
    layer2_outputs(1390) <= not((layer1_outputs(5664)) and (layer1_outputs(2318)));
    layer2_outputs(1391) <= '1';
    layer2_outputs(1392) <= not(layer1_outputs(6641));
    layer2_outputs(1393) <= (layer1_outputs(7449)) and not (layer1_outputs(2346));
    layer2_outputs(1394) <= (layer1_outputs(1053)) and (layer1_outputs(906));
    layer2_outputs(1395) <= '1';
    layer2_outputs(1396) <= not(layer1_outputs(1211)) or (layer1_outputs(4805));
    layer2_outputs(1397) <= '0';
    layer2_outputs(1398) <= layer1_outputs(4985);
    layer2_outputs(1399) <= layer1_outputs(6997);
    layer2_outputs(1400) <= layer1_outputs(654);
    layer2_outputs(1401) <= layer1_outputs(208);
    layer2_outputs(1402) <= not(layer1_outputs(631)) or (layer1_outputs(1210));
    layer2_outputs(1403) <= (layer1_outputs(992)) and not (layer1_outputs(5449));
    layer2_outputs(1404) <= not(layer1_outputs(3407));
    layer2_outputs(1405) <= not((layer1_outputs(4043)) or (layer1_outputs(4081)));
    layer2_outputs(1406) <= not(layer1_outputs(386)) or (layer1_outputs(1184));
    layer2_outputs(1407) <= not((layer1_outputs(5339)) or (layer1_outputs(4206)));
    layer2_outputs(1408) <= not(layer1_outputs(2721)) or (layer1_outputs(2899));
    layer2_outputs(1409) <= not((layer1_outputs(533)) or (layer1_outputs(2028)));
    layer2_outputs(1410) <= layer1_outputs(2106);
    layer2_outputs(1411) <= not((layer1_outputs(1789)) and (layer1_outputs(6875)));
    layer2_outputs(1412) <= not(layer1_outputs(3761));
    layer2_outputs(1413) <= layer1_outputs(2140);
    layer2_outputs(1414) <= '0';
    layer2_outputs(1415) <= not(layer1_outputs(2258));
    layer2_outputs(1416) <= not(layer1_outputs(1941)) or (layer1_outputs(2701));
    layer2_outputs(1417) <= not(layer1_outputs(5670));
    layer2_outputs(1418) <= not((layer1_outputs(5848)) and (layer1_outputs(6661)));
    layer2_outputs(1419) <= (layer1_outputs(1681)) and not (layer1_outputs(7024));
    layer2_outputs(1420) <= layer1_outputs(5154);
    layer2_outputs(1421) <= not((layer1_outputs(3488)) or (layer1_outputs(2975)));
    layer2_outputs(1422) <= not(layer1_outputs(7529));
    layer2_outputs(1423) <= not(layer1_outputs(6236));
    layer2_outputs(1424) <= not((layer1_outputs(3036)) or (layer1_outputs(2766)));
    layer2_outputs(1425) <= (layer1_outputs(4946)) and not (layer1_outputs(4554));
    layer2_outputs(1426) <= layer1_outputs(7208);
    layer2_outputs(1427) <= not(layer1_outputs(6870));
    layer2_outputs(1428) <= layer1_outputs(5249);
    layer2_outputs(1429) <= (layer1_outputs(417)) or (layer1_outputs(2486));
    layer2_outputs(1430) <= layer1_outputs(598);
    layer2_outputs(1431) <= (layer1_outputs(6288)) or (layer1_outputs(846));
    layer2_outputs(1432) <= not(layer1_outputs(1831)) or (layer1_outputs(6926));
    layer2_outputs(1433) <= '1';
    layer2_outputs(1434) <= not(layer1_outputs(5090)) or (layer1_outputs(4538));
    layer2_outputs(1435) <= not((layer1_outputs(442)) and (layer1_outputs(7014)));
    layer2_outputs(1436) <= not(layer1_outputs(1620));
    layer2_outputs(1437) <= not((layer1_outputs(521)) or (layer1_outputs(1558)));
    layer2_outputs(1438) <= (layer1_outputs(947)) or (layer1_outputs(4155));
    layer2_outputs(1439) <= (layer1_outputs(3644)) or (layer1_outputs(2575));
    layer2_outputs(1440) <= not(layer1_outputs(4507)) or (layer1_outputs(6149));
    layer2_outputs(1441) <= not(layer1_outputs(4709));
    layer2_outputs(1442) <= layer1_outputs(2341);
    layer2_outputs(1443) <= layer1_outputs(7533);
    layer2_outputs(1444) <= (layer1_outputs(6599)) or (layer1_outputs(1146));
    layer2_outputs(1445) <= (layer1_outputs(404)) xor (layer1_outputs(3350));
    layer2_outputs(1446) <= not((layer1_outputs(3082)) or (layer1_outputs(7640)));
    layer2_outputs(1447) <= not(layer1_outputs(3558)) or (layer1_outputs(5437));
    layer2_outputs(1448) <= not((layer1_outputs(1875)) and (layer1_outputs(5637)));
    layer2_outputs(1449) <= (layer1_outputs(5061)) and not (layer1_outputs(4906));
    layer2_outputs(1450) <= (layer1_outputs(4009)) and (layer1_outputs(579));
    layer2_outputs(1451) <= layer1_outputs(5990);
    layer2_outputs(1452) <= layer1_outputs(3139);
    layer2_outputs(1453) <= layer1_outputs(3015);
    layer2_outputs(1454) <= not(layer1_outputs(441));
    layer2_outputs(1455) <= '1';
    layer2_outputs(1456) <= layer1_outputs(1074);
    layer2_outputs(1457) <= not(layer1_outputs(5537));
    layer2_outputs(1458) <= (layer1_outputs(1528)) or (layer1_outputs(1470));
    layer2_outputs(1459) <= (layer1_outputs(7231)) and not (layer1_outputs(5686));
    layer2_outputs(1460) <= layer1_outputs(1001);
    layer2_outputs(1461) <= '0';
    layer2_outputs(1462) <= layer1_outputs(6987);
    layer2_outputs(1463) <= '1';
    layer2_outputs(1464) <= not(layer1_outputs(7388)) or (layer1_outputs(6604));
    layer2_outputs(1465) <= not(layer1_outputs(4668));
    layer2_outputs(1466) <= not(layer1_outputs(7257));
    layer2_outputs(1467) <= not(layer1_outputs(6231));
    layer2_outputs(1468) <= not((layer1_outputs(3294)) or (layer1_outputs(1310)));
    layer2_outputs(1469) <= not(layer1_outputs(1880));
    layer2_outputs(1470) <= layer1_outputs(2463);
    layer2_outputs(1471) <= layer1_outputs(4820);
    layer2_outputs(1472) <= (layer1_outputs(2224)) and (layer1_outputs(2805));
    layer2_outputs(1473) <= (layer1_outputs(1042)) and (layer1_outputs(1060));
    layer2_outputs(1474) <= layer1_outputs(4737);
    layer2_outputs(1475) <= (layer1_outputs(281)) and not (layer1_outputs(6176));
    layer2_outputs(1476) <= not((layer1_outputs(7222)) or (layer1_outputs(1550)));
    layer2_outputs(1477) <= not(layer1_outputs(377));
    layer2_outputs(1478) <= not((layer1_outputs(5148)) and (layer1_outputs(7582)));
    layer2_outputs(1479) <= not(layer1_outputs(3698));
    layer2_outputs(1480) <= (layer1_outputs(4753)) and (layer1_outputs(818));
    layer2_outputs(1481) <= (layer1_outputs(7526)) and not (layer1_outputs(436));
    layer2_outputs(1482) <= layer1_outputs(144);
    layer2_outputs(1483) <= not(layer1_outputs(6726));
    layer2_outputs(1484) <= not(layer1_outputs(5871));
    layer2_outputs(1485) <= (layer1_outputs(3467)) and (layer1_outputs(5583));
    layer2_outputs(1486) <= layer1_outputs(6211);
    layer2_outputs(1487) <= not(layer1_outputs(6419));
    layer2_outputs(1488) <= (layer1_outputs(4096)) and (layer1_outputs(7553));
    layer2_outputs(1489) <= not(layer1_outputs(2085));
    layer2_outputs(1490) <= not(layer1_outputs(3907));
    layer2_outputs(1491) <= not((layer1_outputs(6880)) and (layer1_outputs(6432)));
    layer2_outputs(1492) <= not((layer1_outputs(2312)) or (layer1_outputs(302)));
    layer2_outputs(1493) <= not(layer1_outputs(5075)) or (layer1_outputs(595));
    layer2_outputs(1494) <= layer1_outputs(2665);
    layer2_outputs(1495) <= '1';
    layer2_outputs(1496) <= not((layer1_outputs(3961)) and (layer1_outputs(171)));
    layer2_outputs(1497) <= (layer1_outputs(2572)) xor (layer1_outputs(127));
    layer2_outputs(1498) <= (layer1_outputs(5321)) and not (layer1_outputs(4524));
    layer2_outputs(1499) <= not(layer1_outputs(1656)) or (layer1_outputs(4637));
    layer2_outputs(1500) <= not(layer1_outputs(4626)) or (layer1_outputs(1037));
    layer2_outputs(1501) <= layer1_outputs(1487);
    layer2_outputs(1502) <= (layer1_outputs(5801)) or (layer1_outputs(5649));
    layer2_outputs(1503) <= not(layer1_outputs(4720)) or (layer1_outputs(670));
    layer2_outputs(1504) <= not((layer1_outputs(1010)) or (layer1_outputs(2402)));
    layer2_outputs(1505) <= '0';
    layer2_outputs(1506) <= (layer1_outputs(2903)) xor (layer1_outputs(100));
    layer2_outputs(1507) <= '1';
    layer2_outputs(1508) <= not(layer1_outputs(785));
    layer2_outputs(1509) <= (layer1_outputs(2909)) or (layer1_outputs(1192));
    layer2_outputs(1510) <= not((layer1_outputs(3861)) and (layer1_outputs(4569)));
    layer2_outputs(1511) <= (layer1_outputs(5564)) and not (layer1_outputs(5584));
    layer2_outputs(1512) <= not((layer1_outputs(4461)) and (layer1_outputs(5940)));
    layer2_outputs(1513) <= layer1_outputs(486);
    layer2_outputs(1514) <= '1';
    layer2_outputs(1515) <= layer1_outputs(303);
    layer2_outputs(1516) <= layer1_outputs(6168);
    layer2_outputs(1517) <= not(layer1_outputs(3672)) or (layer1_outputs(2283));
    layer2_outputs(1518) <= '0';
    layer2_outputs(1519) <= (layer1_outputs(5876)) and not (layer1_outputs(3976));
    layer2_outputs(1520) <= not(layer1_outputs(3053));
    layer2_outputs(1521) <= not(layer1_outputs(2339)) or (layer1_outputs(4129));
    layer2_outputs(1522) <= layer1_outputs(1900);
    layer2_outputs(1523) <= not(layer1_outputs(2071));
    layer2_outputs(1524) <= (layer1_outputs(258)) and not (layer1_outputs(172));
    layer2_outputs(1525) <= (layer1_outputs(3602)) and not (layer1_outputs(5344));
    layer2_outputs(1526) <= not(layer1_outputs(1753));
    layer2_outputs(1527) <= (layer1_outputs(5659)) and not (layer1_outputs(5049));
    layer2_outputs(1528) <= not(layer1_outputs(360)) or (layer1_outputs(3731));
    layer2_outputs(1529) <= not((layer1_outputs(7367)) or (layer1_outputs(2556)));
    layer2_outputs(1530) <= not(layer1_outputs(3717)) or (layer1_outputs(7332));
    layer2_outputs(1531) <= not(layer1_outputs(4875)) or (layer1_outputs(3157));
    layer2_outputs(1532) <= not(layer1_outputs(1705)) or (layer1_outputs(3682));
    layer2_outputs(1533) <= layer1_outputs(1734);
    layer2_outputs(1534) <= not(layer1_outputs(6048));
    layer2_outputs(1535) <= not((layer1_outputs(6886)) or (layer1_outputs(6797)));
    layer2_outputs(1536) <= not(layer1_outputs(2731)) or (layer1_outputs(4456));
    layer2_outputs(1537) <= (layer1_outputs(5068)) and (layer1_outputs(3676));
    layer2_outputs(1538) <= not(layer1_outputs(2011)) or (layer1_outputs(6618));
    layer2_outputs(1539) <= not(layer1_outputs(279));
    layer2_outputs(1540) <= layer1_outputs(2979);
    layer2_outputs(1541) <= (layer1_outputs(435)) xor (layer1_outputs(7152));
    layer2_outputs(1542) <= (layer1_outputs(5009)) and (layer1_outputs(4697));
    layer2_outputs(1543) <= layer1_outputs(3560);
    layer2_outputs(1544) <= not((layer1_outputs(5255)) and (layer1_outputs(1887)));
    layer2_outputs(1545) <= layer1_outputs(2893);
    layer2_outputs(1546) <= not((layer1_outputs(858)) or (layer1_outputs(3110)));
    layer2_outputs(1547) <= layer1_outputs(6608);
    layer2_outputs(1548) <= '1';
    layer2_outputs(1549) <= not(layer1_outputs(3686)) or (layer1_outputs(2747));
    layer2_outputs(1550) <= '0';
    layer2_outputs(1551) <= not(layer1_outputs(443));
    layer2_outputs(1552) <= (layer1_outputs(6360)) or (layer1_outputs(101));
    layer2_outputs(1553) <= not((layer1_outputs(5578)) and (layer1_outputs(228)));
    layer2_outputs(1554) <= (layer1_outputs(1226)) or (layer1_outputs(6805));
    layer2_outputs(1555) <= (layer1_outputs(2610)) and not (layer1_outputs(2839));
    layer2_outputs(1556) <= '1';
    layer2_outputs(1557) <= not((layer1_outputs(4248)) and (layer1_outputs(2608)));
    layer2_outputs(1558) <= '1';
    layer2_outputs(1559) <= not(layer1_outputs(2095)) or (layer1_outputs(5272));
    layer2_outputs(1560) <= layer1_outputs(6155);
    layer2_outputs(1561) <= (layer1_outputs(5824)) and not (layer1_outputs(1551));
    layer2_outputs(1562) <= (layer1_outputs(5147)) and (layer1_outputs(686));
    layer2_outputs(1563) <= layer1_outputs(3723);
    layer2_outputs(1564) <= (layer1_outputs(4935)) or (layer1_outputs(5264));
    layer2_outputs(1565) <= layer1_outputs(4183);
    layer2_outputs(1566) <= (layer1_outputs(6171)) and not (layer1_outputs(142));
    layer2_outputs(1567) <= (layer1_outputs(7248)) and (layer1_outputs(1361));
    layer2_outputs(1568) <= layer1_outputs(4646);
    layer2_outputs(1569) <= (layer1_outputs(6905)) or (layer1_outputs(260));
    layer2_outputs(1570) <= '0';
    layer2_outputs(1571) <= layer1_outputs(3277);
    layer2_outputs(1572) <= not((layer1_outputs(4333)) xor (layer1_outputs(3873)));
    layer2_outputs(1573) <= not((layer1_outputs(5966)) or (layer1_outputs(3544)));
    layer2_outputs(1574) <= not((layer1_outputs(1792)) and (layer1_outputs(4909)));
    layer2_outputs(1575) <= not(layer1_outputs(4258));
    layer2_outputs(1576) <= (layer1_outputs(2856)) or (layer1_outputs(2039));
    layer2_outputs(1577) <= not((layer1_outputs(1903)) or (layer1_outputs(7579)));
    layer2_outputs(1578) <= not(layer1_outputs(3018));
    layer2_outputs(1579) <= not(layer1_outputs(3041));
    layer2_outputs(1580) <= layer1_outputs(4243);
    layer2_outputs(1581) <= not(layer1_outputs(7628));
    layer2_outputs(1582) <= layer1_outputs(3014);
    layer2_outputs(1583) <= '0';
    layer2_outputs(1584) <= layer1_outputs(7151);
    layer2_outputs(1585) <= not((layer1_outputs(610)) or (layer1_outputs(5254)));
    layer2_outputs(1586) <= layer1_outputs(4109);
    layer2_outputs(1587) <= (layer1_outputs(1359)) and not (layer1_outputs(3769));
    layer2_outputs(1588) <= '0';
    layer2_outputs(1589) <= (layer1_outputs(363)) or (layer1_outputs(7174));
    layer2_outputs(1590) <= (layer1_outputs(5745)) and (layer1_outputs(2294));
    layer2_outputs(1591) <= '0';
    layer2_outputs(1592) <= '0';
    layer2_outputs(1593) <= not(layer1_outputs(4020));
    layer2_outputs(1594) <= not((layer1_outputs(5870)) or (layer1_outputs(5065)));
    layer2_outputs(1595) <= '1';
    layer2_outputs(1596) <= layer1_outputs(3449);
    layer2_outputs(1597) <= '0';
    layer2_outputs(1598) <= not((layer1_outputs(5334)) xor (layer1_outputs(227)));
    layer2_outputs(1599) <= (layer1_outputs(3349)) or (layer1_outputs(2586));
    layer2_outputs(1600) <= '1';
    layer2_outputs(1601) <= layer1_outputs(3093);
    layer2_outputs(1602) <= layer1_outputs(6136);
    layer2_outputs(1603) <= not(layer1_outputs(4300));
    layer2_outputs(1604) <= '0';
    layer2_outputs(1605) <= (layer1_outputs(891)) and (layer1_outputs(2113));
    layer2_outputs(1606) <= '1';
    layer2_outputs(1607) <= layer1_outputs(1639);
    layer2_outputs(1608) <= (layer1_outputs(2459)) and (layer1_outputs(7433));
    layer2_outputs(1609) <= (layer1_outputs(2797)) and (layer1_outputs(5149));
    layer2_outputs(1610) <= not(layer1_outputs(1339));
    layer2_outputs(1611) <= (layer1_outputs(2214)) and not (layer1_outputs(790));
    layer2_outputs(1612) <= not(layer1_outputs(7428));
    layer2_outputs(1613) <= layer1_outputs(1651);
    layer2_outputs(1614) <= (layer1_outputs(5774)) or (layer1_outputs(4138));
    layer2_outputs(1615) <= '0';
    layer2_outputs(1616) <= layer1_outputs(5429);
    layer2_outputs(1617) <= not(layer1_outputs(929)) or (layer1_outputs(4078));
    layer2_outputs(1618) <= layer1_outputs(1302);
    layer2_outputs(1619) <= '1';
    layer2_outputs(1620) <= layer1_outputs(1956);
    layer2_outputs(1621) <= not(layer1_outputs(4849));
    layer2_outputs(1622) <= not(layer1_outputs(3200));
    layer2_outputs(1623) <= (layer1_outputs(6441)) or (layer1_outputs(7443));
    layer2_outputs(1624) <= not(layer1_outputs(2749));
    layer2_outputs(1625) <= not((layer1_outputs(2165)) or (layer1_outputs(6807)));
    layer2_outputs(1626) <= layer1_outputs(4902);
    layer2_outputs(1627) <= not(layer1_outputs(130));
    layer2_outputs(1628) <= layer1_outputs(842);
    layer2_outputs(1629) <= layer1_outputs(5067);
    layer2_outputs(1630) <= (layer1_outputs(3271)) and (layer1_outputs(6983));
    layer2_outputs(1631) <= layer1_outputs(6649);
    layer2_outputs(1632) <= not((layer1_outputs(4124)) or (layer1_outputs(5733)));
    layer2_outputs(1633) <= (layer1_outputs(2640)) xor (layer1_outputs(7678));
    layer2_outputs(1634) <= not(layer1_outputs(685)) or (layer1_outputs(294));
    layer2_outputs(1635) <= (layer1_outputs(3818)) and not (layer1_outputs(868));
    layer2_outputs(1636) <= not((layer1_outputs(741)) or (layer1_outputs(575)));
    layer2_outputs(1637) <= not(layer1_outputs(2128));
    layer2_outputs(1638) <= not(layer1_outputs(7245)) or (layer1_outputs(6086));
    layer2_outputs(1639) <= layer1_outputs(2552);
    layer2_outputs(1640) <= layer1_outputs(902);
    layer2_outputs(1641) <= not(layer1_outputs(650)) or (layer1_outputs(5358));
    layer2_outputs(1642) <= (layer1_outputs(6839)) and (layer1_outputs(5667));
    layer2_outputs(1643) <= not(layer1_outputs(3284)) or (layer1_outputs(2385));
    layer2_outputs(1644) <= layer1_outputs(2720);
    layer2_outputs(1645) <= not((layer1_outputs(4811)) and (layer1_outputs(6214)));
    layer2_outputs(1646) <= '0';
    layer2_outputs(1647) <= (layer1_outputs(5608)) and not (layer1_outputs(4943));
    layer2_outputs(1648) <= (layer1_outputs(1752)) and (layer1_outputs(3609));
    layer2_outputs(1649) <= (layer1_outputs(7531)) and not (layer1_outputs(6202));
    layer2_outputs(1650) <= (layer1_outputs(372)) or (layer1_outputs(5994));
    layer2_outputs(1651) <= '0';
    layer2_outputs(1652) <= '0';
    layer2_outputs(1653) <= not(layer1_outputs(2524)) or (layer1_outputs(6642));
    layer2_outputs(1654) <= layer1_outputs(650);
    layer2_outputs(1655) <= not(layer1_outputs(905)) or (layer1_outputs(326));
    layer2_outputs(1656) <= (layer1_outputs(769)) and (layer1_outputs(6374));
    layer2_outputs(1657) <= (layer1_outputs(1275)) and not (layer1_outputs(2378));
    layer2_outputs(1658) <= not(layer1_outputs(170)) or (layer1_outputs(5379));
    layer2_outputs(1659) <= (layer1_outputs(3078)) and not (layer1_outputs(7528));
    layer2_outputs(1660) <= (layer1_outputs(55)) and not (layer1_outputs(4910));
    layer2_outputs(1661) <= (layer1_outputs(875)) and not (layer1_outputs(3797));
    layer2_outputs(1662) <= layer1_outputs(2399);
    layer2_outputs(1663) <= not(layer1_outputs(3846));
    layer2_outputs(1664) <= not((layer1_outputs(3509)) and (layer1_outputs(6553)));
    layer2_outputs(1665) <= not((layer1_outputs(449)) and (layer1_outputs(6458)));
    layer2_outputs(1666) <= not(layer1_outputs(2197));
    layer2_outputs(1667) <= not((layer1_outputs(3928)) and (layer1_outputs(6584)));
    layer2_outputs(1668) <= layer1_outputs(3778);
    layer2_outputs(1669) <= (layer1_outputs(6869)) or (layer1_outputs(329));
    layer2_outputs(1670) <= '0';
    layer2_outputs(1671) <= not(layer1_outputs(1070)) or (layer1_outputs(512));
    layer2_outputs(1672) <= not(layer1_outputs(5166));
    layer2_outputs(1673) <= '1';
    layer2_outputs(1674) <= not(layer1_outputs(5114));
    layer2_outputs(1675) <= not((layer1_outputs(7556)) and (layer1_outputs(569)));
    layer2_outputs(1676) <= not((layer1_outputs(6242)) xor (layer1_outputs(7605)));
    layer2_outputs(1677) <= (layer1_outputs(3155)) or (layer1_outputs(78));
    layer2_outputs(1678) <= not((layer1_outputs(1859)) and (layer1_outputs(5977)));
    layer2_outputs(1679) <= layer1_outputs(2981);
    layer2_outputs(1680) <= not(layer1_outputs(1337)) or (layer1_outputs(5891));
    layer2_outputs(1681) <= not(layer1_outputs(7253));
    layer2_outputs(1682) <= not(layer1_outputs(1936));
    layer2_outputs(1683) <= not(layer1_outputs(6788));
    layer2_outputs(1684) <= (layer1_outputs(850)) and not (layer1_outputs(7377));
    layer2_outputs(1685) <= not((layer1_outputs(7244)) and (layer1_outputs(3853)));
    layer2_outputs(1686) <= (layer1_outputs(3303)) or (layer1_outputs(5534));
    layer2_outputs(1687) <= not((layer1_outputs(5643)) or (layer1_outputs(2921)));
    layer2_outputs(1688) <= (layer1_outputs(2206)) and not (layer1_outputs(1712));
    layer2_outputs(1689) <= layer1_outputs(1919);
    layer2_outputs(1690) <= '0';
    layer2_outputs(1691) <= (layer1_outputs(6831)) or (layer1_outputs(1289));
    layer2_outputs(1692) <= not((layer1_outputs(5139)) and (layer1_outputs(6901)));
    layer2_outputs(1693) <= not(layer1_outputs(1005));
    layer2_outputs(1694) <= '0';
    layer2_outputs(1695) <= layer1_outputs(7127);
    layer2_outputs(1696) <= (layer1_outputs(4030)) xor (layer1_outputs(3821));
    layer2_outputs(1697) <= not((layer1_outputs(6877)) and (layer1_outputs(3279)));
    layer2_outputs(1698) <= '1';
    layer2_outputs(1699) <= not((layer1_outputs(2453)) and (layer1_outputs(3128)));
    layer2_outputs(1700) <= (layer1_outputs(5540)) and not (layer1_outputs(1172));
    layer2_outputs(1701) <= '1';
    layer2_outputs(1702) <= not(layer1_outputs(1993));
    layer2_outputs(1703) <= layer1_outputs(6287);
    layer2_outputs(1704) <= layer1_outputs(5265);
    layer2_outputs(1705) <= layer1_outputs(254);
    layer2_outputs(1706) <= not((layer1_outputs(2500)) or (layer1_outputs(4136)));
    layer2_outputs(1707) <= not(layer1_outputs(2187));
    layer2_outputs(1708) <= layer1_outputs(529);
    layer2_outputs(1709) <= not((layer1_outputs(5104)) and (layer1_outputs(6210)));
    layer2_outputs(1710) <= not((layer1_outputs(4297)) or (layer1_outputs(6937)));
    layer2_outputs(1711) <= layer1_outputs(6145);
    layer2_outputs(1712) <= not(layer1_outputs(3850)) or (layer1_outputs(4813));
    layer2_outputs(1713) <= '0';
    layer2_outputs(1714) <= '0';
    layer2_outputs(1715) <= '0';
    layer2_outputs(1716) <= layer1_outputs(7079);
    layer2_outputs(1717) <= layer1_outputs(4657);
    layer2_outputs(1718) <= layer1_outputs(7167);
    layer2_outputs(1719) <= not(layer1_outputs(3666)) or (layer1_outputs(108));
    layer2_outputs(1720) <= (layer1_outputs(903)) and not (layer1_outputs(5119));
    layer2_outputs(1721) <= '1';
    layer2_outputs(1722) <= not((layer1_outputs(553)) and (layer1_outputs(4630)));
    layer2_outputs(1723) <= not(layer1_outputs(3076));
    layer2_outputs(1724) <= (layer1_outputs(1205)) and (layer1_outputs(2746));
    layer2_outputs(1725) <= layer1_outputs(2238);
    layer2_outputs(1726) <= not(layer1_outputs(3837)) or (layer1_outputs(1644));
    layer2_outputs(1727) <= layer1_outputs(5792);
    layer2_outputs(1728) <= not((layer1_outputs(5344)) or (layer1_outputs(3524)));
    layer2_outputs(1729) <= not(layer1_outputs(1939));
    layer2_outputs(1730) <= not((layer1_outputs(5093)) and (layer1_outputs(2943)));
    layer2_outputs(1731) <= '0';
    layer2_outputs(1732) <= (layer1_outputs(6101)) or (layer1_outputs(425));
    layer2_outputs(1733) <= layer1_outputs(277);
    layer2_outputs(1734) <= (layer1_outputs(4529)) and not (layer1_outputs(4576));
    layer2_outputs(1735) <= not((layer1_outputs(4851)) or (layer1_outputs(5562)));
    layer2_outputs(1736) <= '0';
    layer2_outputs(1737) <= '0';
    layer2_outputs(1738) <= layer1_outputs(6800);
    layer2_outputs(1739) <= (layer1_outputs(2634)) xor (layer1_outputs(5713));
    layer2_outputs(1740) <= not((layer1_outputs(1237)) or (layer1_outputs(4382)));
    layer2_outputs(1741) <= not(layer1_outputs(3365));
    layer2_outputs(1742) <= not((layer1_outputs(2588)) or (layer1_outputs(5658)));
    layer2_outputs(1743) <= '1';
    layer2_outputs(1744) <= '1';
    layer2_outputs(1745) <= layer1_outputs(3118);
    layer2_outputs(1746) <= '0';
    layer2_outputs(1747) <= layer1_outputs(5152);
    layer2_outputs(1748) <= (layer1_outputs(744)) and not (layer1_outputs(4920));
    layer2_outputs(1749) <= (layer1_outputs(782)) and not (layer1_outputs(3612));
    layer2_outputs(1750) <= '0';
    layer2_outputs(1751) <= not(layer1_outputs(6041)) or (layer1_outputs(1550));
    layer2_outputs(1752) <= '1';
    layer2_outputs(1753) <= layer1_outputs(548);
    layer2_outputs(1754) <= not((layer1_outputs(6396)) xor (layer1_outputs(2490)));
    layer2_outputs(1755) <= (layer1_outputs(2257)) xor (layer1_outputs(4550));
    layer2_outputs(1756) <= not(layer1_outputs(1989)) or (layer1_outputs(867));
    layer2_outputs(1757) <= (layer1_outputs(4380)) and not (layer1_outputs(4385));
    layer2_outputs(1758) <= not(layer1_outputs(4167)) or (layer1_outputs(2279));
    layer2_outputs(1759) <= not((layer1_outputs(6857)) or (layer1_outputs(6716)));
    layer2_outputs(1760) <= not(layer1_outputs(4579));
    layer2_outputs(1761) <= '0';
    layer2_outputs(1762) <= not((layer1_outputs(7435)) or (layer1_outputs(116)));
    layer2_outputs(1763) <= not(layer1_outputs(5991));
    layer2_outputs(1764) <= not(layer1_outputs(7042));
    layer2_outputs(1765) <= layer1_outputs(986);
    layer2_outputs(1766) <= '0';
    layer2_outputs(1767) <= not(layer1_outputs(3478));
    layer2_outputs(1768) <= (layer1_outputs(4192)) or (layer1_outputs(1237));
    layer2_outputs(1769) <= not(layer1_outputs(1054)) or (layer1_outputs(997));
    layer2_outputs(1770) <= not((layer1_outputs(4137)) and (layer1_outputs(6508)));
    layer2_outputs(1771) <= layer1_outputs(1923);
    layer2_outputs(1772) <= layer1_outputs(2793);
    layer2_outputs(1773) <= (layer1_outputs(2634)) and not (layer1_outputs(3481));
    layer2_outputs(1774) <= '1';
    layer2_outputs(1775) <= not(layer1_outputs(1972));
    layer2_outputs(1776) <= (layer1_outputs(525)) and not (layer1_outputs(5246));
    layer2_outputs(1777) <= not(layer1_outputs(5288));
    layer2_outputs(1778) <= not(layer1_outputs(611));
    layer2_outputs(1779) <= not(layer1_outputs(4034));
    layer2_outputs(1780) <= not((layer1_outputs(4705)) and (layer1_outputs(1486)));
    layer2_outputs(1781) <= layer1_outputs(4774);
    layer2_outputs(1782) <= '0';
    layer2_outputs(1783) <= not(layer1_outputs(5528)) or (layer1_outputs(672));
    layer2_outputs(1784) <= not((layer1_outputs(1914)) and (layer1_outputs(1658)));
    layer2_outputs(1785) <= layer1_outputs(1155);
    layer2_outputs(1786) <= layer1_outputs(4613);
    layer2_outputs(1787) <= not(layer1_outputs(4474)) or (layer1_outputs(1384));
    layer2_outputs(1788) <= not((layer1_outputs(5944)) and (layer1_outputs(4730)));
    layer2_outputs(1789) <= '1';
    layer2_outputs(1790) <= '1';
    layer2_outputs(1791) <= '0';
    layer2_outputs(1792) <= not(layer1_outputs(3455));
    layer2_outputs(1793) <= (layer1_outputs(3402)) and not (layer1_outputs(785));
    layer2_outputs(1794) <= (layer1_outputs(6865)) and (layer1_outputs(5686));
    layer2_outputs(1795) <= (layer1_outputs(2253)) or (layer1_outputs(2523));
    layer2_outputs(1796) <= not((layer1_outputs(7438)) or (layer1_outputs(4516)));
    layer2_outputs(1797) <= (layer1_outputs(1102)) and not (layer1_outputs(5255));
    layer2_outputs(1798) <= not((layer1_outputs(5028)) xor (layer1_outputs(6316)));
    layer2_outputs(1799) <= layer1_outputs(3295);
    layer2_outputs(1800) <= '1';
    layer2_outputs(1801) <= not(layer1_outputs(6177));
    layer2_outputs(1802) <= (layer1_outputs(1064)) and not (layer1_outputs(5256));
    layer2_outputs(1803) <= not(layer1_outputs(3971)) or (layer1_outputs(4221));
    layer2_outputs(1804) <= '1';
    layer2_outputs(1805) <= (layer1_outputs(2718)) or (layer1_outputs(3571));
    layer2_outputs(1806) <= (layer1_outputs(5660)) or (layer1_outputs(6388));
    layer2_outputs(1807) <= not(layer1_outputs(2234)) or (layer1_outputs(4343));
    layer2_outputs(1808) <= (layer1_outputs(876)) and (layer1_outputs(3002));
    layer2_outputs(1809) <= layer1_outputs(1515);
    layer2_outputs(1810) <= layer1_outputs(531);
    layer2_outputs(1811) <= (layer1_outputs(27)) and not (layer1_outputs(3346));
    layer2_outputs(1812) <= layer1_outputs(4493);
    layer2_outputs(1813) <= not(layer1_outputs(387)) or (layer1_outputs(231));
    layer2_outputs(1814) <= (layer1_outputs(4024)) and (layer1_outputs(7667));
    layer2_outputs(1815) <= not(layer1_outputs(5710)) or (layer1_outputs(1215));
    layer2_outputs(1816) <= (layer1_outputs(7527)) xor (layer1_outputs(499));
    layer2_outputs(1817) <= not(layer1_outputs(6352));
    layer2_outputs(1818) <= not(layer1_outputs(5309));
    layer2_outputs(1819) <= layer1_outputs(395);
    layer2_outputs(1820) <= '1';
    layer2_outputs(1821) <= (layer1_outputs(2720)) or (layer1_outputs(3773));
    layer2_outputs(1822) <= (layer1_outputs(1990)) and not (layer1_outputs(5261));
    layer2_outputs(1823) <= not((layer1_outputs(2064)) or (layer1_outputs(1309)));
    layer2_outputs(1824) <= not(layer1_outputs(4367)) or (layer1_outputs(7359));
    layer2_outputs(1825) <= not(layer1_outputs(4189));
    layer2_outputs(1826) <= (layer1_outputs(5992)) xor (layer1_outputs(4289));
    layer2_outputs(1827) <= not(layer1_outputs(3441));
    layer2_outputs(1828) <= (layer1_outputs(7054)) and (layer1_outputs(6303));
    layer2_outputs(1829) <= (layer1_outputs(4916)) and (layer1_outputs(419));
    layer2_outputs(1830) <= layer1_outputs(2065);
    layer2_outputs(1831) <= (layer1_outputs(4496)) and (layer1_outputs(4412));
    layer2_outputs(1832) <= layer1_outputs(3574);
    layer2_outputs(1833) <= not(layer1_outputs(2467));
    layer2_outputs(1834) <= (layer1_outputs(4669)) and not (layer1_outputs(2799));
    layer2_outputs(1835) <= not((layer1_outputs(5818)) xor (layer1_outputs(3973)));
    layer2_outputs(1836) <= layer1_outputs(4194);
    layer2_outputs(1837) <= not(layer1_outputs(646));
    layer2_outputs(1838) <= '1';
    layer2_outputs(1839) <= '0';
    layer2_outputs(1840) <= not(layer1_outputs(2347));
    layer2_outputs(1841) <= layer1_outputs(659);
    layer2_outputs(1842) <= '0';
    layer2_outputs(1843) <= '1';
    layer2_outputs(1844) <= not(layer1_outputs(6723)) or (layer1_outputs(7226));
    layer2_outputs(1845) <= not(layer1_outputs(1041)) or (layer1_outputs(3148));
    layer2_outputs(1846) <= not(layer1_outputs(3379)) or (layer1_outputs(4204));
    layer2_outputs(1847) <= not(layer1_outputs(2706)) or (layer1_outputs(467));
    layer2_outputs(1848) <= not(layer1_outputs(7144));
    layer2_outputs(1849) <= not(layer1_outputs(1335));
    layer2_outputs(1850) <= not(layer1_outputs(1954));
    layer2_outputs(1851) <= (layer1_outputs(4594)) and (layer1_outputs(2435));
    layer2_outputs(1852) <= '0';
    layer2_outputs(1853) <= '1';
    layer2_outputs(1854) <= not(layer1_outputs(4449));
    layer2_outputs(1855) <= (layer1_outputs(2331)) and (layer1_outputs(6341));
    layer2_outputs(1856) <= (layer1_outputs(5030)) or (layer1_outputs(7458));
    layer2_outputs(1857) <= layer1_outputs(4992);
    layer2_outputs(1858) <= not(layer1_outputs(5354));
    layer2_outputs(1859) <= (layer1_outputs(5767)) or (layer1_outputs(5233));
    layer2_outputs(1860) <= '1';
    layer2_outputs(1861) <= not(layer1_outputs(3810));
    layer2_outputs(1862) <= layer1_outputs(1436);
    layer2_outputs(1863) <= not(layer1_outputs(1520)) or (layer1_outputs(5104));
    layer2_outputs(1864) <= not(layer1_outputs(1497)) or (layer1_outputs(4598));
    layer2_outputs(1865) <= not(layer1_outputs(4773));
    layer2_outputs(1866) <= not(layer1_outputs(3002)) or (layer1_outputs(2957));
    layer2_outputs(1867) <= not((layer1_outputs(4696)) or (layer1_outputs(3781)));
    layer2_outputs(1868) <= not((layer1_outputs(1203)) or (layer1_outputs(3792)));
    layer2_outputs(1869) <= '0';
    layer2_outputs(1870) <= not((layer1_outputs(7119)) and (layer1_outputs(4322)));
    layer2_outputs(1871) <= not(layer1_outputs(2380));
    layer2_outputs(1872) <= not(layer1_outputs(7622)) or (layer1_outputs(4840));
    layer2_outputs(1873) <= (layer1_outputs(4609)) or (layer1_outputs(2554));
    layer2_outputs(1874) <= layer1_outputs(1996);
    layer2_outputs(1875) <= not(layer1_outputs(6089)) or (layer1_outputs(479));
    layer2_outputs(1876) <= not(layer1_outputs(6294));
    layer2_outputs(1877) <= '1';
    layer2_outputs(1878) <= (layer1_outputs(6348)) and not (layer1_outputs(7294));
    layer2_outputs(1879) <= (layer1_outputs(2157)) and not (layer1_outputs(7272));
    layer2_outputs(1880) <= not(layer1_outputs(6935));
    layer2_outputs(1881) <= not((layer1_outputs(3255)) and (layer1_outputs(3968)));
    layer2_outputs(1882) <= not((layer1_outputs(4069)) or (layer1_outputs(3421)));
    layer2_outputs(1883) <= (layer1_outputs(6348)) and not (layer1_outputs(1333));
    layer2_outputs(1884) <= not((layer1_outputs(5307)) or (layer1_outputs(5365)));
    layer2_outputs(1885) <= '1';
    layer2_outputs(1886) <= not((layer1_outputs(5868)) and (layer1_outputs(2869)));
    layer2_outputs(1887) <= not(layer1_outputs(289)) or (layer1_outputs(6920));
    layer2_outputs(1888) <= not(layer1_outputs(968)) or (layer1_outputs(5627));
    layer2_outputs(1889) <= not(layer1_outputs(4131)) or (layer1_outputs(2458));
    layer2_outputs(1890) <= '0';
    layer2_outputs(1891) <= layer1_outputs(3927);
    layer2_outputs(1892) <= (layer1_outputs(414)) or (layer1_outputs(1011));
    layer2_outputs(1893) <= (layer1_outputs(3796)) and not (layer1_outputs(4801));
    layer2_outputs(1894) <= layer1_outputs(5756);
    layer2_outputs(1895) <= not((layer1_outputs(6878)) or (layer1_outputs(3187)));
    layer2_outputs(1896) <= (layer1_outputs(4803)) and not (layer1_outputs(6759));
    layer2_outputs(1897) <= (layer1_outputs(4142)) or (layer1_outputs(6606));
    layer2_outputs(1898) <= '0';
    layer2_outputs(1899) <= not(layer1_outputs(6147));
    layer2_outputs(1900) <= '0';
    layer2_outputs(1901) <= not(layer1_outputs(5464)) or (layer1_outputs(4944));
    layer2_outputs(1902) <= (layer1_outputs(3461)) or (layer1_outputs(7066));
    layer2_outputs(1903) <= layer1_outputs(7249);
    layer2_outputs(1904) <= not(layer1_outputs(6581)) or (layer1_outputs(4062));
    layer2_outputs(1905) <= '0';
    layer2_outputs(1906) <= '0';
    layer2_outputs(1907) <= layer1_outputs(6987);
    layer2_outputs(1908) <= '0';
    layer2_outputs(1909) <= (layer1_outputs(7516)) and (layer1_outputs(1275));
    layer2_outputs(1910) <= not(layer1_outputs(298));
    layer2_outputs(1911) <= '1';
    layer2_outputs(1912) <= '0';
    layer2_outputs(1913) <= not(layer1_outputs(2806));
    layer2_outputs(1914) <= '0';
    layer2_outputs(1915) <= not((layer1_outputs(5407)) and (layer1_outputs(2419)));
    layer2_outputs(1916) <= '1';
    layer2_outputs(1917) <= layer1_outputs(3014);
    layer2_outputs(1918) <= not(layer1_outputs(6175));
    layer2_outputs(1919) <= not((layer1_outputs(3642)) and (layer1_outputs(3779)));
    layer2_outputs(1920) <= (layer1_outputs(3436)) and not (layer1_outputs(1812));
    layer2_outputs(1921) <= '0';
    layer2_outputs(1922) <= not((layer1_outputs(95)) and (layer1_outputs(45)));
    layer2_outputs(1923) <= not(layer1_outputs(6570)) or (layer1_outputs(300));
    layer2_outputs(1924) <= '0';
    layer2_outputs(1925) <= (layer1_outputs(1823)) and (layer1_outputs(6280));
    layer2_outputs(1926) <= (layer1_outputs(6980)) and not (layer1_outputs(4943));
    layer2_outputs(1927) <= '1';
    layer2_outputs(1928) <= not(layer1_outputs(1352));
    layer2_outputs(1929) <= (layer1_outputs(4702)) and (layer1_outputs(6148));
    layer2_outputs(1930) <= not(layer1_outputs(6071));
    layer2_outputs(1931) <= layer1_outputs(7205);
    layer2_outputs(1932) <= (layer1_outputs(3119)) or (layer1_outputs(1400));
    layer2_outputs(1933) <= not(layer1_outputs(1982));
    layer2_outputs(1934) <= not(layer1_outputs(2155)) or (layer1_outputs(3494));
    layer2_outputs(1935) <= layer1_outputs(6419);
    layer2_outputs(1936) <= (layer1_outputs(217)) or (layer1_outputs(1505));
    layer2_outputs(1937) <= (layer1_outputs(4315)) and (layer1_outputs(3189));
    layer2_outputs(1938) <= not((layer1_outputs(1406)) or (layer1_outputs(511)));
    layer2_outputs(1939) <= layer1_outputs(5975);
    layer2_outputs(1940) <= not(layer1_outputs(1572));
    layer2_outputs(1941) <= layer1_outputs(2464);
    layer2_outputs(1942) <= not(layer1_outputs(4074));
    layer2_outputs(1943) <= layer1_outputs(4091);
    layer2_outputs(1944) <= '0';
    layer2_outputs(1945) <= not(layer1_outputs(2812));
    layer2_outputs(1946) <= not((layer1_outputs(2780)) or (layer1_outputs(213)));
    layer2_outputs(1947) <= not(layer1_outputs(4928));
    layer2_outputs(1948) <= '0';
    layer2_outputs(1949) <= not((layer1_outputs(7575)) or (layer1_outputs(2517)));
    layer2_outputs(1950) <= not(layer1_outputs(6164));
    layer2_outputs(1951) <= '1';
    layer2_outputs(1952) <= not((layer1_outputs(7263)) or (layer1_outputs(2557)));
    layer2_outputs(1953) <= (layer1_outputs(2971)) and not (layer1_outputs(2376));
    layer2_outputs(1954) <= not(layer1_outputs(4389));
    layer2_outputs(1955) <= not((layer1_outputs(1231)) or (layer1_outputs(2049)));
    layer2_outputs(1956) <= (layer1_outputs(2441)) and not (layer1_outputs(4101));
    layer2_outputs(1957) <= layer1_outputs(6241);
    layer2_outputs(1958) <= layer1_outputs(3796);
    layer2_outputs(1959) <= layer1_outputs(660);
    layer2_outputs(1960) <= '1';
    layer2_outputs(1961) <= '1';
    layer2_outputs(1962) <= '0';
    layer2_outputs(1963) <= not(layer1_outputs(2148));
    layer2_outputs(1964) <= layer1_outputs(1856);
    layer2_outputs(1965) <= '1';
    layer2_outputs(1966) <= not(layer1_outputs(5760)) or (layer1_outputs(7670));
    layer2_outputs(1967) <= (layer1_outputs(2611)) xor (layer1_outputs(7131));
    layer2_outputs(1968) <= not(layer1_outputs(7329));
    layer2_outputs(1969) <= (layer1_outputs(5024)) and not (layer1_outputs(7481));
    layer2_outputs(1970) <= not(layer1_outputs(969)) or (layer1_outputs(437));
    layer2_outputs(1971) <= '1';
    layer2_outputs(1972) <= layer1_outputs(5463);
    layer2_outputs(1973) <= (layer1_outputs(4431)) and not (layer1_outputs(3598));
    layer2_outputs(1974) <= not(layer1_outputs(1616)) or (layer1_outputs(3294));
    layer2_outputs(1975) <= not((layer1_outputs(5116)) and (layer1_outputs(6913)));
    layer2_outputs(1976) <= layer1_outputs(5405);
    layer2_outputs(1977) <= not(layer1_outputs(4967));
    layer2_outputs(1978) <= layer1_outputs(5099);
    layer2_outputs(1979) <= not(layer1_outputs(7646)) or (layer1_outputs(3182));
    layer2_outputs(1980) <= not((layer1_outputs(3929)) or (layer1_outputs(5434)));
    layer2_outputs(1981) <= not((layer1_outputs(6786)) or (layer1_outputs(1269)));
    layer2_outputs(1982) <= not(layer1_outputs(6074));
    layer2_outputs(1983) <= '1';
    layer2_outputs(1984) <= (layer1_outputs(385)) and not (layer1_outputs(5731));
    layer2_outputs(1985) <= (layer1_outputs(2198)) or (layer1_outputs(7609));
    layer2_outputs(1986) <= '0';
    layer2_outputs(1987) <= not(layer1_outputs(2769));
    layer2_outputs(1988) <= not(layer1_outputs(6750));
    layer2_outputs(1989) <= not((layer1_outputs(7430)) and (layer1_outputs(4880)));
    layer2_outputs(1990) <= layer1_outputs(6115);
    layer2_outputs(1991) <= layer1_outputs(3762);
    layer2_outputs(1992) <= layer1_outputs(3974);
    layer2_outputs(1993) <= '1';
    layer2_outputs(1994) <= (layer1_outputs(5730)) and not (layer1_outputs(5337));
    layer2_outputs(1995) <= not(layer1_outputs(728));
    layer2_outputs(1996) <= not(layer1_outputs(6196)) or (layer1_outputs(2859));
    layer2_outputs(1997) <= not(layer1_outputs(1305));
    layer2_outputs(1998) <= (layer1_outputs(7340)) and not (layer1_outputs(3775));
    layer2_outputs(1999) <= (layer1_outputs(3172)) or (layer1_outputs(4542));
    layer2_outputs(2000) <= '0';
    layer2_outputs(2001) <= (layer1_outputs(851)) or (layer1_outputs(1793));
    layer2_outputs(2002) <= (layer1_outputs(1177)) and not (layer1_outputs(3984));
    layer2_outputs(2003) <= (layer1_outputs(3592)) or (layer1_outputs(3664));
    layer2_outputs(2004) <= not((layer1_outputs(5300)) xor (layer1_outputs(3779)));
    layer2_outputs(2005) <= layer1_outputs(4311);
    layer2_outputs(2006) <= not(layer1_outputs(6344)) or (layer1_outputs(7000));
    layer2_outputs(2007) <= (layer1_outputs(5639)) and (layer1_outputs(4825));
    layer2_outputs(2008) <= not(layer1_outputs(1123));
    layer2_outputs(2009) <= not(layer1_outputs(6397)) or (layer1_outputs(4301));
    layer2_outputs(2010) <= (layer1_outputs(6388)) or (layer1_outputs(5298));
    layer2_outputs(2011) <= layer1_outputs(6917);
    layer2_outputs(2012) <= layer1_outputs(6709);
    layer2_outputs(2013) <= (layer1_outputs(7179)) and not (layer1_outputs(7182));
    layer2_outputs(2014) <= (layer1_outputs(1216)) and (layer1_outputs(4698));
    layer2_outputs(2015) <= layer1_outputs(3552);
    layer2_outputs(2016) <= not((layer1_outputs(215)) and (layer1_outputs(786)));
    layer2_outputs(2017) <= not((layer1_outputs(5482)) xor (layer1_outputs(6220)));
    layer2_outputs(2018) <= (layer1_outputs(2724)) and not (layer1_outputs(5756));
    layer2_outputs(2019) <= not(layer1_outputs(3209)) or (layer1_outputs(4072));
    layer2_outputs(2020) <= not((layer1_outputs(4274)) and (layer1_outputs(6004)));
    layer2_outputs(2021) <= layer1_outputs(4120);
    layer2_outputs(2022) <= not((layer1_outputs(4539)) or (layer1_outputs(48)));
    layer2_outputs(2023) <= not((layer1_outputs(5503)) or (layer1_outputs(7187)));
    layer2_outputs(2024) <= not(layer1_outputs(2837));
    layer2_outputs(2025) <= (layer1_outputs(578)) and not (layer1_outputs(5016));
    layer2_outputs(2026) <= layer1_outputs(6737);
    layer2_outputs(2027) <= layer1_outputs(687);
    layer2_outputs(2028) <= layer1_outputs(1815);
    layer2_outputs(2029) <= '1';
    layer2_outputs(2030) <= not((layer1_outputs(6225)) and (layer1_outputs(7599)));
    layer2_outputs(2031) <= layer1_outputs(6966);
    layer2_outputs(2032) <= (layer1_outputs(6361)) and not (layer1_outputs(1293));
    layer2_outputs(2033) <= not((layer1_outputs(1981)) and (layer1_outputs(7392)));
    layer2_outputs(2034) <= layer1_outputs(1666);
    layer2_outputs(2035) <= layer1_outputs(1263);
    layer2_outputs(2036) <= layer1_outputs(2343);
    layer2_outputs(2037) <= not(layer1_outputs(1704)) or (layer1_outputs(3101));
    layer2_outputs(2038) <= not(layer1_outputs(3005)) or (layer1_outputs(3256));
    layer2_outputs(2039) <= not((layer1_outputs(4369)) xor (layer1_outputs(5521)));
    layer2_outputs(2040) <= not((layer1_outputs(4122)) or (layer1_outputs(3439)));
    layer2_outputs(2041) <= '0';
    layer2_outputs(2042) <= '0';
    layer2_outputs(2043) <= not(layer1_outputs(7046)) or (layer1_outputs(2493));
    layer2_outputs(2044) <= not((layer1_outputs(1348)) and (layer1_outputs(1476)));
    layer2_outputs(2045) <= not(layer1_outputs(535));
    layer2_outputs(2046) <= '0';
    layer2_outputs(2047) <= (layer1_outputs(523)) and not (layer1_outputs(1936));
    layer2_outputs(2048) <= not(layer1_outputs(2782)) or (layer1_outputs(4922));
    layer2_outputs(2049) <= layer1_outputs(3927);
    layer2_outputs(2050) <= '1';
    layer2_outputs(2051) <= layer1_outputs(5332);
    layer2_outputs(2052) <= layer1_outputs(2247);
    layer2_outputs(2053) <= not(layer1_outputs(2268));
    layer2_outputs(2054) <= (layer1_outputs(1506)) and not (layer1_outputs(7126));
    layer2_outputs(2055) <= (layer1_outputs(688)) or (layer1_outputs(5129));
    layer2_outputs(2056) <= not((layer1_outputs(4847)) or (layer1_outputs(2586)));
    layer2_outputs(2057) <= (layer1_outputs(1326)) and (layer1_outputs(3420));
    layer2_outputs(2058) <= layer1_outputs(3581);
    layer2_outputs(2059) <= '1';
    layer2_outputs(2060) <= layer1_outputs(2436);
    layer2_outputs(2061) <= layer1_outputs(2566);
    layer2_outputs(2062) <= layer1_outputs(5337);
    layer2_outputs(2063) <= (layer1_outputs(225)) or (layer1_outputs(42));
    layer2_outputs(2064) <= not(layer1_outputs(2212)) or (layer1_outputs(5046));
    layer2_outputs(2065) <= not((layer1_outputs(6829)) and (layer1_outputs(4571)));
    layer2_outputs(2066) <= not(layer1_outputs(2426)) or (layer1_outputs(647));
    layer2_outputs(2067) <= layer1_outputs(6479);
    layer2_outputs(2068) <= '1';
    layer2_outputs(2069) <= (layer1_outputs(1252)) xor (layer1_outputs(4393));
    layer2_outputs(2070) <= layer1_outputs(2427);
    layer2_outputs(2071) <= not(layer1_outputs(5506)) or (layer1_outputs(226));
    layer2_outputs(2072) <= (layer1_outputs(3766)) and not (layer1_outputs(3709));
    layer2_outputs(2073) <= not(layer1_outputs(2829)) or (layer1_outputs(2937));
    layer2_outputs(2074) <= (layer1_outputs(2205)) and not (layer1_outputs(6369));
    layer2_outputs(2075) <= not((layer1_outputs(3809)) and (layer1_outputs(6754)));
    layer2_outputs(2076) <= not((layer1_outputs(7658)) and (layer1_outputs(6263)));
    layer2_outputs(2077) <= not(layer1_outputs(3948)) or (layer1_outputs(4193));
    layer2_outputs(2078) <= not((layer1_outputs(6327)) or (layer1_outputs(4409)));
    layer2_outputs(2079) <= not(layer1_outputs(5449));
    layer2_outputs(2080) <= not((layer1_outputs(5582)) or (layer1_outputs(6404)));
    layer2_outputs(2081) <= layer1_outputs(6764);
    layer2_outputs(2082) <= layer1_outputs(683);
    layer2_outputs(2083) <= '0';
    layer2_outputs(2084) <= layer1_outputs(1676);
    layer2_outputs(2085) <= not(layer1_outputs(4654));
    layer2_outputs(2086) <= layer1_outputs(4091);
    layer2_outputs(2087) <= (layer1_outputs(1729)) and not (layer1_outputs(7610));
    layer2_outputs(2088) <= (layer1_outputs(4844)) or (layer1_outputs(6527));
    layer2_outputs(2089) <= not(layer1_outputs(6199));
    layer2_outputs(2090) <= not(layer1_outputs(6107)) or (layer1_outputs(4476));
    layer2_outputs(2091) <= not((layer1_outputs(6361)) or (layer1_outputs(1188)));
    layer2_outputs(2092) <= (layer1_outputs(166)) and not (layer1_outputs(3643));
    layer2_outputs(2093) <= not(layer1_outputs(1097)) or (layer1_outputs(7645));
    layer2_outputs(2094) <= (layer1_outputs(4048)) or (layer1_outputs(7344));
    layer2_outputs(2095) <= (layer1_outputs(4504)) and not (layer1_outputs(5912));
    layer2_outputs(2096) <= (layer1_outputs(2664)) and (layer1_outputs(4606));
    layer2_outputs(2097) <= (layer1_outputs(1635)) or (layer1_outputs(97));
    layer2_outputs(2098) <= not(layer1_outputs(3039));
    layer2_outputs(2099) <= (layer1_outputs(754)) or (layer1_outputs(7117));
    layer2_outputs(2100) <= not(layer1_outputs(4445)) or (layer1_outputs(4628));
    layer2_outputs(2101) <= (layer1_outputs(5604)) and not (layer1_outputs(4088));
    layer2_outputs(2102) <= not(layer1_outputs(1975)) or (layer1_outputs(1200));
    layer2_outputs(2103) <= not(layer1_outputs(6206));
    layer2_outputs(2104) <= '1';
    layer2_outputs(2105) <= not((layer1_outputs(7355)) or (layer1_outputs(6597)));
    layer2_outputs(2106) <= not(layer1_outputs(1578)) or (layer1_outputs(4121));
    layer2_outputs(2107) <= not(layer1_outputs(5892));
    layer2_outputs(2108) <= '0';
    layer2_outputs(2109) <= not(layer1_outputs(1247));
    layer2_outputs(2110) <= '1';
    layer2_outputs(2111) <= '1';
    layer2_outputs(2112) <= not(layer1_outputs(6851)) or (layer1_outputs(1748));
    layer2_outputs(2113) <= '1';
    layer2_outputs(2114) <= not(layer1_outputs(7513));
    layer2_outputs(2115) <= layer1_outputs(4703);
    layer2_outputs(2116) <= '1';
    layer2_outputs(2117) <= '0';
    layer2_outputs(2118) <= not((layer1_outputs(2585)) or (layer1_outputs(3476)));
    layer2_outputs(2119) <= '0';
    layer2_outputs(2120) <= (layer1_outputs(7344)) and (layer1_outputs(4701));
    layer2_outputs(2121) <= layer1_outputs(902);
    layer2_outputs(2122) <= '1';
    layer2_outputs(2123) <= not((layer1_outputs(5616)) and (layer1_outputs(2939)));
    layer2_outputs(2124) <= layer1_outputs(2926);
    layer2_outputs(2125) <= '0';
    layer2_outputs(2126) <= '0';
    layer2_outputs(2127) <= layer1_outputs(913);
    layer2_outputs(2128) <= not((layer1_outputs(2901)) and (layer1_outputs(2446)));
    layer2_outputs(2129) <= (layer1_outputs(3422)) and not (layer1_outputs(6226));
    layer2_outputs(2130) <= not(layer1_outputs(1747));
    layer2_outputs(2131) <= not(layer1_outputs(1082)) or (layer1_outputs(4148));
    layer2_outputs(2132) <= layer1_outputs(4964);
    layer2_outputs(2133) <= (layer1_outputs(6428)) or (layer1_outputs(1315));
    layer2_outputs(2134) <= not(layer1_outputs(3496));
    layer2_outputs(2135) <= not(layer1_outputs(4449));
    layer2_outputs(2136) <= not(layer1_outputs(5683));
    layer2_outputs(2137) <= (layer1_outputs(2395)) and not (layer1_outputs(25));
    layer2_outputs(2138) <= '0';
    layer2_outputs(2139) <= (layer1_outputs(5716)) or (layer1_outputs(5221));
    layer2_outputs(2140) <= (layer1_outputs(264)) or (layer1_outputs(540));
    layer2_outputs(2141) <= layer1_outputs(2303);
    layer2_outputs(2142) <= '1';
    layer2_outputs(2143) <= not(layer1_outputs(4297));
    layer2_outputs(2144) <= not(layer1_outputs(2114)) or (layer1_outputs(468));
    layer2_outputs(2145) <= not((layer1_outputs(5249)) or (layer1_outputs(5707)));
    layer2_outputs(2146) <= not(layer1_outputs(6719)) or (layer1_outputs(661));
    layer2_outputs(2147) <= not((layer1_outputs(474)) or (layer1_outputs(3307)));
    layer2_outputs(2148) <= not(layer1_outputs(6540)) or (layer1_outputs(307));
    layer2_outputs(2149) <= not(layer1_outputs(3439)) or (layer1_outputs(2358));
    layer2_outputs(2150) <= (layer1_outputs(6032)) and (layer1_outputs(3595));
    layer2_outputs(2151) <= (layer1_outputs(2547)) or (layer1_outputs(1235));
    layer2_outputs(2152) <= (layer1_outputs(6285)) and (layer1_outputs(664));
    layer2_outputs(2153) <= layer1_outputs(5929);
    layer2_outputs(2154) <= not(layer1_outputs(2103));
    layer2_outputs(2155) <= not(layer1_outputs(3124));
    layer2_outputs(2156) <= not((layer1_outputs(2663)) or (layer1_outputs(6309)));
    layer2_outputs(2157) <= layer1_outputs(7472);
    layer2_outputs(2158) <= not(layer1_outputs(5717));
    layer2_outputs(2159) <= not(layer1_outputs(1257)) or (layer1_outputs(116));
    layer2_outputs(2160) <= not(layer1_outputs(1502)) or (layer1_outputs(1296));
    layer2_outputs(2161) <= (layer1_outputs(480)) or (layer1_outputs(6027));
    layer2_outputs(2162) <= (layer1_outputs(4834)) and not (layer1_outputs(1949));
    layer2_outputs(2163) <= layer1_outputs(3106);
    layer2_outputs(2164) <= not((layer1_outputs(1674)) or (layer1_outputs(2324)));
    layer2_outputs(2165) <= layer1_outputs(761);
    layer2_outputs(2166) <= not(layer1_outputs(7471));
    layer2_outputs(2167) <= '0';
    layer2_outputs(2168) <= '1';
    layer2_outputs(2169) <= not(layer1_outputs(1768));
    layer2_outputs(2170) <= (layer1_outputs(2348)) and not (layer1_outputs(1731));
    layer2_outputs(2171) <= (layer1_outputs(7482)) or (layer1_outputs(6629));
    layer2_outputs(2172) <= layer1_outputs(2562);
    layer2_outputs(2173) <= '1';
    layer2_outputs(2174) <= layer1_outputs(8);
    layer2_outputs(2175) <= '1';
    layer2_outputs(2176) <= not(layer1_outputs(2293)) or (layer1_outputs(251));
    layer2_outputs(2177) <= layer1_outputs(2752);
    layer2_outputs(2178) <= (layer1_outputs(3200)) and not (layer1_outputs(5453));
    layer2_outputs(2179) <= not(layer1_outputs(5127));
    layer2_outputs(2180) <= not((layer1_outputs(1637)) and (layer1_outputs(3637)));
    layer2_outputs(2181) <= not(layer1_outputs(4177));
    layer2_outputs(2182) <= not(layer1_outputs(4347)) or (layer1_outputs(2821));
    layer2_outputs(2183) <= not((layer1_outputs(3616)) or (layer1_outputs(4026)));
    layer2_outputs(2184) <= not((layer1_outputs(6795)) or (layer1_outputs(5251)));
    layer2_outputs(2185) <= not(layer1_outputs(2709));
    layer2_outputs(2186) <= not(layer1_outputs(1656));
    layer2_outputs(2187) <= layer1_outputs(4367);
    layer2_outputs(2188) <= (layer1_outputs(864)) and not (layer1_outputs(5942));
    layer2_outputs(2189) <= not(layer1_outputs(5730));
    layer2_outputs(2190) <= (layer1_outputs(1006)) and (layer1_outputs(1286));
    layer2_outputs(2191) <= layer1_outputs(4235);
    layer2_outputs(2192) <= not((layer1_outputs(7400)) xor (layer1_outputs(3338)));
    layer2_outputs(2193) <= (layer1_outputs(2231)) and not (layer1_outputs(4193));
    layer2_outputs(2194) <= (layer1_outputs(3143)) and (layer1_outputs(2913));
    layer2_outputs(2195) <= layer1_outputs(118);
    layer2_outputs(2196) <= layer1_outputs(5496);
    layer2_outputs(2197) <= (layer1_outputs(2997)) or (layer1_outputs(1333));
    layer2_outputs(2198) <= layer1_outputs(1585);
    layer2_outputs(2199) <= layer1_outputs(5897);
    layer2_outputs(2200) <= '1';
    layer2_outputs(2201) <= not((layer1_outputs(6307)) and (layer1_outputs(5330)));
    layer2_outputs(2202) <= '1';
    layer2_outputs(2203) <= not(layer1_outputs(5869)) or (layer1_outputs(1888));
    layer2_outputs(2204) <= layer1_outputs(4584);
    layer2_outputs(2205) <= not(layer1_outputs(2852)) or (layer1_outputs(4448));
    layer2_outputs(2206) <= '0';
    layer2_outputs(2207) <= not((layer1_outputs(586)) or (layer1_outputs(7140)));
    layer2_outputs(2208) <= layer1_outputs(2988);
    layer2_outputs(2209) <= layer1_outputs(4163);
    layer2_outputs(2210) <= layer1_outputs(3250);
    layer2_outputs(2211) <= layer1_outputs(6015);
    layer2_outputs(2212) <= layer1_outputs(712);
    layer2_outputs(2213) <= not(layer1_outputs(880));
    layer2_outputs(2214) <= '0';
    layer2_outputs(2215) <= not(layer1_outputs(2161)) or (layer1_outputs(3771));
    layer2_outputs(2216) <= (layer1_outputs(2898)) or (layer1_outputs(1880));
    layer2_outputs(2217) <= not(layer1_outputs(6421));
    layer2_outputs(2218) <= not(layer1_outputs(244)) or (layer1_outputs(4238));
    layer2_outputs(2219) <= (layer1_outputs(1990)) or (layer1_outputs(1845));
    layer2_outputs(2220) <= '1';
    layer2_outputs(2221) <= not(layer1_outputs(2290));
    layer2_outputs(2222) <= (layer1_outputs(4351)) and not (layer1_outputs(1259));
    layer2_outputs(2223) <= (layer1_outputs(3018)) and not (layer1_outputs(2711));
    layer2_outputs(2224) <= '1';
    layer2_outputs(2225) <= not((layer1_outputs(3045)) and (layer1_outputs(7566)));
    layer2_outputs(2226) <= (layer1_outputs(757)) or (layer1_outputs(4896));
    layer2_outputs(2227) <= (layer1_outputs(2334)) and not (layer1_outputs(5662));
    layer2_outputs(2228) <= not(layer1_outputs(5937)) or (layer1_outputs(5206));
    layer2_outputs(2229) <= '0';
    layer2_outputs(2230) <= (layer1_outputs(2072)) and (layer1_outputs(2670));
    layer2_outputs(2231) <= layer1_outputs(7596);
    layer2_outputs(2232) <= not(layer1_outputs(6266));
    layer2_outputs(2233) <= (layer1_outputs(1393)) and not (layer1_outputs(5084));
    layer2_outputs(2234) <= (layer1_outputs(1043)) and not (layer1_outputs(2021));
    layer2_outputs(2235) <= not(layer1_outputs(7175)) or (layer1_outputs(4598));
    layer2_outputs(2236) <= layer1_outputs(4259);
    layer2_outputs(2237) <= not(layer1_outputs(2734));
    layer2_outputs(2238) <= not(layer1_outputs(3321));
    layer2_outputs(2239) <= not(layer1_outputs(3843));
    layer2_outputs(2240) <= layer1_outputs(2652);
    layer2_outputs(2241) <= not((layer1_outputs(5915)) or (layer1_outputs(812)));
    layer2_outputs(2242) <= (layer1_outputs(649)) and not (layer1_outputs(3470));
    layer2_outputs(2243) <= '0';
    layer2_outputs(2244) <= '1';
    layer2_outputs(2245) <= not(layer1_outputs(2349));
    layer2_outputs(2246) <= layer1_outputs(1441);
    layer2_outputs(2247) <= not((layer1_outputs(4218)) or (layer1_outputs(2137)));
    layer2_outputs(2248) <= (layer1_outputs(1409)) and not (layer1_outputs(4132));
    layer2_outputs(2249) <= layer1_outputs(786);
    layer2_outputs(2250) <= layer1_outputs(5047);
    layer2_outputs(2251) <= not(layer1_outputs(7375));
    layer2_outputs(2252) <= (layer1_outputs(541)) or (layer1_outputs(6708));
    layer2_outputs(2253) <= not((layer1_outputs(5059)) xor (layer1_outputs(6001)));
    layer2_outputs(2254) <= not(layer1_outputs(1424));
    layer2_outputs(2255) <= not(layer1_outputs(5831)) or (layer1_outputs(6886));
    layer2_outputs(2256) <= '1';
    layer2_outputs(2257) <= not((layer1_outputs(6079)) and (layer1_outputs(2785)));
    layer2_outputs(2258) <= '0';
    layer2_outputs(2259) <= '0';
    layer2_outputs(2260) <= (layer1_outputs(2788)) and (layer1_outputs(6018));
    layer2_outputs(2261) <= layer1_outputs(5059);
    layer2_outputs(2262) <= not(layer1_outputs(61));
    layer2_outputs(2263) <= layer1_outputs(4997);
    layer2_outputs(2264) <= (layer1_outputs(1096)) and not (layer1_outputs(1921));
    layer2_outputs(2265) <= '0';
    layer2_outputs(2266) <= '0';
    layer2_outputs(2267) <= layer1_outputs(7432);
    layer2_outputs(2268) <= not(layer1_outputs(6083));
    layer2_outputs(2269) <= not(layer1_outputs(5401));
    layer2_outputs(2270) <= not(layer1_outputs(2242)) or (layer1_outputs(4831));
    layer2_outputs(2271) <= not(layer1_outputs(4094));
    layer2_outputs(2272) <= layer1_outputs(2397);
    layer2_outputs(2273) <= layer1_outputs(5106);
    layer2_outputs(2274) <= '0';
    layer2_outputs(2275) <= (layer1_outputs(4803)) and not (layer1_outputs(580));
    layer2_outputs(2276) <= not(layer1_outputs(83));
    layer2_outputs(2277) <= layer1_outputs(4638);
    layer2_outputs(2278) <= (layer1_outputs(4033)) or (layer1_outputs(6625));
    layer2_outputs(2279) <= (layer1_outputs(7403)) or (layer1_outputs(1212));
    layer2_outputs(2280) <= not((layer1_outputs(7600)) or (layer1_outputs(7364)));
    layer2_outputs(2281) <= not(layer1_outputs(4305));
    layer2_outputs(2282) <= (layer1_outputs(6622)) and not (layer1_outputs(2177));
    layer2_outputs(2283) <= layer1_outputs(5906);
    layer2_outputs(2284) <= not((layer1_outputs(653)) or (layer1_outputs(7199)));
    layer2_outputs(2285) <= (layer1_outputs(7309)) and not (layer1_outputs(6796));
    layer2_outputs(2286) <= '1';
    layer2_outputs(2287) <= (layer1_outputs(1719)) and (layer1_outputs(4302));
    layer2_outputs(2288) <= layer1_outputs(7462);
    layer2_outputs(2289) <= (layer1_outputs(2280)) and (layer1_outputs(6410));
    layer2_outputs(2290) <= not(layer1_outputs(4036)) or (layer1_outputs(4200));
    layer2_outputs(2291) <= (layer1_outputs(859)) or (layer1_outputs(6857));
    layer2_outputs(2292) <= (layer1_outputs(3569)) or (layer1_outputs(5792));
    layer2_outputs(2293) <= not(layer1_outputs(7116)) or (layer1_outputs(2496));
    layer2_outputs(2294) <= not(layer1_outputs(6944)) or (layer1_outputs(199));
    layer2_outputs(2295) <= layer1_outputs(252);
    layer2_outputs(2296) <= not(layer1_outputs(1534)) or (layer1_outputs(5262));
    layer2_outputs(2297) <= layer1_outputs(6124);
    layer2_outputs(2298) <= not((layer1_outputs(2349)) and (layer1_outputs(5631)));
    layer2_outputs(2299) <= '0';
    layer2_outputs(2300) <= '1';
    layer2_outputs(2301) <= not((layer1_outputs(4615)) or (layer1_outputs(1385)));
    layer2_outputs(2302) <= (layer1_outputs(2492)) and (layer1_outputs(7676));
    layer2_outputs(2303) <= (layer1_outputs(1749)) or (layer1_outputs(1164));
    layer2_outputs(2304) <= not(layer1_outputs(3191)) or (layer1_outputs(3434));
    layer2_outputs(2305) <= layer1_outputs(7636);
    layer2_outputs(2306) <= not((layer1_outputs(6391)) or (layer1_outputs(7159)));
    layer2_outputs(2307) <= '0';
    layer2_outputs(2308) <= layer1_outputs(164);
    layer2_outputs(2309) <= not((layer1_outputs(2675)) xor (layer1_outputs(1918)));
    layer2_outputs(2310) <= layer1_outputs(2588);
    layer2_outputs(2311) <= not(layer1_outputs(1211));
    layer2_outputs(2312) <= not((layer1_outputs(3339)) and (layer1_outputs(917)));
    layer2_outputs(2313) <= not(layer1_outputs(3220)) or (layer1_outputs(6560));
    layer2_outputs(2314) <= (layer1_outputs(1376)) and not (layer1_outputs(612));
    layer2_outputs(2315) <= not(layer1_outputs(5156)) or (layer1_outputs(6279));
    layer2_outputs(2316) <= not(layer1_outputs(4483)) or (layer1_outputs(2891));
    layer2_outputs(2317) <= (layer1_outputs(702)) and (layer1_outputs(2183));
    layer2_outputs(2318) <= (layer1_outputs(5048)) and (layer1_outputs(4990));
    layer2_outputs(2319) <= not((layer1_outputs(538)) or (layer1_outputs(1217)));
    layer2_outputs(2320) <= not(layer1_outputs(5047));
    layer2_outputs(2321) <= not((layer1_outputs(936)) or (layer1_outputs(6504)));
    layer2_outputs(2322) <= not(layer1_outputs(4181));
    layer2_outputs(2323) <= layer1_outputs(7448);
    layer2_outputs(2324) <= layer1_outputs(4113);
    layer2_outputs(2325) <= not(layer1_outputs(3999));
    layer2_outputs(2326) <= '0';
    layer2_outputs(2327) <= layer1_outputs(4276);
    layer2_outputs(2328) <= layer1_outputs(693);
    layer2_outputs(2329) <= '0';
    layer2_outputs(2330) <= layer1_outputs(3745);
    layer2_outputs(2331) <= not(layer1_outputs(6757));
    layer2_outputs(2332) <= not(layer1_outputs(1637)) or (layer1_outputs(5011));
    layer2_outputs(2333) <= not((layer1_outputs(515)) and (layer1_outputs(4663)));
    layer2_outputs(2334) <= not(layer1_outputs(7301));
    layer2_outputs(2335) <= '0';
    layer2_outputs(2336) <= layer1_outputs(2308);
    layer2_outputs(2337) <= (layer1_outputs(4596)) and not (layer1_outputs(7535));
    layer2_outputs(2338) <= layer1_outputs(6020);
    layer2_outputs(2339) <= not(layer1_outputs(5629)) or (layer1_outputs(3715));
    layer2_outputs(2340) <= not(layer1_outputs(3521));
    layer2_outputs(2341) <= (layer1_outputs(1496)) and not (layer1_outputs(4146));
    layer2_outputs(2342) <= (layer1_outputs(3404)) or (layer1_outputs(5057));
    layer2_outputs(2343) <= (layer1_outputs(2559)) and (layer1_outputs(4730));
    layer2_outputs(2344) <= (layer1_outputs(4573)) and (layer1_outputs(7631));
    layer2_outputs(2345) <= layer1_outputs(311);
    layer2_outputs(2346) <= not(layer1_outputs(4891));
    layer2_outputs(2347) <= (layer1_outputs(2025)) and not (layer1_outputs(5387));
    layer2_outputs(2348) <= (layer1_outputs(5771)) xor (layer1_outputs(5203));
    layer2_outputs(2349) <= '1';
    layer2_outputs(2350) <= not(layer1_outputs(5004));
    layer2_outputs(2351) <= (layer1_outputs(3794)) or (layer1_outputs(7556));
    layer2_outputs(2352) <= not(layer1_outputs(3567)) or (layer1_outputs(3590));
    layer2_outputs(2353) <= not((layer1_outputs(6816)) or (layer1_outputs(6592)));
    layer2_outputs(2354) <= layer1_outputs(5804);
    layer2_outputs(2355) <= layer1_outputs(872);
    layer2_outputs(2356) <= '1';
    layer2_outputs(2357) <= not((layer1_outputs(7222)) xor (layer1_outputs(2281)));
    layer2_outputs(2358) <= not((layer1_outputs(4814)) xor (layer1_outputs(2228)));
    layer2_outputs(2359) <= (layer1_outputs(3802)) and not (layer1_outputs(3649));
    layer2_outputs(2360) <= '1';
    layer2_outputs(2361) <= not(layer1_outputs(6366)) or (layer1_outputs(4733));
    layer2_outputs(2362) <= (layer1_outputs(6422)) and not (layer1_outputs(6480));
    layer2_outputs(2363) <= not((layer1_outputs(973)) or (layer1_outputs(5128)));
    layer2_outputs(2364) <= layer1_outputs(7455);
    layer2_outputs(2365) <= layer1_outputs(1774);
    layer2_outputs(2366) <= (layer1_outputs(4224)) and not (layer1_outputs(2678));
    layer2_outputs(2367) <= (layer1_outputs(7563)) and (layer1_outputs(5093));
    layer2_outputs(2368) <= layer1_outputs(4099);
    layer2_outputs(2369) <= (layer1_outputs(708)) and not (layer1_outputs(1016));
    layer2_outputs(2370) <= (layer1_outputs(3400)) and not (layer1_outputs(7577));
    layer2_outputs(2371) <= layer1_outputs(1396);
    layer2_outputs(2372) <= '1';
    layer2_outputs(2373) <= not((layer1_outputs(4157)) or (layer1_outputs(547)));
    layer2_outputs(2374) <= (layer1_outputs(1459)) and not (layer1_outputs(1371));
    layer2_outputs(2375) <= (layer1_outputs(4023)) and not (layer1_outputs(2819));
    layer2_outputs(2376) <= (layer1_outputs(7256)) and not (layer1_outputs(5379));
    layer2_outputs(2377) <= not(layer1_outputs(3250));
    layer2_outputs(2378) <= layer1_outputs(3581);
    layer2_outputs(2379) <= layer1_outputs(4283);
    layer2_outputs(2380) <= not(layer1_outputs(2559));
    layer2_outputs(2381) <= layer1_outputs(7267);
    layer2_outputs(2382) <= not(layer1_outputs(4826));
    layer2_outputs(2383) <= not(layer1_outputs(6239));
    layer2_outputs(2384) <= (layer1_outputs(3414)) and (layer1_outputs(6378));
    layer2_outputs(2385) <= not(layer1_outputs(57));
    layer2_outputs(2386) <= layer1_outputs(2161);
    layer2_outputs(2387) <= not(layer1_outputs(4556));
    layer2_outputs(2388) <= layer1_outputs(4728);
    layer2_outputs(2389) <= (layer1_outputs(506)) or (layer1_outputs(2745));
    layer2_outputs(2390) <= '0';
    layer2_outputs(2391) <= '1';
    layer2_outputs(2392) <= '1';
    layer2_outputs(2393) <= layer1_outputs(500);
    layer2_outputs(2394) <= not((layer1_outputs(1861)) or (layer1_outputs(3665)));
    layer2_outputs(2395) <= not((layer1_outputs(2587)) and (layer1_outputs(1411)));
    layer2_outputs(2396) <= layer1_outputs(4631);
    layer2_outputs(2397) <= layer1_outputs(1029);
    layer2_outputs(2398) <= layer1_outputs(7604);
    layer2_outputs(2399) <= not(layer1_outputs(3886)) or (layer1_outputs(267));
    layer2_outputs(2400) <= not(layer1_outputs(3519));
    layer2_outputs(2401) <= not((layer1_outputs(6824)) or (layer1_outputs(2788)));
    layer2_outputs(2402) <= not((layer1_outputs(2171)) or (layer1_outputs(2049)));
    layer2_outputs(2403) <= not((layer1_outputs(883)) or (layer1_outputs(5148)));
    layer2_outputs(2404) <= '0';
    layer2_outputs(2405) <= '0';
    layer2_outputs(2406) <= '0';
    layer2_outputs(2407) <= (layer1_outputs(1814)) or (layer1_outputs(752));
    layer2_outputs(2408) <= '1';
    layer2_outputs(2409) <= layer1_outputs(7638);
    layer2_outputs(2410) <= not((layer1_outputs(5972)) or (layer1_outputs(6603)));
    layer2_outputs(2411) <= layer1_outputs(3459);
    layer2_outputs(2412) <= not((layer1_outputs(5689)) or (layer1_outputs(5544)));
    layer2_outputs(2413) <= not(layer1_outputs(6141));
    layer2_outputs(2414) <= not(layer1_outputs(1212));
    layer2_outputs(2415) <= '0';
    layer2_outputs(2416) <= (layer1_outputs(6295)) and not (layer1_outputs(1207));
    layer2_outputs(2417) <= (layer1_outputs(2514)) and (layer1_outputs(2294));
    layer2_outputs(2418) <= not((layer1_outputs(2733)) or (layer1_outputs(2859)));
    layer2_outputs(2419) <= not(layer1_outputs(498));
    layer2_outputs(2420) <= (layer1_outputs(1831)) or (layer1_outputs(3397));
    layer2_outputs(2421) <= layer1_outputs(1176);
    layer2_outputs(2422) <= '0';
    layer2_outputs(2423) <= '1';
    layer2_outputs(2424) <= layer1_outputs(5726);
    layer2_outputs(2425) <= not(layer1_outputs(3720)) or (layer1_outputs(6173));
    layer2_outputs(2426) <= not((layer1_outputs(3554)) or (layer1_outputs(1682)));
    layer2_outputs(2427) <= (layer1_outputs(4771)) and (layer1_outputs(6414));
    layer2_outputs(2428) <= '1';
    layer2_outputs(2429) <= (layer1_outputs(2944)) and not (layer1_outputs(448));
    layer2_outputs(2430) <= not(layer1_outputs(4078)) or (layer1_outputs(5759));
    layer2_outputs(2431) <= not((layer1_outputs(5628)) xor (layer1_outputs(3008)));
    layer2_outputs(2432) <= layer1_outputs(2317);
    layer2_outputs(2433) <= not(layer1_outputs(1670));
    layer2_outputs(2434) <= '1';
    layer2_outputs(2435) <= layer1_outputs(4925);
    layer2_outputs(2436) <= not(layer1_outputs(5327)) or (layer1_outputs(3732));
    layer2_outputs(2437) <= not(layer1_outputs(693)) or (layer1_outputs(1421));
    layer2_outputs(2438) <= '1';
    layer2_outputs(2439) <= layer1_outputs(1180);
    layer2_outputs(2440) <= not(layer1_outputs(811));
    layer2_outputs(2441) <= '0';
    layer2_outputs(2442) <= layer1_outputs(5162);
    layer2_outputs(2443) <= not((layer1_outputs(881)) and (layer1_outputs(3236)));
    layer2_outputs(2444) <= layer1_outputs(4074);
    layer2_outputs(2445) <= '1';
    layer2_outputs(2446) <= not((layer1_outputs(380)) and (layer1_outputs(2251)));
    layer2_outputs(2447) <= (layer1_outputs(3630)) and not (layer1_outputs(5616));
    layer2_outputs(2448) <= '1';
    layer2_outputs(2449) <= (layer1_outputs(3875)) and not (layer1_outputs(2776));
    layer2_outputs(2450) <= not(layer1_outputs(3123));
    layer2_outputs(2451) <= '0';
    layer2_outputs(2452) <= not((layer1_outputs(1131)) and (layer1_outputs(5636)));
    layer2_outputs(2453) <= (layer1_outputs(4480)) and not (layer1_outputs(4452));
    layer2_outputs(2454) <= layer1_outputs(1816);
    layer2_outputs(2455) <= layer1_outputs(6316);
    layer2_outputs(2456) <= not(layer1_outputs(2748));
    layer2_outputs(2457) <= not(layer1_outputs(6783));
    layer2_outputs(2458) <= layer1_outputs(840);
    layer2_outputs(2459) <= not(layer1_outputs(6782));
    layer2_outputs(2460) <= '0';
    layer2_outputs(2461) <= layer1_outputs(3251);
    layer2_outputs(2462) <= not(layer1_outputs(4475)) or (layer1_outputs(6290));
    layer2_outputs(2463) <= not(layer1_outputs(538));
    layer2_outputs(2464) <= not((layer1_outputs(5470)) and (layer1_outputs(2323)));
    layer2_outputs(2465) <= (layer1_outputs(6624)) xor (layer1_outputs(4593));
    layer2_outputs(2466) <= not(layer1_outputs(1622));
    layer2_outputs(2467) <= not(layer1_outputs(1028));
    layer2_outputs(2468) <= layer1_outputs(403);
    layer2_outputs(2469) <= layer1_outputs(4129);
    layer2_outputs(2470) <= not(layer1_outputs(2705)) or (layer1_outputs(1050));
    layer2_outputs(2471) <= layer1_outputs(1928);
    layer2_outputs(2472) <= not(layer1_outputs(2461));
    layer2_outputs(2473) <= not(layer1_outputs(6488));
    layer2_outputs(2474) <= not((layer1_outputs(5929)) or (layer1_outputs(4870)));
    layer2_outputs(2475) <= layer1_outputs(6391);
    layer2_outputs(2476) <= (layer1_outputs(3499)) xor (layer1_outputs(7453));
    layer2_outputs(2477) <= not(layer1_outputs(3094));
    layer2_outputs(2478) <= (layer1_outputs(829)) or (layer1_outputs(4588));
    layer2_outputs(2479) <= (layer1_outputs(5087)) and not (layer1_outputs(3986));
    layer2_outputs(2480) <= '0';
    layer2_outputs(2481) <= not(layer1_outputs(2875)) or (layer1_outputs(3136));
    layer2_outputs(2482) <= (layer1_outputs(4747)) and (layer1_outputs(5866));
    layer2_outputs(2483) <= not(layer1_outputs(7211)) or (layer1_outputs(1239));
    layer2_outputs(2484) <= layer1_outputs(5053);
    layer2_outputs(2485) <= not(layer1_outputs(6720));
    layer2_outputs(2486) <= not(layer1_outputs(2803));
    layer2_outputs(2487) <= not(layer1_outputs(2976)) or (layer1_outputs(1665));
    layer2_outputs(2488) <= '1';
    layer2_outputs(2489) <= not((layer1_outputs(510)) and (layer1_outputs(6778)));
    layer2_outputs(2490) <= not((layer1_outputs(5522)) and (layer1_outputs(1964)));
    layer2_outputs(2491) <= not((layer1_outputs(3820)) or (layer1_outputs(5941)));
    layer2_outputs(2492) <= '1';
    layer2_outputs(2493) <= (layer1_outputs(1559)) or (layer1_outputs(3440));
    layer2_outputs(2494) <= not(layer1_outputs(6651));
    layer2_outputs(2495) <= not(layer1_outputs(1969)) or (layer1_outputs(6291));
    layer2_outputs(2496) <= not((layer1_outputs(3531)) and (layer1_outputs(2194)));
    layer2_outputs(2497) <= not(layer1_outputs(4715)) or (layer1_outputs(6567));
    layer2_outputs(2498) <= (layer1_outputs(3777)) and (layer1_outputs(4126));
    layer2_outputs(2499) <= (layer1_outputs(6910)) and not (layer1_outputs(2116));
    layer2_outputs(2500) <= not(layer1_outputs(4023));
    layer2_outputs(2501) <= not(layer1_outputs(4411)) or (layer1_outputs(5239));
    layer2_outputs(2502) <= (layer1_outputs(7349)) and (layer1_outputs(195));
    layer2_outputs(2503) <= not((layer1_outputs(1566)) or (layer1_outputs(768)));
    layer2_outputs(2504) <= layer1_outputs(4012);
    layer2_outputs(2505) <= not((layer1_outputs(104)) or (layer1_outputs(7643)));
    layer2_outputs(2506) <= not(layer1_outputs(7305)) or (layer1_outputs(2186));
    layer2_outputs(2507) <= (layer1_outputs(4857)) and not (layer1_outputs(6939));
    layer2_outputs(2508) <= not(layer1_outputs(185));
    layer2_outputs(2509) <= (layer1_outputs(2119)) and not (layer1_outputs(1709));
    layer2_outputs(2510) <= not(layer1_outputs(7050)) or (layer1_outputs(5954));
    layer2_outputs(2511) <= (layer1_outputs(3829)) and (layer1_outputs(3933));
    layer2_outputs(2512) <= not(layer1_outputs(4928));
    layer2_outputs(2513) <= not((layer1_outputs(5076)) or (layer1_outputs(5070)));
    layer2_outputs(2514) <= (layer1_outputs(7639)) and not (layer1_outputs(6002));
    layer2_outputs(2515) <= layer1_outputs(4454);
    layer2_outputs(2516) <= (layer1_outputs(4575)) and (layer1_outputs(2602));
    layer2_outputs(2517) <= '0';
    layer2_outputs(2518) <= not(layer1_outputs(1370)) or (layer1_outputs(6190));
    layer2_outputs(2519) <= layer1_outputs(2222);
    layer2_outputs(2520) <= layer1_outputs(93);
    layer2_outputs(2521) <= layer1_outputs(4792);
    layer2_outputs(2522) <= layer1_outputs(3726);
    layer2_outputs(2523) <= (layer1_outputs(129)) and (layer1_outputs(5992));
    layer2_outputs(2524) <= not(layer1_outputs(2260));
    layer2_outputs(2525) <= not(layer1_outputs(2547)) or (layer1_outputs(4113));
    layer2_outputs(2526) <= '0';
    layer2_outputs(2527) <= not((layer1_outputs(3895)) or (layer1_outputs(6213)));
    layer2_outputs(2528) <= '0';
    layer2_outputs(2529) <= '0';
    layer2_outputs(2530) <= layer1_outputs(3813);
    layer2_outputs(2531) <= not((layer1_outputs(7624)) or (layer1_outputs(135)));
    layer2_outputs(2532) <= layer1_outputs(7432);
    layer2_outputs(2533) <= not(layer1_outputs(2241)) or (layer1_outputs(233));
    layer2_outputs(2534) <= not(layer1_outputs(7468));
    layer2_outputs(2535) <= not((layer1_outputs(6542)) and (layer1_outputs(3662)));
    layer2_outputs(2536) <= not((layer1_outputs(4840)) or (layer1_outputs(6739)));
    layer2_outputs(2537) <= not(layer1_outputs(7069));
    layer2_outputs(2538) <= not(layer1_outputs(5642));
    layer2_outputs(2539) <= not(layer1_outputs(230));
    layer2_outputs(2540) <= not(layer1_outputs(398));
    layer2_outputs(2541) <= (layer1_outputs(771)) and (layer1_outputs(2986));
    layer2_outputs(2542) <= (layer1_outputs(7135)) and (layer1_outputs(5019));
    layer2_outputs(2543) <= layer1_outputs(6418);
    layer2_outputs(2544) <= not(layer1_outputs(1807));
    layer2_outputs(2545) <= not((layer1_outputs(1085)) or (layer1_outputs(3503)));
    layer2_outputs(2546) <= layer1_outputs(4743);
    layer2_outputs(2547) <= not(layer1_outputs(1703)) or (layer1_outputs(3653));
    layer2_outputs(2548) <= (layer1_outputs(3089)) and not (layer1_outputs(1166));
    layer2_outputs(2549) <= not(layer1_outputs(7660)) or (layer1_outputs(5112));
    layer2_outputs(2550) <= '0';
    layer2_outputs(2551) <= not((layer1_outputs(7639)) and (layer1_outputs(2965)));
    layer2_outputs(2552) <= layer1_outputs(7425);
    layer2_outputs(2553) <= not(layer1_outputs(11));
    layer2_outputs(2554) <= not((layer1_outputs(2672)) or (layer1_outputs(5572)));
    layer2_outputs(2555) <= layer1_outputs(3856);
    layer2_outputs(2556) <= not(layer1_outputs(7241));
    layer2_outputs(2557) <= not(layer1_outputs(1380));
    layer2_outputs(2558) <= not(layer1_outputs(6675));
    layer2_outputs(2559) <= layer1_outputs(7537);
    layer2_outputs(2560) <= not(layer1_outputs(4115)) or (layer1_outputs(5352));
    layer2_outputs(2561) <= (layer1_outputs(5997)) and not (layer1_outputs(3313));
    layer2_outputs(2562) <= not(layer1_outputs(4597)) or (layer1_outputs(5267));
    layer2_outputs(2563) <= (layer1_outputs(2323)) and not (layer1_outputs(1796));
    layer2_outputs(2564) <= not((layer1_outputs(3610)) or (layer1_outputs(6430)));
    layer2_outputs(2565) <= not(layer1_outputs(4204)) or (layer1_outputs(5706));
    layer2_outputs(2566) <= (layer1_outputs(3554)) and not (layer1_outputs(1640));
    layer2_outputs(2567) <= '0';
    layer2_outputs(2568) <= not(layer1_outputs(5508));
    layer2_outputs(2569) <= not(layer1_outputs(3583));
    layer2_outputs(2570) <= '1';
    layer2_outputs(2571) <= '0';
    layer2_outputs(2572) <= (layer1_outputs(1832)) and not (layer1_outputs(4779));
    layer2_outputs(2573) <= not(layer1_outputs(3714));
    layer2_outputs(2574) <= '1';
    layer2_outputs(2575) <= (layer1_outputs(4707)) xor (layer1_outputs(2172));
    layer2_outputs(2576) <= '1';
    layer2_outputs(2577) <= (layer1_outputs(3342)) and not (layer1_outputs(6881));
    layer2_outputs(2578) <= not(layer1_outputs(5832)) or (layer1_outputs(5417));
    layer2_outputs(2579) <= layer1_outputs(4800);
    layer2_outputs(2580) <= layer1_outputs(1439);
    layer2_outputs(2581) <= (layer1_outputs(5894)) and (layer1_outputs(1812));
    layer2_outputs(2582) <= (layer1_outputs(320)) and (layer1_outputs(1042));
    layer2_outputs(2583) <= (layer1_outputs(3028)) and not (layer1_outputs(6170));
    layer2_outputs(2584) <= not(layer1_outputs(2915)) or (layer1_outputs(5042));
    layer2_outputs(2585) <= '1';
    layer2_outputs(2586) <= '0';
    layer2_outputs(2587) <= '0';
    layer2_outputs(2588) <= (layer1_outputs(3209)) and (layer1_outputs(4929));
    layer2_outputs(2589) <= not(layer1_outputs(5195)) or (layer1_outputs(457));
    layer2_outputs(2590) <= (layer1_outputs(7006)) or (layer1_outputs(7018));
    layer2_outputs(2591) <= (layer1_outputs(3786)) and not (layer1_outputs(2332));
    layer2_outputs(2592) <= not((layer1_outputs(7322)) or (layer1_outputs(560)));
    layer2_outputs(2593) <= layer1_outputs(3096);
    layer2_outputs(2594) <= layer1_outputs(3597);
    layer2_outputs(2595) <= not(layer1_outputs(7341));
    layer2_outputs(2596) <= layer1_outputs(4425);
    layer2_outputs(2597) <= (layer1_outputs(5153)) and not (layer1_outputs(2624));
    layer2_outputs(2598) <= not(layer1_outputs(5821));
    layer2_outputs(2599) <= layer1_outputs(5813);
    layer2_outputs(2600) <= not(layer1_outputs(2310)) or (layer1_outputs(1340));
    layer2_outputs(2601) <= not(layer1_outputs(1802));
    layer2_outputs(2602) <= not(layer1_outputs(4047)) or (layer1_outputs(2651));
    layer2_outputs(2603) <= '0';
    layer2_outputs(2604) <= not(layer1_outputs(2337)) or (layer1_outputs(4342));
    layer2_outputs(2605) <= layer1_outputs(3903);
    layer2_outputs(2606) <= (layer1_outputs(2181)) or (layer1_outputs(4609));
    layer2_outputs(2607) <= not((layer1_outputs(5357)) or (layer1_outputs(672)));
    layer2_outputs(2608) <= not(layer1_outputs(616)) or (layer1_outputs(559));
    layer2_outputs(2609) <= '0';
    layer2_outputs(2610) <= (layer1_outputs(5424)) and not (layer1_outputs(4993));
    layer2_outputs(2611) <= not(layer1_outputs(2973));
    layer2_outputs(2612) <= '1';
    layer2_outputs(2613) <= layer1_outputs(6232);
    layer2_outputs(2614) <= (layer1_outputs(7401)) and (layer1_outputs(6677));
    layer2_outputs(2615) <= layer1_outputs(2387);
    layer2_outputs(2616) <= '0';
    layer2_outputs(2617) <= (layer1_outputs(446)) and (layer1_outputs(4689));
    layer2_outputs(2618) <= '0';
    layer2_outputs(2619) <= (layer1_outputs(1111)) and not (layer1_outputs(4191));
    layer2_outputs(2620) <= '1';
    layer2_outputs(2621) <= layer1_outputs(5867);
    layer2_outputs(2622) <= not(layer1_outputs(4538));
    layer2_outputs(2623) <= (layer1_outputs(4581)) and not (layer1_outputs(4401));
    layer2_outputs(2624) <= (layer1_outputs(7098)) and not (layer1_outputs(5516));
    layer2_outputs(2625) <= not(layer1_outputs(6532)) or (layer1_outputs(7627));
    layer2_outputs(2626) <= not(layer1_outputs(6562));
    layer2_outputs(2627) <= (layer1_outputs(4846)) or (layer1_outputs(3891));
    layer2_outputs(2628) <= not(layer1_outputs(1523));
    layer2_outputs(2629) <= not(layer1_outputs(1715)) or (layer1_outputs(526));
    layer2_outputs(2630) <= (layer1_outputs(2654)) and not (layer1_outputs(6505));
    layer2_outputs(2631) <= not((layer1_outputs(6249)) and (layer1_outputs(4409)));
    layer2_outputs(2632) <= not(layer1_outputs(3026)) or (layer1_outputs(3215));
    layer2_outputs(2633) <= not(layer1_outputs(468)) or (layer1_outputs(297));
    layer2_outputs(2634) <= (layer1_outputs(1771)) xor (layer1_outputs(3805));
    layer2_outputs(2635) <= '1';
    layer2_outputs(2636) <= not(layer1_outputs(4964)) or (layer1_outputs(2468));
    layer2_outputs(2637) <= not(layer1_outputs(6528)) or (layer1_outputs(5414));
    layer2_outputs(2638) <= '0';
    layer2_outputs(2639) <= '1';
    layer2_outputs(2640) <= (layer1_outputs(2613)) and not (layer1_outputs(2370));
    layer2_outputs(2641) <= not(layer1_outputs(5611)) or (layer1_outputs(168));
    layer2_outputs(2642) <= not(layer1_outputs(4957)) or (layer1_outputs(2242));
    layer2_outputs(2643) <= '1';
    layer2_outputs(2644) <= layer1_outputs(4628);
    layer2_outputs(2645) <= not(layer1_outputs(5575)) or (layer1_outputs(684));
    layer2_outputs(2646) <= not(layer1_outputs(2566));
    layer2_outputs(2647) <= '1';
    layer2_outputs(2648) <= (layer1_outputs(1085)) and not (layer1_outputs(4219));
    layer2_outputs(2649) <= (layer1_outputs(488)) and (layer1_outputs(2168));
    layer2_outputs(2650) <= layer1_outputs(4901);
    layer2_outputs(2651) <= not(layer1_outputs(6986)) or (layer1_outputs(1195));
    layer2_outputs(2652) <= not(layer1_outputs(2570)) or (layer1_outputs(6564));
    layer2_outputs(2653) <= '1';
    layer2_outputs(2654) <= layer1_outputs(5560);
    layer2_outputs(2655) <= (layer1_outputs(1088)) xor (layer1_outputs(6851));
    layer2_outputs(2656) <= layer1_outputs(5754);
    layer2_outputs(2657) <= (layer1_outputs(5841)) and not (layer1_outputs(5181));
    layer2_outputs(2658) <= layer1_outputs(7504);
    layer2_outputs(2659) <= (layer1_outputs(4358)) or (layer1_outputs(961));
    layer2_outputs(2660) <= (layer1_outputs(5943)) and not (layer1_outputs(272));
    layer2_outputs(2661) <= not((layer1_outputs(2212)) or (layer1_outputs(7390)));
    layer2_outputs(2662) <= not(layer1_outputs(1767));
    layer2_outputs(2663) <= (layer1_outputs(5124)) and not (layer1_outputs(3071));
    layer2_outputs(2664) <= not(layer1_outputs(749)) or (layer1_outputs(6645));
    layer2_outputs(2665) <= (layer1_outputs(4119)) and (layer1_outputs(6824));
    layer2_outputs(2666) <= (layer1_outputs(6320)) and not (layer1_outputs(7284));
    layer2_outputs(2667) <= (layer1_outputs(2476)) and not (layer1_outputs(5922));
    layer2_outputs(2668) <= not(layer1_outputs(3498));
    layer2_outputs(2669) <= layer1_outputs(5776);
    layer2_outputs(2670) <= not(layer1_outputs(5636)) or (layer1_outputs(7020));
    layer2_outputs(2671) <= not((layer1_outputs(7473)) or (layer1_outputs(6346)));
    layer2_outputs(2672) <= not((layer1_outputs(7314)) or (layer1_outputs(822)));
    layer2_outputs(2673) <= not((layer1_outputs(7477)) or (layer1_outputs(895)));
    layer2_outputs(2674) <= layer1_outputs(173);
    layer2_outputs(2675) <= layer1_outputs(3217);
    layer2_outputs(2676) <= layer1_outputs(2399);
    layer2_outputs(2677) <= (layer1_outputs(62)) and not (layer1_outputs(6813));
    layer2_outputs(2678) <= (layer1_outputs(5193)) and not (layer1_outputs(360));
    layer2_outputs(2679) <= (layer1_outputs(948)) and not (layer1_outputs(6922));
    layer2_outputs(2680) <= not(layer1_outputs(704));
    layer2_outputs(2681) <= not((layer1_outputs(4274)) or (layer1_outputs(6498)));
    layer2_outputs(2682) <= not(layer1_outputs(7538)) or (layer1_outputs(1392));
    layer2_outputs(2683) <= not(layer1_outputs(3100));
    layer2_outputs(2684) <= not(layer1_outputs(3092)) or (layer1_outputs(4984));
    layer2_outputs(2685) <= not(layer1_outputs(7030));
    layer2_outputs(2686) <= '0';
    layer2_outputs(2687) <= (layer1_outputs(3173)) and not (layer1_outputs(7086));
    layer2_outputs(2688) <= not(layer1_outputs(234));
    layer2_outputs(2689) <= (layer1_outputs(4117)) and not (layer1_outputs(3635));
    layer2_outputs(2690) <= '0';
    layer2_outputs(2691) <= layer1_outputs(409);
    layer2_outputs(2692) <= layer1_outputs(117);
    layer2_outputs(2693) <= not(layer1_outputs(743)) or (layer1_outputs(6977));
    layer2_outputs(2694) <= not((layer1_outputs(3831)) and (layer1_outputs(656)));
    layer2_outputs(2695) <= (layer1_outputs(6172)) and (layer1_outputs(4523));
    layer2_outputs(2696) <= not(layer1_outputs(7122));
    layer2_outputs(2697) <= (layer1_outputs(4633)) and not (layer1_outputs(7638));
    layer2_outputs(2698) <= '1';
    layer2_outputs(2699) <= not((layer1_outputs(1274)) and (layer1_outputs(2581)));
    layer2_outputs(2700) <= layer1_outputs(4119);
    layer2_outputs(2701) <= (layer1_outputs(1245)) and not (layer1_outputs(6865));
    layer2_outputs(2702) <= not(layer1_outputs(1813));
    layer2_outputs(2703) <= '0';
    layer2_outputs(2704) <= (layer1_outputs(1671)) and (layer1_outputs(2875));
    layer2_outputs(2705) <= (layer1_outputs(6476)) or (layer1_outputs(4725));
    layer2_outputs(2706) <= not((layer1_outputs(6024)) or (layer1_outputs(1012)));
    layer2_outputs(2707) <= not(layer1_outputs(5368));
    layer2_outputs(2708) <= '1';
    layer2_outputs(2709) <= '1';
    layer2_outputs(2710) <= (layer1_outputs(6525)) and not (layer1_outputs(3731));
    layer2_outputs(2711) <= (layer1_outputs(755)) and not (layer1_outputs(2468));
    layer2_outputs(2712) <= not(layer1_outputs(3388)) or (layer1_outputs(1108));
    layer2_outputs(2713) <= not((layer1_outputs(1626)) and (layer1_outputs(1530)));
    layer2_outputs(2714) <= not(layer1_outputs(6131));
    layer2_outputs(2715) <= layer1_outputs(39);
    layer2_outputs(2716) <= '0';
    layer2_outputs(2717) <= not(layer1_outputs(7271));
    layer2_outputs(2718) <= not(layer1_outputs(3238));
    layer2_outputs(2719) <= '1';
    layer2_outputs(2720) <= '0';
    layer2_outputs(2721) <= not(layer1_outputs(3044)) or (layer1_outputs(7407));
    layer2_outputs(2722) <= (layer1_outputs(833)) and (layer1_outputs(4337));
    layer2_outputs(2723) <= (layer1_outputs(7580)) or (layer1_outputs(1916));
    layer2_outputs(2724) <= not(layer1_outputs(2638));
    layer2_outputs(2725) <= (layer1_outputs(5591)) and (layer1_outputs(7417));
    layer2_outputs(2726) <= not(layer1_outputs(2542));
    layer2_outputs(2727) <= (layer1_outputs(3866)) and (layer1_outputs(125));
    layer2_outputs(2728) <= not(layer1_outputs(5742)) or (layer1_outputs(4182));
    layer2_outputs(2729) <= not(layer1_outputs(6838));
    layer2_outputs(2730) <= (layer1_outputs(4795)) or (layer1_outputs(1358));
    layer2_outputs(2731) <= not(layer1_outputs(978)) or (layer1_outputs(7054));
    layer2_outputs(2732) <= not((layer1_outputs(2230)) and (layer1_outputs(1225)));
    layer2_outputs(2733) <= not((layer1_outputs(4974)) and (layer1_outputs(5436)));
    layer2_outputs(2734) <= (layer1_outputs(4141)) and (layer1_outputs(6655));
    layer2_outputs(2735) <= not(layer1_outputs(1284)) or (layer1_outputs(2038));
    layer2_outputs(2736) <= (layer1_outputs(4795)) and not (layer1_outputs(7306));
    layer2_outputs(2737) <= (layer1_outputs(6254)) and (layer1_outputs(6769));
    layer2_outputs(2738) <= (layer1_outputs(4536)) and not (layer1_outputs(270));
    layer2_outputs(2739) <= not(layer1_outputs(5954));
    layer2_outputs(2740) <= (layer1_outputs(4214)) and not (layer1_outputs(3792));
    layer2_outputs(2741) <= (layer1_outputs(7540)) or (layer1_outputs(343));
    layer2_outputs(2742) <= layer1_outputs(6595);
    layer2_outputs(2743) <= not(layer1_outputs(3147)) or (layer1_outputs(1536));
    layer2_outputs(2744) <= not((layer1_outputs(7)) and (layer1_outputs(2679)));
    layer2_outputs(2745) <= not(layer1_outputs(2464)) or (layer1_outputs(3145));
    layer2_outputs(2746) <= '1';
    layer2_outputs(2747) <= (layer1_outputs(1023)) and not (layer1_outputs(1242));
    layer2_outputs(2748) <= not(layer1_outputs(3824));
    layer2_outputs(2749) <= not((layer1_outputs(1600)) and (layer1_outputs(1886)));
    layer2_outputs(2750) <= not(layer1_outputs(7606));
    layer2_outputs(2751) <= '1';
    layer2_outputs(2752) <= '0';
    layer2_outputs(2753) <= (layer1_outputs(1005)) and (layer1_outputs(414));
    layer2_outputs(2754) <= '0';
    layer2_outputs(2755) <= layer1_outputs(6765);
    layer2_outputs(2756) <= not(layer1_outputs(6465));
    layer2_outputs(2757) <= layer1_outputs(3915);
    layer2_outputs(2758) <= layer1_outputs(3604);
    layer2_outputs(2759) <= not(layer1_outputs(504)) or (layer1_outputs(4923));
    layer2_outputs(2760) <= not(layer1_outputs(5192));
    layer2_outputs(2761) <= not(layer1_outputs(2644));
    layer2_outputs(2762) <= layer1_outputs(4545);
    layer2_outputs(2763) <= not(layer1_outputs(2180)) or (layer1_outputs(455));
    layer2_outputs(2764) <= '1';
    layer2_outputs(2765) <= (layer1_outputs(4764)) and not (layer1_outputs(7093));
    layer2_outputs(2766) <= '0';
    layer2_outputs(2767) <= layer1_outputs(477);
    layer2_outputs(2768) <= (layer1_outputs(6404)) and not (layer1_outputs(6770));
    layer2_outputs(2769) <= layer1_outputs(1010);
    layer2_outputs(2770) <= (layer1_outputs(6398)) and not (layer1_outputs(1508));
    layer2_outputs(2771) <= not(layer1_outputs(1780));
    layer2_outputs(2772) <= not((layer1_outputs(3573)) or (layer1_outputs(2847)));
    layer2_outputs(2773) <= layer1_outputs(534);
    layer2_outputs(2774) <= (layer1_outputs(3869)) or (layer1_outputs(3546));
    layer2_outputs(2775) <= layer1_outputs(6240);
    layer2_outputs(2776) <= not(layer1_outputs(7521)) or (layer1_outputs(7465));
    layer2_outputs(2777) <= not(layer1_outputs(7118));
    layer2_outputs(2778) <= (layer1_outputs(6906)) and (layer1_outputs(7237));
    layer2_outputs(2779) <= '1';
    layer2_outputs(2780) <= (layer1_outputs(4095)) and not (layer1_outputs(6898));
    layer2_outputs(2781) <= (layer1_outputs(6282)) and (layer1_outputs(2164));
    layer2_outputs(2782) <= '0';
    layer2_outputs(2783) <= not(layer1_outputs(2001));
    layer2_outputs(2784) <= '1';
    layer2_outputs(2785) <= (layer1_outputs(3914)) or (layer1_outputs(271));
    layer2_outputs(2786) <= (layer1_outputs(4767)) or (layer1_outputs(6855));
    layer2_outputs(2787) <= '0';
    layer2_outputs(2788) <= not((layer1_outputs(2449)) or (layer1_outputs(2838)));
    layer2_outputs(2789) <= not(layer1_outputs(6946));
    layer2_outputs(2790) <= not(layer1_outputs(3399)) or (layer1_outputs(216));
    layer2_outputs(2791) <= '1';
    layer2_outputs(2792) <= layer1_outputs(2494);
    layer2_outputs(2793) <= not(layer1_outputs(2680)) or (layer1_outputs(4608));
    layer2_outputs(2794) <= not(layer1_outputs(1457)) or (layer1_outputs(4578));
    layer2_outputs(2795) <= not((layer1_outputs(6114)) and (layer1_outputs(1707)));
    layer2_outputs(2796) <= (layer1_outputs(4355)) and (layer1_outputs(7365));
    layer2_outputs(2797) <= layer1_outputs(2627);
    layer2_outputs(2798) <= (layer1_outputs(2516)) and not (layer1_outputs(2373));
    layer2_outputs(2799) <= (layer1_outputs(4665)) and not (layer1_outputs(128));
    layer2_outputs(2800) <= not(layer1_outputs(4948));
    layer2_outputs(2801) <= layer1_outputs(6624);
    layer2_outputs(2802) <= '0';
    layer2_outputs(2803) <= not(layer1_outputs(6699));
    layer2_outputs(2804) <= layer1_outputs(3162);
    layer2_outputs(2805) <= '1';
    layer2_outputs(2806) <= not(layer1_outputs(2502));
    layer2_outputs(2807) <= (layer1_outputs(1116)) and (layer1_outputs(2512));
    layer2_outputs(2808) <= (layer1_outputs(364)) and (layer1_outputs(6110));
    layer2_outputs(2809) <= (layer1_outputs(6506)) and (layer1_outputs(1352));
    layer2_outputs(2810) <= not(layer1_outputs(6579));
    layer2_outputs(2811) <= layer1_outputs(5185);
    layer2_outputs(2812) <= '0';
    layer2_outputs(2813) <= layer1_outputs(6169);
    layer2_outputs(2814) <= (layer1_outputs(6846)) and not (layer1_outputs(5142));
    layer2_outputs(2815) <= not(layer1_outputs(3613)) or (layer1_outputs(1222));
    layer2_outputs(2816) <= not(layer1_outputs(7356)) or (layer1_outputs(6600));
    layer2_outputs(2817) <= '1';
    layer2_outputs(2818) <= '1';
    layer2_outputs(2819) <= layer1_outputs(5664);
    layer2_outputs(2820) <= (layer1_outputs(7676)) and not (layer1_outputs(1003));
    layer2_outputs(2821) <= not(layer1_outputs(484)) or (layer1_outputs(2208));
    layer2_outputs(2822) <= not(layer1_outputs(1046));
    layer2_outputs(2823) <= layer1_outputs(3024);
    layer2_outputs(2824) <= (layer1_outputs(7520)) or (layer1_outputs(3848));
    layer2_outputs(2825) <= '0';
    layer2_outputs(2826) <= (layer1_outputs(4931)) and not (layer1_outputs(98));
    layer2_outputs(2827) <= (layer1_outputs(6244)) and not (layer1_outputs(3431));
    layer2_outputs(2828) <= (layer1_outputs(1359)) and not (layer1_outputs(6183));
    layer2_outputs(2829) <= layer1_outputs(4230);
    layer2_outputs(2830) <= not(layer1_outputs(716));
    layer2_outputs(2831) <= '1';
    layer2_outputs(2832) <= not((layer1_outputs(3908)) and (layer1_outputs(1482)));
    layer2_outputs(2833) <= (layer1_outputs(5951)) and (layer1_outputs(5116));
    layer2_outputs(2834) <= layer1_outputs(7173);
    layer2_outputs(2835) <= not(layer1_outputs(5421)) or (layer1_outputs(1265));
    layer2_outputs(2836) <= (layer1_outputs(6898)) and not (layer1_outputs(3536));
    layer2_outputs(2837) <= (layer1_outputs(5585)) or (layer1_outputs(4180));
    layer2_outputs(2838) <= not(layer1_outputs(3276));
    layer2_outputs(2839) <= not(layer1_outputs(6490)) or (layer1_outputs(2012));
    layer2_outputs(2840) <= not(layer1_outputs(4330));
    layer2_outputs(2841) <= not(layer1_outputs(6270));
    layer2_outputs(2842) <= not((layer1_outputs(7119)) xor (layer1_outputs(1999)));
    layer2_outputs(2843) <= not(layer1_outputs(3714)) or (layer1_outputs(1185));
    layer2_outputs(2844) <= not(layer1_outputs(695));
    layer2_outputs(2845) <= (layer1_outputs(7256)) and not (layer1_outputs(1071));
    layer2_outputs(2846) <= layer1_outputs(7277);
    layer2_outputs(2847) <= (layer1_outputs(241)) and not (layer1_outputs(5454));
    layer2_outputs(2848) <= layer1_outputs(7532);
    layer2_outputs(2849) <= (layer1_outputs(5176)) or (layer1_outputs(1657));
    layer2_outputs(2850) <= not(layer1_outputs(6389)) or (layer1_outputs(3569));
    layer2_outputs(2851) <= not(layer1_outputs(6122)) or (layer1_outputs(1459));
    layer2_outputs(2852) <= not((layer1_outputs(7371)) or (layer1_outputs(5541)));
    layer2_outputs(2853) <= not(layer1_outputs(6333)) or (layer1_outputs(7663));
    layer2_outputs(2854) <= '0';
    layer2_outputs(2855) <= (layer1_outputs(3828)) and (layer1_outputs(7158));
    layer2_outputs(2856) <= layer1_outputs(6133);
    layer2_outputs(2857) <= '0';
    layer2_outputs(2858) <= not((layer1_outputs(7515)) and (layer1_outputs(6023)));
    layer2_outputs(2859) <= (layer1_outputs(3149)) and not (layer1_outputs(3754));
    layer2_outputs(2860) <= not(layer1_outputs(4161)) or (layer1_outputs(7623));
    layer2_outputs(2861) <= not((layer1_outputs(6908)) and (layer1_outputs(6752)));
    layer2_outputs(2862) <= (layer1_outputs(1926)) and not (layer1_outputs(2703));
    layer2_outputs(2863) <= '0';
    layer2_outputs(2864) <= (layer1_outputs(5284)) or (layer1_outputs(4898));
    layer2_outputs(2865) <= not((layer1_outputs(1022)) or (layer1_outputs(4558)));
    layer2_outputs(2866) <= '0';
    layer2_outputs(2867) <= not(layer1_outputs(385));
    layer2_outputs(2868) <= not(layer1_outputs(1448)) or (layer1_outputs(2118));
    layer2_outputs(2869) <= not(layer1_outputs(711));
    layer2_outputs(2870) <= not(layer1_outputs(5552)) or (layer1_outputs(4655));
    layer2_outputs(2871) <= (layer1_outputs(1625)) and not (layer1_outputs(3487));
    layer2_outputs(2872) <= '1';
    layer2_outputs(2873) <= '0';
    layer2_outputs(2874) <= not(layer1_outputs(2339)) or (layer1_outputs(7629));
    layer2_outputs(2875) <= not(layer1_outputs(1084));
    layer2_outputs(2876) <= not(layer1_outputs(3094)) or (layer1_outputs(5489));
    layer2_outputs(2877) <= (layer1_outputs(6387)) and not (layer1_outputs(6350));
    layer2_outputs(2878) <= (layer1_outputs(5539)) and not (layer1_outputs(3211));
    layer2_outputs(2879) <= '1';
    layer2_outputs(2880) <= layer1_outputs(3233);
    layer2_outputs(2881) <= (layer1_outputs(660)) and not (layer1_outputs(2449));
    layer2_outputs(2882) <= '1';
    layer2_outputs(2883) <= layer1_outputs(6814);
    layer2_outputs(2884) <= not(layer1_outputs(5879));
    layer2_outputs(2885) <= layer1_outputs(1503);
    layer2_outputs(2886) <= not((layer1_outputs(115)) xor (layer1_outputs(597)));
    layer2_outputs(2887) <= not((layer1_outputs(3989)) or (layer1_outputs(3154)));
    layer2_outputs(2888) <= not((layer1_outputs(6971)) and (layer1_outputs(5637)));
    layer2_outputs(2889) <= not((layer1_outputs(7589)) or (layer1_outputs(3660)));
    layer2_outputs(2890) <= not(layer1_outputs(3331));
    layer2_outputs(2891) <= layer1_outputs(6595);
    layer2_outputs(2892) <= (layer1_outputs(3754)) and (layer1_outputs(2846));
    layer2_outputs(2893) <= not((layer1_outputs(3736)) or (layer1_outputs(322)));
    layer2_outputs(2894) <= (layer1_outputs(4236)) and (layer1_outputs(1090));
    layer2_outputs(2895) <= not(layer1_outputs(1366));
    layer2_outputs(2896) <= layer1_outputs(5094);
    layer2_outputs(2897) <= (layer1_outputs(2838)) and (layer1_outputs(2995));
    layer2_outputs(2898) <= (layer1_outputs(7627)) and not (layer1_outputs(6111));
    layer2_outputs(2899) <= '0';
    layer2_outputs(2900) <= not(layer1_outputs(4201));
    layer2_outputs(2901) <= (layer1_outputs(1273)) or (layer1_outputs(2015));
    layer2_outputs(2902) <= (layer1_outputs(4235)) and not (layer1_outputs(649));
    layer2_outputs(2903) <= not(layer1_outputs(2270)) or (layer1_outputs(2104));
    layer2_outputs(2904) <= not((layer1_outputs(4121)) or (layer1_outputs(5702)));
    layer2_outputs(2905) <= not(layer1_outputs(7620)) or (layer1_outputs(1383));
    layer2_outputs(2906) <= not(layer1_outputs(5117));
    layer2_outputs(2907) <= not(layer1_outputs(7661));
    layer2_outputs(2908) <= (layer1_outputs(1949)) and not (layer1_outputs(6129));
    layer2_outputs(2909) <= not(layer1_outputs(1154));
    layer2_outputs(2910) <= not(layer1_outputs(1325));
    layer2_outputs(2911) <= '0';
    layer2_outputs(2912) <= not(layer1_outputs(7431));
    layer2_outputs(2913) <= layer1_outputs(2496);
    layer2_outputs(2914) <= '1';
    layer2_outputs(2915) <= not((layer1_outputs(5243)) or (layer1_outputs(7612)));
    layer2_outputs(2916) <= layer1_outputs(1407);
    layer2_outputs(2917) <= not((layer1_outputs(7125)) and (layer1_outputs(2120)));
    layer2_outputs(2918) <= not((layer1_outputs(1287)) or (layer1_outputs(1633)));
    layer2_outputs(2919) <= not(layer1_outputs(3604)) or (layer1_outputs(3181));
    layer2_outputs(2920) <= '0';
    layer2_outputs(2921) <= layer1_outputs(2710);
    layer2_outputs(2922) <= not(layer1_outputs(1130));
    layer2_outputs(2923) <= (layer1_outputs(2193)) or (layer1_outputs(4845));
    layer2_outputs(2924) <= layer1_outputs(1363);
    layer2_outputs(2925) <= (layer1_outputs(6135)) and (layer1_outputs(7567));
    layer2_outputs(2926) <= '1';
    layer2_outputs(2927) <= layer1_outputs(3022);
    layer2_outputs(2928) <= not(layer1_outputs(5240));
    layer2_outputs(2929) <= not(layer1_outputs(6901));
    layer2_outputs(2930) <= (layer1_outputs(5033)) and not (layer1_outputs(3855));
    layer2_outputs(2931) <= not(layer1_outputs(1318));
    layer2_outputs(2932) <= '1';
    layer2_outputs(2933) <= not(layer1_outputs(2934));
    layer2_outputs(2934) <= not((layer1_outputs(5633)) xor (layer1_outputs(5791)));
    layer2_outputs(2935) <= not(layer1_outputs(1133)) or (layer1_outputs(1618));
    layer2_outputs(2936) <= layer1_outputs(1153);
    layer2_outputs(2937) <= not((layer1_outputs(6362)) and (layer1_outputs(5589)));
    layer2_outputs(2938) <= '1';
    layer2_outputs(2939) <= layer1_outputs(819);
    layer2_outputs(2940) <= not(layer1_outputs(6353));
    layer2_outputs(2941) <= layer1_outputs(265);
    layer2_outputs(2942) <= not(layer1_outputs(1426));
    layer2_outputs(2943) <= not(layer1_outputs(5900));
    layer2_outputs(2944) <= '0';
    layer2_outputs(2945) <= not(layer1_outputs(2841));
    layer2_outputs(2946) <= (layer1_outputs(3812)) or (layer1_outputs(5069));
    layer2_outputs(2947) <= layer1_outputs(6147);
    layer2_outputs(2948) <= '0';
    layer2_outputs(2949) <= not((layer1_outputs(1511)) or (layer1_outputs(20)));
    layer2_outputs(2950) <= not(layer1_outputs(690));
    layer2_outputs(2951) <= not(layer1_outputs(4459)) or (layer1_outputs(5445));
    layer2_outputs(2952) <= layer1_outputs(2626);
    layer2_outputs(2953) <= layer1_outputs(6552);
    layer2_outputs(2954) <= layer1_outputs(528);
    layer2_outputs(2955) <= '0';
    layer2_outputs(2956) <= '0';
    layer2_outputs(2957) <= not((layer1_outputs(5590)) or (layer1_outputs(7072)));
    layer2_outputs(2958) <= not(layer1_outputs(3423)) or (layer1_outputs(2122));
    layer2_outputs(2959) <= '1';
    layer2_outputs(2960) <= '1';
    layer2_outputs(2961) <= (layer1_outputs(4762)) and not (layer1_outputs(494));
    layer2_outputs(2962) <= not((layer1_outputs(2828)) xor (layer1_outputs(6646)));
    layer2_outputs(2963) <= layer1_outputs(2406);
    layer2_outputs(2964) <= not((layer1_outputs(7427)) or (layer1_outputs(7209)));
    layer2_outputs(2965) <= '1';
    layer2_outputs(2966) <= (layer1_outputs(2668)) and not (layer1_outputs(3127));
    layer2_outputs(2967) <= layer1_outputs(3082);
    layer2_outputs(2968) <= (layer1_outputs(6223)) and not (layer1_outputs(6663));
    layer2_outputs(2969) <= (layer1_outputs(4480)) or (layer1_outputs(865));
    layer2_outputs(2970) <= '0';
    layer2_outputs(2971) <= (layer1_outputs(4294)) and not (layer1_outputs(2584));
    layer2_outputs(2972) <= layer1_outputs(3777);
    layer2_outputs(2973) <= layer1_outputs(5652);
    layer2_outputs(2974) <= (layer1_outputs(5734)) and (layer1_outputs(1186));
    layer2_outputs(2975) <= '1';
    layer2_outputs(2976) <= '0';
    layer2_outputs(2977) <= (layer1_outputs(5703)) xor (layer1_outputs(6417));
    layer2_outputs(2978) <= layer1_outputs(1228);
    layer2_outputs(2979) <= (layer1_outputs(6934)) or (layer1_outputs(3563));
    layer2_outputs(2980) <= (layer1_outputs(1072)) and not (layer1_outputs(4234));
    layer2_outputs(2981) <= not((layer1_outputs(938)) xor (layer1_outputs(6601)));
    layer2_outputs(2982) <= (layer1_outputs(6714)) and (layer1_outputs(3584));
    layer2_outputs(2983) <= '1';
    layer2_outputs(2984) <= not(layer1_outputs(3450)) or (layer1_outputs(1997));
    layer2_outputs(2985) <= not((layer1_outputs(5133)) and (layer1_outputs(3028)));
    layer2_outputs(2986) <= '1';
    layer2_outputs(2987) <= '1';
    layer2_outputs(2988) <= layer1_outputs(5390);
    layer2_outputs(2989) <= layer1_outputs(4281);
    layer2_outputs(2990) <= '0';
    layer2_outputs(2991) <= layer1_outputs(471);
    layer2_outputs(2992) <= not(layer1_outputs(2975)) or (layer1_outputs(7037));
    layer2_outputs(2993) <= '1';
    layer2_outputs(2994) <= '1';
    layer2_outputs(2995) <= not(layer1_outputs(4679));
    layer2_outputs(2996) <= (layer1_outputs(4056)) and not (layer1_outputs(7492));
    layer2_outputs(2997) <= '1';
    layer2_outputs(2998) <= '0';
    layer2_outputs(2999) <= not(layer1_outputs(1683));
    layer2_outputs(3000) <= not(layer1_outputs(6625)) or (layer1_outputs(3711));
    layer2_outputs(3001) <= (layer1_outputs(4691)) and not (layer1_outputs(7138));
    layer2_outputs(3002) <= not((layer1_outputs(5967)) and (layer1_outputs(7656)));
    layer2_outputs(3003) <= '1';
    layer2_outputs(3004) <= not((layer1_outputs(6230)) or (layer1_outputs(6067)));
    layer2_outputs(3005) <= (layer1_outputs(2895)) and not (layer1_outputs(4052));
    layer2_outputs(3006) <= not(layer1_outputs(6949));
    layer2_outputs(3007) <= not((layer1_outputs(5393)) or (layer1_outputs(4232)));
    layer2_outputs(3008) <= (layer1_outputs(6247)) and (layer1_outputs(7177));
    layer2_outputs(3009) <= (layer1_outputs(2311)) and (layer1_outputs(6833));
    layer2_outputs(3010) <= (layer1_outputs(2598)) xor (layer1_outputs(2444));
    layer2_outputs(3011) <= (layer1_outputs(1590)) or (layer1_outputs(1098));
    layer2_outputs(3012) <= (layer1_outputs(1587)) and (layer1_outputs(2328));
    layer2_outputs(3013) <= (layer1_outputs(255)) and (layer1_outputs(7519));
    layer2_outputs(3014) <= '0';
    layer2_outputs(3015) <= layer1_outputs(7085);
    layer2_outputs(3016) <= (layer1_outputs(4307)) or (layer1_outputs(1978));
    layer2_outputs(3017) <= layer1_outputs(1149);
    layer2_outputs(3018) <= layer1_outputs(2390);
    layer2_outputs(3019) <= (layer1_outputs(6697)) or (layer1_outputs(356));
    layer2_outputs(3020) <= not((layer1_outputs(5598)) and (layer1_outputs(172)));
    layer2_outputs(3021) <= not(layer1_outputs(3571));
    layer2_outputs(3022) <= not((layer1_outputs(5269)) and (layer1_outputs(3272)));
    layer2_outputs(3023) <= not((layer1_outputs(7353)) and (layer1_outputs(5851)));
    layer2_outputs(3024) <= layer1_outputs(5737);
    layer2_outputs(3025) <= (layer1_outputs(6098)) and not (layer1_outputs(5600));
    layer2_outputs(3026) <= not((layer1_outputs(6025)) or (layer1_outputs(648)));
    layer2_outputs(3027) <= not(layer1_outputs(3804));
    layer2_outputs(3028) <= (layer1_outputs(6182)) and (layer1_outputs(4976));
    layer2_outputs(3029) <= not((layer1_outputs(3370)) xor (layer1_outputs(3337)));
    layer2_outputs(3030) <= not(layer1_outputs(4513)) or (layer1_outputs(4629));
    layer2_outputs(3031) <= not(layer1_outputs(7438)) or (layer1_outputs(6909));
    layer2_outputs(3032) <= (layer1_outputs(6591)) or (layer1_outputs(2252));
    layer2_outputs(3033) <= layer1_outputs(3638);
    layer2_outputs(3034) <= layer1_outputs(5088);
    layer2_outputs(3035) <= (layer1_outputs(3357)) and not (layer1_outputs(4155));
    layer2_outputs(3036) <= (layer1_outputs(212)) and not (layer1_outputs(466));
    layer2_outputs(3037) <= not(layer1_outputs(489)) or (layer1_outputs(3259));
    layer2_outputs(3038) <= not((layer1_outputs(1652)) and (layer1_outputs(4294)));
    layer2_outputs(3039) <= not((layer1_outputs(5787)) or (layer1_outputs(5348)));
    layer2_outputs(3040) <= (layer1_outputs(6036)) and (layer1_outputs(1083));
    layer2_outputs(3041) <= '1';
    layer2_outputs(3042) <= (layer1_outputs(568)) and not (layer1_outputs(4618));
    layer2_outputs(3043) <= not((layer1_outputs(4327)) or (layer1_outputs(3261)));
    layer2_outputs(3044) <= (layer1_outputs(1136)) and not (layer1_outputs(6680));
    layer2_outputs(3045) <= (layer1_outputs(2360)) and not (layer1_outputs(7284));
    layer2_outputs(3046) <= not(layer1_outputs(6296)) or (layer1_outputs(3280));
    layer2_outputs(3047) <= layer1_outputs(5106);
    layer2_outputs(3048) <= not(layer1_outputs(4280));
    layer2_outputs(3049) <= not(layer1_outputs(1901)) or (layer1_outputs(5287));
    layer2_outputs(3050) <= '0';
    layer2_outputs(3051) <= (layer1_outputs(3462)) or (layer1_outputs(3888));
    layer2_outputs(3052) <= '0';
    layer2_outputs(3053) <= '1';
    layer2_outputs(3054) <= '1';
    layer2_outputs(3055) <= not(layer1_outputs(7209)) or (layer1_outputs(2249));
    layer2_outputs(3056) <= '1';
    layer2_outputs(3057) <= not((layer1_outputs(3335)) or (layer1_outputs(4089)));
    layer2_outputs(3058) <= '1';
    layer2_outputs(3059) <= not(layer1_outputs(4194)) or (layer1_outputs(710));
    layer2_outputs(3060) <= (layer1_outputs(2248)) and (layer1_outputs(2469));
    layer2_outputs(3061) <= not(layer1_outputs(186));
    layer2_outputs(3062) <= '1';
    layer2_outputs(3063) <= (layer1_outputs(3159)) and not (layer1_outputs(4549));
    layer2_outputs(3064) <= (layer1_outputs(1526)) and not (layer1_outputs(6792));
    layer2_outputs(3065) <= not(layer1_outputs(7382));
    layer2_outputs(3066) <= '0';
    layer2_outputs(3067) <= layer1_outputs(6471);
    layer2_outputs(3068) <= not(layer1_outputs(1472));
    layer2_outputs(3069) <= not(layer1_outputs(1490));
    layer2_outputs(3070) <= not((layer1_outputs(71)) and (layer1_outputs(5837)));
    layer2_outputs(3071) <= (layer1_outputs(5610)) or (layer1_outputs(5586));
    layer2_outputs(3072) <= '0';
    layer2_outputs(3073) <= not(layer1_outputs(6866));
    layer2_outputs(3074) <= not(layer1_outputs(827)) or (layer1_outputs(6838));
    layer2_outputs(3075) <= '0';
    layer2_outputs(3076) <= not(layer1_outputs(2384));
    layer2_outputs(3077) <= not((layer1_outputs(1703)) and (layer1_outputs(6102)));
    layer2_outputs(3078) <= layer1_outputs(2972);
    layer2_outputs(3079) <= not(layer1_outputs(3770)) or (layer1_outputs(2699));
    layer2_outputs(3080) <= not(layer1_outputs(5883)) or (layer1_outputs(5270));
    layer2_outputs(3081) <= (layer1_outputs(3235)) and not (layer1_outputs(6861));
    layer2_outputs(3082) <= '0';
    layer2_outputs(3083) <= '1';
    layer2_outputs(3084) <= '0';
    layer2_outputs(3085) <= not(layer1_outputs(3663));
    layer2_outputs(3086) <= (layer1_outputs(7273)) and (layer1_outputs(934));
    layer2_outputs(3087) <= '1';
    layer2_outputs(3088) <= not(layer1_outputs(3897));
    layer2_outputs(3089) <= layer1_outputs(5609);
    layer2_outputs(3090) <= layer1_outputs(259);
    layer2_outputs(3091) <= not(layer1_outputs(3411)) or (layer1_outputs(3719));
    layer2_outputs(3092) <= not((layer1_outputs(5185)) and (layer1_outputs(2768)));
    layer2_outputs(3093) <= '0';
    layer2_outputs(3094) <= layer1_outputs(4370);
    layer2_outputs(3095) <= '1';
    layer2_outputs(3096) <= (layer1_outputs(1296)) or (layer1_outputs(7570));
    layer2_outputs(3097) <= (layer1_outputs(2083)) or (layer1_outputs(4646));
    layer2_outputs(3098) <= not((layer1_outputs(4834)) and (layer1_outputs(6296)));
    layer2_outputs(3099) <= '1';
    layer2_outputs(3100) <= (layer1_outputs(1693)) and (layer1_outputs(1877));
    layer2_outputs(3101) <= '0';
    layer2_outputs(3102) <= layer1_outputs(7155);
    layer2_outputs(3103) <= (layer1_outputs(5838)) or (layer1_outputs(1450));
    layer2_outputs(3104) <= '0';
    layer2_outputs(3105) <= layer1_outputs(4430);
    layer2_outputs(3106) <= layer1_outputs(394);
    layer2_outputs(3107) <= (layer1_outputs(4054)) xor (layer1_outputs(7495));
    layer2_outputs(3108) <= not(layer1_outputs(6398)) or (layer1_outputs(5957));
    layer2_outputs(3109) <= (layer1_outputs(7613)) xor (layer1_outputs(5392));
    layer2_outputs(3110) <= not(layer1_outputs(3257));
    layer2_outputs(3111) <= layer1_outputs(2887);
    layer2_outputs(3112) <= '0';
    layer2_outputs(3113) <= layer1_outputs(2074);
    layer2_outputs(3114) <= not(layer1_outputs(134)) or (layer1_outputs(1970));
    layer2_outputs(3115) <= not(layer1_outputs(2050)) or (layer1_outputs(6712));
    layer2_outputs(3116) <= '0';
    layer2_outputs(3117) <= layer1_outputs(5123);
    layer2_outputs(3118) <= not(layer1_outputs(3319));
    layer2_outputs(3119) <= '1';
    layer2_outputs(3120) <= (layer1_outputs(6537)) and not (layer1_outputs(3325));
    layer2_outputs(3121) <= (layer1_outputs(3932)) and (layer1_outputs(501));
    layer2_outputs(3122) <= not(layer1_outputs(1463)) or (layer1_outputs(7062));
    layer2_outputs(3123) <= not(layer1_outputs(3134)) or (layer1_outputs(359));
    layer2_outputs(3124) <= '0';
    layer2_outputs(3125) <= (layer1_outputs(1694)) and not (layer1_outputs(3487));
    layer2_outputs(3126) <= not((layer1_outputs(1617)) and (layer1_outputs(2989)));
    layer2_outputs(3127) <= not(layer1_outputs(124));
    layer2_outputs(3128) <= layer1_outputs(1177);
    layer2_outputs(3129) <= not(layer1_outputs(7590));
    layer2_outputs(3130) <= layer1_outputs(1281);
    layer2_outputs(3131) <= not((layer1_outputs(5916)) and (layer1_outputs(2273)));
    layer2_outputs(3132) <= not((layer1_outputs(6895)) or (layer1_outputs(1002)));
    layer2_outputs(3133) <= layer1_outputs(2199);
    layer2_outputs(3134) <= layer1_outputs(1592);
    layer2_outputs(3135) <= '1';
    layer2_outputs(3136) <= (layer1_outputs(6982)) or (layer1_outputs(1840));
    layer2_outputs(3137) <= '1';
    layer2_outputs(3138) <= (layer1_outputs(6067)) and not (layer1_outputs(6306));
    layer2_outputs(3139) <= layer1_outputs(156);
    layer2_outputs(3140) <= layer1_outputs(921);
    layer2_outputs(3141) <= not(layer1_outputs(6454));
    layer2_outputs(3142) <= not(layer1_outputs(3451)) or (layer1_outputs(700));
    layer2_outputs(3143) <= not(layer1_outputs(150));
    layer2_outputs(3144) <= layer1_outputs(3826);
    layer2_outputs(3145) <= not(layer1_outputs(5532)) or (layer1_outputs(2289));
    layer2_outputs(3146) <= (layer1_outputs(1736)) and not (layer1_outputs(2772));
    layer2_outputs(3147) <= not((layer1_outputs(7028)) or (layer1_outputs(6456)));
    layer2_outputs(3148) <= layer1_outputs(3424);
    layer2_outputs(3149) <= not((layer1_outputs(7010)) and (layer1_outputs(1504)));
    layer2_outputs(3150) <= not(layer1_outputs(1029));
    layer2_outputs(3151) <= not((layer1_outputs(806)) or (layer1_outputs(1579)));
    layer2_outputs(3152) <= not(layer1_outputs(5796)) or (layer1_outputs(4789));
    layer2_outputs(3153) <= '0';
    layer2_outputs(3154) <= layer1_outputs(7325);
    layer2_outputs(3155) <= layer1_outputs(2418);
    layer2_outputs(3156) <= not((layer1_outputs(7619)) or (layer1_outputs(4392)));
    layer2_outputs(3157) <= (layer1_outputs(5259)) and not (layer1_outputs(3384));
    layer2_outputs(3158) <= (layer1_outputs(5939)) and not (layer1_outputs(144));
    layer2_outputs(3159) <= '1';
    layer2_outputs(3160) <= layer1_outputs(661);
    layer2_outputs(3161) <= (layer1_outputs(5145)) or (layer1_outputs(2440));
    layer2_outputs(3162) <= (layer1_outputs(7022)) and not (layer1_outputs(5466));
    layer2_outputs(3163) <= layer1_outputs(3370);
    layer2_outputs(3164) <= not(layer1_outputs(5131));
    layer2_outputs(3165) <= not((layer1_outputs(3222)) or (layer1_outputs(1420)));
    layer2_outputs(3166) <= layer1_outputs(6832);
    layer2_outputs(3167) <= (layer1_outputs(1008)) and not (layer1_outputs(75));
    layer2_outputs(3168) <= layer1_outputs(6586);
    layer2_outputs(3169) <= not(layer1_outputs(317));
    layer2_outputs(3170) <= not(layer1_outputs(6338));
    layer2_outputs(3171) <= '0';
    layer2_outputs(3172) <= not((layer1_outputs(2319)) and (layer1_outputs(5625)));
    layer2_outputs(3173) <= '0';
    layer2_outputs(3174) <= not((layer1_outputs(6725)) or (layer1_outputs(2100)));
    layer2_outputs(3175) <= '1';
    layer2_outputs(3176) <= (layer1_outputs(6582)) xor (layer1_outputs(2450));
    layer2_outputs(3177) <= '1';
    layer2_outputs(3178) <= layer1_outputs(5744);
    layer2_outputs(3179) <= not(layer1_outputs(9));
    layer2_outputs(3180) <= (layer1_outputs(2532)) or (layer1_outputs(2222));
    layer2_outputs(3181) <= not(layer1_outputs(5418)) or (layer1_outputs(7016));
    layer2_outputs(3182) <= layer1_outputs(493);
    layer2_outputs(3183) <= layer1_outputs(5199);
    layer2_outputs(3184) <= (layer1_outputs(5297)) and not (layer1_outputs(3957));
    layer2_outputs(3185) <= '0';
    layer2_outputs(3186) <= layer1_outputs(4161);
    layer2_outputs(3187) <= '1';
    layer2_outputs(3188) <= '1';
    layer2_outputs(3189) <= not(layer1_outputs(1447)) or (layer1_outputs(5241));
    layer2_outputs(3190) <= layer1_outputs(4732);
    layer2_outputs(3191) <= '0';
    layer2_outputs(3192) <= (layer1_outputs(2230)) and not (layer1_outputs(6260));
    layer2_outputs(3193) <= (layer1_outputs(4722)) or (layer1_outputs(799));
    layer2_outputs(3194) <= not(layer1_outputs(2004));
    layer2_outputs(3195) <= not(layer1_outputs(1931));
    layer2_outputs(3196) <= not(layer1_outputs(6465));
    layer2_outputs(3197) <= (layer1_outputs(845)) and not (layer1_outputs(2575));
    layer2_outputs(3198) <= not(layer1_outputs(7358));
    layer2_outputs(3199) <= (layer1_outputs(6455)) xor (layer1_outputs(5961));
    layer2_outputs(3200) <= not(layer1_outputs(3540));
    layer2_outputs(3201) <= not(layer1_outputs(7274));
    layer2_outputs(3202) <= not((layer1_outputs(4653)) or (layer1_outputs(7562)));
    layer2_outputs(3203) <= (layer1_outputs(4954)) and not (layer1_outputs(4244));
    layer2_outputs(3204) <= not(layer1_outputs(112)) or (layer1_outputs(519));
    layer2_outputs(3205) <= (layer1_outputs(4595)) or (layer1_outputs(5108));
    layer2_outputs(3206) <= not(layer1_outputs(5224)) or (layer1_outputs(7100));
    layer2_outputs(3207) <= not(layer1_outputs(1512));
    layer2_outputs(3208) <= not((layer1_outputs(4501)) or (layer1_outputs(1556)));
    layer2_outputs(3209) <= (layer1_outputs(2066)) or (layer1_outputs(4812));
    layer2_outputs(3210) <= not(layer1_outputs(1935));
    layer2_outputs(3211) <= not(layer1_outputs(5601));
    layer2_outputs(3212) <= not(layer1_outputs(3160));
    layer2_outputs(3213) <= '0';
    layer2_outputs(3214) <= (layer1_outputs(6497)) xor (layer1_outputs(397));
    layer2_outputs(3215) <= '1';
    layer2_outputs(3216) <= not(layer1_outputs(3272));
    layer2_outputs(3217) <= not(layer1_outputs(2641));
    layer2_outputs(3218) <= not((layer1_outputs(1750)) or (layer1_outputs(4819)));
    layer2_outputs(3219) <= not((layer1_outputs(2368)) and (layer1_outputs(7135)));
    layer2_outputs(3220) <= (layer1_outputs(2059)) and not (layer1_outputs(6290));
    layer2_outputs(3221) <= not(layer1_outputs(6668));
    layer2_outputs(3222) <= not(layer1_outputs(42)) or (layer1_outputs(3176));
    layer2_outputs(3223) <= not((layer1_outputs(7270)) and (layer1_outputs(1108)));
    layer2_outputs(3224) <= not(layer1_outputs(1387));
    layer2_outputs(3225) <= layer1_outputs(1314);
    layer2_outputs(3226) <= not(layer1_outputs(3533));
    layer2_outputs(3227) <= (layer1_outputs(6606)) and (layer1_outputs(2844));
    layer2_outputs(3228) <= layer1_outputs(749);
    layer2_outputs(3229) <= (layer1_outputs(3174)) and not (layer1_outputs(7246));
    layer2_outputs(3230) <= '0';
    layer2_outputs(3231) <= not(layer1_outputs(5195)) or (layer1_outputs(1891));
    layer2_outputs(3232) <= '1';
    layer2_outputs(3233) <= layer1_outputs(2315);
    layer2_outputs(3234) <= not((layer1_outputs(6940)) or (layer1_outputs(1267)));
    layer2_outputs(3235) <= not(layer1_outputs(4403)) or (layer1_outputs(6780));
    layer2_outputs(3236) <= not((layer1_outputs(5645)) xor (layer1_outputs(893)));
    layer2_outputs(3237) <= layer1_outputs(2736);
    layer2_outputs(3238) <= not(layer1_outputs(6272));
    layer2_outputs(3239) <= '1';
    layer2_outputs(3240) <= not(layer1_outputs(5302));
    layer2_outputs(3241) <= (layer1_outputs(982)) and not (layer1_outputs(601));
    layer2_outputs(3242) <= layer1_outputs(3150);
    layer2_outputs(3243) <= not(layer1_outputs(3302));
    layer2_outputs(3244) <= '1';
    layer2_outputs(3245) <= (layer1_outputs(3102)) and (layer1_outputs(1577));
    layer2_outputs(3246) <= not(layer1_outputs(2055)) or (layer1_outputs(371));
    layer2_outputs(3247) <= (layer1_outputs(3775)) xor (layer1_outputs(2642));
    layer2_outputs(3248) <= (layer1_outputs(5455)) and not (layer1_outputs(3715));
    layer2_outputs(3249) <= not((layer1_outputs(5671)) or (layer1_outputs(3265)));
    layer2_outputs(3250) <= '0';
    layer2_outputs(3251) <= not(layer1_outputs(6567));
    layer2_outputs(3252) <= (layer1_outputs(4410)) and (layer1_outputs(7074));
    layer2_outputs(3253) <= (layer1_outputs(6274)) and (layer1_outputs(5512));
    layer2_outputs(3254) <= '1';
    layer2_outputs(3255) <= not(layer1_outputs(1081)) or (layer1_outputs(6643));
    layer2_outputs(3256) <= (layer1_outputs(6415)) and not (layer1_outputs(1467));
    layer2_outputs(3257) <= (layer1_outputs(1156)) or (layer1_outputs(4415));
    layer2_outputs(3258) <= not((layer1_outputs(1851)) and (layer1_outputs(2908)));
    layer2_outputs(3259) <= (layer1_outputs(1567)) and (layer1_outputs(1279));
    layer2_outputs(3260) <= not((layer1_outputs(1971)) or (layer1_outputs(2786)));
    layer2_outputs(3261) <= (layer1_outputs(2079)) and (layer1_outputs(5613));
    layer2_outputs(3262) <= '1';
    layer2_outputs(3263) <= '1';
    layer2_outputs(3264) <= layer1_outputs(1940);
    layer2_outputs(3265) <= not(layer1_outputs(4755)) or (layer1_outputs(7358));
    layer2_outputs(3266) <= '0';
    layer2_outputs(3267) <= not(layer1_outputs(6495));
    layer2_outputs(3268) <= not(layer1_outputs(3387)) or (layer1_outputs(4508));
    layer2_outputs(3269) <= (layer1_outputs(2206)) and not (layer1_outputs(1088));
    layer2_outputs(3270) <= not(layer1_outputs(4708));
    layer2_outputs(3271) <= not((layer1_outputs(2640)) or (layer1_outputs(2040)));
    layer2_outputs(3272) <= not((layer1_outputs(2833)) and (layer1_outputs(4535)));
    layer2_outputs(3273) <= not(layer1_outputs(3495));
    layer2_outputs(3274) <= layer1_outputs(4963);
    layer2_outputs(3275) <= (layer1_outputs(353)) and (layer1_outputs(6462));
    layer2_outputs(3276) <= layer1_outputs(2989);
    layer2_outputs(3277) <= (layer1_outputs(6346)) xor (layer1_outputs(1798));
    layer2_outputs(3278) <= not(layer1_outputs(1255));
    layer2_outputs(3279) <= (layer1_outputs(1224)) and not (layer1_outputs(5663));
    layer2_outputs(3280) <= not(layer1_outputs(176)) or (layer1_outputs(3456));
    layer2_outputs(3281) <= '1';
    layer2_outputs(3282) <= not(layer1_outputs(200)) or (layer1_outputs(1521));
    layer2_outputs(3283) <= '1';
    layer2_outputs(3284) <= not(layer1_outputs(7649)) or (layer1_outputs(7494));
    layer2_outputs(3285) <= (layer1_outputs(5197)) and (layer1_outputs(6830));
    layer2_outputs(3286) <= not(layer1_outputs(5762)) or (layer1_outputs(3288));
    layer2_outputs(3287) <= (layer1_outputs(2132)) and not (layer1_outputs(6680));
    layer2_outputs(3288) <= not(layer1_outputs(373));
    layer2_outputs(3289) <= not(layer1_outputs(2653)) or (layer1_outputs(5184));
    layer2_outputs(3290) <= not((layer1_outputs(2839)) and (layer1_outputs(3361)));
    layer2_outputs(3291) <= (layer1_outputs(877)) and (layer1_outputs(6180));
    layer2_outputs(3292) <= (layer1_outputs(1865)) or (layer1_outputs(2717));
    layer2_outputs(3293) <= '0';
    layer2_outputs(3294) <= not((layer1_outputs(6557)) and (layer1_outputs(4956)));
    layer2_outputs(3295) <= not((layer1_outputs(6243)) or (layer1_outputs(6184)));
    layer2_outputs(3296) <= not((layer1_outputs(1714)) and (layer1_outputs(2098)));
    layer2_outputs(3297) <= '1';
    layer2_outputs(3298) <= '0';
    layer2_outputs(3299) <= (layer1_outputs(529)) and (layer1_outputs(911));
    layer2_outputs(3300) <= '0';
    layer2_outputs(3301) <= not(layer1_outputs(6591));
    layer2_outputs(3302) <= not((layer1_outputs(6384)) and (layer1_outputs(2543)));
    layer2_outputs(3303) <= not((layer1_outputs(4262)) or (layer1_outputs(2628)));
    layer2_outputs(3304) <= not(layer1_outputs(2998));
    layer2_outputs(3305) <= not((layer1_outputs(222)) or (layer1_outputs(1860)));
    layer2_outputs(3306) <= (layer1_outputs(3852)) or (layer1_outputs(2583));
    layer2_outputs(3307) <= not(layer1_outputs(3188)) or (layer1_outputs(6325));
    layer2_outputs(3308) <= not(layer1_outputs(1987));
    layer2_outputs(3309) <= (layer1_outputs(7419)) and not (layer1_outputs(2911));
    layer2_outputs(3310) <= not(layer1_outputs(2917)) or (layer1_outputs(5815));
    layer2_outputs(3311) <= layer1_outputs(23);
    layer2_outputs(3312) <= not(layer1_outputs(3108));
    layer2_outputs(3313) <= layer1_outputs(3647);
    layer2_outputs(3314) <= (layer1_outputs(1466)) and not (layer1_outputs(2395));
    layer2_outputs(3315) <= not((layer1_outputs(7180)) and (layer1_outputs(7202)));
    layer2_outputs(3316) <= '1';
    layer2_outputs(3317) <= '1';
    layer2_outputs(3318) <= layer1_outputs(7287);
    layer2_outputs(3319) <= not((layer1_outputs(3206)) and (layer1_outputs(5294)));
    layer2_outputs(3320) <= not((layer1_outputs(2055)) xor (layer1_outputs(2552)));
    layer2_outputs(3321) <= layer1_outputs(6534);
    layer2_outputs(3322) <= layer1_outputs(870);
    layer2_outputs(3323) <= not(layer1_outputs(926)) or (layer1_outputs(7120));
    layer2_outputs(3324) <= layer1_outputs(5253);
    layer2_outputs(3325) <= not(layer1_outputs(2893));
    layer2_outputs(3326) <= not(layer1_outputs(5813));
    layer2_outputs(3327) <= (layer1_outputs(4819)) or (layer1_outputs(5872));
    layer2_outputs(3328) <= layer1_outputs(3442);
    layer2_outputs(3329) <= not(layer1_outputs(5015)) or (layer1_outputs(4627));
    layer2_outputs(3330) <= not((layer1_outputs(7313)) or (layer1_outputs(5875)));
    layer2_outputs(3331) <= (layer1_outputs(7002)) or (layer1_outputs(6676));
    layer2_outputs(3332) <= not(layer1_outputs(3486)) or (layer1_outputs(3198));
    layer2_outputs(3333) <= (layer1_outputs(724)) and not (layer1_outputs(3347));
    layer2_outputs(3334) <= '1';
    layer2_outputs(3335) <= layer1_outputs(4477);
    layer2_outputs(3336) <= (layer1_outputs(7179)) and not (layer1_outputs(7175));
    layer2_outputs(3337) <= not(layer1_outputs(5943));
    layer2_outputs(3338) <= (layer1_outputs(5201)) and not (layer1_outputs(1787));
    layer2_outputs(3339) <= layer1_outputs(226);
    layer2_outputs(3340) <= (layer1_outputs(1799)) and (layer1_outputs(7671));
    layer2_outputs(3341) <= not(layer1_outputs(6575));
    layer2_outputs(3342) <= (layer1_outputs(7160)) and not (layer1_outputs(1417));
    layer2_outputs(3343) <= not(layer1_outputs(5977));
    layer2_outputs(3344) <= not(layer1_outputs(4879)) or (layer1_outputs(4540));
    layer2_outputs(3345) <= '1';
    layer2_outputs(3346) <= not((layer1_outputs(1412)) xor (layer1_outputs(2126)));
    layer2_outputs(3347) <= not(layer1_outputs(5797));
    layer2_outputs(3348) <= '0';
    layer2_outputs(3349) <= layer1_outputs(695);
    layer2_outputs(3350) <= not(layer1_outputs(6305)) or (layer1_outputs(7147));
    layer2_outputs(3351) <= (layer1_outputs(2678)) and not (layer1_outputs(6759));
    layer2_outputs(3352) <= '1';
    layer2_outputs(3353) <= not((layer1_outputs(4436)) or (layer1_outputs(966)));
    layer2_outputs(3354) <= '0';
    layer2_outputs(3355) <= not(layer1_outputs(4551)) or (layer1_outputs(1894));
    layer2_outputs(3356) <= layer1_outputs(6183);
    layer2_outputs(3357) <= (layer1_outputs(587)) and not (layer1_outputs(3332));
    layer2_outputs(3358) <= layer1_outputs(5535);
    layer2_outputs(3359) <= not(layer1_outputs(4286));
    layer2_outputs(3360) <= layer1_outputs(113);
    layer2_outputs(3361) <= (layer1_outputs(3992)) and not (layer1_outputs(6616));
    layer2_outputs(3362) <= not((layer1_outputs(1905)) or (layer1_outputs(4144)));
    layer2_outputs(3363) <= '1';
    layer2_outputs(3364) <= '1';
    layer2_outputs(3365) <= (layer1_outputs(976)) and (layer1_outputs(7510));
    layer2_outputs(3366) <= (layer1_outputs(4396)) and (layer1_outputs(2110));
    layer2_outputs(3367) <= not(layer1_outputs(5769)) or (layer1_outputs(5548));
    layer2_outputs(3368) <= not(layer1_outputs(71));
    layer2_outputs(3369) <= not(layer1_outputs(3500)) or (layer1_outputs(6083));
    layer2_outputs(3370) <= '1';
    layer2_outputs(3371) <= layer1_outputs(4019);
    layer2_outputs(3372) <= (layer1_outputs(1425)) or (layer1_outputs(5758));
    layer2_outputs(3373) <= (layer1_outputs(2422)) or (layer1_outputs(6722));
    layer2_outputs(3374) <= (layer1_outputs(1302)) and not (layer1_outputs(5298));
    layer2_outputs(3375) <= (layer1_outputs(1754)) or (layer1_outputs(949));
    layer2_outputs(3376) <= (layer1_outputs(3142)) and not (layer1_outputs(5293));
    layer2_outputs(3377) <= not(layer1_outputs(1929));
    layer2_outputs(3378) <= not((layer1_outputs(6421)) xor (layer1_outputs(524)));
    layer2_outputs(3379) <= '0';
    layer2_outputs(3380) <= layer1_outputs(2899);
    layer2_outputs(3381) <= not(layer1_outputs(3429)) or (layer1_outputs(2142));
    layer2_outputs(3382) <= not(layer1_outputs(6631));
    layer2_outputs(3383) <= (layer1_outputs(7451)) and not (layer1_outputs(5246));
    layer2_outputs(3384) <= (layer1_outputs(4768)) and not (layer1_outputs(2639));
    layer2_outputs(3385) <= not(layer1_outputs(1043));
    layer2_outputs(3386) <= (layer1_outputs(5526)) xor (layer1_outputs(4419));
    layer2_outputs(3387) <= not(layer1_outputs(3316)) or (layer1_outputs(5055));
    layer2_outputs(3388) <= layer1_outputs(3385);
    layer2_outputs(3389) <= layer1_outputs(6535);
    layer2_outputs(3390) <= (layer1_outputs(4939)) and not (layer1_outputs(6513));
    layer2_outputs(3391) <= '1';
    layer2_outputs(3392) <= not((layer1_outputs(2968)) or (layer1_outputs(5964)));
    layer2_outputs(3393) <= layer1_outputs(5504);
    layer2_outputs(3394) <= not(layer1_outputs(139));
    layer2_outputs(3395) <= '0';
    layer2_outputs(3396) <= (layer1_outputs(6937)) and not (layer1_outputs(3361));
    layer2_outputs(3397) <= not(layer1_outputs(2568));
    layer2_outputs(3398) <= (layer1_outputs(3656)) and (layer1_outputs(4590));
    layer2_outputs(3399) <= '1';
    layer2_outputs(3400) <= layer1_outputs(3687);
    layer2_outputs(3401) <= not(layer1_outputs(824)) or (layer1_outputs(1760));
    layer2_outputs(3402) <= (layer1_outputs(6220)) and not (layer1_outputs(6154));
    layer2_outputs(3403) <= not(layer1_outputs(3923)) or (layer1_outputs(4178));
    layer2_outputs(3404) <= (layer1_outputs(4660)) xor (layer1_outputs(406));
    layer2_outputs(3405) <= '0';
    layer2_outputs(3406) <= (layer1_outputs(2810)) and (layer1_outputs(7255));
    layer2_outputs(3407) <= not(layer1_outputs(3098)) or (layer1_outputs(4168));
    layer2_outputs(3408) <= (layer1_outputs(36)) and not (layer1_outputs(4980));
    layer2_outputs(3409) <= (layer1_outputs(6798)) and not (layer1_outputs(1925));
    layer2_outputs(3410) <= not(layer1_outputs(3484)) or (layer1_outputs(7112));
    layer2_outputs(3411) <= '0';
    layer2_outputs(3412) <= not((layer1_outputs(2967)) and (layer1_outputs(7310)));
    layer2_outputs(3413) <= '0';
    layer2_outputs(3414) <= not(layer1_outputs(5318)) or (layer1_outputs(3073));
    layer2_outputs(3415) <= '0';
    layer2_outputs(3416) <= not(layer1_outputs(4600));
    layer2_outputs(3417) <= not((layer1_outputs(6721)) or (layer1_outputs(1781)));
    layer2_outputs(3418) <= not(layer1_outputs(2413));
    layer2_outputs(3419) <= (layer1_outputs(7323)) and not (layer1_outputs(5380));
    layer2_outputs(3420) <= (layer1_outputs(7218)) and not (layer1_outputs(1963));
    layer2_outputs(3421) <= '0';
    layer2_outputs(3422) <= not((layer1_outputs(3727)) and (layer1_outputs(5276)));
    layer2_outputs(3423) <= (layer1_outputs(6634)) or (layer1_outputs(7654));
    layer2_outputs(3424) <= (layer1_outputs(6945)) and not (layer1_outputs(3264));
    layer2_outputs(3425) <= not(layer1_outputs(5853)) or (layer1_outputs(4822));
    layer2_outputs(3426) <= layer1_outputs(1980);
    layer2_outputs(3427) <= (layer1_outputs(7168)) and not (layer1_outputs(4848));
    layer2_outputs(3428) <= not((layer1_outputs(3475)) or (layer1_outputs(3212)));
    layer2_outputs(3429) <= layer1_outputs(154);
    layer2_outputs(3430) <= not((layer1_outputs(4931)) or (layer1_outputs(1161)));
    layer2_outputs(3431) <= not((layer1_outputs(998)) or (layer1_outputs(5851)));
    layer2_outputs(3432) <= layer1_outputs(1127);
    layer2_outputs(3433) <= (layer1_outputs(4852)) xor (layer1_outputs(3017));
    layer2_outputs(3434) <= not(layer1_outputs(5550)) or (layer1_outputs(1491));
    layer2_outputs(3435) <= layer1_outputs(6979);
    layer2_outputs(3436) <= '1';
    layer2_outputs(3437) <= layer1_outputs(7421);
    layer2_outputs(3438) <= '0';
    layer2_outputs(3439) <= not(layer1_outputs(5893));
    layer2_outputs(3440) <= not(layer1_outputs(6648));
    layer2_outputs(3441) <= layer1_outputs(5342);
    layer2_outputs(3442) <= layer1_outputs(4384);
    layer2_outputs(3443) <= layer1_outputs(1989);
    layer2_outputs(3444) <= (layer1_outputs(3710)) and not (layer1_outputs(6447));
    layer2_outputs(3445) <= not(layer1_outputs(2923));
    layer2_outputs(3446) <= not((layer1_outputs(1593)) and (layer1_outputs(1032)));
    layer2_outputs(3447) <= layer1_outputs(4572);
    layer2_outputs(3448) <= layer1_outputs(7336);
    layer2_outputs(3449) <= not(layer1_outputs(163)) or (layer1_outputs(7073));
    layer2_outputs(3450) <= layer1_outputs(7466);
    layer2_outputs(3451) <= not((layer1_outputs(4263)) and (layer1_outputs(792)));
    layer2_outputs(3452) <= not(layer1_outputs(740));
    layer2_outputs(3453) <= not(layer1_outputs(5369));
    layer2_outputs(3454) <= not(layer1_outputs(5248)) or (layer1_outputs(5395));
    layer2_outputs(3455) <= not(layer1_outputs(3878));
    layer2_outputs(3456) <= not(layer1_outputs(6929));
    layer2_outputs(3457) <= layer1_outputs(1968);
    layer2_outputs(3458) <= not(layer1_outputs(1452)) or (layer1_outputs(1832));
    layer2_outputs(3459) <= (layer1_outputs(2131)) and (layer1_outputs(1228));
    layer2_outputs(3460) <= (layer1_outputs(6060)) or (layer1_outputs(4082));
    layer2_outputs(3461) <= (layer1_outputs(4905)) and (layer1_outputs(6856));
    layer2_outputs(3462) <= '1';
    layer2_outputs(3463) <= '1';
    layer2_outputs(3464) <= '0';
    layer2_outputs(3465) <= '1';
    layer2_outputs(3466) <= not(layer1_outputs(2040));
    layer2_outputs(3467) <= (layer1_outputs(3060)) and (layer1_outputs(2821));
    layer2_outputs(3468) <= not((layer1_outputs(1517)) or (layer1_outputs(3920)));
    layer2_outputs(3469) <= not((layer1_outputs(7374)) and (layer1_outputs(7394)));
    layer2_outputs(3470) <= not(layer1_outputs(4724)) or (layer1_outputs(7148));
    layer2_outputs(3471) <= layer1_outputs(4084);
    layer2_outputs(3472) <= not(layer1_outputs(4581)) or (layer1_outputs(443));
    layer2_outputs(3473) <= not((layer1_outputs(6382)) and (layer1_outputs(305)));
    layer2_outputs(3474) <= layer1_outputs(7434);
    layer2_outputs(3475) <= not((layer1_outputs(2383)) and (layer1_outputs(2863)));
    layer2_outputs(3476) <= not(layer1_outputs(2578)) or (layer1_outputs(4640));
    layer2_outputs(3477) <= not(layer1_outputs(6320)) or (layer1_outputs(402));
    layer2_outputs(3478) <= layer1_outputs(6264);
    layer2_outputs(3479) <= (layer1_outputs(4605)) and (layer1_outputs(6559));
    layer2_outputs(3480) <= not(layer1_outputs(1689)) or (layer1_outputs(598));
    layer2_outputs(3481) <= '0';
    layer2_outputs(3482) <= not(layer1_outputs(3359)) or (layer1_outputs(1273));
    layer2_outputs(3483) <= (layer1_outputs(4349)) and not (layer1_outputs(1769));
    layer2_outputs(3484) <= layer1_outputs(4662);
    layer2_outputs(3485) <= not(layer1_outputs(5032));
    layer2_outputs(3486) <= (layer1_outputs(3962)) and not (layer1_outputs(5701));
    layer2_outputs(3487) <= not(layer1_outputs(5777));
    layer2_outputs(3488) <= not(layer1_outputs(3409));
    layer2_outputs(3489) <= not(layer1_outputs(3406));
    layer2_outputs(3490) <= not(layer1_outputs(4223));
    layer2_outputs(3491) <= (layer1_outputs(7101)) and not (layer1_outputs(5506));
    layer2_outputs(3492) <= not(layer1_outputs(6520)) or (layer1_outputs(1547));
    layer2_outputs(3493) <= (layer1_outputs(6975)) and (layer1_outputs(3981));
    layer2_outputs(3494) <= (layer1_outputs(2350)) and not (layer1_outputs(2697));
    layer2_outputs(3495) <= layer1_outputs(1862);
    layer2_outputs(3496) <= not(layer1_outputs(1431));
    layer2_outputs(3497) <= '1';
    layer2_outputs(3498) <= not(layer1_outputs(1337)) or (layer1_outputs(6370));
    layer2_outputs(3499) <= (layer1_outputs(4413)) xor (layer1_outputs(691));
    layer2_outputs(3500) <= (layer1_outputs(380)) and not (layer1_outputs(6988));
    layer2_outputs(3501) <= '0';
    layer2_outputs(3502) <= not(layer1_outputs(438));
    layer2_outputs(3503) <= not(layer1_outputs(2614)) or (layer1_outputs(886));
    layer2_outputs(3504) <= '0';
    layer2_outputs(3505) <= (layer1_outputs(4227)) and (layer1_outputs(728));
    layer2_outputs(3506) <= (layer1_outputs(6337)) and not (layer1_outputs(2667));
    layer2_outputs(3507) <= not((layer1_outputs(5169)) and (layer1_outputs(6047)));
    layer2_outputs(3508) <= not(layer1_outputs(3784));
    layer2_outputs(3509) <= (layer1_outputs(3695)) and not (layer1_outputs(2876));
    layer2_outputs(3510) <= '1';
    layer2_outputs(3511) <= (layer1_outputs(5859)) and (layer1_outputs(1464));
    layer2_outputs(3512) <= layer1_outputs(6961);
    layer2_outputs(3513) <= not(layer1_outputs(7649));
    layer2_outputs(3514) <= '0';
    layer2_outputs(3515) <= not(layer1_outputs(5094));
    layer2_outputs(3516) <= layer1_outputs(2870);
    layer2_outputs(3517) <= not(layer1_outputs(3953));
    layer2_outputs(3518) <= layer1_outputs(927);
    layer2_outputs(3519) <= layer1_outputs(5226);
    layer2_outputs(3520) <= not(layer1_outputs(843)) or (layer1_outputs(1888));
    layer2_outputs(3521) <= (layer1_outputs(3136)) and not (layer1_outputs(6112));
    layer2_outputs(3522) <= not(layer1_outputs(141));
    layer2_outputs(3523) <= (layer1_outputs(4951)) and (layer1_outputs(574));
    layer2_outputs(3524) <= '1';
    layer2_outputs(3525) <= not(layer1_outputs(1318)) or (layer1_outputs(5765));
    layer2_outputs(3526) <= not(layer1_outputs(4261)) or (layer1_outputs(1920));
    layer2_outputs(3527) <= '0';
    layer2_outputs(3528) <= layer1_outputs(5072);
    layer2_outputs(3529) <= not((layer1_outputs(1646)) and (layer1_outputs(6308)));
    layer2_outputs(3530) <= layer1_outputs(1404);
    layer2_outputs(3531) <= not(layer1_outputs(2041)) or (layer1_outputs(633));
    layer2_outputs(3532) <= (layer1_outputs(2389)) and (layer1_outputs(1402));
    layer2_outputs(3533) <= (layer1_outputs(6815)) and (layer1_outputs(2540));
    layer2_outputs(3534) <= '0';
    layer2_outputs(3535) <= not(layer1_outputs(3219)) or (layer1_outputs(3904));
    layer2_outputs(3536) <= not(layer1_outputs(5037)) or (layer1_outputs(4429));
    layer2_outputs(3537) <= (layer1_outputs(5693)) and not (layer1_outputs(2555));
    layer2_outputs(3538) <= '0';
    layer2_outputs(3539) <= '1';
    layer2_outputs(3540) <= layer1_outputs(721);
    layer2_outputs(3541) <= (layer1_outputs(6757)) and not (layer1_outputs(2673));
    layer2_outputs(3542) <= not((layer1_outputs(4651)) xor (layer1_outputs(837)));
    layer2_outputs(3543) <= not(layer1_outputs(2555));
    layer2_outputs(3544) <= not(layer1_outputs(2351));
    layer2_outputs(3545) <= (layer1_outputs(5257)) and not (layer1_outputs(187));
    layer2_outputs(3546) <= '0';
    layer2_outputs(3547) <= not((layer1_outputs(2430)) and (layer1_outputs(6181)));
    layer2_outputs(3548) <= layer1_outputs(6390);
    layer2_outputs(3549) <= not((layer1_outputs(3835)) and (layer1_outputs(709)));
    layer2_outputs(3550) <= not(layer1_outputs(1541)) or (layer1_outputs(3336));
    layer2_outputs(3551) <= '1';
    layer2_outputs(3552) <= layer1_outputs(3616);
    layer2_outputs(3553) <= layer1_outputs(1191);
    layer2_outputs(3554) <= (layer1_outputs(4046)) and (layer1_outputs(5652));
    layer2_outputs(3555) <= not(layer1_outputs(7455)) or (layer1_outputs(4399));
    layer2_outputs(3556) <= (layer1_outputs(4191)) or (layer1_outputs(6592));
    layer2_outputs(3557) <= not(layer1_outputs(2666)) or (layer1_outputs(4838));
    layer2_outputs(3558) <= layer1_outputs(4616);
    layer2_outputs(3559) <= not(layer1_outputs(7512));
    layer2_outputs(3560) <= (layer1_outputs(805)) and not (layer1_outputs(3772));
    layer2_outputs(3561) <= not(layer1_outputs(5861));
    layer2_outputs(3562) <= not(layer1_outputs(2299));
    layer2_outputs(3563) <= not(layer1_outputs(7246));
    layer2_outputs(3564) <= not((layer1_outputs(5566)) and (layer1_outputs(1876)));
    layer2_outputs(3565) <= layer1_outputs(1119);
    layer2_outputs(3566) <= (layer1_outputs(2509)) and not (layer1_outputs(3935));
    layer2_outputs(3567) <= not(layer1_outputs(4941)) or (layer1_outputs(3552));
    layer2_outputs(3568) <= '1';
    layer2_outputs(3569) <= not(layer1_outputs(4602)) or (layer1_outputs(3040));
    layer2_outputs(3570) <= (layer1_outputs(2403)) and not (layer1_outputs(3685));
    layer2_outputs(3571) <= not(layer1_outputs(2355));
    layer2_outputs(3572) <= not((layer1_outputs(4381)) and (layer1_outputs(2335)));
    layer2_outputs(3573) <= layer1_outputs(3042);
    layer2_outputs(3574) <= (layer1_outputs(5483)) and (layer1_outputs(1411));
    layer2_outputs(3575) <= '0';
    layer2_outputs(3576) <= '1';
    layer2_outputs(3577) <= not((layer1_outputs(2374)) or (layer1_outputs(4275)));
    layer2_outputs(3578) <= '0';
    layer2_outputs(3579) <= not(layer1_outputs(5885)) or (layer1_outputs(6165));
    layer2_outputs(3580) <= '1';
    layer2_outputs(3581) <= not((layer1_outputs(1202)) or (layer1_outputs(2271)));
    layer2_outputs(3582) <= (layer1_outputs(3239)) and not (layer1_outputs(3721));
    layer2_outputs(3583) <= '0';
    layer2_outputs(3584) <= not(layer1_outputs(3841)) or (layer1_outputs(7630));
    layer2_outputs(3585) <= not(layer1_outputs(2604));
    layer2_outputs(3586) <= not(layer1_outputs(6695));
    layer2_outputs(3587) <= not((layer1_outputs(6487)) and (layer1_outputs(6152)));
    layer2_outputs(3588) <= not(layer1_outputs(658)) or (layer1_outputs(5439));
    layer2_outputs(3589) <= not(layer1_outputs(1734)) or (layer1_outputs(4870));
    layer2_outputs(3590) <= '0';
    layer2_outputs(3591) <= (layer1_outputs(267)) and not (layer1_outputs(5923));
    layer2_outputs(3592) <= (layer1_outputs(2216)) and not (layer1_outputs(6572));
    layer2_outputs(3593) <= (layer1_outputs(5376)) and not (layer1_outputs(5419));
    layer2_outputs(3594) <= not((layer1_outputs(2520)) or (layer1_outputs(3027)));
    layer2_outputs(3595) <= not(layer1_outputs(879)) or (layer1_outputs(6293));
    layer2_outputs(3596) <= (layer1_outputs(6308)) and (layer1_outputs(4599));
    layer2_outputs(3597) <= not(layer1_outputs(4750)) or (layer1_outputs(2525));
    layer2_outputs(3598) <= not(layer1_outputs(7211));
    layer2_outputs(3599) <= not(layer1_outputs(3632));
    layer2_outputs(3600) <= layer1_outputs(4582);
    layer2_outputs(3601) <= layer1_outputs(6888);
    layer2_outputs(3602) <= '0';
    layer2_outputs(3603) <= '1';
    layer2_outputs(3604) <= (layer1_outputs(3707)) or (layer1_outputs(4969));
    layer2_outputs(3605) <= '1';
    layer2_outputs(3606) <= (layer1_outputs(6537)) or (layer1_outputs(5815));
    layer2_outputs(3607) <= not(layer1_outputs(6756));
    layer2_outputs(3608) <= not(layer1_outputs(5672)) or (layer1_outputs(4467));
    layer2_outputs(3609) <= (layer1_outputs(3628)) xor (layer1_outputs(4438));
    layer2_outputs(3610) <= not((layer1_outputs(7499)) xor (layer1_outputs(4758)));
    layer2_outputs(3611) <= not(layer1_outputs(1643)) or (layer1_outputs(78));
    layer2_outputs(3612) <= '1';
    layer2_outputs(3613) <= (layer1_outputs(5234)) or (layer1_outputs(754));
    layer2_outputs(3614) <= layer1_outputs(4100);
    layer2_outputs(3615) <= (layer1_outputs(1500)) or (layer1_outputs(3416));
    layer2_outputs(3616) <= not((layer1_outputs(5998)) or (layer1_outputs(441)));
    layer2_outputs(3617) <= not((layer1_outputs(2843)) xor (layer1_outputs(5016)));
    layer2_outputs(3618) <= not(layer1_outputs(1874)) or (layer1_outputs(154));
    layer2_outputs(3619) <= (layer1_outputs(1811)) xor (layer1_outputs(5008));
    layer2_outputs(3620) <= not(layer1_outputs(1240)) or (layer1_outputs(1632));
    layer2_outputs(3621) <= layer1_outputs(7546);
    layer2_outputs(3622) <= (layer1_outputs(1080)) and not (layer1_outputs(5006));
    layer2_outputs(3623) <= (layer1_outputs(735)) and (layer1_outputs(6889));
    layer2_outputs(3624) <= not(layer1_outputs(3225)) or (layer1_outputs(4785));
    layer2_outputs(3625) <= not(layer1_outputs(7277)) or (layer1_outputs(7356));
    layer2_outputs(3626) <= not((layer1_outputs(2942)) xor (layer1_outputs(7098)));
    layer2_outputs(3627) <= not((layer1_outputs(5771)) and (layer1_outputs(6489)));
    layer2_outputs(3628) <= (layer1_outputs(1354)) and (layer1_outputs(1445));
    layer2_outputs(3629) <= (layer1_outputs(1821)) or (layer1_outputs(2373));
    layer2_outputs(3630) <= not(layer1_outputs(3859)) or (layer1_outputs(6253));
    layer2_outputs(3631) <= '1';
    layer2_outputs(3632) <= layer1_outputs(900);
    layer2_outputs(3633) <= '1';
    layer2_outputs(3634) <= not(layer1_outputs(85));
    layer2_outputs(3635) <= (layer1_outputs(7132)) and not (layer1_outputs(2447));
    layer2_outputs(3636) <= layer1_outputs(1197);
    layer2_outputs(3637) <= not((layer1_outputs(5740)) or (layer1_outputs(5030)));
    layer2_outputs(3638) <= layer1_outputs(5045);
    layer2_outputs(3639) <= not(layer1_outputs(4084));
    layer2_outputs(3640) <= (layer1_outputs(602)) and not (layer1_outputs(1239));
    layer2_outputs(3641) <= '1';
    layer2_outputs(3642) <= layer1_outputs(4280);
    layer2_outputs(3643) <= (layer1_outputs(2331)) and (layer1_outputs(2990));
    layer2_outputs(3644) <= not(layer1_outputs(4827));
    layer2_outputs(3645) <= not(layer1_outputs(6834));
    layer2_outputs(3646) <= not((layer1_outputs(2526)) and (layer1_outputs(4317)));
    layer2_outputs(3647) <= not(layer1_outputs(5420));
    layer2_outputs(3648) <= (layer1_outputs(7536)) and (layer1_outputs(7393));
    layer2_outputs(3649) <= layer1_outputs(6623);
    layer2_outputs(3650) <= not(layer1_outputs(4960)) or (layer1_outputs(5168));
    layer2_outputs(3651) <= '0';
    layer2_outputs(3652) <= not(layer1_outputs(4446)) or (layer1_outputs(4880));
    layer2_outputs(3653) <= (layer1_outputs(1388)) and not (layer1_outputs(6742));
    layer2_outputs(3654) <= (layer1_outputs(5746)) or (layer1_outputs(5752));
    layer2_outputs(3655) <= (layer1_outputs(2244)) and not (layer1_outputs(6576));
    layer2_outputs(3656) <= not(layer1_outputs(1966)) or (layer1_outputs(2925));
    layer2_outputs(3657) <= (layer1_outputs(1859)) and not (layer1_outputs(7588));
    layer2_outputs(3658) <= (layer1_outputs(5559)) and not (layer1_outputs(6734));
    layer2_outputs(3659) <= (layer1_outputs(5442)) and not (layer1_outputs(7368));
    layer2_outputs(3660) <= not(layer1_outputs(4975));
    layer2_outputs(3661) <= '0';
    layer2_outputs(3662) <= not(layer1_outputs(5316)) or (layer1_outputs(4372));
    layer2_outputs(3663) <= not(layer1_outputs(3559)) or (layer1_outputs(5415));
    layer2_outputs(3664) <= not(layer1_outputs(2803));
    layer2_outputs(3665) <= '1';
    layer2_outputs(3666) <= not(layer1_outputs(7024)) or (layer1_outputs(2797));
    layer2_outputs(3667) <= not((layer1_outputs(3299)) or (layer1_outputs(1506)));
    layer2_outputs(3668) <= (layer1_outputs(6541)) and (layer1_outputs(6820));
    layer2_outputs(3669) <= not((layer1_outputs(2157)) or (layer1_outputs(2305)));
    layer2_outputs(3670) <= (layer1_outputs(3493)) and (layer1_outputs(1144));
    layer2_outputs(3671) <= not((layer1_outputs(4856)) or (layer1_outputs(77)));
    layer2_outputs(3672) <= not((layer1_outputs(832)) and (layer1_outputs(33)));
    layer2_outputs(3673) <= not(layer1_outputs(1103));
    layer2_outputs(3674) <= layer1_outputs(7105);
    layer2_outputs(3675) <= not(layer1_outputs(5260));
    layer2_outputs(3676) <= not(layer1_outputs(6811));
    layer2_outputs(3677) <= (layer1_outputs(4256)) and not (layer1_outputs(5720));
    layer2_outputs(3678) <= not((layer1_outputs(5459)) or (layer1_outputs(2127)));
    layer2_outputs(3679) <= layer1_outputs(3791);
    layer2_outputs(3680) <= not(layer1_outputs(2139)) or (layer1_outputs(6214));
    layer2_outputs(3681) <= not(layer1_outputs(1266));
    layer2_outputs(3682) <= not(layer1_outputs(6375)) or (layer1_outputs(4008));
    layer2_outputs(3683) <= '1';
    layer2_outputs(3684) <= (layer1_outputs(3473)) and not (layer1_outputs(5188));
    layer2_outputs(3685) <= (layer1_outputs(7039)) and not (layer1_outputs(2491));
    layer2_outputs(3686) <= not(layer1_outputs(5958));
    layer2_outputs(3687) <= layer1_outputs(6341);
    layer2_outputs(3688) <= not(layer1_outputs(6088)) or (layer1_outputs(5300));
    layer2_outputs(3689) <= (layer1_outputs(7185)) and (layer1_outputs(7226));
    layer2_outputs(3690) <= not((layer1_outputs(1872)) or (layer1_outputs(898)));
    layer2_outputs(3691) <= not(layer1_outputs(1262)) or (layer1_outputs(2623));
    layer2_outputs(3692) <= (layer1_outputs(2736)) or (layer1_outputs(678));
    layer2_outputs(3693) <= (layer1_outputs(4644)) and not (layer1_outputs(757));
    layer2_outputs(3694) <= not((layer1_outputs(2023)) xor (layer1_outputs(6688)));
    layer2_outputs(3695) <= (layer1_outputs(4515)) and (layer1_outputs(3618));
    layer2_outputs(3696) <= (layer1_outputs(526)) or (layer1_outputs(1348));
    layer2_outputs(3697) <= not(layer1_outputs(7386));
    layer2_outputs(3698) <= layer1_outputs(1009);
    layer2_outputs(3699) <= '0';
    layer2_outputs(3700) <= '1';
    layer2_outputs(3701) <= '0';
    layer2_outputs(3702) <= not(layer1_outputs(4648));
    layer2_outputs(3703) <= not(layer1_outputs(345)) or (layer1_outputs(1143));
    layer2_outputs(3704) <= not((layer1_outputs(6795)) and (layer1_outputs(2340)));
    layer2_outputs(3705) <= not(layer1_outputs(3106));
    layer2_outputs(3706) <= (layer1_outputs(6611)) or (layer1_outputs(2619));
    layer2_outputs(3707) <= not(layer1_outputs(5554)) or (layer1_outputs(7319));
    layer2_outputs(3708) <= not(layer1_outputs(4142));
    layer2_outputs(3709) <= layer1_outputs(4767);
    layer2_outputs(3710) <= (layer1_outputs(2967)) and (layer1_outputs(4277));
    layer2_outputs(3711) <= layer1_outputs(7581);
    layer2_outputs(3712) <= not((layer1_outputs(2918)) and (layer1_outputs(6906)));
    layer2_outputs(3713) <= not(layer1_outputs(4747)) or (layer1_outputs(800));
    layer2_outputs(3714) <= not((layer1_outputs(7568)) or (layer1_outputs(4963)));
    layer2_outputs(3715) <= layer1_outputs(1571);
    layer2_outputs(3716) <= layer1_outputs(2101);
    layer2_outputs(3717) <= not((layer1_outputs(2621)) and (layer1_outputs(1539)));
    layer2_outputs(3718) <= not(layer1_outputs(4750));
    layer2_outputs(3719) <= '1';
    layer2_outputs(3720) <= not((layer1_outputs(2874)) or (layer1_outputs(4992)));
    layer2_outputs(3721) <= not(layer1_outputs(5198));
    layer2_outputs(3722) <= layer1_outputs(6015);
    layer2_outputs(3723) <= (layer1_outputs(7162)) or (layer1_outputs(2231));
    layer2_outputs(3724) <= (layer1_outputs(5890)) and (layer1_outputs(1064));
    layer2_outputs(3725) <= not(layer1_outputs(4396));
    layer2_outputs(3726) <= not((layer1_outputs(4153)) or (layer1_outputs(930)));
    layer2_outputs(3727) <= (layer1_outputs(7004)) and not (layer1_outputs(5804));
    layer2_outputs(3728) <= not(layer1_outputs(3687)) or (layer1_outputs(2776));
    layer2_outputs(3729) <= not(layer1_outputs(6253));
    layer2_outputs(3730) <= not(layer1_outputs(420)) or (layer1_outputs(794));
    layer2_outputs(3731) <= (layer1_outputs(2123)) and (layer1_outputs(6075));
    layer2_outputs(3732) <= (layer1_outputs(7546)) or (layer1_outputs(4005));
    layer2_outputs(3733) <= not(layer1_outputs(5218));
    layer2_outputs(3734) <= '1';
    layer2_outputs(3735) <= not((layer1_outputs(734)) and (layer1_outputs(3619)));
    layer2_outputs(3736) <= (layer1_outputs(6903)) or (layer1_outputs(2340));
    layer2_outputs(3737) <= '0';
    layer2_outputs(3738) <= not(layer1_outputs(4608)) or (layer1_outputs(2635));
    layer2_outputs(3739) <= not(layer1_outputs(2514)) or (layer1_outputs(6289));
    layer2_outputs(3740) <= not(layer1_outputs(263));
    layer2_outputs(3741) <= not(layer1_outputs(1816)) or (layer1_outputs(6096));
    layer2_outputs(3742) <= '1';
    layer2_outputs(3743) <= (layer1_outputs(3471)) or (layer1_outputs(4169));
    layer2_outputs(3744) <= (layer1_outputs(6245)) and not (layer1_outputs(502));
    layer2_outputs(3745) <= not((layer1_outputs(4359)) or (layer1_outputs(1732)));
    layer2_outputs(3746) <= not((layer1_outputs(993)) xor (layer1_outputs(1579)));
    layer2_outputs(3747) <= not(layer1_outputs(4981));
    layer2_outputs(3748) <= (layer1_outputs(4029)) and not (layer1_outputs(4150));
    layer2_outputs(3749) <= layer1_outputs(1379);
    layer2_outputs(3750) <= not(layer1_outputs(5593));
    layer2_outputs(3751) <= not(layer1_outputs(1511));
    layer2_outputs(3752) <= not((layer1_outputs(892)) and (layer1_outputs(5933)));
    layer2_outputs(3753) <= not(layer1_outputs(1376));
    layer2_outputs(3754) <= layer1_outputs(5083);
    layer2_outputs(3755) <= (layer1_outputs(4514)) and not (layer1_outputs(7532));
    layer2_outputs(3756) <= (layer1_outputs(7615)) and (layer1_outputs(4135));
    layer2_outputs(3757) <= (layer1_outputs(4615)) and not (layer1_outputs(1574));
    layer2_outputs(3758) <= not(layer1_outputs(243)) or (layer1_outputs(2655));
    layer2_outputs(3759) <= (layer1_outputs(1775)) and not (layer1_outputs(498));
    layer2_outputs(3760) <= layer1_outputs(6312);
    layer2_outputs(3761) <= (layer1_outputs(73)) and not (layer1_outputs(2026));
    layer2_outputs(3762) <= not(layer1_outputs(1458)) or (layer1_outputs(2163));
    layer2_outputs(3763) <= not(layer1_outputs(2203)) or (layer1_outputs(3911));
    layer2_outputs(3764) <= not(layer1_outputs(1434));
    layer2_outputs(3765) <= (layer1_outputs(4881)) and not (layer1_outputs(7362));
    layer2_outputs(3766) <= not(layer1_outputs(2942)) or (layer1_outputs(2877));
    layer2_outputs(3767) <= not(layer1_outputs(5497)) or (layer1_outputs(4518));
    layer2_outputs(3768) <= not(layer1_outputs(6744));
    layer2_outputs(3769) <= (layer1_outputs(5063)) and not (layer1_outputs(6701));
    layer2_outputs(3770) <= not(layer1_outputs(889)) or (layer1_outputs(3568));
    layer2_outputs(3771) <= not(layer1_outputs(5501)) or (layer1_outputs(6331));
    layer2_outputs(3772) <= (layer1_outputs(3023)) xor (layer1_outputs(5257));
    layer2_outputs(3773) <= (layer1_outputs(3374)) and not (layer1_outputs(5377));
    layer2_outputs(3774) <= not((layer1_outputs(19)) xor (layer1_outputs(431)));
    layer2_outputs(3775) <= (layer1_outputs(4688)) and (layer1_outputs(3146));
    layer2_outputs(3776) <= layer1_outputs(6409);
    layer2_outputs(3777) <= (layer1_outputs(2663)) and not (layer1_outputs(3058));
    layer2_outputs(3778) <= '1';
    layer2_outputs(3779) <= not((layer1_outputs(7047)) and (layer1_outputs(5487)));
    layer2_outputs(3780) <= (layer1_outputs(1103)) and not (layer1_outputs(4640));
    layer2_outputs(3781) <= not((layer1_outputs(2479)) or (layer1_outputs(2533)));
    layer2_outputs(3782) <= not(layer1_outputs(5688)) or (layer1_outputs(4746));
    layer2_outputs(3783) <= not(layer1_outputs(4365));
    layer2_outputs(3784) <= layer1_outputs(3811);
    layer2_outputs(3785) <= not((layer1_outputs(5781)) and (layer1_outputs(4322)));
    layer2_outputs(3786) <= not((layer1_outputs(2237)) or (layer1_outputs(637)));
    layer2_outputs(3787) <= '1';
    layer2_outputs(3788) <= (layer1_outputs(5274)) or (layer1_outputs(1786));
    layer2_outputs(3789) <= not((layer1_outputs(5283)) and (layer1_outputs(7239)));
    layer2_outputs(3790) <= not(layer1_outputs(3371));
    layer2_outputs(3791) <= (layer1_outputs(5437)) and not (layer1_outputs(5931));
    layer2_outputs(3792) <= not((layer1_outputs(6213)) or (layer1_outputs(162)));
    layer2_outputs(3793) <= (layer1_outputs(2704)) and (layer1_outputs(5790));
    layer2_outputs(3794) <= not(layer1_outputs(3517));
    layer2_outputs(3795) <= '0';
    layer2_outputs(3796) <= (layer1_outputs(618)) and not (layer1_outputs(7035));
    layer2_outputs(3797) <= layer1_outputs(2979);
    layer2_outputs(3798) <= not((layer1_outputs(4045)) and (layer1_outputs(536)));
    layer2_outputs(3799) <= (layer1_outputs(5431)) or (layer1_outputs(3458));
    layer2_outputs(3800) <= not(layer1_outputs(4053)) or (layer1_outputs(523));
    layer2_outputs(3801) <= (layer1_outputs(2958)) and not (layer1_outputs(2590));
    layer2_outputs(3802) <= not(layer1_outputs(3852)) or (layer1_outputs(7180));
    layer2_outputs(3803) <= not(layer1_outputs(580)) or (layer1_outputs(3003));
    layer2_outputs(3804) <= not((layer1_outputs(4213)) or (layer1_outputs(2585)));
    layer2_outputs(3805) <= layer1_outputs(4313);
    layer2_outputs(3806) <= not(layer1_outputs(7139));
    layer2_outputs(3807) <= '1';
    layer2_outputs(3808) <= (layer1_outputs(5031)) and (layer1_outputs(6780));
    layer2_outputs(3809) <= not(layer1_outputs(5896)) or (layer1_outputs(1697));
    layer2_outputs(3810) <= not(layer1_outputs(5033)) or (layer1_outputs(3589));
    layer2_outputs(3811) <= not(layer1_outputs(5653)) or (layer1_outputs(6751));
    layer2_outputs(3812) <= (layer1_outputs(4210)) and not (layer1_outputs(4816));
    layer2_outputs(3813) <= (layer1_outputs(591)) or (layer1_outputs(2584));
    layer2_outputs(3814) <= '1';
    layer2_outputs(3815) <= layer1_outputs(4517);
    layer2_outputs(3816) <= not(layer1_outputs(4330));
    layer2_outputs(3817) <= not(layer1_outputs(6867));
    layer2_outputs(3818) <= not((layer1_outputs(6538)) and (layer1_outputs(3863)));
    layer2_outputs(3819) <= layer1_outputs(4466);
    layer2_outputs(3820) <= '1';
    layer2_outputs(3821) <= not(layer1_outputs(7033)) or (layer1_outputs(4682));
    layer2_outputs(3822) <= not(layer1_outputs(1055));
    layer2_outputs(3823) <= not((layer1_outputs(5845)) and (layer1_outputs(699)));
    layer2_outputs(3824) <= layer1_outputs(5360);
    layer2_outputs(3825) <= (layer1_outputs(7095)) and not (layer1_outputs(4723));
    layer2_outputs(3826) <= not((layer1_outputs(5567)) and (layer1_outputs(6350)));
    layer2_outputs(3827) <= not((layer1_outputs(1251)) or (layer1_outputs(287)));
    layer2_outputs(3828) <= not(layer1_outputs(1035)) or (layer1_outputs(3001));
    layer2_outputs(3829) <= '1';
    layer2_outputs(3830) <= not(layer1_outputs(2996)) or (layer1_outputs(417));
    layer2_outputs(3831) <= not(layer1_outputs(283)) or (layer1_outputs(1367));
    layer2_outputs(3832) <= not(layer1_outputs(1441));
    layer2_outputs(3833) <= not(layer1_outputs(4660)) or (layer1_outputs(1271));
    layer2_outputs(3834) <= '1';
    layer2_outputs(3835) <= (layer1_outputs(2174)) xor (layer1_outputs(4752));
    layer2_outputs(3836) <= (layer1_outputs(1278)) and (layer1_outputs(1882));
    layer2_outputs(3837) <= layer1_outputs(1133);
    layer2_outputs(3838) <= '1';
    layer2_outputs(3839) <= not(layer1_outputs(5447));
    layer2_outputs(3840) <= not((layer1_outputs(6964)) or (layer1_outputs(2735)));
    layer2_outputs(3841) <= not(layer1_outputs(889)) or (layer1_outputs(3906));
    layer2_outputs(3842) <= (layer1_outputs(496)) or (layer1_outputs(4790));
    layer2_outputs(3843) <= not(layer1_outputs(4612));
    layer2_outputs(3844) <= layer1_outputs(5003);
    layer2_outputs(3845) <= (layer1_outputs(5835)) and not (layer1_outputs(6915));
    layer2_outputs(3846) <= layer1_outputs(5630);
    layer2_outputs(3847) <= '1';
    layer2_outputs(3848) <= (layer1_outputs(5624)) and not (layer1_outputs(6226));
    layer2_outputs(3849) <= not(layer1_outputs(1394));
    layer2_outputs(3850) <= (layer1_outputs(938)) or (layer1_outputs(5323));
    layer2_outputs(3851) <= not((layer1_outputs(7396)) xor (layer1_outputs(394)));
    layer2_outputs(3852) <= layer1_outputs(5934);
    layer2_outputs(3853) <= '1';
    layer2_outputs(3854) <= not(layer1_outputs(2429));
    layer2_outputs(3855) <= (layer1_outputs(5443)) and not (layer1_outputs(1720));
    layer2_outputs(3856) <= (layer1_outputs(1612)) or (layer1_outputs(3104));
    layer2_outputs(3857) <= (layer1_outputs(5984)) and (layer1_outputs(1504));
    layer2_outputs(3858) <= not(layer1_outputs(2564));
    layer2_outputs(3859) <= '1';
    layer2_outputs(3860) <= layer1_outputs(698);
    layer2_outputs(3861) <= '0';
    layer2_outputs(3862) <= (layer1_outputs(2553)) and (layer1_outputs(4921));
    layer2_outputs(3863) <= not((layer1_outputs(383)) and (layer1_outputs(5488)));
    layer2_outputs(3864) <= '1';
    layer2_outputs(3865) <= '0';
    layer2_outputs(3866) <= not(layer1_outputs(1131)) or (layer1_outputs(7283));
    layer2_outputs(3867) <= (layer1_outputs(2874)) or (layer1_outputs(352));
    layer2_outputs(3868) <= not(layer1_outputs(1806));
    layer2_outputs(3869) <= (layer1_outputs(689)) and (layer1_outputs(1787));
    layer2_outputs(3870) <= layer1_outputs(6573);
    layer2_outputs(3871) <= not(layer1_outputs(6323));
    layer2_outputs(3872) <= not((layer1_outputs(7152)) and (layer1_outputs(6674)));
    layer2_outputs(3873) <= (layer1_outputs(6070)) and not (layer1_outputs(4130));
    layer2_outputs(3874) <= not((layer1_outputs(5327)) xor (layer1_outputs(7668)));
    layer2_outputs(3875) <= not((layer1_outputs(4208)) and (layer1_outputs(1911)));
    layer2_outputs(3876) <= not(layer1_outputs(7365)) or (layer1_outputs(2276));
    layer2_outputs(3877) <= not(layer1_outputs(7033));
    layer2_outputs(3878) <= layer1_outputs(4569);
    layer2_outputs(3879) <= not(layer1_outputs(7060)) or (layer1_outputs(4962));
    layer2_outputs(3880) <= '1';
    layer2_outputs(3881) <= (layer1_outputs(6221)) and not (layer1_outputs(5085));
    layer2_outputs(3882) <= not(layer1_outputs(4868));
    layer2_outputs(3883) <= (layer1_outputs(7144)) or (layer1_outputs(5623));
    layer2_outputs(3884) <= not(layer1_outputs(5098));
    layer2_outputs(3885) <= (layer1_outputs(798)) and not (layer1_outputs(3795));
    layer2_outputs(3886) <= not(layer1_outputs(4990)) or (layer1_outputs(3547));
    layer2_outputs(3887) <= '0';
    layer2_outputs(3888) <= not((layer1_outputs(4462)) and (layer1_outputs(2408)));
    layer2_outputs(3889) <= (layer1_outputs(7323)) or (layer1_outputs(5176));
    layer2_outputs(3890) <= '1';
    layer2_outputs(3891) <= (layer1_outputs(2847)) and not (layer1_outputs(3103));
    layer2_outputs(3892) <= not(layer1_outputs(6923)) or (layer1_outputs(7491));
    layer2_outputs(3893) <= not(layer1_outputs(7593)) or (layer1_outputs(2361));
    layer2_outputs(3894) <= (layer1_outputs(1722)) and (layer1_outputs(1274));
    layer2_outputs(3895) <= '1';
    layer2_outputs(3896) <= '1';
    layer2_outputs(3897) <= not(layer1_outputs(6604));
    layer2_outputs(3898) <= (layer1_outputs(2561)) and not (layer1_outputs(2598));
    layer2_outputs(3899) <= '0';
    layer2_outputs(3900) <= '0';
    layer2_outputs(3901) <= not(layer1_outputs(1926)) or (layer1_outputs(2267));
    layer2_outputs(3902) <= '0';
    layer2_outputs(3903) <= not((layer1_outputs(3260)) or (layer1_outputs(613)));
    layer2_outputs(3904) <= not(layer1_outputs(1));
    layer2_outputs(3905) <= layer1_outputs(4215);
    layer2_outputs(3906) <= not(layer1_outputs(3580));
    layer2_outputs(3907) <= '0';
    layer2_outputs(3908) <= not((layer1_outputs(722)) or (layer1_outputs(530)));
    layer2_outputs(3909) <= '0';
    layer2_outputs(3910) <= (layer1_outputs(4937)) and (layer1_outputs(6494));
    layer2_outputs(3911) <= not(layer1_outputs(3463)) or (layer1_outputs(1061));
    layer2_outputs(3912) <= not(layer1_outputs(2152));
    layer2_outputs(3913) <= '0';
    layer2_outputs(3914) <= layer1_outputs(3926);
    layer2_outputs(3915) <= not(layer1_outputs(1792));
    layer2_outputs(3916) <= not((layer1_outputs(6804)) and (layer1_outputs(5783)));
    layer2_outputs(3917) <= not(layer1_outputs(1738));
    layer2_outputs(3918) <= '0';
    layer2_outputs(3919) <= '0';
    layer2_outputs(3920) <= (layer1_outputs(3753)) or (layer1_outputs(5589));
    layer2_outputs(3921) <= '0';
    layer2_outputs(3922) <= not(layer1_outputs(4391)) or (layer1_outputs(1480));
    layer2_outputs(3923) <= not(layer1_outputs(7509));
    layer2_outputs(3924) <= not((layer1_outputs(651)) or (layer1_outputs(6799)));
    layer2_outputs(3925) <= not((layer1_outputs(4787)) or (layer1_outputs(1260)));
    layer2_outputs(3926) <= '0';
    layer2_outputs(3927) <= not((layer1_outputs(3229)) or (layer1_outputs(5608)));
    layer2_outputs(3928) <= not((layer1_outputs(645)) or (layer1_outputs(1498)));
    layer2_outputs(3929) <= '0';
    layer2_outputs(3930) <= (layer1_outputs(4291)) and (layer1_outputs(5120));
    layer2_outputs(3931) <= (layer1_outputs(224)) and not (layer1_outputs(2147));
    layer2_outputs(3932) <= (layer1_outputs(6233)) and not (layer1_outputs(6053));
    layer2_outputs(3933) <= not((layer1_outputs(1852)) or (layer1_outputs(6345)));
    layer2_outputs(3934) <= (layer1_outputs(5755)) and not (layer1_outputs(5213));
    layer2_outputs(3935) <= (layer1_outputs(6180)) or (layer1_outputs(161));
    layer2_outputs(3936) <= not(layer1_outputs(5974));
    layer2_outputs(3937) <= layer1_outputs(3228);
    layer2_outputs(3938) <= (layer1_outputs(3228)) and (layer1_outputs(6493));
    layer2_outputs(3939) <= not((layer1_outputs(6671)) and (layer1_outputs(5704)));
    layer2_outputs(3940) <= not(layer1_outputs(275));
    layer2_outputs(3941) <= (layer1_outputs(5982)) and not (layer1_outputs(2985));
    layer2_outputs(3942) <= not(layer1_outputs(7637));
    layer2_outputs(3943) <= (layer1_outputs(3846)) or (layer1_outputs(6492));
    layer2_outputs(3944) <= (layer1_outputs(6965)) or (layer1_outputs(629));
    layer2_outputs(3945) <= not(layer1_outputs(6685));
    layer2_outputs(3946) <= (layer1_outputs(100)) or (layer1_outputs(2618));
    layer2_outputs(3947) <= '1';
    layer2_outputs(3948) <= (layer1_outputs(3016)) and not (layer1_outputs(3065));
    layer2_outputs(3949) <= not(layer1_outputs(6957));
    layer2_outputs(3950) <= not((layer1_outputs(2879)) and (layer1_outputs(813)));
    layer2_outputs(3951) <= '0';
    layer2_outputs(3952) <= '1';
    layer2_outputs(3953) <= not(layer1_outputs(3607));
    layer2_outputs(3954) <= (layer1_outputs(6523)) and (layer1_outputs(5));
    layer2_outputs(3955) <= layer1_outputs(1046);
    layer2_outputs(3956) <= not((layer1_outputs(3239)) and (layer1_outputs(3188)));
    layer2_outputs(3957) <= not(layer1_outputs(1773)) or (layer1_outputs(4114));
    layer2_outputs(3958) <= (layer1_outputs(1313)) and not (layer1_outputs(4112));
    layer2_outputs(3959) <= (layer1_outputs(368)) and (layer1_outputs(2022));
    layer2_outputs(3960) <= '0';
    layer2_outputs(3961) <= '0';
    layer2_outputs(3962) <= '1';
    layer2_outputs(3963) <= '1';
    layer2_outputs(3964) <= not((layer1_outputs(1113)) or (layer1_outputs(274)));
    layer2_outputs(3965) <= not((layer1_outputs(6303)) or (layer1_outputs(2897)));
    layer2_outputs(3966) <= not(layer1_outputs(5405));
    layer2_outputs(3967) <= (layer1_outputs(3591)) and not (layer1_outputs(3430));
    layer2_outputs(3968) <= (layer1_outputs(3221)) and (layer1_outputs(2195));
    layer2_outputs(3969) <= (layer1_outputs(4421)) and not (layer1_outputs(4541));
    layer2_outputs(3970) <= (layer1_outputs(2708)) and not (layer1_outputs(7456));
    layer2_outputs(3971) <= not(layer1_outputs(5557)) or (layer1_outputs(5136));
    layer2_outputs(3972) <= not((layer1_outputs(2125)) or (layer1_outputs(601)));
    layer2_outputs(3973) <= not(layer1_outputs(4471));
    layer2_outputs(3974) <= not(layer1_outputs(2881)) or (layer1_outputs(3985));
    layer2_outputs(3975) <= (layer1_outputs(600)) or (layer1_outputs(4788));
    layer2_outputs(3976) <= not(layer1_outputs(5788));
    layer2_outputs(3977) <= '1';
    layer2_outputs(3978) <= not(layer1_outputs(262));
    layer2_outputs(3979) <= '0';
    layer2_outputs(3980) <= not(layer1_outputs(21));
    layer2_outputs(3981) <= not(layer1_outputs(3728));
    layer2_outputs(3982) <= not((layer1_outputs(331)) and (layer1_outputs(5732)));
    layer2_outputs(3983) <= (layer1_outputs(5023)) and not (layer1_outputs(5660));
    layer2_outputs(3984) <= (layer1_outputs(6613)) and not (layer1_outputs(5400));
    layer2_outputs(3985) <= not(layer1_outputs(2489)) or (layer1_outputs(278));
    layer2_outputs(3986) <= not(layer1_outputs(238)) or (layer1_outputs(4841));
    layer2_outputs(3987) <= not((layer1_outputs(4296)) and (layer1_outputs(1619)));
    layer2_outputs(3988) <= not(layer1_outputs(4201)) or (layer1_outputs(6466));
    layer2_outputs(3989) <= (layer1_outputs(5286)) and (layer1_outputs(1551));
    layer2_outputs(3990) <= (layer1_outputs(5066)) and (layer1_outputs(1770));
    layer2_outputs(3991) <= '0';
    layer2_outputs(3992) <= layer1_outputs(6278);
    layer2_outputs(3993) <= not((layer1_outputs(4570)) or (layer1_outputs(2291)));
    layer2_outputs(3994) <= (layer1_outputs(4978)) and not (layer1_outputs(7626));
    layer2_outputs(3995) <= not(layer1_outputs(840));
    layer2_outputs(3996) <= not(layer1_outputs(91));
    layer2_outputs(3997) <= not(layer1_outputs(506)) or (layer1_outputs(1811));
    layer2_outputs(3998) <= not(layer1_outputs(4065)) or (layer1_outputs(6123));
    layer2_outputs(3999) <= layer1_outputs(4794);
    layer2_outputs(4000) <= (layer1_outputs(5545)) and not (layer1_outputs(1621));
    layer2_outputs(4001) <= '0';
    layer2_outputs(4002) <= (layer1_outputs(4217)) and not (layer1_outputs(5435));
    layer2_outputs(4003) <= (layer1_outputs(23)) and not (layer1_outputs(3355));
    layer2_outputs(4004) <= layer1_outputs(2908);
    layer2_outputs(4005) <= not((layer1_outputs(4453)) xor (layer1_outputs(6917)));
    layer2_outputs(4006) <= (layer1_outputs(6933)) and (layer1_outputs(3695));
    layer2_outputs(4007) <= not(layer1_outputs(5005));
    layer2_outputs(4008) <= not((layer1_outputs(4919)) or (layer1_outputs(4288)));
    layer2_outputs(4009) <= not(layer1_outputs(5159));
    layer2_outputs(4010) <= layer1_outputs(4738);
    layer2_outputs(4011) <= (layer1_outputs(5163)) or (layer1_outputs(6681));
    layer2_outputs(4012) <= (layer1_outputs(3897)) or (layer1_outputs(2861));
    layer2_outputs(4013) <= layer1_outputs(5498);
    layer2_outputs(4014) <= not(layer1_outputs(259));
    layer2_outputs(4015) <= not((layer1_outputs(285)) xor (layer1_outputs(5812)));
    layer2_outputs(4016) <= (layer1_outputs(645)) or (layer1_outputs(3256));
    layer2_outputs(4017) <= layer1_outputs(5857);
    layer2_outputs(4018) <= not(layer1_outputs(4371));
    layer2_outputs(4019) <= not(layer1_outputs(5496));
    layer2_outputs(4020) <= (layer1_outputs(3234)) xor (layer1_outputs(2354));
    layer2_outputs(4021) <= not((layer1_outputs(3561)) and (layer1_outputs(37)));
    layer2_outputs(4022) <= (layer1_outputs(7429)) and not (layer1_outputs(6043));
    layer2_outputs(4023) <= not(layer1_outputs(2402)) or (layer1_outputs(319));
    layer2_outputs(4024) <= not(layer1_outputs(457));
    layer2_outputs(4025) <= '1';
    layer2_outputs(4026) <= (layer1_outputs(5700)) and not (layer1_outputs(3839));
    layer2_outputs(4027) <= (layer1_outputs(1052)) or (layer1_outputs(2204));
    layer2_outputs(4028) <= (layer1_outputs(6744)) xor (layer1_outputs(1146));
    layer2_outputs(4029) <= not((layer1_outputs(1498)) or (layer1_outputs(6766)));
    layer2_outputs(4030) <= not((layer1_outputs(4058)) and (layer1_outputs(3338)));
    layer2_outputs(4031) <= not(layer1_outputs(7203));
    layer2_outputs(4032) <= (layer1_outputs(6276)) and not (layer1_outputs(1234));
    layer2_outputs(4033) <= (layer1_outputs(674)) or (layer1_outputs(1984));
    layer2_outputs(4034) <= not(layer1_outputs(5478)) or (layer1_outputs(6701));
    layer2_outputs(4035) <= '1';
    layer2_outputs(4036) <= '1';
    layer2_outputs(4037) <= layer1_outputs(7107);
    layer2_outputs(4038) <= (layer1_outputs(4954)) or (layer1_outputs(4988));
    layer2_outputs(4039) <= not((layer1_outputs(4118)) or (layer1_outputs(6312)));
    layer2_outputs(4040) <= not(layer1_outputs(3410)) or (layer1_outputs(1118));
    layer2_outputs(4041) <= not(layer1_outputs(3513)) or (layer1_outputs(1048));
    layer2_outputs(4042) <= (layer1_outputs(3939)) and not (layer1_outputs(6640));
    layer2_outputs(4043) <= (layer1_outputs(2013)) or (layer1_outputs(561));
    layer2_outputs(4044) <= '0';
    layer2_outputs(4045) <= (layer1_outputs(6638)) xor (layer1_outputs(4666));
    layer2_outputs(4046) <= not(layer1_outputs(1293)) or (layer1_outputs(1405));
    layer2_outputs(4047) <= not(layer1_outputs(315));
    layer2_outputs(4048) <= (layer1_outputs(643)) and (layer1_outputs(6992));
    layer2_outputs(4049) <= (layer1_outputs(1272)) or (layer1_outputs(4939));
    layer2_outputs(4050) <= not(layer1_outputs(4437));
    layer2_outputs(4051) <= (layer1_outputs(3711)) and (layer1_outputs(6234));
    layer2_outputs(4052) <= not(layer1_outputs(1858)) or (layer1_outputs(4884));
    layer2_outputs(4053) <= not((layer1_outputs(6543)) or (layer1_outputs(1481)));
    layer2_outputs(4054) <= not(layer1_outputs(6946));
    layer2_outputs(4055) <= not(layer1_outputs(6965));
    layer2_outputs(4056) <= '1';
    layer2_outputs(4057) <= (layer1_outputs(2314)) and not (layer1_outputs(2199));
    layer2_outputs(4058) <= '1';
    layer2_outputs(4059) <= (layer1_outputs(1022)) and not (layer1_outputs(5450));
    layer2_outputs(4060) <= not((layer1_outputs(2947)) or (layer1_outputs(2237)));
    layer2_outputs(4061) <= not(layer1_outputs(6389));
    layer2_outputs(4062) <= layer1_outputs(4299);
    layer2_outputs(4063) <= (layer1_outputs(3025)) and not (layer1_outputs(2962));
    layer2_outputs(4064) <= layer1_outputs(6132);
    layer2_outputs(4065) <= layer1_outputs(2420);
    layer2_outputs(4066) <= not(layer1_outputs(6875)) or (layer1_outputs(2669));
    layer2_outputs(4067) <= (layer1_outputs(6981)) or (layer1_outputs(5911));
    layer2_outputs(4068) <= not(layer1_outputs(1965)) or (layer1_outputs(483));
    layer2_outputs(4069) <= (layer1_outputs(6403)) or (layer1_outputs(2992));
    layer2_outputs(4070) <= '1';
    layer2_outputs(4071) <= (layer1_outputs(4043)) and not (layer1_outputs(970));
    layer2_outputs(4072) <= not((layer1_outputs(5177)) and (layer1_outputs(5826)));
    layer2_outputs(4073) <= not(layer1_outputs(1902));
    layer2_outputs(4074) <= not((layer1_outputs(6242)) or (layer1_outputs(324)));
    layer2_outputs(4075) <= '0';
    layer2_outputs(4076) <= not(layer1_outputs(4793));
    layer2_outputs(4077) <= (layer1_outputs(3980)) and not (layer1_outputs(1258));
    layer2_outputs(4078) <= not(layer1_outputs(4977));
    layer2_outputs(4079) <= not((layer1_outputs(4083)) and (layer1_outputs(1055)));
    layer2_outputs(4080) <= (layer1_outputs(5864)) and (layer1_outputs(15));
    layer2_outputs(4081) <= layer1_outputs(763);
    layer2_outputs(4082) <= not((layer1_outputs(3864)) and (layer1_outputs(3445)));
    layer2_outputs(4083) <= not(layer1_outputs(5910));
    layer2_outputs(4084) <= layer1_outputs(7424);
    layer2_outputs(4085) <= not((layer1_outputs(3392)) and (layer1_outputs(379)));
    layer2_outputs(4086) <= not((layer1_outputs(5042)) xor (layer1_outputs(90)));
    layer2_outputs(4087) <= '0';
    layer2_outputs(4088) <= not(layer1_outputs(2342)) or (layer1_outputs(2982));
    layer2_outputs(4089) <= (layer1_outputs(3216)) and not (layer1_outputs(453));
    layer2_outputs(4090) <= (layer1_outputs(623)) and (layer1_outputs(3910));
    layer2_outputs(4091) <= not((layer1_outputs(133)) or (layer1_outputs(6454)));
    layer2_outputs(4092) <= not((layer1_outputs(5291)) and (layer1_outputs(6651)));
    layer2_outputs(4093) <= (layer1_outputs(1263)) xor (layer1_outputs(148));
    layer2_outputs(4094) <= '0';
    layer2_outputs(4095) <= not(layer1_outputs(5286));
    layer2_outputs(4096) <= not((layer1_outputs(4399)) or (layer1_outputs(7232)));
    layer2_outputs(4097) <= not(layer1_outputs(4505));
    layer2_outputs(4098) <= (layer1_outputs(6011)) and not (layer1_outputs(6484));
    layer2_outputs(4099) <= layer1_outputs(5124);
    layer2_outputs(4100) <= not(layer1_outputs(1363));
    layer2_outputs(4101) <= not(layer1_outputs(4249));
    layer2_outputs(4102) <= not(layer1_outputs(4491)) or (layer1_outputs(1860));
    layer2_outputs(4103) <= (layer1_outputs(2262)) and not (layer1_outputs(4561));
    layer2_outputs(4104) <= (layer1_outputs(3892)) and not (layer1_outputs(4907));
    layer2_outputs(4105) <= not(layer1_outputs(4645));
    layer2_outputs(4106) <= '0';
    layer2_outputs(4107) <= (layer1_outputs(5206)) xor (layer1_outputs(5441));
    layer2_outputs(4108) <= not(layer1_outputs(1513)) or (layer1_outputs(6684));
    layer2_outputs(4109) <= not((layer1_outputs(4414)) or (layer1_outputs(5435)));
    layer2_outputs(4110) <= (layer1_outputs(3533)) and (layer1_outputs(1282));
    layer2_outputs(4111) <= layer1_outputs(675);
    layer2_outputs(4112) <= '0';
    layer2_outputs(4113) <= layer1_outputs(1687);
    layer2_outputs(4114) <= not(layer1_outputs(7188));
    layer2_outputs(4115) <= not((layer1_outputs(2638)) and (layer1_outputs(3991)));
    layer2_outputs(4116) <= '1';
    layer2_outputs(4117) <= layer1_outputs(3708);
    layer2_outputs(4118) <= not(layer1_outputs(1896));
    layer2_outputs(4119) <= '1';
    layer2_outputs(4120) <= not((layer1_outputs(3508)) and (layer1_outputs(2802)));
    layer2_outputs(4121) <= (layer1_outputs(804)) and not (layer1_outputs(2362));
    layer2_outputs(4122) <= not(layer1_outputs(3934));
    layer2_outputs(4123) <= not((layer1_outputs(7312)) and (layer1_outputs(2832)));
    layer2_outputs(4124) <= not(layer1_outputs(7372));
    layer2_outputs(4125) <= (layer1_outputs(400)) or (layer1_outputs(5146));
    layer2_outputs(4126) <= layer1_outputs(2970);
    layer2_outputs(4127) <= '0';
    layer2_outputs(4128) <= (layer1_outputs(1060)) and not (layer1_outputs(3007));
    layer2_outputs(4129) <= '1';
    layer2_outputs(4130) <= (layer1_outputs(6882)) or (layer1_outputs(1633));
    layer2_outputs(4131) <= not(layer1_outputs(1912));
    layer2_outputs(4132) <= (layer1_outputs(7134)) and not (layer1_outputs(3894));
    layer2_outputs(4133) <= not(layer1_outputs(5741));
    layer2_outputs(4134) <= '1';
    layer2_outputs(4135) <= layer1_outputs(1415);
    layer2_outputs(4136) <= not(layer1_outputs(4152));
    layer2_outputs(4137) <= (layer1_outputs(879)) and not (layer1_outputs(854));
    layer2_outputs(4138) <= not(layer1_outputs(4955));
    layer2_outputs(4139) <= (layer1_outputs(3013)) and (layer1_outputs(3528));
    layer2_outputs(4140) <= (layer1_outputs(4755)) and (layer1_outputs(2192));
    layer2_outputs(4141) <= not(layer1_outputs(2364)) or (layer1_outputs(7064));
    layer2_outputs(4142) <= (layer1_outputs(2023)) and not (layer1_outputs(3049));
    layer2_outputs(4143) <= not(layer1_outputs(4589)) or (layer1_outputs(4149));
    layer2_outputs(4144) <= not(layer1_outputs(5955));
    layer2_outputs(4145) <= (layer1_outputs(691)) and not (layer1_outputs(1488));
    layer2_outputs(4146) <= not(layer1_outputs(582)) or (layer1_outputs(6507));
    layer2_outputs(4147) <= not((layer1_outputs(1821)) or (layer1_outputs(2615)));
    layer2_outputs(4148) <= '1';
    layer2_outputs(4149) <= not((layer1_outputs(7583)) and (layer1_outputs(975)));
    layer2_outputs(4150) <= '1';
    layer2_outputs(4151) <= layer1_outputs(4035);
    layer2_outputs(4152) <= (layer1_outputs(2889)) and not (layer1_outputs(932));
    layer2_outputs(4153) <= layer1_outputs(5865);
    layer2_outputs(4154) <= (layer1_outputs(5372)) and (layer1_outputs(5843));
    layer2_outputs(4155) <= (layer1_outputs(1609)) and not (layer1_outputs(2107));
    layer2_outputs(4156) <= not(layer1_outputs(841));
    layer2_outputs(4157) <= layer1_outputs(955);
    layer2_outputs(4158) <= (layer1_outputs(5241)) and (layer1_outputs(7518));
    layer2_outputs(4159) <= layer1_outputs(3298);
    layer2_outputs(4160) <= layer1_outputs(1510);
    layer2_outputs(4161) <= (layer1_outputs(3307)) or (layer1_outputs(2105));
    layer2_outputs(4162) <= not(layer1_outputs(6847)) or (layer1_outputs(149));
    layer2_outputs(4163) <= layer1_outputs(3311);
    layer2_outputs(4164) <= not((layer1_outputs(1291)) or (layer1_outputs(6251)));
    layer2_outputs(4165) <= (layer1_outputs(6003)) or (layer1_outputs(1947));
    layer2_outputs(4166) <= layer1_outputs(1558);
    layer2_outputs(4167) <= layer1_outputs(4124);
    layer2_outputs(4168) <= layer1_outputs(7067);
    layer2_outputs(4169) <= not((layer1_outputs(2198)) xor (layer1_outputs(5491)));
    layer2_outputs(4170) <= layer1_outputs(50);
    layer2_outputs(4171) <= not((layer1_outputs(1158)) and (layer1_outputs(1058)));
    layer2_outputs(4172) <= (layer1_outputs(2203)) and not (layer1_outputs(3669));
    layer2_outputs(4173) <= layer1_outputs(3290);
    layer2_outputs(4174) <= layer1_outputs(5980);
    layer2_outputs(4175) <= '0';
    layer2_outputs(4176) <= not(layer1_outputs(3593)) or (layer1_outputs(2268));
    layer2_outputs(4177) <= not(layer1_outputs(3706));
    layer2_outputs(4178) <= layer1_outputs(265);
    layer2_outputs(4179) <= layer1_outputs(7295);
    layer2_outputs(4180) <= (layer1_outputs(752)) or (layer1_outputs(4658));
    layer2_outputs(4181) <= (layer1_outputs(2359)) and (layer1_outputs(5301));
    layer2_outputs(4182) <= '0';
    layer2_outputs(4183) <= not((layer1_outputs(720)) and (layer1_outputs(1570)));
    layer2_outputs(4184) <= '1';
    layer2_outputs(4185) <= not(layer1_outputs(4415));
    layer2_outputs(4186) <= not(layer1_outputs(4951)) or (layer1_outputs(1294));
    layer2_outputs(4187) <= layer1_outputs(7387);
    layer2_outputs(4188) <= '0';
    layer2_outputs(4189) <= layer1_outputs(4589);
    layer2_outputs(4190) <= not(layer1_outputs(137)) or (layer1_outputs(2169));
    layer2_outputs(4191) <= '0';
    layer2_outputs(4192) <= (layer1_outputs(7544)) and not (layer1_outputs(856));
    layer2_outputs(4193) <= (layer1_outputs(2545)) and not (layer1_outputs(6879));
    layer2_outputs(4194) <= not((layer1_outputs(1721)) or (layer1_outputs(7476)));
    layer2_outputs(4195) <= '0';
    layer2_outputs(4196) <= not((layer1_outputs(451)) and (layer1_outputs(4520)));
    layer2_outputs(4197) <= layer1_outputs(3739);
    layer2_outputs(4198) <= not(layer1_outputs(4527)) or (layer1_outputs(1314));
    layer2_outputs(4199) <= '0';
    layer2_outputs(4200) <= (layer1_outputs(2610)) or (layer1_outputs(6037));
    layer2_outputs(4201) <= layer1_outputs(7636);
    layer2_outputs(4202) <= layer1_outputs(5668);
    layer2_outputs(4203) <= '0';
    layer2_outputs(4204) <= (layer1_outputs(44)) and not (layer1_outputs(3172));
    layer2_outputs(4205) <= not((layer1_outputs(5397)) and (layer1_outputs(1409)));
    layer2_outputs(4206) <= '1';
    layer2_outputs(4207) <= not(layer1_outputs(2424));
    layer2_outputs(4208) <= not(layer1_outputs(577)) or (layer1_outputs(7203));
    layer2_outputs(4209) <= not(layer1_outputs(7440));
    layer2_outputs(4210) <= not(layer1_outputs(5878)) or (layer1_outputs(2002));
    layer2_outputs(4211) <= not(layer1_outputs(4325)) or (layer1_outputs(5258));
    layer2_outputs(4212) <= layer1_outputs(3633);
    layer2_outputs(4213) <= not(layer1_outputs(1426));
    layer2_outputs(4214) <= '0';
    layer2_outputs(4215) <= not(layer1_outputs(577)) or (layer1_outputs(2749));
    layer2_outputs(4216) <= '1';
    layer2_outputs(4217) <= '0';
    layer2_outputs(4218) <= layer1_outputs(954);
    layer2_outputs(4219) <= (layer1_outputs(3405)) and (layer1_outputs(3849));
    layer2_outputs(4220) <= '1';
    layer2_outputs(4221) <= not(layer1_outputs(849));
    layer2_outputs(4222) <= not(layer1_outputs(6271)) or (layer1_outputs(3738));
    layer2_outputs(4223) <= layer1_outputs(6546);
    layer2_outputs(4224) <= (layer1_outputs(4255)) and not (layer1_outputs(7539));
    layer2_outputs(4225) <= (layer1_outputs(903)) or (layer1_outputs(7196));
    layer2_outputs(4226) <= not((layer1_outputs(1203)) or (layer1_outputs(4606)));
    layer2_outputs(4227) <= not(layer1_outputs(317));
    layer2_outputs(4228) <= '1';
    layer2_outputs(4229) <= layer1_outputs(575);
    layer2_outputs(4230) <= not((layer1_outputs(2679)) or (layer1_outputs(2492)));
    layer2_outputs(4231) <= not(layer1_outputs(1386));
    layer2_outputs(4232) <= not((layer1_outputs(3146)) or (layer1_outputs(1752)));
    layer2_outputs(4233) <= '1';
    layer2_outputs(4234) <= not(layer1_outputs(5518));
    layer2_outputs(4235) <= '0';
    layer2_outputs(4236) <= (layer1_outputs(3537)) and not (layer1_outputs(1628));
    layer2_outputs(4237) <= not(layer1_outputs(2654));
    layer2_outputs(4238) <= (layer1_outputs(7068)) and not (layer1_outputs(5525));
    layer2_outputs(4239) <= not(layer1_outputs(1563)) or (layer1_outputs(688));
    layer2_outputs(4240) <= '1';
    layer2_outputs(4241) <= '0';
    layer2_outputs(4242) <= layer1_outputs(4702);
    layer2_outputs(4243) <= not((layer1_outputs(5294)) or (layer1_outputs(2482)));
    layer2_outputs(4244) <= not(layer1_outputs(3314)) or (layer1_outputs(6202));
    layer2_outputs(4245) <= not(layer1_outputs(4833)) or (layer1_outputs(212));
    layer2_outputs(4246) <= layer1_outputs(327);
    layer2_outputs(4247) <= '0';
    layer2_outputs(4248) <= '0';
    layer2_outputs(4249) <= (layer1_outputs(551)) or (layer1_outputs(3262));
    layer2_outputs(4250) <= not(layer1_outputs(3286));
    layer2_outputs(4251) <= not(layer1_outputs(3245)) or (layer1_outputs(2953));
    layer2_outputs(4252) <= (layer1_outputs(6806)) or (layer1_outputs(1549));
    layer2_outputs(4253) <= (layer1_outputs(125)) and not (layer1_outputs(3170));
    layer2_outputs(4254) <= (layer1_outputs(739)) and (layer1_outputs(426));
    layer2_outputs(4255) <= layer1_outputs(2591);
    layer2_outputs(4256) <= (layer1_outputs(5074)) and not (layer1_outputs(1447));
    layer2_outputs(4257) <= not(layer1_outputs(7377));
    layer2_outputs(4258) <= '1';
    layer2_outputs(4259) <= not((layer1_outputs(5000)) and (layer1_outputs(2506)));
    layer2_outputs(4260) <= '1';
    layer2_outputs(4261) <= (layer1_outputs(4507)) and (layer1_outputs(3204));
    layer2_outputs(4262) <= not(layer1_outputs(7200)) or (layer1_outputs(4722));
    layer2_outputs(4263) <= not(layer1_outputs(2999));
    layer2_outputs(4264) <= layer1_outputs(965);
    layer2_outputs(4265) <= not((layer1_outputs(5273)) and (layer1_outputs(7439)));
    layer2_outputs(4266) <= layer1_outputs(7183);
    layer2_outputs(4267) <= not(layer1_outputs(5099));
    layer2_outputs(4268) <= (layer1_outputs(1469)) and not (layer1_outputs(4823));
    layer2_outputs(4269) <= not((layer1_outputs(1149)) and (layer1_outputs(4440)));
    layer2_outputs(4270) <= layer1_outputs(7538);
    layer2_outputs(4271) <= (layer1_outputs(7650)) and not (layer1_outputs(6558));
    layer2_outputs(4272) <= not(layer1_outputs(5012));
    layer2_outputs(4273) <= '0';
    layer2_outputs(4274) <= not(layer1_outputs(1313));
    layer2_outputs(4275) <= layer1_outputs(6240);
    layer2_outputs(4276) <= (layer1_outputs(3965)) and (layer1_outputs(7386));
    layer2_outputs(4277) <= layer1_outputs(4259);
    layer2_outputs(4278) <= not((layer1_outputs(1992)) and (layer1_outputs(1167)));
    layer2_outputs(4279) <= not(layer1_outputs(3293)) or (layer1_outputs(2557));
    layer2_outputs(4280) <= '0';
    layer2_outputs(4281) <= (layer1_outputs(5794)) and (layer1_outputs(3410));
    layer2_outputs(4282) <= not(layer1_outputs(1080));
    layer2_outputs(4283) <= (layer1_outputs(3959)) and (layer1_outputs(336));
    layer2_outputs(4284) <= (layer1_outputs(3437)) and not (layer1_outputs(4775));
    layer2_outputs(4285) <= '0';
    layer2_outputs(4286) <= '0';
    layer2_outputs(4287) <= '0';
    layer2_outputs(4288) <= layer1_outputs(2216);
    layer2_outputs(4289) <= not(layer1_outputs(6241));
    layer2_outputs(4290) <= not(layer1_outputs(1399)) or (layer1_outputs(7275));
    layer2_outputs(4291) <= layer1_outputs(1957);
    layer2_outputs(4292) <= layer1_outputs(4184);
    layer2_outputs(4293) <= layer1_outputs(777);
    layer2_outputs(4294) <= layer1_outputs(5134);
    layer2_outputs(4295) <= layer1_outputs(1727);
    layer2_outputs(4296) <= not((layer1_outputs(3237)) or (layer1_outputs(4042)));
    layer2_outputs(4297) <= '1';
    layer2_outputs(4298) <= not(layer1_outputs(5250)) or (layer1_outputs(1761));
    layer2_outputs(4299) <= not(layer1_outputs(5074)) or (layer1_outputs(6292));
    layer2_outputs(4300) <= (layer1_outputs(5609)) and not (layer1_outputs(6536));
    layer2_outputs(4301) <= layer1_outputs(7021);
    layer2_outputs(4302) <= not(layer1_outputs(2785));
    layer2_outputs(4303) <= not((layer1_outputs(4962)) or (layer1_outputs(43)));
    layer2_outputs(4304) <= (layer1_outputs(1221)) and not (layer1_outputs(6407));
    layer2_outputs(4305) <= not((layer1_outputs(178)) xor (layer1_outputs(6283)));
    layer2_outputs(4306) <= not(layer1_outputs(6163));
    layer2_outputs(4307) <= layer1_outputs(3351);
    layer2_outputs(4308) <= not((layer1_outputs(7574)) or (layer1_outputs(1889)));
    layer2_outputs(4309) <= not(layer1_outputs(5133)) or (layer1_outputs(1794));
    layer2_outputs(4310) <= (layer1_outputs(3736)) and not (layer1_outputs(2195));
    layer2_outputs(4311) <= not((layer1_outputs(261)) or (layer1_outputs(907)));
    layer2_outputs(4312) <= not((layer1_outputs(437)) or (layer1_outputs(2659)));
    layer2_outputs(4313) <= not(layer1_outputs(6394)) or (layer1_outputs(2810));
    layer2_outputs(4314) <= (layer1_outputs(733)) and not (layer1_outputs(5226));
    layer2_outputs(4315) <= (layer1_outputs(7238)) or (layer1_outputs(4386));
    layer2_outputs(4316) <= (layer1_outputs(6297)) xor (layer1_outputs(344));
    layer2_outputs(4317) <= '1';
    layer2_outputs(4318) <= not(layer1_outputs(4532)) or (layer1_outputs(3073));
    layer2_outputs(4319) <= not(layer1_outputs(1867));
    layer2_outputs(4320) <= not((layer1_outputs(138)) or (layer1_outputs(1198)));
    layer2_outputs(4321) <= not(layer1_outputs(1421));
    layer2_outputs(4322) <= (layer1_outputs(617)) or (layer1_outputs(2385));
    layer2_outputs(4323) <= not((layer1_outputs(3066)) or (layer1_outputs(6529)));
    layer2_outputs(4324) <= not((layer1_outputs(4957)) or (layer1_outputs(5895)));
    layer2_outputs(4325) <= '0';
    layer2_outputs(4326) <= (layer1_outputs(5847)) and (layer1_outputs(668));
    layer2_outputs(4327) <= '1';
    layer2_outputs(4328) <= not(layer1_outputs(5393));
    layer2_outputs(4329) <= not((layer1_outputs(7523)) or (layer1_outputs(3289)));
    layer2_outputs(4330) <= '0';
    layer2_outputs(4331) <= '1';
    layer2_outputs(4332) <= layer1_outputs(5433);
    layer2_outputs(4333) <= layer1_outputs(2338);
    layer2_outputs(4334) <= not(layer1_outputs(3034));
    layer2_outputs(4335) <= layer1_outputs(4670);
    layer2_outputs(4336) <= (layer1_outputs(5465)) or (layer1_outputs(6169));
    layer2_outputs(4337) <= layer1_outputs(3427);
    layer2_outputs(4338) <= not((layer1_outputs(6954)) or (layer1_outputs(1036)));
    layer2_outputs(4339) <= (layer1_outputs(3025)) and (layer1_outputs(3963));
    layer2_outputs(4340) <= layer1_outputs(6853);
    layer2_outputs(4341) <= (layer1_outputs(6167)) and not (layer1_outputs(1869));
    layer2_outputs(4342) <= layer1_outputs(5978);
    layer2_outputs(4343) <= (layer1_outputs(396)) and not (layer1_outputs(2467));
    layer2_outputs(4344) <= layer1_outputs(1336);
    layer2_outputs(4345) <= not(layer1_outputs(7013));
    layer2_outputs(4346) <= not(layer1_outputs(5862));
    layer2_outputs(4347) <= not(layer1_outputs(3438)) or (layer1_outputs(5523));
    layer2_outputs(4348) <= not(layer1_outputs(1243));
    layer2_outputs(4349) <= not((layer1_outputs(5371)) and (layer1_outputs(5082)));
    layer2_outputs(4350) <= not(layer1_outputs(7161)) or (layer1_outputs(4314));
    layer2_outputs(4351) <= not((layer1_outputs(6108)) and (layer1_outputs(2453)));
    layer2_outputs(4352) <= not((layer1_outputs(1342)) or (layer1_outputs(904)));
    layer2_outputs(4353) <= not((layer1_outputs(6146)) and (layer1_outputs(4309)));
    layer2_outputs(4354) <= layer1_outputs(4320);
    layer2_outputs(4355) <= not((layer1_outputs(1560)) or (layer1_outputs(2753)));
    layer2_outputs(4356) <= (layer1_outputs(2629)) xor (layer1_outputs(6550));
    layer2_outputs(4357) <= (layer1_outputs(4340)) and (layer1_outputs(1908));
    layer2_outputs(4358) <= not(layer1_outputs(7447)) or (layer1_outputs(4544));
    layer2_outputs(4359) <= not(layer1_outputs(7173));
    layer2_outputs(4360) <= (layer1_outputs(7324)) and not (layer1_outputs(6966));
    layer2_outputs(4361) <= layer1_outputs(918);
    layer2_outputs(4362) <= not((layer1_outputs(5904)) and (layer1_outputs(5604)));
    layer2_outputs(4363) <= '0';
    layer2_outputs(4364) <= layer1_outputs(4534);
    layer2_outputs(4365) <= (layer1_outputs(3764)) or (layer1_outputs(5902));
    layer2_outputs(4366) <= '0';
    layer2_outputs(4367) <= (layer1_outputs(3473)) and (layer1_outputs(7057));
    layer2_outputs(4368) <= '0';
    layer2_outputs(4369) <= not((layer1_outputs(1764)) or (layer1_outputs(3800)));
    layer2_outputs(4370) <= (layer1_outputs(4034)) and not (layer1_outputs(3414));
    layer2_outputs(4371) <= not(layer1_outputs(1495));
    layer2_outputs(4372) <= (layer1_outputs(6659)) and not (layer1_outputs(2916));
    layer2_outputs(4373) <= (layer1_outputs(4164)) and (layer1_outputs(6431));
    layer2_outputs(4374) <= (layer1_outputs(5384)) and not (layer1_outputs(990));
    layer2_outputs(4375) <= not((layer1_outputs(1248)) and (layer1_outputs(5947)));
    layer2_outputs(4376) <= (layer1_outputs(2579)) or (layer1_outputs(3368));
    layer2_outputs(4377) <= layer1_outputs(1875);
    layer2_outputs(4378) <= layer1_outputs(427);
    layer2_outputs(4379) <= not(layer1_outputs(4368));
    layer2_outputs(4380) <= layer1_outputs(1420);
    layer2_outputs(4381) <= (layer1_outputs(745)) and not (layer1_outputs(3226));
    layer2_outputs(4382) <= (layer1_outputs(6121)) and not (layer1_outputs(1377));
    layer2_outputs(4383) <= (layer1_outputs(2815)) and not (layer1_outputs(4734));
    layer2_outputs(4384) <= not((layer1_outputs(6925)) and (layer1_outputs(4290)));
    layer2_outputs(4385) <= (layer1_outputs(7383)) and not (layer1_outputs(1232));
    layer2_outputs(4386) <= layer1_outputs(1048);
    layer2_outputs(4387) <= layer1_outputs(776);
    layer2_outputs(4388) <= '1';
    layer2_outputs(4389) <= not(layer1_outputs(2811));
    layer2_outputs(4390) <= not(layer1_outputs(1557)) or (layer1_outputs(3586));
    layer2_outputs(4391) <= (layer1_outputs(6488)) and (layer1_outputs(2603));
    layer2_outputs(4392) <= (layer1_outputs(802)) and not (layer1_outputs(7457));
    layer2_outputs(4393) <= '1';
    layer2_outputs(4394) <= not((layer1_outputs(2225)) and (layer1_outputs(2840)));
    layer2_outputs(4395) <= layer1_outputs(3976);
    layer2_outputs(4396) <= '0';
    layer2_outputs(4397) <= (layer1_outputs(4717)) or (layer1_outputs(725));
    layer2_outputs(4398) <= (layer1_outputs(1645)) and not (layer1_outputs(5574));
    layer2_outputs(4399) <= layer1_outputs(4005);
    layer2_outputs(4400) <= '0';
    layer2_outputs(4401) <= (layer1_outputs(1045)) and not (layer1_outputs(3074));
    layer2_outputs(4402) <= layer1_outputs(7198);
    layer2_outputs(4403) <= '0';
    layer2_outputs(4404) <= not(layer1_outputs(4551)) or (layer1_outputs(6491));
    layer2_outputs(4405) <= '1';
    layer2_outputs(4406) <= layer1_outputs(6686);
    layer2_outputs(4407) <= not((layer1_outputs(197)) and (layer1_outputs(4799)));
    layer2_outputs(4408) <= (layer1_outputs(192)) and not (layer1_outputs(4070));
    layer2_outputs(4409) <= layer1_outputs(7489);
    layer2_outputs(4410) <= layer1_outputs(224);
    layer2_outputs(4411) <= '0';
    layer2_outputs(4412) <= not(layer1_outputs(5024));
    layer2_outputs(4413) <= (layer1_outputs(5324)) xor (layer1_outputs(4032));
    layer2_outputs(4414) <= '0';
    layer2_outputs(4415) <= '1';
    layer2_outputs(4416) <= (layer1_outputs(5465)) and (layer1_outputs(6974));
    layer2_outputs(4417) <= not(layer1_outputs(1505)) or (layer1_outputs(5550));
    layer2_outputs(4418) <= layer1_outputs(5650);
    layer2_outputs(4419) <= '0';
    layer2_outputs(4420) <= layer1_outputs(3324);
    layer2_outputs(4421) <= (layer1_outputs(2014)) and (layer1_outputs(2716));
    layer2_outputs(4422) <= '1';
    layer2_outputs(4423) <= layer1_outputs(2657);
    layer2_outputs(4424) <= layer1_outputs(7107);
    layer2_outputs(4425) <= not((layer1_outputs(680)) or (layer1_outputs(1327)));
    layer2_outputs(4426) <= not((layer1_outputs(3572)) or (layer1_outputs(2392)));
    layer2_outputs(4427) <= not(layer1_outputs(6413)) or (layer1_outputs(1660));
    layer2_outputs(4428) <= '0';
    layer2_outputs(4429) <= layer1_outputs(1751);
    layer2_outputs(4430) <= not((layer1_outputs(3226)) or (layer1_outputs(3481)));
    layer2_outputs(4431) <= not(layer1_outputs(3380)) or (layer1_outputs(1672));
    layer2_outputs(4432) <= not(layer1_outputs(4873));
    layer2_outputs(4433) <= '1';
    layer2_outputs(4434) <= (layer1_outputs(6449)) and not (layer1_outputs(6919));
    layer2_outputs(4435) <= (layer1_outputs(6285)) and not (layer1_outputs(6223));
    layer2_outputs(4436) <= layer1_outputs(5726);
    layer2_outputs(4437) <= not(layer1_outputs(2027)) or (layer1_outputs(7420));
    layer2_outputs(4438) <= (layer1_outputs(2302)) or (layer1_outputs(3271));
    layer2_outputs(4439) <= layer1_outputs(3816);
    layer2_outputs(4440) <= not((layer1_outputs(3420)) and (layer1_outputs(3769)));
    layer2_outputs(4441) <= (layer1_outputs(2593)) and not (layer1_outputs(7476));
    layer2_outputs(4442) <= not(layer1_outputs(4427));
    layer2_outputs(4443) <= (layer1_outputs(4565)) and (layer1_outputs(2034));
    layer2_outputs(4444) <= (layer1_outputs(268)) or (layer1_outputs(2297));
    layer2_outputs(4445) <= layer1_outputs(1946);
    layer2_outputs(4446) <= (layer1_outputs(3756)) or (layer1_outputs(3579));
    layer2_outputs(4447) <= (layer1_outputs(6985)) and not (layer1_outputs(1035));
    layer2_outputs(4448) <= layer1_outputs(5350);
    layer2_outputs(4449) <= (layer1_outputs(6149)) and not (layer1_outputs(4192));
    layer2_outputs(4450) <= not((layer1_outputs(4068)) or (layer1_outputs(1912)));
    layer2_outputs(4451) <= (layer1_outputs(594)) or (layer1_outputs(5802));
    layer2_outputs(4452) <= (layer1_outputs(6656)) and not (layer1_outputs(2462));
    layer2_outputs(4453) <= layer1_outputs(6321);
    layer2_outputs(4454) <= not(layer1_outputs(7097)) or (layer1_outputs(605));
    layer2_outputs(4455) <= (layer1_outputs(7286)) and not (layer1_outputs(4003));
    layer2_outputs(4456) <= '0';
    layer2_outputs(4457) <= not(layer1_outputs(419)) or (layer1_outputs(3510));
    layer2_outputs(4458) <= layer1_outputs(6310);
    layer2_outputs(4459) <= not((layer1_outputs(1898)) and (layer1_outputs(6803)));
    layer2_outputs(4460) <= (layer1_outputs(4611)) and (layer1_outputs(7555));
    layer2_outputs(4461) <= not((layer1_outputs(2934)) or (layer1_outputs(4271)));
    layer2_outputs(4462) <= layer1_outputs(3126);
    layer2_outputs(4463) <= (layer1_outputs(934)) and not (layer1_outputs(4923));
    layer2_outputs(4464) <= layer1_outputs(3515);
    layer2_outputs(4465) <= (layer1_outputs(2830)) and not (layer1_outputs(4051));
    layer2_outputs(4466) <= layer1_outputs(7597);
    layer2_outputs(4467) <= layer1_outputs(5779);
    layer2_outputs(4468) <= not((layer1_outputs(3132)) and (layer1_outputs(3564)));
    layer2_outputs(4469) <= layer1_outputs(5973);
    layer2_outputs(4470) <= layer1_outputs(7428);
    layer2_outputs(4471) <= (layer1_outputs(6895)) and (layer1_outputs(3245));
    layer2_outputs(4472) <= not(layer1_outputs(3594)) or (layer1_outputs(6647));
    layer2_outputs(4473) <= not((layer1_outputs(5786)) or (layer1_outputs(1836)));
    layer2_outputs(4474) <= layer1_outputs(581);
    layer2_outputs(4475) <= '0';
    layer2_outputs(4476) <= (layer1_outputs(7268)) and (layer1_outputs(2004));
    layer2_outputs(4477) <= layer1_outputs(1122);
    layer2_outputs(4478) <= '0';
    layer2_outputs(4479) <= not((layer1_outputs(5336)) and (layer1_outputs(4710)));
    layer2_outputs(4480) <= not((layer1_outputs(83)) and (layer1_outputs(7192)));
    layer2_outputs(4481) <= (layer1_outputs(5715)) and not (layer1_outputs(5382));
    layer2_outputs(4482) <= (layer1_outputs(5931)) and (layer1_outputs(3512));
    layer2_outputs(4483) <= not(layer1_outputs(690)) or (layer1_outputs(912));
    layer2_outputs(4484) <= '0';
    layer2_outputs(4485) <= not((layer1_outputs(2930)) or (layer1_outputs(5140)));
    layer2_outputs(4486) <= layer1_outputs(4478);
    layer2_outputs(4487) <= '0';
    layer2_outputs(4488) <= not(layer1_outputs(6785));
    layer2_outputs(4489) <= layer1_outputs(3015);
    layer2_outputs(4490) <= not((layer1_outputs(7194)) or (layer1_outputs(1171)));
    layer2_outputs(4491) <= (layer1_outputs(1567)) and (layer1_outputs(305));
    layer2_outputs(4492) <= not(layer1_outputs(2352));
    layer2_outputs(4493) <= (layer1_outputs(1251)) and (layer1_outputs(7506));
    layer2_outputs(4494) <= '1';
    layer2_outputs(4495) <= layer1_outputs(1546);
    layer2_outputs(4496) <= layer1_outputs(1286);
    layer2_outputs(4497) <= not(layer1_outputs(4710)) or (layer1_outputs(5478));
    layer2_outputs(4498) <= not(layer1_outputs(5541)) or (layer1_outputs(6358));
    layer2_outputs(4499) <= not((layer1_outputs(6924)) or (layer1_outputs(1609)));
    layer2_outputs(4500) <= layer1_outputs(3905);
    layer2_outputs(4501) <= not((layer1_outputs(4892)) and (layer1_outputs(3750)));
    layer2_outputs(4502) <= not(layer1_outputs(4021));
    layer2_outputs(4503) <= not(layer1_outputs(1864));
    layer2_outputs(4504) <= not(layer1_outputs(4357));
    layer2_outputs(4505) <= layer1_outputs(1543);
    layer2_outputs(4506) <= (layer1_outputs(3641)) and (layer1_outputs(3048));
    layer2_outputs(4507) <= not((layer1_outputs(4495)) or (layer1_outputs(7591)));
    layer2_outputs(4508) <= not(layer1_outputs(7379));
    layer2_outputs(4509) <= not((layer1_outputs(2527)) or (layer1_outputs(3356)));
    layer2_outputs(4510) <= not((layer1_outputs(4060)) and (layer1_outputs(7457)));
    layer2_outputs(4511) <= (layer1_outputs(293)) and not (layer1_outputs(5711));
    layer2_outputs(4512) <= (layer1_outputs(6237)) or (layer1_outputs(852));
    layer2_outputs(4513) <= layer1_outputs(7050);
    layer2_outputs(4514) <= not(layer1_outputs(1542));
    layer2_outputs(4515) <= not(layer1_outputs(346));
    layer2_outputs(4516) <= not(layer1_outputs(7481));
    layer2_outputs(4517) <= not(layer1_outputs(6617)) or (layer1_outputs(7615));
    layer2_outputs(4518) <= not(layer1_outputs(6019)) or (layer1_outputs(7053));
    layer2_outputs(4519) <= not((layer1_outputs(2854)) or (layer1_outputs(7009)));
    layer2_outputs(4520) <= layer1_outputs(180);
    layer2_outputs(4521) <= layer1_outputs(5292);
    layer2_outputs(4522) <= (layer1_outputs(4978)) and not (layer1_outputs(390));
    layer2_outputs(4523) <= not((layer1_outputs(6084)) and (layer1_outputs(5998)));
    layer2_outputs(4524) <= '1';
    layer2_outputs(4525) <= layer1_outputs(6271);
    layer2_outputs(4526) <= (layer1_outputs(6395)) or (layer1_outputs(4825));
    layer2_outputs(4527) <= '1';
    layer2_outputs(4528) <= '1';
    layer2_outputs(4529) <= layer1_outputs(4405);
    layer2_outputs(4530) <= not((layer1_outputs(7297)) and (layer1_outputs(2236)));
    layer2_outputs(4531) <= layer1_outputs(3033);
    layer2_outputs(4532) <= not(layer1_outputs(1419)) or (layer1_outputs(5123));
    layer2_outputs(4533) <= '0';
    layer2_outputs(4534) <= not(layer1_outputs(3881));
    layer2_outputs(4535) <= not((layer1_outputs(6100)) xor (layer1_outputs(1951)));
    layer2_outputs(4536) <= not((layer1_outputs(4956)) or (layer1_outputs(3034)));
    layer2_outputs(4537) <= layer1_outputs(1298);
    layer2_outputs(4538) <= (layer1_outputs(7052)) or (layer1_outputs(6104));
    layer2_outputs(4539) <= (layer1_outputs(6116)) and not (layer1_outputs(1216));
    layer2_outputs(4540) <= layer1_outputs(1342);
    layer2_outputs(4541) <= layer1_outputs(4543);
    layer2_outputs(4542) <= '0';
    layer2_outputs(4543) <= not((layer1_outputs(5567)) and (layer1_outputs(483)));
    layer2_outputs(4544) <= layer1_outputs(6843);
    layer2_outputs(4545) <= not(layer1_outputs(3648));
    layer2_outputs(4546) <= not((layer1_outputs(1271)) and (layer1_outputs(673)));
    layer2_outputs(4547) <= (layer1_outputs(1219)) and (layer1_outputs(5584));
    layer2_outputs(4548) <= not(layer1_outputs(2841)) or (layer1_outputs(945));
    layer2_outputs(4549) <= not((layer1_outputs(4818)) and (layer1_outputs(6386)));
    layer2_outputs(4550) <= '1';
    layer2_outputs(4551) <= not(layer1_outputs(7578));
    layer2_outputs(4552) <= not((layer1_outputs(4998)) or (layer1_outputs(4364)));
    layer2_outputs(4553) <= '1';
    layer2_outputs(4554) <= not(layer1_outputs(3585));
    layer2_outputs(4555) <= layer1_outputs(5551);
    layer2_outputs(4556) <= layer1_outputs(6610);
    layer2_outputs(4557) <= not(layer1_outputs(6091)) or (layer1_outputs(5555));
    layer2_outputs(4558) <= layer1_outputs(1440);
    layer2_outputs(4559) <= (layer1_outputs(4802)) or (layer1_outputs(594));
    layer2_outputs(4560) <= not(layer1_outputs(58));
    layer2_outputs(4561) <= (layer1_outputs(549)) and not (layer1_outputs(291));
    layer2_outputs(4562) <= not(layer1_outputs(6823));
    layer2_outputs(4563) <= layer1_outputs(2725);
    layer2_outputs(4564) <= not((layer1_outputs(527)) and (layer1_outputs(3623)));
    layer2_outputs(4565) <= (layer1_outputs(6345)) and (layer1_outputs(4624));
    layer2_outputs(4566) <= not(layer1_outputs(6445));
    layer2_outputs(4567) <= not(layer1_outputs(5563)) or (layer1_outputs(365));
    layer2_outputs(4568) <= not(layer1_outputs(5329));
    layer2_outputs(4569) <= (layer1_outputs(1361)) or (layer1_outputs(3022));
    layer2_outputs(4570) <= layer1_outputs(3242);
    layer2_outputs(4571) <= not(layer1_outputs(1739));
    layer2_outputs(4572) <= not(layer1_outputs(4140));
    layer2_outputs(4573) <= (layer1_outputs(6127)) and (layer1_outputs(5515));
    layer2_outputs(4574) <= layer1_outputs(2960);
    layer2_outputs(4575) <= not(layer1_outputs(1659)) or (layer1_outputs(6930));
    layer2_outputs(4576) <= (layer1_outputs(1658)) or (layer1_outputs(5983));
    layer2_outputs(4577) <= layer1_outputs(7228);
    layer2_outputs(4578) <= not(layer1_outputs(6884)) or (layer1_outputs(4172));
    layer2_outputs(4579) <= layer1_outputs(2213);
    layer2_outputs(4580) <= '0';
    layer2_outputs(4581) <= layer1_outputs(481);
    layer2_outputs(4582) <= (layer1_outputs(6808)) xor (layer1_outputs(4911));
    layer2_outputs(4583) <= not(layer1_outputs(1196)) or (layer1_outputs(328));
    layer2_outputs(4584) <= not(layer1_outputs(6060)) or (layer1_outputs(5510));
    layer2_outputs(4585) <= layer1_outputs(6327);
    layer2_outputs(4586) <= not(layer1_outputs(3913));
    layer2_outputs(4587) <= layer1_outputs(4770);
    layer2_outputs(4588) <= not(layer1_outputs(5015));
    layer2_outputs(4589) <= layer1_outputs(1673);
    layer2_outputs(4590) <= not(layer1_outputs(6773));
    layer2_outputs(4591) <= (layer1_outputs(6859)) and not (layer1_outputs(3213));
    layer2_outputs(4592) <= not(layer1_outputs(5474)) or (layer1_outputs(3207));
    layer2_outputs(4593) <= '1';
    layer2_outputs(4594) <= not(layer1_outputs(537));
    layer2_outputs(4595) <= not(layer1_outputs(2209)) or (layer1_outputs(685));
    layer2_outputs(4596) <= not((layer1_outputs(1344)) or (layer1_outputs(7187)));
    layer2_outputs(4597) <= layer1_outputs(7510);
    layer2_outputs(4598) <= not((layer1_outputs(4635)) or (layer1_outputs(3151)));
    layer2_outputs(4599) <= layer1_outputs(7027);
    layer2_outputs(4600) <= not((layer1_outputs(7445)) and (layer1_outputs(6602)));
    layer2_outputs(4601) <= not(layer1_outputs(4184));
    layer2_outputs(4602) <= (layer1_outputs(2531)) or (layer1_outputs(3598));
    layer2_outputs(4603) <= not((layer1_outputs(2478)) or (layer1_outputs(2594)));
    layer2_outputs(4604) <= (layer1_outputs(4153)) and not (layer1_outputs(4239));
    layer2_outputs(4605) <= '1';
    layer2_outputs(4606) <= not(layer1_outputs(2179));
    layer2_outputs(4607) <= not((layer1_outputs(6848)) or (layer1_outputs(1974)));
    layer2_outputs(4608) <= '1';
    layer2_outputs(4609) <= not((layer1_outputs(272)) and (layer1_outputs(6812)));
    layer2_outputs(4610) <= (layer1_outputs(4011)) or (layer1_outputs(3304));
    layer2_outputs(4611) <= layer1_outputs(151);
    layer2_outputs(4612) <= layer1_outputs(2410);
    layer2_outputs(4613) <= layer1_outputs(3490);
    layer2_outputs(4614) <= (layer1_outputs(5516)) and not (layer1_outputs(2782));
    layer2_outputs(4615) <= (layer1_outputs(4416)) and not (layer1_outputs(5025));
    layer2_outputs(4616) <= '0';
    layer2_outputs(4617) <= (layer1_outputs(3799)) or (layer1_outputs(2419));
    layer2_outputs(4618) <= layer1_outputs(6117);
    layer2_outputs(4619) <= not((layer1_outputs(7025)) or (layer1_outputs(509)));
    layer2_outputs(4620) <= (layer1_outputs(567)) and (layer1_outputs(4379));
    layer2_outputs(4621) <= '1';
    layer2_outputs(4622) <= layer1_outputs(6835);
    layer2_outputs(4623) <= '0';
    layer2_outputs(4624) <= (layer1_outputs(7215)) and not (layer1_outputs(3833));
    layer2_outputs(4625) <= layer1_outputs(3032);
    layer2_outputs(4626) <= not(layer1_outputs(2279)) or (layer1_outputs(658));
    layer2_outputs(4627) <= not(layer1_outputs(38));
    layer2_outputs(4628) <= not((layer1_outputs(4876)) or (layer1_outputs(2823)));
    layer2_outputs(4629) <= (layer1_outputs(1791)) or (layer1_outputs(94));
    layer2_outputs(4630) <= layer1_outputs(5798);
    layer2_outputs(4631) <= layer1_outputs(722);
    layer2_outputs(4632) <= layer1_outputs(3087);
    layer2_outputs(4633) <= not(layer1_outputs(7005)) or (layer1_outputs(7335));
    layer2_outputs(4634) <= not(layer1_outputs(3403)) or (layer1_outputs(7579));
    layer2_outputs(4635) <= not(layer1_outputs(3316)) or (layer1_outputs(3254));
    layer2_outputs(4636) <= layer1_outputs(486);
    layer2_outputs(4637) <= '1';
    layer2_outputs(4638) <= '1';
    layer2_outputs(4639) <= not(layer1_outputs(5745)) or (layer1_outputs(475));
    layer2_outputs(4640) <= (layer1_outputs(2224)) and not (layer1_outputs(1631));
    layer2_outputs(4641) <= '1';
    layer2_outputs(4642) <= (layer1_outputs(434)) and not (layer1_outputs(807));
    layer2_outputs(4643) <= not(layer1_outputs(5753));
    layer2_outputs(4644) <= '1';
    layer2_outputs(4645) <= (layer1_outputs(4412)) and (layer1_outputs(6941));
    layer2_outputs(4646) <= (layer1_outputs(228)) and not (layer1_outputs(6342));
    layer2_outputs(4647) <= not(layer1_outputs(1199));
    layer2_outputs(4648) <= (layer1_outputs(6568)) and not (layer1_outputs(7370));
    layer2_outputs(4649) <= (layer1_outputs(5053)) and not (layer1_outputs(6847));
    layer2_outputs(4650) <= not(layer1_outputs(7504));
    layer2_outputs(4651) <= (layer1_outputs(2768)) xor (layer1_outputs(4178));
    layer2_outputs(4652) <= not((layer1_outputs(957)) and (layer1_outputs(4650)));
    layer2_outputs(4653) <= not((layer1_outputs(6354)) and (layer1_outputs(4202)));
    layer2_outputs(4654) <= '1';
    layer2_outputs(4655) <= (layer1_outputs(2303)) and (layer1_outputs(5326));
    layer2_outputs(4656) <= (layer1_outputs(1529)) and not (layer1_outputs(1344));
    layer2_outputs(4657) <= not(layer1_outputs(4075));
    layer2_outputs(4658) <= not(layer1_outputs(983)) or (layer1_outputs(59));
    layer2_outputs(4659) <= not((layer1_outputs(1746)) and (layer1_outputs(201)));
    layer2_outputs(4660) <= (layer1_outputs(6836)) or (layer1_outputs(1474));
    layer2_outputs(4661) <= not((layer1_outputs(3926)) or (layer1_outputs(2912)));
    layer2_outputs(4662) <= (layer1_outputs(545)) or (layer1_outputs(6503));
    layer2_outputs(4663) <= (layer1_outputs(5539)) or (layer1_outputs(66));
    layer2_outputs(4664) <= (layer1_outputs(5868)) and not (layer1_outputs(82));
    layer2_outputs(4665) <= (layer1_outputs(6343)) and (layer1_outputs(2437));
    layer2_outputs(4666) <= layer1_outputs(5492);
    layer2_outputs(4667) <= not(layer1_outputs(5505));
    layer2_outputs(4668) <= (layer1_outputs(1276)) and not (layer1_outputs(5588));
    layer2_outputs(4669) <= not(layer1_outputs(3648)) or (layer1_outputs(3969));
    layer2_outputs(4670) <= (layer1_outputs(5893)) and not (layer1_outputs(1308));
    layer2_outputs(4671) <= not((layer1_outputs(5353)) or (layer1_outputs(3477)));
    layer2_outputs(4672) <= not(layer1_outputs(6227)) or (layer1_outputs(952));
    layer2_outputs(4673) <= layer1_outputs(5648);
    layer2_outputs(4674) <= (layer1_outputs(5896)) or (layer1_outputs(59));
    layer2_outputs(4675) <= '1';
    layer2_outputs(4676) <= not(layer1_outputs(5772));
    layer2_outputs(4677) <= '0';
    layer2_outputs(4678) <= not((layer1_outputs(1113)) and (layer1_outputs(5768)));
    layer2_outputs(4679) <= (layer1_outputs(3453)) and (layer1_outputs(5252));
    layer2_outputs(4680) <= layer1_outputs(2388);
    layer2_outputs(4681) <= not((layer1_outputs(3099)) or (layer1_outputs(3601)));
    layer2_outputs(4682) <= '1';
    layer2_outputs(4683) <= (layer1_outputs(3917)) and not (layer1_outputs(5050));
    layer2_outputs(4684) <= not((layer1_outputs(2497)) and (layer1_outputs(4066)));
    layer2_outputs(4685) <= (layer1_outputs(6809)) and not (layer1_outputs(250));
    layer2_outputs(4686) <= (layer1_outputs(5281)) and (layer1_outputs(4007));
    layer2_outputs(4687) <= not((layer1_outputs(6082)) and (layer1_outputs(5828)));
    layer2_outputs(4688) <= not(layer1_outputs(3697));
    layer2_outputs(4689) <= not((layer1_outputs(6335)) xor (layer1_outputs(6762)));
    layer2_outputs(4690) <= not(layer1_outputs(851)) or (layer1_outputs(1373));
    layer2_outputs(4691) <= layer1_outputs(3900);
    layer2_outputs(4692) <= not(layer1_outputs(6444)) or (layer1_outputs(5013));
    layer2_outputs(4693) <= not(layer1_outputs(1183)) or (layer1_outputs(2221));
    layer2_outputs(4694) <= (layer1_outputs(5569)) and (layer1_outputs(3566));
    layer2_outputs(4695) <= not(layer1_outputs(6993)) or (layer1_outputs(4934));
    layer2_outputs(4696) <= not(layer1_outputs(7130)) or (layer1_outputs(1830));
    layer2_outputs(4697) <= not((layer1_outputs(7560)) and (layer1_outputs(3141)));
    layer2_outputs(4698) <= not(layer1_outputs(731)) or (layer1_outputs(769));
    layer2_outputs(4699) <= (layer1_outputs(7378)) and not (layer1_outputs(7286));
    layer2_outputs(4700) <= not(layer1_outputs(6259));
    layer2_outputs(4701) <= not(layer1_outputs(7047));
    layer2_outputs(4702) <= not(layer1_outputs(3438));
    layer2_outputs(4703) <= (layer1_outputs(367)) and not (layer1_outputs(648));
    layer2_outputs(4704) <= not(layer1_outputs(1889));
    layer2_outputs(4705) <= (layer1_outputs(890)) and not (layer1_outputs(2314));
    layer2_outputs(4706) <= (layer1_outputs(7592)) and not (layer1_outputs(5385));
    layer2_outputs(4707) <= '0';
    layer2_outputs(4708) <= not(layer1_outputs(2032));
    layer2_outputs(4709) <= (layer1_outputs(5965)) and not (layer1_outputs(6666));
    layer2_outputs(4710) <= layer1_outputs(4889);
    layer2_outputs(4711) <= layer1_outputs(7319);
    layer2_outputs(4712) <= (layer1_outputs(2428)) xor (layer1_outputs(1820));
    layer2_outputs(4713) <= (layer1_outputs(5933)) and (layer1_outputs(4887));
    layer2_outputs(4714) <= not(layer1_outputs(1640));
    layer2_outputs(4715) <= (layer1_outputs(1740)) and not (layer1_outputs(7651));
    layer2_outputs(4716) <= not(layer1_outputs(6063)) or (layer1_outputs(5542));
    layer2_outputs(4717) <= layer1_outputs(2415);
    layer2_outputs(4718) <= layer1_outputs(333);
    layer2_outputs(4719) <= not(layer1_outputs(3369)) or (layer1_outputs(4429));
    layer2_outputs(4720) <= layer1_outputs(7251);
    layer2_outputs(4721) <= layer1_outputs(5275);
    layer2_outputs(4722) <= '0';
    layer2_outputs(4723) <= '1';
    layer2_outputs(4724) <= not(layer1_outputs(7348)) or (layer1_outputs(3415));
    layer2_outputs(4725) <= not(layer1_outputs(4576));
    layer2_outputs(4726) <= (layer1_outputs(1777)) and (layer1_outputs(7113));
    layer2_outputs(4727) <= not(layer1_outputs(5854));
    layer2_outputs(4728) <= not((layer1_outputs(644)) and (layer1_outputs(4800)));
    layer2_outputs(4729) <= layer1_outputs(6661);
    layer2_outputs(4730) <= '0';
    layer2_outputs(4731) <= not(layer1_outputs(4678)) or (layer1_outputs(68));
    layer2_outputs(4732) <= not((layer1_outputs(7163)) and (layer1_outputs(4497)));
    layer2_outputs(4733) <= layer1_outputs(1739);
    layer2_outputs(4734) <= (layer1_outputs(2403)) or (layer1_outputs(1483));
    layer2_outputs(4735) <= not(layer1_outputs(5527));
    layer2_outputs(4736) <= (layer1_outputs(256)) or (layer1_outputs(3273));
    layer2_outputs(4737) <= not(layer1_outputs(3885));
    layer2_outputs(4738) <= (layer1_outputs(7411)) and not (layer1_outputs(7133));
    layer2_outputs(4739) <= layer1_outputs(6429);
    layer2_outputs(4740) <= (layer1_outputs(5816)) or (layer1_outputs(5460));
    layer2_outputs(4741) <= not(layer1_outputs(3542));
    layer2_outputs(4742) <= layer1_outputs(3490);
    layer2_outputs(4743) <= not(layer1_outputs(3548));
    layer2_outputs(4744) <= layer1_outputs(3596);
    layer2_outputs(4745) <= '1';
    layer2_outputs(4746) <= (layer1_outputs(1139)) and not (layer1_outputs(1397));
    layer2_outputs(4747) <= layer1_outputs(871);
    layer2_outputs(4748) <= (layer1_outputs(1099)) and not (layer1_outputs(5032));
    layer2_outputs(4749) <= not(layer1_outputs(6565));
    layer2_outputs(4750) <= (layer1_outputs(2155)) and not (layer1_outputs(3669));
    layer2_outputs(4751) <= not(layer1_outputs(2959));
    layer2_outputs(4752) <= (layer1_outputs(3416)) or (layer1_outputs(3262));
    layer2_outputs(4753) <= (layer1_outputs(2456)) and (layer1_outputs(5856));
    layer2_outputs(4754) <= layer1_outputs(459);
    layer2_outputs(4755) <= not(layer1_outputs(2897));
    layer2_outputs(4756) <= (layer1_outputs(3635)) and not (layer1_outputs(5208));
    layer2_outputs(4757) <= not((layer1_outputs(1655)) xor (layer1_outputs(2734)));
    layer2_outputs(4758) <= layer1_outputs(1051);
    layer2_outputs(4759) <= '0';
    layer2_outputs(4760) <= (layer1_outputs(798)) and (layer1_outputs(1709));
    layer2_outputs(4761) <= '1';
    layer2_outputs(4762) <= not(layer1_outputs(4851)) or (layer1_outputs(4583));
    layer2_outputs(4763) <= '0';
    layer2_outputs(4764) <= not(layer1_outputs(1223)) or (layer1_outputs(5010));
    layer2_outputs(4765) <= not(layer1_outputs(4029));
    layer2_outputs(4766) <= not(layer1_outputs(7001)) or (layer1_outputs(2300));
    layer2_outputs(4767) <= layer1_outputs(5901);
    layer2_outputs(4768) <= (layer1_outputs(2723)) and not (layer1_outputs(7501));
    layer2_outputs(4769) <= not(layer1_outputs(5005)) or (layer1_outputs(3468));
    layer2_outputs(4770) <= not(layer1_outputs(2511));
    layer2_outputs(4771) <= not(layer1_outputs(2903));
    layer2_outputs(4772) <= '1';
    layer2_outputs(4773) <= not(layer1_outputs(6721));
    layer2_outputs(4774) <= not(layer1_outputs(5729)) or (layer1_outputs(3765));
    layer2_outputs(4775) <= not(layer1_outputs(1776)) or (layer1_outputs(5157));
    layer2_outputs(4776) <= layer1_outputs(6845);
    layer2_outputs(4777) <= layer1_outputs(6192);
    layer2_outputs(4778) <= (layer1_outputs(2622)) or (layer1_outputs(3023));
    layer2_outputs(4779) <= not((layer1_outputs(554)) or (layer1_outputs(2210)));
    layer2_outputs(4780) <= layer1_outputs(5448);
    layer2_outputs(4781) <= (layer1_outputs(3194)) and not (layer1_outputs(1983));
    layer2_outputs(4782) <= not(layer1_outputs(3270));
    layer2_outputs(4783) <= not((layer1_outputs(5500)) or (layer1_outputs(4179)));
    layer2_outputs(4784) <= (layer1_outputs(4860)) and (layer1_outputs(1129));
    layer2_outputs(4785) <= not(layer1_outputs(814));
    layer2_outputs(4786) <= (layer1_outputs(7201)) and not (layer1_outputs(4332));
    layer2_outputs(4787) <= (layer1_outputs(7385)) and not (layer1_outputs(3894));
    layer2_outputs(4788) <= '1';
    layer2_outputs(4789) <= not(layer1_outputs(2006)) or (layer1_outputs(4705));
    layer2_outputs(4790) <= not(layer1_outputs(1408)) or (layer1_outputs(2404));
    layer2_outputs(4791) <= not((layer1_outputs(251)) and (layer1_outputs(2948)));
    layer2_outputs(4792) <= '1';
    layer2_outputs(4793) <= (layer1_outputs(4038)) and not (layer1_outputs(4974));
    layer2_outputs(4794) <= not(layer1_outputs(5959));
    layer2_outputs(4795) <= '0';
    layer2_outputs(4796) <= (layer1_outputs(2925)) and (layer1_outputs(4404));
    layer2_outputs(4797) <= not(layer1_outputs(5518));
    layer2_outputs(4798) <= '1';
    layer2_outputs(4799) <= layer1_outputs(6596);
    layer2_outputs(4800) <= not(layer1_outputs(2416));
    layer2_outputs(4801) <= not(layer1_outputs(1575)) or (layer1_outputs(2244));
    layer2_outputs(4802) <= '1';
    layer2_outputs(4803) <= not(layer1_outputs(6915));
    layer2_outputs(4804) <= not((layer1_outputs(1121)) xor (layer1_outputs(564)));
    layer2_outputs(4805) <= (layer1_outputs(2174)) and not (layer1_outputs(3712));
    layer2_outputs(4806) <= not((layer1_outputs(202)) or (layer1_outputs(7381)));
    layer2_outputs(4807) <= not(layer1_outputs(5718));
    layer2_outputs(4808) <= not(layer1_outputs(3851)) or (layer1_outputs(4695));
    layer2_outputs(4809) <= not(layer1_outputs(1666)) or (layer1_outputs(74));
    layer2_outputs(4810) <= layer1_outputs(1078);
    layer2_outputs(4811) <= not(layer1_outputs(3038));
    layer2_outputs(4812) <= not((layer1_outputs(3197)) or (layer1_outputs(7572)));
    layer2_outputs(4813) <= not(layer1_outputs(4729));
    layer2_outputs(4814) <= '0';
    layer2_outputs(4815) <= not((layer1_outputs(6005)) or (layer1_outputs(183)));
    layer2_outputs(4816) <= '1';
    layer2_outputs(4817) <= (layer1_outputs(1979)) xor (layer1_outputs(7210));
    layer2_outputs(4818) <= (layer1_outputs(3930)) and (layer1_outputs(180));
    layer2_outputs(4819) <= not((layer1_outputs(7607)) and (layer1_outputs(6814)));
    layer2_outputs(4820) <= '0';
    layer2_outputs(4821) <= not(layer1_outputs(1853));
    layer2_outputs(4822) <= layer1_outputs(340);
    layer2_outputs(4823) <= not(layer1_outputs(6882));
    layer2_outputs(4824) <= '0';
    layer2_outputs(4825) <= layer1_outputs(6817);
    layer2_outputs(4826) <= (layer1_outputs(4526)) xor (layer1_outputs(2794));
    layer2_outputs(4827) <= not(layer1_outputs(5910)) or (layer1_outputs(3074));
    layer2_outputs(4828) <= '1';
    layer2_outputs(4829) <= (layer1_outputs(4072)) and not (layer1_outputs(3019));
    layer2_outputs(4830) <= not((layer1_outputs(932)) or (layer1_outputs(6867)));
    layer2_outputs(4831) <= not(layer1_outputs(4402));
    layer2_outputs(4832) <= not(layer1_outputs(4843));
    layer2_outputs(4833) <= (layer1_outputs(7657)) and not (layer1_outputs(6737));
    layer2_outputs(4834) <= '0';
    layer2_outputs(4835) <= layer1_outputs(565);
    layer2_outputs(4836) <= not(layer1_outputs(6714));
    layer2_outputs(4837) <= not(layer1_outputs(3135));
    layer2_outputs(4838) <= not(layer1_outputs(3585));
    layer2_outputs(4839) <= (layer1_outputs(6059)) or (layer1_outputs(7251));
    layer2_outputs(4840) <= (layer1_outputs(5625)) and not (layer1_outputs(4000));
    layer2_outputs(4841) <= layer1_outputs(386);
    layer2_outputs(4842) <= not(layer1_outputs(476));
    layer2_outputs(4843) <= (layer1_outputs(6039)) or (layer1_outputs(2873));
    layer2_outputs(4844) <= layer1_outputs(1250);
    layer2_outputs(4845) <= layer1_outputs(5526);
    layer2_outputs(4846) <= not(layer1_outputs(5118));
    layer2_outputs(4847) <= (layer1_outputs(2858)) and not (layer1_outputs(57));
    layer2_outputs(4848) <= not(layer1_outputs(5806));
    layer2_outputs(4849) <= not(layer1_outputs(771));
    layer2_outputs(4850) <= (layer1_outputs(4712)) and not (layer1_outputs(5200));
    layer2_outputs(4851) <= layer1_outputs(6206);
    layer2_outputs(4852) <= layer1_outputs(4826);
    layer2_outputs(4853) <= not(layer1_outputs(2139)) or (layer1_outputs(6163));
    layer2_outputs(4854) <= not((layer1_outputs(4132)) and (layer1_outputs(3283)));
    layer2_outputs(4855) <= not(layer1_outputs(6328)) or (layer1_outputs(3868));
    layer2_outputs(4856) <= (layer1_outputs(940)) and (layer1_outputs(474));
    layer2_outputs(4857) <= not(layer1_outputs(4433)) or (layer1_outputs(1589));
    layer2_outputs(4858) <= not(layer1_outputs(5245));
    layer2_outputs(4859) <= '0';
    layer2_outputs(4860) <= (layer1_outputs(6292)) or (layer1_outputs(5534));
    layer2_outputs(4861) <= not((layer1_outputs(348)) and (layer1_outputs(6577)));
    layer2_outputs(4862) <= (layer1_outputs(3699)) and not (layer1_outputs(6704));
    layer2_outputs(4863) <= not(layer1_outputs(5981)) or (layer1_outputs(7516));
    layer2_outputs(4864) <= layer1_outputs(5368);
    layer2_outputs(4865) <= layer1_outputs(1758);
    layer2_outputs(4866) <= (layer1_outputs(5568)) and not (layer1_outputs(4295));
    layer2_outputs(4867) <= (layer1_outputs(5874)) or (layer1_outputs(7536));
    layer2_outputs(4868) <= not(layer1_outputs(1999)) or (layer1_outputs(6144));
    layer2_outputs(4869) <= not(layer1_outputs(3345)) or (layer1_outputs(6589));
    layer2_outputs(4870) <= not(layer1_outputs(184));
    layer2_outputs(4871) <= not(layer1_outputs(3900));
    layer2_outputs(4872) <= not((layer1_outputs(7067)) or (layer1_outputs(3444)));
    layer2_outputs(4873) <= layer1_outputs(3692);
    layer2_outputs(4874) <= not((layer1_outputs(6249)) or (layer1_outputs(4063)));
    layer2_outputs(4875) <= not((layer1_outputs(3303)) or (layer1_outputs(3745)));
    layer2_outputs(4876) <= not(layer1_outputs(1873)) or (layer1_outputs(4190));
    layer2_outputs(4877) <= not(layer1_outputs(2017)) or (layer1_outputs(7279));
    layer2_outputs(4878) <= not((layer1_outputs(488)) and (layer1_outputs(7527)));
    layer2_outputs(4879) <= (layer1_outputs(4176)) or (layer1_outputs(3329));
    layer2_outputs(4880) <= '1';
    layer2_outputs(4881) <= not(layer1_outputs(5028));
    layer2_outputs(4882) <= not((layer1_outputs(4107)) or (layer1_outputs(1586)));
    layer2_outputs(4883) <= not((layer1_outputs(5444)) and (layer1_outputs(205)));
    layer2_outputs(4884) <= not((layer1_outputs(7529)) and (layer1_outputs(861)));
    layer2_outputs(4885) <= '1';
    layer2_outputs(4886) <= (layer1_outputs(4754)) and not (layer1_outputs(989));
    layer2_outputs(4887) <= (layer1_outputs(176)) and not (layer1_outputs(778));
    layer2_outputs(4888) <= not(layer1_outputs(6017)) or (layer1_outputs(682));
    layer2_outputs(4889) <= not(layer1_outputs(219)) or (layer1_outputs(6621));
    layer2_outputs(4890) <= (layer1_outputs(1552)) or (layer1_outputs(6800));
    layer2_outputs(4891) <= '1';
    layer2_outputs(4892) <= (layer1_outputs(6684)) and (layer1_outputs(4914));
    layer2_outputs(4893) <= (layer1_outputs(1031)) and (layer1_outputs(3149));
    layer2_outputs(4894) <= layer1_outputs(6092);
    layer2_outputs(4895) <= '1';
    layer2_outputs(4896) <= not(layer1_outputs(5595)) or (layer1_outputs(4292));
    layer2_outputs(4897) <= not(layer1_outputs(4594));
    layer2_outputs(4898) <= not(layer1_outputs(203));
    layer2_outputs(4899) <= layer1_outputs(5579);
    layer2_outputs(4900) <= (layer1_outputs(3713)) and (layer1_outputs(6588));
    layer2_outputs(4901) <= not(layer1_outputs(7623));
    layer2_outputs(4902) <= layer1_outputs(3324);
    layer2_outputs(4903) <= (layer1_outputs(3600)) and not (layer1_outputs(4506));
    layer2_outputs(4904) <= layer1_outputs(7207);
    layer2_outputs(4905) <= not(layer1_outputs(3725)) or (layer1_outputs(7032));
    layer2_outputs(4906) <= '1';
    layer2_outputs(4907) <= (layer1_outputs(6490)) or (layer1_outputs(233));
    layer2_outputs(4908) <= not((layer1_outputs(3387)) and (layer1_outputs(6486)));
    layer2_outputs(4909) <= not((layer1_outputs(362)) or (layer1_outputs(6692)));
    layer2_outputs(4910) <= (layer1_outputs(6414)) and (layer1_outputs(2659));
    layer2_outputs(4911) <= not(layer1_outputs(3160));
    layer2_outputs(4912) <= (layer1_outputs(6278)) and (layer1_outputs(7264));
    layer2_outputs(4913) <= (layer1_outputs(2683)) xor (layer1_outputs(730));
    layer2_outputs(4914) <= (layer1_outputs(703)) and (layer1_outputs(4017));
    layer2_outputs(4915) <= not(layer1_outputs(168));
    layer2_outputs(4916) <= '0';
    layer2_outputs(4917) <= (layer1_outputs(2277)) xor (layer1_outputs(1243));
    layer2_outputs(4918) <= (layer1_outputs(3670)) or (layer1_outputs(350));
    layer2_outputs(4919) <= (layer1_outputs(4218)) and not (layer1_outputs(3563));
    layer2_outputs(4920) <= not((layer1_outputs(1193)) and (layer1_outputs(2701)));
    layer2_outputs(4921) <= layer1_outputs(7399);
    layer2_outputs(4922) <= not(layer1_outputs(3197));
    layer2_outputs(4923) <= '1';
    layer2_outputs(4924) <= not(layer1_outputs(2502));
    layer2_outputs(4925) <= '1';
    layer2_outputs(4926) <= (layer1_outputs(924)) or (layer1_outputs(4687));
    layer2_outputs(4927) <= not(layer1_outputs(1661)) or (layer1_outputs(4839));
    layer2_outputs(4928) <= layer1_outputs(4858);
    layer2_outputs(4929) <= (layer1_outputs(4571)) or (layer1_outputs(1785));
    layer2_outputs(4930) <= not((layer1_outputs(1927)) xor (layer1_outputs(289)));
    layer2_outputs(4931) <= not((layer1_outputs(2497)) or (layer1_outputs(2050)));
    layer2_outputs(4932) <= not(layer1_outputs(6099));
    layer2_outputs(4933) <= not((layer1_outputs(4920)) and (layer1_outputs(5840)));
    layer2_outputs(4934) <= layer1_outputs(190);
    layer2_outputs(4935) <= layer1_outputs(3480);
    layer2_outputs(4936) <= not(layer1_outputs(5409)) or (layer1_outputs(2931));
    layer2_outputs(4937) <= not(layer1_outputs(5687)) or (layer1_outputs(6054));
    layer2_outputs(4938) <= (layer1_outputs(3806)) and (layer1_outputs(4605));
    layer2_outputs(4939) <= layer1_outputs(4298);
    layer2_outputs(4940) <= '0';
    layer2_outputs(4941) <= layer1_outputs(7469);
    layer2_outputs(4942) <= not(layer1_outputs(7405));
    layer2_outputs(4943) <= layer1_outputs(6541);
    layer2_outputs(4944) <= not(layer1_outputs(7533));
    layer2_outputs(4945) <= (layer1_outputs(5397)) and not (layer1_outputs(7669));
    layer2_outputs(4946) <= not(layer1_outputs(46));
    layer2_outputs(4947) <= not((layer1_outputs(5433)) and (layer1_outputs(6844)));
    layer2_outputs(4948) <= (layer1_outputs(4335)) or (layer1_outputs(7647));
    layer2_outputs(4949) <= (layer1_outputs(5480)) and not (layer1_outputs(4683));
    layer2_outputs(4950) <= (layer1_outputs(1317)) and not (layer1_outputs(2849));
    layer2_outputs(4951) <= (layer1_outputs(4672)) or (layer1_outputs(1394));
    layer2_outputs(4952) <= '0';
    layer2_outputs(4953) <= not((layer1_outputs(7270)) or (layer1_outputs(5996)));
    layer2_outputs(4954) <= layer1_outputs(3062);
    layer2_outputs(4955) <= '0';
    layer2_outputs(4956) <= (layer1_outputs(2439)) and not (layer1_outputs(1002));
    layer2_outputs(4957) <= (layer1_outputs(5150)) or (layer1_outputs(2968));
    layer2_outputs(4958) <= not(layer1_outputs(6832));
    layer2_outputs(4959) <= (layer1_outputs(3103)) or (layer1_outputs(1015));
    layer2_outputs(4960) <= not(layer1_outputs(7585));
    layer2_outputs(4961) <= not(layer1_outputs(4971)) or (layer1_outputs(2661));
    layer2_outputs(4962) <= not((layer1_outputs(3492)) and (layer1_outputs(1355)));
    layer2_outputs(4963) <= (layer1_outputs(2892)) and (layer1_outputs(614));
    layer2_outputs(4964) <= not(layer1_outputs(6982));
    layer2_outputs(4965) <= layer1_outputs(5088);
    layer2_outputs(4966) <= layer1_outputs(1638);
    layer2_outputs(4967) <= layer1_outputs(341);
    layer2_outputs(4968) <= (layer1_outputs(779)) and (layer1_outputs(805));
    layer2_outputs(4969) <= layer1_outputs(1708);
    layer2_outputs(4970) <= layer1_outputs(5678);
    layer2_outputs(4971) <= not(layer1_outputs(1580));
    layer2_outputs(4972) <= not((layer1_outputs(52)) and (layer1_outputs(831)));
    layer2_outputs(4973) <= '0';
    layer2_outputs(4974) <= not(layer1_outputs(190));
    layer2_outputs(4975) <= (layer1_outputs(7257)) xor (layer1_outputs(2999));
    layer2_outputs(4976) <= layer1_outputs(5551);
    layer2_outputs(4977) <= layer1_outputs(983);
    layer2_outputs(4978) <= (layer1_outputs(3784)) or (layer1_outputs(6942));
    layer2_outputs(4979) <= '1';
    layer2_outputs(4980) <= not(layer1_outputs(4340));
    layer2_outputs(4981) <= '0';
    layer2_outputs(4982) <= '0';
    layer2_outputs(4983) <= (layer1_outputs(977)) or (layer1_outputs(5378));
    layer2_outputs(4984) <= not((layer1_outputs(6657)) or (layer1_outputs(7401)));
    layer2_outputs(4985) <= not((layer1_outputs(5155)) and (layer1_outputs(1719)));
    layer2_outputs(4986) <= '1';
    layer2_outputs(4987) <= (layer1_outputs(1695)) or (layer1_outputs(1541));
    layer2_outputs(4988) <= '0';
    layer2_outputs(4989) <= not(layer1_outputs(5749));
    layer2_outputs(4990) <= not(layer1_outputs(139));
    layer2_outputs(4991) <= not(layer1_outputs(2823)) or (layer1_outputs(2791));
    layer2_outputs(4992) <= (layer1_outputs(5073)) or (layer1_outputs(7176));
    layer2_outputs(4993) <= '1';
    layer2_outputs(4994) <= (layer1_outputs(761)) or (layer1_outputs(6593));
    layer2_outputs(4995) <= (layer1_outputs(2833)) and not (layer1_outputs(2093));
    layer2_outputs(4996) <= '1';
    layer2_outputs(4997) <= (layer1_outputs(5811)) and not (layer1_outputs(4343));
    layer2_outputs(4998) <= layer1_outputs(6501);
    layer2_outputs(4999) <= (layer1_outputs(604)) and not (layer1_outputs(2741));
    layer2_outputs(5000) <= '0';
    layer2_outputs(5001) <= (layer1_outputs(7427)) and not (layer1_outputs(4635));
    layer2_outputs(5002) <= (layer1_outputs(5889)) and (layer1_outputs(837));
    layer2_outputs(5003) <= layer1_outputs(6093);
    layer2_outputs(5004) <= '1';
    layer2_outputs(5005) <= '0';
    layer2_outputs(5006) <= '0';
    layer2_outputs(5007) <= layer1_outputs(5763);
    layer2_outputs(5008) <= not(layer1_outputs(6116)) or (layer1_outputs(7213));
    layer2_outputs(5009) <= (layer1_outputs(5564)) and (layer1_outputs(7653));
    layer2_outputs(5010) <= not(layer1_outputs(3279));
    layer2_outputs(5011) <= (layer1_outputs(5023)) and (layer1_outputs(668));
    layer2_outputs(5012) <= not(layer1_outputs(6485));
    layer2_outputs(5013) <= '0';
    layer2_outputs(5014) <= '1';
    layer2_outputs(5015) <= not(layer1_outputs(6961));
    layer2_outputs(5016) <= (layer1_outputs(6841)) and not (layer1_outputs(4808));
    layer2_outputs(5017) <= not(layer1_outputs(5336)) or (layer1_outputs(3815));
    layer2_outputs(5018) <= layer1_outputs(5230);
    layer2_outputs(5019) <= layer1_outputs(16);
    layer2_outputs(5020) <= layer1_outputs(4089);
    layer2_outputs(5021) <= not(layer1_outputs(6530));
    layer2_outputs(5022) <= (layer1_outputs(3828)) or (layer1_outputs(1389));
    layer2_outputs(5023) <= not(layer1_outputs(6822)) or (layer1_outputs(5881));
    layer2_outputs(5024) <= (layer1_outputs(5754)) and not (layer1_outputs(1053));
    layer2_outputs(5025) <= '1';
    layer2_outputs(5026) <= (layer1_outputs(1720)) and not (layer1_outputs(6909));
    layer2_outputs(5027) <= (layer1_outputs(1253)) and not (layer1_outputs(3326));
    layer2_outputs(5028) <= not(layer1_outputs(4237));
    layer2_outputs(5029) <= (layer1_outputs(6081)) and not (layer1_outputs(366));
    layer2_outputs(5030) <= not(layer1_outputs(5867)) or (layer1_outputs(3182));
    layer2_outputs(5031) <= '0';
    layer2_outputs(5032) <= not(layer1_outputs(3230)) or (layer1_outputs(3388));
    layer2_outputs(5033) <= not((layer1_outputs(1390)) or (layer1_outputs(7558)));
    layer2_outputs(5034) <= not(layer1_outputs(1175));
    layer2_outputs(5035) <= (layer1_outputs(6700)) and not (layer1_outputs(3098));
    layer2_outputs(5036) <= layer1_outputs(5627);
    layer2_outputs(5037) <= '1';
    layer2_outputs(5038) <= not(layer1_outputs(2369));
    layer2_outputs(5039) <= (layer1_outputs(4746)) or (layer1_outputs(3790));
    layer2_outputs(5040) <= '1';
    layer2_outputs(5041) <= not(layer1_outputs(3427));
    layer2_outputs(5042) <= (layer1_outputs(3955)) and not (layer1_outputs(6887));
    layer2_outputs(5043) <= (layer1_outputs(493)) or (layer1_outputs(2457));
    layer2_outputs(5044) <= layer1_outputs(6110);
    layer2_outputs(5045) <= not((layer1_outputs(7049)) and (layer1_outputs(7576)));
    layer2_outputs(5046) <= '1';
    layer2_outputs(5047) <= not(layer1_outputs(4125)) or (layer1_outputs(7379));
    layer2_outputs(5048) <= not(layer1_outputs(2181)) or (layer1_outputs(4389));
    layer2_outputs(5049) <= (layer1_outputs(1300)) and not (layer1_outputs(2539));
    layer2_outputs(5050) <= '0';
    layer2_outputs(5051) <= (layer1_outputs(3990)) and not (layer1_outputs(2830));
    layer2_outputs(5052) <= '1';
    layer2_outputs(5053) <= (layer1_outputs(5845)) and not (layer1_outputs(5778));
    layer2_outputs(5054) <= (layer1_outputs(1050)) and (layer1_outputs(5738));
    layer2_outputs(5055) <= layer1_outputs(1173);
    layer2_outputs(5056) <= layer1_outputs(4587);
    layer2_outputs(5057) <= not(layer1_outputs(1257)) or (layer1_outputs(5065));
    layer2_outputs(5058) <= (layer1_outputs(4857)) and not (layer1_outputs(5354));
    layer2_outputs(5059) <= not(layer1_outputs(7005)) or (layer1_outputs(3799));
    layer2_outputs(5060) <= (layer1_outputs(7276)) and not (layer1_outputs(1006));
    layer2_outputs(5061) <= not(layer1_outputs(5772));
    layer2_outputs(5062) <= not(layer1_outputs(374));
    layer2_outputs(5063) <= not((layer1_outputs(4789)) and (layer1_outputs(2209)));
    layer2_outputs(5064) <= not(layer1_outputs(7409));
    layer2_outputs(5065) <= '0';
    layer2_outputs(5066) <= not(layer1_outputs(2376)) or (layer1_outputs(4426));
    layer2_outputs(5067) <= (layer1_outputs(3748)) or (layer1_outputs(3575));
    layer2_outputs(5068) <= not((layer1_outputs(6859)) and (layer1_outputs(6198)));
    layer2_outputs(5069) <= not(layer1_outputs(765));
    layer2_outputs(5070) <= (layer1_outputs(2783)) and not (layer1_outputs(6791));
    layer2_outputs(5071) <= (layer1_outputs(5)) or (layer1_outputs(428));
    layer2_outputs(5072) <= (layer1_outputs(6791)) and not (layer1_outputs(5280));
    layer2_outputs(5073) <= not((layer1_outputs(4525)) or (layer1_outputs(6968)));
    layer2_outputs(5074) <= layer1_outputs(3584);
    layer2_outputs(5075) <= (layer1_outputs(2211)) and not (layer1_outputs(4624));
    layer2_outputs(5076) <= layer1_outputs(6425);
    layer2_outputs(5077) <= (layer1_outputs(2058)) and (layer1_outputs(2844));
    layer2_outputs(5078) <= not(layer1_outputs(6753)) or (layer1_outputs(931));
    layer2_outputs(5079) <= layer1_outputs(2662);
    layer2_outputs(5080) <= (layer1_outputs(1514)) or (layer1_outputs(4732));
    layer2_outputs(5081) <= layer1_outputs(338);
    layer2_outputs(5082) <= not(layer1_outputs(2636)) or (layer1_outputs(2269));
    layer2_outputs(5083) <= not((layer1_outputs(7215)) and (layer1_outputs(6555)));
    layer2_outputs(5084) <= layer1_outputs(268);
    layer2_outputs(5085) <= (layer1_outputs(715)) and not (layer1_outputs(2361));
    layer2_outputs(5086) <= not((layer1_outputs(4830)) or (layer1_outputs(6772)));
    layer2_outputs(5087) <= '1';
    layer2_outputs(5088) <= (layer1_outputs(5913)) or (layer1_outputs(1619));
    layer2_outputs(5089) <= not((layer1_outputs(3930)) and (layer1_outputs(5193)));
    layer2_outputs(5090) <= not((layer1_outputs(4123)) or (layer1_outputs(3527)));
    layer2_outputs(5091) <= (layer1_outputs(4077)) and not (layer1_outputs(1449));
    layer2_outputs(5092) <= '0';
    layer2_outputs(5093) <= '1';
    layer2_outputs(5094) <= not((layer1_outputs(4440)) or (layer1_outputs(1000)));
    layer2_outputs(5095) <= not(layer1_outputs(1083));
    layer2_outputs(5096) <= not(layer1_outputs(1343));
    layer2_outputs(5097) <= '0';
    layer2_outputs(5098) <= (layer1_outputs(2536)) or (layer1_outputs(1795));
    layer2_outputs(5099) <= layer1_outputs(826);
    layer2_outputs(5100) <= layer1_outputs(4950);
    layer2_outputs(5101) <= not(layer1_outputs(7296)) or (layer1_outputs(5438));
    layer2_outputs(5102) <= (layer1_outputs(5819)) or (layer1_outputs(2672));
    layer2_outputs(5103) <= (layer1_outputs(5568)) and not (layer1_outputs(6080));
    layer2_outputs(5104) <= '0';
    layer2_outputs(5105) <= (layer1_outputs(7534)) and (layer1_outputs(6962));
    layer2_outputs(5106) <= not(layer1_outputs(2629));
    layer2_outputs(5107) <= (layer1_outputs(6378)) and not (layer1_outputs(6607));
    layer2_outputs(5108) <= not(layer1_outputs(2902));
    layer2_outputs(5109) <= (layer1_outputs(7197)) and (layer1_outputs(3680));
    layer2_outputs(5110) <= layer1_outputs(4528);
    layer2_outputs(5111) <= (layer1_outputs(2564)) and not (layer1_outputs(7235));
    layer2_outputs(5112) <= not(layer1_outputs(1265)) or (layer1_outputs(1630));
    layer2_outputs(5113) <= not(layer1_outputs(447));
    layer2_outputs(5114) <= not(layer1_outputs(2504));
    layer2_outputs(5115) <= not((layer1_outputs(2500)) and (layer1_outputs(175)));
    layer2_outputs(5116) <= '0';
    layer2_outputs(5117) <= '1';
    layer2_outputs(5118) <= (layer1_outputs(5750)) and not (layer1_outputs(425));
    layer2_outputs(5119) <= not(layer1_outputs(384));
    layer2_outputs(5120) <= layer1_outputs(4894);
    layer2_outputs(5121) <= not((layer1_outputs(148)) and (layer1_outputs(554)));
    layer2_outputs(5122) <= not((layer1_outputs(4659)) or (layer1_outputs(5963)));
    layer2_outputs(5123) <= not(layer1_outputs(1607));
    layer2_outputs(5124) <= not((layer1_outputs(1601)) or (layer1_outputs(5573)));
    layer2_outputs(5125) <= (layer1_outputs(4070)) and (layer1_outputs(916));
    layer2_outputs(5126) <= not(layer1_outputs(5111)) or (layer1_outputs(3913));
    layer2_outputs(5127) <= not(layer1_outputs(7524)) or (layer1_outputs(2320));
    layer2_outputs(5128) <= (layer1_outputs(121)) or (layer1_outputs(1893));
    layer2_outputs(5129) <= not(layer1_outputs(376));
    layer2_outputs(5130) <= not(layer1_outputs(1075)) or (layer1_outputs(1884));
    layer2_outputs(5131) <= not(layer1_outputs(4366)) or (layer1_outputs(5603));
    layer2_outputs(5132) <= (layer1_outputs(845)) or (layer1_outputs(3348));
    layer2_outputs(5133) <= (layer1_outputs(484)) and not (layer1_outputs(4843));
    layer2_outputs(5134) <= not((layer1_outputs(4141)) and (layer1_outputs(6756)));
    layer2_outputs(5135) <= '1';
    layer2_outputs(5136) <= not(layer1_outputs(3479));
    layer2_outputs(5137) <= (layer1_outputs(1073)) or (layer1_outputs(4519));
    layer2_outputs(5138) <= layer1_outputs(7650);
    layer2_outputs(5139) <= '1';
    layer2_outputs(5140) <= (layer1_outputs(6068)) and not (layer1_outputs(1644));
    layer2_outputs(5141) <= '0';
    layer2_outputs(5142) <= not(layer1_outputs(5364));
    layer2_outputs(5143) <= (layer1_outputs(1104)) and not (layer1_outputs(608));
    layer2_outputs(5144) <= not(layer1_outputs(3933)) or (layer1_outputs(5322));
    layer2_outputs(5145) <= (layer1_outputs(552)) and not (layer1_outputs(5219));
    layer2_outputs(5146) <= not((layer1_outputs(5045)) or (layer1_outputs(3802)));
    layer2_outputs(5147) <= (layer1_outputs(6151)) or (layer1_outputs(6626));
    layer2_outputs(5148) <= (layer1_outputs(357)) or (layer1_outputs(4753));
    layer2_outputs(5149) <= (layer1_outputs(86)) and not (layer1_outputs(415));
    layer2_outputs(5150) <= layer1_outputs(5800);
    layer2_outputs(5151) <= layer1_outputs(740);
    layer2_outputs(5152) <= (layer1_outputs(5146)) or (layer1_outputs(5445));
    layer2_outputs(5153) <= not((layer1_outputs(5912)) and (layer1_outputs(4669)));
    layer2_outputs(5154) <= not((layer1_outputs(6135)) or (layer1_outputs(4854)));
    layer2_outputs(5155) <= (layer1_outputs(3666)) and not (layer1_outputs(856));
    layer2_outputs(5156) <= not(layer1_outputs(5850)) or (layer1_outputs(5741));
    layer2_outputs(5157) <= layer1_outputs(1169);
    layer2_outputs(5158) <= layer1_outputs(638);
    layer2_outputs(5159) <= layer1_outputs(2358);
    layer2_outputs(5160) <= layer1_outputs(258);
    layer2_outputs(5161) <= (layer1_outputs(3285)) and (layer1_outputs(7414));
    layer2_outputs(5162) <= '1';
    layer2_outputs(5163) <= not(layer1_outputs(4055));
    layer2_outputs(5164) <= not((layer1_outputs(4944)) or (layer1_outputs(5493)));
    layer2_outputs(5165) <= layer1_outputs(2941);
    layer2_outputs(5166) <= '1';
    layer2_outputs(5167) <= not((layer1_outputs(5844)) and (layer1_outputs(1058)));
    layer2_outputs(5168) <= not(layer1_outputs(2580));
    layer2_outputs(5169) <= (layer1_outputs(6730)) or (layer1_outputs(7666));
    layer2_outputs(5170) <= '1';
    layer2_outputs(5171) <= (layer1_outputs(3760)) and not (layer1_outputs(505));
    layer2_outputs(5172) <= '1';
    layer2_outputs(5173) <= '1';
    layer2_outputs(5174) <= not(layer1_outputs(4704));
    layer2_outputs(5175) <= '0';
    layer2_outputs(5176) <= '1';
    layer2_outputs(5177) <= not(layer1_outputs(4975));
    layer2_outputs(5178) <= layer1_outputs(4022);
    layer2_outputs(5179) <= '0';
    layer2_outputs(5180) <= layer1_outputs(3052);
    layer2_outputs(5181) <= not(layer1_outputs(4836)) or (layer1_outputs(5661));
    layer2_outputs(5182) <= not((layer1_outputs(7305)) or (layer1_outputs(4407)));
    layer2_outputs(5183) <= layer1_outputs(2084);
    layer2_outputs(5184) <= '0';
    layer2_outputs(5185) <= layer1_outputs(5212);
    layer2_outputs(5186) <= not(layer1_outputs(6478));
    layer2_outputs(5187) <= '0';
    layer2_outputs(5188) <= not(layer1_outputs(816));
    layer2_outputs(5189) <= layer1_outputs(6156);
    layer2_outputs(5190) <= not(layer1_outputs(7634));
    layer2_outputs(5191) <= not(layer1_outputs(4744)) or (layer1_outputs(3397));
    layer2_outputs(5192) <= not(layer1_outputs(4738));
    layer2_outputs(5193) <= '1';
    layer2_outputs(5194) <= not(layer1_outputs(6549));
    layer2_outputs(5195) <= layer1_outputs(2503);
    layer2_outputs(5196) <= (layer1_outputs(7551)) or (layer1_outputs(4761));
    layer2_outputs(5197) <= not(layer1_outputs(5655)) or (layer1_outputs(4982));
    layer2_outputs(5198) <= not((layer1_outputs(3260)) and (layer1_outputs(6010)));
    layer2_outputs(5199) <= (layer1_outputs(221)) or (layer1_outputs(5886));
    layer2_outputs(5200) <= not((layer1_outputs(6767)) and (layer1_outputs(2606)));
    layer2_outputs(5201) <= (layer1_outputs(2758)) and not (layer1_outputs(633));
    layer2_outputs(5202) <= (layer1_outputs(3890)) and not (layer1_outputs(1413));
    layer2_outputs(5203) <= not(layer1_outputs(3781)) or (layer1_outputs(1414));
    layer2_outputs(5204) <= (layer1_outputs(7354)) or (layer1_outputs(1788));
    layer2_outputs(5205) <= (layer1_outputs(5830)) and not (layer1_outputs(5591));
    layer2_outputs(5206) <= '0';
    layer2_outputs(5207) <= not(layer1_outputs(1955)) or (layer1_outputs(1843));
    layer2_outputs(5208) <= (layer1_outputs(17)) and not (layer1_outputs(5462));
    layer2_outputs(5209) <= layer1_outputs(2866);
    layer2_outputs(5210) <= not(layer1_outputs(7464)) or (layer1_outputs(1262));
    layer2_outputs(5211) <= layer1_outputs(1677);
    layer2_outputs(5212) <= not(layer1_outputs(1885));
    layer2_outputs(5213) <= (layer1_outputs(6922)) and not (layer1_outputs(5924));
    layer2_outputs(5214) <= '1';
    layer2_outputs(5215) <= (layer1_outputs(336)) and not (layer1_outputs(4772));
    layer2_outputs(5216) <= layer1_outputs(316);
    layer2_outputs(5217) <= (layer1_outputs(2037)) and (layer1_outputs(3922));
    layer2_outputs(5218) <= '1';
    layer2_outputs(5219) <= (layer1_outputs(4444)) and (layer1_outputs(1456));
    layer2_outputs(5220) <= not(layer1_outputs(6696)) or (layer1_outputs(4102));
    layer2_outputs(5221) <= (layer1_outputs(3911)) and not (layer1_outputs(1074));
    layer2_outputs(5222) <= '1';
    layer2_outputs(5223) <= not(layer1_outputs(2938));
    layer2_outputs(5224) <= layer1_outputs(2748);
    layer2_outputs(5225) <= (layer1_outputs(6514)) and (layer1_outputs(2285));
    layer2_outputs(5226) <= layer1_outputs(4886);
    layer2_outputs(5227) <= not((layer1_outputs(2536)) and (layer1_outputs(381)));
    layer2_outputs(5228) <= '1';
    layer2_outputs(5229) <= not((layer1_outputs(5583)) or (layer1_outputs(3797)));
    layer2_outputs(5230) <= not(layer1_outputs(2549));
    layer2_outputs(5231) <= not(layer1_outputs(5283));
    layer2_outputs(5232) <= layer1_outputs(2397);
    layer2_outputs(5233) <= layer1_outputs(2455);
    layer2_outputs(5234) <= not(layer1_outputs(7224)) or (layer1_outputs(6029));
    layer2_outputs(5235) <= layer1_outputs(5260);
    layer2_outputs(5236) <= (layer1_outputs(1605)) or (layer1_outputs(3627));
    layer2_outputs(5237) <= not(layer1_outputs(4363)) or (layer1_outputs(570));
    layer2_outputs(5238) <= not(layer1_outputs(2677)) or (layer1_outputs(5861));
    layer2_outputs(5239) <= layer1_outputs(1116);
    layer2_outputs(5240) <= layer1_outputs(7621);
    layer2_outputs(5241) <= not((layer1_outputs(274)) and (layer1_outputs(3918)));
    layer2_outputs(5242) <= (layer1_outputs(6570)) and (layer1_outputs(4393));
    layer2_outputs(5243) <= not(layer1_outputs(5317)) or (layer1_outputs(7183));
    layer2_outputs(5244) <= not(layer1_outputs(4390));
    layer2_outputs(5245) <= '1';
    layer2_outputs(5246) <= not(layer1_outputs(6588));
    layer2_outputs(5247) <= (layer1_outputs(5085)) and not (layer1_outputs(7412));
    layer2_outputs(5248) <= (layer1_outputs(4786)) and not (layer1_outputs(1898));
    layer2_outputs(5249) <= not(layer1_outputs(6994)) or (layer1_outputs(2012));
    layer2_outputs(5250) <= layer1_outputs(406);
    layer2_outputs(5251) <= layer1_outputs(6368);
    layer2_outputs(5252) <= layer1_outputs(4898);
    layer2_outputs(5253) <= (layer1_outputs(3627)) and (layer1_outputs(1094));
    layer2_outputs(5254) <= layer1_outputs(7298);
    layer2_outputs(5255) <= not(layer1_outputs(3376));
    layer2_outputs(5256) <= not((layer1_outputs(5268)) and (layer1_outputs(4535)));
    layer2_outputs(5257) <= not(layer1_outputs(5266)) or (layer1_outputs(5536));
    layer2_outputs(5258) <= not(layer1_outputs(4240));
    layer2_outputs(5259) <= layer1_outputs(186);
    layer2_outputs(5260) <= (layer1_outputs(5243)) and not (layer1_outputs(6890));
    layer2_outputs(5261) <= (layer1_outputs(1455)) and not (layer1_outputs(3305));
    layer2_outputs(5262) <= not(layer1_outputs(4068));
    layer2_outputs(5263) <= not(layer1_outputs(5352));
    layer2_outputs(5264) <= (layer1_outputs(6105)) and not (layer1_outputs(4621));
    layer2_outputs(5265) <= (layer1_outputs(364)) and not (layer1_outputs(2016));
    layer2_outputs(5266) <= not((layer1_outputs(3825)) and (layer1_outputs(3443)));
    layer2_outputs(5267) <= not(layer1_outputs(6968)) or (layer1_outputs(6482));
    layer2_outputs(5268) <= layer1_outputs(3068);
    layer2_outputs(5269) <= (layer1_outputs(6787)) and not (layer1_outputs(400));
    layer2_outputs(5270) <= (layer1_outputs(5220)) and not (layer1_outputs(382));
    layer2_outputs(5271) <= not(layer1_outputs(1917)) or (layer1_outputs(4094));
    layer2_outputs(5272) <= not(layer1_outputs(770));
    layer2_outputs(5273) <= not(layer1_outputs(4260)) or (layer1_outputs(3683));
    layer2_outputs(5274) <= (layer1_outputs(1904)) and (layer1_outputs(4210));
    layer2_outputs(5275) <= layer1_outputs(3296);
    layer2_outputs(5276) <= not(layer1_outputs(2773));
    layer2_outputs(5277) <= (layer1_outputs(6319)) and (layer1_outputs(3915));
    layer2_outputs(5278) <= '1';
    layer2_outputs(5279) <= layer1_outputs(5556);
    layer2_outputs(5280) <= not(layer1_outputs(7265)) or (layer1_outputs(1045));
    layer2_outputs(5281) <= '1';
    layer2_outputs(5282) <= (layer1_outputs(7367)) or (layer1_outputs(3339));
    layer2_outputs(5283) <= not(layer1_outputs(6713));
    layer2_outputs(5284) <= not((layer1_outputs(3835)) or (layer1_outputs(4108)));
    layer2_outputs(5285) <= (layer1_outputs(3309)) and not (layer1_outputs(132));
    layer2_outputs(5286) <= not(layer1_outputs(3625));
    layer2_outputs(5287) <= (layer1_outputs(3382)) and (layer1_outputs(3230));
    layer2_outputs(5288) <= not(layer1_outputs(2455));
    layer2_outputs(5289) <= layer1_outputs(5775);
    layer2_outputs(5290) <= (layer1_outputs(1513)) and not (layer1_outputs(743));
    layer2_outputs(5291) <= (layer1_outputs(1747)) or (layer1_outputs(3333));
    layer2_outputs(5292) <= '1';
    layer2_outputs(5293) <= (layer1_outputs(2024)) or (layer1_outputs(4162));
    layer2_outputs(5294) <= not(layer1_outputs(4817));
    layer2_outputs(5295) <= not(layer1_outputs(583));
    layer2_outputs(5296) <= not(layer1_outputs(6372)) or (layer1_outputs(3199));
    layer2_outputs(5297) <= '1';
    layer2_outputs(5298) <= not((layer1_outputs(342)) or (layer1_outputs(6049)));
    layer2_outputs(5299) <= layer1_outputs(1547);
    layer2_outputs(5300) <= layer1_outputs(1668);
    layer2_outputs(5301) <= (layer1_outputs(933)) and (layer1_outputs(7057));
    layer2_outputs(5302) <= (layer1_outputs(2722)) and not (layer1_outputs(4915));
    layer2_outputs(5303) <= not((layer1_outputs(5258)) or (layer1_outputs(2193)));
    layer2_outputs(5304) <= '1';
    layer2_outputs(5305) <= '1';
    layer2_outputs(5306) <= '1';
    layer2_outputs(5307) <= layer1_outputs(4264);
    layer2_outputs(5308) <= layer1_outputs(2210);
    layer2_outputs(5309) <= layer1_outputs(5062);
    layer2_outputs(5310) <= not(layer1_outputs(3304)) or (layer1_outputs(6583));
    layer2_outputs(5311) <= '1';
    layer2_outputs(5312) <= not(layer1_outputs(4134));
    layer2_outputs(5313) <= not(layer1_outputs(6957)) or (layer1_outputs(1279));
    layer2_outputs(5314) <= '0';
    layer2_outputs(5315) <= '0';
    layer2_outputs(5316) <= layer1_outputs(3578);
    layer2_outputs(5317) <= layer1_outputs(5955);
    layer2_outputs(5318) <= not(layer1_outputs(6644));
    layer2_outputs(5319) <= layer1_outputs(3086);
    layer2_outputs(5320) <= not(layer1_outputs(3951));
    layer2_outputs(5321) <= not(layer1_outputs(96));
    layer2_outputs(5322) <= not((layer1_outputs(5341)) and (layer1_outputs(7535)));
    layer2_outputs(5323) <= (layer1_outputs(5719)) or (layer1_outputs(5930));
    layer2_outputs(5324) <= not(layer1_outputs(4946));
    layer2_outputs(5325) <= not((layer1_outputs(1872)) or (layer1_outputs(6818)));
    layer2_outputs(5326) <= '0';
    layer2_outputs(5327) <= '1';
    layer2_outputs(5328) <= (layer1_outputs(1254)) and not (layer1_outputs(2019));
    layer2_outputs(5329) <= layer1_outputs(99);
    layer2_outputs(5330) <= not((layer1_outputs(565)) or (layer1_outputs(5755)));
    layer2_outputs(5331) <= not(layer1_outputs(1416)) or (layer1_outputs(6698));
    layer2_outputs(5332) <= (layer1_outputs(7103)) and not (layer1_outputs(1209));
    layer2_outputs(5333) <= (layer1_outputs(5525)) and (layer1_outputs(3317));
    layer2_outputs(5334) <= '0';
    layer2_outputs(5335) <= not(layer1_outputs(470)) or (layer1_outputs(7633));
    layer2_outputs(5336) <= not((layer1_outputs(7587)) or (layer1_outputs(1295)));
    layer2_outputs(5337) <= '1';
    layer2_outputs(5338) <= not(layer1_outputs(5510));
    layer2_outputs(5339) <= (layer1_outputs(2322)) or (layer1_outputs(1096));
    layer2_outputs(5340) <= (layer1_outputs(1785)) or (layer1_outputs(5859));
    layer2_outputs(5341) <= (layer1_outputs(6817)) and not (layer1_outputs(4796));
    layer2_outputs(5342) <= layer1_outputs(1606);
    layer2_outputs(5343) <= '0';
    layer2_outputs(5344) <= (layer1_outputs(2434)) xor (layer1_outputs(4224));
    layer2_outputs(5345) <= '1';
    layer2_outputs(5346) <= layer1_outputs(7357);
    layer2_outputs(5347) <= layer1_outputs(5304);
    layer2_outputs(5348) <= (layer1_outputs(4610)) or (layer1_outputs(2020));
    layer2_outputs(5349) <= not(layer1_outputs(5552)) or (layer1_outputs(4891));
    layer2_outputs(5350) <= layer1_outputs(7280);
    layer2_outputs(5351) <= not(layer1_outputs(3166)) or (layer1_outputs(736));
    layer2_outputs(5352) <= not(layer1_outputs(1624));
    layer2_outputs(5353) <= '1';
    layer2_outputs(5354) <= layer1_outputs(273);
    layer2_outputs(5355) <= not((layer1_outputs(6634)) and (layer1_outputs(2621)));
    layer2_outputs(5356) <= (layer1_outputs(5428)) and (layer1_outputs(1114));
    layer2_outputs(5357) <= (layer1_outputs(7279)) and not (layer1_outputs(1954));
    layer2_outputs(5358) <= layer1_outputs(102);
    layer2_outputs(5359) <= not(layer1_outputs(2440));
    layer2_outputs(5360) <= '1';
    layer2_outputs(5361) <= not((layer1_outputs(4163)) xor (layer1_outputs(1582)));
    layer2_outputs(5362) <= not((layer1_outputs(2341)) and (layer1_outputs(1650)));
    layer2_outputs(5363) <= layer1_outputs(6210);
    layer2_outputs(5364) <= not((layer1_outputs(4486)) or (layer1_outputs(174)));
    layer2_outputs(5365) <= (layer1_outputs(7281)) and not (layer1_outputs(3898));
    layer2_outputs(5366) <= layer1_outputs(1950);
    layer2_outputs(5367) <= '0';
    layer2_outputs(5368) <= not(layer1_outputs(3751));
    layer2_outputs(5369) <= '1';
    layer2_outputs(5370) <= '1';
    layer2_outputs(5371) <= (layer1_outputs(6916)) or (layer1_outputs(5225));
    layer2_outputs(5372) <= '1';
    layer2_outputs(5373) <= layer1_outputs(7003);
    layer2_outputs(5374) <= not(layer1_outputs(871));
    layer2_outputs(5375) <= '0';
    layer2_outputs(5376) <= (layer1_outputs(6586)) and not (layer1_outputs(3038));
    layer2_outputs(5377) <= not(layer1_outputs(7519));
    layer2_outputs(5378) <= layer1_outputs(4251);
    layer2_outputs(5379) <= not((layer1_outputs(5378)) or (layer1_outputs(3489)));
    layer2_outputs(5380) <= not(layer1_outputs(2307));
    layer2_outputs(5381) <= not((layer1_outputs(548)) and (layer1_outputs(4252)));
    layer2_outputs(5382) <= layer1_outputs(5120);
    layer2_outputs(5383) <= (layer1_outputs(4980)) and not (layer1_outputs(3042));
    layer2_outputs(5384) <= (layer1_outputs(7059)) and (layer1_outputs(4925));
    layer2_outputs(5385) <= not(layer1_outputs(6939));
    layer2_outputs(5386) <= layer1_outputs(6433);
    layer2_outputs(5387) <= (layer1_outputs(2130)) or (layer1_outputs(3601));
    layer2_outputs(5388) <= not((layer1_outputs(4566)) or (layer1_outputs(1802)));
    layer2_outputs(5389) <= '0';
    layer2_outputs(5390) <= (layer1_outputs(3059)) and (layer1_outputs(1365));
    layer2_outputs(5391) <= (layer1_outputs(3599)) and (layer1_outputs(900));
    layer2_outputs(5392) <= (layer1_outputs(951)) and (layer1_outputs(6509));
    layer2_outputs(5393) <= not(layer1_outputs(3322));
    layer2_outputs(5394) <= (layer1_outputs(1488)) and not (layer1_outputs(571));
    layer2_outputs(5395) <= '1';
    layer2_outputs(5396) <= (layer1_outputs(5173)) and not (layer1_outputs(7602));
    layer2_outputs(5397) <= not(layer1_outputs(6876)) or (layer1_outputs(3068));
    layer2_outputs(5398) <= layer1_outputs(1232);
    layer2_outputs(5399) <= (layer1_outputs(6564)) or (layer1_outputs(6741));
    layer2_outputs(5400) <= (layer1_outputs(3817)) and not (layer1_outputs(3475));
    layer2_outputs(5401) <= not((layer1_outputs(6164)) and (layer1_outputs(3344)));
    layer2_outputs(5402) <= not((layer1_outputs(6222)) and (layer1_outputs(2852)));
    layer2_outputs(5403) <= not(layer1_outputs(5593)) or (layer1_outputs(6749));
    layer2_outputs(5404) <= not((layer1_outputs(5061)) or (layer1_outputs(3588)));
    layer2_outputs(5405) <= not((layer1_outputs(3829)) or (layer1_outputs(4470)));
    layer2_outputs(5406) <= not(layer1_outputs(3433)) or (layer1_outputs(6511));
    layer2_outputs(5407) <= not(layer1_outputs(3918)) or (layer1_outputs(6440));
    layer2_outputs(5408) <= not(layer1_outputs(3586));
    layer2_outputs(5409) <= '1';
    layer2_outputs(5410) <= '1';
    layer2_outputs(5411) <= (layer1_outputs(1679)) and not (layer1_outputs(6911));
    layer2_outputs(5412) <= not(layer1_outputs(157)) or (layer1_outputs(158));
    layer2_outputs(5413) <= (layer1_outputs(5349)) or (layer1_outputs(4806));
    layer2_outputs(5414) <= not(layer1_outputs(4466));
    layer2_outputs(5415) <= not(layer1_outputs(2347)) or (layer1_outputs(2077));
    layer2_outputs(5416) <= '0';
    layer2_outputs(5417) <= layer1_outputs(3039);
    layer2_outputs(5418) <= not(layer1_outputs(5532)) or (layer1_outputs(5773));
    layer2_outputs(5419) <= not(layer1_outputs(30));
    layer2_outputs(5420) <= not((layer1_outputs(7469)) xor (layer1_outputs(3978)));
    layer2_outputs(5421) <= (layer1_outputs(1335)) and not (layer1_outputs(5313));
    layer2_outputs(5422) <= not(layer1_outputs(3705)) or (layer1_outputs(1487));
    layer2_outputs(5423) <= not((layer1_outputs(6527)) or (layer1_outputs(7090)));
    layer2_outputs(5424) <= not((layer1_outputs(1648)) and (layer1_outputs(5635)));
    layer2_outputs(5425) <= '0';
    layer2_outputs(5426) <= not((layer1_outputs(1346)) or (layer1_outputs(597)));
    layer2_outputs(5427) <= layer1_outputs(4370);
    layer2_outputs(5428) <= layer1_outputs(3943);
    layer2_outputs(5429) <= not(layer1_outputs(3085)) or (layer1_outputs(3861));
    layer2_outputs(5430) <= '0';
    layer2_outputs(5431) <= layer1_outputs(6510);
    layer2_outputs(5432) <= not(layer1_outputs(6897)) or (layer1_outputs(2450));
    layer2_outputs(5433) <= not(layer1_outputs(6437)) or (layer1_outputs(6073));
    layer2_outputs(5434) <= not((layer1_outputs(1835)) and (layer1_outputs(4254)));
    layer2_outputs(5435) <= not(layer1_outputs(3));
    layer2_outputs(5436) <= '1';
    layer2_outputs(5437) <= (layer1_outputs(1969)) and (layer1_outputs(4304));
    layer2_outputs(5438) <= '0';
    layer2_outputs(5439) <= not(layer1_outputs(391));
    layer2_outputs(5440) <= '0';
    layer2_outputs(5441) <= not(layer1_outputs(4411)) or (layer1_outputs(3942));
    layer2_outputs(5442) <= not(layer1_outputs(1970));
    layer2_outputs(5443) <= layer1_outputs(4394);
    layer2_outputs(5444) <= not(layer1_outputs(6354)) or (layer1_outputs(2400));
    layer2_outputs(5445) <= not(layer1_outputs(3158));
    layer2_outputs(5446) <= not(layer1_outputs(6200)) or (layer1_outputs(1126));
    layer2_outputs(5447) <= not(layer1_outputs(513)) or (layer1_outputs(1998));
    layer2_outputs(5448) <= not(layer1_outputs(3252)) or (layer1_outputs(4682));
    layer2_outputs(5449) <= (layer1_outputs(1066)) and not (layer1_outputs(5599));
    layer2_outputs(5450) <= not((layer1_outputs(2401)) or (layer1_outputs(4701)));
    layer2_outputs(5451) <= not(layer1_outputs(7585));
    layer2_outputs(5452) <= not(layer1_outputs(5823)) or (layer1_outputs(6524));
    layer2_outputs(5453) <= layer1_outputs(2163);
    layer2_outputs(5454) <= not((layer1_outputs(591)) or (layer1_outputs(3334)));
    layer2_outputs(5455) <= layer1_outputs(4288);
    layer2_outputs(5456) <= not(layer1_outputs(6016));
    layer2_outputs(5457) <= not(layer1_outputs(1366)) or (layer1_outputs(2814));
    layer2_outputs(5458) <= '1';
    layer2_outputs(5459) <= '1';
    layer2_outputs(5460) <= not(layer1_outputs(4345)) or (layer1_outputs(6442));
    layer2_outputs(5461) <= (layer1_outputs(6277)) or (layer1_outputs(1100));
    layer2_outputs(5462) <= not(layer1_outputs(6329));
    layer2_outputs(5463) <= layer1_outputs(5385);
    layer2_outputs(5464) <= not(layer1_outputs(2306));
    layer2_outputs(5465) <= not(layer1_outputs(2190)) or (layer1_outputs(4823));
    layer2_outputs(5466) <= not((layer1_outputs(2202)) xor (layer1_outputs(3300)));
    layer2_outputs(5467) <= not(layer1_outputs(3095)) or (layer1_outputs(6840));
    layer2_outputs(5468) <= layer1_outputs(5060);
    layer2_outputs(5469) <= (layer1_outputs(1160)) or (layer1_outputs(7446));
    layer2_outputs(5470) <= (layer1_outputs(4293)) and not (layer1_outputs(5612));
    layer2_outputs(5471) <= not((layer1_outputs(7522)) or (layer1_outputs(5554)));
    layer2_outputs(5472) <= layer1_outputs(7131);
    layer2_outputs(5473) <= layer1_outputs(5838);
    layer2_outputs(5474) <= not((layer1_outputs(6467)) and (layer1_outputs(4617)));
    layer2_outputs(5475) <= not(layer1_outputs(43)) or (layer1_outputs(2836));
    layer2_outputs(5476) <= not(layer1_outputs(446));
    layer2_outputs(5477) <= not(layer1_outputs(1007)) or (layer1_outputs(1130));
    layer2_outputs(5478) <= not(layer1_outputs(6077));
    layer2_outputs(5479) <= layer1_outputs(7214);
    layer2_outputs(5480) <= (layer1_outputs(1877)) and (layer1_outputs(1662));
    layer2_outputs(5481) <= (layer1_outputs(418)) and (layer1_outputs(4229));
    layer2_outputs(5482) <= (layer1_outputs(4287)) and not (layer1_outputs(922));
    layer2_outputs(5483) <= '1';
    layer2_outputs(5484) <= not((layer1_outputs(6397)) and (layer1_outputs(6660)));
    layer2_outputs(5485) <= (layer1_outputs(1066)) and not (layer1_outputs(4333));
    layer2_outputs(5486) <= not(layer1_outputs(6868));
    layer2_outputs(5487) <= '0';
    layer2_outputs(5488) <= not((layer1_outputs(5095)) and (layer1_outputs(3658)));
    layer2_outputs(5489) <= '0';
    layer2_outputs(5490) <= layer1_outputs(6890);
    layer2_outputs(5491) <= not(layer1_outputs(7612)) or (layer1_outputs(875));
    layer2_outputs(5492) <= not((layer1_outputs(5287)) and (layer1_outputs(3317)));
    layer2_outputs(5493) <= not(layer1_outputs(6952));
    layer2_outputs(5494) <= '1';
    layer2_outputs(5495) <= '1';
    layer2_outputs(5496) <= '0';
    layer2_outputs(5497) <= not((layer1_outputs(287)) or (layer1_outputs(1675)));
    layer2_outputs(5498) <= not(layer1_outputs(1569)) or (layer1_outputs(898));
    layer2_outputs(5499) <= (layer1_outputs(2170)) and not (layer1_outputs(3223));
    layer2_outputs(5500) <= not((layer1_outputs(1303)) and (layer1_outputs(2196)));
    layer2_outputs(5501) <= not((layer1_outputs(7486)) or (layer1_outputs(6860)));
    layer2_outputs(5502) <= '1';
    layer2_outputs(5503) <= not(layer1_outputs(5488));
    layer2_outputs(5504) <= not(layer1_outputs(1301)) or (layer1_outputs(2063));
    layer2_outputs(5505) <= '0';
    layer2_outputs(5506) <= (layer1_outputs(3465)) or (layer1_outputs(2735));
    layer2_outputs(5507) <= '1';
    layer2_outputs(5508) <= not(layer1_outputs(6472)) or (layer1_outputs(401));
    layer2_outputs(5509) <= '0';
    layer2_outputs(5510) <= layer1_outputs(3813);
    layer2_outputs(5511) <= (layer1_outputs(482)) and not (layer1_outputs(1857));
    layer2_outputs(5512) <= (layer1_outputs(6452)) or (layer1_outputs(7315));
    layer2_outputs(5513) <= not(layer1_outputs(1121)) or (layer1_outputs(5103));
    layer2_outputs(5514) <= (layer1_outputs(857)) or (layer1_outputs(6158));
    layer2_outputs(5515) <= (layer1_outputs(1391)) and not (layer1_outputs(2935));
    layer2_outputs(5516) <= layer1_outputs(4625);
    layer2_outputs(5517) <= not(layer1_outputs(4744)) or (layer1_outputs(7465));
    layer2_outputs(5518) <= (layer1_outputs(7218)) and not (layer1_outputs(3865));
    layer2_outputs(5519) <= '0';
    layer2_outputs(5520) <= not((layer1_outputs(5430)) or (layer1_outputs(6658)));
    layer2_outputs(5521) <= '1';
    layer2_outputs(5522) <= (layer1_outputs(314)) and not (layer1_outputs(916));
    layer2_outputs(5523) <= '0';
    layer2_outputs(5524) <= layer1_outputs(1475);
    layer2_outputs(5525) <= '1';
    layer2_outputs(5526) <= not(layer1_outputs(5818));
    layer2_outputs(5527) <= not((layer1_outputs(5519)) or (layer1_outputs(4099)));
    layer2_outputs(5528) <= layer1_outputs(5238);
    layer2_outputs(5529) <= not((layer1_outputs(5719)) and (layer1_outputs(5078)));
    layer2_outputs(5530) <= not(layer1_outputs(967));
    layer2_outputs(5531) <= not((layer1_outputs(6130)) or (layer1_outputs(3350)));
    layer2_outputs(5532) <= not(layer1_outputs(1987));
    layer2_outputs(5533) <= '1';
    layer2_outputs(5534) <= layer1_outputs(7507);
    layer2_outputs(5535) <= '0';
    layer2_outputs(5536) <= (layer1_outputs(5647)) and not (layer1_outputs(92));
    layer2_outputs(5537) <= '0';
    layer2_outputs(5538) <= not(layer1_outputs(5546));
    layer2_outputs(5539) <= '0';
    layer2_outputs(5540) <= '1';
    layer2_outputs(5541) <= '0';
    layer2_outputs(5542) <= not((layer1_outputs(1179)) or (layer1_outputs(416)));
    layer2_outputs(5543) <= (layer1_outputs(5302)) and (layer1_outputs(5161));
    layer2_outputs(5544) <= not(layer1_outputs(1932));
    layer2_outputs(5545) <= '1';
    layer2_outputs(5546) <= '0';
    layer2_outputs(5547) <= '1';
    layer2_outputs(5548) <= not(layer1_outputs(103)) or (layer1_outputs(5734));
    layer2_outputs(5549) <= layer1_outputs(1038);
    layer2_outputs(5550) <= (layer1_outputs(5039)) and not (layer1_outputs(2264));
    layer2_outputs(5551) <= (layer1_outputs(203)) and not (layer1_outputs(6191));
    layer2_outputs(5552) <= (layer1_outputs(6455)) and not (layer1_outputs(3451));
    layer2_outputs(5553) <= (layer1_outputs(3830)) and (layer1_outputs(4406));
    layer2_outputs(5554) <= not(layer1_outputs(177));
    layer2_outputs(5555) <= '0';
    layer2_outputs(5556) <= layer1_outputs(1261);
    layer2_outputs(5557) <= (layer1_outputs(4691)) and (layer1_outputs(4700));
    layer2_outputs(5558) <= (layer1_outputs(5153)) and (layer1_outputs(2609));
    layer2_outputs(5559) <= (layer1_outputs(2001)) xor (layer1_outputs(4788));
    layer2_outputs(5560) <= not(layer1_outputs(1746));
    layer2_outputs(5561) <= (layer1_outputs(5250)) or (layer1_outputs(6631));
    layer2_outputs(5562) <= not(layer1_outputs(2176));
    layer2_outputs(5563) <= not(layer1_outputs(979));
    layer2_outputs(5564) <= '1';
    layer2_outputs(5565) <= not(layer1_outputs(6357)) or (layer1_outputs(4651));
    layer2_outputs(5566) <= not(layer1_outputs(919)) or (layer1_outputs(1110));
    layer2_outputs(5567) <= not((layer1_outputs(3922)) or (layer1_outputs(1244)));
    layer2_outputs(5568) <= layer1_outputs(4168);
    layer2_outputs(5569) <= layer1_outputs(865);
    layer2_outputs(5570) <= not(layer1_outputs(4815));
    layer2_outputs(5571) <= layer1_outputs(1881);
    layer2_outputs(5572) <= not((layer1_outputs(4269)) and (layer1_outputs(1499)));
    layer2_outputs(5573) <= '0';
    layer2_outputs(5574) <= not(layer1_outputs(5100)) or (layer1_outputs(4748));
    layer2_outputs(5575) <= (layer1_outputs(7644)) xor (layer1_outputs(1639));
    layer2_outputs(5576) <= not((layer1_outputs(7353)) and (layer1_outputs(509)));
    layer2_outputs(5577) <= not(layer1_outputs(4841));
    layer2_outputs(5578) <= not(layer1_outputs(7614)) or (layer1_outputs(7157));
    layer2_outputs(5579) <= not(layer1_outputs(4435));
    layer2_outputs(5580) <= layer1_outputs(838);
    layer2_outputs(5581) <= not(layer1_outputs(517)) or (layer1_outputs(5236));
    layer2_outputs(5582) <= not((layer1_outputs(184)) or (layer1_outputs(2479)));
    layer2_outputs(5583) <= layer1_outputs(1673);
    layer2_outputs(5584) <= (layer1_outputs(3305)) xor (layer1_outputs(2739));
    layer2_outputs(5585) <= not(layer1_outputs(6134)) or (layer1_outputs(6045));
    layer2_outputs(5586) <= (layer1_outputs(5252)) and not (layer1_outputs(3544));
    layer2_outputs(5587) <= '1';
    layer2_outputs(5588) <= not(layer1_outputs(6972)) or (layer1_outputs(1805));
    layer2_outputs(5589) <= not(layer1_outputs(7019)) or (layer1_outputs(732));
    layer2_outputs(5590) <= layer1_outputs(72);
    layer2_outputs(5591) <= layer1_outputs(2109);
    layer2_outputs(5592) <= '1';
    layer2_outputs(5593) <= not(layer1_outputs(6672));
    layer2_outputs(5594) <= not((layer1_outputs(7496)) or (layer1_outputs(7598)));
    layer2_outputs(5595) <= not(layer1_outputs(3798));
    layer2_outputs(5596) <= not(layer1_outputs(795));
    layer2_outputs(5597) <= (layer1_outputs(3227)) xor (layer1_outputs(7354));
    layer2_outputs(5598) <= (layer1_outputs(1442)) and not (layer1_outputs(6274));
    layer2_outputs(5599) <= '1';
    layer2_outputs(5600) <= not((layer1_outputs(4977)) and (layer1_outputs(7304)));
    layer2_outputs(5601) <= layer1_outputs(3756);
    layer2_outputs(5602) <= (layer1_outputs(4427)) and (layer1_outputs(2765));
    layer2_outputs(5603) <= (layer1_outputs(7384)) and (layer1_outputs(2070));
    layer2_outputs(5604) <= (layer1_outputs(2172)) and not (layer1_outputs(1397));
    layer2_outputs(5605) <= (layer1_outputs(2683)) and (layer1_outputs(7634));
    layer2_outputs(5606) <= '0';
    layer2_outputs(5607) <= (layer1_outputs(6367)) and (layer1_outputs(114));
    layer2_outputs(5608) <= '1';
    layer2_outputs(5609) <= not((layer1_outputs(1448)) or (layer1_outputs(726)));
    layer2_outputs(5610) <= '1';
    layer2_outputs(5611) <= not(layer1_outputs(182));
    layer2_outputs(5612) <= not((layer1_outputs(53)) or (layer1_outputs(3091)));
    layer2_outputs(5613) <= (layer1_outputs(2150)) and (layer1_outputs(140));
    layer2_outputs(5614) <= not(layer1_outputs(5365)) or (layer1_outputs(2656));
    layer2_outputs(5615) <= layer1_outputs(2922);
    layer2_outputs(5616) <= not((layer1_outputs(5248)) or (layer1_outputs(5021)));
    layer2_outputs(5617) <= (layer1_outputs(6764)) and not (layer1_outputs(1422));
    layer2_outputs(5618) <= (layer1_outputs(3428)) and not (layer1_outputs(2236));
    layer2_outputs(5619) <= '0';
    layer2_outputs(5620) <= (layer1_outputs(3174)) and (layer1_outputs(5412));
    layer2_outputs(5621) <= (layer1_outputs(5218)) and not (layer1_outputs(7480));
    layer2_outputs(5622) <= '1';
    layer2_outputs(5623) <= not(layer1_outputs(640));
    layer2_outputs(5624) <= '1';
    layer2_outputs(5625) <= (layer1_outputs(942)) xor (layer1_outputs(1918));
    layer2_outputs(5626) <= (layer1_outputs(438)) or (layer1_outputs(2137));
    layer2_outputs(5627) <= '0';
    layer2_outputs(5628) <= not((layer1_outputs(907)) and (layer1_outputs(4465)));
    layer2_outputs(5629) <= not(layer1_outputs(2475)) or (layer1_outputs(3417));
    layer2_outputs(5630) <= (layer1_outputs(3161)) or (layer1_outputs(2618));
    layer2_outputs(5631) <= layer1_outputs(620);
    layer2_outputs(5632) <= not(layer1_outputs(2215)) or (layer1_outputs(6409));
    layer2_outputs(5633) <= layer1_outputs(4305);
    layer2_outputs(5634) <= layer1_outputs(6377);
    layer2_outputs(5635) <= layer1_outputs(2851);
    layer2_outputs(5636) <= not((layer1_outputs(4299)) xor (layer1_outputs(2652)));
    layer2_outputs(5637) <= '1';
    layer2_outputs(5638) <= not(layer1_outputs(4166)) or (layer1_outputs(3340));
    layer2_outputs(5639) <= (layer1_outputs(5632)) and (layer1_outputs(7562));
    layer2_outputs(5640) <= not((layer1_outputs(6512)) or (layer1_outputs(2205)));
    layer2_outputs(5641) <= not(layer1_outputs(117));
    layer2_outputs(5642) <= (layer1_outputs(7216)) and not (layer1_outputs(4257));
    layer2_outputs(5643) <= '1';
    layer2_outputs(5644) <= not(layer1_outputs(1943));
    layer2_outputs(5645) <= (layer1_outputs(5126)) and not (layer1_outputs(1768));
    layer2_outputs(5646) <= not(layer1_outputs(6376));
    layer2_outputs(5647) <= not(layer1_outputs(4015)) or (layer1_outputs(3019));
    layer2_outputs(5648) <= '0';
    layer2_outputs(5649) <= layer1_outputs(2072);
    layer2_outputs(5650) <= (layer1_outputs(4039)) and not (layer1_outputs(85));
    layer2_outputs(5651) <= (layer1_outputs(6513)) or (layer1_outputs(1897));
    layer2_outputs(5652) <= layer1_outputs(3594);
    layer2_outputs(5653) <= not((layer1_outputs(4316)) and (layer1_outputs(3618)));
    layer2_outputs(5654) <= layer1_outputs(5067);
    layer2_outputs(5655) <= not((layer1_outputs(6450)) or (layer1_outputs(974)));
    layer2_outputs(5656) <= not(layer1_outputs(6402));
    layer2_outputs(5657) <= not(layer1_outputs(7383));
    layer2_outputs(5658) <= layer1_outputs(2520);
    layer2_outputs(5659) <= layer1_outputs(5214);
    layer2_outputs(5660) <= (layer1_outputs(663)) and not (layer1_outputs(3511));
    layer2_outputs(5661) <= not(layer1_outputs(4087)) or (layer1_outputs(7492));
    layer2_outputs(5662) <= layer1_outputs(6808);
    layer2_outputs(5663) <= not(layer1_outputs(492));
    layer2_outputs(5664) <= (layer1_outputs(1214)) xor (layer1_outputs(5383));
    layer2_outputs(5665) <= '0';
    layer2_outputs(5666) <= layer1_outputs(5090);
    layer2_outputs(5667) <= (layer1_outputs(7644)) and not (layer1_outputs(6934));
    layer2_outputs(5668) <= not((layer1_outputs(3988)) or (layer1_outputs(3080)));
    layer2_outputs(5669) <= not(layer1_outputs(4675));
    layer2_outputs(5670) <= not((layer1_outputs(5938)) or (layer1_outputs(5973)));
    layer2_outputs(5671) <= (layer1_outputs(2913)) or (layer1_outputs(3757));
    layer2_outputs(5672) <= (layer1_outputs(689)) and (layer1_outputs(1516));
    layer2_outputs(5673) <= layer1_outputs(6436);
    layer2_outputs(5674) <= not((layer1_outputs(7302)) and (layer1_outputs(5702)));
    layer2_outputs(5675) <= '0';
    layer2_outputs(5676) <= not(layer1_outputs(1256)) or (layer1_outputs(7610));
    layer2_outputs(5677) <= not((layer1_outputs(1095)) and (layer1_outputs(5709)));
    layer2_outputs(5678) <= (layer1_outputs(6481)) and (layer1_outputs(1319));
    layer2_outputs(5679) <= (layer1_outputs(7355)) and (layer1_outputs(7264));
    layer2_outputs(5680) <= not((layer1_outputs(756)) and (layer1_outputs(3854)));
    layer2_outputs(5681) <= not((layer1_outputs(3950)) or (layer1_outputs(3311)));
    layer2_outputs(5682) <= (layer1_outputs(5035)) or (layer1_outputs(1195));
    layer2_outputs(5683) <= '0';
    layer2_outputs(5684) <= '1';
    layer2_outputs(5685) <= (layer1_outputs(6078)) and (layer1_outputs(6995));
    layer2_outputs(5686) <= not(layer1_outputs(5982));
    layer2_outputs(5687) <= '0';
    layer2_outputs(5688) <= (layer1_outputs(4909)) and not (layer1_outputs(1833));
    layer2_outputs(5689) <= not(layer1_outputs(4533));
    layer2_outputs(5690) <= '1';
    layer2_outputs(5691) <= not(layer1_outputs(4933)) or (layer1_outputs(7273));
    layer2_outputs(5692) <= not(layer1_outputs(3278));
    layer2_outputs(5693) <= not(layer1_outputs(2446)) or (layer1_outputs(2885));
    layer2_outputs(5694) <= not(layer1_outputs(6902));
    layer2_outputs(5695) <= layer1_outputs(7501);
    layer2_outputs(5696) <= (layer1_outputs(5598)) or (layer1_outputs(7063));
    layer2_outputs(5697) <= not((layer1_outputs(6881)) or (layer1_outputs(2005)));
    layer2_outputs(5698) <= not(layer1_outputs(1627)) or (layer1_outputs(4283));
    layer2_outputs(5699) <= layer1_outputs(2534);
    layer2_outputs(5700) <= not(layer1_outputs(5403));
    layer2_outputs(5701) <= not(layer1_outputs(7008)) or (layer1_outputs(2377));
    layer2_outputs(5702) <= (layer1_outputs(567)) and not (layer1_outputs(2778));
    layer2_outputs(5703) <= not((layer1_outputs(4716)) or (layer1_outputs(4498)));
    layer2_outputs(5704) <= layer1_outputs(4708);
    layer2_outputs(5705) <= '0';
    layer2_outputs(5706) <= not(layer1_outputs(6125)) or (layer1_outputs(285));
    layer2_outputs(5707) <= (layer1_outputs(6277)) and (layer1_outputs(778));
    layer2_outputs(5708) <= layer1_outputs(6959);
    layer2_outputs(5709) <= (layer1_outputs(2490)) xor (layer1_outputs(3543));
    layer2_outputs(5710) <= not((layer1_outputs(5675)) and (layer1_outputs(6681)));
    layer2_outputs(5711) <= '1';
    layer2_outputs(5712) <= not(layer1_outputs(2000));
    layer2_outputs(5713) <= not((layer1_outputs(5892)) or (layer1_outputs(874)));
    layer2_outputs(5714) <= layer1_outputs(2507);
    layer2_outputs(5715) <= (layer1_outputs(5620)) or (layer1_outputs(1597));
    layer2_outputs(5716) <= not(layer1_outputs(6656)) or (layer1_outputs(7543));
    layer2_outputs(5717) <= not(layer1_outputs(3746));
    layer2_outputs(5718) <= (layer1_outputs(6690)) and not (layer1_outputs(4949));
    layer2_outputs(5719) <= not((layer1_outputs(5572)) or (layer1_outputs(7065)));
    layer2_outputs(5720) <= not(layer1_outputs(2211));
    layer2_outputs(5721) <= not(layer1_outputs(6120)) or (layer1_outputs(7325));
    layer2_outputs(5722) <= '0';
    layer2_outputs(5723) <= (layer1_outputs(6545)) and not (layer1_outputs(4634));
    layer2_outputs(5724) <= not(layer1_outputs(1934)) or (layer1_outputs(392));
    layer2_outputs(5725) <= (layer1_outputs(2761)) and not (layer1_outputs(7148));
    layer2_outputs(5726) <= not(layer1_outputs(1701)) or (layer1_outputs(5958));
    layer2_outputs(5727) <= not(layer1_outputs(1588));
    layer2_outputs(5728) <= (layer1_outputs(107)) and not (layer1_outputs(775));
    layer2_outputs(5729) <= not(layer1_outputs(6893)) or (layer1_outputs(6284));
    layer2_outputs(5730) <= (layer1_outputs(3232)) and not (layer1_outputs(3706));
    layer2_outputs(5731) <= not((layer1_outputs(3803)) and (layer1_outputs(2582)));
    layer2_outputs(5732) <= not((layer1_outputs(6002)) and (layer1_outputs(4378)));
    layer2_outputs(5733) <= not(layer1_outputs(6336)) or (layer1_outputs(1148));
    layer2_outputs(5734) <= not((layer1_outputs(7633)) or (layer1_outputs(4970)));
    layer2_outputs(5735) <= not(layer1_outputs(3346)) or (layer1_outputs(6009));
    layer2_outputs(5736) <= layer1_outputs(4592);
    layer2_outputs(5737) <= not((layer1_outputs(5871)) and (layer1_outputs(7669)));
    layer2_outputs(5738) <= (layer1_outputs(2432)) or (layer1_outputs(6201));
    layer2_outputs(5739) <= not(layer1_outputs(6514)) or (layer1_outputs(2978));
    layer2_outputs(5740) <= not((layer1_outputs(6334)) or (layer1_outputs(2601)));
    layer2_outputs(5741) <= layer1_outputs(4877);
    layer2_outputs(5742) <= not(layer1_outputs(7167));
    layer2_outputs(5743) <= not(layer1_outputs(2499));
    layer2_outputs(5744) <= layer1_outputs(1647);
    layer2_outputs(5745) <= not((layer1_outputs(7262)) and (layer1_outputs(4207)));
    layer2_outputs(5746) <= not((layer1_outputs(2377)) and (layer1_outputs(3790)));
    layer2_outputs(5747) <= not(layer1_outputs(3943)) or (layer1_outputs(3061));
    layer2_outputs(5748) <= layer1_outputs(461);
    layer2_outputs(5749) <= not((layer1_outputs(6499)) and (layer1_outputs(5182)));
    layer2_outputs(5750) <= not((layer1_outputs(6420)) xor (layer1_outputs(1120)));
    layer2_outputs(5751) <= (layer1_outputs(3006)) and (layer1_outputs(7120));
    layer2_outputs(5752) <= not(layer1_outputs(24));
    layer2_outputs(5753) <= not(layer1_outputs(4894)) or (layer1_outputs(3524));
    layer2_outputs(5754) <= '1';
    layer2_outputs(5755) <= layer1_outputs(6317);
    layer2_outputs(5756) <= (layer1_outputs(3482)) and (layer1_outputs(6370));
    layer2_outputs(5757) <= not(layer1_outputs(3696)) or (layer1_outputs(2293));
    layer2_outputs(5758) <= not((layer1_outputs(7361)) and (layer1_outputs(4871)));
    layer2_outputs(5759) <= '1';
    layer2_outputs(5760) <= (layer1_outputs(4159)) and not (layer1_outputs(6998));
    layer2_outputs(5761) <= layer1_outputs(6740);
    layer2_outputs(5762) <= not((layer1_outputs(6399)) and (layer1_outputs(820)));
    layer2_outputs(5763) <= layer1_outputs(3572);
    layer2_outputs(5764) <= not((layer1_outputs(109)) and (layer1_outputs(2738)));
    layer2_outputs(5765) <= not(layer1_outputs(7014));
    layer2_outputs(5766) <= (layer1_outputs(3937)) xor (layer1_outputs(1015));
    layer2_outputs(5767) <= not((layer1_outputs(7252)) and (layer1_outputs(6888)));
    layer2_outputs(5768) <= not(layer1_outputs(7049));
    layer2_outputs(5769) <= not(layer1_outputs(7573)) or (layer1_outputs(5997));
    layer2_outputs(5770) <= '1';
    layer2_outputs(5771) <= not(layer1_outputs(7486));
    layer2_outputs(5772) <= not(layer1_outputs(3973)) or (layer1_outputs(4733));
    layer2_outputs(5773) <= (layer1_outputs(1381)) and not (layer1_outputs(3413));
    layer2_outputs(5774) <= (layer1_outputs(787)) and not (layer1_outputs(5921));
    layer2_outputs(5775) <= '1';
    layer2_outputs(5776) <= layer1_outputs(5761);
    layer2_outputs(5777) <= '1';
    layer2_outputs(5778) <= not((layer1_outputs(1018)) or (layer1_outputs(170)));
    layer2_outputs(5779) <= layer1_outputs(963);
    layer2_outputs(5780) <= (layer1_outputs(4961)) and (layer1_outputs(3145));
    layer2_outputs(5781) <= not(layer1_outputs(4422));
    layer2_outputs(5782) <= not(layer1_outputs(2616));
    layer2_outputs(5783) <= '1';
    layer2_outputs(5784) <= (layer1_outputs(6232)) and not (layer1_outputs(5177));
    layer2_outputs(5785) <= layer1_outputs(6777);
    layer2_outputs(5786) <= not(layer1_outputs(1667));
    layer2_outputs(5787) <= (layer1_outputs(415)) or (layer1_outputs(1122));
    layer2_outputs(5788) <= (layer1_outputs(6072)) and (layer1_outputs(4328));
    layer2_outputs(5789) <= (layer1_outputs(7537)) and not (layer1_outputs(196));
    layer2_outputs(5790) <= not(layer1_outputs(3354));
    layer2_outputs(5791) <= layer1_outputs(2167);
    layer2_outputs(5792) <= (layer1_outputs(2613)) or (layer1_outputs(4938));
    layer2_outputs(5793) <= '1';
    layer2_outputs(5794) <= layer1_outputs(5275);
    layer2_outputs(5795) <= '1';
    layer2_outputs(5796) <= not(layer1_outputs(290)) or (layer1_outputs(7253));
    layer2_outputs(5797) <= '0';
    layer2_outputs(5798) <= not((layer1_outputs(593)) and (layer1_outputs(3292)));
    layer2_outputs(5799) <= not(layer1_outputs(6371)) or (layer1_outputs(378));
    layer2_outputs(5800) <= not((layer1_outputs(888)) and (layer1_outputs(1661)));
    layer2_outputs(5801) <= (layer1_outputs(3599)) and (layer1_outputs(4003));
    layer2_outputs(5802) <= (layer1_outputs(3223)) xor (layer1_outputs(1418));
    layer2_outputs(5803) <= not((layer1_outputs(6980)) or (layer1_outputs(4075)));
    layer2_outputs(5804) <= layer1_outputs(2561);
    layer2_outputs(5805) <= (layer1_outputs(2524)) and not (layer1_outputs(7517));
    layer2_outputs(5806) <= layer1_outputs(1540);
    layer2_outputs(5807) <= not((layer1_outputs(2630)) or (layer1_outputs(6861)));
    layer2_outputs(5808) <= not(layer1_outputs(5952));
    layer2_outputs(5809) <= not(layer1_outputs(3576));
    layer2_outputs(5810) <= (layer1_outputs(1674)) and not (layer1_outputs(5182));
    layer2_outputs(5811) <= not(layer1_outputs(3789));
    layer2_outputs(5812) <= layer1_outputs(2615);
    layer2_outputs(5813) <= '0';
    layer2_outputs(5814) <= not(layer1_outputs(1798)) or (layer1_outputs(1135));
    layer2_outputs(5815) <= not(layer1_outputs(3902)) or (layer1_outputs(6142));
    layer2_outputs(5816) <= layer1_outputs(2612);
    layer2_outputs(5817) <= (layer1_outputs(2120)) and (layer1_outputs(7278));
    layer2_outputs(5818) <= layer1_outputs(2207);
    layer2_outputs(5819) <= not(layer1_outputs(3702)) or (layer1_outputs(1935));
    layer2_outputs(5820) <= (layer1_outputs(355)) and not (layer1_outputs(1501));
    layer2_outputs(5821) <= not(layer1_outputs(4171)) or (layer1_outputs(2386));
    layer2_outputs(5822) <= (layer1_outputs(54)) and not (layer1_outputs(5849));
    layer2_outputs(5823) <= not(layer1_outputs(3899));
    layer2_outputs(5824) <= (layer1_outputs(1364)) and not (layer1_outputs(1021));
    layer2_outputs(5825) <= not(layer1_outputs(4326)) or (layer1_outputs(5457));
    layer2_outputs(5826) <= not(layer1_outputs(4236));
    layer2_outputs(5827) <= not((layer1_outputs(7447)) or (layer1_outputs(600)));
    layer2_outputs(5828) <= layer1_outputs(3924);
    layer2_outputs(5829) <= layer1_outputs(4659);
    layer2_outputs(5830) <= not((layer1_outputs(5796)) and (layer1_outputs(3773)));
    layer2_outputs(5831) <= not(layer1_outputs(2184));
    layer2_outputs(5832) <= (layer1_outputs(217)) and not (layer1_outputs(5432));
    layer2_outputs(5833) <= '1';
    layer2_outputs(5834) <= (layer1_outputs(4647)) or (layer1_outputs(2436));
    layer2_outputs(5835) <= not(layer1_outputs(5331));
    layer2_outputs(5836) <= layer1_outputs(3224);
    layer2_outputs(5837) <= '1';
    layer2_outputs(5838) <= layer1_outputs(2027);
    layer2_outputs(5839) <= not(layer1_outputs(1135)) or (layer1_outputs(844));
    layer2_outputs(5840) <= layer1_outputs(4419);
    layer2_outputs(5841) <= not((layer1_outputs(4791)) or (layer1_outputs(1892)));
    layer2_outputs(5842) <= '1';
    layer2_outputs(5843) <= layer1_outputs(7677);
    layer2_outputs(5844) <= (layer1_outputs(4560)) and (layer1_outputs(7423));
    layer2_outputs(5845) <= (layer1_outputs(5687)) and not (layer1_outputs(7573));
    layer2_outputs(5846) <= '0';
    layer2_outputs(5847) <= (layer1_outputs(4116)) xor (layer1_outputs(596));
    layer2_outputs(5848) <= not(layer1_outputs(475)) or (layer1_outputs(5553));
    layer2_outputs(5849) <= not((layer1_outputs(1753)) or (layer1_outputs(1662)));
    layer2_outputs(5850) <= not(layer1_outputs(1680)) or (layer1_outputs(1157));
    layer2_outputs(5851) <= layer1_outputs(4715);
    layer2_outputs(5852) <= not((layer1_outputs(7329)) or (layer1_outputs(5623)));
    layer2_outputs(5853) <= (layer1_outputs(7601)) or (layer1_outputs(2036));
    layer2_outputs(5854) <= (layer1_outputs(4897)) or (layer1_outputs(7082));
    layer2_outputs(5855) <= (layer1_outputs(2270)) and not (layer1_outputs(5292));
    layer2_outputs(5856) <= (layer1_outputs(118)) and (layer1_outputs(4872));
    layer2_outputs(5857) <= (layer1_outputs(5166)) xor (layer1_outputs(863));
    layer2_outputs(5858) <= (layer1_outputs(1011)) and not (layer1_outputs(3787));
    layer2_outputs(5859) <= not((layer1_outputs(1157)) or (layer1_outputs(4600)));
    layer2_outputs(5860) <= not(layer1_outputs(5212));
    layer2_outputs(5861) <= not(layer1_outputs(7191));
    layer2_outputs(5862) <= layer1_outputs(1139);
    layer2_outputs(5863) <= layer1_outputs(4377);
    layer2_outputs(5864) <= not(layer1_outputs(6694));
    layer2_outputs(5865) <= not(layer1_outputs(2002)) or (layer1_outputs(7266));
    layer2_outputs(5866) <= layer1_outputs(959);
    layer2_outputs(5867) <= (layer1_outputs(3241)) and not (layer1_outputs(3100));
    layer2_outputs(5868) <= (layer1_outputs(4801)) or (layer1_outputs(7278));
    layer2_outputs(5869) <= (layer1_outputs(4213)) and not (layer1_outputs(5932));
    layer2_outputs(5870) <= layer1_outputs(4724);
    layer2_outputs(5871) <= not(layer1_outputs(3871));
    layer2_outputs(5872) <= (layer1_outputs(1374)) and (layer1_outputs(1584));
    layer2_outputs(5873) <= not(layer1_outputs(5951)) or (layer1_outputs(4835));
    layer2_outputs(5874) <= layer1_outputs(2099);
    layer2_outputs(5875) <= (layer1_outputs(935)) and (layer1_outputs(5905));
    layer2_outputs(5876) <= '0';
    layer2_outputs(5877) <= not((layer1_outputs(6086)) xor (layer1_outputs(3477)));
    layer2_outputs(5878) <= not(layer1_outputs(2141));
    layer2_outputs(5879) <= (layer1_outputs(7043)) xor (layer1_outputs(5520));
    layer2_outputs(5880) <= '0';
    layer2_outputs(5881) <= '1';
    layer2_outputs(5882) <= (layer1_outputs(2465)) and not (layer1_outputs(721));
    layer2_outputs(5883) <= not(layer1_outputs(6740));
    layer2_outputs(5884) <= not(layer1_outputs(1867));
    layer2_outputs(5885) <= not(layer1_outputs(4400));
    layer2_outputs(5886) <= not(layer1_outputs(2405)) or (layer1_outputs(2101));
    layer2_outputs(5887) <= not(layer1_outputs(4058));
    layer2_outputs(5888) <= (layer1_outputs(1072)) or (layer1_outputs(7240));
    layer2_outputs(5889) <= not(layer1_outputs(2977));
    layer2_outputs(5890) <= (layer1_outputs(2872)) and not (layer1_outputs(5464));
    layer2_outputs(5891) <= '1';
    layer2_outputs(5892) <= not(layer1_outputs(2461)) or (layer1_outputs(2363));
    layer2_outputs(5893) <= layer1_outputs(4601);
    layer2_outputs(5894) <= not((layer1_outputs(5648)) or (layer1_outputs(6238)));
    layer2_outputs(5895) <= layer1_outputs(2920);
    layer2_outputs(5896) <= '1';
    layer2_outputs(5897) <= (layer1_outputs(5390)) or (layer1_outputs(7478));
    layer2_outputs(5898) <= (layer1_outputs(1948)) and (layer1_outputs(4927));
    layer2_outputs(5899) <= '1';
    layer2_outputs(5900) <= layer1_outputs(781);
    layer2_outputs(5901) <= (layer1_outputs(2345)) and not (layer1_outputs(7002));
    layer2_outputs(5902) <= '1';
    layer2_outputs(5903) <= not(layer1_outputs(3950)) or (layer1_outputs(2097));
    layer2_outputs(5904) <= '0';
    layer2_outputs(5905) <= (layer1_outputs(2842)) and not (layer1_outputs(5315));
    layer2_outputs(5906) <= (layer1_outputs(1896)) and (layer1_outputs(4478));
    layer2_outputs(5907) <= '1';
    layer2_outputs(5908) <= (layer1_outputs(3411)) xor (layer1_outputs(3529));
    layer2_outputs(5909) <= (layer1_outputs(7608)) or (layer1_outputs(7335));
    layer2_outputs(5910) <= layer1_outputs(4879);
    layer2_outputs(5911) <= (layer1_outputs(6571)) and not (layer1_outputs(4062));
    layer2_outputs(5912) <= (layer1_outputs(2570)) and not (layer1_outputs(422));
    layer2_outputs(5913) <= (layer1_outputs(6810)) and (layer1_outputs(3055));
    layer2_outputs(5914) <= not(layer1_outputs(5870)) or (layer1_outputs(1531));
    layer2_outputs(5915) <= not(layer1_outputs(6672));
    layer2_outputs(5916) <= '1';
    layer2_outputs(5917) <= (layer1_outputs(4038)) and not (layer1_outputs(2795));
    layer2_outputs(5918) <= layer1_outputs(7007);
    layer2_outputs(5919) <= layer1_outputs(3588);
    layer2_outputs(5920) <= not(layer1_outputs(7081));
    layer2_outputs(5921) <= not(layer1_outputs(4953)) or (layer1_outputs(5357));
    layer2_outputs(5922) <= not(layer1_outputs(1206)) or (layer1_outputs(3676));
    layer2_outputs(5923) <= (layer1_outputs(6188)) and not (layer1_outputs(7394));
    layer2_outputs(5924) <= not((layer1_outputs(2282)) or (layer1_outputs(4824)));
    layer2_outputs(5925) <= not(layer1_outputs(4422));
    layer2_outputs(5926) <= not(layer1_outputs(3667)) or (layer1_outputs(5865));
    layer2_outputs(5927) <= (layer1_outputs(52)) and not (layer1_outputs(3530));
    layer2_outputs(5928) <= not((layer1_outputs(110)) and (layer1_outputs(3984)));
    layer2_outputs(5929) <= layer1_outputs(4949);
    layer2_outputs(5930) <= '1';
    layer2_outputs(5931) <= (layer1_outputs(3215)) and not (layer1_outputs(1117));
    layer2_outputs(5932) <= not((layer1_outputs(2232)) and (layer1_outputs(863)));
    layer2_outputs(5933) <= not(layer1_outputs(1801));
    layer2_outputs(5934) <= not((layer1_outputs(3497)) and (layer1_outputs(3500)));
    layer2_outputs(5935) <= (layer1_outputs(3030)) or (layer1_outputs(1041));
    layer2_outputs(5936) <= (layer1_outputs(1910)) and not (layer1_outputs(5830));
    layer2_outputs(5937) <= (layer1_outputs(315)) and not (layer1_outputs(897));
    layer2_outputs(5938) <= '0';
    layer2_outputs(5939) <= not(layer1_outputs(892)) or (layer1_outputs(6173));
    layer2_outputs(5940) <= not(layer1_outputs(6339));
    layer2_outputs(5941) <= '1';
    layer2_outputs(5942) <= layer1_outputs(7037);
    layer2_outputs(5943) <= not(layer1_outputs(4815)) or (layer1_outputs(5778));
    layer2_outputs(5944) <= (layer1_outputs(5398)) and not (layer1_outputs(1017));
    layer2_outputs(5945) <= (layer1_outputs(1178)) and not (layer1_outputs(700));
    layer2_outputs(5946) <= (layer1_outputs(5682)) and not (layer1_outputs(3193));
    layer2_outputs(5947) <= not(layer1_outputs(4588));
    layer2_outputs(5948) <= not((layer1_outputs(7321)) or (layer1_outputs(4869)));
    layer2_outputs(5949) <= not((layer1_outputs(4938)) xor (layer1_outputs(4364)));
    layer2_outputs(5950) <= '0';
    layer2_outputs(5951) <= (layer1_outputs(1698)) and not (layer1_outputs(2544));
    layer2_outputs(5952) <= layer1_outputs(1381);
    layer2_outputs(5953) <= (layer1_outputs(6992)) and not (layer1_outputs(6109));
    layer2_outputs(5954) <= not(layer1_outputs(1182));
    layer2_outputs(5955) <= not(layer1_outputs(5268)) or (layer1_outputs(2285));
    layer2_outputs(5956) <= not((layer1_outputs(7283)) or (layer1_outputs(5293)));
    layer2_outputs(5957) <= not(layer1_outputs(2775));
    layer2_outputs(5958) <= layer1_outputs(6066);
    layer2_outputs(5959) <= layer1_outputs(7041);
    layer2_outputs(5960) <= not(layer1_outputs(3328)) or (layer1_outputs(5717));
    layer2_outputs(5961) <= layer1_outputs(3127);
    layer2_outputs(5962) <= not(layer1_outputs(7440));
    layer2_outputs(5963) <= layer1_outputs(2771);
    layer2_outputs(5964) <= (layer1_outputs(50)) and not (layer1_outputs(1110));
    layer2_outputs(5965) <= not((layer1_outputs(7387)) or (layer1_outputs(5217)));
    layer2_outputs(5966) <= (layer1_outputs(2445)) and not (layer1_outputs(84));
    layer2_outputs(5967) <= '0';
    layer2_outputs(5968) <= '0';
    layer2_outputs(5969) <= layer1_outputs(7388);
    layer2_outputs(5970) <= (layer1_outputs(608)) and not (layer1_outputs(1346));
    layer2_outputs(5971) <= '1';
    layer2_outputs(5972) <= not(layer1_outputs(1065));
    layer2_outputs(5973) <= not(layer1_outputs(3995)) or (layer1_outputs(2149));
    layer2_outputs(5974) <= layer1_outputs(6437);
    layer2_outputs(5975) <= not(layer1_outputs(3997));
    layer2_outputs(5976) <= '1';
    layer2_outputs(5977) <= not(layer1_outputs(4625));
    layer2_outputs(5978) <= not((layer1_outputs(936)) or (layer1_outputs(4181)));
    layer2_outputs(5979) <= layer1_outputs(3639);
    layer2_outputs(5980) <= not(layer1_outputs(4130));
    layer2_outputs(5981) <= (layer1_outputs(4167)) or (layer1_outputs(2220));
    layer2_outputs(5982) <= not(layer1_outputs(3675)) or (layer1_outputs(3783));
    layer2_outputs(5983) <= not(layer1_outputs(5602));
    layer2_outputs(5984) <= layer1_outputs(2731);
    layer2_outputs(5985) <= not((layer1_outputs(818)) and (layer1_outputs(6081)));
    layer2_outputs(5986) <= (layer1_outputs(3954)) and not (layer1_outputs(1328));
    layer2_outputs(5987) <= not(layer1_outputs(411));
    layer2_outputs(5988) <= not((layer1_outputs(7227)) or (layer1_outputs(3608)));
    layer2_outputs(5989) <= (layer1_outputs(7405)) and (layer1_outputs(4448));
    layer2_outputs(5990) <= layer1_outputs(4490);
    layer2_outputs(5991) <= (layer1_outputs(6068)) and (layer1_outputs(7621));
    layer2_outputs(5992) <= not(layer1_outputs(4339)) or (layer1_outputs(2245));
    layer2_outputs(5993) <= not((layer1_outputs(402)) and (layer1_outputs(3570)));
    layer2_outputs(5994) <= '1';
    layer2_outputs(5995) <= not(layer1_outputs(3309));
    layer2_outputs(5996) <= not(layer1_outputs(6464)) or (layer1_outputs(4718));
    layer2_outputs(5997) <= '1';
    layer2_outputs(5998) <= not((layer1_outputs(6639)) or (layer1_outputs(5097)));
    layer2_outputs(5999) <= not(layer1_outputs(3326));
    layer2_outputs(6000) <= layer1_outputs(4172);
    layer2_outputs(6001) <= (layer1_outputs(3026)) and not (layer1_outputs(1845));
    layer2_outputs(6002) <= not(layer1_outputs(521));
    layer2_outputs(6003) <= (layer1_outputs(5001)) and not (layer1_outputs(5703));
    layer2_outputs(6004) <= not(layer1_outputs(5485));
    layer2_outputs(6005) <= not(layer1_outputs(2265));
    layer2_outputs(6006) <= not(layer1_outputs(653));
    layer2_outputs(6007) <= not(layer1_outputs(4000));
    layer2_outputs(6008) <= not(layer1_outputs(6506));
    layer2_outputs(6009) <= not((layer1_outputs(6476)) or (layer1_outputs(6434)));
    layer2_outputs(6010) <= (layer1_outputs(4829)) or (layer1_outputs(107));
    layer2_outputs(6011) <= not(layer1_outputs(6182));
    layer2_outputs(6012) <= (layer1_outputs(7084)) and (layer1_outputs(2931));
    layer2_outputs(6013) <= layer1_outputs(857);
    layer2_outputs(6014) <= layer1_outputs(5721);
    layer2_outputs(6015) <= not(layer1_outputs(2780));
    layer2_outputs(6016) <= '1';
    layer2_outputs(6017) <= layer1_outputs(7298);
    layer2_outputs(6018) <= not((layer1_outputs(5305)) or (layer1_outputs(4999)));
    layer2_outputs(6019) <= (layer1_outputs(1477)) and not (layer1_outputs(1696));
    layer2_outputs(6020) <= not(layer1_outputs(528));
    layer2_outputs(6021) <= '0';
    layer2_outputs(6022) <= not(layer1_outputs(5732)) or (layer1_outputs(1213));
    layer2_outputs(6023) <= not((layer1_outputs(1882)) or (layer1_outputs(6084)));
    layer2_outputs(6024) <= layer1_outputs(3759);
    layer2_outputs(6025) <= (layer1_outputs(4512)) and not (layer1_outputs(5242));
    layer2_outputs(6026) <= (layer1_outputs(1593)) or (layer1_outputs(6178));
    layer2_outputs(6027) <= not(layer1_outputs(777));
    layer2_outputs(6028) <= '1';
    layer2_outputs(6029) <= not(layer1_outputs(3807));
    layer2_outputs(6030) <= layer1_outputs(3467);
    layer2_outputs(6031) <= not((layer1_outputs(334)) xor (layer1_outputs(1679)));
    layer2_outputs(6032) <= not(layer1_outputs(4885)) or (layer1_outputs(7291));
    layer2_outputs(6033) <= (layer1_outputs(26)) or (layer1_outputs(7140));
    layer2_outputs(6034) <= not(layer1_outputs(60));
    layer2_outputs(6035) <= (layer1_outputs(4577)) xor (layer1_outputs(7108));
    layer2_outputs(6036) <= not(layer1_outputs(5620));
    layer2_outputs(6037) <= layer1_outputs(4580);
    layer2_outputs(6038) <= not(layer1_outputs(4108));
    layer2_outputs(6039) <= layer1_outputs(5440);
    layer2_outputs(6040) <= not(layer1_outputs(5619)) or (layer1_outputs(2035));
    layer2_outputs(6041) <= layer1_outputs(5208);
    layer2_outputs(6042) <= (layer1_outputs(1624)) and not (layer1_outputs(4057));
    layer2_outputs(6043) <= not(layer1_outputs(7312));
    layer2_outputs(6044) <= '0';
    layer2_outputs(6045) <= not(layer1_outputs(2020));
    layer2_outputs(6046) <= not(layer1_outputs(1515));
    layer2_outputs(6047) <= not((layer1_outputs(3412)) xor (layer1_outputs(4817)));
    layer2_outputs(6048) <= layer1_outputs(3472);
    layer2_outputs(6049) <= (layer1_outputs(3003)) or (layer1_outputs(4871));
    layer2_outputs(6050) <= not(layer1_outputs(3168));
    layer2_outputs(6051) <= not(layer1_outputs(5303)) or (layer1_outputs(3787));
    layer2_outputs(6052) <= not(layer1_outputs(3392)) or (layer1_outputs(2784));
    layer2_outputs(6053) <= (layer1_outputs(832)) and not (layer1_outputs(1247));
    layer2_outputs(6054) <= not(layer1_outputs(1548));
    layer2_outputs(6055) <= not(layer1_outputs(2818)) or (layer1_outputs(7619));
    layer2_outputs(6056) <= (layer1_outputs(1261)) and not (layer1_outputs(5103));
    layer2_outputs(6057) <= (layer1_outputs(4437)) and (layer1_outputs(6267));
    layer2_outputs(6058) <= layer1_outputs(7299);
    layer2_outputs(6059) <= (layer1_outputs(7184)) and (layer1_outputs(1461));
    layer2_outputs(6060) <= layer1_outputs(3185);
    layer2_outputs(6061) <= not((layer1_outputs(2043)) or (layer1_outputs(2190)));
    layer2_outputs(6062) <= '1';
    layer2_outputs(6063) <= not(layer1_outputs(3631));
    layer2_outputs(6064) <= not(layer1_outputs(159));
    layer2_outputs(6065) <= '0';
    layer2_outputs(6066) <= not(layer1_outputs(6989));
    layer2_outputs(6067) <= not(layer1_outputs(98)) or (layer1_outputs(901));
    layer2_outputs(6068) <= not(layer1_outputs(3114));
    layer2_outputs(6069) <= '1';
    layer2_outputs(6070) <= layer1_outputs(2792);
    layer2_outputs(6071) <= (layer1_outputs(10)) or (layer1_outputs(7104));
    layer2_outputs(6072) <= not(layer1_outputs(7239)) or (layer1_outputs(5555));
    layer2_outputs(6073) <= '1';
    layer2_outputs(6074) <= (layer1_outputs(1922)) or (layer1_outputs(5158));
    layer2_outputs(6075) <= layer1_outputs(376);
    layer2_outputs(6076) <= layer1_outputs(4464);
    layer2_outputs(6077) <= layer1_outputs(4875);
    layer2_outputs(6078) <= layer1_outputs(6013);
    layer2_outputs(6079) <= not(layer1_outputs(3167));
    layer2_outputs(6080) <= not(layer1_outputs(4942)) or (layer1_outputs(4205));
    layer2_outputs(6081) <= not(layer1_outputs(4272));
    layer2_outputs(6082) <= not((layer1_outputs(5048)) and (layer1_outputs(405)));
    layer2_outputs(6083) <= layer1_outputs(2118);
    layer2_outputs(6084) <= (layer1_outputs(5320)) and not (layer1_outputs(5181));
    layer2_outputs(6085) <= '0';
    layer2_outputs(6086) <= not(layer1_outputs(7539));
    layer2_outputs(6087) <= '1';
    layer2_outputs(6088) <= layer1_outputs(6785);
    layer2_outputs(6089) <= not(layer1_outputs(6844));
    layer2_outputs(6090) <= layer1_outputs(87);
    layer2_outputs(6091) <= not((layer1_outputs(3556)) or (layer1_outputs(456)));
    layer2_outputs(6092) <= layer1_outputs(2984);
    layer2_outputs(6093) <= not((layer1_outputs(5643)) or (layer1_outputs(2646)));
    layer2_outputs(6094) <= (layer1_outputs(1723)) and not (layer1_outputs(583));
    layer2_outputs(6095) <= (layer1_outputs(5373)) and (layer1_outputs(6983));
    layer2_outputs(6096) <= not(layer1_outputs(4985)) or (layer1_outputs(6003));
    layer2_outputs(6097) <= not((layer1_outputs(3895)) and (layer1_outputs(7236)));
    layer2_outputs(6098) <= (layer1_outputs(976)) and (layer1_outputs(2684));
    layer2_outputs(6099) <= not(layer1_outputs(1763)) or (layer1_outputs(2046));
    layer2_outputs(6100) <= not((layer1_outputs(4088)) and (layer1_outputs(3962)));
    layer2_outputs(6101) <= not((layer1_outputs(1013)) and (layer1_outputs(3062)));
    layer2_outputs(6102) <= (layer1_outputs(1436)) and not (layer1_outputs(3880));
    layer2_outputs(6103) <= not((layer1_outputs(2429)) or (layer1_outputs(5269)));
    layer2_outputs(6104) <= (layer1_outputs(3296)) and not (layer1_outputs(2153));
    layer2_outputs(6105) <= (layer1_outputs(6904)) and not (layer1_outputs(1729));
    layer2_outputs(6106) <= not((layer1_outputs(3657)) xor (layer1_outputs(697)));
    layer2_outputs(6107) <= (layer1_outputs(458)) and not (layer1_outputs(6258));
    layer2_outputs(6108) <= not(layer1_outputs(3683)) or (layer1_outputs(1642));
    layer2_outputs(6109) <= not(layer1_outputs(2694));
    layer2_outputs(6110) <= not(layer1_outputs(1573)) or (layer1_outputs(4227));
    layer2_outputs(6111) <= (layer1_outputs(271)) and not (layer1_outputs(313));
    layer2_outputs(6112) <= not((layer1_outputs(1602)) or (layer1_outputs(2184)));
    layer2_outputs(6113) <= not(layer1_outputs(195)) or (layer1_outputs(3165));
    layer2_outputs(6114) <= not(layer1_outputs(4718)) or (layer1_outputs(5455));
    layer2_outputs(6115) <= not(layer1_outputs(6878)) or (layer1_outputs(2334));
    layer2_outputs(6116) <= (layer1_outputs(3734)) or (layer1_outputs(2421));
    layer2_outputs(6117) <= layer1_outputs(3917);
    layer2_outputs(6118) <= not((layer1_outputs(2522)) xor (layer1_outputs(3454)));
    layer2_outputs(6119) <= layer1_outputs(5263);
    layer2_outputs(6120) <= '1';
    layer2_outputs(6121) <= (layer1_outputs(1573)) and not (layer1_outputs(3936));
    layer2_outputs(6122) <= not(layer1_outputs(105));
    layer2_outputs(6123) <= '0';
    layer2_outputs(6124) <= (layer1_outputs(6269)) and (layer1_outputs(4509));
    layer2_outputs(6125) <= (layer1_outputs(6166)) and not (layer1_outputs(1226));
    layer2_outputs(6126) <= (layer1_outputs(3171)) and not (layer1_outputs(6117));
    layer2_outputs(6127) <= not(layer1_outputs(5328));
    layer2_outputs(6128) <= '1';
    layer2_outputs(6129) <= '0';
    layer2_outputs(6130) <= not(layer1_outputs(5793));
    layer2_outputs(6131) <= not((layer1_outputs(2759)) or (layer1_outputs(4387)));
    layer2_outputs(6132) <= '1';
    layer2_outputs(6133) <= not(layer1_outputs(6679));
    layer2_outputs(6134) <= (layer1_outputs(6416)) and (layer1_outputs(4874));
    layer2_outputs(6135) <= not(layer1_outputs(1784));
    layer2_outputs(6136) <= not((layer1_outputs(1189)) and (layer1_outputs(3285)));
    layer2_outputs(6137) <= (layer1_outputs(3358)) and not (layer1_outputs(5356));
    layer2_outputs(6138) <= (layer1_outputs(4809)) and not (layer1_outputs(6468));
    layer2_outputs(6139) <= not((layer1_outputs(954)) or (layer1_outputs(3867)));
    layer2_outputs(6140) <= layer1_outputs(3000);
    layer2_outputs(6141) <= not(layer1_outputs(3700));
    layer2_outputs(6142) <= not(layer1_outputs(1268));
    layer2_outputs(6143) <= '0';
    layer2_outputs(6144) <= (layer1_outputs(558)) or (layer1_outputs(335));
    layer2_outputs(6145) <= layer1_outputs(7422);
    layer2_outputs(6146) <= not(layer1_outputs(676));
    layer2_outputs(6147) <= not(layer1_outputs(6021)) or (layer1_outputs(6365));
    layer2_outputs(6148) <= not(layer1_outputs(2567));
    layer2_outputs(6149) <= not((layer1_outputs(1347)) or (layer1_outputs(5086)));
    layer2_outputs(6150) <= '1';
    layer2_outputs(6151) <= '0';
    layer2_outputs(6152) <= (layer1_outputs(3155)) or (layer1_outputs(3043));
    layer2_outputs(6153) <= '1';
    layer2_outputs(6154) <= not(layer1_outputs(3951));
    layer2_outputs(6155) <= (layer1_outputs(6033)) or (layer1_outputs(2260));
    layer2_outputs(6156) <= not(layer1_outputs(1568));
    layer2_outputs(6157) <= not((layer1_outputs(6400)) or (layer1_outputs(4331)));
    layer2_outputs(6158) <= layer1_outputs(755);
    layer2_outputs(6159) <= (layer1_outputs(6124)) and not (layer1_outputs(7011));
    layer2_outputs(6160) <= not(layer1_outputs(5597));
    layer2_outputs(6161) <= (layer1_outputs(5080)) and not (layer1_outputs(4952));
    layer2_outputs(6162) <= not(layer1_outputs(5469)) or (layer1_outputs(4884));
    layer2_outputs(6163) <= not(layer1_outputs(1890)) or (layer1_outputs(2108));
    layer2_outputs(6164) <= not((layer1_outputs(207)) and (layer1_outputs(1287)));
    layer2_outputs(6165) <= not(layer1_outputs(2517)) or (layer1_outputs(4421));
    layer2_outputs(6166) <= (layer1_outputs(5684)) xor (layer1_outputs(5080));
    layer2_outputs(6167) <= not(layer1_outputs(4907));
    layer2_outputs(6168) <= '1';
    layer2_outputs(6169) <= not(layer1_outputs(4831));
    layer2_outputs(6170) <= '0';
    layer2_outputs(6171) <= not(layer1_outputs(6056)) or (layer1_outputs(2178));
    layer2_outputs(6172) <= layer1_outputs(2316);
    layer2_outputs(6173) <= layer1_outputs(4741);
    layer2_outputs(6174) <= not(layer1_outputs(5508));
    layer2_outputs(6175) <= '0';
    layer2_outputs(6176) <= (layer1_outputs(667)) and not (layer1_outputs(2973));
    layer2_outputs(6177) <= not(layer1_outputs(6967));
    layer2_outputs(6178) <= '1';
    layer2_outputs(6179) <= (layer1_outputs(454)) or (layer1_outputs(1438));
    layer2_outputs(6180) <= not(layer1_outputs(1180));
    layer2_outputs(6181) <= (layer1_outputs(3898)) and not (layer1_outputs(147));
    layer2_outputs(6182) <= not(layer1_outputs(2396));
    layer2_outputs(6183) <= layer1_outputs(2189);
    layer2_outputs(6184) <= '1';
    layer2_outputs(6185) <= not(layer1_outputs(2274));
    layer2_outputs(6186) <= not((layer1_outputs(3470)) or (layer1_outputs(4289)));
    layer2_outputs(6187) <= (layer1_outputs(3617)) or (layer1_outputs(5374));
    layer2_outputs(6188) <= not((layer1_outputs(4174)) or (layer1_outputs(5677)));
    layer2_outputs(6189) <= (layer1_outputs(1779)) and not (layer1_outputs(2298));
    layer2_outputs(6190) <= not(layer1_outputs(941));
    layer2_outputs(6191) <= not(layer1_outputs(202));
    layer2_outputs(6192) <= (layer1_outputs(3814)) xor (layer1_outputs(6079));
    layer2_outputs(6193) <= (layer1_outputs(6984)) and (layer1_outputs(6051));
    layer2_outputs(6194) <= (layer1_outputs(2715)) and (layer1_outputs(41));
    layer2_outputs(6195) <= not((layer1_outputs(2147)) and (layer1_outputs(49)));
    layer2_outputs(6196) <= layer1_outputs(7603);
    layer2_outputs(6197) <= not(layer1_outputs(32)) or (layer1_outputs(5895));
    layer2_outputs(6198) <= layer1_outputs(7375);
    layer2_outputs(6199) <= (layer1_outputs(7281)) and not (layer1_outputs(4373));
    layer2_outputs(6200) <= not(layer1_outputs(4611)) or (layer1_outputs(1192));
    layer2_outputs(6201) <= (layer1_outputs(4092)) and (layer1_outputs(3408));
    layer2_outputs(6202) <= '1';
    layer2_outputs(6203) <= not(layer1_outputs(3834)) or (layer1_outputs(7525));
    layer2_outputs(6204) <= not((layer1_outputs(1835)) and (layer1_outputs(2320)));
    layer2_outputs(6205) <= (layer1_outputs(6578)) xor (layer1_outputs(2481));
    layer2_outputs(6206) <= not(layer1_outputs(2949));
    layer2_outputs(6207) <= not((layer1_outputs(3352)) or (layer1_outputs(6479)));
    layer2_outputs(6208) <= layer1_outputs(7317);
    layer2_outputs(6209) <= (layer1_outputs(4855)) and not (layer1_outputs(4366));
    layer2_outputs(6210) <= '1';
    layer2_outputs(6211) <= layer1_outputs(1144);
    layer2_outputs(6212) <= not(layer1_outputs(2232)) or (layer1_outputs(5882));
    layer2_outputs(6213) <= not(layer1_outputs(7310)) or (layer1_outputs(7521));
    layer2_outputs(6214) <= not(layer1_outputs(6423)) or (layer1_outputs(4620));
    layer2_outputs(6215) <= (layer1_outputs(1292)) or (layer1_outputs(1598));
    layer2_outputs(6216) <= '1';
    layer2_outputs(6217) <= (layer1_outputs(1834)) or (layer1_outputs(6622));
    layer2_outputs(6218) <= not((layer1_outputs(3266)) or (layer1_outputs(6698)));
    layer2_outputs(6219) <= '0';
    layer2_outputs(6220) <= not((layer1_outputs(3623)) and (layer1_outputs(7213)));
    layer2_outputs(6221) <= not(layer1_outputs(6059));
    layer2_outputs(6222) <= not(layer1_outputs(6362)) or (layer1_outputs(7296));
    layer2_outputs(6223) <= not((layer1_outputs(3012)) and (layer1_outputs(146)));
    layer2_outputs(6224) <= not((layer1_outputs(5113)) or (layer1_outputs(3747)));
    layer2_outputs(6225) <= not((layer1_outputs(6194)) xor (layer1_outputs(1396)));
    layer2_outputs(6226) <= (layer1_outputs(4433)) and not (layer1_outputs(2312));
    layer2_outputs(6227) <= layer1_outputs(4361);
    layer2_outputs(6228) <= not(layer1_outputs(2688)) or (layer1_outputs(4680));
    layer2_outputs(6229) <= not(layer1_outputs(5427));
    layer2_outputs(6230) <= layer1_outputs(3175);
    layer2_outputs(6231) <= not((layer1_outputs(3446)) or (layer1_outputs(5371)));
    layer2_outputs(6232) <= layer1_outputs(2696);
    layer2_outputs(6233) <= (layer1_outputs(1104)) and not (layer1_outputs(5086));
    layer2_outputs(6234) <= not(layer1_outputs(6456));
    layer2_outputs(6235) <= not((layer1_outputs(1857)) and (layer1_outputs(4573)));
    layer2_outputs(6236) <= (layer1_outputs(4637)) or (layer1_outputs(2573));
    layer2_outputs(6237) <= layer1_outputs(3649);
    layer2_outputs(6238) <= not(layer1_outputs(1490));
    layer2_outputs(6239) <= '0';
    layer2_outputs(6240) <= '1';
    layer2_outputs(6241) <= not(layer1_outputs(3021));
    layer2_outputs(6242) <= not(layer1_outputs(2261));
    layer2_outputs(6243) <= not((layer1_outputs(1101)) and (layer1_outputs(2423)));
    layer2_outputs(6244) <= (layer1_outputs(6085)) or (layer1_outputs(6204));
    layer2_outputs(6245) <= not(layer1_outputs(2911));
    layer2_outputs(6246) <= not((layer1_outputs(7133)) and (layer1_outputs(5762)));
    layer2_outputs(6247) <= not(layer1_outputs(381));
    layer2_outputs(6248) <= '1';
    layer2_outputs(6249) <= (layer1_outputs(5839)) and not (layer1_outputs(2325));
    layer2_outputs(6250) <= layer1_outputs(1562);
    layer2_outputs(6251) <= not(layer1_outputs(3661));
    layer2_outputs(6252) <= (layer1_outputs(5484)) and not (layer1_outputs(7138));
    layer2_outputs(6253) <= not(layer1_outputs(2614));
    layer2_outputs(6254) <= (layer1_outputs(2143)) xor (layer1_outputs(6538));
    layer2_outputs(6255) <= (layer1_outputs(568)) or (layer1_outputs(6031));
    layer2_outputs(6256) <= (layer1_outputs(5324)) and not (layer1_outputs(5334));
    layer2_outputs(6257) <= not(layer1_outputs(4468)) or (layer1_outputs(7193));
    layer2_outputs(6258) <= not((layer1_outputs(2499)) or (layer1_outputs(1863)));
    layer2_outputs(6259) <= (layer1_outputs(1837)) and not (layer1_outputs(1425));
    layer2_outputs(6260) <= '0';
    layer2_outputs(6261) <= (layer1_outputs(491)) and not (layer1_outputs(5826));
    layer2_outputs(6262) <= layer1_outputs(72);
    layer2_outputs(6263) <= layer1_outputs(5383);
    layer2_outputs(6264) <= layer1_outputs(4965);
    layer2_outputs(6265) <= (layer1_outputs(2442)) and not (layer1_outputs(6056));
    layer2_outputs(6266) <= '0';
    layer2_outputs(6267) <= layer1_outputs(3629);
    layer2_outputs(6268) <= not(layer1_outputs(5971)) or (layer1_outputs(5559));
    layer2_outputs(6269) <= not(layer1_outputs(2309)) or (layer1_outputs(2820));
    layer2_outputs(6270) <= (layer1_outputs(803)) and (layer1_outputs(2117));
    layer2_outputs(6271) <= not(layer1_outputs(5736));
    layer2_outputs(6272) <= not(layer1_outputs(3474)) or (layer1_outputs(4548));
    layer2_outputs(6273) <= (layer1_outputs(1955)) and not (layer1_outputs(1174));
    layer2_outputs(6274) <= layer1_outputs(2330);
    layer2_outputs(6275) <= (layer1_outputs(882)) or (layer1_outputs(6275));
    layer2_outputs(6276) <= (layer1_outputs(6907)) and not (layer1_outputs(1942));
    layer2_outputs(6277) <= '0';
    layer2_outputs(6278) <= (layer1_outputs(2888)) and (layer1_outputs(2117));
    layer2_outputs(6279) <= not(layer1_outputs(13)) or (layer1_outputs(797));
    layer2_outputs(6280) <= (layer1_outputs(2233)) and (layer1_outputs(6028));
    layer2_outputs(6281) <= not(layer1_outputs(3434));
    layer2_outputs(6282) <= not((layer1_outputs(6615)) and (layer1_outputs(1093)));
    layer2_outputs(6283) <= not(layer1_outputs(3248)) or (layer1_outputs(2078));
    layer2_outputs(6284) <= (layer1_outputs(4514)) or (layer1_outputs(5391));
    layer2_outputs(6285) <= layer1_outputs(3265);
    layer2_outputs(6286) <= '0';
    layer2_outputs(6287) <= layer1_outputs(2239);
    layer2_outputs(6288) <= (layer1_outputs(5019)) and (layer1_outputs(4232));
    layer2_outputs(6289) <= (layer1_outputs(5459)) and not (layer1_outputs(2083));
    layer2_outputs(6290) <= not(layer1_outputs(4743)) or (layer1_outputs(7205));
    layer2_outputs(6291) <= (layer1_outputs(2439)) and not (layer1_outputs(3096));
    layer2_outputs(6292) <= not(layer1_outputs(1915));
    layer2_outputs(6293) <= (layer1_outputs(445)) and not (layer1_outputs(5187));
    layer2_outputs(6294) <= (layer1_outputs(1583)) and not (layer1_outputs(5064));
    layer2_outputs(6295) <= '1';
    layer2_outputs(6296) <= not(layer1_outputs(1044)) or (layer1_outputs(3072));
    layer2_outputs(6297) <= not((layer1_outputs(7105)) and (layer1_outputs(2538)));
    layer2_outputs(6298) <= not((layer1_outputs(6069)) or (layer1_outputs(6930)));
    layer2_outputs(6299) <= '0';
    layer2_outputs(6300) <= (layer1_outputs(3301)) and not (layer1_outputs(339));
    layer2_outputs(6301) <= not((layer1_outputs(1013)) and (layer1_outputs(3138)));
    layer2_outputs(6302) <= not(layer1_outputs(5628));
    layer2_outputs(6303) <= (layer1_outputs(4067)) and not (layer1_outputs(6623));
    layer2_outputs(6304) <= (layer1_outputs(5549)) and not (layer1_outputs(9));
    layer2_outputs(6305) <= (layer1_outputs(2390)) and not (layer1_outputs(2213));
    layer2_outputs(6306) <= (layer1_outputs(6324)) and (layer1_outputs(7352));
    layer2_outputs(6307) <= (layer1_outputs(2938)) and (layer1_outputs(6300));
    layer2_outputs(6308) <= not(layer1_outputs(4296));
    layer2_outputs(6309) <= '0';
    layer2_outputs(6310) <= (layer1_outputs(1892)) and not (layer1_outputs(7416));
    layer2_outputs(6311) <= (layer1_outputs(878)) and not (layer1_outputs(7463));
    layer2_outputs(6312) <= layer1_outputs(7338);
    layer2_outputs(6313) <= layer1_outputs(616);
    layer2_outputs(6314) <= not((layer1_outputs(5223)) or (layer1_outputs(7306)));
    layer2_outputs(6315) <= (layer1_outputs(6775)) and not (layer1_outputs(4933));
    layer2_outputs(6316) <= not((layer1_outputs(756)) or (layer1_outputs(282)));
    layer2_outputs(6317) <= (layer1_outputs(1373)) xor (layer1_outputs(6138));
    layer2_outputs(6318) <= layer1_outputs(5751);
    layer2_outputs(6319) <= not(layer1_outputs(6298));
    layer2_outputs(6320) <= not(layer1_outputs(673)) or (layer1_outputs(2329));
    layer2_outputs(6321) <= layer1_outputs(318);
    layer2_outputs(6322) <= not(layer1_outputs(3395));
    layer2_outputs(6323) <= '1';
    layer2_outputs(6324) <= not(layer1_outputs(2014)) or (layer1_outputs(6798));
    layer2_outputs(6325) <= (layer1_outputs(2326)) or (layer1_outputs(1864));
    layer2_outputs(6326) <= not(layer1_outputs(6369)) or (layer1_outputs(1710));
    layer2_outputs(6327) <= (layer1_outputs(2306)) and (layer1_outputs(1718));
    layer2_outputs(6328) <= '0';
    layer2_outputs(6329) <= not(layer1_outputs(2728));
    layer2_outputs(6330) <= not(layer1_outputs(3056));
    layer2_outputs(6331) <= not(layer1_outputs(4458));
    layer2_outputs(6332) <= not(layer1_outputs(3832)) or (layer1_outputs(968));
    layer2_outputs(6333) <= not((layer1_outputs(562)) or (layer1_outputs(160)));
    layer2_outputs(6334) <= layer1_outputs(7670);
    layer2_outputs(6335) <= layer1_outputs(2865);
    layer2_outputs(6336) <= (layer1_outputs(2986)) and not (layer1_outputs(4877));
    layer2_outputs(6337) <= (layer1_outputs(337)) and not (layer1_outputs(5158));
    layer2_outputs(6338) <= not(layer1_outputs(5018));
    layer2_outputs(6339) <= not(layer1_outputs(6754));
    layer2_outputs(6340) <= '1';
    layer2_outputs(6341) <= '0';
    layer2_outputs(6342) <= not((layer1_outputs(4562)) and (layer1_outputs(6601)));
    layer2_outputs(6343) <= not(layer1_outputs(6896));
    layer2_outputs(6344) <= not(layer1_outputs(3921));
    layer2_outputs(6345) <= layer1_outputs(763);
    layer2_outputs(6346) <= layer1_outputs(1152);
    layer2_outputs(6347) <= not((layer1_outputs(58)) xor (layer1_outputs(7667)));
    layer2_outputs(6348) <= (layer1_outputs(143)) and (layer1_outputs(6208));
    layer2_outputs(6349) <= layer1_outputs(334);
    layer2_outputs(6350) <= '0';
    layer2_outputs(6351) <= not(layer1_outputs(675)) or (layer1_outputs(7095));
    layer2_outputs(6352) <= not(layer1_outputs(5729)) or (layer1_outputs(5947));
    layer2_outputs(6353) <= not(layer1_outputs(6283));
    layer2_outputs(6354) <= layer1_outputs(5451);
    layer2_outputs(6355) <= not((layer1_outputs(2944)) and (layer1_outputs(7295)));
    layer2_outputs(6356) <= layer1_outputs(6191);
    layer2_outputs(6357) <= not(layer1_outputs(1345));
    layer2_outputs(6358) <= layer1_outputs(3455);
    layer2_outputs(6359) <= layer1_outputs(4481);
    layer2_outputs(6360) <= not(layer1_outputs(3862)) or (layer1_outputs(6852));
    layer2_outputs(6361) <= (layer1_outputs(4627)) xor (layer1_outputs(3685));
    layer2_outputs(6362) <= (layer1_outputs(3713)) xor (layer1_outputs(4362));
    layer2_outputs(6363) <= layer1_outputs(989);
    layer2_outputs(6364) <= not(layer1_outputs(6518)) or (layer1_outputs(7134));
    layer2_outputs(6365) <= not((layer1_outputs(38)) and (layer1_outputs(1939)));
    layer2_outputs(6366) <= (layer1_outputs(4597)) and (layer1_outputs(4494));
    layer2_outputs(6367) <= not((layer1_outputs(2269)) or (layer1_outputs(2255)));
    layer2_outputs(6368) <= layer1_outputs(340);
    layer2_outputs(6369) <= (layer1_outputs(1069)) and not (layer1_outputs(2964));
    layer2_outputs(6370) <= not(layer1_outputs(4426)) or (layer1_outputs(4822));
    layer2_outputs(6371) <= not((layer1_outputs(4560)) and (layer1_outputs(2687)));
    layer2_outputs(6372) <= (layer1_outputs(7320)) or (layer1_outputs(3721));
    layer2_outputs(6373) <= not(layer1_outputs(6955));
    layer2_outputs(6374) <= not(layer1_outputs(6741)) or (layer1_outputs(6359));
    layer2_outputs(6375) <= layer1_outputs(436);
    layer2_outputs(6376) <= not(layer1_outputs(1443)) or (layer1_outputs(458));
    layer2_outputs(6377) <= not(layer1_outputs(404));
    layer2_outputs(6378) <= (layer1_outputs(2356)) and not (layer1_outputs(3561));
    layer2_outputs(6379) <= (layer1_outputs(5897)) and not (layer1_outputs(6585));
    layer2_outputs(6380) <= '0';
    layer2_outputs(6381) <= layer1_outputs(2981);
    layer2_outputs(6382) <= layer1_outputs(6228);
    layer2_outputs(6383) <= not(layer1_outputs(5728)) or (layer1_outputs(657));
    layer2_outputs(6384) <= layer1_outputs(4631);
    layer2_outputs(6385) <= '0';
    layer2_outputs(6386) <= not((layer1_outputs(7625)) or (layer1_outputs(7414)));
    layer2_outputs(6387) <= (layer1_outputs(4006)) and (layer1_outputs(1615));
    layer2_outputs(6388) <= layer1_outputs(1417);
    layer2_outputs(6389) <= (layer1_outputs(4527)) and not (layer1_outputs(7366));
    layer2_outputs(6390) <= (layer1_outputs(3060)) and not (layer1_outputs(1385));
    layer2_outputs(6391) <= '1';
    layer2_outputs(6392) <= not((layer1_outputs(6062)) and (layer1_outputs(5332)));
    layer2_outputs(6393) <= (layer1_outputs(5949)) or (layer1_outputs(6633));
    layer2_outputs(6394) <= not((layer1_outputs(3534)) or (layer1_outputs(3011)));
    layer2_outputs(6395) <= '0';
    layer2_outputs(6396) <= (layer1_outputs(1462)) and not (layer1_outputs(666));
    layer2_outputs(6397) <= (layer1_outputs(1863)) and (layer1_outputs(5978));
    layer2_outputs(6398) <= layer1_outputs(7157);
    layer2_outputs(6399) <= not(layer1_outputs(2717)) or (layer1_outputs(3882));
    layer2_outputs(6400) <= not(layer1_outputs(273));
    layer2_outputs(6401) <= not(layer1_outputs(544)) or (layer1_outputs(473));
    layer2_outputs(6402) <= not(layer1_outputs(7530));
    layer2_outputs(6403) <= not(layer1_outputs(4578));
    layer2_outputs(6404) <= layer1_outputs(6013);
    layer2_outputs(6405) <= (layer1_outputs(723)) or (layer1_outputs(7373));
    layer2_outputs(6406) <= '0';
    layer2_outputs(6407) <= (layer1_outputs(1828)) and not (layer1_outputs(7078));
    layer2_outputs(6408) <= '0';
    layer2_outputs(6409) <= (layer1_outputs(6748)) xor (layer1_outputs(2493));
    layer2_outputs(6410) <= layer1_outputs(5151);
    layer2_outputs(6411) <= not(layer1_outputs(3525));
    layer2_outputs(6412) <= not(layer1_outputs(6960));
    layer2_outputs(6413) <= not((layer1_outputs(2017)) and (layer1_outputs(2682)));
    layer2_outputs(6414) <= layer1_outputs(6069);
    layer2_outputs(6415) <= not((layer1_outputs(5321)) and (layer1_outputs(5645)));
    layer2_outputs(6416) <= (layer1_outputs(7334)) and not (layer1_outputs(3153));
    layer2_outputs(6417) <= not(layer1_outputs(2674));
    layer2_outputs(6418) <= (layer1_outputs(4093)) or (layer1_outputs(6340));
    layer2_outputs(6419) <= '1';
    layer2_outputs(6420) <= '0';
    layer2_outputs(6421) <= not(layer1_outputs(2590)) or (layer1_outputs(5240));
    layer2_outputs(6422) <= not((layer1_outputs(161)) or (layer1_outputs(4268)));
    layer2_outputs(6423) <= layer1_outputs(4771);
    layer2_outputs(6424) <= (layer1_outputs(7229)) and not (layer1_outputs(5960));
    layer2_outputs(6425) <= (layer1_outputs(2761)) and (layer1_outputs(6835));
    layer2_outputs(6426) <= not(layer1_outputs(5957)) or (layer1_outputs(6357));
    layer2_outputs(6427) <= layer1_outputs(1429);
    layer2_outputs(6428) <= (layer1_outputs(5361)) and (layer1_outputs(2112));
    layer2_outputs(6429) <= '1';
    layer2_outputs(6430) <= not(layer1_outputs(4829));
    layer2_outputs(6431) <= not(layer1_outputs(3547));
    layer2_outputs(6432) <= not(layer1_outputs(4908)) or (layer1_outputs(3452));
    layer2_outputs(6433) <= (layer1_outputs(4863)) and not (layer1_outputs(920));
    layer2_outputs(6434) <= not(layer1_outputs(512)) or (layer1_outputs(2078));
    layer2_outputs(6435) <= '0';
    layer2_outputs(6436) <= '1';
    layer2_outputs(6437) <= not(layer1_outputs(3881)) or (layer1_outputs(5473));
    layer2_outputs(6438) <= layer1_outputs(56);
    layer2_outputs(6439) <= (layer1_outputs(1428)) and not (layer1_outputs(7660));
    layer2_outputs(6440) <= not(layer1_outputs(7395)) or (layer1_outputs(2750));
    layer2_outputs(6441) <= not((layer1_outputs(6201)) and (layer1_outputs(88)));
    layer2_outputs(6442) <= '1';
    layer2_outputs(6443) <= (layer1_outputs(4709)) and not (layer1_outputs(2046));
    layer2_outputs(6444) <= not(layer1_outputs(5641)) or (layer1_outputs(6333));
    layer2_outputs(6445) <= '0';
    layer2_outputs(6446) <= not(layer1_outputs(2473));
    layer2_outputs(6447) <= (layer1_outputs(237)) and (layer1_outputs(2071));
    layer2_outputs(6448) <= (layer1_outputs(1087)) and not (layer1_outputs(4770));
    layer2_outputs(6449) <= not(layer1_outputs(7679));
    layer2_outputs(6450) <= '1';
    layer2_outputs(6451) <= not((layer1_outputs(1453)) or (layer1_outputs(6309)));
    layer2_outputs(6452) <= (layer1_outputs(1223)) and not (layer1_outputs(3505));
    layer2_outputs(6453) <= (layer1_outputs(5483)) and not (layer1_outputs(6994));
    layer2_outputs(6454) <= (layer1_outputs(2868)) and not (layer1_outputs(5711));
    layer2_outputs(6455) <= (layer1_outputs(1978)) and not (layer1_outputs(2443));
    layer2_outputs(6456) <= layer1_outputs(3998);
    layer2_outputs(6457) <= (layer1_outputs(1737)) or (layer1_outputs(2218));
    layer2_outputs(6458) <= (layer1_outputs(3982)) and (layer1_outputs(1649));
    layer2_outputs(6459) <= (layer1_outputs(7303)) or (layer1_outputs(539));
    layer2_outputs(6460) <= (layer1_outputs(6392)) and (layer1_outputs(3701));
    layer2_outputs(6461) <= not((layer1_outputs(6952)) and (layer1_outputs(2817)));
    layer2_outputs(6462) <= not(layer1_outputs(1032));
    layer2_outputs(6463) <= '0';
    layer2_outputs(6464) <= layer1_outputs(5312);
    layer2_outputs(6465) <= (layer1_outputs(2313)) and not (layer1_outputs(3010));
    layer2_outputs(6466) <= '0';
    layer2_outputs(6467) <= not(layer1_outputs(6162)) or (layer1_outputs(1422));
    layer2_outputs(6468) <= (layer1_outputs(4731)) or (layer1_outputs(5945));
    layer2_outputs(6469) <= layer1_outputs(1685);
    layer2_outputs(6470) <= not((layer1_outputs(7201)) or (layer1_outputs(4643)));
    layer2_outputs(6471) <= not((layer1_outputs(4626)) or (layer1_outputs(5313)));
    layer2_outputs(6472) <= layer1_outputs(2351);
    layer2_outputs(6473) <= not(layer1_outputs(6863));
    layer2_outputs(6474) <= '0';
    layer2_outputs(6475) <= layer1_outputs(6729);
    layer2_outputs(6476) <= layer1_outputs(6748);
    layer2_outputs(6477) <= not(layer1_outputs(5884)) or (layer1_outputs(231));
    layer2_outputs(6478) <= layer1_outputs(2215);
    layer2_outputs(6479) <= not(layer1_outputs(7498));
    layer2_outputs(6480) <= (layer1_outputs(815)) and (layer1_outputs(510));
    layer2_outputs(6481) <= not((layer1_outputs(5480)) and (layer1_outputs(4028)));
    layer2_outputs(6482) <= (layer1_outputs(6548)) and not (layer1_outputs(4890));
    layer2_outputs(6483) <= not(layer1_outputs(1742));
    layer2_outputs(6484) <= (layer1_outputs(6542)) and not (layer1_outputs(6846));
    layer2_outputs(6485) <= (layer1_outputs(2121)) or (layer1_outputs(207));
    layer2_outputs(6486) <= not(layer1_outputs(876)) or (layer1_outputs(3375));
    layer2_outputs(6487) <= not(layer1_outputs(5209));
    layer2_outputs(6488) <= (layer1_outputs(6697)) or (layer1_outputs(4453));
    layer2_outputs(6489) <= layer1_outputs(3716);
    layer2_outputs(6490) <= '1';
    layer2_outputs(6491) <= '1';
    layer2_outputs(6492) <= layer1_outputs(7028);
    layer2_outputs(6493) <= (layer1_outputs(6198)) and not (layer1_outputs(293));
    layer2_outputs(6494) <= not(layer1_outputs(5634)) or (layer1_outputs(3050));
    layer2_outputs(6495) <= (layer1_outputs(5130)) or (layer1_outputs(1623));
    layer2_outputs(6496) <= not(layer1_outputs(5420));
    layer2_outputs(6497) <= not(layer1_outputs(4612));
    layer2_outputs(6498) <= not(layer1_outputs(1524));
    layer2_outputs(6499) <= not((layer1_outputs(3375)) and (layer1_outputs(6411)));
    layer2_outputs(6500) <= (layer1_outputs(445)) and (layer1_outputs(7299));
    layer2_outputs(6501) <= (layer1_outputs(2804)) and not (layer1_outputs(3113));
    layer2_outputs(6502) <= (layer1_outputs(5367)) and not (layer1_outputs(373));
    layer2_outputs(6503) <= (layer1_outputs(3402)) and (layer1_outputs(7111));
    layer2_outputs(6504) <= layer1_outputs(3);
    layer2_outputs(6505) <= not((layer1_outputs(2433)) or (layer1_outputs(7629)));
    layer2_outputs(6506) <= '0';
    layer2_outputs(6507) <= layer1_outputs(5549);
    layer2_outputs(6508) <= not((layer1_outputs(6417)) and (layer1_outputs(3176)));
    layer2_outputs(6509) <= (layer1_outputs(3677)) and (layer1_outputs(2131));
    layer2_outputs(6510) <= not((layer1_outputs(6821)) and (layer1_outputs(5186)));
    layer2_outputs(6511) <= not((layer1_outputs(4945)) or (layer1_outputs(4582)));
    layer2_outputs(6512) <= '0';
    layer2_outputs(6513) <= (layer1_outputs(5844)) xor (layer1_outputs(6055));
    layer2_outputs(6514) <= (layer1_outputs(3678)) and not (layer1_outputs(5367));
    layer2_outputs(6515) <= (layer1_outputs(3993)) and (layer1_outputs(88));
    layer2_outputs(6516) <= (layer1_outputs(5102)) and not (layer1_outputs(3975));
    layer2_outputs(6517) <= not(layer1_outputs(4809)) or (layer1_outputs(6394));
    layer2_outputs(6518) <= not(layer1_outputs(6894));
    layer2_outputs(6519) <= not((layer1_outputs(6405)) or (layer1_outputs(3243)));
    layer2_outputs(6520) <= not(layer1_outputs(1900));
    layer2_outputs(6521) <= '0';
    layer2_outputs(6522) <= not(layer1_outputs(3696)) or (layer1_outputs(5373));
    layer2_outputs(6523) <= not((layer1_outputs(5079)) and (layer1_outputs(1227)));
    layer2_outputs(6524) <= (layer1_outputs(2756)) and not (layer1_outputs(1204));
    layer2_outputs(6525) <= layer1_outputs(1353);
    layer2_outputs(6526) <= not(layer1_outputs(4423));
    layer2_outputs(6527) <= not(layer1_outputs(382));
    layer2_outputs(6528) <= layer1_outputs(5098);
    layer2_outputs(6529) <= '1';
    layer2_outputs(6530) <= '1';
    layer2_outputs(6531) <= not(layer1_outputs(3610));
    layer2_outputs(6532) <= not((layer1_outputs(5699)) or (layer1_outputs(4293)));
    layer2_outputs(6533) <= not((layer1_outputs(7474)) and (layer1_outputs(6040)));
    layer2_outputs(6534) <= '1';
    layer2_outputs(6535) <= (layer1_outputs(4493)) and not (layer1_outputs(985));
    layer2_outputs(6536) <= not(layer1_outputs(4151));
    layer2_outputs(6537) <= not(layer1_outputs(5202)) or (layer1_outputs(3626));
    layer2_outputs(6538) <= '0';
    layer2_outputs(6539) <= layer1_outputs(5911);
    layer2_outputs(6540) <= not(layer1_outputs(3612));
    layer2_outputs(6541) <= not((layer1_outputs(5423)) and (layer1_outputs(725)));
    layer2_outputs(6542) <= (layer1_outputs(3063)) or (layer1_outputs(6768));
    layer2_outputs(6543) <= (layer1_outputs(2597)) or (layer1_outputs(6677));
    layer2_outputs(6544) <= '1';
    layer2_outputs(6545) <= '0';
    layer2_outputs(6546) <= '1';
    layer2_outputs(6547) <= (layer1_outputs(6373)) and (layer1_outputs(6763));
    layer2_outputs(6548) <= not(layer1_outputs(1233));
    layer2_outputs(6549) <= '0';
    layer2_outputs(6550) <= layer1_outputs(3204);
    layer2_outputs(6551) <= not(layer1_outputs(1913));
    layer2_outputs(6552) <= not(layer1_outputs(4375));
    layer2_outputs(6553) <= not(layer1_outputs(6749));
    layer2_outputs(6554) <= (layer1_outputs(3040)) xor (layer1_outputs(6374));
    layer2_outputs(6555) <= (layer1_outputs(7483)) xor (layer1_outputs(5366));
    layer2_outputs(6556) <= not((layer1_outputs(2344)) or (layer1_outputs(4760)));
    layer2_outputs(6557) <= not((layer1_outputs(2696)) and (layer1_outputs(1151)));
    layer2_outputs(6558) <= (layer1_outputs(5066)) and not (layer1_outputs(2956));
    layer2_outputs(6559) <= '0';
    layer2_outputs(6560) <= layer1_outputs(2541);
    layer2_outputs(6561) <= layer1_outputs(2353);
    layer2_outputs(6562) <= '0';
    layer2_outputs(6563) <= not(layer1_outputs(4031));
    layer2_outputs(6564) <= not(layer1_outputs(7553)) or (layer1_outputs(211));
    layer2_outputs(6565) <= (layer1_outputs(4336)) and (layer1_outputs(1584));
    layer2_outputs(6566) <= (layer1_outputs(4059)) and (layer1_outputs(6563));
    layer2_outputs(6567) <= (layer1_outputs(6850)) and (layer1_outputs(3953));
    layer2_outputs(6568) <= not(layer1_outputs(3539)) or (layer1_outputs(7069));
    layer2_outputs(6569) <= (layer1_outputs(7254)) xor (layer1_outputs(585));
    layer2_outputs(6570) <= (layer1_outputs(6811)) or (layer1_outputs(4511));
    layer2_outputs(6571) <= layer1_outputs(3184);
    layer2_outputs(6572) <= not((layer1_outputs(7431)) or (layer1_outputs(3865)));
    layer2_outputs(6573) <= layer1_outputs(7398);
    layer2_outputs(6574) <= layer1_outputs(1562);
    layer2_outputs(6575) <= layer1_outputs(6796);
    layer2_outputs(6576) <= not(layer1_outputs(1047)) or (layer1_outputs(6556));
    layer2_outputs(6577) <= not((layer1_outputs(6745)) and (layer1_outputs(7280)));
    layer2_outputs(6578) <= not(layer1_outputs(2380)) or (layer1_outputs(6123));
    layer2_outputs(6579) <= '0';
    layer2_outputs(6580) <= layer1_outputs(2867);
    layer2_outputs(6581) <= layer1_outputs(7177);
    layer2_outputs(6582) <= layer1_outputs(110);
    layer2_outputs(6583) <= not(layer1_outputs(4714)) or (layer1_outputs(28));
    layer2_outputs(6584) <= not(layer1_outputs(788));
    layer2_outputs(6585) <= (layer1_outputs(5950)) and not (layer1_outputs(858));
    layer2_outputs(6586) <= not((layer1_outputs(2396)) and (layer1_outputs(6008)));
    layer2_outputs(6587) <= (layer1_outputs(6038)) and not (layer1_outputs(3577));
    layer2_outputs(6588) <= layer1_outputs(5184);
    layer2_outputs(6589) <= (layer1_outputs(6022)) xor (layer1_outputs(6658));
    layer2_outputs(6590) <= layer1_outputs(6579);
    layer2_outputs(6591) <= '0';
    layer2_outputs(6592) <= not(layer1_outputs(3076)) or (layer1_outputs(6143));
    layer2_outputs(6593) <= layer1_outputs(2709);
    layer2_outputs(6594) <= not(layer1_outputs(5253));
    layer2_outputs(6595) <= (layer1_outputs(6891)) or (layer1_outputs(3398));
    layer2_outputs(6596) <= not(layer1_outputs(2469));
    layer2_outputs(6597) <= not(layer1_outputs(62)) or (layer1_outputs(3117));
    layer2_outputs(6598) <= not(layer1_outputs(4797)) or (layer1_outputs(90));
    layer2_outputs(6599) <= not(layer1_outputs(3684));
    layer2_outputs(6600) <= '0';
    layer2_outputs(6601) <= not((layer1_outputs(7413)) or (layer1_outputs(69)));
    layer2_outputs(6602) <= (layer1_outputs(1627)) or (layer1_outputs(6933));
    layer2_outputs(6603) <= (layer1_outputs(308)) or (layer1_outputs(7630));
    layer2_outputs(6604) <= not(layer1_outputs(4456));
    layer2_outputs(6605) <= not((layer1_outputs(4742)) or (layer1_outputs(5917)));
    layer2_outputs(6606) <= not(layer1_outputs(4408)) or (layer1_outputs(7609));
    layer2_outputs(6607) <= not(layer1_outputs(6673));
    layer2_outputs(6608) <= (layer1_outputs(3527)) and (layer1_outputs(4325));
    layer2_outputs(6609) <= layer1_outputs(5247);
    layer2_outputs(6610) <= '0';
    layer2_outputs(6611) <= not(layer1_outputs(596));
    layer2_outputs(6612) <= not((layer1_outputs(4500)) and (layer1_outputs(2410)));
    layer2_outputs(6613) <= not(layer1_outputs(5899));
    layer2_outputs(6614) <= not(layer1_outputs(1201)) or (layer1_outputs(6644));
    layer2_outputs(6615) <= not(layer1_outputs(5743)) or (layer1_outputs(6605));
    layer2_outputs(6616) <= not(layer1_outputs(4820));
    layer2_outputs(6617) <= '1';
    layer2_outputs(6618) <= (layer1_outputs(7009)) or (layer1_outputs(4544));
    layer2_outputs(6619) <= not(layer1_outputs(6268));
    layer2_outputs(6620) <= layer1_outputs(1920);
    layer2_outputs(6621) <= not((layer1_outputs(5817)) or (layer1_outputs(4008)));
    layer2_outputs(6622) <= not(layer1_outputs(68));
    layer2_outputs(6623) <= (layer1_outputs(6628)) or (layer1_outputs(5505));
    layer2_outputs(6624) <= layer1_outputs(1404);
    layer2_outputs(6625) <= (layer1_outputs(5335)) and not (layer1_outputs(1435));
    layer2_outputs(6626) <= not((layer1_outputs(7554)) or (layer1_outputs(3557)));
    layer2_outputs(6627) <= (layer1_outputs(7385)) and not (layer1_outputs(996));
    layer2_outputs(6628) <= not((layer1_outputs(4258)) or (layer1_outputs(1415)));
    layer2_outputs(6629) <= (layer1_outputs(5138)) and not (layer1_outputs(3511));
    layer2_outputs(6630) <= (layer1_outputs(2343)) and not (layer1_outputs(5310));
    layer2_outputs(6631) <= (layer1_outputs(6035)) and not (layer1_outputs(56));
    layer2_outputs(6632) <= '1';
    layer2_outputs(6633) <= not((layer1_outputs(6044)) and (layer1_outputs(4503)));
    layer2_outputs(6634) <= layer1_outputs(770);
    layer2_outputs(6635) <= not(layer1_outputs(6530));
    layer2_outputs(6636) <= '1';
    layer2_outputs(6637) <= not(layer1_outputs(5290)) or (layer1_outputs(1305));
    layer2_outputs(6638) <= '1';
    layer2_outputs(6639) <= '0';
    layer2_outputs(6640) <= '0';
    layer2_outputs(6641) <= not(layer1_outputs(4337));
    layer2_outputs(6642) <= (layer1_outputs(3218)) and (layer1_outputs(5926));
    layer2_outputs(6643) <= layer1_outputs(2412);
    layer2_outputs(6644) <= layer1_outputs(3207);
    layer2_outputs(6645) <= not((layer1_outputs(1822)) and (layer1_outputs(3281)));
    layer2_outputs(6646) <= '1';
    layer2_outputs(6647) <= '1';
    layer2_outputs(6648) <= not(layer1_outputs(193));
    layer2_outputs(6649) <= not(layer1_outputs(3086));
    layer2_outputs(6650) <= (layer1_outputs(3426)) or (layer1_outputs(2528));
    layer2_outputs(6651) <= not(layer1_outputs(4658)) or (layer1_outputs(1176));
    layer2_outputs(6652) <= not(layer1_outputs(5789)) or (layer1_outputs(4737));
    layer2_outputs(6653) <= '1';
    layer2_outputs(6654) <= not((layer1_outputs(7450)) xor (layer1_outputs(4014)));
    layer2_outputs(6655) <= not((layer1_outputs(5370)) and (layer1_outputs(4151)));
    layer2_outputs(6656) <= layer1_outputs(2162);
    layer2_outputs(6657) <= layer1_outputs(3225);
    layer2_outputs(6658) <= not(layer1_outputs(827)) or (layer1_outputs(5221));
    layer2_outputs(6659) <= not((layer1_outputs(5051)) or (layer1_outputs(3780)));
    layer2_outputs(6660) <= layer1_outputs(5236);
    layer2_outputs(6661) <= layer1_outputs(3611);
    layer2_outputs(6662) <= not(layer1_outputs(2201)) or (layer1_outputs(1626));
    layer2_outputs(6663) <= not(layer1_outputs(3863)) or (layer1_outputs(3280));
    layer2_outputs(6664) <= not(layer1_outputs(6641));
    layer2_outputs(6665) <= not(layer1_outputs(1427)) or (layer1_outputs(6536));
    layer2_outputs(6666) <= layer1_outputs(3443);
    layer2_outputs(6667) <= '1';
    layer2_outputs(6668) <= not(layer1_outputs(533)) or (layer1_outputs(1581));
    layer2_outputs(6669) <= (layer1_outputs(2617)) or (layer1_outputs(3020));
    layer2_outputs(6670) <= not(layer1_outputs(7487)) or (layer1_outputs(4479));
    layer2_outputs(6671) <= (layer1_outputs(2563)) or (layer1_outputs(3611));
    layer2_outputs(6672) <= '1';
    layer2_outputs(6673) <= not(layer1_outputs(4901)) or (layer1_outputs(3507));
    layer2_outputs(6674) <= (layer1_outputs(2327)) and not (layer1_outputs(1453));
    layer2_outputs(6675) <= not(layer1_outputs(3659));
    layer2_outputs(6676) <= (layer1_outputs(4336)) and not (layer1_outputs(4144));
    layer2_outputs(6677) <= not(layer1_outputs(1372));
    layer2_outputs(6678) <= layer1_outputs(929);
    layer2_outputs(6679) <= '1';
    layer2_outputs(6680) <= not(layer1_outputs(1956));
    layer2_outputs(6681) <= not((layer1_outputs(4850)) or (layer1_outputs(6255)));
    layer2_outputs(6682) <= not(layer1_outputs(2760));
    layer2_outputs(6683) <= not(layer1_outputs(3944)) or (layer1_outputs(563));
    layer2_outputs(6684) <= not(layer1_outputs(4066));
    layer2_outputs(6685) <= '0';
    layer2_outputs(6686) <= '1';
    layer2_outputs(6687) <= (layer1_outputs(6058)) or (layer1_outputs(128));
    layer2_outputs(6688) <= (layer1_outputs(7068)) or (layer1_outputs(6927));
    layer2_outputs(6689) <= '0';
    layer2_outputs(6690) <= not((layer1_outputs(7031)) or (layer1_outputs(6693)));
    layer2_outputs(6691) <= layer1_outputs(5669);
    layer2_outputs(6692) <= '1';
    layer2_outputs(6693) <= not((layer1_outputs(3814)) and (layer1_outputs(573)));
    layer2_outputs(6694) <= '0';
    layer2_outputs(6695) <= '1';
    layer2_outputs(6696) <= layer1_outputs(7123);
    layer2_outputs(6697) <= not(layer1_outputs(6627)) or (layer1_outputs(2809));
    layer2_outputs(6698) <= (layer1_outputs(1343)) and not (layer1_outputs(3740));
    layer2_outputs(6699) <= (layer1_outputs(1466)) and not (layer1_outputs(1921));
    layer2_outputs(6700) <= '1';
    layer2_outputs(6701) <= not(layer1_outputs(4090)) or (layer1_outputs(1307));
    layer2_outputs(6702) <= '1';
    layer2_outputs(6703) <= (layer1_outputs(7034)) and not (layer1_outputs(7560));
    layer2_outputs(6704) <= not(layer1_outputs(5003)) or (layer1_outputs(2812));
    layer2_outputs(6705) <= (layer1_outputs(6958)) and not (layer1_outputs(772));
    layer2_outputs(6706) <= layer1_outputs(3526);
    layer2_outputs(6707) <= '0';
    layer2_outputs(6708) <= (layer1_outputs(2166)) and not (layer1_outputs(7096));
    layer2_outputs(6709) <= not(layer1_outputs(2657)) or (layer1_outputs(6593));
    layer2_outputs(6710) <= not(layer1_outputs(6654));
    layer2_outputs(6711) <= (layer1_outputs(7433)) or (layer1_outputs(816));
    layer2_outputs(6712) <= '0';
    layer2_outputs(6713) <= (layer1_outputs(1150)) and (layer1_outputs(6355));
    layer2_outputs(6714) <= layer1_outputs(3896);
    layer2_outputs(6715) <= not(layer1_outputs(103)) or (layer1_outputs(6288));
    layer2_outputs(6716) <= not(layer1_outputs(2904));
    layer2_outputs(6717) <= not(layer1_outputs(3308)) or (layer1_outputs(1356));
    layer2_outputs(6718) <= (layer1_outputs(3867)) and not (layer1_outputs(6137));
    layer2_outputs(6719) <= layer1_outputs(7088);
    layer2_outputs(6720) <= not(layer1_outputs(5507)) or (layer1_outputs(4905));
    layer2_outputs(6721) <= '1';
    layer2_outputs(6722) <= (layer1_outputs(1486)) and (layer1_outputs(2871));
    layer2_outputs(6723) <= not(layer1_outputs(3224));
    layer2_outputs(6724) <= layer1_outputs(5173);
    layer2_outputs(6725) <= not((layer1_outputs(4233)) and (layer1_outputs(6384)));
    layer2_outputs(6726) <= '1';
    layer2_outputs(6727) <= '1';
    layer2_outputs(6728) <= (layer1_outputs(4149)) or (layer1_outputs(4420));
    layer2_outputs(6729) <= '1';
    layer2_outputs(6730) <= not(layer1_outputs(3776));
    layer2_outputs(6731) <= not(layer1_outputs(5209)) or (layer1_outputs(3433));
    layer2_outputs(6732) <= not(layer1_outputs(2772));
    layer2_outputs(6733) <= not(layer1_outputs(5333));
    layer2_outputs(6734) <= '0';
    layer2_outputs(6735) <= (layer1_outputs(163)) and (layer1_outputs(3624));
    layer2_outputs(6736) <= '0';
    layer2_outputs(6737) <= '1';
    layer2_outputs(6738) <= '0';
    layer2_outputs(6739) <= (layer1_outputs(4154)) or (layer1_outputs(4656));
    layer2_outputs(6740) <= not(layer1_outputs(6314));
    layer2_outputs(6741) <= not(layer1_outputs(5902)) or (layer1_outputs(7502));
    layer2_outputs(6742) <= not(layer1_outputs(3850)) or (layer1_outputs(2912));
    layer2_outputs(6743) <= not((layer1_outputs(1841)) or (layer1_outputs(2273)));
    layer2_outputs(6744) <= (layer1_outputs(3678)) and not (layer1_outputs(7389));
    layer2_outputs(6745) <= not(layer1_outputs(5489));
    layer2_outputs(6746) <= (layer1_outputs(4351)) or (layer1_outputs(5946));
    layer2_outputs(6747) <= not(layer1_outputs(3037)) or (layer1_outputs(626));
    layer2_outputs(6748) <= (layer1_outputs(1561)) and not (layer1_outputs(1169));
    layer2_outputs(6749) <= not(layer1_outputs(6186));
    layer2_outputs(6750) <= (layer1_outputs(2470)) and (layer1_outputs(5530));
    layer2_outputs(6751) <= (layer1_outputs(2241)) and not (layer1_outputs(7227));
    layer2_outputs(6752) <= layer1_outputs(7324);
    layer2_outputs(6753) <= (layer1_outputs(7477)) and not (layer1_outputs(1068));
    layer2_outputs(6754) <= not((layer1_outputs(6630)) or (layer1_outputs(67)));
    layer2_outputs(6755) <= not(layer1_outputs(2976));
    layer2_outputs(6756) <= not((layer1_outputs(714)) and (layer1_outputs(3480)));
    layer2_outputs(6757) <= layer1_outputs(5341);
    layer2_outputs(6758) <= (layer1_outputs(3786)) or (layer1_outputs(5475));
    layer2_outputs(6759) <= '0';
    layer2_outputs(6760) <= (layer1_outputs(2784)) and (layer1_outputs(3892));
    layer2_outputs(6761) <= (layer1_outputs(375)) or (layer1_outputs(7345));
    layer2_outputs(6762) <= not(layer1_outputs(6587));
    layer2_outputs(6763) <= not((layer1_outputs(6689)) and (layer1_outputs(681)));
    layer2_outputs(6764) <= '0';
    layer2_outputs(6765) <= not(layer1_outputs(1866));
    layer2_outputs(6766) <= not(layer1_outputs(2544)) or (layer1_outputs(4128));
    layer2_outputs(6767) <= (layer1_outputs(6105)) and not (layer1_outputs(3625));
    layer2_outputs(6768) <= (layer1_outputs(3667)) and not (layer1_outputs(1610));
    layer2_outputs(6769) <= not(layer1_outputs(3164));
    layer2_outputs(6770) <= not(layer1_outputs(2471)) or (layer1_outputs(2955));
    layer2_outputs(6771) <= layer1_outputs(514);
    layer2_outputs(6772) <= not(layer1_outputs(4357));
    layer2_outputs(6773) <= (layer1_outputs(1145)) and (layer1_outputs(2698));
    layer2_outputs(6774) <= layer1_outputs(3551);
    layer2_outputs(6775) <= layer1_outputs(5785);
    layer2_outputs(6776) <= not(layer1_outputs(5199));
    layer2_outputs(6777) <= not(layer1_outputs(817));
    layer2_outputs(6778) <= layer1_outputs(996);
    layer2_outputs(6779) <= (layer1_outputs(5661)) or (layer1_outputs(3195));
    layer2_outputs(6780) <= '0';
    layer2_outputs(6781) <= (layer1_outputs(2779)) and not (layer1_outputs(4350));
    layer2_outputs(6782) <= '0';
    layer2_outputs(6783) <= layer1_outputs(5935);
    layer2_outputs(6784) <= (layer1_outputs(1953)) and not (layer1_outputs(6259));
    layer2_outputs(6785) <= not(layer1_outputs(2695)) or (layer1_outputs(4479));
    layer2_outputs(6786) <= not(layer1_outputs(397)) or (layer1_outputs(4721));
    layer2_outputs(6787) <= (layer1_outputs(5562)) and (layer1_outputs(6042));
    layer2_outputs(6788) <= layer1_outputs(7059);
    layer2_outputs(6789) <= not((layer1_outputs(6589)) or (layer1_outputs(7013)));
    layer2_outputs(6790) <= layer1_outputs(2656);
    layer2_outputs(6791) <= layer1_outputs(2970);
    layer2_outputs(6792) <= (layer1_outputs(2034)) and (layer1_outputs(4379));
    layer2_outputs(6793) <= layer1_outputs(477);
    layer2_outputs(6794) <= not(layer1_outputs(5105));
    layer2_outputs(6795) <= not(layer1_outputs(7540));
    layer2_outputs(6796) <= not(layer1_outputs(3655));
    layer2_outputs(6797) <= (layer1_outputs(6552)) or (layer1_outputs(4593));
    layer2_outputs(6798) <= not(layer1_outputs(637)) or (layer1_outputs(4906));
    layer2_outputs(6799) <= '0';
    layer2_outputs(6800) <= not(layer1_outputs(6157));
    layer2_outputs(6801) <= not(layer1_outputs(6275));
    layer2_outputs(6802) <= '1';
    layer2_outputs(6803) <= (layer1_outputs(7620)) and (layer1_outputs(3965));
    layer2_outputs(6804) <= (layer1_outputs(126)) and not (layer1_outputs(1215));
    layer2_outputs(6805) <= not(layer1_outputs(149));
    layer2_outputs(6806) <= (layer1_outputs(1496)) xor (layer1_outputs(6166));
    layer2_outputs(6807) <= (layer1_outputs(3720)) and (layer1_outputs(4488));
    layer2_outputs(6808) <= not((layer1_outputs(7584)) or (layer1_outputs(4913)));
    layer2_outputs(6809) <= (layer1_outputs(2309)) and not (layer1_outputs(1809));
    layer2_outputs(6810) <= not(layer1_outputs(5326));
    layer2_outputs(6811) <= layer1_outputs(7282);
    layer2_outputs(6812) <= '1';
    layer2_outputs(6813) <= not((layer1_outputs(7602)) and (layer1_outputs(6215)));
    layer2_outputs(6814) <= '0';
    layer2_outputs(6815) <= not(layer1_outputs(3244)) or (layer1_outputs(1945));
    layer2_outputs(6816) <= layer1_outputs(904);
    layer2_outputs(6817) <= (layer1_outputs(1838)) and (layer1_outputs(2862));
    layer2_outputs(6818) <= (layer1_outputs(6912)) and not (layer1_outputs(6866));
    layer2_outputs(6819) <= not(layer1_outputs(5901));
    layer2_outputs(6820) <= '1';
    layer2_outputs(6821) <= not(layer1_outputs(4932));
    layer2_outputs(6822) <= '1';
    layer2_outputs(6823) <= not(layer1_outputs(1520));
    layer2_outputs(6824) <= not(layer1_outputs(254));
    layer2_outputs(6825) <= not(layer1_outputs(2712)) or (layer1_outputs(6707));
    layer2_outputs(6826) <= not(layer1_outputs(1595));
    layer2_outputs(6827) <= (layer1_outputs(6237)) and not (layer1_outputs(3555));
    layer2_outputs(6828) <= layer1_outputs(5079);
    layer2_outputs(6829) <= not(layer1_outputs(1290)) or (layer1_outputs(2952));
    layer2_outputs(6830) <= not(layer1_outputs(6855));
    layer2_outputs(6831) <= layer1_outputs(5657);
    layer2_outputs(6832) <= not(layer1_outputs(1542));
    layer2_outputs(6833) <= '0';
    layer2_outputs(6834) <= layer1_outputs(2290);
    layer2_outputs(6835) <= (layer1_outputs(6204)) xor (layer1_outputs(264));
    layer2_outputs(6836) <= layer1_outputs(3516);
    layer2_outputs(6837) <= '1';
    layer2_outputs(6838) <= '1';
    layer2_outputs(6839) <= (layer1_outputs(6207)) or (layer1_outputs(5569));
    layer2_outputs(6840) <= '0';
    layer2_outputs(6841) <= not(layer1_outputs(1878));
    layer2_outputs(6842) <= layer1_outputs(1201);
    layer2_outputs(6843) <= not(layer1_outputs(4503)) or (layer1_outputs(3553));
    layer2_outputs(6844) <= not(layer1_outputs(3936));
    layer2_outputs(6845) <= not(layer1_outputs(4139));
    layer2_outputs(6846) <= (layer1_outputs(1026)) and not (layer1_outputs(6505));
    layer2_outputs(6847) <= (layer1_outputs(408)) or (layer1_outputs(7616));
    layer2_outputs(6848) <= '0';
    layer2_outputs(6849) <= not(layer1_outputs(947));
    layer2_outputs(6850) <= not(layer1_outputs(7150));
    layer2_outputs(6851) <= (layer1_outputs(490)) or (layer1_outputs(5477));
    layer2_outputs(6852) <= (layer1_outputs(7370)) and not (layer1_outputs(796));
    layer2_outputs(6853) <= not(layer1_outputs(6408));
    layer2_outputs(6854) <= not(layer1_outputs(7230)) or (layer1_outputs(6137));
    layer2_outputs(6855) <= (layer1_outputs(1268)) and not (layer1_outputs(1186));
    layer2_outputs(6856) <= layer1_outputs(2649);
    layer2_outputs(6857) <= not(layer1_outputs(2577)) or (layer1_outputs(5846));
    layer2_outputs(6858) <= not((layer1_outputs(1187)) and (layer1_outputs(7544)));
    layer2_outputs(6859) <= not(layer1_outputs(742));
    layer2_outputs(6860) <= not(layer1_outputs(5263)) or (layer1_outputs(6111));
    layer2_outputs(6861) <= not(layer1_outputs(1433));
    layer2_outputs(6862) <= (layer1_outputs(2675)) or (layer1_outputs(387));
    layer2_outputs(6863) <= not((layer1_outputs(599)) and (layer1_outputs(3429)));
    layer2_outputs(6864) <= (layer1_outputs(1450)) and not (layer1_outputs(4952));
    layer2_outputs(6865) <= layer1_outputs(7099);
    layer2_outputs(6866) <= layer1_outputs(247);
    layer2_outputs(6867) <= not(layer1_outputs(4471));
    layer2_outputs(6868) <= (layer1_outputs(4882)) and (layer1_outputs(655));
    layer2_outputs(6869) <= not(layer1_outputs(4313)) or (layer1_outputs(5708));
    layer2_outputs(6870) <= not(layer1_outputs(2650));
    layer2_outputs(6871) <= not((layer1_outputs(6705)) or (layer1_outputs(3373)));
    layer2_outputs(6872) <= not((layer1_outputs(2432)) and (layer1_outputs(4780)));
    layer2_outputs(6873) <= (layer1_outputs(2313)) or (layer1_outputs(3698));
    layer2_outputs(6874) <= not(layer1_outputs(942)) or (layer1_outputs(3033));
    layer2_outputs(6875) <= not((layer1_outputs(3412)) and (layer1_outputs(7564)));
    layer2_outputs(6876) <= layer1_outputs(5877);
    layer2_outputs(6877) <= not(layer1_outputs(447)) or (layer1_outputs(5724));
    layer2_outputs(6878) <= not(layer1_outputs(5986));
    layer2_outputs(6879) <= (layer1_outputs(6112)) or (layer1_outputs(4991));
    layer2_outputs(6880) <= (layer1_outputs(7403)) or (layer1_outputs(81));
    layer2_outputs(6881) <= not(layer1_outputs(1632));
    layer2_outputs(6882) <= not((layer1_outputs(6981)) and (layer1_outputs(6724)));
    layer2_outputs(6883) <= (layer1_outputs(3575)) and not (layer1_outputs(1590));
    layer2_outputs(6884) <= '1';
    layer2_outputs(6885) <= not(layer1_outputs(3116)) or (layer1_outputs(3372));
    layer2_outputs(6886) <= '1';
    layer2_outputs(6887) <= not((layer1_outputs(3344)) or (layer1_outputs(566)));
    layer2_outputs(6888) <= (layer1_outputs(5672)) or (layer1_outputs(896));
    layer2_outputs(6889) <= not(layer1_outputs(6788)) or (layer1_outputs(1717));
    layer2_outputs(6890) <= not(layer1_outputs(7677)) or (layer1_outputs(2790));
    layer2_outputs(6891) <= not(layer1_outputs(1587)) or (layer1_outputs(1044));
    layer2_outputs(6892) <= not(layer1_outputs(55));
    layer2_outputs(6893) <= not(layer1_outputs(4125));
    layer2_outputs(6894) <= not(layer1_outputs(4837));
    layer2_outputs(6895) <= (layer1_outputs(7268)) and not (layer1_outputs(3476));
    layer2_outputs(6896) <= not((layer1_outputs(6821)) or (layer1_outputs(1207)));
    layer2_outputs(6897) <= not(layer1_outputs(6121));
    layer2_outputs(6898) <= not(layer1_outputs(4692)) or (layer1_outputs(2872));
    layer2_outputs(6899) <= '1';
    layer2_outputs(6900) <= not(layer1_outputs(4443)) or (layer1_outputs(7679));
    layer2_outputs(6901) <= layer1_outputs(3960);
    layer2_outputs(6902) <= (layer1_outputs(490)) and not (layer1_outputs(2573));
    layer2_outputs(6903) <= (layer1_outputs(7347)) and not (layer1_outputs(541));
    layer2_outputs(6904) <= (layer1_outputs(776)) and (layer1_outputs(4861));
    layer2_outputs(6905) <= layer1_outputs(6969);
    layer2_outputs(6906) <= not((layer1_outputs(4186)) and (layer1_outputs(7035)));
    layer2_outputs(6907) <= (layer1_outputs(4685)) and (layer1_outputs(6526));
    layer2_outputs(6908) <= (layer1_outputs(7101)) and (layer1_outputs(5819));
    layer2_outputs(6909) <= (layer1_outputs(2509)) and not (layer1_outputs(4281));
    layer2_outputs(6910) <= not(layer1_outputs(6834)) or (layer1_outputs(1737));
    layer2_outputs(6911) <= layer1_outputs(5396);
    layer2_outputs(6912) <= (layer1_outputs(3826)) and not (layer1_outputs(2884));
    layer2_outputs(6913) <= not((layer1_outputs(6576)) and (layer1_outputs(7563)));
    layer2_outputs(6914) <= '0';
    layer2_outputs(6915) <= (layer1_outputs(6118)) and not (layer1_outputs(7408));
    layer2_outputs(6916) <= layer1_outputs(3441);
    layer2_outputs(6917) <= not((layer1_outputs(2053)) xor (layer1_outputs(253)));
    layer2_outputs(6918) <= (layer1_outputs(4749)) and not (layer1_outputs(6955));
    layer2_outputs(6919) <= (layer1_outputs(4720)) and (layer1_outputs(3729));
    layer2_outputs(6920) <= not((layer1_outputs(3562)) and (layer1_outputs(5614)));
    layer2_outputs(6921) <= not(layer1_outputs(2691));
    layer2_outputs(6922) <= layer1_outputs(5051);
    layer2_outputs(6923) <= '0';
    layer2_outputs(6924) <= not((layer1_outputs(1552)) or (layer1_outputs(2623)));
    layer2_outputs(6925) <= (layer1_outputs(6126)) and (layer1_outputs(2827));
    layer2_outputs(6926) <= not((layer1_outputs(5211)) and (layer1_outputs(5160)));
    layer2_outputs(6927) <= layer1_outputs(6762);
    layer2_outputs(6928) <= not((layer1_outputs(2051)) or (layer1_outputs(1576)));
    layer2_outputs(6929) <= (layer1_outputs(6072)) and not (layer1_outputs(6630));
    layer2_outputs(6930) <= '0';
    layer2_outputs(6931) <= (layer1_outputs(6330)) or (layer1_outputs(1047));
    layer2_outputs(6932) <= '0';
    layer2_outputs(6933) <= (layer1_outputs(3371)) and not (layer1_outputs(1154));
    layer2_outputs(6934) <= (layer1_outputs(3986)) and not (layer1_outputs(5513));
    layer2_outputs(6935) <= not((layer1_outputs(2022)) and (layer1_outputs(7076)));
    layer2_outputs(6936) <= layer1_outputs(1536);
    layer2_outputs(6937) <= not(layer1_outputs(1030));
    layer2_outputs(6938) <= not(layer1_outputs(713));
    layer2_outputs(6939) <= not((layer1_outputs(6235)) and (layer1_outputs(7443)));
    layer2_outputs(6940) <= layer1_outputs(3901);
    layer2_outputs(6941) <= (layer1_outputs(6224)) and (layer1_outputs(3173));
    layer2_outputs(6942) <= layer1_outputs(4666);
    layer2_outputs(6943) <= not((layer1_outputs(6645)) and (layer1_outputs(6399)));
    layer2_outputs(6944) <= (layer1_outputs(5617)) and not (layer1_outputs(5113));
    layer2_outputs(6945) <= not((layer1_outputs(6931)) and (layer1_outputs(152)));
    layer2_outputs(6946) <= not(layer1_outputs(2091)) or (layer1_outputs(3983));
    layer2_outputs(6947) <= '0';
    layer2_outputs(6948) <= not(layer1_outputs(3896));
    layer2_outputs(6949) <= (layer1_outputs(1522)) or (layer1_outputs(4862));
    layer2_outputs(6950) <= layer1_outputs(6229);
    layer2_outputs(6951) <= (layer1_outputs(1836)) and not (layer1_outputs(4245));
    layer2_outputs(6952) <= not(layer1_outputs(3576));
    layer2_outputs(6953) <= not((layer1_outputs(5050)) or (layer1_outputs(6561)));
    layer2_outputs(6954) <= not(layer1_outputs(5898));
    layer2_outputs(6955) <= layer1_outputs(3733);
    layer2_outputs(6956) <= layer1_outputs(5342);
    layer2_outputs(6957) <= '1';
    layer2_outputs(6958) <= not((layer1_outputs(4408)) or (layer1_outputs(4156)));
    layer2_outputs(6959) <= '0';
    layer2_outputs(6960) <= (layer1_outputs(1183)) and not (layer1_outputs(2433));
    layer2_outputs(6961) <= not((layer1_outputs(867)) or (layer1_outputs(7291)));
    layer2_outputs(6962) <= (layer1_outputs(3461)) or (layer1_outputs(3432));
    layer2_outputs(6963) <= not(layer1_outputs(7261)) or (layer1_outputs(6080));
    layer2_outputs(6964) <= not((layer1_outputs(2792)) xor (layer1_outputs(6521)));
    layer2_outputs(6965) <= (layer1_outputs(3384)) and not (layer1_outputs(2087));
    layer2_outputs(6966) <= not(layer1_outputs(1676));
    layer2_outputs(6967) <= (layer1_outputs(2546)) and not (layer1_outputs(4116));
    layer2_outputs(6968) <= (layer1_outputs(7672)) or (layer1_outputs(2243));
    layer2_outputs(6969) <= '1';
    layer2_outputs(6970) <= not(layer1_outputs(4865)) or (layer1_outputs(7503));
    layer2_outputs(6971) <= layer1_outputs(1509);
    layer2_outputs(6972) <= (layer1_outputs(4833)) and (layer1_outputs(5194));
    layer2_outputs(6973) <= not(layer1_outputs(4312)) or (layer1_outputs(4037));
    layer2_outputs(6974) <= not((layer1_outputs(6755)) xor (layer1_outputs(278)));
    layer2_outputs(6975) <= not(layer1_outputs(3614));
    layer2_outputs(6976) <= not((layer1_outputs(7223)) and (layer1_outputs(1977)));
    layer2_outputs(6977) <= (layer1_outputs(7235)) or (layer1_outputs(1437));
    layer2_outputs(6978) <= (layer1_outputs(1986)) and not (layer1_outputs(3762));
    layer2_outputs(6979) <= (layer1_outputs(2000)) or (layer1_outputs(5934));
    layer2_outputs(6980) <= not(layer1_outputs(410)) or (layer1_outputs(1672));
    layer2_outputs(6981) <= not(layer1_outputs(3743));
    layer2_outputs(6982) <= not(layer1_outputs(2177));
    layer2_outputs(6983) <= (layer1_outputs(1967)) and (layer1_outputs(5304));
    layer2_outputs(6984) <= '1';
    layer2_outputs(6985) <= not(layer1_outputs(2745)) or (layer1_outputs(7655));
    layer2_outputs(6986) <= '0';
    layer2_outputs(6987) <= layer1_outputs(4150);
    layer2_outputs(6988) <= not(layer1_outputs(3622)) or (layer1_outputs(6336));
    layer2_outputs(6989) <= not((layer1_outputs(1020)) and (layer1_outputs(2115)));
    layer2_outputs(6990) <= (layer1_outputs(3869)) or (layer1_outputs(886));
    layer2_outputs(6991) <= not((layer1_outputs(6951)) or (layer1_outputs(987)));
    layer2_outputs(6992) <= layer1_outputs(6962);
    layer2_outputs(6993) <= not(layer1_outputs(1158));
    layer2_outputs(6994) <= layer1_outputs(6773);
    layer2_outputs(6995) <= (layer1_outputs(7577)) and not (layer1_outputs(6194));
    layer2_outputs(6996) <= (layer1_outputs(1465)) and not (layer1_outputs(2936));
    layer2_outputs(6997) <= not(layer1_outputs(920));
    layer2_outputs(6998) <= (layer1_outputs(1702)) and not (layer1_outputs(3701));
    layer2_outputs(6999) <= '1';
    layer2_outputs(7000) <= layer1_outputs(3967);
    layer2_outputs(7001) <= (layer1_outputs(4475)) or (layer1_outputs(3653));
    layer2_outputs(7002) <= (layer1_outputs(5183)) xor (layer1_outputs(6452));
    layer2_outputs(7003) <= not(layer1_outputs(4531));
    layer2_outputs(7004) <= (layer1_outputs(7231)) xor (layer1_outputs(2130));
    layer2_outputs(7005) <= '0';
    layer2_outputs(7006) <= (layer1_outputs(6261)) or (layer1_outputs(1199));
    layer2_outputs(7007) <= not(layer1_outputs(1664)) or (layer1_outputs(4860));
    layer2_outputs(7008) <= not(layer1_outputs(5416));
    layer2_outputs(7009) <= layer1_outputs(1200);
    layer2_outputs(7010) <= '0';
    layer2_outputs(7011) <= not(layer1_outputs(1700));
    layer2_outputs(7012) <= (layer1_outputs(982)) and not (layer1_outputs(351));
    layer2_outputs(7013) <= not(layer1_outputs(6106)) or (layer1_outputs(5701));
    layer2_outputs(7014) <= not(layer1_outputs(1071));
    layer2_outputs(7015) <= (layer1_outputs(2876)) and not (layer1_outputs(5244));
    layer2_outputs(7016) <= layer1_outputs(4360);
    layer2_outputs(7017) <= not((layer1_outputs(6945)) and (layer1_outputs(3718)));
    layer2_outputs(7018) <= layer1_outputs(7479);
    layer2_outputs(7019) <= not(layer1_outputs(2692));
    layer2_outputs(7020) <= not(layer1_outputs(7542));
    layer2_outputs(7021) <= not((layer1_outputs(4404)) and (layer1_outputs(1378)));
    layer2_outputs(7022) <= layer1_outputs(2271);
    layer2_outputs(7023) <= '1';
    layer2_outputs(7024) <= '1';
    layer2_outputs(7025) <= not(layer1_outputs(6940));
    layer2_outputs(7026) <= layer1_outputs(1079);
    layer2_outputs(7027) <= not(layer1_outputs(5215));
    layer2_outputs(7028) <= not(layer1_outputs(5988));
    layer2_outputs(7029) <= not(layer1_outputs(237)) or (layer1_outputs(33));
    layer2_outputs(7030) <= layer1_outputs(6412);
    layer2_outputs(7031) <= (layer1_outputs(1254)) and not (layer1_outputs(6281));
    layer2_outputs(7032) <= (layer1_outputs(1968)) and (layer1_outputs(5710));
    layer2_outputs(7033) <= '0';
    layer2_outputs(7034) <= not(layer1_outputs(3347));
    layer2_outputs(7035) <= not(layer1_outputs(4888)) or (layer1_outputs(3057));
    layer2_outputs(7036) <= '1';
    layer2_outputs(7037) <= (layer1_outputs(5581)) and not (layer1_outputs(4031));
    layer2_outputs(7038) <= not(layer1_outputs(221));
    layer2_outputs(7039) <= not(layer1_outputs(4639)) or (layer1_outputs(671));
    layer2_outputs(7040) <= not((layer1_outputs(6474)) and (layer1_outputs(7089)));
    layer2_outputs(7041) <= not(layer1_outputs(4893)) or (layer1_outputs(834));
    layer2_outputs(7042) <= (layer1_outputs(4104)) or (layer1_outputs(5522));
    layer2_outputs(7043) <= not((layer1_outputs(6457)) or (layer1_outputs(3758)));
    layer2_outputs(7044) <= not(layer1_outputs(1173));
    layer2_outputs(7045) <= not((layer1_outputs(1106)) or (layer1_outputs(2081)));
    layer2_outputs(7046) <= layer1_outputs(341);
    layer2_outputs(7047) <= (layer1_outputs(5611)) or (layer1_outputs(5429));
    layer2_outputs(7048) <= not((layer1_outputs(2077)) or (layer1_outputs(7505)));
    layer2_outputs(7049) <= layer1_outputs(5138);
    layer2_outputs(7050) <= '1';
    layer2_outputs(7051) <= layer1_outputs(4959);
    layer2_outputs(7052) <= (layer1_outputs(6407)) xor (layer1_outputs(4727));
    layer2_outputs(7053) <= not(layer1_outputs(5140));
    layer2_outputs(7054) <= layer1_outputs(3887);
    layer2_outputs(7055) <= not((layer1_outputs(6596)) or (layer1_outputs(4587)));
    layer2_outputs(7056) <= not(layer1_outputs(6038)) or (layer1_outputs(4441));
    layer2_outputs(7057) <= (layer1_outputs(1805)) and not (layer1_outputs(4735));
    layer2_outputs(7058) <= (layer1_outputs(7330)) and (layer1_outputs(3415));
    layer2_outputs(7059) <= '0';
    layer2_outputs(7060) <= (layer1_outputs(3365)) xor (layer1_outputs(3345));
    layer2_outputs(7061) <= layer1_outputs(2929);
    layer2_outputs(7062) <= not((layer1_outputs(4959)) or (layer1_outputs(1430)));
    layer2_outputs(7063) <= (layer1_outputs(4253)) and (layer1_outputs(451));
    layer2_outputs(7064) <= (layer1_outputs(6893)) or (layer1_outputs(7261));
    layer2_outputs(7065) <= (layer1_outputs(4186)) and (layer1_outputs(465));
    layer2_outputs(7066) <= not(layer1_outputs(2528)) or (layer1_outputs(6082));
    layer2_outputs(7067) <= (layer1_outputs(2235)) and not (layer1_outputs(5676));
    layer2_outputs(7068) <= '1';
    layer2_outputs(7069) <= (layer1_outputs(1742)) or (layer1_outputs(4176));
    layer2_outputs(7070) <= '1';
    layer2_outputs(7071) <= '1';
    layer2_outputs(7072) <= (layer1_outputs(2472)) and (layer1_outputs(1750));
    layer2_outputs(7073) <= not((layer1_outputs(5742)) and (layer1_outputs(3693)));
    layer2_outputs(7074) <= '1';
    layer2_outputs(7075) <= not((layer1_outputs(3342)) or (layer1_outputs(134)));
    layer2_outputs(7076) <= (layer1_outputs(3842)) and not (layer1_outputs(6896));
    layer2_outputs(7077) <= (layer1_outputs(6928)) and not (layer1_outputs(767));
    layer2_outputs(7078) <= not((layer1_outputs(494)) xor (layer1_outputs(6224)));
    layer2_outputs(7079) <= not(layer1_outputs(6197));
    layer2_outputs(7080) <= (layer1_outputs(6119)) and not (layer1_outputs(2256));
    layer2_outputs(7081) <= (layer1_outputs(980)) and not (layer1_outputs(3539));
    layer2_outputs(7082) <= not(layer1_outputs(2929));
    layer2_outputs(7083) <= (layer1_outputs(3377)) and not (layer1_outputs(5662));
    layer2_outputs(7084) <= layer1_outputs(6159);
    layer2_outputs(7085) <= not(layer1_outputs(7373));
    layer2_outputs(7086) <= not(layer1_outputs(2563));
    layer2_outputs(7087) <= not(layer1_outputs(389));
    layer2_outputs(7088) <= '1';
    layer2_outputs(7089) <= not(layer1_outputs(4269));
    layer2_outputs(7090) <= (layer1_outputs(260)) and (layer1_outputs(4332));
    layer2_outputs(7091) <= '1';
    layer2_outputs(7092) <= not(layer1_outputs(5056));
    layer2_outputs(7093) <= layer1_outputs(7548);
    layer2_outputs(7094) <= (layer1_outputs(944)) or (layer1_outputs(6920));
    layer2_outputs(7095) <= not((layer1_outputs(4487)) and (layer1_outputs(3821)));
    layer2_outputs(7096) <= (layer1_outputs(4859)) and not (layer1_outputs(2044));
    layer2_outputs(7097) <= (layer1_outputs(3707)) and not (layer1_outputs(4439));
    layer2_outputs(7098) <= not(layer1_outputs(1555)) or (layer1_outputs(5311));
    layer2_outputs(7099) <= not((layer1_outputs(2756)) and (layer1_outputs(1351)));
    layer2_outputs(7100) <= '0';
    layer2_outputs(7101) <= not(layer1_outputs(5805));
    layer2_outputs(7102) <= (layer1_outputs(5204)) or (layer1_outputs(713));
    layer2_outputs(7103) <= not(layer1_outputs(4649)) or (layer1_outputs(4642));
    layer2_outputs(7104) <= (layer1_outputs(1846)) and not (layer1_outputs(5476));
    layer2_outputs(7105) <= not((layer1_outputs(4647)) or (layer1_outputs(4553)));
    layer2_outputs(7106) <= '1';
    layer2_outputs(7107) <= not((layer1_outputs(99)) or (layer1_outputs(6583)));
    layer2_outputs(7108) <= '1';
    layer2_outputs(7109) <= '1';
    layer2_outputs(7110) <= '0';
    layer2_outputs(7111) <= layer1_outputs(1040);
    layer2_outputs(7112) <= not(layer1_outputs(5949));
    layer2_outputs(7113) <= layer1_outputs(1539);
    layer2_outputs(7114) <= (layer1_outputs(1507)) and not (layer1_outputs(586));
    layer2_outputs(7115) <= not((layer1_outputs(7045)) and (layer1_outputs(2048)));
    layer2_outputs(7116) <= not(layer1_outputs(1738));
    layer2_outputs(7117) <= not((layer1_outputs(664)) or (layer1_outputs(6122)));
    layer2_outputs(7118) <= (layer1_outputs(2183)) and not (layer1_outputs(5481));
    layer2_outputs(7119) <= (layer1_outputs(7015)) and not (layer1_outputs(2084));
    layer2_outputs(7120) <= not(layer1_outputs(6119)) or (layer1_outputs(6446));
    layer2_outputs(7121) <= not((layer1_outputs(1003)) and (layer1_outputs(5499)));
    layer2_outputs(7122) <= (layer1_outputs(642)) and not (layer1_outputs(2624));
    layer2_outputs(7123) <= not(layer1_outputs(3310)) or (layer1_outputs(6534));
    layer2_outputs(7124) <= not(layer1_outputs(5466));
    layer2_outputs(7125) <= not(layer1_outputs(1432)) or (layer1_outputs(4134));
    layer2_outputs(7126) <= layer1_outputs(2056);
    layer2_outputs(7127) <= not((layer1_outputs(4653)) or (layer1_outputs(634)));
    layer2_outputs(7128) <= not(layer1_outputs(3631));
    layer2_outputs(7129) <= (layer1_outputs(5347)) and not (layer1_outputs(3815));
    layer2_outputs(7130) <= layer1_outputs(6365);
    layer2_outputs(7131) <= (layer1_outputs(747)) xor (layer1_outputs(1145));
    layer2_outputs(7132) <= not(layer1_outputs(762));
    layer2_outputs(7133) <= layer1_outputs(2642);
    layer2_outputs(7134) <= (layer1_outputs(4603)) and not (layer1_outputs(2596));
    layer2_outputs(7135) <= not(layer1_outputs(748));
    layer2_outputs(7136) <= layer1_outputs(7463);
    layer2_outputs(7137) <= '1';
    layer2_outputs(7138) <= (layer1_outputs(6727)) and (layer1_outputs(1503));
    layer2_outputs(7139) <= layer1_outputs(4097);
    layer2_outputs(7140) <= (layer1_outputs(6682)) and not (layer1_outputs(686));
    layer2_outputs(7141) <= not(layer1_outputs(1962));
    layer2_outputs(7142) <= not(layer1_outputs(6535)) or (layer1_outputs(3920));
    layer2_outputs(7143) <= (layer1_outputs(2029)) and not (layer1_outputs(1599));
    layer2_outputs(7144) <= (layer1_outputs(1849)) and not (layer1_outputs(3923));
    layer2_outputs(7145) <= (layer1_outputs(5922)) and not (layer1_outputs(880));
    layer2_outputs(7146) <= not(layer1_outputs(1256)) or (layer1_outputs(1684));
    layer2_outputs(7147) <= '0';
    layer2_outputs(7148) <= (layer1_outputs(2957)) and (layer1_outputs(3198));
    layer2_outputs(7149) <= (layer1_outputs(2916)) and not (layer1_outputs(3704));
    layer2_outputs(7150) <= (layer1_outputs(2721)) and not (layer1_outputs(6379));
    layer2_outputs(7151) <= (layer1_outputs(2501)) and not (layer1_outputs(4418));
    layer2_outputs(7152) <= (layer1_outputs(2608)) or (layer1_outputs(4984));
    layer2_outputs(7153) <= layer1_outputs(5602);
    layer2_outputs(7154) <= '0';
    layer2_outputs(7155) <= layer1_outputs(7249);
    layer2_outputs(7156) <= '0';
    layer2_outputs(7157) <= layer1_outputs(1654);
    layer2_outputs(7158) <= '0';
    layer2_outputs(7159) <= not(layer1_outputs(508));
    layer2_outputs(7160) <= not((layer1_outputs(7624)) and (layer1_outputs(4914)));
    layer2_outputs(7161) <= layer1_outputs(5691);
    layer2_outputs(7162) <= not(layer1_outputs(7578));
    layer2_outputs(7163) <= not(layer1_outputs(4136)) or (layer1_outputs(836));
    layer2_outputs(7164) <= not(layer1_outputs(7269));
    layer2_outputs(7165) <= not((layer1_outputs(1766)) or (layer1_outputs(5533)));
    layer2_outputs(7166) <= not((layer1_outputs(3491)) or (layer1_outputs(6340)));
    layer2_outputs(7167) <= (layer1_outputs(6528)) or (layer1_outputs(884));
    layer2_outputs(7168) <= '1';
    layer2_outputs(7169) <= (layer1_outputs(2276)) and not (layer1_outputs(7569));
    layer2_outputs(7170) <= (layer1_outputs(4494)) and not (layer1_outputs(6660));
    layer2_outputs(7171) <= not((layer1_outputs(7346)) or (layer1_outputs(6143)));
    layer2_outputs(7172) <= not(layer1_outputs(6161));
    layer2_outputs(7173) <= '0';
    layer2_outputs(7174) <= not(layer1_outputs(5513));
    layer2_outputs(7175) <= not(layer1_outputs(2906));
    layer2_outputs(7176) <= '1';
    layer2_outputs(7177) <= not((layer1_outputs(5479)) or (layer1_outputs(6998)));
    layer2_outputs(7178) <= (layer1_outputs(5179)) and not (layer1_outputs(569));
    layer2_outputs(7179) <= not((layer1_outputs(7318)) and (layer1_outputs(1458)));
    layer2_outputs(7180) <= not(layer1_outputs(3431));
    layer2_outputs(7181) <= not(layer1_outputs(935)) or (layer1_outputs(5766));
    layer2_outputs(7182) <= not(layer1_outputs(1856));
    layer2_outputs(7183) <= layer1_outputs(1395);
    layer2_outputs(7184) <= not(layer1_outputs(5739));
    layer2_outputs(7185) <= not(layer1_outputs(4858));
    layer2_outputs(7186) <= layer1_outputs(2977);
    layer2_outputs(7187) <= '0';
    layer2_outputs(7188) <= not(layer1_outputs(6188)) or (layer1_outputs(5656));
    layer2_outputs(7189) <= not(layer1_outputs(6004));
    layer2_outputs(7190) <= not(layer1_outputs(5576)) or (layer1_outputs(4028));
    layer2_outputs(7191) <= layer1_outputs(309);
    layer2_outputs(7192) <= not(layer1_outputs(2755)) or (layer1_outputs(7435));
    layer2_outputs(7193) <= '0';
    layer2_outputs(7194) <= not(layer1_outputs(517));
    layer2_outputs(7195) <= not((layer1_outputs(1248)) and (layer1_outputs(3097)));
    layer2_outputs(7196) <= layer1_outputs(6133);
    layer2_outputs(7197) <= '0';
    layer2_outputs(7198) <= not(layer1_outputs(2950));
    layer2_outputs(7199) <= not(layer1_outputs(2092));
    layer2_outputs(7200) <= not(layer1_outputs(1178)) or (layer1_outputs(3647));
    layer2_outputs(7201) <= '1';
    layer2_outputs(7202) <= not(layer1_outputs(4229));
    layer2_outputs(7203) <= not(layer1_outputs(4873)) or (layer1_outputs(3738));
    layer2_outputs(7204) <= not(layer1_outputs(7186)) or (layer1_outputs(424));
    layer2_outputs(7205) <= layer1_outputs(189);
    layer2_outputs(7206) <= (layer1_outputs(4463)) and not (layer1_outputs(5265));
    layer2_outputs(7207) <= layer1_outputs(2031);
    layer2_outputs(7208) <= (layer1_outputs(7191)) and not (layer1_outputs(7318));
    layer2_outputs(7209) <= (layer1_outputs(5017)) xor (layer1_outputs(4350));
    layer2_outputs(7210) <= (layer1_outputs(1034)) and not (layer1_outputs(1651));
    layer2_outputs(7211) <= (layer1_outputs(3830)) and (layer1_outputs(1613));
    layer2_outputs(7212) <= not(layer1_outputs(6217)) or (layer1_outputs(3947));
    layer2_outputs(7213) <= (layer1_outputs(3634)) and not (layer1_outputs(808));
    layer2_outputs(7214) <= (layer1_outputs(6243)) and not (layer1_outputs(2617));
    layer2_outputs(7215) <= not(layer1_outputs(5769)) or (layer1_outputs(971));
    layer2_outputs(7216) <= not(layer1_outputs(3319));
    layer2_outputs(7217) <= layer1_outputs(5995);
    layer2_outputs(7218) <= (layer1_outputs(2505)) and not (layer1_outputs(3284));
    layer2_outputs(7219) <= not(layer1_outputs(1950));
    layer2_outputs(7220) <= not(layer1_outputs(7269));
    layer2_outputs(7221) <= (layer1_outputs(416)) and not (layer1_outputs(950));
    layer2_outputs(7222) <= '1';
    layer2_outputs(7223) <= not((layer1_outputs(5237)) and (layer1_outputs(4650)));
    layer2_outputs(7224) <= not((layer1_outputs(3840)) and (layer1_outputs(5705)));
    layer2_outputs(7225) <= not(layer1_outputs(815));
    layer2_outputs(7226) <= layer1_outputs(316);
    layer2_outputs(7227) <= (layer1_outputs(702)) or (layer1_outputs(1323));
    layer2_outputs(7228) <= (layer1_outputs(6597)) and not (layer1_outputs(2927));
    layer2_outputs(7229) <= (layer1_outputs(5941)) and not (layer1_outputs(4717));
    layer2_outputs(7230) <= (layer1_outputs(7523)) and not (layer1_outputs(7204));
    layer2_outputs(7231) <= '0';
    layer2_outputs(7232) <= '1';
    layer2_outputs(7233) <= not(layer1_outputs(590)) or (layer1_outputs(6892));
    layer2_outputs(7234) <= '0';
    layer2_outputs(7235) <= (layer1_outputs(6184)) and (layer1_outputs(6639));
    layer2_outputs(7236) <= (layer1_outputs(3066)) xor (layer1_outputs(4784));
    layer2_outputs(7237) <= layer1_outputs(7506);
    layer2_outputs(7238) <= (layer1_outputs(6179)) and not (layer1_outputs(6519));
    layer2_outputs(7239) <= not((layer1_outputs(7234)) or (layer1_outputs(1634)));
    layer2_outputs(7240) <= layer1_outputs(60);
    layer2_outputs(7241) <= not((layer1_outputs(5402)) or (layer1_outputs(5142)));
    layer2_outputs(7242) <= '0';
    layer2_outputs(7243) <= layer1_outputs(3849);
    layer2_outputs(7244) <= not(layer1_outputs(5607));
    layer2_outputs(7245) <= layer1_outputs(1555);
    layer2_outputs(7246) <= not(layer1_outputs(3067)) or (layer1_outputs(1566));
    layer2_outputs(7247) <= (layer1_outputs(6652)) and (layer1_outputs(2096));
    layer2_outputs(7248) <= (layer1_outputs(625)) and (layer1_outputs(3526));
    layer2_outputs(7249) <= not(layer1_outputs(4146));
    layer2_outputs(7250) <= '1';
    layer2_outputs(7251) <= '0';
    layer2_outputs(7252) <= '0';
    layer2_outputs(7253) <= '0';
    layer2_outputs(7254) <= layer1_outputs(7308);
    layer2_outputs(7255) <= '0';
    layer2_outputs(7256) <= not(layer1_outputs(7115));
    layer2_outputs(7257) <= (layer1_outputs(4619)) and not (layer1_outputs(5318));
    layer2_outputs(7258) <= (layer1_outputs(5282)) and (layer1_outputs(2150));
    layer2_outputs(7259) <= not((layer1_outputs(3004)) or (layer1_outputs(2483)));
    layer2_outputs(7260) <= '1';
    layer2_outputs(7261) <= not(layer1_outputs(5376)) or (layer1_outputs(5295));
    layer2_outputs(7262) <= not(layer1_outputs(7111));
    layer2_outputs(7263) <= not(layer1_outputs(3283)) or (layer1_outputs(5753));
    layer2_outputs(7264) <= (layer1_outputs(5810)) and not (layer1_outputs(518));
    layer2_outputs(7265) <= not(layer1_outputs(6061)) or (layer1_outputs(7169));
    layer2_outputs(7266) <= not((layer1_outputs(7392)) or (layer1_outputs(662)));
    layer2_outputs(7267) <= (layer1_outputs(787)) or (layer1_outputs(6439));
    layer2_outputs(7268) <= '0';
    layer2_outputs(7269) <= not(layer1_outputs(5521)) or (layer1_outputs(7038));
    layer2_outputs(7270) <= (layer1_outputs(6412)) and not (layer1_outputs(1663));
    layer2_outputs(7271) <= not(layer1_outputs(4960));
    layer2_outputs(7272) <= '0';
    layer2_outputs(7273) <= not(layer1_outputs(3697));
    layer2_outputs(7274) <= '1';
    layer2_outputs(7275) <= (layer1_outputs(1322)) or (layer1_outputs(4472));
    layer2_outputs(7276) <= '1';
    layer2_outputs(7277) <= layer1_outputs(2774);
    layer2_outputs(7278) <= not(layer1_outputs(5898));
    layer2_outputs(7279) <= not(layer1_outputs(1284));
    layer2_outputs(7280) <= not(layer1_outputs(6007));
    layer2_outputs(7281) <= (layer1_outputs(0)) and (layer1_outputs(2354));
    layer2_outputs(7282) <= '0';
    layer2_outputs(7283) <= '0';
    layer2_outputs(7284) <= not((layer1_outputs(711)) or (layer1_outputs(6159)));
    layer2_outputs(7285) <= not(layer1_outputs(6825)) or (layer1_outputs(2737));
    layer2_outputs(7286) <= not(layer1_outputs(2542)) or (layer1_outputs(3705));
    layer2_outputs(7287) <= not(layer1_outputs(454));
    layer2_outputs(7288) <= not(layer1_outputs(1290));
    layer2_outputs(7289) <= layer1_outputs(2622);
    layer2_outputs(7290) <= not(layer1_outputs(5440));
    layer2_outputs(7291) <= not(layer1_outputs(3559)) or (layer1_outputs(6363));
    layer2_outputs(7292) <= not(layer1_outputs(7062));
    layer2_outputs(7293) <= not((layer1_outputs(1297)) xor (layer1_outputs(4971)));
    layer2_outputs(7294) <= (layer1_outputs(4537)) and (layer1_outputs(5817));
    layer2_outputs(7295) <= not((layer1_outputs(3333)) and (layer1_outputs(6331)));
    layer2_outputs(7296) <= (layer1_outputs(2175)) and (layer1_outputs(5121));
    layer2_outputs(7297) <= layer1_outputs(869);
    layer2_outputs(7298) <= '0';
    layer2_outputs(7299) <= '1';
    layer2_outputs(7300) <= not(layer1_outputs(2473));
    layer2_outputs(7301) <= '1';
    layer2_outputs(7302) <= (layer1_outputs(7591)) and not (layer1_outputs(3064));
    layer2_outputs(7303) <= '0';
    layer2_outputs(7304) <= layer1_outputs(5966);
    layer2_outputs(7305) <= (layer1_outputs(4813)) or (layer1_outputs(1478));
    layer2_outputs(7306) <= '0';
    layer2_outputs(7307) <= layer1_outputs(2080);
    layer2_outputs(7308) <= not(layer1_outputs(873)) or (layer1_outputs(5682));
    layer2_outputs(7309) <= not(layer1_outputs(7483)) or (layer1_outputs(830));
    layer2_outputs(7310) <= not(layer1_outputs(3177));
    layer2_outputs(7311) <= not((layer1_outputs(440)) and (layer1_outputs(3286)));
    layer2_outputs(7312) <= (layer1_outputs(4469)) or (layer1_outputs(7116));
    layer2_outputs(7313) <= not(layer1_outputs(7106)) or (layer1_outputs(5360));
    layer2_outputs(7314) <= (layer1_outputs(7030)) and not (layer1_outputs(3636));
    layer2_outputs(7315) <= (layer1_outputs(2707)) or (layer1_outputs(6727));
    layer2_outputs(7316) <= (layer1_outputs(2154)) and not (layer1_outputs(1906));
    layer2_outputs(7317) <= not(layer1_outputs(2765)) or (layer1_outputs(6711));
    layer2_outputs(7318) <= (layer1_outputs(5052)) and not (layer1_outputs(3542));
    layer2_outputs(7319) <= '0';
    layer2_outputs(7320) <= (layer1_outputs(3916)) and (layer1_outputs(6098));
    layer2_outputs(7321) <= (layer1_outputs(5277)) and not (layer1_outputs(6162));
    layer2_outputs(7322) <= (layer1_outputs(6154)) and not (layer1_outputs(439));
    layer2_outputs(7323) <= (layer1_outputs(3320)) and not (layer1_outputs(1914));
    layer2_outputs(7324) <= layer1_outputs(611);
    layer2_outputs(7325) <= '1';
    layer2_outputs(7326) <= (layer1_outputs(4104)) and (layer1_outputs(5036));
    layer2_outputs(7327) <= layer1_outputs(5575);
    layer2_outputs(7328) <= (layer1_outputs(531)) and (layer1_outputs(247));
    layer2_outputs(7329) <= not(layer1_outputs(2010)) or (layer1_outputs(388));
    layer2_outputs(7330) <= not(layer1_outputs(5561));
    layer2_outputs(7331) <= (layer1_outputs(6120)) and not (layer1_outputs(2835));
    layer2_outputs(7332) <= not(layer1_outputs(1677)) or (layer1_outputs(5203));
    layer2_outputs(7333) <= '1';
    layer2_outputs(7334) <= layer1_outputs(855);
    layer2_outputs(7335) <= layer1_outputs(6101);
    layer2_outputs(7336) <= not((layer1_outputs(5530)) or (layer1_outputs(4742)));
    layer2_outputs(7337) <= not(layer1_outputs(5600)) or (layer1_outputs(4729));
    layer2_outputs(7338) <= not((layer1_outputs(7470)) or (layer1_outputs(7113)));
    layer2_outputs(7339) <= not(layer1_outputs(5841));
    layer2_outputs(7340) <= not(layer1_outputs(5196)) or (layer1_outputs(1788));
    layer2_outputs(7341) <= '1';
    layer2_outputs(7342) <= not(layer1_outputs(2945));
    layer2_outputs(7343) <= not(layer1_outputs(7262)) or (layer1_outputs(4042));
    layer2_outputs(7344) <= not((layer1_outputs(3024)) xor (layer1_outputs(3860)));
    layer2_outputs(7345) <= not((layer1_outputs(324)) and (layer1_outputs(1693)));
    layer2_outputs(7346) <= '0';
    layer2_outputs(7347) <= layer1_outputs(1755);
    layer2_outputs(7348) <= layer1_outputs(1557);
    layer2_outputs(7349) <= '1';
    layer2_outputs(7350) <= layer1_outputs(2080);
    layer2_outputs(7351) <= (layer1_outputs(588)) or (layer1_outputs(736));
    layer2_outputs(7352) <= (layer1_outputs(2963)) and not (layer1_outputs(5468));
    layer2_outputs(7353) <= not(layer1_outputs(5529));
    layer2_outputs(7354) <= '0';
    layer2_outputs(7355) <= not((layer1_outputs(4947)) xor (layer1_outputs(1181)));
    layer2_outputs(7356) <= layer1_outputs(6678);
    layer2_outputs(7357) <= (layer1_outputs(1849)) or (layer1_outputs(3282));
    layer2_outputs(7358) <= layer1_outputs(5511);
    layer2_outputs(7359) <= (layer1_outputs(970)) or (layer1_outputs(5695));
    layer2_outputs(7360) <= not((layer1_outputs(7485)) or (layer1_outputs(2348)));
    layer2_outputs(7361) <= not(layer1_outputs(5708)) or (layer1_outputs(2556));
    layer2_outputs(7362) <= layer1_outputs(6469);
    layer2_outputs(7363) <= layer1_outputs(7605);
    layer2_outputs(7364) <= (layer1_outputs(3440)) and not (layer1_outputs(958));
    layer2_outputs(7365) <= (layer1_outputs(3988)) and (layer1_outputs(1908));
    layer2_outputs(7366) <= (layer1_outputs(6862)) and not (layer1_outputs(7206));
    layer2_outputs(7367) <= (layer1_outputs(1716)) and not (layer1_outputs(2135));
    layer2_outputs(7368) <= layer1_outputs(4810);
    layer2_outputs(7369) <= not(layer1_outputs(1283));
    layer2_outputs(7370) <= not(layer1_outputs(2151));
    layer2_outputs(7371) <= (layer1_outputs(2090)) and not (layer1_outputs(6359));
    layer2_outputs(7372) <= not(layer1_outputs(2355)) or (layer1_outputs(1521));
    layer2_outputs(7373) <= not(layer1_outputs(2098));
    layer2_outputs(7374) <= not((layer1_outputs(5493)) and (layer1_outputs(32)));
    layer2_outputs(7375) <= layer1_outputs(2813);
    layer2_outputs(7376) <= not(layer1_outputs(1280)) or (layer1_outputs(3551));
    layer2_outputs(7377) <= not(layer1_outputs(2577));
    layer2_outputs(7378) <= (layer1_outputs(3690)) and (layer1_outputs(2379));
    layer2_outputs(7379) <= '1';
    layer2_outputs(7380) <= layer1_outputs(2400);
    layer2_outputs(7381) <= not(layer1_outputs(1980));
    layer2_outputs(7382) <= not((layer1_outputs(3966)) and (layer1_outputs(1976)));
    layer2_outputs(7383) <= not(layer1_outputs(7117)) or (layer1_outputs(1138));
    layer2_outputs(7384) <= not(layer1_outputs(5038));
    layer2_outputs(7385) <= (layer1_outputs(5063)) and not (layer1_outputs(6239));
    layer2_outputs(7386) <= (layer1_outputs(6055)) and not (layer1_outputs(379));
    layer2_outputs(7387) <= not(layer1_outputs(6424)) or (layer1_outputs(607));
    layer2_outputs(7388) <= '1';
    layer2_outputs(7389) <= (layer1_outputs(642)) and (layer1_outputs(5409));
    layer2_outputs(7390) <= '0';
    layer2_outputs(7391) <= not(layer1_outputs(3658)) or (layer1_outputs(3408));
    layer2_outputs(7392) <= (layer1_outputs(3801)) or (layer1_outputs(5974));
    layer2_outputs(7393) <= not((layer1_outputs(5422)) or (layer1_outputs(6021)));
    layer2_outputs(7394) <= not(layer1_outputs(1357));
    layer2_outputs(7395) <= not((layer1_outputs(5842)) or (layer1_outputs(3751)));
    layer2_outputs(7396) <= not(layer1_outputs(4546));
    layer2_outputs(7397) <= (layer1_outputs(2592)) or (layer1_outputs(7454));
    layer2_outputs(7398) <= layer1_outputs(4439);
    layer2_outputs(7399) <= '0';
    layer2_outputs(7400) <= (layer1_outputs(5296)) or (layer1_outputs(1594));
    layer2_outputs(7401) <= not((layer1_outputs(6671)) or (layer1_outputs(4526)));
    layer2_outputs(7402) <= (layer1_outputs(1570)) and not (layer1_outputs(6029));
    layer2_outputs(7403) <= (layer1_outputs(5857)) and (layer1_outputs(6257));
    layer2_outputs(7404) <= '1';
    layer2_outputs(7405) <= not(layer1_outputs(4327)) or (layer1_outputs(774));
    layer2_outputs(7406) <= '0';
    layer2_outputs(7407) <= (layer1_outputs(242)) and not (layer1_outputs(6950));
    layer2_outputs(7408) <= '0';
    layer2_outputs(7409) <= (layer1_outputs(6687)) and not (layer1_outputs(6460));
    layer2_outputs(7410) <= not(layer1_outputs(6559));
    layer2_outputs(7411) <= not(layer1_outputs(401));
    layer2_outputs(7412) <= (layer1_outputs(3449)) and not (layer1_outputs(5814));
    layer2_outputs(7413) <= layer1_outputs(960);
    layer2_outputs(7414) <= not((layer1_outputs(5254)) and (layer1_outputs(6228)));
    layer2_outputs(7415) <= not(layer1_outputs(3258)) or (layer1_outputs(230));
    layer2_outputs(7416) <= not(layer1_outputs(991)) or (layer1_outputs(733));
    layer2_outputs(7417) <= '0';
    layer2_outputs(7418) <= layer1_outputs(1375);
    layer2_outputs(7419) <= layer1_outputs(6150);
    layer2_outputs(7420) <= (layer1_outputs(2115)) or (layer1_outputs(2867));
    layer2_outputs(7421) <= not(layer1_outputs(2798));
    layer2_outputs(7422) <= layer1_outputs(5888);
    layer2_outputs(7423) <= layer1_outputs(1249);
    layer2_outputs(7424) <= not(layer1_outputs(720)) or (layer1_outputs(2498));
    layer2_outputs(7425) <= layer1_outputs(5725);
    layer2_outputs(7426) <= (layer1_outputs(3582)) and (layer1_outputs(1118));
    layer2_outputs(7427) <= not(layer1_outputs(4147));
    layer2_outputs(7428) <= not((layer1_outputs(2997)) or (layer1_outputs(4739)));
    layer2_outputs(7429) <= not(layer1_outputs(3063));
    layer2_outputs(7430) <= (layer1_outputs(4665)) or (layer1_outputs(6565));
    layer2_outputs(7431) <= layer1_outputs(1250);
    layer2_outputs(7432) <= not(layer1_outputs(2855)) or (layer1_outputs(1481));
    layer2_outputs(7433) <= '1';
    layer2_outputs(7434) <= (layer1_outputs(6212)) or (layer1_outputs(4298));
    layer2_outputs(7435) <= not(layer1_outputs(6750)) or (layer1_outputs(1164));
    layer2_outputs(7436) <= layer1_outputs(6526);
    layer2_outputs(7437) <= (layer1_outputs(6466)) and not (layer1_outputs(5500));
    layer2_outputs(7438) <= layer1_outputs(3684);
    layer2_outputs(7439) <= '1';
    layer2_outputs(7440) <= not(layer1_outputs(3343));
    layer2_outputs(7441) <= not((layer1_outputs(6212)) or (layer1_outputs(7446)));
    layer2_outputs(7442) <= '0';
    layer2_outputs(7443) <= layer1_outputs(495);
    layer2_outputs(7444) <= not(layer1_outputs(5077)) or (layer1_outputs(599));
    layer2_outputs(7445) <= layer1_outputs(1021);
    layer2_outputs(7446) <= not(layer1_outputs(1797)) or (layer1_outputs(3393));
    layer2_outputs(7447) <= '1';
    layer2_outputs(7448) <= not((layer1_outputs(1569)) and (layer1_outputs(6297)));
    layer2_outputs(7449) <= (layer1_outputs(5847)) or (layer1_outputs(825));
    layer2_outputs(7450) <= layer1_outputs(1595);
    layer2_outputs(7451) <= '0';
    layer2_outputs(7452) <= (layer1_outputs(7287)) and not (layer1_outputs(6636));
    layer2_outputs(7453) <= (layer1_outputs(4486)) and not (layer1_outputs(6037));
    layer2_outputs(7454) <= not(layer1_outputs(3369)) or (layer1_outputs(911));
    layer2_outputs(7455) <= not(layer1_outputs(3903)) or (layer1_outputs(89));
    layer2_outputs(7456) <= '1';
    layer2_outputs(7457) <= not(layer1_outputs(7043));
    layer2_outputs(7458) <= (layer1_outputs(194)) and not (layer1_outputs(2247));
    layer2_outputs(7459) <= (layer1_outputs(1899)) or (layer1_outputs(5680));
    layer2_outputs(7460) <= not(layer1_outputs(7470));
    layer2_outputs(7461) <= not(layer1_outputs(1151)) or (layer1_outputs(7357));
    layer2_outputs(7462) <= layer1_outputs(5083);
    layer2_outputs(7463) <= (layer1_outputs(5822)) or (layer1_outputs(5961));
    layer2_outputs(7464) <= layer1_outputs(4726);
    layer2_outputs(7465) <= not(layer1_outputs(4321)) or (layer1_outputs(6428));
    layer2_outputs(7466) <= (layer1_outputs(2667)) or (layer1_outputs(1091));
    layer2_outputs(7467) <= (layer1_outputs(655)) and not (layer1_outputs(2822));
    layer2_outputs(7468) <= not((layer1_outputs(1442)) or (layer1_outputs(5621)));
    layer2_outputs(7469) <= '0';
    layer2_outputs(7470) <= not((layer1_outputs(6295)) and (layer1_outputs(7225)));
    layer2_outputs(7471) <= not((layer1_outputs(5996)) and (layer1_outputs(160)));
    layer2_outputs(7472) <= (layer1_outputs(4285)) or (layer1_outputs(3503));
    layer2_outputs(7473) <= not(layer1_outputs(7594));
    layer2_outputs(7474) <= (layer1_outputs(2824)) or (layer1_outputs(2250));
    layer2_outputs(7475) <= not((layer1_outputs(6581)) and (layer1_outputs(5685)));
    layer2_outputs(7476) <= '1';
    layer2_outputs(7477) <= not(layer1_outputs(6614)) or (layer1_outputs(1774));
    layer2_outputs(7478) <= not((layer1_outputs(3921)) or (layer1_outputs(7468)));
    layer2_outputs(7479) <= not(layer1_outputs(424)) or (layer1_outputs(2045));
    layer2_outputs(7480) <= not(layer1_outputs(1485));
    layer2_outputs(7481) <= not((layer1_outputs(731)) xor (layer1_outputs(2644)));
    layer2_outputs(7482) <= (layer1_outputs(2506)) and not (layer1_outputs(1518));
    layer2_outputs(7483) <= layer1_outputs(1669);
    layer2_outputs(7484) <= (layer1_outputs(3457)) and (layer1_outputs(1014));
    layer2_outputs(7485) <= not(layer1_outputs(5043)) or (layer1_outputs(4824));
    layer2_outputs(7486) <= layer1_outputs(5874);
    layer2_outputs(7487) <= layer1_outputs(946);
    layer2_outputs(7488) <= not(layer1_outputs(2760));
    layer2_outputs(7489) <= not(layer1_outputs(5962)) or (layer1_outputs(3161));
    layer2_outputs(7490) <= not(layer1_outputs(5002)) or (layer1_outputs(2746));
    layer2_outputs(7491) <= (layer1_outputs(5432)) and not (layer1_outputs(462));
    layer2_outputs(7492) <= layer1_outputs(5112);
    layer2_outputs(7493) <= '0';
    layer2_outputs(7494) <= not((layer1_outputs(870)) or (layer1_outputs(1264)));
    layer2_outputs(7495) <= (layer1_outputs(6028)) and (layer1_outputs(209));
    layer2_outputs(7496) <= not(layer1_outputs(4520));
    layer2_outputs(7497) <= not(layer1_outputs(3606));
    layer2_outputs(7498) <= not(layer1_outputs(3274));
    layer2_outputs(7499) <= not(layer1_outputs(5797)) or (layer1_outputs(5151));
    layer2_outputs(7500) <= '0';
    layer2_outputs(7501) <= (layer1_outputs(366)) or (layer1_outputs(6030));
    layer2_outputs(7502) <= not(layer1_outputs(3520));
    layer2_outputs(7503) <= not((layer1_outputs(113)) or (layer1_outputs(6914)));
    layer2_outputs(7504) <= not(layer1_outputs(4726)) or (layer1_outputs(4391));
    layer2_outputs(7505) <= layer1_outputs(6323);
    layer2_outputs(7506) <= (layer1_outputs(5872)) and not (layer1_outputs(7618));
    layer2_outputs(7507) <= not(layer1_outputs(6580)) or (layer1_outputs(1227));
    layer2_outputs(7508) <= layer1_outputs(4169);
    layer2_outputs(7509) <= not(layer1_outputs(167));
    layer2_outputs(7510) <= not(layer1_outputs(2409));
    layer2_outputs(7511) <= (layer1_outputs(1772)) and (layer1_outputs(5913));
    layer2_outputs(7512) <= layer1_outputs(5803);
    layer2_outputs(7513) <= (layer1_outputs(2226)) xor (layer1_outputs(4562));
    layer2_outputs(7514) <= (layer1_outputs(7250)) and not (layer1_outputs(607));
    layer2_outputs(7515) <= (layer1_outputs(269)) and not (layer1_outputs(6301));
    layer2_outputs(7516) <= layer1_outputs(3378);
    layer2_outputs(7517) <= '0';
    layer2_outputs(7518) <= layer1_outputs(5230);
    layer2_outputs(7519) <= not(layer1_outputs(663));
    layer2_outputs(7520) <= '1';
    layer2_outputs(7521) <= (layer1_outputs(6027)) and not (layer1_outputs(5727));
    layer2_outputs(7522) <= '0';
    layer2_outputs(7523) <= not(layer1_outputs(209)) or (layer1_outputs(6792));
    layer2_outputs(7524) <= (layer1_outputs(6629)) and not (layer1_outputs(4011));
    layer2_outputs(7525) <= layer1_outputs(644);
    layer2_outputs(7526) <= (layer1_outputs(6841)) or (layer1_outputs(919));
    layer2_outputs(7527) <= '1';
    layer2_outputs(7528) <= (layer1_outputs(4883)) and not (layer1_outputs(5361));
    layer2_outputs(7529) <= not(layer1_outputs(1084)) or (layer1_outputs(4899));
    layer2_outputs(7530) <= '1';
    layer2_outputs(7531) <= (layer1_outputs(2483)) and not (layer1_outputs(7466));
    layer2_outputs(7532) <= not(layer1_outputs(3530));
    layer2_outputs(7533) <= layer1_outputs(3122);
    layer2_outputs(7534) <= (layer1_outputs(3847)) and (layer1_outputs(1423));
    layer2_outputs(7535) <= (layer1_outputs(5533)) and (layer1_outputs(698));
    layer2_outputs(7536) <= layer1_outputs(6199);
    layer2_outputs(7537) <= layer1_outputs(4623);
    layer2_outputs(7538) <= not((layer1_outputs(2550)) or (layer1_outputs(3948)));
    layer2_outputs(7539) <= (layer1_outputs(1123)) and not (layer1_outputs(6862));
    layer2_outputs(7540) <= (layer1_outputs(7092)) and not (layer1_outputs(263));
    layer2_outputs(7541) <= layer1_outputs(4532);
    layer2_outputs(7542) <= (layer1_outputs(5747)) and not (layer1_outputs(4292));
    layer2_outputs(7543) <= layer1_outputs(4908);
    layer2_outputs(7544) <= '0';
    layer2_outputs(7545) <= '1';
    layer2_outputs(7546) <= not(layer1_outputs(3080)) or (layer1_outputs(5406));
    layer2_outputs(7547) <= layer1_outputs(3699);
    layer2_outputs(7548) <= not((layer1_outputs(3879)) or (layer1_outputs(1510)));
    layer2_outputs(7549) <= '0';
    layer2_outputs(7550) <= layer1_outputs(6219);
    layer2_outputs(7551) <= '0';
    layer2_outputs(7552) <= layer1_outputs(6473);
    layer2_outputs(7553) <= layer1_outputs(1601);
    layer2_outputs(7554) <= (layer1_outputs(3134)) and not (layer1_outputs(2006));
    layer2_outputs(7555) <= (layer1_outputs(635)) or (layer1_outputs(4361));
    layer2_outputs(7556) <= '0';
    layer2_outputs(7557) <= (layer1_outputs(1931)) and (layer1_outputs(4403));
    layer2_outputs(7558) <= '0';
    layer2_outputs(7559) <= '0';
    layer2_outputs(7560) <= not((layer1_outputs(2905)) or (layer1_outputs(5441)));
    layer2_outputs(7561) <= not(layer1_outputs(7525)) or (layer1_outputs(1759));
    layer2_outputs(7562) <= '1';
    layer2_outputs(7563) <= (layer1_outputs(6233)) and (layer1_outputs(1794));
    layer2_outputs(7564) <= not(layer1_outputs(1444));
    layer2_outputs(7565) <= (layer1_outputs(7314)) or (layer1_outputs(3137));
    layer2_outputs(7566) <= (layer1_outputs(5350)) and not (layer1_outputs(641));
    layer2_outputs(7567) <= layer1_outputs(182);
    layer2_outputs(7568) <= not(layer1_outputs(5428)) or (layer1_outputs(1580));
    layer2_outputs(7569) <= layer1_outputs(6007);
    layer2_outputs(7570) <= (layer1_outputs(2325)) and not (layer1_outputs(2864));
    layer2_outputs(7571) <= not(layer1_outputs(296)) or (layer1_outputs(1825));
    layer2_outputs(7572) <= not(layer1_outputs(831));
    layer2_outputs(7573) <= not(layer1_outputs(6435)) or (layer1_outputs(89));
    layer2_outputs(7574) <= not((layer1_outputs(3291)) and (layer1_outputs(4515)));
    layer2_outputs(7575) <= layer1_outputs(4798);
    layer2_outputs(7576) <= layer1_outputs(4013);
    layer2_outputs(7577) <= layer1_outputs(4782);
    layer2_outputs(7578) <= (layer1_outputs(2452)) or (layer1_outputs(5462));
    layer2_outputs(7579) <= not(layer1_outputs(4110));
    layer2_outputs(7580) <= (layer1_outputs(566)) and not (layer1_outputs(5785));
    layer2_outputs(7581) <= (layer1_outputs(7480)) and not (layer1_outputs(3424));
    layer2_outputs(7582) <= not(layer1_outputs(610));
    layer2_outputs(7583) <= not((layer1_outputs(2189)) and (layer1_outputs(2813)));
    layer2_outputs(7584) <= (layer1_outputs(2533)) xor (layer1_outputs(4245));
    layer2_outputs(7585) <= layer1_outputs(1903);
    layer2_outputs(7586) <= not(layer1_outputs(4549));
    layer2_outputs(7587) <= not((layer1_outputs(5986)) and (layer1_outputs(2917)));
    layer2_outputs(7588) <= layer1_outputs(3748);
    layer2_outputs(7589) <= (layer1_outputs(5214)) or (layer1_outputs(2160));
    layer2_outputs(7590) <= not(layer1_outputs(4189));
    layer2_outputs(7591) <= not(layer1_outputs(5175));
    layer2_outputs(7592) <= not(layer1_outputs(2513));
    layer2_outputs(7593) <= (layer1_outputs(1948)) and (layer1_outputs(4329));
    layer2_outputs(7594) <= not((layer1_outputs(552)) or (layer1_outputs(2719)));
    layer2_outputs(7595) <= not((layer1_outputs(3372)) and (layer1_outputs(1092)));
    layer2_outputs(7596) <= (layer1_outputs(3293)) and not (layer1_outputs(6118));
    layer2_outputs(7597) <= layer1_outputs(2238);
    layer2_outputs(7598) <= (layer1_outputs(1971)) and not (layer1_outputs(79));
    layer2_outputs(7599) <= (layer1_outputs(1771)) and not (layer1_outputs(604));
    layer2_outputs(7600) <= not(layer1_outputs(696));
    layer2_outputs(7601) <= not(layer1_outputs(4085));
    layer2_outputs(7602) <= '1';
    layer2_outputs(7603) <= (layer1_outputs(3843)) and not (layer1_outputs(3247));
    layer2_outputs(7604) <= (layer1_outputs(7228)) and not (layer1_outputs(81));
    layer2_outputs(7605) <= layer1_outputs(4932);
    layer2_outputs(7606) <= (layer1_outputs(2092)) and (layer1_outputs(213));
    layer2_outputs(7607) <= (layer1_outputs(3514)) and (layer1_outputs(4751));
    layer2_outputs(7608) <= '0';
    layer2_outputs(7609) <= (layer1_outputs(2699)) and not (layer1_outputs(7450));
    layer2_outputs(7610) <= '0';
    layer2_outputs(7611) <= (layer1_outputs(6246)) or (layer1_outputs(6326));
    layer2_outputs(7612) <= not(layer1_outputs(4310)) or (layer1_outputs(2425));
    layer2_outputs(7613) <= layer1_outputs(2726);
    layer2_outputs(7614) <= '0';
    layer2_outputs(7615) <= (layer1_outputs(2173)) and not (layer1_outputs(4081));
    layer2_outputs(7616) <= not(layer1_outputs(6153));
    layer2_outputs(7617) <= not(layer1_outputs(4900)) or (layer1_outputs(3462));
    layer2_outputs(7618) <= not(layer1_outputs(2658));
    layer2_outputs(7619) <= (layer1_outputs(3969)) or (layer1_outputs(5436));
    layer2_outputs(7620) <= not(layer1_outputs(6710));
    layer2_outputs(7621) <= layer1_outputs(362);
    layer2_outputs(7622) <= not(layer1_outputs(5807));
    layer2_outputs(7623) <= '1';
    layer2_outputs(7624) <= layer1_outputs(310);
    layer2_outputs(7625) <= not(layer1_outputs(555)) or (layer1_outputs(1675));
    layer2_outputs(7626) <= not((layer1_outputs(2378)) or (layer1_outputs(1395)));
    layer2_outputs(7627) <= layer1_outputs(7380);
    layer2_outputs(7628) <= not(layer1_outputs(292)) or (layer1_outputs(1890));
    layer2_outputs(7629) <= not(layer1_outputs(1605));
    layer2_outputs(7630) <= (layer1_outputs(5700)) and not (layer1_outputs(7031));
    layer2_outputs(7631) <= not((layer1_outputs(6833)) and (layer1_outputs(2227)));
    layer2_outputs(7632) <= (layer1_outputs(2668)) and not (layer1_outputs(6889));
    layer2_outputs(7633) <= layer1_outputs(1009);
    layer2_outputs(7634) <= (layer1_outputs(3141)) and not (layer1_outputs(4924));
    layer2_outputs(7635) <= '0';
    layer2_outputs(7636) <= '1';
    layer2_outputs(7637) <= (layer1_outputs(5125)) and not (layer1_outputs(2589));
    layer2_outputs(7638) <= (layer1_outputs(1909)) and (layer1_outputs(6330));
    layer2_outputs(7639) <= (layer1_outputs(5885)) and not (layer1_outputs(5418));
    layer2_outputs(7640) <= '0';
    layer2_outputs(7641) <= not((layer1_outputs(304)) or (layer1_outputs(1109)));
    layer2_outputs(7642) <= (layer1_outputs(1476)) or (layer1_outputs(1051));
    layer2_outputs(7643) <= layer1_outputs(4678);
    layer2_outputs(7644) <= not((layer1_outputs(4548)) and (layer1_outputs(3987)));
    layer2_outputs(7645) <= (layer1_outputs(2121)) and not (layer1_outputs(4864));
    layer2_outputs(7646) <= not((layer1_outputs(3323)) or (layer1_outputs(7234)));
    layer2_outputs(7647) <= '0';
    layer2_outputs(7648) <= '0';
    layer2_outputs(7649) <= not(layer1_outputs(1778));
    layer2_outputs(7650) <= '1';
    layer2_outputs(7651) <= (layer1_outputs(1855)) and (layer1_outputs(1713));
    layer2_outputs(7652) <= (layer1_outputs(232)) and not (layer1_outputs(6302));
    layer2_outputs(7653) <= not(layer1_outputs(4256));
    layer2_outputs(7654) <= not((layer1_outputs(3932)) or (layer1_outputs(4048)));
    layer2_outputs(7655) <= not(layer1_outputs(3782)) or (layer1_outputs(3591));
    layer2_outputs(7656) <= layer1_outputs(6664);
    layer2_outputs(7657) <= (layer1_outputs(1285)) and not (layer1_outputs(783));
    layer2_outputs(7658) <= not(layer1_outputs(3423)) or (layer1_outputs(4216));
    layer2_outputs(7659) <= not((layer1_outputs(5679)) and (layer1_outputs(6512)));
    layer2_outputs(7660) <= not(layer1_outputs(7145));
    layer2_outputs(7661) <= not(layer1_outputs(7426)) or (layer1_outputs(6207));
    layer2_outputs(7662) <= (layer1_outputs(327)) and not (layer1_outputs(5712));
    layer2_outputs(7663) <= (layer1_outputs(3550)) and not (layer1_outputs(5956));
    layer2_outputs(7664) <= (layer1_outputs(396)) or (layer1_outputs(5319));
    layer2_outputs(7665) <= (layer1_outputs(6999)) and (layer1_outputs(6774));
    layer2_outputs(7666) <= not(layer1_outputs(7665)) or (layer1_outputs(47));
    layer2_outputs(7667) <= (layer1_outputs(350)) and not (layer1_outputs(1711));
    layer2_outputs(7668) <= not(layer1_outputs(3112)) or (layer1_outputs(503));
    layer2_outputs(7669) <= '1';
    layer2_outputs(7670) <= not(layer1_outputs(4277)) or (layer1_outputs(3491));
    layer2_outputs(7671) <= not(layer1_outputs(3734)) or (layer1_outputs(5222));
    layer2_outputs(7672) <= not(layer1_outputs(5887));
    layer2_outputs(7673) <= not((layer1_outputs(2993)) or (layer1_outputs(248)));
    layer2_outputs(7674) <= '0';
    layer2_outputs(7675) <= layer1_outputs(4633);
    layer2_outputs(7676) <= layer1_outputs(4912);
    layer2_outputs(7677) <= '0';
    layer2_outputs(7678) <= not(layer1_outputs(2987)) or (layer1_outputs(7350));
    layer2_outputs(7679) <= not(layer1_outputs(1913)) or (layer1_outputs(956));
    layer3_outputs(0) <= (layer2_outputs(811)) or (layer2_outputs(5625));
    layer3_outputs(1) <= not((layer2_outputs(951)) or (layer2_outputs(3786)));
    layer3_outputs(2) <= not((layer2_outputs(1689)) or (layer2_outputs(5071)));
    layer3_outputs(3) <= (layer2_outputs(19)) or (layer2_outputs(7211));
    layer3_outputs(4) <= (layer2_outputs(702)) and (layer2_outputs(1708));
    layer3_outputs(5) <= not(layer2_outputs(2604));
    layer3_outputs(6) <= '1';
    layer3_outputs(7) <= '0';
    layer3_outputs(8) <= not(layer2_outputs(7185));
    layer3_outputs(9) <= not(layer2_outputs(1094)) or (layer2_outputs(2087));
    layer3_outputs(10) <= layer2_outputs(166);
    layer3_outputs(11) <= not(layer2_outputs(6098));
    layer3_outputs(12) <= not(layer2_outputs(3482)) or (layer2_outputs(1976));
    layer3_outputs(13) <= layer2_outputs(5365);
    layer3_outputs(14) <= not(layer2_outputs(6711)) or (layer2_outputs(5223));
    layer3_outputs(15) <= not((layer2_outputs(3919)) and (layer2_outputs(77)));
    layer3_outputs(16) <= (layer2_outputs(5102)) or (layer2_outputs(5069));
    layer3_outputs(17) <= (layer2_outputs(2222)) or (layer2_outputs(663));
    layer3_outputs(18) <= (layer2_outputs(3445)) and not (layer2_outputs(6603));
    layer3_outputs(19) <= not(layer2_outputs(6024));
    layer3_outputs(20) <= not((layer2_outputs(6380)) and (layer2_outputs(31)));
    layer3_outputs(21) <= layer2_outputs(6011);
    layer3_outputs(22) <= not((layer2_outputs(3936)) and (layer2_outputs(5005)));
    layer3_outputs(23) <= not(layer2_outputs(4270));
    layer3_outputs(24) <= not(layer2_outputs(6272));
    layer3_outputs(25) <= (layer2_outputs(5369)) xor (layer2_outputs(570));
    layer3_outputs(26) <= layer2_outputs(7377);
    layer3_outputs(27) <= not(layer2_outputs(5192)) or (layer2_outputs(7143));
    layer3_outputs(28) <= not(layer2_outputs(4292));
    layer3_outputs(29) <= (layer2_outputs(3173)) and (layer2_outputs(234));
    layer3_outputs(30) <= not(layer2_outputs(1540));
    layer3_outputs(31) <= not(layer2_outputs(3694)) or (layer2_outputs(3328));
    layer3_outputs(32) <= (layer2_outputs(5421)) and not (layer2_outputs(4615));
    layer3_outputs(33) <= (layer2_outputs(5314)) and (layer2_outputs(192));
    layer3_outputs(34) <= layer2_outputs(1044);
    layer3_outputs(35) <= (layer2_outputs(3422)) and not (layer2_outputs(1393));
    layer3_outputs(36) <= layer2_outputs(5237);
    layer3_outputs(37) <= '1';
    layer3_outputs(38) <= not(layer2_outputs(5631));
    layer3_outputs(39) <= not(layer2_outputs(883));
    layer3_outputs(40) <= (layer2_outputs(4172)) and not (layer2_outputs(5218));
    layer3_outputs(41) <= (layer2_outputs(1549)) or (layer2_outputs(2318));
    layer3_outputs(42) <= not((layer2_outputs(284)) or (layer2_outputs(906)));
    layer3_outputs(43) <= not((layer2_outputs(4863)) and (layer2_outputs(940)));
    layer3_outputs(44) <= not(layer2_outputs(6762));
    layer3_outputs(45) <= not((layer2_outputs(1927)) or (layer2_outputs(2852)));
    layer3_outputs(46) <= not((layer2_outputs(6770)) and (layer2_outputs(4561)));
    layer3_outputs(47) <= layer2_outputs(2730);
    layer3_outputs(48) <= not(layer2_outputs(7616));
    layer3_outputs(49) <= not((layer2_outputs(4950)) or (layer2_outputs(6652)));
    layer3_outputs(50) <= not(layer2_outputs(1287)) or (layer2_outputs(2785));
    layer3_outputs(51) <= layer2_outputs(540);
    layer3_outputs(52) <= '0';
    layer3_outputs(53) <= not((layer2_outputs(3644)) or (layer2_outputs(949)));
    layer3_outputs(54) <= not(layer2_outputs(4218));
    layer3_outputs(55) <= (layer2_outputs(7162)) and not (layer2_outputs(6283));
    layer3_outputs(56) <= not(layer2_outputs(7365));
    layer3_outputs(57) <= layer2_outputs(182);
    layer3_outputs(58) <= not(layer2_outputs(3811)) or (layer2_outputs(5946));
    layer3_outputs(59) <= layer2_outputs(4520);
    layer3_outputs(60) <= (layer2_outputs(833)) xor (layer2_outputs(4257));
    layer3_outputs(61) <= '1';
    layer3_outputs(62) <= not(layer2_outputs(2864)) or (layer2_outputs(5678));
    layer3_outputs(63) <= layer2_outputs(6125);
    layer3_outputs(64) <= not(layer2_outputs(4628));
    layer3_outputs(65) <= (layer2_outputs(4716)) xor (layer2_outputs(3764));
    layer3_outputs(66) <= layer2_outputs(1348);
    layer3_outputs(67) <= (layer2_outputs(7071)) and not (layer2_outputs(3258));
    layer3_outputs(68) <= (layer2_outputs(996)) xor (layer2_outputs(5316));
    layer3_outputs(69) <= not(layer2_outputs(2652));
    layer3_outputs(70) <= (layer2_outputs(5362)) or (layer2_outputs(4889));
    layer3_outputs(71) <= not(layer2_outputs(2940));
    layer3_outputs(72) <= not(layer2_outputs(3830));
    layer3_outputs(73) <= '1';
    layer3_outputs(74) <= (layer2_outputs(3500)) xor (layer2_outputs(5890));
    layer3_outputs(75) <= not(layer2_outputs(2806));
    layer3_outputs(76) <= '0';
    layer3_outputs(77) <= not(layer2_outputs(3664));
    layer3_outputs(78) <= not(layer2_outputs(966));
    layer3_outputs(79) <= (layer2_outputs(5877)) and not (layer2_outputs(3257));
    layer3_outputs(80) <= (layer2_outputs(4709)) xor (layer2_outputs(1829));
    layer3_outputs(81) <= '1';
    layer3_outputs(82) <= layer2_outputs(3593);
    layer3_outputs(83) <= (layer2_outputs(3053)) and (layer2_outputs(4309));
    layer3_outputs(84) <= '1';
    layer3_outputs(85) <= not((layer2_outputs(4262)) or (layer2_outputs(913)));
    layer3_outputs(86) <= not((layer2_outputs(3431)) xor (layer2_outputs(2661)));
    layer3_outputs(87) <= not((layer2_outputs(6025)) and (layer2_outputs(963)));
    layer3_outputs(88) <= layer2_outputs(5586);
    layer3_outputs(89) <= layer2_outputs(2091);
    layer3_outputs(90) <= not(layer2_outputs(5563));
    layer3_outputs(91) <= not(layer2_outputs(5502));
    layer3_outputs(92) <= not(layer2_outputs(2302)) or (layer2_outputs(7588));
    layer3_outputs(93) <= not(layer2_outputs(1856));
    layer3_outputs(94) <= not(layer2_outputs(3184)) or (layer2_outputs(6529));
    layer3_outputs(95) <= (layer2_outputs(5478)) and (layer2_outputs(2322));
    layer3_outputs(96) <= not((layer2_outputs(5353)) or (layer2_outputs(4895)));
    layer3_outputs(97) <= not(layer2_outputs(6201)) or (layer2_outputs(1744));
    layer3_outputs(98) <= not((layer2_outputs(6688)) or (layer2_outputs(3568)));
    layer3_outputs(99) <= '0';
    layer3_outputs(100) <= (layer2_outputs(4936)) and (layer2_outputs(880));
    layer3_outputs(101) <= layer2_outputs(6061);
    layer3_outputs(102) <= layer2_outputs(1753);
    layer3_outputs(103) <= layer2_outputs(94);
    layer3_outputs(104) <= not((layer2_outputs(6233)) or (layer2_outputs(2762)));
    layer3_outputs(105) <= '1';
    layer3_outputs(106) <= (layer2_outputs(1077)) and (layer2_outputs(4395));
    layer3_outputs(107) <= layer2_outputs(4898);
    layer3_outputs(108) <= layer2_outputs(1995);
    layer3_outputs(109) <= not(layer2_outputs(2612));
    layer3_outputs(110) <= '0';
    layer3_outputs(111) <= not(layer2_outputs(7481));
    layer3_outputs(112) <= layer2_outputs(4277);
    layer3_outputs(113) <= (layer2_outputs(2866)) xor (layer2_outputs(327));
    layer3_outputs(114) <= (layer2_outputs(7361)) and not (layer2_outputs(5868));
    layer3_outputs(115) <= (layer2_outputs(925)) xor (layer2_outputs(7222));
    layer3_outputs(116) <= '1';
    layer3_outputs(117) <= (layer2_outputs(3211)) and not (layer2_outputs(3339));
    layer3_outputs(118) <= not((layer2_outputs(5178)) or (layer2_outputs(396)));
    layer3_outputs(119) <= (layer2_outputs(7402)) and not (layer2_outputs(5893));
    layer3_outputs(120) <= (layer2_outputs(2846)) or (layer2_outputs(5666));
    layer3_outputs(121) <= (layer2_outputs(6848)) and not (layer2_outputs(4263));
    layer3_outputs(122) <= not((layer2_outputs(1576)) and (layer2_outputs(2577)));
    layer3_outputs(123) <= layer2_outputs(4762);
    layer3_outputs(124) <= not((layer2_outputs(6004)) or (layer2_outputs(2664)));
    layer3_outputs(125) <= not((layer2_outputs(6056)) and (layer2_outputs(3446)));
    layer3_outputs(126) <= '0';
    layer3_outputs(127) <= '1';
    layer3_outputs(128) <= not((layer2_outputs(2602)) or (layer2_outputs(5263)));
    layer3_outputs(129) <= not((layer2_outputs(4986)) or (layer2_outputs(5134)));
    layer3_outputs(130) <= layer2_outputs(4126);
    layer3_outputs(131) <= '0';
    layer3_outputs(132) <= not((layer2_outputs(2616)) xor (layer2_outputs(5101)));
    layer3_outputs(133) <= not((layer2_outputs(1292)) and (layer2_outputs(3971)));
    layer3_outputs(134) <= (layer2_outputs(7433)) and (layer2_outputs(1131));
    layer3_outputs(135) <= not(layer2_outputs(995));
    layer3_outputs(136) <= layer2_outputs(6524);
    layer3_outputs(137) <= (layer2_outputs(5500)) and (layer2_outputs(6778));
    layer3_outputs(138) <= not(layer2_outputs(3421)) or (layer2_outputs(6763));
    layer3_outputs(139) <= '0';
    layer3_outputs(140) <= layer2_outputs(5501);
    layer3_outputs(141) <= not(layer2_outputs(2496)) or (layer2_outputs(2786));
    layer3_outputs(142) <= (layer2_outputs(244)) or (layer2_outputs(4685));
    layer3_outputs(143) <= (layer2_outputs(3711)) and (layer2_outputs(5955));
    layer3_outputs(144) <= not((layer2_outputs(4514)) or (layer2_outputs(4666)));
    layer3_outputs(145) <= layer2_outputs(3114);
    layer3_outputs(146) <= not((layer2_outputs(2606)) and (layer2_outputs(783)));
    layer3_outputs(147) <= '0';
    layer3_outputs(148) <= not(layer2_outputs(3499));
    layer3_outputs(149) <= layer2_outputs(7498);
    layer3_outputs(150) <= '1';
    layer3_outputs(151) <= layer2_outputs(5676);
    layer3_outputs(152) <= not((layer2_outputs(5783)) or (layer2_outputs(2006)));
    layer3_outputs(153) <= layer2_outputs(3667);
    layer3_outputs(154) <= '1';
    layer3_outputs(155) <= not(layer2_outputs(7281));
    layer3_outputs(156) <= (layer2_outputs(4753)) and not (layer2_outputs(7310));
    layer3_outputs(157) <= not(layer2_outputs(2467));
    layer3_outputs(158) <= not((layer2_outputs(4180)) and (layer2_outputs(2357)));
    layer3_outputs(159) <= not((layer2_outputs(933)) and (layer2_outputs(4575)));
    layer3_outputs(160) <= not(layer2_outputs(5148));
    layer3_outputs(161) <= (layer2_outputs(6669)) or (layer2_outputs(4228));
    layer3_outputs(162) <= layer2_outputs(6604);
    layer3_outputs(163) <= layer2_outputs(5596);
    layer3_outputs(164) <= not(layer2_outputs(1985)) or (layer2_outputs(396));
    layer3_outputs(165) <= not((layer2_outputs(5127)) or (layer2_outputs(6324)));
    layer3_outputs(166) <= not(layer2_outputs(3546));
    layer3_outputs(167) <= '0';
    layer3_outputs(168) <= not(layer2_outputs(7641));
    layer3_outputs(169) <= not((layer2_outputs(4778)) and (layer2_outputs(3189)));
    layer3_outputs(170) <= not(layer2_outputs(1012)) or (layer2_outputs(6038));
    layer3_outputs(171) <= (layer2_outputs(4139)) and not (layer2_outputs(3187));
    layer3_outputs(172) <= not(layer2_outputs(7048));
    layer3_outputs(173) <= not(layer2_outputs(3877));
    layer3_outputs(174) <= (layer2_outputs(1515)) or (layer2_outputs(458));
    layer3_outputs(175) <= (layer2_outputs(7026)) and not (layer2_outputs(4561));
    layer3_outputs(176) <= '0';
    layer3_outputs(177) <= not(layer2_outputs(3870));
    layer3_outputs(178) <= '0';
    layer3_outputs(179) <= layer2_outputs(1296);
    layer3_outputs(180) <= layer2_outputs(5017);
    layer3_outputs(181) <= layer2_outputs(5490);
    layer3_outputs(182) <= not((layer2_outputs(4725)) and (layer2_outputs(4337)));
    layer3_outputs(183) <= layer2_outputs(6664);
    layer3_outputs(184) <= (layer2_outputs(7169)) and not (layer2_outputs(1892));
    layer3_outputs(185) <= not(layer2_outputs(4343));
    layer3_outputs(186) <= not(layer2_outputs(179));
    layer3_outputs(187) <= not(layer2_outputs(880));
    layer3_outputs(188) <= (layer2_outputs(2843)) and not (layer2_outputs(124));
    layer3_outputs(189) <= layer2_outputs(3776);
    layer3_outputs(190) <= (layer2_outputs(1369)) or (layer2_outputs(7186));
    layer3_outputs(191) <= '0';
    layer3_outputs(192) <= (layer2_outputs(6865)) or (layer2_outputs(7459));
    layer3_outputs(193) <= layer2_outputs(1893);
    layer3_outputs(194) <= not(layer2_outputs(1164));
    layer3_outputs(195) <= (layer2_outputs(4258)) and not (layer2_outputs(581));
    layer3_outputs(196) <= layer2_outputs(2891);
    layer3_outputs(197) <= (layer2_outputs(4940)) and not (layer2_outputs(2043));
    layer3_outputs(198) <= layer2_outputs(2568);
    layer3_outputs(199) <= layer2_outputs(1558);
    layer3_outputs(200) <= not((layer2_outputs(1278)) and (layer2_outputs(2327)));
    layer3_outputs(201) <= '0';
    layer3_outputs(202) <= not(layer2_outputs(1627)) or (layer2_outputs(7496));
    layer3_outputs(203) <= not((layer2_outputs(2476)) or (layer2_outputs(307)));
    layer3_outputs(204) <= not((layer2_outputs(3637)) and (layer2_outputs(3689)));
    layer3_outputs(205) <= not(layer2_outputs(5943));
    layer3_outputs(206) <= (layer2_outputs(462)) and (layer2_outputs(5573));
    layer3_outputs(207) <= not(layer2_outputs(501));
    layer3_outputs(208) <= not(layer2_outputs(967)) or (layer2_outputs(7523));
    layer3_outputs(209) <= not(layer2_outputs(4525)) or (layer2_outputs(5905));
    layer3_outputs(210) <= (layer2_outputs(1708)) and not (layer2_outputs(813));
    layer3_outputs(211) <= not(layer2_outputs(3155));
    layer3_outputs(212) <= '1';
    layer3_outputs(213) <= layer2_outputs(7027);
    layer3_outputs(214) <= not(layer2_outputs(5241));
    layer3_outputs(215) <= (layer2_outputs(7258)) and not (layer2_outputs(3364));
    layer3_outputs(216) <= not(layer2_outputs(5231)) or (layer2_outputs(3828));
    layer3_outputs(217) <= '1';
    layer3_outputs(218) <= (layer2_outputs(1827)) and (layer2_outputs(4825));
    layer3_outputs(219) <= not(layer2_outputs(4192)) or (layer2_outputs(1235));
    layer3_outputs(220) <= not(layer2_outputs(1501));
    layer3_outputs(221) <= (layer2_outputs(5724)) and not (layer2_outputs(6589));
    layer3_outputs(222) <= (layer2_outputs(5565)) or (layer2_outputs(4926));
    layer3_outputs(223) <= layer2_outputs(1208);
    layer3_outputs(224) <= not((layer2_outputs(4958)) or (layer2_outputs(2579)));
    layer3_outputs(225) <= layer2_outputs(4510);
    layer3_outputs(226) <= (layer2_outputs(2105)) and not (layer2_outputs(7394));
    layer3_outputs(227) <= not(layer2_outputs(686));
    layer3_outputs(228) <= layer2_outputs(5634);
    layer3_outputs(229) <= (layer2_outputs(5793)) or (layer2_outputs(4454));
    layer3_outputs(230) <= not((layer2_outputs(4494)) and (layer2_outputs(440)));
    layer3_outputs(231) <= '0';
    layer3_outputs(232) <= layer2_outputs(7043);
    layer3_outputs(233) <= layer2_outputs(392);
    layer3_outputs(234) <= not((layer2_outputs(4515)) xor (layer2_outputs(2970)));
    layer3_outputs(235) <= not(layer2_outputs(5630));
    layer3_outputs(236) <= not(layer2_outputs(4152));
    layer3_outputs(237) <= layer2_outputs(915);
    layer3_outputs(238) <= '1';
    layer3_outputs(239) <= (layer2_outputs(6644)) and not (layer2_outputs(6698));
    layer3_outputs(240) <= (layer2_outputs(90)) and not (layer2_outputs(4041));
    layer3_outputs(241) <= not(layer2_outputs(1620));
    layer3_outputs(242) <= layer2_outputs(6900);
    layer3_outputs(243) <= layer2_outputs(5914);
    layer3_outputs(244) <= (layer2_outputs(122)) or (layer2_outputs(4248));
    layer3_outputs(245) <= layer2_outputs(7286);
    layer3_outputs(246) <= layer2_outputs(4780);
    layer3_outputs(247) <= (layer2_outputs(3252)) xor (layer2_outputs(5370));
    layer3_outputs(248) <= '0';
    layer3_outputs(249) <= not(layer2_outputs(2777));
    layer3_outputs(250) <= layer2_outputs(4113);
    layer3_outputs(251) <= (layer2_outputs(4074)) and not (layer2_outputs(2566));
    layer3_outputs(252) <= layer2_outputs(4734);
    layer3_outputs(253) <= not(layer2_outputs(6881));
    layer3_outputs(254) <= layer2_outputs(4259);
    layer3_outputs(255) <= not(layer2_outputs(2648));
    layer3_outputs(256) <= (layer2_outputs(1850)) or (layer2_outputs(3190));
    layer3_outputs(257) <= not(layer2_outputs(4627)) or (layer2_outputs(6072));
    layer3_outputs(258) <= not(layer2_outputs(359));
    layer3_outputs(259) <= (layer2_outputs(6348)) or (layer2_outputs(5204));
    layer3_outputs(260) <= (layer2_outputs(749)) and not (layer2_outputs(1697));
    layer3_outputs(261) <= not((layer2_outputs(3989)) and (layer2_outputs(2826)));
    layer3_outputs(262) <= '0';
    layer3_outputs(263) <= '1';
    layer3_outputs(264) <= layer2_outputs(2684);
    layer3_outputs(265) <= layer2_outputs(4601);
    layer3_outputs(266) <= layer2_outputs(380);
    layer3_outputs(267) <= layer2_outputs(169);
    layer3_outputs(268) <= not((layer2_outputs(1742)) xor (layer2_outputs(2426)));
    layer3_outputs(269) <= not(layer2_outputs(6381));
    layer3_outputs(270) <= (layer2_outputs(4215)) or (layer2_outputs(2392));
    layer3_outputs(271) <= not(layer2_outputs(1354)) or (layer2_outputs(1082));
    layer3_outputs(272) <= not((layer2_outputs(2503)) and (layer2_outputs(5937)));
    layer3_outputs(273) <= (layer2_outputs(5583)) or (layer2_outputs(6762));
    layer3_outputs(274) <= (layer2_outputs(1548)) or (layer2_outputs(2935));
    layer3_outputs(275) <= not(layer2_outputs(7627));
    layer3_outputs(276) <= layer2_outputs(702);
    layer3_outputs(277) <= not(layer2_outputs(7259));
    layer3_outputs(278) <= layer2_outputs(1987);
    layer3_outputs(279) <= '0';
    layer3_outputs(280) <= not(layer2_outputs(5288)) or (layer2_outputs(3326));
    layer3_outputs(281) <= (layer2_outputs(7172)) and (layer2_outputs(297));
    layer3_outputs(282) <= (layer2_outputs(6903)) and not (layer2_outputs(6571));
    layer3_outputs(283) <= (layer2_outputs(3570)) or (layer2_outputs(2037));
    layer3_outputs(284) <= not((layer2_outputs(7181)) or (layer2_outputs(1057)));
    layer3_outputs(285) <= layer2_outputs(2414);
    layer3_outputs(286) <= not(layer2_outputs(3756));
    layer3_outputs(287) <= not(layer2_outputs(1333));
    layer3_outputs(288) <= layer2_outputs(5585);
    layer3_outputs(289) <= (layer2_outputs(954)) and not (layer2_outputs(2793));
    layer3_outputs(290) <= (layer2_outputs(775)) or (layer2_outputs(5566));
    layer3_outputs(291) <= not((layer2_outputs(2667)) or (layer2_outputs(1931)));
    layer3_outputs(292) <= layer2_outputs(5363);
    layer3_outputs(293) <= not((layer2_outputs(4629)) or (layer2_outputs(5781)));
    layer3_outputs(294) <= not(layer2_outputs(3141)) or (layer2_outputs(6870));
    layer3_outputs(295) <= not(layer2_outputs(5034));
    layer3_outputs(296) <= (layer2_outputs(2161)) and not (layer2_outputs(6471));
    layer3_outputs(297) <= not(layer2_outputs(7154)) or (layer2_outputs(1216));
    layer3_outputs(298) <= layer2_outputs(2714);
    layer3_outputs(299) <= '1';
    layer3_outputs(300) <= layer2_outputs(4944);
    layer3_outputs(301) <= (layer2_outputs(4020)) and (layer2_outputs(5839));
    layer3_outputs(302) <= not((layer2_outputs(5124)) or (layer2_outputs(7020)));
    layer3_outputs(303) <= (layer2_outputs(206)) or (layer2_outputs(5589));
    layer3_outputs(304) <= (layer2_outputs(3460)) and not (layer2_outputs(384));
    layer3_outputs(305) <= not((layer2_outputs(6750)) or (layer2_outputs(4476)));
    layer3_outputs(306) <= (layer2_outputs(4479)) or (layer2_outputs(6641));
    layer3_outputs(307) <= layer2_outputs(2967);
    layer3_outputs(308) <= (layer2_outputs(2665)) and (layer2_outputs(5485));
    layer3_outputs(309) <= not(layer2_outputs(5100));
    layer3_outputs(310) <= layer2_outputs(5136);
    layer3_outputs(311) <= layer2_outputs(5800);
    layer3_outputs(312) <= layer2_outputs(4103);
    layer3_outputs(313) <= not(layer2_outputs(5970)) or (layer2_outputs(956));
    layer3_outputs(314) <= (layer2_outputs(2794)) or (layer2_outputs(3108));
    layer3_outputs(315) <= layer2_outputs(4727);
    layer3_outputs(316) <= '1';
    layer3_outputs(317) <= layer2_outputs(2340);
    layer3_outputs(318) <= not(layer2_outputs(3485)) or (layer2_outputs(471));
    layer3_outputs(319) <= '0';
    layer3_outputs(320) <= (layer2_outputs(1785)) and not (layer2_outputs(1884));
    layer3_outputs(321) <= (layer2_outputs(3819)) and not (layer2_outputs(3556));
    layer3_outputs(322) <= (layer2_outputs(4216)) or (layer2_outputs(5157));
    layer3_outputs(323) <= (layer2_outputs(2252)) or (layer2_outputs(2244));
    layer3_outputs(324) <= not((layer2_outputs(311)) or (layer2_outputs(3419)));
    layer3_outputs(325) <= layer2_outputs(7359);
    layer3_outputs(326) <= not(layer2_outputs(5305)) or (layer2_outputs(5186));
    layer3_outputs(327) <= layer2_outputs(1962);
    layer3_outputs(328) <= not(layer2_outputs(6924));
    layer3_outputs(329) <= (layer2_outputs(3231)) and not (layer2_outputs(3892));
    layer3_outputs(330) <= not((layer2_outputs(2767)) and (layer2_outputs(1958)));
    layer3_outputs(331) <= not((layer2_outputs(3686)) and (layer2_outputs(6735)));
    layer3_outputs(332) <= not(layer2_outputs(7368));
    layer3_outputs(333) <= (layer2_outputs(1976)) and not (layer2_outputs(2226));
    layer3_outputs(334) <= '0';
    layer3_outputs(335) <= (layer2_outputs(6116)) and not (layer2_outputs(2632));
    layer3_outputs(336) <= not(layer2_outputs(4839));
    layer3_outputs(337) <= (layer2_outputs(5252)) and (layer2_outputs(3171));
    layer3_outputs(338) <= (layer2_outputs(2574)) or (layer2_outputs(6726));
    layer3_outputs(339) <= layer2_outputs(2579);
    layer3_outputs(340) <= '0';
    layer3_outputs(341) <= layer2_outputs(6171);
    layer3_outputs(342) <= not(layer2_outputs(2804)) or (layer2_outputs(4423));
    layer3_outputs(343) <= (layer2_outputs(1832)) and not (layer2_outputs(5490));
    layer3_outputs(344) <= (layer2_outputs(7333)) and (layer2_outputs(3234));
    layer3_outputs(345) <= not((layer2_outputs(4491)) and (layer2_outputs(2041)));
    layer3_outputs(346) <= not(layer2_outputs(68));
    layer3_outputs(347) <= layer2_outputs(2052);
    layer3_outputs(348) <= layer2_outputs(319);
    layer3_outputs(349) <= not(layer2_outputs(6551));
    layer3_outputs(350) <= (layer2_outputs(6031)) and (layer2_outputs(2921));
    layer3_outputs(351) <= not((layer2_outputs(1480)) or (layer2_outputs(6959)));
    layer3_outputs(352) <= layer2_outputs(770);
    layer3_outputs(353) <= (layer2_outputs(1428)) xor (layer2_outputs(5083));
    layer3_outputs(354) <= not(layer2_outputs(6509));
    layer3_outputs(355) <= not(layer2_outputs(2819));
    layer3_outputs(356) <= (layer2_outputs(6869)) or (layer2_outputs(7341));
    layer3_outputs(357) <= (layer2_outputs(3137)) xor (layer2_outputs(6049));
    layer3_outputs(358) <= (layer2_outputs(7528)) xor (layer2_outputs(3006));
    layer3_outputs(359) <= not((layer2_outputs(5602)) and (layer2_outputs(6435)));
    layer3_outputs(360) <= not(layer2_outputs(1166));
    layer3_outputs(361) <= not(layer2_outputs(6303));
    layer3_outputs(362) <= (layer2_outputs(6112)) and (layer2_outputs(3112));
    layer3_outputs(363) <= layer2_outputs(4932);
    layer3_outputs(364) <= layer2_outputs(2139);
    layer3_outputs(365) <= not((layer2_outputs(4075)) and (layer2_outputs(1578)));
    layer3_outputs(366) <= layer2_outputs(1283);
    layer3_outputs(367) <= layer2_outputs(3067);
    layer3_outputs(368) <= '0';
    layer3_outputs(369) <= not(layer2_outputs(716));
    layer3_outputs(370) <= not((layer2_outputs(5077)) or (layer2_outputs(1513)));
    layer3_outputs(371) <= not(layer2_outputs(3163));
    layer3_outputs(372) <= layer2_outputs(4265);
    layer3_outputs(373) <= (layer2_outputs(6769)) and (layer2_outputs(5827));
    layer3_outputs(374) <= not(layer2_outputs(1399));
    layer3_outputs(375) <= not((layer2_outputs(5140)) and (layer2_outputs(4028)));
    layer3_outputs(376) <= not(layer2_outputs(2263)) or (layer2_outputs(3200));
    layer3_outputs(377) <= '1';
    layer3_outputs(378) <= '0';
    layer3_outputs(379) <= (layer2_outputs(1123)) xor (layer2_outputs(3513));
    layer3_outputs(380) <= '0';
    layer3_outputs(381) <= '0';
    layer3_outputs(382) <= layer2_outputs(7544);
    layer3_outputs(383) <= (layer2_outputs(1540)) and not (layer2_outputs(5275));
    layer3_outputs(384) <= layer2_outputs(4935);
    layer3_outputs(385) <= not(layer2_outputs(3651));
    layer3_outputs(386) <= not((layer2_outputs(7589)) and (layer2_outputs(71)));
    layer3_outputs(387) <= (layer2_outputs(5277)) and not (layer2_outputs(3226));
    layer3_outputs(388) <= layer2_outputs(6148);
    layer3_outputs(389) <= not((layer2_outputs(344)) or (layer2_outputs(5217)));
    layer3_outputs(390) <= not(layer2_outputs(3382));
    layer3_outputs(391) <= layer2_outputs(5339);
    layer3_outputs(392) <= not((layer2_outputs(5562)) or (layer2_outputs(7668)));
    layer3_outputs(393) <= not(layer2_outputs(6575));
    layer3_outputs(394) <= not(layer2_outputs(1668));
    layer3_outputs(395) <= '1';
    layer3_outputs(396) <= (layer2_outputs(6165)) and (layer2_outputs(1052));
    layer3_outputs(397) <= layer2_outputs(7672);
    layer3_outputs(398) <= not(layer2_outputs(1546));
    layer3_outputs(399) <= (layer2_outputs(5041)) and not (layer2_outputs(4697));
    layer3_outputs(400) <= not(layer2_outputs(5909));
    layer3_outputs(401) <= not((layer2_outputs(3502)) or (layer2_outputs(2435)));
    layer3_outputs(402) <= '0';
    layer3_outputs(403) <= not((layer2_outputs(3222)) or (layer2_outputs(5925)));
    layer3_outputs(404) <= not(layer2_outputs(4852));
    layer3_outputs(405) <= not(layer2_outputs(6786));
    layer3_outputs(406) <= not(layer2_outputs(690));
    layer3_outputs(407) <= not(layer2_outputs(5418));
    layer3_outputs(408) <= '1';
    layer3_outputs(409) <= (layer2_outputs(7207)) and not (layer2_outputs(5552));
    layer3_outputs(410) <= not(layer2_outputs(2697)) or (layer2_outputs(6564));
    layer3_outputs(411) <= '1';
    layer3_outputs(412) <= layer2_outputs(7679);
    layer3_outputs(413) <= not(layer2_outputs(5489)) or (layer2_outputs(1790));
    layer3_outputs(414) <= (layer2_outputs(5083)) and not (layer2_outputs(4513));
    layer3_outputs(415) <= layer2_outputs(3360);
    layer3_outputs(416) <= '1';
    layer3_outputs(417) <= (layer2_outputs(2761)) and not (layer2_outputs(4710));
    layer3_outputs(418) <= not((layer2_outputs(5555)) and (layer2_outputs(3089)));
    layer3_outputs(419) <= (layer2_outputs(2268)) xor (layer2_outputs(7296));
    layer3_outputs(420) <= (layer2_outputs(3687)) and not (layer2_outputs(7261));
    layer3_outputs(421) <= not(layer2_outputs(6290));
    layer3_outputs(422) <= (layer2_outputs(4344)) and (layer2_outputs(3860));
    layer3_outputs(423) <= not(layer2_outputs(2638)) or (layer2_outputs(1201));
    layer3_outputs(424) <= (layer2_outputs(1861)) and not (layer2_outputs(6577));
    layer3_outputs(425) <= not(layer2_outputs(5468)) or (layer2_outputs(2100));
    layer3_outputs(426) <= layer2_outputs(918);
    layer3_outputs(427) <= not((layer2_outputs(5265)) and (layer2_outputs(6662)));
    layer3_outputs(428) <= not(layer2_outputs(2163));
    layer3_outputs(429) <= (layer2_outputs(5172)) or (layer2_outputs(2612));
    layer3_outputs(430) <= layer2_outputs(5417);
    layer3_outputs(431) <= (layer2_outputs(3215)) and not (layer2_outputs(3042));
    layer3_outputs(432) <= (layer2_outputs(3196)) xor (layer2_outputs(2835));
    layer3_outputs(433) <= '1';
    layer3_outputs(434) <= (layer2_outputs(1982)) or (layer2_outputs(6515));
    layer3_outputs(435) <= not((layer2_outputs(7663)) and (layer2_outputs(1981)));
    layer3_outputs(436) <= '0';
    layer3_outputs(437) <= not(layer2_outputs(6680));
    layer3_outputs(438) <= not(layer2_outputs(7411));
    layer3_outputs(439) <= not((layer2_outputs(6346)) or (layer2_outputs(4183)));
    layer3_outputs(440) <= (layer2_outputs(4646)) or (layer2_outputs(6621));
    layer3_outputs(441) <= not((layer2_outputs(332)) and (layer2_outputs(1671)));
    layer3_outputs(442) <= not(layer2_outputs(119));
    layer3_outputs(443) <= not(layer2_outputs(1552));
    layer3_outputs(444) <= not(layer2_outputs(2134)) or (layer2_outputs(7333));
    layer3_outputs(445) <= (layer2_outputs(4567)) and not (layer2_outputs(473));
    layer3_outputs(446) <= not(layer2_outputs(4533)) or (layer2_outputs(2967));
    layer3_outputs(447) <= not(layer2_outputs(2671)) or (layer2_outputs(4826));
    layer3_outputs(448) <= layer2_outputs(1226);
    layer3_outputs(449) <= layer2_outputs(1076);
    layer3_outputs(450) <= not(layer2_outputs(4037)) or (layer2_outputs(6704));
    layer3_outputs(451) <= layer2_outputs(651);
    layer3_outputs(452) <= not(layer2_outputs(52)) or (layer2_outputs(1277));
    layer3_outputs(453) <= not((layer2_outputs(1017)) or (layer2_outputs(1719)));
    layer3_outputs(454) <= (layer2_outputs(4109)) and not (layer2_outputs(2625));
    layer3_outputs(455) <= not(layer2_outputs(6330));
    layer3_outputs(456) <= not(layer2_outputs(4345));
    layer3_outputs(457) <= not(layer2_outputs(7247)) or (layer2_outputs(2950));
    layer3_outputs(458) <= not(layer2_outputs(5486));
    layer3_outputs(459) <= not(layer2_outputs(3660));
    layer3_outputs(460) <= not(layer2_outputs(4375)) or (layer2_outputs(7637));
    layer3_outputs(461) <= not((layer2_outputs(5002)) or (layer2_outputs(1602)));
    layer3_outputs(462) <= '1';
    layer3_outputs(463) <= not((layer2_outputs(6208)) or (layer2_outputs(4793)));
    layer3_outputs(464) <= not(layer2_outputs(6303)) or (layer2_outputs(634));
    layer3_outputs(465) <= (layer2_outputs(1246)) and not (layer2_outputs(7486));
    layer3_outputs(466) <= not((layer2_outputs(4318)) or (layer2_outputs(467)));
    layer3_outputs(467) <= not((layer2_outputs(348)) or (layer2_outputs(2345)));
    layer3_outputs(468) <= not(layer2_outputs(5327));
    layer3_outputs(469) <= layer2_outputs(4390);
    layer3_outputs(470) <= not(layer2_outputs(5188));
    layer3_outputs(471) <= (layer2_outputs(5197)) and not (layer2_outputs(542));
    layer3_outputs(472) <= '1';
    layer3_outputs(473) <= (layer2_outputs(1023)) and not (layer2_outputs(3103));
    layer3_outputs(474) <= layer2_outputs(1163);
    layer3_outputs(475) <= (layer2_outputs(5112)) or (layer2_outputs(5018));
    layer3_outputs(476) <= layer2_outputs(4455);
    layer3_outputs(477) <= not(layer2_outputs(2680)) or (layer2_outputs(415));
    layer3_outputs(478) <= not((layer2_outputs(6049)) or (layer2_outputs(2874)));
    layer3_outputs(479) <= '1';
    layer3_outputs(480) <= not((layer2_outputs(6893)) or (layer2_outputs(5428)));
    layer3_outputs(481) <= '0';
    layer3_outputs(482) <= not(layer2_outputs(7561));
    layer3_outputs(483) <= layer2_outputs(6259);
    layer3_outputs(484) <= not(layer2_outputs(6886)) or (layer2_outputs(6317));
    layer3_outputs(485) <= layer2_outputs(3555);
    layer3_outputs(486) <= not(layer2_outputs(3400));
    layer3_outputs(487) <= not(layer2_outputs(2745)) or (layer2_outputs(950));
    layer3_outputs(488) <= not(layer2_outputs(2770));
    layer3_outputs(489) <= layer2_outputs(1134);
    layer3_outputs(490) <= '0';
    layer3_outputs(491) <= not(layer2_outputs(1490)) or (layer2_outputs(2276));
    layer3_outputs(492) <= not(layer2_outputs(1470)) or (layer2_outputs(3845));
    layer3_outputs(493) <= (layer2_outputs(1276)) or (layer2_outputs(1849));
    layer3_outputs(494) <= layer2_outputs(6410);
    layer3_outputs(495) <= not((layer2_outputs(6080)) or (layer2_outputs(4433)));
    layer3_outputs(496) <= not(layer2_outputs(3781)) or (layer2_outputs(4565));
    layer3_outputs(497) <= not(layer2_outputs(34)) or (layer2_outputs(1869));
    layer3_outputs(498) <= not(layer2_outputs(941));
    layer3_outputs(499) <= layer2_outputs(51);
    layer3_outputs(500) <= not(layer2_outputs(6580));
    layer3_outputs(501) <= not(layer2_outputs(4261)) or (layer2_outputs(7232));
    layer3_outputs(502) <= not((layer2_outputs(1682)) and (layer2_outputs(4543)));
    layer3_outputs(503) <= layer2_outputs(5960);
    layer3_outputs(504) <= layer2_outputs(539);
    layer3_outputs(505) <= not(layer2_outputs(3138)) or (layer2_outputs(7235));
    layer3_outputs(506) <= not(layer2_outputs(1713));
    layer3_outputs(507) <= not(layer2_outputs(5727)) or (layer2_outputs(7080));
    layer3_outputs(508) <= layer2_outputs(5990);
    layer3_outputs(509) <= not((layer2_outputs(1431)) or (layer2_outputs(3498)));
    layer3_outputs(510) <= not(layer2_outputs(1380));
    layer3_outputs(511) <= '0';
    layer3_outputs(512) <= (layer2_outputs(4925)) and not (layer2_outputs(4198));
    layer3_outputs(513) <= not(layer2_outputs(4628));
    layer3_outputs(514) <= (layer2_outputs(349)) xor (layer2_outputs(1654));
    layer3_outputs(515) <= not(layer2_outputs(4836)) or (layer2_outputs(7289));
    layer3_outputs(516) <= not(layer2_outputs(5951));
    layer3_outputs(517) <= (layer2_outputs(3622)) and not (layer2_outputs(1419));
    layer3_outputs(518) <= not((layer2_outputs(7062)) and (layer2_outputs(2112)));
    layer3_outputs(519) <= not(layer2_outputs(1647)) or (layer2_outputs(7465));
    layer3_outputs(520) <= layer2_outputs(6395);
    layer3_outputs(521) <= '1';
    layer3_outputs(522) <= (layer2_outputs(1923)) and (layer2_outputs(7204));
    layer3_outputs(523) <= '1';
    layer3_outputs(524) <= (layer2_outputs(3120)) and (layer2_outputs(3635));
    layer3_outputs(525) <= '0';
    layer3_outputs(526) <= not(layer2_outputs(1686));
    layer3_outputs(527) <= not(layer2_outputs(7678));
    layer3_outputs(528) <= (layer2_outputs(4896)) and (layer2_outputs(6144));
    layer3_outputs(529) <= (layer2_outputs(1437)) and not (layer2_outputs(4464));
    layer3_outputs(530) <= (layer2_outputs(6508)) and (layer2_outputs(3745));
    layer3_outputs(531) <= not((layer2_outputs(4667)) and (layer2_outputs(617)));
    layer3_outputs(532) <= not(layer2_outputs(3700));
    layer3_outputs(533) <= not(layer2_outputs(5400));
    layer3_outputs(534) <= (layer2_outputs(2392)) and not (layer2_outputs(6898));
    layer3_outputs(535) <= not(layer2_outputs(70));
    layer3_outputs(536) <= not(layer2_outputs(4993)) or (layer2_outputs(4833));
    layer3_outputs(537) <= (layer2_outputs(777)) and not (layer2_outputs(2514));
    layer3_outputs(538) <= not(layer2_outputs(7350));
    layer3_outputs(539) <= not(layer2_outputs(6919));
    layer3_outputs(540) <= layer2_outputs(6064);
    layer3_outputs(541) <= (layer2_outputs(4399)) and not (layer2_outputs(3004));
    layer3_outputs(542) <= (layer2_outputs(399)) or (layer2_outputs(3895));
    layer3_outputs(543) <= not((layer2_outputs(5224)) or (layer2_outputs(4387)));
    layer3_outputs(544) <= (layer2_outputs(5729)) xor (layer2_outputs(7513));
    layer3_outputs(545) <= not(layer2_outputs(6396));
    layer3_outputs(546) <= not(layer2_outputs(3230)) or (layer2_outputs(4731));
    layer3_outputs(547) <= not(layer2_outputs(4406));
    layer3_outputs(548) <= (layer2_outputs(4243)) or (layer2_outputs(1627));
    layer3_outputs(549) <= (layer2_outputs(6177)) and not (layer2_outputs(3688));
    layer3_outputs(550) <= (layer2_outputs(1366)) xor (layer2_outputs(1261));
    layer3_outputs(551) <= '1';
    layer3_outputs(552) <= not((layer2_outputs(3324)) and (layer2_outputs(333)));
    layer3_outputs(553) <= layer2_outputs(2069);
    layer3_outputs(554) <= not(layer2_outputs(5058));
    layer3_outputs(555) <= (layer2_outputs(1779)) and (layer2_outputs(3567));
    layer3_outputs(556) <= '0';
    layer3_outputs(557) <= not(layer2_outputs(924)) or (layer2_outputs(6822));
    layer3_outputs(558) <= not(layer2_outputs(6147)) or (layer2_outputs(3081));
    layer3_outputs(559) <= (layer2_outputs(5691)) or (layer2_outputs(1071));
    layer3_outputs(560) <= layer2_outputs(2199);
    layer3_outputs(561) <= (layer2_outputs(614)) or (layer2_outputs(3866));
    layer3_outputs(562) <= layer2_outputs(5717);
    layer3_outputs(563) <= (layer2_outputs(6298)) and (layer2_outputs(4063));
    layer3_outputs(564) <= '1';
    layer3_outputs(565) <= '0';
    layer3_outputs(566) <= not((layer2_outputs(2495)) and (layer2_outputs(2352)));
    layer3_outputs(567) <= layer2_outputs(1214);
    layer3_outputs(568) <= not(layer2_outputs(7577)) or (layer2_outputs(7235));
    layer3_outputs(569) <= (layer2_outputs(5741)) and (layer2_outputs(4710));
    layer3_outputs(570) <= layer2_outputs(5851);
    layer3_outputs(571) <= not((layer2_outputs(7394)) or (layer2_outputs(7225)));
    layer3_outputs(572) <= not(layer2_outputs(4310)) or (layer2_outputs(6773));
    layer3_outputs(573) <= layer2_outputs(4516);
    layer3_outputs(574) <= '0';
    layer3_outputs(575) <= not((layer2_outputs(3274)) or (layer2_outputs(5119)));
    layer3_outputs(576) <= (layer2_outputs(2317)) and not (layer2_outputs(5958));
    layer3_outputs(577) <= (layer2_outputs(5314)) and not (layer2_outputs(906));
    layer3_outputs(578) <= not(layer2_outputs(6724));
    layer3_outputs(579) <= (layer2_outputs(6876)) and not (layer2_outputs(1613));
    layer3_outputs(580) <= not(layer2_outputs(3097));
    layer3_outputs(581) <= not(layer2_outputs(6535));
    layer3_outputs(582) <= layer2_outputs(5393);
    layer3_outputs(583) <= not(layer2_outputs(5750));
    layer3_outputs(584) <= not(layer2_outputs(1807));
    layer3_outputs(585) <= not((layer2_outputs(1834)) and (layer2_outputs(7365)));
    layer3_outputs(586) <= '1';
    layer3_outputs(587) <= not(layer2_outputs(330)) or (layer2_outputs(1609));
    layer3_outputs(588) <= not(layer2_outputs(5299));
    layer3_outputs(589) <= layer2_outputs(1903);
    layer3_outputs(590) <= not(layer2_outputs(1651)) or (layer2_outputs(5976));
    layer3_outputs(591) <= layer2_outputs(4034);
    layer3_outputs(592) <= (layer2_outputs(643)) and not (layer2_outputs(3926));
    layer3_outputs(593) <= not(layer2_outputs(1367));
    layer3_outputs(594) <= layer2_outputs(6893);
    layer3_outputs(595) <= not(layer2_outputs(2037));
    layer3_outputs(596) <= not(layer2_outputs(5186));
    layer3_outputs(597) <= layer2_outputs(3014);
    layer3_outputs(598) <= (layer2_outputs(2145)) and not (layer2_outputs(5203));
    layer3_outputs(599) <= not((layer2_outputs(5380)) xor (layer2_outputs(6180)));
    layer3_outputs(600) <= (layer2_outputs(229)) and not (layer2_outputs(6469));
    layer3_outputs(601) <= not((layer2_outputs(7455)) or (layer2_outputs(4322)));
    layer3_outputs(602) <= not((layer2_outputs(3858)) or (layer2_outputs(5945)));
    layer3_outputs(603) <= layer2_outputs(4161);
    layer3_outputs(604) <= (layer2_outputs(3476)) or (layer2_outputs(6780));
    layer3_outputs(605) <= '0';
    layer3_outputs(606) <= (layer2_outputs(5882)) or (layer2_outputs(1158));
    layer3_outputs(607) <= '1';
    layer3_outputs(608) <= not(layer2_outputs(5467));
    layer3_outputs(609) <= layer2_outputs(2088);
    layer3_outputs(610) <= (layer2_outputs(209)) and (layer2_outputs(2805));
    layer3_outputs(611) <= not(layer2_outputs(2010));
    layer3_outputs(612) <= layer2_outputs(900);
    layer3_outputs(613) <= '0';
    layer3_outputs(614) <= not(layer2_outputs(6541)) or (layer2_outputs(7281));
    layer3_outputs(615) <= (layer2_outputs(1816)) and not (layer2_outputs(5998));
    layer3_outputs(616) <= (layer2_outputs(6719)) and (layer2_outputs(4523));
    layer3_outputs(617) <= not(layer2_outputs(715));
    layer3_outputs(618) <= layer2_outputs(1974);
    layer3_outputs(619) <= '1';
    layer3_outputs(620) <= layer2_outputs(105);
    layer3_outputs(621) <= (layer2_outputs(5614)) or (layer2_outputs(4435));
    layer3_outputs(622) <= not(layer2_outputs(6461));
    layer3_outputs(623) <= (layer2_outputs(5384)) and (layer2_outputs(2447));
    layer3_outputs(624) <= layer2_outputs(4380);
    layer3_outputs(625) <= layer2_outputs(3861);
    layer3_outputs(626) <= (layer2_outputs(2707)) and not (layer2_outputs(6670));
    layer3_outputs(627) <= not(layer2_outputs(4309)) or (layer2_outputs(2219));
    layer3_outputs(628) <= layer2_outputs(6597);
    layer3_outputs(629) <= layer2_outputs(2722);
    layer3_outputs(630) <= '1';
    layer3_outputs(631) <= layer2_outputs(5981);
    layer3_outputs(632) <= (layer2_outputs(6925)) or (layer2_outputs(5113));
    layer3_outputs(633) <= '0';
    layer3_outputs(634) <= (layer2_outputs(3695)) and not (layer2_outputs(1645));
    layer3_outputs(635) <= layer2_outputs(3871);
    layer3_outputs(636) <= not(layer2_outputs(2972)) or (layer2_outputs(3851));
    layer3_outputs(637) <= (layer2_outputs(1055)) and not (layer2_outputs(7166));
    layer3_outputs(638) <= '1';
    layer3_outputs(639) <= (layer2_outputs(5446)) and not (layer2_outputs(609));
    layer3_outputs(640) <= '0';
    layer3_outputs(641) <= (layer2_outputs(3399)) and (layer2_outputs(2902));
    layer3_outputs(642) <= '1';
    layer3_outputs(643) <= '1';
    layer3_outputs(644) <= not(layer2_outputs(127));
    layer3_outputs(645) <= not((layer2_outputs(3250)) and (layer2_outputs(6455)));
    layer3_outputs(646) <= '0';
    layer3_outputs(647) <= layer2_outputs(4410);
    layer3_outputs(648) <= not((layer2_outputs(2586)) or (layer2_outputs(6335)));
    layer3_outputs(649) <= (layer2_outputs(4406)) and not (layer2_outputs(6554));
    layer3_outputs(650) <= not((layer2_outputs(7389)) and (layer2_outputs(5375)));
    layer3_outputs(651) <= not(layer2_outputs(3054));
    layer3_outputs(652) <= not(layer2_outputs(2426)) or (layer2_outputs(6684));
    layer3_outputs(653) <= not(layer2_outputs(422));
    layer3_outputs(654) <= not(layer2_outputs(7366));
    layer3_outputs(655) <= layer2_outputs(4661);
    layer3_outputs(656) <= layer2_outputs(1136);
    layer3_outputs(657) <= (layer2_outputs(4351)) and (layer2_outputs(2532));
    layer3_outputs(658) <= not((layer2_outputs(5681)) and (layer2_outputs(7049)));
    layer3_outputs(659) <= not(layer2_outputs(583)) or (layer2_outputs(5458));
    layer3_outputs(660) <= not((layer2_outputs(2288)) xor (layer2_outputs(4247)));
    layer3_outputs(661) <= not((layer2_outputs(6160)) and (layer2_outputs(2588)));
    layer3_outputs(662) <= (layer2_outputs(4596)) or (layer2_outputs(5538));
    layer3_outputs(663) <= (layer2_outputs(6417)) and not (layer2_outputs(1758));
    layer3_outputs(664) <= (layer2_outputs(6033)) and not (layer2_outputs(3261));
    layer3_outputs(665) <= layer2_outputs(6403);
    layer3_outputs(666) <= not(layer2_outputs(6126));
    layer3_outputs(667) <= (layer2_outputs(1259)) and (layer2_outputs(5556));
    layer3_outputs(668) <= not(layer2_outputs(7432));
    layer3_outputs(669) <= not(layer2_outputs(6350)) or (layer2_outputs(734));
    layer3_outputs(670) <= not(layer2_outputs(7176));
    layer3_outputs(671) <= not((layer2_outputs(3571)) or (layer2_outputs(1865)));
    layer3_outputs(672) <= not(layer2_outputs(1670));
    layer3_outputs(673) <= not(layer2_outputs(1801));
    layer3_outputs(674) <= (layer2_outputs(2721)) or (layer2_outputs(4889));
    layer3_outputs(675) <= layer2_outputs(533);
    layer3_outputs(676) <= layer2_outputs(2054);
    layer3_outputs(677) <= not(layer2_outputs(4878)) or (layer2_outputs(2462));
    layer3_outputs(678) <= not((layer2_outputs(2576)) or (layer2_outputs(5436)));
    layer3_outputs(679) <= not(layer2_outputs(169));
    layer3_outputs(680) <= '0';
    layer3_outputs(681) <= layer2_outputs(6324);
    layer3_outputs(682) <= not((layer2_outputs(1906)) and (layer2_outputs(2374)));
    layer3_outputs(683) <= layer2_outputs(7588);
    layer3_outputs(684) <= not(layer2_outputs(5152));
    layer3_outputs(685) <= (layer2_outputs(950)) and not (layer2_outputs(1141));
    layer3_outputs(686) <= (layer2_outputs(6649)) and (layer2_outputs(5067));
    layer3_outputs(687) <= not(layer2_outputs(2598));
    layer3_outputs(688) <= layer2_outputs(6543);
    layer3_outputs(689) <= not(layer2_outputs(4720));
    layer3_outputs(690) <= (layer2_outputs(446)) and (layer2_outputs(2013));
    layer3_outputs(691) <= '0';
    layer3_outputs(692) <= (layer2_outputs(6634)) and not (layer2_outputs(5903));
    layer3_outputs(693) <= (layer2_outputs(7179)) and not (layer2_outputs(5346));
    layer3_outputs(694) <= not(layer2_outputs(6235));
    layer3_outputs(695) <= not(layer2_outputs(6198));
    layer3_outputs(696) <= layer2_outputs(1328);
    layer3_outputs(697) <= not((layer2_outputs(1496)) or (layer2_outputs(4134)));
    layer3_outputs(698) <= layer2_outputs(5342);
    layer3_outputs(699) <= (layer2_outputs(1800)) and (layer2_outputs(3765));
    layer3_outputs(700) <= layer2_outputs(5319);
    layer3_outputs(701) <= not(layer2_outputs(4374));
    layer3_outputs(702) <= (layer2_outputs(6825)) or (layer2_outputs(6657));
    layer3_outputs(703) <= layer2_outputs(1775);
    layer3_outputs(704) <= not(layer2_outputs(1174));
    layer3_outputs(705) <= not(layer2_outputs(1855));
    layer3_outputs(706) <= not(layer2_outputs(4827));
    layer3_outputs(707) <= not(layer2_outputs(5607)) or (layer2_outputs(1201));
    layer3_outputs(708) <= not((layer2_outputs(7032)) or (layer2_outputs(2262)));
    layer3_outputs(709) <= not(layer2_outputs(656)) or (layer2_outputs(6665));
    layer3_outputs(710) <= not((layer2_outputs(306)) or (layer2_outputs(654)));
    layer3_outputs(711) <= not((layer2_outputs(6486)) and (layer2_outputs(7227)));
    layer3_outputs(712) <= not((layer2_outputs(4773)) or (layer2_outputs(1676)));
    layer3_outputs(713) <= (layer2_outputs(4042)) and (layer2_outputs(6425));
    layer3_outputs(714) <= not((layer2_outputs(1496)) and (layer2_outputs(3780)));
    layer3_outputs(715) <= not(layer2_outputs(1827)) or (layer2_outputs(7355));
    layer3_outputs(716) <= not((layer2_outputs(2861)) or (layer2_outputs(4809)));
    layer3_outputs(717) <= '1';
    layer3_outputs(718) <= not(layer2_outputs(4573));
    layer3_outputs(719) <= not(layer2_outputs(286));
    layer3_outputs(720) <= not(layer2_outputs(6570));
    layer3_outputs(721) <= not(layer2_outputs(6182));
    layer3_outputs(722) <= '0';
    layer3_outputs(723) <= (layer2_outputs(701)) and not (layer2_outputs(7652));
    layer3_outputs(724) <= not(layer2_outputs(4022)) or (layer2_outputs(2668));
    layer3_outputs(725) <= (layer2_outputs(6008)) and (layer2_outputs(6170));
    layer3_outputs(726) <= layer2_outputs(285);
    layer3_outputs(727) <= not((layer2_outputs(1867)) xor (layer2_outputs(7268)));
    layer3_outputs(728) <= not((layer2_outputs(3816)) xor (layer2_outputs(6294)));
    layer3_outputs(729) <= not((layer2_outputs(1135)) or (layer2_outputs(1626)));
    layer3_outputs(730) <= (layer2_outputs(2259)) and not (layer2_outputs(3922));
    layer3_outputs(731) <= (layer2_outputs(1228)) or (layer2_outputs(459));
    layer3_outputs(732) <= (layer2_outputs(3675)) or (layer2_outputs(7470));
    layer3_outputs(733) <= (layer2_outputs(3050)) and not (layer2_outputs(5842));
    layer3_outputs(734) <= not(layer2_outputs(3216)) or (layer2_outputs(6017));
    layer3_outputs(735) <= not(layer2_outputs(7385));
    layer3_outputs(736) <= not(layer2_outputs(5333));
    layer3_outputs(737) <= not((layer2_outputs(2925)) and (layer2_outputs(7321)));
    layer3_outputs(738) <= (layer2_outputs(3879)) or (layer2_outputs(2702));
    layer3_outputs(739) <= not((layer2_outputs(647)) or (layer2_outputs(2173)));
    layer3_outputs(740) <= not((layer2_outputs(5181)) or (layer2_outputs(1464)));
    layer3_outputs(741) <= (layer2_outputs(3639)) and not (layer2_outputs(4768));
    layer3_outputs(742) <= not(layer2_outputs(4967)) or (layer2_outputs(6227));
    layer3_outputs(743) <= (layer2_outputs(378)) and not (layer2_outputs(3313));
    layer3_outputs(744) <= layer2_outputs(2867);
    layer3_outputs(745) <= (layer2_outputs(6774)) and not (layer2_outputs(5901));
    layer3_outputs(746) <= not(layer2_outputs(6958));
    layer3_outputs(747) <= layer2_outputs(326);
    layer3_outputs(748) <= layer2_outputs(2676);
    layer3_outputs(749) <= layer2_outputs(4211);
    layer3_outputs(750) <= layer2_outputs(1691);
    layer3_outputs(751) <= (layer2_outputs(3463)) or (layer2_outputs(2549));
    layer3_outputs(752) <= layer2_outputs(1886);
    layer3_outputs(753) <= (layer2_outputs(943)) and not (layer2_outputs(3595));
    layer3_outputs(754) <= '0';
    layer3_outputs(755) <= '0';
    layer3_outputs(756) <= layer2_outputs(1161);
    layer3_outputs(757) <= layer2_outputs(3001);
    layer3_outputs(758) <= (layer2_outputs(6610)) and not (layer2_outputs(445));
    layer3_outputs(759) <= not(layer2_outputs(1267)) or (layer2_outputs(6716));
    layer3_outputs(760) <= (layer2_outputs(6015)) and not (layer2_outputs(5565));
    layer3_outputs(761) <= not((layer2_outputs(5964)) and (layer2_outputs(7202)));
    layer3_outputs(762) <= (layer2_outputs(3500)) and (layer2_outputs(1643));
    layer3_outputs(763) <= (layer2_outputs(7253)) and not (layer2_outputs(3683));
    layer3_outputs(764) <= not(layer2_outputs(7078));
    layer3_outputs(765) <= not((layer2_outputs(3225)) or (layer2_outputs(1611)));
    layer3_outputs(766) <= not((layer2_outputs(3876)) and (layer2_outputs(7324)));
    layer3_outputs(767) <= layer2_outputs(4068);
    layer3_outputs(768) <= (layer2_outputs(3428)) and not (layer2_outputs(5511));
    layer3_outputs(769) <= not(layer2_outputs(3225));
    layer3_outputs(770) <= layer2_outputs(573);
    layer3_outputs(771) <= not(layer2_outputs(586));
    layer3_outputs(772) <= layer2_outputs(7550);
    layer3_outputs(773) <= (layer2_outputs(1905)) or (layer2_outputs(1851));
    layer3_outputs(774) <= (layer2_outputs(6934)) and not (layer2_outputs(2382));
    layer3_outputs(775) <= not(layer2_outputs(1403));
    layer3_outputs(776) <= not(layer2_outputs(5797)) or (layer2_outputs(4678));
    layer3_outputs(777) <= not((layer2_outputs(2025)) or (layer2_outputs(1300)));
    layer3_outputs(778) <= not(layer2_outputs(364)) or (layer2_outputs(577));
    layer3_outputs(779) <= not((layer2_outputs(6622)) or (layer2_outputs(1229)));
    layer3_outputs(780) <= not(layer2_outputs(6897));
    layer3_outputs(781) <= not(layer2_outputs(6041));
    layer3_outputs(782) <= (layer2_outputs(1542)) or (layer2_outputs(4505));
    layer3_outputs(783) <= (layer2_outputs(27)) xor (layer2_outputs(1363));
    layer3_outputs(784) <= layer2_outputs(4098);
    layer3_outputs(785) <= not((layer2_outputs(1442)) and (layer2_outputs(7009)));
    layer3_outputs(786) <= '0';
    layer3_outputs(787) <= layer2_outputs(2588);
    layer3_outputs(788) <= (layer2_outputs(4887)) and not (layer2_outputs(4897));
    layer3_outputs(789) <= '1';
    layer3_outputs(790) <= layer2_outputs(6672);
    layer3_outputs(791) <= not(layer2_outputs(3488)) or (layer2_outputs(7245));
    layer3_outputs(792) <= (layer2_outputs(3260)) and not (layer2_outputs(4913));
    layer3_outputs(793) <= layer2_outputs(263);
    layer3_outputs(794) <= (layer2_outputs(4107)) and (layer2_outputs(4237));
    layer3_outputs(795) <= not((layer2_outputs(7292)) and (layer2_outputs(4832)));
    layer3_outputs(796) <= layer2_outputs(2174);
    layer3_outputs(797) <= layer2_outputs(4957);
    layer3_outputs(798) <= not((layer2_outputs(6563)) and (layer2_outputs(5683)));
    layer3_outputs(799) <= not(layer2_outputs(3482)) or (layer2_outputs(5150));
    layer3_outputs(800) <= (layer2_outputs(5029)) or (layer2_outputs(63));
    layer3_outputs(801) <= '0';
    layer3_outputs(802) <= not(layer2_outputs(761));
    layer3_outputs(803) <= not(layer2_outputs(5543)) or (layer2_outputs(723));
    layer3_outputs(804) <= layer2_outputs(2623);
    layer3_outputs(805) <= '0';
    layer3_outputs(806) <= not(layer2_outputs(23));
    layer3_outputs(807) <= not(layer2_outputs(4625));
    layer3_outputs(808) <= (layer2_outputs(5402)) and not (layer2_outputs(5336));
    layer3_outputs(809) <= (layer2_outputs(5658)) and not (layer2_outputs(3694));
    layer3_outputs(810) <= '1';
    layer3_outputs(811) <= not((layer2_outputs(2871)) and (layer2_outputs(5967)));
    layer3_outputs(812) <= not(layer2_outputs(5412));
    layer3_outputs(813) <= '0';
    layer3_outputs(814) <= not(layer2_outputs(4059));
    layer3_outputs(815) <= layer2_outputs(313);
    layer3_outputs(816) <= not(layer2_outputs(7215));
    layer3_outputs(817) <= layer2_outputs(5626);
    layer3_outputs(818) <= not((layer2_outputs(4742)) or (layer2_outputs(3923)));
    layer3_outputs(819) <= not(layer2_outputs(6236)) or (layer2_outputs(1575));
    layer3_outputs(820) <= not(layer2_outputs(2410));
    layer3_outputs(821) <= not(layer2_outputs(3117)) or (layer2_outputs(1339));
    layer3_outputs(822) <= layer2_outputs(5655);
    layer3_outputs(823) <= not((layer2_outputs(5962)) or (layer2_outputs(85)));
    layer3_outputs(824) <= not(layer2_outputs(44));
    layer3_outputs(825) <= not(layer2_outputs(5255)) or (layer2_outputs(1168));
    layer3_outputs(826) <= (layer2_outputs(483)) and not (layer2_outputs(2484));
    layer3_outputs(827) <= '1';
    layer3_outputs(828) <= not(layer2_outputs(1642));
    layer3_outputs(829) <= not(layer2_outputs(1233));
    layer3_outputs(830) <= not(layer2_outputs(5443));
    layer3_outputs(831) <= '1';
    layer3_outputs(832) <= (layer2_outputs(7384)) and not (layer2_outputs(4934));
    layer3_outputs(833) <= not((layer2_outputs(3844)) and (layer2_outputs(3749)));
    layer3_outputs(834) <= not(layer2_outputs(2093));
    layer3_outputs(835) <= (layer2_outputs(7173)) and not (layer2_outputs(2240));
    layer3_outputs(836) <= not(layer2_outputs(1773));
    layer3_outputs(837) <= '0';
    layer3_outputs(838) <= (layer2_outputs(4740)) and (layer2_outputs(7236));
    layer3_outputs(839) <= '0';
    layer3_outputs(840) <= not(layer2_outputs(1825));
    layer3_outputs(841) <= not(layer2_outputs(6354));
    layer3_outputs(842) <= layer2_outputs(2840);
    layer3_outputs(843) <= not(layer2_outputs(272));
    layer3_outputs(844) <= not(layer2_outputs(4464)) or (layer2_outputs(2431));
    layer3_outputs(845) <= not(layer2_outputs(7632));
    layer3_outputs(846) <= not(layer2_outputs(2002));
    layer3_outputs(847) <= not((layer2_outputs(5276)) xor (layer2_outputs(6111)));
    layer3_outputs(848) <= (layer2_outputs(1205)) or (layer2_outputs(7076));
    layer3_outputs(849) <= not((layer2_outputs(3058)) or (layer2_outputs(2563)));
    layer3_outputs(850) <= not(layer2_outputs(6066));
    layer3_outputs(851) <= '0';
    layer3_outputs(852) <= layer2_outputs(409);
    layer3_outputs(853) <= not(layer2_outputs(4179)) or (layer2_outputs(7574));
    layer3_outputs(854) <= (layer2_outputs(5147)) or (layer2_outputs(2887));
    layer3_outputs(855) <= not(layer2_outputs(5692));
    layer3_outputs(856) <= layer2_outputs(3220);
    layer3_outputs(857) <= not(layer2_outputs(6860));
    layer3_outputs(858) <= layer2_outputs(6083);
    layer3_outputs(859) <= not((layer2_outputs(3246)) and (layer2_outputs(76)));
    layer3_outputs(860) <= not((layer2_outputs(3933)) xor (layer2_outputs(2917)));
    layer3_outputs(861) <= layer2_outputs(5271);
    layer3_outputs(862) <= '1';
    layer3_outputs(863) <= not(layer2_outputs(7009));
    layer3_outputs(864) <= (layer2_outputs(7590)) and not (layer2_outputs(6810));
    layer3_outputs(865) <= not((layer2_outputs(4272)) and (layer2_outputs(4471)));
    layer3_outputs(866) <= not((layer2_outputs(503)) or (layer2_outputs(2573)));
    layer3_outputs(867) <= layer2_outputs(3385);
    layer3_outputs(868) <= not(layer2_outputs(3614));
    layer3_outputs(869) <= not(layer2_outputs(4541));
    layer3_outputs(870) <= (layer2_outputs(7581)) and (layer2_outputs(7593));
    layer3_outputs(871) <= not(layer2_outputs(3242)) or (layer2_outputs(3258));
    layer3_outputs(872) <= not(layer2_outputs(5445));
    layer3_outputs(873) <= not(layer2_outputs(2281)) or (layer2_outputs(565));
    layer3_outputs(874) <= not(layer2_outputs(4332));
    layer3_outputs(875) <= layer2_outputs(1416);
    layer3_outputs(876) <= layer2_outputs(5979);
    layer3_outputs(877) <= not(layer2_outputs(5710));
    layer3_outputs(878) <= '1';
    layer3_outputs(879) <= '1';
    layer3_outputs(880) <= not(layer2_outputs(5541)) or (layer2_outputs(3317));
    layer3_outputs(881) <= layer2_outputs(383);
    layer3_outputs(882) <= (layer2_outputs(1283)) and not (layer2_outputs(7017));
    layer3_outputs(883) <= (layer2_outputs(186)) and not (layer2_outputs(1973));
    layer3_outputs(884) <= (layer2_outputs(6370)) or (layer2_outputs(6839));
    layer3_outputs(885) <= (layer2_outputs(96)) xor (layer2_outputs(3805));
    layer3_outputs(886) <= not(layer2_outputs(7040));
    layer3_outputs(887) <= layer2_outputs(5871);
    layer3_outputs(888) <= not(layer2_outputs(4093));
    layer3_outputs(889) <= not(layer2_outputs(6336));
    layer3_outputs(890) <= layer2_outputs(438);
    layer3_outputs(891) <= (layer2_outputs(4723)) and (layer2_outputs(2324));
    layer3_outputs(892) <= '0';
    layer3_outputs(893) <= not((layer2_outputs(1814)) or (layer2_outputs(5418)));
    layer3_outputs(894) <= '0';
    layer3_outputs(895) <= not(layer2_outputs(5459));
    layer3_outputs(896) <= not(layer2_outputs(2031)) or (layer2_outputs(2028));
    layer3_outputs(897) <= layer2_outputs(502);
    layer3_outputs(898) <= layer2_outputs(1003);
    layer3_outputs(899) <= (layer2_outputs(1939)) and not (layer2_outputs(4303));
    layer3_outputs(900) <= (layer2_outputs(4111)) and not (layer2_outputs(7381));
    layer3_outputs(901) <= (layer2_outputs(4724)) and not (layer2_outputs(5513));
    layer3_outputs(902) <= '0';
    layer3_outputs(903) <= layer2_outputs(6360);
    layer3_outputs(904) <= not(layer2_outputs(1043)) or (layer2_outputs(3368));
    layer3_outputs(905) <= not((layer2_outputs(3329)) and (layer2_outputs(733)));
    layer3_outputs(906) <= not((layer2_outputs(2873)) or (layer2_outputs(2130)));
    layer3_outputs(907) <= (layer2_outputs(3261)) and not (layer2_outputs(2039));
    layer3_outputs(908) <= (layer2_outputs(6074)) and not (layer2_outputs(4141));
    layer3_outputs(909) <= layer2_outputs(2851);
    layer3_outputs(910) <= not(layer2_outputs(890)) or (layer2_outputs(4568));
    layer3_outputs(911) <= not((layer2_outputs(4229)) or (layer2_outputs(25)));
    layer3_outputs(912) <= not(layer2_outputs(2689)) or (layer2_outputs(2132));
    layer3_outputs(913) <= not((layer2_outputs(4244)) and (layer2_outputs(1466)));
    layer3_outputs(914) <= (layer2_outputs(7437)) xor (layer2_outputs(3175));
    layer3_outputs(915) <= (layer2_outputs(6650)) and not (layer2_outputs(6555));
    layer3_outputs(916) <= (layer2_outputs(3121)) and not (layer2_outputs(982));
    layer3_outputs(917) <= layer2_outputs(3427);
    layer3_outputs(918) <= not(layer2_outputs(1401));
    layer3_outputs(919) <= '0';
    layer3_outputs(920) <= not((layer2_outputs(5348)) or (layer2_outputs(936)));
    layer3_outputs(921) <= (layer2_outputs(2525)) and not (layer2_outputs(4606));
    layer3_outputs(922) <= not(layer2_outputs(6040));
    layer3_outputs(923) <= not(layer2_outputs(5586)) or (layer2_outputs(7180));
    layer3_outputs(924) <= layer2_outputs(6357);
    layer3_outputs(925) <= (layer2_outputs(5434)) and not (layer2_outputs(4791));
    layer3_outputs(926) <= '1';
    layer3_outputs(927) <= layer2_outputs(991);
    layer3_outputs(928) <= layer2_outputs(5151);
    layer3_outputs(929) <= '0';
    layer3_outputs(930) <= '0';
    layer3_outputs(931) <= '0';
    layer3_outputs(932) <= (layer2_outputs(6258)) and not (layer2_outputs(6647));
    layer3_outputs(933) <= (layer2_outputs(4793)) and (layer2_outputs(7339));
    layer3_outputs(934) <= not(layer2_outputs(1415));
    layer3_outputs(935) <= layer2_outputs(6081);
    layer3_outputs(936) <= '1';
    layer3_outputs(937) <= not(layer2_outputs(3265));
    layer3_outputs(938) <= not(layer2_outputs(5095));
    layer3_outputs(939) <= (layer2_outputs(41)) and (layer2_outputs(7550));
    layer3_outputs(940) <= not(layer2_outputs(3359));
    layer3_outputs(941) <= not((layer2_outputs(1735)) or (layer2_outputs(5692)));
    layer3_outputs(942) <= (layer2_outputs(3336)) or (layer2_outputs(3408));
    layer3_outputs(943) <= not(layer2_outputs(7457));
    layer3_outputs(944) <= '0';
    layer3_outputs(945) <= not((layer2_outputs(418)) or (layer2_outputs(3166)));
    layer3_outputs(946) <= (layer2_outputs(1037)) and (layer2_outputs(2250));
    layer3_outputs(947) <= (layer2_outputs(2133)) and (layer2_outputs(4113));
    layer3_outputs(948) <= '1';
    layer3_outputs(949) <= (layer2_outputs(1189)) and (layer2_outputs(1200));
    layer3_outputs(950) <= '0';
    layer3_outputs(951) <= layer2_outputs(2464);
    layer3_outputs(952) <= not(layer2_outputs(1397)) or (layer2_outputs(1102));
    layer3_outputs(953) <= (layer2_outputs(1028)) and not (layer2_outputs(6634));
    layer3_outputs(954) <= not((layer2_outputs(5835)) or (layer2_outputs(5396)));
    layer3_outputs(955) <= (layer2_outputs(1341)) and (layer2_outputs(3150));
    layer3_outputs(956) <= layer2_outputs(7250);
    layer3_outputs(957) <= not(layer2_outputs(742)) or (layer2_outputs(6658));
    layer3_outputs(958) <= not(layer2_outputs(3008)) or (layer2_outputs(934));
    layer3_outputs(959) <= not((layer2_outputs(3449)) and (layer2_outputs(3594)));
    layer3_outputs(960) <= not(layer2_outputs(3920));
    layer3_outputs(961) <= not(layer2_outputs(540)) or (layer2_outputs(6094));
    layer3_outputs(962) <= (layer2_outputs(5503)) and (layer2_outputs(1349));
    layer3_outputs(963) <= '0';
    layer3_outputs(964) <= layer2_outputs(652);
    layer3_outputs(965) <= (layer2_outputs(2478)) xor (layer2_outputs(3172));
    layer3_outputs(966) <= (layer2_outputs(6268)) or (layer2_outputs(3761));
    layer3_outputs(967) <= (layer2_outputs(2521)) and not (layer2_outputs(3432));
    layer3_outputs(968) <= layer2_outputs(4508);
    layer3_outputs(969) <= not(layer2_outputs(7431));
    layer3_outputs(970) <= not(layer2_outputs(3110));
    layer3_outputs(971) <= layer2_outputs(1126);
    layer3_outputs(972) <= '0';
    layer3_outputs(973) <= (layer2_outputs(5733)) and (layer2_outputs(2148));
    layer3_outputs(974) <= (layer2_outputs(4210)) and not (layer2_outputs(1358));
    layer3_outputs(975) <= not(layer2_outputs(5755)) or (layer2_outputs(84));
    layer3_outputs(976) <= (layer2_outputs(6792)) or (layer2_outputs(1172));
    layer3_outputs(977) <= '0';
    layer3_outputs(978) <= not(layer2_outputs(5022));
    layer3_outputs(979) <= not(layer2_outputs(1152));
    layer3_outputs(980) <= layer2_outputs(7448);
    layer3_outputs(981) <= not(layer2_outputs(6999));
    layer3_outputs(982) <= not(layer2_outputs(663));
    layer3_outputs(983) <= not(layer2_outputs(3435));
    layer3_outputs(984) <= layer2_outputs(2879);
    layer3_outputs(985) <= not(layer2_outputs(7589));
    layer3_outputs(986) <= layer2_outputs(4970);
    layer3_outputs(987) <= not(layer2_outputs(6519)) or (layer2_outputs(2622));
    layer3_outputs(988) <= not(layer2_outputs(453)) or (layer2_outputs(2296));
    layer3_outputs(989) <= not(layer2_outputs(1551)) or (layer2_outputs(1812));
    layer3_outputs(990) <= layer2_outputs(1773);
    layer3_outputs(991) <= layer2_outputs(3656);
    layer3_outputs(992) <= not((layer2_outputs(6949)) xor (layer2_outputs(6538)));
    layer3_outputs(993) <= not((layer2_outputs(3383)) and (layer2_outputs(6556)));
    layer3_outputs(994) <= layer2_outputs(1129);
    layer3_outputs(995) <= (layer2_outputs(6902)) and (layer2_outputs(1896));
    layer3_outputs(996) <= not(layer2_outputs(4991)) or (layer2_outputs(1509));
    layer3_outputs(997) <= not((layer2_outputs(3138)) xor (layer2_outputs(2799)));
    layer3_outputs(998) <= (layer2_outputs(1528)) and (layer2_outputs(6557));
    layer3_outputs(999) <= not((layer2_outputs(4158)) xor (layer2_outputs(2821)));
    layer3_outputs(1000) <= not(layer2_outputs(2409)) or (layer2_outputs(3944));
    layer3_outputs(1001) <= not(layer2_outputs(3061));
    layer3_outputs(1002) <= not(layer2_outputs(1784)) or (layer2_outputs(69));
    layer3_outputs(1003) <= layer2_outputs(7216);
    layer3_outputs(1004) <= (layer2_outputs(5295)) or (layer2_outputs(1012));
    layer3_outputs(1005) <= not((layer2_outputs(6187)) or (layer2_outputs(4837)));
    layer3_outputs(1006) <= layer2_outputs(4835);
    layer3_outputs(1007) <= (layer2_outputs(3804)) and not (layer2_outputs(4356));
    layer3_outputs(1008) <= (layer2_outputs(2912)) and not (layer2_outputs(2974));
    layer3_outputs(1009) <= not(layer2_outputs(4269)) or (layer2_outputs(5308));
    layer3_outputs(1010) <= layer2_outputs(3665);
    layer3_outputs(1011) <= layer2_outputs(3185);
    layer3_outputs(1012) <= (layer2_outputs(1142)) xor (layer2_outputs(5942));
    layer3_outputs(1013) <= '1';
    layer3_outputs(1014) <= not(layer2_outputs(4420));
    layer3_outputs(1015) <= '0';
    layer3_outputs(1016) <= not(layer2_outputs(6422)) or (layer2_outputs(1411));
    layer3_outputs(1017) <= not(layer2_outputs(2922));
    layer3_outputs(1018) <= (layer2_outputs(7213)) and (layer2_outputs(97));
    layer3_outputs(1019) <= '0';
    layer3_outputs(1020) <= (layer2_outputs(4994)) and not (layer2_outputs(933));
    layer3_outputs(1021) <= not(layer2_outputs(701)) or (layer2_outputs(7372));
    layer3_outputs(1022) <= layer2_outputs(5202);
    layer3_outputs(1023) <= not(layer2_outputs(6296)) or (layer2_outputs(3028));
    layer3_outputs(1024) <= '0';
    layer3_outputs(1025) <= (layer2_outputs(4499)) and (layer2_outputs(5674));
    layer3_outputs(1026) <= not(layer2_outputs(4169)) or (layer2_outputs(5403));
    layer3_outputs(1027) <= '1';
    layer3_outputs(1028) <= not((layer2_outputs(1179)) or (layer2_outputs(6897)));
    layer3_outputs(1029) <= (layer2_outputs(6095)) and not (layer2_outputs(6197));
    layer3_outputs(1030) <= layer2_outputs(4288);
    layer3_outputs(1031) <= not(layer2_outputs(7299)) or (layer2_outputs(5974));
    layer3_outputs(1032) <= not((layer2_outputs(2603)) and (layer2_outputs(2252)));
    layer3_outputs(1033) <= not((layer2_outputs(4454)) and (layer2_outputs(2536)));
    layer3_outputs(1034) <= not((layer2_outputs(649)) or (layer2_outputs(486)));
    layer3_outputs(1035) <= layer2_outputs(5856);
    layer3_outputs(1036) <= (layer2_outputs(5212)) and not (layer2_outputs(937));
    layer3_outputs(1037) <= layer2_outputs(2797);
    layer3_outputs(1038) <= (layer2_outputs(5133)) or (layer2_outputs(4178));
    layer3_outputs(1039) <= '0';
    layer3_outputs(1040) <= layer2_outputs(633);
    layer3_outputs(1041) <= (layer2_outputs(6052)) and not (layer2_outputs(5745));
    layer3_outputs(1042) <= not((layer2_outputs(4451)) or (layer2_outputs(5634)));
    layer3_outputs(1043) <= '1';
    layer3_outputs(1044) <= not((layer2_outputs(7668)) or (layer2_outputs(6935)));
    layer3_outputs(1045) <= (layer2_outputs(4598)) and not (layer2_outputs(7424));
    layer3_outputs(1046) <= not(layer2_outputs(5146));
    layer3_outputs(1047) <= layer2_outputs(817);
    layer3_outputs(1048) <= (layer2_outputs(2469)) and not (layer2_outputs(3031));
    layer3_outputs(1049) <= not((layer2_outputs(4441)) and (layer2_outputs(2000)));
    layer3_outputs(1050) <= layer2_outputs(5506);
    layer3_outputs(1051) <= layer2_outputs(4727);
    layer3_outputs(1052) <= (layer2_outputs(1353)) or (layer2_outputs(2741));
    layer3_outputs(1053) <= not((layer2_outputs(6621)) or (layer2_outputs(838)));
    layer3_outputs(1054) <= (layer2_outputs(3284)) and not (layer2_outputs(4665));
    layer3_outputs(1055) <= not(layer2_outputs(2109));
    layer3_outputs(1056) <= not(layer2_outputs(765)) or (layer2_outputs(123));
    layer3_outputs(1057) <= (layer2_outputs(4875)) and not (layer2_outputs(3542));
    layer3_outputs(1058) <= not((layer2_outputs(4726)) or (layer2_outputs(5843)));
    layer3_outputs(1059) <= not(layer2_outputs(5762)) or (layer2_outputs(6627));
    layer3_outputs(1060) <= not((layer2_outputs(7153)) or (layer2_outputs(6816)));
    layer3_outputs(1061) <= (layer2_outputs(4570)) and not (layer2_outputs(6591));
    layer3_outputs(1062) <= layer2_outputs(2411);
    layer3_outputs(1063) <= (layer2_outputs(7145)) and (layer2_outputs(7631));
    layer3_outputs(1064) <= layer2_outputs(6443);
    layer3_outputs(1065) <= layer2_outputs(1943);
    layer3_outputs(1066) <= (layer2_outputs(2188)) and (layer2_outputs(4226));
    layer3_outputs(1067) <= not(layer2_outputs(7375));
    layer3_outputs(1068) <= not(layer2_outputs(4800)) or (layer2_outputs(7524));
    layer3_outputs(1069) <= layer2_outputs(7563);
    layer3_outputs(1070) <= (layer2_outputs(2849)) and not (layer2_outputs(4510));
    layer3_outputs(1071) <= not((layer2_outputs(1387)) and (layer2_outputs(4603)));
    layer3_outputs(1072) <= layer2_outputs(5600);
    layer3_outputs(1073) <= (layer2_outputs(1519)) or (layer2_outputs(337));
    layer3_outputs(1074) <= '1';
    layer3_outputs(1075) <= (layer2_outputs(2486)) and not (layer2_outputs(1251));
    layer3_outputs(1076) <= not(layer2_outputs(5611)) or (layer2_outputs(3527));
    layer3_outputs(1077) <= '1';
    layer3_outputs(1078) <= layer2_outputs(5954);
    layer3_outputs(1079) <= (layer2_outputs(5866)) or (layer2_outputs(1275));
    layer3_outputs(1080) <= '0';
    layer3_outputs(1081) <= (layer2_outputs(1497)) and not (layer2_outputs(535));
    layer3_outputs(1082) <= layer2_outputs(2268);
    layer3_outputs(1083) <= not(layer2_outputs(1958));
    layer3_outputs(1084) <= (layer2_outputs(2332)) or (layer2_outputs(6534));
    layer3_outputs(1085) <= not((layer2_outputs(1511)) xor (layer2_outputs(6164)));
    layer3_outputs(1086) <= not((layer2_outputs(6951)) and (layer2_outputs(7574)));
    layer3_outputs(1087) <= not((layer2_outputs(567)) or (layer2_outputs(2099)));
    layer3_outputs(1088) <= '1';
    layer3_outputs(1089) <= (layer2_outputs(6243)) and (layer2_outputs(3615));
    layer3_outputs(1090) <= not((layer2_outputs(5897)) and (layer2_outputs(1159)));
    layer3_outputs(1091) <= '1';
    layer3_outputs(1092) <= layer2_outputs(1913);
    layer3_outputs(1093) <= layer2_outputs(7);
    layer3_outputs(1094) <= '0';
    layer3_outputs(1095) <= (layer2_outputs(6257)) and (layer2_outputs(6921));
    layer3_outputs(1096) <= (layer2_outputs(6359)) and not (layer2_outputs(5036));
    layer3_outputs(1097) <= not(layer2_outputs(3589));
    layer3_outputs(1098) <= (layer2_outputs(267)) and not (layer2_outputs(5930));
    layer3_outputs(1099) <= layer2_outputs(1402);
    layer3_outputs(1100) <= layer2_outputs(4087);
    layer3_outputs(1101) <= (layer2_outputs(5993)) and (layer2_outputs(161));
    layer3_outputs(1102) <= layer2_outputs(4176);
    layer3_outputs(1103) <= (layer2_outputs(3575)) and not (layer2_outputs(6630));
    layer3_outputs(1104) <= not((layer2_outputs(5767)) or (layer2_outputs(2655)));
    layer3_outputs(1105) <= not(layer2_outputs(7249));
    layer3_outputs(1106) <= (layer2_outputs(2402)) and not (layer2_outputs(1292));
    layer3_outputs(1107) <= (layer2_outputs(4824)) and (layer2_outputs(6301));
    layer3_outputs(1108) <= layer2_outputs(3023);
    layer3_outputs(1109) <= '1';
    layer3_outputs(1110) <= (layer2_outputs(1793)) and not (layer2_outputs(7002));
    layer3_outputs(1111) <= (layer2_outputs(1622)) and (layer2_outputs(2811));
    layer3_outputs(1112) <= not(layer2_outputs(4156));
    layer3_outputs(1113) <= not(layer2_outputs(4783)) or (layer2_outputs(5985));
    layer3_outputs(1114) <= layer2_outputs(6905);
    layer3_outputs(1115) <= layer2_outputs(3430);
    layer3_outputs(1116) <= '0';
    layer3_outputs(1117) <= (layer2_outputs(1132)) or (layer2_outputs(7210));
    layer3_outputs(1118) <= (layer2_outputs(2748)) and not (layer2_outputs(512));
    layer3_outputs(1119) <= layer2_outputs(7029);
    layer3_outputs(1120) <= layer2_outputs(7596);
    layer3_outputs(1121) <= '0';
    layer3_outputs(1122) <= not(layer2_outputs(599));
    layer3_outputs(1123) <= not(layer2_outputs(3772)) or (layer2_outputs(1600));
    layer3_outputs(1124) <= '0';
    layer3_outputs(1125) <= not((layer2_outputs(1509)) or (layer2_outputs(4920)));
    layer3_outputs(1126) <= layer2_outputs(785);
    layer3_outputs(1127) <= '0';
    layer3_outputs(1128) <= not(layer2_outputs(2450)) or (layer2_outputs(4746));
    layer3_outputs(1129) <= not((layer2_outputs(2104)) or (layer2_outputs(7571)));
    layer3_outputs(1130) <= not((layer2_outputs(1742)) and (layer2_outputs(1386)));
    layer3_outputs(1131) <= not(layer2_outputs(4647));
    layer3_outputs(1132) <= not(layer2_outputs(2724));
    layer3_outputs(1133) <= layer2_outputs(1221);
    layer3_outputs(1134) <= not(layer2_outputs(5304));
    layer3_outputs(1135) <= not((layer2_outputs(5261)) and (layer2_outputs(2004)));
    layer3_outputs(1136) <= not(layer2_outputs(5331)) or (layer2_outputs(2466));
    layer3_outputs(1137) <= not((layer2_outputs(5663)) or (layer2_outputs(6095)));
    layer3_outputs(1138) <= layer2_outputs(3096);
    layer3_outputs(1139) <= (layer2_outputs(7136)) or (layer2_outputs(4078));
    layer3_outputs(1140) <= (layer2_outputs(4603)) and not (layer2_outputs(3492));
    layer3_outputs(1141) <= (layer2_outputs(6938)) and not (layer2_outputs(1709));
    layer3_outputs(1142) <= layer2_outputs(4751);
    layer3_outputs(1143) <= layer2_outputs(6239);
    layer3_outputs(1144) <= not((layer2_outputs(5013)) or (layer2_outputs(3190)));
    layer3_outputs(1145) <= '1';
    layer3_outputs(1146) <= not((layer2_outputs(2902)) or (layer2_outputs(5533)));
    layer3_outputs(1147) <= '0';
    layer3_outputs(1148) <= layer2_outputs(1111);
    layer3_outputs(1149) <= not(layer2_outputs(7345));
    layer3_outputs(1150) <= not((layer2_outputs(1595)) and (layer2_outputs(5899)));
    layer3_outputs(1151) <= not(layer2_outputs(6388));
    layer3_outputs(1152) <= layer2_outputs(3235);
    layer3_outputs(1153) <= not(layer2_outputs(5401));
    layer3_outputs(1154) <= (layer2_outputs(3136)) and (layer2_outputs(605));
    layer3_outputs(1155) <= not(layer2_outputs(1));
    layer3_outputs(1156) <= not((layer2_outputs(2144)) or (layer2_outputs(2001)));
    layer3_outputs(1157) <= not(layer2_outputs(2212)) or (layer2_outputs(1897));
    layer3_outputs(1158) <= not(layer2_outputs(5802));
    layer3_outputs(1159) <= layer2_outputs(7420);
    layer3_outputs(1160) <= (layer2_outputs(908)) and (layer2_outputs(5943));
    layer3_outputs(1161) <= not(layer2_outputs(4689)) or (layer2_outputs(4887));
    layer3_outputs(1162) <= not((layer2_outputs(407)) and (layer2_outputs(7438)));
    layer3_outputs(1163) <= (layer2_outputs(2670)) and not (layer2_outputs(1923));
    layer3_outputs(1164) <= '0';
    layer3_outputs(1165) <= (layer2_outputs(4170)) and (layer2_outputs(7197));
    layer3_outputs(1166) <= not(layer2_outputs(4174));
    layer3_outputs(1167) <= (layer2_outputs(6565)) and (layer2_outputs(6618));
    layer3_outputs(1168) <= not((layer2_outputs(7545)) or (layer2_outputs(148)));
    layer3_outputs(1169) <= not(layer2_outputs(2837));
    layer3_outputs(1170) <= not(layer2_outputs(3449)) or (layer2_outputs(5979));
    layer3_outputs(1171) <= (layer2_outputs(1210)) and not (layer2_outputs(317));
    layer3_outputs(1172) <= (layer2_outputs(6488)) and not (layer2_outputs(398));
    layer3_outputs(1173) <= (layer2_outputs(3402)) and not (layer2_outputs(4669));
    layer3_outputs(1174) <= not(layer2_outputs(1818));
    layer3_outputs(1175) <= not((layer2_outputs(2653)) and (layer2_outputs(3894)));
    layer3_outputs(1176) <= not((layer2_outputs(3378)) and (layer2_outputs(2281)));
    layer3_outputs(1177) <= not(layer2_outputs(2176)) or (layer2_outputs(2608));
    layer3_outputs(1178) <= not((layer2_outputs(1898)) xor (layer2_outputs(347)));
    layer3_outputs(1179) <= (layer2_outputs(3188)) or (layer2_outputs(3));
    layer3_outputs(1180) <= not(layer2_outputs(2312)) or (layer2_outputs(6803));
    layer3_outputs(1181) <= not(layer2_outputs(2649));
    layer3_outputs(1182) <= not(layer2_outputs(5840));
    layer3_outputs(1183) <= layer2_outputs(7182);
    layer3_outputs(1184) <= '1';
    layer3_outputs(1185) <= not(layer2_outputs(2692)) or (layer2_outputs(413));
    layer3_outputs(1186) <= not((layer2_outputs(329)) xor (layer2_outputs(7021)));
    layer3_outputs(1187) <= layer2_outputs(4347);
    layer3_outputs(1188) <= '0';
    layer3_outputs(1189) <= not(layer2_outputs(331));
    layer3_outputs(1190) <= not(layer2_outputs(3130));
    layer3_outputs(1191) <= not(layer2_outputs(3255)) or (layer2_outputs(959));
    layer3_outputs(1192) <= not(layer2_outputs(3318)) or (layer2_outputs(2380));
    layer3_outputs(1193) <= not((layer2_outputs(3515)) and (layer2_outputs(1410)));
    layer3_outputs(1194) <= (layer2_outputs(754)) or (layer2_outputs(3326));
    layer3_outputs(1195) <= not(layer2_outputs(4207)) or (layer2_outputs(6272));
    layer3_outputs(1196) <= not(layer2_outputs(590));
    layer3_outputs(1197) <= '0';
    layer3_outputs(1198) <= '1';
    layer3_outputs(1199) <= layer2_outputs(1309);
    layer3_outputs(1200) <= layer2_outputs(5143);
    layer3_outputs(1201) <= not((layer2_outputs(1039)) and (layer2_outputs(650)));
    layer3_outputs(1202) <= (layer2_outputs(3468)) and not (layer2_outputs(4521));
    layer3_outputs(1203) <= not(layer2_outputs(2685));
    layer3_outputs(1204) <= layer2_outputs(4304);
    layer3_outputs(1205) <= not(layer2_outputs(1118));
    layer3_outputs(1206) <= not(layer2_outputs(1491));
    layer3_outputs(1207) <= not(layer2_outputs(2441));
    layer3_outputs(1208) <= not(layer2_outputs(2646));
    layer3_outputs(1209) <= '1';
    layer3_outputs(1210) <= (layer2_outputs(3002)) and (layer2_outputs(5649));
    layer3_outputs(1211) <= '1';
    layer3_outputs(1212) <= layer2_outputs(6326);
    layer3_outputs(1213) <= (layer2_outputs(506)) and (layer2_outputs(385));
    layer3_outputs(1214) <= (layer2_outputs(2834)) or (layer2_outputs(6697));
    layer3_outputs(1215) <= not(layer2_outputs(2278)) or (layer2_outputs(2435));
    layer3_outputs(1216) <= not(layer2_outputs(6387));
    layer3_outputs(1217) <= not(layer2_outputs(3057));
    layer3_outputs(1218) <= not((layer2_outputs(7537)) and (layer2_outputs(4610)));
    layer3_outputs(1219) <= (layer2_outputs(6655)) and not (layer2_outputs(449));
    layer3_outputs(1220) <= not(layer2_outputs(4956)) or (layer2_outputs(4112));
    layer3_outputs(1221) <= '1';
    layer3_outputs(1222) <= (layer2_outputs(2261)) and not (layer2_outputs(6856));
    layer3_outputs(1223) <= not(layer2_outputs(439)) or (layer2_outputs(4574));
    layer3_outputs(1224) <= not(layer2_outputs(1089));
    layer3_outputs(1225) <= '1';
    layer3_outputs(1226) <= layer2_outputs(7261);
    layer3_outputs(1227) <= not(layer2_outputs(1282));
    layer3_outputs(1228) <= not(layer2_outputs(1943)) or (layer2_outputs(3028));
    layer3_outputs(1229) <= (layer2_outputs(262)) or (layer2_outputs(6518));
    layer3_outputs(1230) <= layer2_outputs(2236);
    layer3_outputs(1231) <= not((layer2_outputs(1072)) xor (layer2_outputs(5533)));
    layer3_outputs(1232) <= not((layer2_outputs(213)) or (layer2_outputs(7405)));
    layer3_outputs(1233) <= (layer2_outputs(2727)) and (layer2_outputs(1457));
    layer3_outputs(1234) <= (layer2_outputs(2568)) and not (layer2_outputs(3554));
    layer3_outputs(1235) <= (layer2_outputs(3843)) and not (layer2_outputs(7163));
    layer3_outputs(1236) <= not(layer2_outputs(1864));
    layer3_outputs(1237) <= not(layer2_outputs(825)) or (layer2_outputs(7217));
    layer3_outputs(1238) <= (layer2_outputs(1096)) and (layer2_outputs(4132));
    layer3_outputs(1239) <= '1';
    layer3_outputs(1240) <= (layer2_outputs(2125)) and not (layer2_outputs(759));
    layer3_outputs(1241) <= '0';
    layer3_outputs(1242) <= layer2_outputs(357);
    layer3_outputs(1243) <= not(layer2_outputs(6043));
    layer3_outputs(1244) <= '1';
    layer3_outputs(1245) <= layer2_outputs(6956);
    layer3_outputs(1246) <= not((layer2_outputs(197)) and (layer2_outputs(7210)));
    layer3_outputs(1247) <= not(layer2_outputs(6349));
    layer3_outputs(1248) <= layer2_outputs(5114);
    layer3_outputs(1249) <= (layer2_outputs(7520)) and (layer2_outputs(5471));
    layer3_outputs(1250) <= not(layer2_outputs(397));
    layer3_outputs(1251) <= '1';
    layer3_outputs(1252) <= (layer2_outputs(2601)) and (layer2_outputs(4607));
    layer3_outputs(1253) <= not(layer2_outputs(167)) or (layer2_outputs(2918));
    layer3_outputs(1254) <= (layer2_outputs(5746)) and not (layer2_outputs(121));
    layer3_outputs(1255) <= '1';
    layer3_outputs(1256) <= not((layer2_outputs(6065)) xor (layer2_outputs(3793)));
    layer3_outputs(1257) <= not((layer2_outputs(3950)) or (layer2_outputs(4017)));
    layer3_outputs(1258) <= not(layer2_outputs(5569));
    layer3_outputs(1259) <= not(layer2_outputs(5354)) or (layer2_outputs(4939));
    layer3_outputs(1260) <= layer2_outputs(6346);
    layer3_outputs(1261) <= layer2_outputs(4539);
    layer3_outputs(1262) <= layer2_outputs(1056);
    layer3_outputs(1263) <= not((layer2_outputs(4254)) xor (layer2_outputs(2373)));
    layer3_outputs(1264) <= not((layer2_outputs(1673)) or (layer2_outputs(4583)));
    layer3_outputs(1265) <= layer2_outputs(4900);
    layer3_outputs(1266) <= not(layer2_outputs(6264));
    layer3_outputs(1267) <= not(layer2_outputs(4261)) or (layer2_outputs(5340));
    layer3_outputs(1268) <= not(layer2_outputs(4765)) or (layer2_outputs(395));
    layer3_outputs(1269) <= not((layer2_outputs(3448)) and (layer2_outputs(3748)));
    layer3_outputs(1270) <= not(layer2_outputs(3809));
    layer3_outputs(1271) <= not(layer2_outputs(7440));
    layer3_outputs(1272) <= layer2_outputs(5917);
    layer3_outputs(1273) <= layer2_outputs(3423);
    layer3_outputs(1274) <= layer2_outputs(5827);
    layer3_outputs(1275) <= (layer2_outputs(7651)) and not (layer2_outputs(26));
    layer3_outputs(1276) <= (layer2_outputs(4934)) and not (layer2_outputs(2412));
    layer3_outputs(1277) <= (layer2_outputs(7237)) and not (layer2_outputs(2875));
    layer3_outputs(1278) <= layer2_outputs(4500);
    layer3_outputs(1279) <= (layer2_outputs(1580)) and not (layer2_outputs(5558));
    layer3_outputs(1280) <= not(layer2_outputs(1743));
    layer3_outputs(1281) <= not(layer2_outputs(6892));
    layer3_outputs(1282) <= (layer2_outputs(17)) and (layer2_outputs(5820));
    layer3_outputs(1283) <= layer2_outputs(4573);
    layer3_outputs(1284) <= not(layer2_outputs(5545));
    layer3_outputs(1285) <= not(layer2_outputs(5099));
    layer3_outputs(1286) <= layer2_outputs(6251);
    layer3_outputs(1287) <= (layer2_outputs(5462)) and (layer2_outputs(1045));
    layer3_outputs(1288) <= layer2_outputs(862);
    layer3_outputs(1289) <= (layer2_outputs(7073)) or (layer2_outputs(4327));
    layer3_outputs(1290) <= layer2_outputs(2231);
    layer3_outputs(1291) <= not(layer2_outputs(6962)) or (layer2_outputs(3766));
    layer3_outputs(1292) <= not(layer2_outputs(7188));
    layer3_outputs(1293) <= '0';
    layer3_outputs(1294) <= layer2_outputs(5808);
    layer3_outputs(1295) <= layer2_outputs(1910);
    layer3_outputs(1296) <= not((layer2_outputs(6274)) or (layer2_outputs(1343)));
    layer3_outputs(1297) <= not(layer2_outputs(4915));
    layer3_outputs(1298) <= not((layer2_outputs(3164)) or (layer2_outputs(1080)));
    layer3_outputs(1299) <= not(layer2_outputs(5427)) or (layer2_outputs(2491));
    layer3_outputs(1300) <= not(layer2_outputs(1068)) or (layer2_outputs(5504));
    layer3_outputs(1301) <= not(layer2_outputs(1260)) or (layer2_outputs(1711));
    layer3_outputs(1302) <= not(layer2_outputs(1662));
    layer3_outputs(1303) <= not((layer2_outputs(6568)) xor (layer2_outputs(1151)));
    layer3_outputs(1304) <= (layer2_outputs(3531)) and (layer2_outputs(62));
    layer3_outputs(1305) <= (layer2_outputs(5527)) and not (layer2_outputs(5782));
    layer3_outputs(1306) <= not((layer2_outputs(834)) and (layer2_outputs(291)));
    layer3_outputs(1307) <= not((layer2_outputs(5107)) xor (layer2_outputs(4013)));
    layer3_outputs(1308) <= (layer2_outputs(4562)) or (layer2_outputs(3292));
    layer3_outputs(1309) <= not(layer2_outputs(2688));
    layer3_outputs(1310) <= not((layer2_outputs(7052)) and (layer2_outputs(7303)));
    layer3_outputs(1311) <= layer2_outputs(642);
    layer3_outputs(1312) <= (layer2_outputs(4595)) and not (layer2_outputs(5630));
    layer3_outputs(1313) <= layer2_outputs(6263);
    layer3_outputs(1314) <= layer2_outputs(2560);
    layer3_outputs(1315) <= not(layer2_outputs(6453)) or (layer2_outputs(2026));
    layer3_outputs(1316) <= '1';
    layer3_outputs(1317) <= layer2_outputs(1193);
    layer3_outputs(1318) <= layer2_outputs(6671);
    layer3_outputs(1319) <= (layer2_outputs(5118)) and (layer2_outputs(5811));
    layer3_outputs(1320) <= not(layer2_outputs(5426)) or (layer2_outputs(1356));
    layer3_outputs(1321) <= not((layer2_outputs(6072)) and (layer2_outputs(52)));
    layer3_outputs(1322) <= not(layer2_outputs(6345));
    layer3_outputs(1323) <= '1';
    layer3_outputs(1324) <= not(layer2_outputs(2536)) or (layer2_outputs(866));
    layer3_outputs(1325) <= '1';
    layer3_outputs(1326) <= (layer2_outputs(4636)) and not (layer2_outputs(6819));
    layer3_outputs(1327) <= not((layer2_outputs(2187)) or (layer2_outputs(3207)));
    layer3_outputs(1328) <= (layer2_outputs(433)) and not (layer2_outputs(362));
    layer3_outputs(1329) <= (layer2_outputs(6391)) or (layer2_outputs(2323));
    layer3_outputs(1330) <= not(layer2_outputs(1435));
    layer3_outputs(1331) <= not((layer2_outputs(7194)) xor (layer2_outputs(3277)));
    layer3_outputs(1332) <= not(layer2_outputs(769));
    layer3_outputs(1333) <= '0';
    layer3_outputs(1334) <= not(layer2_outputs(4124)) or (layer2_outputs(6187));
    layer3_outputs(1335) <= (layer2_outputs(5062)) and (layer2_outputs(926));
    layer3_outputs(1336) <= layer2_outputs(51);
    layer3_outputs(1337) <= not(layer2_outputs(4342));
    layer3_outputs(1338) <= layer2_outputs(1683);
    layer3_outputs(1339) <= not(layer2_outputs(6070));
    layer3_outputs(1340) <= '0';
    layer3_outputs(1341) <= not(layer2_outputs(2644)) or (layer2_outputs(56));
    layer3_outputs(1342) <= layer2_outputs(4480);
    layer3_outputs(1343) <= not(layer2_outputs(3093)) or (layer2_outputs(2349));
    layer3_outputs(1344) <= (layer2_outputs(4136)) and not (layer2_outputs(3469));
    layer3_outputs(1345) <= layer2_outputs(3371);
    layer3_outputs(1346) <= (layer2_outputs(6129)) and not (layer2_outputs(7072));
    layer3_outputs(1347) <= (layer2_outputs(993)) and not (layer2_outputs(4765));
    layer3_outputs(1348) <= (layer2_outputs(1762)) and not (layer2_outputs(4832));
    layer3_outputs(1349) <= '0';
    layer3_outputs(1350) <= (layer2_outputs(3062)) xor (layer2_outputs(2424));
    layer3_outputs(1351) <= not(layer2_outputs(3061)) or (layer2_outputs(1732));
    layer3_outputs(1352) <= layer2_outputs(416);
    layer3_outputs(1353) <= not(layer2_outputs(2890));
    layer3_outputs(1354) <= not(layer2_outputs(5048)) or (layer2_outputs(7286));
    layer3_outputs(1355) <= layer2_outputs(129);
    layer3_outputs(1356) <= '0';
    layer3_outputs(1357) <= not(layer2_outputs(6948));
    layer3_outputs(1358) <= not(layer2_outputs(4614)) or (layer2_outputs(3824));
    layer3_outputs(1359) <= not(layer2_outputs(6021)) or (layer2_outputs(3150));
    layer3_outputs(1360) <= not(layer2_outputs(6234));
    layer3_outputs(1361) <= '1';
    layer3_outputs(1362) <= (layer2_outputs(5434)) or (layer2_outputs(4388));
    layer3_outputs(1363) <= '1';
    layer3_outputs(1364) <= not(layer2_outputs(5306));
    layer3_outputs(1365) <= not(layer2_outputs(7533));
    layer3_outputs(1366) <= (layer2_outputs(6661)) and not (layer2_outputs(3850));
    layer3_outputs(1367) <= '1';
    layer3_outputs(1368) <= (layer2_outputs(2814)) or (layer2_outputs(4612));
    layer3_outputs(1369) <= '0';
    layer3_outputs(1370) <= (layer2_outputs(7083)) and not (layer2_outputs(6997));
    layer3_outputs(1371) <= (layer2_outputs(6950)) or (layer2_outputs(1061));
    layer3_outputs(1372) <= not((layer2_outputs(2697)) or (layer2_outputs(6601)));
    layer3_outputs(1373) <= '0';
    layer3_outputs(1374) <= (layer2_outputs(4813)) and (layer2_outputs(4141));
    layer3_outputs(1375) <= layer2_outputs(3277);
    layer3_outputs(1376) <= '1';
    layer3_outputs(1377) <= not((layer2_outputs(6886)) and (layer2_outputs(4350)));
    layer3_outputs(1378) <= not((layer2_outputs(6092)) or (layer2_outputs(5253)));
    layer3_outputs(1379) <= (layer2_outputs(465)) and not (layer2_outputs(7396));
    layer3_outputs(1380) <= '1';
    layer3_outputs(1381) <= layer2_outputs(6655);
    layer3_outputs(1382) <= not((layer2_outputs(4704)) and (layer2_outputs(5721)));
    layer3_outputs(1383) <= layer2_outputs(2230);
    layer3_outputs(1384) <= not((layer2_outputs(756)) and (layer2_outputs(4693)));
    layer3_outputs(1385) <= '1';
    layer3_outputs(1386) <= not((layer2_outputs(6279)) or (layer2_outputs(201)));
    layer3_outputs(1387) <= layer2_outputs(3638);
    layer3_outputs(1388) <= (layer2_outputs(2862)) and not (layer2_outputs(1498));
    layer3_outputs(1389) <= (layer2_outputs(6157)) xor (layer2_outputs(5020));
    layer3_outputs(1390) <= layer2_outputs(356);
    layer3_outputs(1391) <= not(layer2_outputs(125)) or (layer2_outputs(524));
    layer3_outputs(1392) <= not(layer2_outputs(2169));
    layer3_outputs(1393) <= '1';
    layer3_outputs(1394) <= (layer2_outputs(5983)) and not (layer2_outputs(3517));
    layer3_outputs(1395) <= layer2_outputs(1465);
    layer3_outputs(1396) <= '0';
    layer3_outputs(1397) <= (layer2_outputs(3355)) and not (layer2_outputs(5386));
    layer3_outputs(1398) <= not(layer2_outputs(5071)) or (layer2_outputs(2283));
    layer3_outputs(1399) <= layer2_outputs(5238);
    layer3_outputs(1400) <= (layer2_outputs(7197)) and (layer2_outputs(1937));
    layer3_outputs(1401) <= not(layer2_outputs(5621)) or (layer2_outputs(375));
    layer3_outputs(1402) <= not(layer2_outputs(7568));
    layer3_outputs(1403) <= layer2_outputs(6720);
    layer3_outputs(1404) <= (layer2_outputs(4933)) and (layer2_outputs(1834));
    layer3_outputs(1405) <= (layer2_outputs(5968)) and (layer2_outputs(2194));
    layer3_outputs(1406) <= layer2_outputs(2388);
    layer3_outputs(1407) <= not((layer2_outputs(6659)) or (layer2_outputs(1453)));
    layer3_outputs(1408) <= (layer2_outputs(870)) and (layer2_outputs(2442));
    layer3_outputs(1409) <= (layer2_outputs(4908)) or (layer2_outputs(4891));
    layer3_outputs(1410) <= (layer2_outputs(1293)) and (layer2_outputs(4135));
    layer3_outputs(1411) <= not(layer2_outputs(4466));
    layer3_outputs(1412) <= layer2_outputs(2109);
    layer3_outputs(1413) <= (layer2_outputs(4000)) and (layer2_outputs(5064));
    layer3_outputs(1414) <= layer2_outputs(5472);
    layer3_outputs(1415) <= layer2_outputs(5900);
    layer3_outputs(1416) <= layer2_outputs(6891);
    layer3_outputs(1417) <= not((layer2_outputs(132)) or (layer2_outputs(4946)));
    layer3_outputs(1418) <= (layer2_outputs(3627)) and not (layer2_outputs(4233));
    layer3_outputs(1419) <= not(layer2_outputs(2936));
    layer3_outputs(1420) <= not((layer2_outputs(6824)) xor (layer2_outputs(3145)));
    layer3_outputs(1421) <= (layer2_outputs(3327)) and not (layer2_outputs(291));
    layer3_outputs(1422) <= not((layer2_outputs(3969)) and (layer2_outputs(457)));
    layer3_outputs(1423) <= not(layer2_outputs(5440)) or (layer2_outputs(812));
    layer3_outputs(1424) <= not(layer2_outputs(1069));
    layer3_outputs(1425) <= (layer2_outputs(536)) and not (layer2_outputs(7089));
    layer3_outputs(1426) <= layer2_outputs(4009);
    layer3_outputs(1427) <= not(layer2_outputs(6033)) or (layer2_outputs(5795));
    layer3_outputs(1428) <= not(layer2_outputs(28));
    layer3_outputs(1429) <= not(layer2_outputs(6594)) or (layer2_outputs(4846));
    layer3_outputs(1430) <= (layer2_outputs(7591)) and not (layer2_outputs(3670));
    layer3_outputs(1431) <= not(layer2_outputs(5698));
    layer3_outputs(1432) <= '1';
    layer3_outputs(1433) <= (layer2_outputs(5432)) and (layer2_outputs(3543));
    layer3_outputs(1434) <= '1';
    layer3_outputs(1435) <= (layer2_outputs(2083)) and (layer2_outputs(872));
    layer3_outputs(1436) <= layer2_outputs(7338);
    layer3_outputs(1437) <= not(layer2_outputs(5131));
    layer3_outputs(1438) <= not((layer2_outputs(3709)) or (layer2_outputs(6674)));
    layer3_outputs(1439) <= (layer2_outputs(3514)) and not (layer2_outputs(1901));
    layer3_outputs(1440) <= layer2_outputs(7380);
    layer3_outputs(1441) <= (layer2_outputs(772)) and not (layer2_outputs(1104));
    layer3_outputs(1442) <= not(layer2_outputs(823));
    layer3_outputs(1443) <= '1';
    layer3_outputs(1444) <= not((layer2_outputs(7010)) or (layer2_outputs(5700)));
    layer3_outputs(1445) <= layer2_outputs(4143);
    layer3_outputs(1446) <= not(layer2_outputs(6656));
    layer3_outputs(1447) <= '0';
    layer3_outputs(1448) <= not((layer2_outputs(6750)) and (layer2_outputs(3320)));
    layer3_outputs(1449) <= '1';
    layer3_outputs(1450) <= '0';
    layer3_outputs(1451) <= layer2_outputs(6172);
    layer3_outputs(1452) <= (layer2_outputs(352)) or (layer2_outputs(7201));
    layer3_outputs(1453) <= not(layer2_outputs(1312));
    layer3_outputs(1454) <= not((layer2_outputs(6317)) or (layer2_outputs(6708)));
    layer3_outputs(1455) <= not(layer2_outputs(340));
    layer3_outputs(1456) <= layer2_outputs(4373);
    layer3_outputs(1457) <= layer2_outputs(1817);
    layer3_outputs(1458) <= (layer2_outputs(5243)) and not (layer2_outputs(1503));
    layer3_outputs(1459) <= layer2_outputs(2807);
    layer3_outputs(1460) <= layer2_outputs(1826);
    layer3_outputs(1461) <= not(layer2_outputs(4197));
    layer3_outputs(1462) <= not((layer2_outputs(3079)) or (layer2_outputs(3555)));
    layer3_outputs(1463) <= not(layer2_outputs(2419)) or (layer2_outputs(7590));
    layer3_outputs(1464) <= not(layer2_outputs(6375)) or (layer2_outputs(5658));
    layer3_outputs(1465) <= not(layer2_outputs(816)) or (layer2_outputs(1730));
    layer3_outputs(1466) <= (layer2_outputs(5580)) and not (layer2_outputs(7133));
    layer3_outputs(1467) <= layer2_outputs(4740);
    layer3_outputs(1468) <= layer2_outputs(2637);
    layer3_outputs(1469) <= (layer2_outputs(7426)) and not (layer2_outputs(4693));
    layer3_outputs(1470) <= layer2_outputs(5984);
    layer3_outputs(1471) <= (layer2_outputs(4185)) and not (layer2_outputs(5930));
    layer3_outputs(1472) <= layer2_outputs(366);
    layer3_outputs(1473) <= not(layer2_outputs(6034));
    layer3_outputs(1474) <= not((layer2_outputs(6880)) or (layer2_outputs(5860)));
    layer3_outputs(1475) <= not(layer2_outputs(673)) or (layer2_outputs(7204));
    layer3_outputs(1476) <= not(layer2_outputs(4493));
    layer3_outputs(1477) <= not(layer2_outputs(2317));
    layer3_outputs(1478) <= not(layer2_outputs(1641));
    layer3_outputs(1479) <= not((layer2_outputs(840)) or (layer2_outputs(1685)));
    layer3_outputs(1480) <= (layer2_outputs(6733)) or (layer2_outputs(5810));
    layer3_outputs(1481) <= not(layer2_outputs(6998));
    layer3_outputs(1482) <= not((layer2_outputs(5971)) or (layer2_outputs(7447)));
    layer3_outputs(1483) <= layer2_outputs(3959);
    layer3_outputs(1484) <= (layer2_outputs(4315)) and (layer2_outputs(7114));
    layer3_outputs(1485) <= not((layer2_outputs(4672)) xor (layer2_outputs(6629)));
    layer3_outputs(1486) <= '1';
    layer3_outputs(1487) <= layer2_outputs(5862);
    layer3_outputs(1488) <= not((layer2_outputs(3024)) and (layer2_outputs(5912)));
    layer3_outputs(1489) <= (layer2_outputs(3749)) and not (layer2_outputs(948));
    layer3_outputs(1490) <= (layer2_outputs(4401)) and not (layer2_outputs(7503));
    layer3_outputs(1491) <= layer2_outputs(4886);
    layer3_outputs(1492) <= layer2_outputs(6956);
    layer3_outputs(1493) <= not(layer2_outputs(3864)) or (layer2_outputs(594));
    layer3_outputs(1494) <= layer2_outputs(563);
    layer3_outputs(1495) <= (layer2_outputs(763)) and (layer2_outputs(4806));
    layer3_outputs(1496) <= layer2_outputs(4754);
    layer3_outputs(1497) <= (layer2_outputs(1487)) and not (layer2_outputs(3751));
    layer3_outputs(1498) <= not(layer2_outputs(1428)) or (layer2_outputs(778));
    layer3_outputs(1499) <= layer2_outputs(1861);
    layer3_outputs(1500) <= (layer2_outputs(4218)) and not (layer2_outputs(5636));
    layer3_outputs(1501) <= (layer2_outputs(6436)) and not (layer2_outputs(3756));
    layer3_outputs(1502) <= (layer2_outputs(742)) and not (layer2_outputs(5320));
    layer3_outputs(1503) <= not((layer2_outputs(5988)) or (layer2_outputs(3181)));
    layer3_outputs(1504) <= layer2_outputs(5386);
    layer3_outputs(1505) <= not(layer2_outputs(836));
    layer3_outputs(1506) <= '0';
    layer3_outputs(1507) <= not((layer2_outputs(3828)) or (layer2_outputs(2985)));
    layer3_outputs(1508) <= layer2_outputs(4242);
    layer3_outputs(1509) <= (layer2_outputs(984)) and not (layer2_outputs(4801));
    layer3_outputs(1510) <= not(layer2_outputs(6321));
    layer3_outputs(1511) <= not(layer2_outputs(3549));
    layer3_outputs(1512) <= layer2_outputs(552);
    layer3_outputs(1513) <= not(layer2_outputs(6894)) or (layer2_outputs(1725));
    layer3_outputs(1514) <= layer2_outputs(5529);
    layer3_outputs(1515) <= not((layer2_outputs(6480)) or (layer2_outputs(7222)));
    layer3_outputs(1516) <= '1';
    layer3_outputs(1517) <= not(layer2_outputs(6161)) or (layer2_outputs(4259));
    layer3_outputs(1518) <= layer2_outputs(182);
    layer3_outputs(1519) <= (layer2_outputs(804)) and not (layer2_outputs(7620));
    layer3_outputs(1520) <= not(layer2_outputs(7679));
    layer3_outputs(1521) <= not(layer2_outputs(4275));
    layer3_outputs(1522) <= not(layer2_outputs(3124)) or (layer2_outputs(5745));
    layer3_outputs(1523) <= layer2_outputs(26);
    layer3_outputs(1524) <= not(layer2_outputs(5244));
    layer3_outputs(1525) <= not(layer2_outputs(3443));
    layer3_outputs(1526) <= not((layer2_outputs(5222)) and (layer2_outputs(3242)));
    layer3_outputs(1527) <= not(layer2_outputs(7473));
    layer3_outputs(1528) <= layer2_outputs(239);
    layer3_outputs(1529) <= (layer2_outputs(4008)) and (layer2_outputs(732));
    layer3_outputs(1530) <= not(layer2_outputs(2995));
    layer3_outputs(1531) <= '0';
    layer3_outputs(1532) <= layer2_outputs(7280);
    layer3_outputs(1533) <= '1';
    layer3_outputs(1534) <= '1';
    layer3_outputs(1535) <= (layer2_outputs(1978)) xor (layer2_outputs(648));
    layer3_outputs(1536) <= (layer2_outputs(5391)) and not (layer2_outputs(1863));
    layer3_outputs(1537) <= not(layer2_outputs(3849)) or (layer2_outputs(4397));
    layer3_outputs(1538) <= not(layer2_outputs(2840));
    layer3_outputs(1539) <= not((layer2_outputs(4346)) or (layer2_outputs(5403)));
    layer3_outputs(1540) <= (layer2_outputs(3604)) and not (layer2_outputs(7468));
    layer3_outputs(1541) <= '1';
    layer3_outputs(1542) <= '1';
    layer3_outputs(1543) <= not((layer2_outputs(6286)) xor (layer2_outputs(1721)));
    layer3_outputs(1544) <= layer2_outputs(3579);
    layer3_outputs(1545) <= not(layer2_outputs(310)) or (layer2_outputs(2400));
    layer3_outputs(1546) <= (layer2_outputs(6807)) and not (layer2_outputs(6613));
    layer3_outputs(1547) <= not(layer2_outputs(153));
    layer3_outputs(1548) <= '1';
    layer3_outputs(1549) <= not(layer2_outputs(5111)) or (layer2_outputs(501));
    layer3_outputs(1550) <= (layer2_outputs(4517)) and not (layer2_outputs(4481));
    layer3_outputs(1551) <= layer2_outputs(219);
    layer3_outputs(1552) <= not(layer2_outputs(2573)) or (layer2_outputs(5096));
    layer3_outputs(1553) <= layer2_outputs(2396);
    layer3_outputs(1554) <= not((layer2_outputs(6431)) and (layer2_outputs(4563)));
    layer3_outputs(1555) <= (layer2_outputs(1840)) and not (layer2_outputs(4231));
    layer3_outputs(1556) <= '1';
    layer3_outputs(1557) <= '1';
    layer3_outputs(1558) <= (layer2_outputs(3016)) or (layer2_outputs(5749));
    layer3_outputs(1559) <= (layer2_outputs(3626)) and not (layer2_outputs(1251));
    layer3_outputs(1560) <= not(layer2_outputs(6988));
    layer3_outputs(1561) <= not(layer2_outputs(405));
    layer3_outputs(1562) <= '0';
    layer3_outputs(1563) <= '0';
    layer3_outputs(1564) <= not((layer2_outputs(6134)) or (layer2_outputs(3471)));
    layer3_outputs(1565) <= (layer2_outputs(764)) xor (layer2_outputs(5072));
    layer3_outputs(1566) <= (layer2_outputs(7487)) or (layer2_outputs(3731));
    layer3_outputs(1567) <= (layer2_outputs(2677)) and not (layer2_outputs(5890));
    layer3_outputs(1568) <= (layer2_outputs(213)) and not (layer2_outputs(7116));
    layer3_outputs(1569) <= not(layer2_outputs(57));
    layer3_outputs(1570) <= '0';
    layer3_outputs(1571) <= not(layer2_outputs(2742)) or (layer2_outputs(5105));
    layer3_outputs(1572) <= layer2_outputs(6267);
    layer3_outputs(1573) <= not(layer2_outputs(6395));
    layer3_outputs(1574) <= layer2_outputs(6390);
    layer3_outputs(1575) <= layer2_outputs(3152);
    layer3_outputs(1576) <= (layer2_outputs(1154)) and not (layer2_outputs(7527));
    layer3_outputs(1577) <= not(layer2_outputs(1095));
    layer3_outputs(1578) <= not(layer2_outputs(4795)) or (layer2_outputs(4925));
    layer3_outputs(1579) <= not(layer2_outputs(5287));
    layer3_outputs(1580) <= (layer2_outputs(1234)) or (layer2_outputs(5275));
    layer3_outputs(1581) <= layer2_outputs(2563);
    layer3_outputs(1582) <= (layer2_outputs(2942)) and (layer2_outputs(4274));
    layer3_outputs(1583) <= (layer2_outputs(1117)) or (layer2_outputs(163));
    layer3_outputs(1584) <= not(layer2_outputs(3817));
    layer3_outputs(1585) <= not(layer2_outputs(7420)) or (layer2_outputs(7047));
    layer3_outputs(1586) <= (layer2_outputs(6799)) and not (layer2_outputs(6179));
    layer3_outputs(1587) <= not(layer2_outputs(983));
    layer3_outputs(1588) <= layer2_outputs(11);
    layer3_outputs(1589) <= not(layer2_outputs(3018));
    layer3_outputs(1590) <= not(layer2_outputs(5365)) or (layer2_outputs(2430));
    layer3_outputs(1591) <= (layer2_outputs(5373)) or (layer2_outputs(7564));
    layer3_outputs(1592) <= not(layer2_outputs(517)) or (layer2_outputs(679));
    layer3_outputs(1593) <= '1';
    layer3_outputs(1594) <= layer2_outputs(2319);
    layer3_outputs(1595) <= layer2_outputs(715);
    layer3_outputs(1596) <= not(layer2_outputs(1501));
    layer3_outputs(1597) <= (layer2_outputs(7097)) and not (layer2_outputs(1326));
    layer3_outputs(1598) <= '0';
    layer3_outputs(1599) <= (layer2_outputs(7297)) and not (layer2_outputs(5736));
    layer3_outputs(1600) <= '1';
    layer3_outputs(1601) <= not(layer2_outputs(2838)) or (layer2_outputs(504));
    layer3_outputs(1602) <= not((layer2_outputs(4582)) or (layer2_outputs(892)));
    layer3_outputs(1603) <= layer2_outputs(3905);
    layer3_outputs(1604) <= layer2_outputs(5975);
    layer3_outputs(1605) <= (layer2_outputs(3305)) and (layer2_outputs(2242));
    layer3_outputs(1606) <= (layer2_outputs(6748)) and not (layer2_outputs(1548));
    layer3_outputs(1607) <= not(layer2_outputs(1030));
    layer3_outputs(1608) <= (layer2_outputs(1737)) or (layer2_outputs(2873));
    layer3_outputs(1609) <= (layer2_outputs(6188)) and not (layer2_outputs(1716));
    layer3_outputs(1610) <= not(layer2_outputs(47));
    layer3_outputs(1611) <= '1';
    layer3_outputs(1612) <= layer2_outputs(3512);
    layer3_outputs(1613) <= (layer2_outputs(529)) or (layer2_outputs(5823));
    layer3_outputs(1614) <= not(layer2_outputs(6658));
    layer3_outputs(1615) <= not(layer2_outputs(2453)) or (layer2_outputs(707));
    layer3_outputs(1616) <= not(layer2_outputs(2));
    layer3_outputs(1617) <= layer2_outputs(6316);
    layer3_outputs(1618) <= layer2_outputs(2673);
    layer3_outputs(1619) <= not((layer2_outputs(5758)) or (layer2_outputs(7328)));
    layer3_outputs(1620) <= (layer2_outputs(1589)) or (layer2_outputs(263));
    layer3_outputs(1621) <= (layer2_outputs(4416)) xor (layer2_outputs(5575));
    layer3_outputs(1622) <= not(layer2_outputs(5701)) or (layer2_outputs(5551));
    layer3_outputs(1623) <= (layer2_outputs(3578)) and (layer2_outputs(2260));
    layer3_outputs(1624) <= (layer2_outputs(7093)) and not (layer2_outputs(7472));
    layer3_outputs(1625) <= (layer2_outputs(788)) and (layer2_outputs(2471));
    layer3_outputs(1626) <= (layer2_outputs(6374)) and not (layer2_outputs(5399));
    layer3_outputs(1627) <= not(layer2_outputs(5939)) or (layer2_outputs(2085));
    layer3_outputs(1628) <= not(layer2_outputs(4159));
    layer3_outputs(1629) <= (layer2_outputs(1521)) or (layer2_outputs(7071));
    layer3_outputs(1630) <= not(layer2_outputs(549));
    layer3_outputs(1631) <= not(layer2_outputs(14));
    layer3_outputs(1632) <= layer2_outputs(6606);
    layer3_outputs(1633) <= not((layer2_outputs(974)) and (layer2_outputs(6277)));
    layer3_outputs(1634) <= layer2_outputs(3084);
    layer3_outputs(1635) <= (layer2_outputs(2522)) or (layer2_outputs(1843));
    layer3_outputs(1636) <= '1';
    layer3_outputs(1637) <= layer2_outputs(3458);
    layer3_outputs(1638) <= not(layer2_outputs(410));
    layer3_outputs(1639) <= (layer2_outputs(6754)) or (layer2_outputs(1633));
    layer3_outputs(1640) <= not((layer2_outputs(554)) and (layer2_outputs(3998)));
    layer3_outputs(1641) <= layer2_outputs(3335);
    layer3_outputs(1642) <= not(layer2_outputs(6453));
    layer3_outputs(1643) <= not(layer2_outputs(6334));
    layer3_outputs(1644) <= not((layer2_outputs(7170)) or (layer2_outputs(7159)));
    layer3_outputs(1645) <= (layer2_outputs(22)) xor (layer2_outputs(3364));
    layer3_outputs(1646) <= not(layer2_outputs(6027));
    layer3_outputs(1647) <= layer2_outputs(5641);
    layer3_outputs(1648) <= (layer2_outputs(6477)) or (layer2_outputs(4815));
    layer3_outputs(1649) <= (layer2_outputs(2669)) xor (layer2_outputs(3473));
    layer3_outputs(1650) <= not(layer2_outputs(3736));
    layer3_outputs(1651) <= (layer2_outputs(7397)) or (layer2_outputs(5732));
    layer3_outputs(1652) <= (layer2_outputs(2993)) and not (layer2_outputs(3165));
    layer3_outputs(1653) <= not((layer2_outputs(2468)) and (layer2_outputs(7624)));
    layer3_outputs(1654) <= not((layer2_outputs(2629)) and (layer2_outputs(3201)));
    layer3_outputs(1655) <= not(layer2_outputs(1700));
    layer3_outputs(1656) <= (layer2_outputs(2768)) or (layer2_outputs(3252));
    layer3_outputs(1657) <= layer2_outputs(6196);
    layer3_outputs(1658) <= not(layer2_outputs(190)) or (layer2_outputs(3060));
    layer3_outputs(1659) <= '1';
    layer3_outputs(1660) <= not(layer2_outputs(1912)) or (layer2_outputs(2299));
    layer3_outputs(1661) <= (layer2_outputs(2310)) xor (layer2_outputs(5668));
    layer3_outputs(1662) <= (layer2_outputs(7452)) and not (layer2_outputs(6647));
    layer3_outputs(1663) <= (layer2_outputs(414)) or (layer2_outputs(514));
    layer3_outputs(1664) <= (layer2_outputs(4788)) and not (layer2_outputs(3717));
    layer3_outputs(1665) <= layer2_outputs(6012);
    layer3_outputs(1666) <= not(layer2_outputs(6034));
    layer3_outputs(1667) <= layer2_outputs(4465);
    layer3_outputs(1668) <= layer2_outputs(7183);
    layer3_outputs(1669) <= layer2_outputs(372);
    layer3_outputs(1670) <= '0';
    layer3_outputs(1671) <= not(layer2_outputs(1475));
    layer3_outputs(1672) <= not((layer2_outputs(4608)) xor (layer2_outputs(6642)));
    layer3_outputs(1673) <= (layer2_outputs(5293)) or (layer2_outputs(3704));
    layer3_outputs(1674) <= '1';
    layer3_outputs(1675) <= (layer2_outputs(6282)) or (layer2_outputs(758));
    layer3_outputs(1676) <= not((layer2_outputs(7074)) or (layer2_outputs(1803)));
    layer3_outputs(1677) <= (layer2_outputs(1685)) and not (layer2_outputs(7547));
    layer3_outputs(1678) <= not(layer2_outputs(2347));
    layer3_outputs(1679) <= layer2_outputs(3489);
    layer3_outputs(1680) <= '0';
    layer3_outputs(1681) <= not((layer2_outputs(236)) or (layer2_outputs(2395)));
    layer3_outputs(1682) <= '0';
    layer3_outputs(1683) <= not(layer2_outputs(2614)) or (layer2_outputs(6276));
    layer3_outputs(1684) <= not(layer2_outputs(3962));
    layer3_outputs(1685) <= '1';
    layer3_outputs(1686) <= not((layer2_outputs(6226)) xor (layer2_outputs(1256)));
    layer3_outputs(1687) <= not(layer2_outputs(4870));
    layer3_outputs(1688) <= not((layer2_outputs(6702)) or (layer2_outputs(319)));
    layer3_outputs(1689) <= not((layer2_outputs(5350)) or (layer2_outputs(1959)));
    layer3_outputs(1690) <= not((layer2_outputs(1295)) and (layer2_outputs(7599)));
    layer3_outputs(1691) <= (layer2_outputs(7636)) or (layer2_outputs(5084));
    layer3_outputs(1692) <= layer2_outputs(2893);
    layer3_outputs(1693) <= not((layer2_outputs(5)) or (layer2_outputs(1965)));
    layer3_outputs(1694) <= (layer2_outputs(5430)) xor (layer2_outputs(5836));
    layer3_outputs(1695) <= (layer2_outputs(4119)) and not (layer2_outputs(789));
    layer3_outputs(1696) <= not(layer2_outputs(339));
    layer3_outputs(1697) <= not(layer2_outputs(5619)) or (layer2_outputs(602));
    layer3_outputs(1698) <= layer2_outputs(1523);
    layer3_outputs(1699) <= not(layer2_outputs(1107));
    layer3_outputs(1700) <= (layer2_outputs(2593)) and (layer2_outputs(4818));
    layer3_outputs(1701) <= layer2_outputs(7494);
    layer3_outputs(1702) <= not((layer2_outputs(5123)) or (layer2_outputs(5099)));
    layer3_outputs(1703) <= not(layer2_outputs(4974)) or (layer2_outputs(755));
    layer3_outputs(1704) <= '1';
    layer3_outputs(1705) <= layer2_outputs(5574);
    layer3_outputs(1706) <= (layer2_outputs(637)) and (layer2_outputs(734));
    layer3_outputs(1707) <= (layer2_outputs(3657)) or (layer2_outputs(3434));
    layer3_outputs(1708) <= '0';
    layer3_outputs(1709) <= layer2_outputs(3908);
    layer3_outputs(1710) <= not(layer2_outputs(4146));
    layer3_outputs(1711) <= (layer2_outputs(7528)) and (layer2_outputs(5687));
    layer3_outputs(1712) <= '1';
    layer3_outputs(1713) <= layer2_outputs(4611);
    layer3_outputs(1714) <= (layer2_outputs(5178)) and (layer2_outputs(3899));
    layer3_outputs(1715) <= not(layer2_outputs(686));
    layer3_outputs(1716) <= not(layer2_outputs(6539)) or (layer2_outputs(6700));
    layer3_outputs(1717) <= not(layer2_outputs(7521));
    layer3_outputs(1718) <= not((layer2_outputs(1147)) or (layer2_outputs(1615)));
    layer3_outputs(1719) <= (layer2_outputs(6404)) and not (layer2_outputs(3550));
    layer3_outputs(1720) <= not(layer2_outputs(2713));
    layer3_outputs(1721) <= not(layer2_outputs(755));
    layer3_outputs(1722) <= not((layer2_outputs(3977)) xor (layer2_outputs(4590)));
    layer3_outputs(1723) <= layer2_outputs(74);
    layer3_outputs(1724) <= not(layer2_outputs(1603)) or (layer2_outputs(687));
    layer3_outputs(1725) <= (layer2_outputs(2721)) and (layer2_outputs(6614));
    layer3_outputs(1726) <= not(layer2_outputs(1904)) or (layer2_outputs(4767));
    layer3_outputs(1727) <= '0';
    layer3_outputs(1728) <= (layer2_outputs(7195)) and not (layer2_outputs(3554));
    layer3_outputs(1729) <= not(layer2_outputs(1170)) or (layer2_outputs(1746));
    layer3_outputs(1730) <= not((layer2_outputs(2350)) xor (layer2_outputs(6925)));
    layer3_outputs(1731) <= not(layer2_outputs(4440)) or (layer2_outputs(4549));
    layer3_outputs(1732) <= (layer2_outputs(2249)) or (layer2_outputs(1503));
    layer3_outputs(1733) <= layer2_outputs(851);
    layer3_outputs(1734) <= '1';
    layer3_outputs(1735) <= not(layer2_outputs(2437));
    layer3_outputs(1736) <= not(layer2_outputs(2290));
    layer3_outputs(1737) <= not((layer2_outputs(7395)) or (layer2_outputs(1622)));
    layer3_outputs(1738) <= '1';
    layer3_outputs(1739) <= layer2_outputs(6988);
    layer3_outputs(1740) <= not(layer2_outputs(4913)) or (layer2_outputs(4446));
    layer3_outputs(1741) <= '1';
    layer3_outputs(1742) <= layer2_outputs(5878);
    layer3_outputs(1743) <= not((layer2_outputs(38)) xor (layer2_outputs(6127)));
    layer3_outputs(1744) <= not(layer2_outputs(5773));
    layer3_outputs(1745) <= not(layer2_outputs(3928)) or (layer2_outputs(3498));
    layer3_outputs(1746) <= (layer2_outputs(4829)) or (layer2_outputs(3249));
    layer3_outputs(1747) <= (layer2_outputs(7068)) or (layer2_outputs(7163));
    layer3_outputs(1748) <= not(layer2_outputs(1280)) or (layer2_outputs(5936));
    layer3_outputs(1749) <= not(layer2_outputs(7259)) or (layer2_outputs(4679));
    layer3_outputs(1750) <= (layer2_outputs(1254)) and not (layer2_outputs(4315));
    layer3_outputs(1751) <= (layer2_outputs(2904)) or (layer2_outputs(5568));
    layer3_outputs(1752) <= not(layer2_outputs(3588));
    layer3_outputs(1753) <= not((layer2_outputs(6192)) and (layer2_outputs(7560)));
    layer3_outputs(1754) <= not(layer2_outputs(791));
    layer3_outputs(1755) <= not((layer2_outputs(7193)) and (layer2_outputs(406)));
    layer3_outputs(1756) <= not((layer2_outputs(3827)) xor (layer2_outputs(4868)));
    layer3_outputs(1757) <= not(layer2_outputs(1175));
    layer3_outputs(1758) <= (layer2_outputs(5824)) and not (layer2_outputs(5532));
    layer3_outputs(1759) <= not((layer2_outputs(370)) or (layer2_outputs(6080)));
    layer3_outputs(1760) <= not(layer2_outputs(1531)) or (layer2_outputs(5036));
    layer3_outputs(1761) <= not((layer2_outputs(1796)) or (layer2_outputs(5569)));
    layer3_outputs(1762) <= not(layer2_outputs(6590)) or (layer2_outputs(3513));
    layer3_outputs(1763) <= layer2_outputs(443);
    layer3_outputs(1764) <= not(layer2_outputs(312)) or (layer2_outputs(7444));
    layer3_outputs(1765) <= (layer2_outputs(4502)) and (layer2_outputs(3722));
    layer3_outputs(1766) <= not((layer2_outputs(2946)) and (layer2_outputs(5644)));
    layer3_outputs(1767) <= layer2_outputs(5614);
    layer3_outputs(1768) <= not(layer2_outputs(5073)) or (layer2_outputs(731));
    layer3_outputs(1769) <= layer2_outputs(3007);
    layer3_outputs(1770) <= '0';
    layer3_outputs(1771) <= not(layer2_outputs(4036)) or (layer2_outputs(4932));
    layer3_outputs(1772) <= (layer2_outputs(7056)) or (layer2_outputs(7631));
    layer3_outputs(1773) <= not((layer2_outputs(3368)) or (layer2_outputs(2756)));
    layer3_outputs(1774) <= '0';
    layer3_outputs(1775) <= layer2_outputs(2841);
    layer3_outputs(1776) <= not(layer2_outputs(2631)) or (layer2_outputs(2223));
    layer3_outputs(1777) <= (layer2_outputs(7277)) or (layer2_outputs(1483));
    layer3_outputs(1778) <= '0';
    layer3_outputs(1779) <= not(layer2_outputs(7128)) or (layer2_outputs(4513));
    layer3_outputs(1780) <= layer2_outputs(590);
    layer3_outputs(1781) <= not(layer2_outputs(2025));
    layer3_outputs(1782) <= layer2_outputs(5396);
    layer3_outputs(1783) <= (layer2_outputs(824)) or (layer2_outputs(1845));
    layer3_outputs(1784) <= '0';
    layer3_outputs(1785) <= not((layer2_outputs(3011)) or (layer2_outputs(307)));
    layer3_outputs(1786) <= not(layer2_outputs(7099));
    layer3_outputs(1787) <= not(layer2_outputs(1671)) or (layer2_outputs(2905));
    layer3_outputs(1788) <= layer2_outputs(1383);
    layer3_outputs(1789) <= not(layer2_outputs(6449));
    layer3_outputs(1790) <= not((layer2_outputs(3770)) and (layer2_outputs(1536)));
    layer3_outputs(1791) <= (layer2_outputs(1267)) and not (layer2_outputs(3047));
    layer3_outputs(1792) <= not(layer2_outputs(1737)) or (layer2_outputs(1934));
    layer3_outputs(1793) <= not((layer2_outputs(5481)) xor (layer2_outputs(1893)));
    layer3_outputs(1794) <= layer2_outputs(3068);
    layer3_outputs(1795) <= not(layer2_outputs(4750)) or (layer2_outputs(819));
    layer3_outputs(1796) <= layer2_outputs(4255);
    layer3_outputs(1797) <= not(layer2_outputs(6987));
    layer3_outputs(1798) <= not(layer2_outputs(3559)) or (layer2_outputs(1090));
    layer3_outputs(1799) <= not(layer2_outputs(4029));
    layer3_outputs(1800) <= '0';
    layer3_outputs(1801) <= not(layer2_outputs(732));
    layer3_outputs(1802) <= not(layer2_outputs(1022));
    layer3_outputs(1803) <= (layer2_outputs(1516)) or (layer2_outputs(3754));
    layer3_outputs(1804) <= (layer2_outputs(56)) xor (layer2_outputs(6838));
    layer3_outputs(1805) <= '0';
    layer3_outputs(1806) <= (layer2_outputs(4046)) and not (layer2_outputs(1256));
    layer3_outputs(1807) <= not(layer2_outputs(5286));
    layer3_outputs(1808) <= not(layer2_outputs(4314)) or (layer2_outputs(1718));
    layer3_outputs(1809) <= layer2_outputs(2569);
    layer3_outputs(1810) <= not((layer2_outputs(339)) and (layer2_outputs(159)));
    layer3_outputs(1811) <= not((layer2_outputs(5735)) or (layer2_outputs(7274)));
    layer3_outputs(1812) <= not(layer2_outputs(1178));
    layer3_outputs(1813) <= not(layer2_outputs(1579));
    layer3_outputs(1814) <= (layer2_outputs(4364)) xor (layer2_outputs(2405));
    layer3_outputs(1815) <= not(layer2_outputs(4200));
    layer3_outputs(1816) <= not(layer2_outputs(2554));
    layer3_outputs(1817) <= not(layer2_outputs(272));
    layer3_outputs(1818) <= not(layer2_outputs(1313)) or (layer2_outputs(738));
    layer3_outputs(1819) <= not(layer2_outputs(5808));
    layer3_outputs(1820) <= not(layer2_outputs(4882));
    layer3_outputs(1821) <= not((layer2_outputs(4465)) xor (layer2_outputs(1804)));
    layer3_outputs(1822) <= (layer2_outputs(1868)) and not (layer2_outputs(2041));
    layer3_outputs(1823) <= not(layer2_outputs(6058)) or (layer2_outputs(6827));
    layer3_outputs(1824) <= '0';
    layer3_outputs(1825) <= layer2_outputs(2399);
    layer3_outputs(1826) <= layer2_outputs(4777);
    layer3_outputs(1827) <= not(layer2_outputs(3067)) or (layer2_outputs(1778));
    layer3_outputs(1828) <= not(layer2_outputs(5391));
    layer3_outputs(1829) <= layer2_outputs(7144);
    layer3_outputs(1830) <= (layer2_outputs(6082)) xor (layer2_outputs(3878));
    layer3_outputs(1831) <= not(layer2_outputs(3484));
    layer3_outputs(1832) <= not(layer2_outputs(4564));
    layer3_outputs(1833) <= (layer2_outputs(2254)) and (layer2_outputs(1888));
    layer3_outputs(1834) <= not(layer2_outputs(4752));
    layer3_outputs(1835) <= layer2_outputs(1208);
    layer3_outputs(1836) <= layer2_outputs(5623);
    layer3_outputs(1837) <= '0';
    layer3_outputs(1838) <= not(layer2_outputs(6448));
    layer3_outputs(1839) <= not(layer2_outputs(2626));
    layer3_outputs(1840) <= not((layer2_outputs(3524)) or (layer2_outputs(7031)));
    layer3_outputs(1841) <= (layer2_outputs(1624)) and not (layer2_outputs(656));
    layer3_outputs(1842) <= (layer2_outputs(1450)) and not (layer2_outputs(5637));
    layer3_outputs(1843) <= not((layer2_outputs(3917)) xor (layer2_outputs(4778)));
    layer3_outputs(1844) <= layer2_outputs(430);
    layer3_outputs(1845) <= not((layer2_outputs(6596)) or (layer2_outputs(2390)));
    layer3_outputs(1846) <= not(layer2_outputs(1565));
    layer3_outputs(1847) <= not((layer2_outputs(1199)) or (layer2_outputs(3271)));
    layer3_outputs(1848) <= not(layer2_outputs(3064)) or (layer2_outputs(7554));
    layer3_outputs(1849) <= not(layer2_outputs(3369));
    layer3_outputs(1850) <= (layer2_outputs(3990)) and (layer2_outputs(2929));
    layer3_outputs(1851) <= not(layer2_outputs(4634)) or (layer2_outputs(219));
    layer3_outputs(1852) <= (layer2_outputs(5995)) or (layer2_outputs(4323));
    layer3_outputs(1853) <= layer2_outputs(1845);
    layer3_outputs(1854) <= '0';
    layer3_outputs(1855) <= not((layer2_outputs(5066)) xor (layer2_outputs(979)));
    layer3_outputs(1856) <= not((layer2_outputs(2065)) or (layer2_outputs(3721)));
    layer3_outputs(1857) <= (layer2_outputs(5441)) or (layer2_outputs(5663));
    layer3_outputs(1858) <= (layer2_outputs(7105)) and (layer2_outputs(2167));
    layer3_outputs(1859) <= '0';
    layer3_outputs(1860) <= not((layer2_outputs(2149)) and (layer2_outputs(276)));
    layer3_outputs(1861) <= (layer2_outputs(3960)) and (layer2_outputs(2024));
    layer3_outputs(1862) <= not((layer2_outputs(3228)) or (layer2_outputs(3665)));
    layer3_outputs(1863) <= not(layer2_outputs(3945));
    layer3_outputs(1864) <= layer2_outputs(5157);
    layer3_outputs(1865) <= '1';
    layer3_outputs(1866) <= (layer2_outputs(302)) and (layer2_outputs(7391));
    layer3_outputs(1867) <= not((layer2_outputs(1140)) or (layer2_outputs(1087)));
    layer3_outputs(1868) <= layer2_outputs(6941);
    layer3_outputs(1869) <= not((layer2_outputs(1302)) or (layer2_outputs(1303)));
    layer3_outputs(1870) <= not(layer2_outputs(7464));
    layer3_outputs(1871) <= not((layer2_outputs(6920)) or (layer2_outputs(7318)));
    layer3_outputs(1872) <= not((layer2_outputs(3796)) xor (layer2_outputs(6195)));
    layer3_outputs(1873) <= not(layer2_outputs(3314)) or (layer2_outputs(4677));
    layer3_outputs(1874) <= not(layer2_outputs(3762));
    layer3_outputs(1875) <= layer2_outputs(627);
    layer3_outputs(1876) <= not((layer2_outputs(3188)) or (layer2_outputs(5112)));
    layer3_outputs(1877) <= not((layer2_outputs(945)) and (layer2_outputs(5411)));
    layer3_outputs(1878) <= (layer2_outputs(2233)) xor (layer2_outputs(7118));
    layer3_outputs(1879) <= not(layer2_outputs(4980));
    layer3_outputs(1880) <= not(layer2_outputs(1918)) or (layer2_outputs(3137));
    layer3_outputs(1881) <= layer2_outputs(3932);
    layer3_outputs(1882) <= not((layer2_outputs(6768)) xor (layer2_outputs(7182)));
    layer3_outputs(1883) <= not((layer2_outputs(7081)) or (layer2_outputs(3822)));
    layer3_outputs(1884) <= (layer2_outputs(7273)) and (layer2_outputs(2662));
    layer3_outputs(1885) <= not(layer2_outputs(4149));
    layer3_outputs(1886) <= not(layer2_outputs(3591));
    layer3_outputs(1887) <= (layer2_outputs(639)) or (layer2_outputs(2787));
    layer3_outputs(1888) <= not(layer2_outputs(7605));
    layer3_outputs(1889) <= layer2_outputs(6340);
    layer3_outputs(1890) <= not((layer2_outputs(6281)) xor (layer2_outputs(1240)));
    layer3_outputs(1891) <= not(layer2_outputs(4374)) or (layer2_outputs(152));
    layer3_outputs(1892) <= (layer2_outputs(4569)) and not (layer2_outputs(5811));
    layer3_outputs(1893) <= not(layer2_outputs(3478)) or (layer2_outputs(6866));
    layer3_outputs(1894) <= layer2_outputs(299);
    layer3_outputs(1895) <= layer2_outputs(2534);
    layer3_outputs(1896) <= not(layer2_outputs(5913)) or (layer2_outputs(1358));
    layer3_outputs(1897) <= not(layer2_outputs(1340)) or (layer2_outputs(526));
    layer3_outputs(1898) <= not(layer2_outputs(2033));
    layer3_outputs(1899) <= '0';
    layer3_outputs(1900) <= not(layer2_outputs(2294)) or (layer2_outputs(2182));
    layer3_outputs(1901) <= layer2_outputs(6717);
    layer3_outputs(1902) <= not(layer2_outputs(5449)) or (layer2_outputs(4193));
    layer3_outputs(1903) <= not(layer2_outputs(7198));
    layer3_outputs(1904) <= '1';
    layer3_outputs(1905) <= (layer2_outputs(1552)) and (layer2_outputs(3376));
    layer3_outputs(1906) <= (layer2_outputs(2982)) and not (layer2_outputs(3966));
    layer3_outputs(1907) <= '0';
    layer3_outputs(1908) <= not((layer2_outputs(4862)) xor (layer2_outputs(2045)));
    layer3_outputs(1909) <= (layer2_outputs(1924)) and not (layer2_outputs(2578));
    layer3_outputs(1910) <= not((layer2_outputs(7357)) or (layer2_outputs(6940)));
    layer3_outputs(1911) <= (layer2_outputs(4851)) or (layer2_outputs(2751));
    layer3_outputs(1912) <= (layer2_outputs(230)) and not (layer2_outputs(5374));
    layer3_outputs(1913) <= '0';
    layer3_outputs(1914) <= layer2_outputs(7593);
    layer3_outputs(1915) <= not(layer2_outputs(4604));
    layer3_outputs(1916) <= layer2_outputs(5323);
    layer3_outputs(1917) <= not(layer2_outputs(2087)) or (layer2_outputs(1894));
    layer3_outputs(1918) <= (layer2_outputs(5671)) or (layer2_outputs(3070));
    layer3_outputs(1919) <= not(layer2_outputs(3564)) or (layer2_outputs(6105));
    layer3_outputs(1920) <= (layer2_outputs(6687)) or (layer2_outputs(5461));
    layer3_outputs(1921) <= not(layer2_outputs(1596));
    layer3_outputs(1922) <= not((layer2_outputs(2371)) or (layer2_outputs(3330)));
    layer3_outputs(1923) <= (layer2_outputs(43)) and not (layer2_outputs(402));
    layer3_outputs(1924) <= not(layer2_outputs(6654));
    layer3_outputs(1925) <= not(layer2_outputs(3912));
    layer3_outputs(1926) <= (layer2_outputs(7642)) or (layer2_outputs(4755));
    layer3_outputs(1927) <= not((layer2_outputs(1454)) or (layer2_outputs(3944)));
    layer3_outputs(1928) <= '0';
    layer3_outputs(1929) <= layer2_outputs(7353);
    layer3_outputs(1930) <= not(layer2_outputs(3251)) or (layer2_outputs(5415));
    layer3_outputs(1931) <= (layer2_outputs(3999)) and (layer2_outputs(297));
    layer3_outputs(1932) <= not((layer2_outputs(3587)) or (layer2_outputs(918)));
    layer3_outputs(1933) <= not((layer2_outputs(3135)) or (layer2_outputs(1464)));
    layer3_outputs(1934) <= '1';
    layer3_outputs(1935) <= (layer2_outputs(3987)) and not (layer2_outputs(5407));
    layer3_outputs(1936) <= not(layer2_outputs(114));
    layer3_outputs(1937) <= not(layer2_outputs(7219));
    layer3_outputs(1938) <= (layer2_outputs(3478)) and not (layer2_outputs(3103));
    layer3_outputs(1939) <= layer2_outputs(2271);
    layer3_outputs(1940) <= not(layer2_outputs(7407));
    layer3_outputs(1941) <= not(layer2_outputs(7504)) or (layer2_outputs(6635));
    layer3_outputs(1942) <= layer2_outputs(4006);
    layer3_outputs(1943) <= (layer2_outputs(2663)) and not (layer2_outputs(3822));
    layer3_outputs(1944) <= not(layer2_outputs(6078));
    layer3_outputs(1945) <= not(layer2_outputs(736));
    layer3_outputs(1946) <= not(layer2_outputs(4770));
    layer3_outputs(1947) <= not(layer2_outputs(7327));
    layer3_outputs(1948) <= (layer2_outputs(3515)) or (layer2_outputs(680));
    layer3_outputs(1949) <= (layer2_outputs(976)) and not (layer2_outputs(2118));
    layer3_outputs(1950) <= layer2_outputs(4285);
    layer3_outputs(1951) <= not(layer2_outputs(767));
    layer3_outputs(1952) <= (layer2_outputs(5235)) xor (layer2_outputs(3821));
    layer3_outputs(1953) <= layer2_outputs(5841);
    layer3_outputs(1954) <= not(layer2_outputs(2534)) or (layer2_outputs(553));
    layer3_outputs(1955) <= not(layer2_outputs(2247));
    layer3_outputs(1956) <= not((layer2_outputs(6670)) or (layer2_outputs(5327)));
    layer3_outputs(1957) <= not(layer2_outputs(5066)) or (layer2_outputs(4031));
    layer3_outputs(1958) <= layer2_outputs(4647);
    layer3_outputs(1959) <= (layer2_outputs(2048)) and not (layer2_outputs(5028));
    layer3_outputs(1960) <= (layer2_outputs(5129)) and not (layer2_outputs(1686));
    layer3_outputs(1961) <= (layer2_outputs(5666)) and not (layer2_outputs(4023));
    layer3_outputs(1962) <= not(layer2_outputs(5755));
    layer3_outputs(1963) <= not((layer2_outputs(360)) or (layer2_outputs(6685)));
    layer3_outputs(1964) <= (layer2_outputs(591)) and not (layer2_outputs(3222));
    layer3_outputs(1965) <= layer2_outputs(3609);
    layer3_outputs(1966) <= not((layer2_outputs(730)) xor (layer2_outputs(269)));
    layer3_outputs(1967) <= not((layer2_outputs(900)) or (layer2_outputs(1449)));
    layer3_outputs(1968) <= not(layer2_outputs(2086)) or (layer2_outputs(5574));
    layer3_outputs(1969) <= layer2_outputs(6372);
    layer3_outputs(1970) <= (layer2_outputs(6319)) and (layer2_outputs(2300));
    layer3_outputs(1971) <= layer2_outputs(986);
    layer3_outputs(1972) <= not(layer2_outputs(666)) or (layer2_outputs(7056));
    layer3_outputs(1973) <= not((layer2_outputs(7072)) xor (layer2_outputs(3223)));
    layer3_outputs(1974) <= not(layer2_outputs(1679));
    layer3_outputs(1975) <= not(layer2_outputs(7109));
    layer3_outputs(1976) <= not(layer2_outputs(2314));
    layer3_outputs(1977) <= (layer2_outputs(6545)) and not (layer2_outputs(3923));
    layer3_outputs(1978) <= not(layer2_outputs(121)) or (layer2_outputs(4408));
    layer3_outputs(1979) <= not(layer2_outputs(2594));
    layer3_outputs(1980) <= not((layer2_outputs(6875)) or (layer2_outputs(1216)));
    layer3_outputs(1981) <= not(layer2_outputs(5875));
    layer3_outputs(1982) <= not(layer2_outputs(5033)) or (layer2_outputs(1780));
    layer3_outputs(1983) <= '1';
    layer3_outputs(1984) <= layer2_outputs(3955);
    layer3_outputs(1985) <= not(layer2_outputs(3803));
    layer3_outputs(1986) <= (layer2_outputs(6458)) or (layer2_outputs(7505));
    layer3_outputs(1987) <= layer2_outputs(4316);
    layer3_outputs(1988) <= (layer2_outputs(4297)) or (layer2_outputs(961));
    layer3_outputs(1989) <= not(layer2_outputs(902));
    layer3_outputs(1990) <= not(layer2_outputs(4823)) or (layer2_outputs(5497));
    layer3_outputs(1991) <= not((layer2_outputs(2515)) and (layer2_outputs(4507)));
    layer3_outputs(1992) <= not(layer2_outputs(6318)) or (layer2_outputs(3733));
    layer3_outputs(1993) <= not(layer2_outputs(5244));
    layer3_outputs(1994) <= (layer2_outputs(314)) and not (layer2_outputs(1724));
    layer3_outputs(1995) <= layer2_outputs(6854);
    layer3_outputs(1996) <= layer2_outputs(7238);
    layer3_outputs(1997) <= not(layer2_outputs(601));
    layer3_outputs(1998) <= not(layer2_outputs(3693));
    layer3_outputs(1999) <= not(layer2_outputs(5898)) or (layer2_outputs(4802));
    layer3_outputs(2000) <= layer2_outputs(2971);
    layer3_outputs(2001) <= layer2_outputs(3216);
    layer3_outputs(2002) <= (layer2_outputs(4447)) and not (layer2_outputs(7441));
    layer3_outputs(2003) <= layer2_outputs(3815);
    layer3_outputs(2004) <= (layer2_outputs(2445)) and not (layer2_outputs(644));
    layer3_outputs(2005) <= not((layer2_outputs(5082)) xor (layer2_outputs(2292)));
    layer3_outputs(2006) <= not((layer2_outputs(7649)) or (layer2_outputs(6031)));
    layer3_outputs(2007) <= (layer2_outputs(7228)) and (layer2_outputs(5404));
    layer3_outputs(2008) <= (layer2_outputs(6474)) and not (layer2_outputs(4816));
    layer3_outputs(2009) <= layer2_outputs(2239);
    layer3_outputs(2010) <= not((layer2_outputs(3769)) and (layer2_outputs(2971)));
    layer3_outputs(2011) <= '1';
    layer3_outputs(2012) <= '1';
    layer3_outputs(2013) <= '1';
    layer3_outputs(2014) <= not(layer2_outputs(3200)) or (layer2_outputs(6216));
    layer3_outputs(2015) <= (layer2_outputs(7064)) and not (layer2_outputs(4056));
    layer3_outputs(2016) <= '1';
    layer3_outputs(2017) <= not((layer2_outputs(6416)) xor (layer2_outputs(2124)));
    layer3_outputs(2018) <= (layer2_outputs(223)) and not (layer2_outputs(4638));
    layer3_outputs(2019) <= not((layer2_outputs(4250)) or (layer2_outputs(4100)));
    layer3_outputs(2020) <= layer2_outputs(5089);
    layer3_outputs(2021) <= not(layer2_outputs(6788));
    layer3_outputs(2022) <= layer2_outputs(7269);
    layer3_outputs(2023) <= not((layer2_outputs(5328)) or (layer2_outputs(5492)));
    layer3_outputs(2024) <= layer2_outputs(932);
    layer3_outputs(2025) <= (layer2_outputs(967)) and not (layer2_outputs(7326));
    layer3_outputs(2026) <= not(layer2_outputs(210)) or (layer2_outputs(3672));
    layer3_outputs(2027) <= (layer2_outputs(6270)) and not (layer2_outputs(1013));
    layer3_outputs(2028) <= (layer2_outputs(5341)) and not (layer2_outputs(4215));
    layer3_outputs(2029) <= not(layer2_outputs(6552));
    layer3_outputs(2030) <= '0';
    layer3_outputs(2031) <= not(layer2_outputs(4611)) or (layer2_outputs(1668));
    layer3_outputs(2032) <= (layer2_outputs(6528)) and not (layer2_outputs(7328));
    layer3_outputs(2033) <= layer2_outputs(766);
    layer3_outputs(2034) <= layer2_outputs(7621);
    layer3_outputs(2035) <= not(layer2_outputs(4741));
    layer3_outputs(2036) <= not(layer2_outputs(857)) or (layer2_outputs(4660));
    layer3_outputs(2037) <= not((layer2_outputs(6205)) or (layer2_outputs(3954)));
    layer3_outputs(2038) <= not(layer2_outputs(678)) or (layer2_outputs(1758));
    layer3_outputs(2039) <= not(layer2_outputs(5915));
    layer3_outputs(2040) <= '1';
    layer3_outputs(2041) <= '0';
    layer3_outputs(2042) <= not((layer2_outputs(729)) and (layer2_outputs(6794)));
    layer3_outputs(2043) <= not(layer2_outputs(6801)) or (layer2_outputs(2403));
    layer3_outputs(2044) <= not(layer2_outputs(4383));
    layer3_outputs(2045) <= (layer2_outputs(6771)) and not (layer2_outputs(4317));
    layer3_outputs(2046) <= not(layer2_outputs(2659)) or (layer2_outputs(1196));
    layer3_outputs(2047) <= (layer2_outputs(4456)) and not (layer2_outputs(1833));
    layer3_outputs(2048) <= not(layer2_outputs(1125));
    layer3_outputs(2049) <= not(layer2_outputs(5200)) or (layer2_outputs(3679));
    layer3_outputs(2050) <= not(layer2_outputs(4203));
    layer3_outputs(2051) <= not(layer2_outputs(6906)) or (layer2_outputs(7047));
    layer3_outputs(2052) <= not((layer2_outputs(7170)) or (layer2_outputs(6977)));
    layer3_outputs(2053) <= (layer2_outputs(3288)) and not (layer2_outputs(7305));
    layer3_outputs(2054) <= not(layer2_outputs(1377));
    layer3_outputs(2055) <= '1';
    layer3_outputs(2056) <= not((layer2_outputs(6231)) xor (layer2_outputs(5249)));
    layer3_outputs(2057) <= (layer2_outputs(3532)) and (layer2_outputs(4750));
    layer3_outputs(2058) <= not(layer2_outputs(3311));
    layer3_outputs(2059) <= layer2_outputs(4370);
    layer3_outputs(2060) <= not((layer2_outputs(767)) or (layer2_outputs(2221)));
    layer3_outputs(2061) <= layer2_outputs(4450);
    layer3_outputs(2062) <= not(layer2_outputs(2283));
    layer3_outputs(2063) <= (layer2_outputs(2125)) and (layer2_outputs(6691));
    layer3_outputs(2064) <= (layer2_outputs(3371)) and not (layer2_outputs(3046));
    layer3_outputs(2065) <= (layer2_outputs(5577)) and not (layer2_outputs(440));
    layer3_outputs(2066) <= '1';
    layer3_outputs(2067) <= '1';
    layer3_outputs(2068) <= '0';
    layer3_outputs(2069) <= (layer2_outputs(1906)) and (layer2_outputs(7220));
    layer3_outputs(2070) <= (layer2_outputs(267)) and not (layer2_outputs(3126));
    layer3_outputs(2071) <= layer2_outputs(5838);
    layer3_outputs(2072) <= not(layer2_outputs(2636));
    layer3_outputs(2073) <= '1';
    layer3_outputs(2074) <= not(layer2_outputs(3625));
    layer3_outputs(2075) <= not(layer2_outputs(420)) or (layer2_outputs(5194));
    layer3_outputs(2076) <= '1';
    layer3_outputs(2077) <= not(layer2_outputs(2047)) or (layer2_outputs(1194));
    layer3_outputs(2078) <= (layer2_outputs(3848)) and not (layer2_outputs(3582));
    layer3_outputs(2079) <= (layer2_outputs(6219)) and not (layer2_outputs(3462));
    layer3_outputs(2080) <= not(layer2_outputs(5283));
    layer3_outputs(2081) <= '0';
    layer3_outputs(2082) <= (layer2_outputs(433)) and not (layer2_outputs(3000));
    layer3_outputs(2083) <= (layer2_outputs(6302)) and not (layer2_outputs(818));
    layer3_outputs(2084) <= layer2_outputs(3818);
    layer3_outputs(2085) <= '0';
    layer3_outputs(2086) <= not((layer2_outputs(6076)) xor (layer2_outputs(2132)));
    layer3_outputs(2087) <= (layer2_outputs(368)) and (layer2_outputs(3270));
    layer3_outputs(2088) <= not((layer2_outputs(1105)) xor (layer2_outputs(7247)));
    layer3_outputs(2089) <= (layer2_outputs(7502)) and (layer2_outputs(5332));
    layer3_outputs(2090) <= '0';
    layer3_outputs(2091) <= '0';
    layer3_outputs(2092) <= (layer2_outputs(4139)) or (layer2_outputs(1995));
    layer3_outputs(2093) <= not((layer2_outputs(6709)) xor (layer2_outputs(2813)));
    layer3_outputs(2094) <= not(layer2_outputs(4720));
    layer3_outputs(2095) <= (layer2_outputs(5572)) or (layer2_outputs(516));
    layer3_outputs(2096) <= not(layer2_outputs(189));
    layer3_outputs(2097) <= layer2_outputs(3377);
    layer3_outputs(2098) <= (layer2_outputs(4805)) or (layer2_outputs(4597));
    layer3_outputs(2099) <= layer2_outputs(2286);
    layer3_outputs(2100) <= '1';
    layer3_outputs(2101) <= not(layer2_outputs(6310));
    layer3_outputs(2102) <= (layer2_outputs(7278)) and not (layer2_outputs(6297));
    layer3_outputs(2103) <= (layer2_outputs(3092)) and not (layer2_outputs(1280));
    layer3_outputs(2104) <= (layer2_outputs(2696)) and not (layer2_outputs(4371));
    layer3_outputs(2105) <= (layer2_outputs(2002)) or (layer2_outputs(4629));
    layer3_outputs(2106) <= layer2_outputs(5199);
    layer3_outputs(2107) <= layer2_outputs(1516);
    layer3_outputs(2108) <= layer2_outputs(5806);
    layer3_outputs(2109) <= layer2_outputs(4125);
    layer3_outputs(2110) <= layer2_outputs(205);
    layer3_outputs(2111) <= layer2_outputs(1150);
    layer3_outputs(2112) <= '0';
    layer3_outputs(2113) <= not(layer2_outputs(3938));
    layer3_outputs(2114) <= '1';
    layer3_outputs(2115) <= not((layer2_outputs(1811)) or (layer2_outputs(5928)));
    layer3_outputs(2116) <= not((layer2_outputs(454)) and (layer2_outputs(5288)));
    layer3_outputs(2117) <= '0';
    layer3_outputs(2118) <= not((layer2_outputs(1460)) and (layer2_outputs(2217)));
    layer3_outputs(2119) <= (layer2_outputs(4469)) and (layer2_outputs(1544));
    layer3_outputs(2120) <= not(layer2_outputs(316));
    layer3_outputs(2121) <= '0';
    layer3_outputs(2122) <= not(layer2_outputs(6898));
    layer3_outputs(2123) <= layer2_outputs(6110);
    layer3_outputs(2124) <= '1';
    layer3_outputs(2125) <= '0';
    layer3_outputs(2126) <= not(layer2_outputs(6305));
    layer3_outputs(2127) <= not(layer2_outputs(7248));
    layer3_outputs(2128) <= '0';
    layer3_outputs(2129) <= not((layer2_outputs(560)) or (layer2_outputs(3977)));
    layer3_outputs(2130) <= not(layer2_outputs(7622));
    layer3_outputs(2131) <= layer2_outputs(6410);
    layer3_outputs(2132) <= layer2_outputs(1760);
    layer3_outputs(2133) <= '0';
    layer3_outputs(2134) <= not(layer2_outputs(6960)) or (layer2_outputs(1744));
    layer3_outputs(2135) <= (layer2_outputs(3437)) and (layer2_outputs(2329));
    layer3_outputs(2136) <= not(layer2_outputs(2820));
    layer3_outputs(2137) <= not(layer2_outputs(4972));
    layer3_outputs(2138) <= not(layer2_outputs(583));
    layer3_outputs(2139) <= layer2_outputs(4225);
    layer3_outputs(2140) <= (layer2_outputs(7214)) and not (layer2_outputs(2172));
    layer3_outputs(2141) <= (layer2_outputs(3387)) or (layer2_outputs(5524));
    layer3_outputs(2142) <= layer2_outputs(1572);
    layer3_outputs(2143) <= not(layer2_outputs(1329));
    layer3_outputs(2144) <= (layer2_outputs(3111)) or (layer2_outputs(6519));
    layer3_outputs(2145) <= not(layer2_outputs(558));
    layer3_outputs(2146) <= layer2_outputs(5226);
    layer3_outputs(2147) <= not(layer2_outputs(3392)) or (layer2_outputs(904));
    layer3_outputs(2148) <= (layer2_outputs(6464)) and not (layer2_outputs(6514));
    layer3_outputs(2149) <= not(layer2_outputs(7317)) or (layer2_outputs(1602));
    layer3_outputs(2150) <= not(layer2_outputs(796));
    layer3_outputs(2151) <= not(layer2_outputs(2227));
    layer3_outputs(2152) <= (layer2_outputs(2583)) or (layer2_outputs(6469));
    layer3_outputs(2153) <= not((layer2_outputs(4389)) and (layer2_outputs(1726)));
    layer3_outputs(2154) <= (layer2_outputs(5849)) and not (layer2_outputs(4236));
    layer3_outputs(2155) <= (layer2_outputs(2120)) and not (layer2_outputs(1270));
    layer3_outputs(2156) <= (layer2_outputs(2589)) xor (layer2_outputs(1782));
    layer3_outputs(2157) <= (layer2_outputs(131)) and (layer2_outputs(6889));
    layer3_outputs(2158) <= (layer2_outputs(1738)) or (layer2_outputs(960));
    layer3_outputs(2159) <= (layer2_outputs(288)) and not (layer2_outputs(6163));
    layer3_outputs(2160) <= not(layer2_outputs(1148)) or (layer2_outputs(6196));
    layer3_outputs(2161) <= layer2_outputs(426);
    layer3_outputs(2162) <= '0';
    layer3_outputs(2163) <= not((layer2_outputs(3038)) and (layer2_outputs(6765)));
    layer3_outputs(2164) <= not(layer2_outputs(1433));
    layer3_outputs(2165) <= not(layer2_outputs(5439)) or (layer2_outputs(6363));
    layer3_outputs(2166) <= layer2_outputs(1285);
    layer3_outputs(2167) <= (layer2_outputs(258)) or (layer2_outputs(2291));
    layer3_outputs(2168) <= not(layer2_outputs(1777));
    layer3_outputs(2169) <= layer2_outputs(4165);
    layer3_outputs(2170) <= layer2_outputs(1462);
    layer3_outputs(2171) <= not((layer2_outputs(6039)) or (layer2_outputs(7453)));
    layer3_outputs(2172) <= not(layer2_outputs(3774)) or (layer2_outputs(6775));
    layer3_outputs(2173) <= '0';
    layer3_outputs(2174) <= not((layer2_outputs(6903)) or (layer2_outputs(5705)));
    layer3_outputs(2175) <= (layer2_outputs(5820)) xor (layer2_outputs(3519));
    layer3_outputs(2176) <= not(layer2_outputs(5727)) or (layer2_outputs(4308));
    layer3_outputs(2177) <= not(layer2_outputs(6596));
    layer3_outputs(2178) <= (layer2_outputs(858)) or (layer2_outputs(4501));
    layer3_outputs(2179) <= not((layer2_outputs(694)) or (layer2_outputs(919)));
    layer3_outputs(2180) <= not(layer2_outputs(2794));
    layer3_outputs(2181) <= '1';
    layer3_outputs(2182) <= (layer2_outputs(2045)) xor (layer2_outputs(2278));
    layer3_outputs(2183) <= not(layer2_outputs(547));
    layer3_outputs(2184) <= not(layer2_outputs(3675));
    layer3_outputs(2185) <= not(layer2_outputs(6441)) or (layer2_outputs(4784));
    layer3_outputs(2186) <= '1';
    layer3_outputs(2187) <= not(layer2_outputs(5947));
    layer3_outputs(2188) <= (layer2_outputs(1143)) and not (layer2_outputs(3732));
    layer3_outputs(2189) <= layer2_outputs(6160);
    layer3_outputs(2190) <= not(layer2_outputs(3924)) or (layer2_outputs(3962));
    layer3_outputs(2191) <= (layer2_outputs(3321)) or (layer2_outputs(5756));
    layer3_outputs(2192) <= (layer2_outputs(1915)) or (layer2_outputs(5684));
    layer3_outputs(2193) <= (layer2_outputs(3598)) and not (layer2_outputs(3405));
    layer3_outputs(2194) <= layer2_outputs(7639);
    layer3_outputs(2195) <= not(layer2_outputs(1979));
    layer3_outputs(2196) <= not((layer2_outputs(5501)) and (layer2_outputs(5624)));
    layer3_outputs(2197) <= (layer2_outputs(2153)) and (layer2_outputs(6855));
    layer3_outputs(2198) <= (layer2_outputs(6156)) and (layer2_outputs(2898));
    layer3_outputs(2199) <= not(layer2_outputs(4841)) or (layer2_outputs(7287));
    layer3_outputs(2200) <= not(layer2_outputs(1672));
    layer3_outputs(2201) <= (layer2_outputs(6768)) and (layer2_outputs(5080));
    layer3_outputs(2202) <= not(layer2_outputs(7025));
    layer3_outputs(2203) <= not(layer2_outputs(703));
    layer3_outputs(2204) <= not(layer2_outputs(2295)) or (layer2_outputs(1186));
    layer3_outputs(2205) <= not((layer2_outputs(7539)) and (layer2_outputs(2500)));
    layer3_outputs(2206) <= not(layer2_outputs(3949)) or (layer2_outputs(1451));
    layer3_outputs(2207) <= not((layer2_outputs(3972)) and (layer2_outputs(1306)));
    layer3_outputs(2208) <= layer2_outputs(6475);
    layer3_outputs(2209) <= (layer2_outputs(1736)) and not (layer2_outputs(3170));
    layer3_outputs(2210) <= layer2_outputs(5864);
    layer3_outputs(2211) <= not((layer2_outputs(4668)) xor (layer2_outputs(4254)));
    layer3_outputs(2212) <= '0';
    layer3_outputs(2213) <= layer2_outputs(4046);
    layer3_outputs(2214) <= not((layer2_outputs(4038)) xor (layer2_outputs(3077)));
    layer3_outputs(2215) <= layer2_outputs(3817);
    layer3_outputs(2216) <= (layer2_outputs(6004)) and not (layer2_outputs(4857));
    layer3_outputs(2217) <= not((layer2_outputs(1721)) or (layer2_outputs(555)));
    layer3_outputs(2218) <= not(layer2_outputs(1546)) or (layer2_outputs(3586));
    layer3_outputs(2219) <= (layer2_outputs(4154)) and (layer2_outputs(5717));
    layer3_outputs(2220) <= '0';
    layer3_outputs(2221) <= not(layer2_outputs(6249));
    layer3_outputs(2222) <= not(layer2_outputs(716));
    layer3_outputs(2223) <= '0';
    layer3_outputs(2224) <= '1';
    layer3_outputs(2225) <= not(layer2_outputs(1853));
    layer3_outputs(2226) <= not(layer2_outputs(2512));
    layer3_outputs(2227) <= (layer2_outputs(6507)) and (layer2_outputs(1683));
    layer3_outputs(2228) <= not((layer2_outputs(1504)) and (layer2_outputs(2687)));
    layer3_outputs(2229) <= layer2_outputs(4917);
    layer3_outputs(2230) <= not((layer2_outputs(2529)) and (layer2_outputs(1162)));
    layer3_outputs(2231) <= layer2_outputs(7552);
    layer3_outputs(2232) <= (layer2_outputs(896)) and (layer2_outputs(4086));
    layer3_outputs(2233) <= not(layer2_outputs(3550)) or (layer2_outputs(7546));
    layer3_outputs(2234) <= '1';
    layer3_outputs(2235) <= not(layer2_outputs(282)) or (layer2_outputs(3331));
    layer3_outputs(2236) <= layer2_outputs(6868);
    layer3_outputs(2237) <= not((layer2_outputs(4857)) or (layer2_outputs(4185)));
    layer3_outputs(2238) <= not((layer2_outputs(657)) or (layer2_outputs(7288)));
    layer3_outputs(2239) <= not((layer2_outputs(3020)) or (layer2_outputs(7425)));
    layer3_outputs(2240) <= not(layer2_outputs(5982));
    layer3_outputs(2241) <= not(layer2_outputs(2980)) or (layer2_outputs(5520));
    layer3_outputs(2242) <= not(layer2_outputs(655));
    layer3_outputs(2243) <= not((layer2_outputs(1230)) and (layer2_outputs(2638)));
    layer3_outputs(2244) <= layer2_outputs(917);
    layer3_outputs(2245) <= (layer2_outputs(1886)) and not (layer2_outputs(4969));
    layer3_outputs(2246) <= not(layer2_outputs(157));
    layer3_outputs(2247) <= '1';
    layer3_outputs(2248) <= not((layer2_outputs(6705)) and (layer2_outputs(6278)));
    layer3_outputs(2249) <= not(layer2_outputs(5312)) or (layer2_outputs(67));
    layer3_outputs(2250) <= not((layer2_outputs(3995)) or (layer2_outputs(5657)));
    layer3_outputs(2251) <= not(layer2_outputs(2757));
    layer3_outputs(2252) <= (layer2_outputs(1056)) or (layer2_outputs(3257));
    layer3_outputs(2253) <= not(layer2_outputs(2335)) or (layer2_outputs(5994));
    layer3_outputs(2254) <= not(layer2_outputs(7290));
    layer3_outputs(2255) <= layer2_outputs(672);
    layer3_outputs(2256) <= (layer2_outputs(5419)) and not (layer2_outputs(1971));
    layer3_outputs(2257) <= (layer2_outputs(2607)) and not (layer2_outputs(5000));
    layer3_outputs(2258) <= (layer2_outputs(6976)) or (layer2_outputs(5570));
    layer3_outputs(2259) <= '0';
    layer3_outputs(2260) <= not(layer2_outputs(3248)) or (layer2_outputs(7251));
    layer3_outputs(2261) <= not(layer2_outputs(6687));
    layer3_outputs(2262) <= '0';
    layer3_outputs(2263) <= (layer2_outputs(7276)) and (layer2_outputs(1738));
    layer3_outputs(2264) <= not(layer2_outputs(3910)) or (layer2_outputs(3148));
    layer3_outputs(2265) <= '1';
    layer3_outputs(2266) <= (layer2_outputs(3247)) and (layer2_outputs(406));
    layer3_outputs(2267) <= not(layer2_outputs(6358)) or (layer2_outputs(6090));
    layer3_outputs(2268) <= (layer2_outputs(6457)) and not (layer2_outputs(2884));
    layer3_outputs(2269) <= (layer2_outputs(6500)) and (layer2_outputs(3416));
    layer3_outputs(2270) <= (layer2_outputs(1643)) and not (layer2_outputs(891));
    layer3_outputs(2271) <= '0';
    layer3_outputs(2272) <= (layer2_outputs(7652)) xor (layer2_outputs(7093));
    layer3_outputs(2273) <= '0';
    layer3_outputs(2274) <= '0';
    layer3_outputs(2275) <= not(layer2_outputs(2021));
    layer3_outputs(2276) <= not((layer2_outputs(32)) xor (layer2_outputs(1928)));
    layer3_outputs(2277) <= not(layer2_outputs(5593));
    layer3_outputs(2278) <= not(layer2_outputs(2272));
    layer3_outputs(2279) <= layer2_outputs(6255);
    layer3_outputs(2280) <= not((layer2_outputs(3015)) and (layer2_outputs(6844)));
    layer3_outputs(2281) <= not(layer2_outputs(2527));
    layer3_outputs(2282) <= layer2_outputs(4890);
    layer3_outputs(2283) <= not(layer2_outputs(6811));
    layer3_outputs(2284) <= not(layer2_outputs(7008));
    layer3_outputs(2285) <= layer2_outputs(1186);
    layer3_outputs(2286) <= layer2_outputs(6574);
    layer3_outputs(2287) <= not(layer2_outputs(4174));
    layer3_outputs(2288) <= not(layer2_outputs(6452)) or (layer2_outputs(3524));
    layer3_outputs(2289) <= (layer2_outputs(6240)) and not (layer2_outputs(3146));
    layer3_outputs(2290) <= layer2_outputs(3836);
    layer3_outputs(2291) <= (layer2_outputs(3914)) and not (layer2_outputs(6306));
    layer3_outputs(2292) <= (layer2_outputs(1224)) or (layer2_outputs(4748));
    layer3_outputs(2293) <= (layer2_outputs(4955)) or (layer2_outputs(661));
    layer3_outputs(2294) <= not(layer2_outputs(4026)) or (layer2_outputs(4796));
    layer3_outputs(2295) <= layer2_outputs(6598);
    layer3_outputs(2296) <= (layer2_outputs(7194)) and not (layer2_outputs(4439));
    layer3_outputs(2297) <= (layer2_outputs(3790)) and (layer2_outputs(3398));
    layer3_outputs(2298) <= not(layer2_outputs(234)) or (layer2_outputs(5043));
    layer3_outputs(2299) <= not(layer2_outputs(6019));
    layer3_outputs(2300) <= not(layer2_outputs(4649)) or (layer2_outputs(3029));
    layer3_outputs(2301) <= not(layer2_outputs(3673)) or (layer2_outputs(800));
    layer3_outputs(2302) <= layer2_outputs(747);
    layer3_outputs(2303) <= (layer2_outputs(3389)) and not (layer2_outputs(2282));
    layer3_outputs(2304) <= not((layer2_outputs(6313)) and (layer2_outputs(6794)));
    layer3_outputs(2305) <= (layer2_outputs(4566)) and not (layer2_outputs(3492));
    layer3_outputs(2306) <= not(layer2_outputs(587)) or (layer2_outputs(2498));
    layer3_outputs(2307) <= not((layer2_outputs(3323)) and (layer2_outputs(6855)));
    layer3_outputs(2308) <= not(layer2_outputs(7344)) or (layer2_outputs(191));
    layer3_outputs(2309) <= not((layer2_outputs(5520)) or (layer2_outputs(5796)));
    layer3_outputs(2310) <= (layer2_outputs(2816)) or (layer2_outputs(6002));
    layer3_outputs(2311) <= not(layer2_outputs(7641));
    layer3_outputs(2312) <= not(layer2_outputs(7510));
    layer3_outputs(2313) <= not(layer2_outputs(232));
    layer3_outputs(2314) <= (layer2_outputs(4282)) and not (layer2_outputs(3486));
    layer3_outputs(2315) <= (layer2_outputs(5880)) and (layer2_outputs(7370));
    layer3_outputs(2316) <= not((layer2_outputs(2081)) and (layer2_outputs(2679)));
    layer3_outputs(2317) <= not((layer2_outputs(9)) or (layer2_outputs(3534)));
    layer3_outputs(2318) <= not(layer2_outputs(4614)) or (layer2_outputs(2363));
    layer3_outputs(2319) <= not(layer2_outputs(7552));
    layer3_outputs(2320) <= layer2_outputs(4503);
    layer3_outputs(2321) <= '1';
    layer3_outputs(2322) <= not(layer2_outputs(4263));
    layer3_outputs(2323) <= not(layer2_outputs(6850)) or (layer2_outputs(4475));
    layer3_outputs(2324) <= (layer2_outputs(271)) and not (layer2_outputs(6968));
    layer3_outputs(2325) <= (layer2_outputs(5347)) or (layer2_outputs(1760));
    layer3_outputs(2326) <= not(layer2_outputs(4473));
    layer3_outputs(2327) <= not((layer2_outputs(1840)) or (layer2_outputs(1831)));
    layer3_outputs(2328) <= not(layer2_outputs(3234));
    layer3_outputs(2329) <= (layer2_outputs(3397)) and not (layer2_outputs(2976));
    layer3_outputs(2330) <= '1';
    layer3_outputs(2331) <= not(layer2_outputs(5114));
    layer3_outputs(2332) <= (layer2_outputs(464)) and (layer2_outputs(984));
    layer3_outputs(2333) <= not(layer2_outputs(5944)) or (layer2_outputs(2156));
    layer3_outputs(2334) <= not(layer2_outputs(6394));
    layer3_outputs(2335) <= not(layer2_outputs(3048));
    layer3_outputs(2336) <= not((layer2_outputs(828)) or (layer2_outputs(1038)));
    layer3_outputs(2337) <= layer2_outputs(2343);
    layer3_outputs(2338) <= not(layer2_outputs(1321)) or (layer2_outputs(2061));
    layer3_outputs(2339) <= not(layer2_outputs(5364));
    layer3_outputs(2340) <= not(layer2_outputs(6974));
    layer3_outputs(2341) <= layer2_outputs(3838);
    layer3_outputs(2342) <= layer2_outputs(5612);
    layer3_outputs(2343) <= not(layer2_outputs(5649));
    layer3_outputs(2344) <= '1';
    layer3_outputs(2345) <= not(layer2_outputs(3505));
    layer3_outputs(2346) <= not((layer2_outputs(5662)) xor (layer2_outputs(6489)));
    layer3_outputs(2347) <= layer2_outputs(7191);
    layer3_outputs(2348) <= layer2_outputs(6836);
    layer3_outputs(2349) <= (layer2_outputs(5956)) and not (layer2_outputs(5696));
    layer3_outputs(2350) <= layer2_outputs(1006);
    layer3_outputs(2351) <= '1';
    layer3_outputs(2352) <= layer2_outputs(3797);
    layer3_outputs(2353) <= layer2_outputs(1715);
    layer3_outputs(2354) <= layer2_outputs(3331);
    layer3_outputs(2355) <= layer2_outputs(5765);
    layer3_outputs(2356) <= not((layer2_outputs(3785)) or (layer2_outputs(1059)));
    layer3_outputs(2357) <= '0';
    layer3_outputs(2358) <= not(layer2_outputs(1155));
    layer3_outputs(2359) <= not((layer2_outputs(1188)) and (layer2_outputs(4759)));
    layer3_outputs(2360) <= (layer2_outputs(3996)) and (layer2_outputs(614));
    layer3_outputs(2361) <= (layer2_outputs(6137)) or (layer2_outputs(2540));
    layer3_outputs(2362) <= layer2_outputs(3886);
    layer3_outputs(2363) <= (layer2_outputs(5557)) or (layer2_outputs(5925));
    layer3_outputs(2364) <= (layer2_outputs(3973)) and (layer2_outputs(1036));
    layer3_outputs(2365) <= not((layer2_outputs(4307)) and (layer2_outputs(521)));
    layer3_outputs(2366) <= not(layer2_outputs(4437));
    layer3_outputs(2367) <= not(layer2_outputs(2019)) or (layer2_outputs(3931));
    layer3_outputs(2368) <= '1';
    layer3_outputs(2369) <= layer2_outputs(2895);
    layer3_outputs(2370) <= not((layer2_outputs(7178)) and (layer2_outputs(7138)));
    layer3_outputs(2371) <= not((layer2_outputs(6665)) and (layer2_outputs(5393)));
    layer3_outputs(2372) <= (layer2_outputs(5991)) xor (layer2_outputs(2703));
    layer3_outputs(2373) <= '0';
    layer3_outputs(2374) <= not(layer2_outputs(5613)) or (layer2_outputs(3753));
    layer3_outputs(2375) <= not(layer2_outputs(5659));
    layer3_outputs(2376) <= not(layer2_outputs(706));
    layer3_outputs(2377) <= not(layer2_outputs(5919));
    layer3_outputs(2378) <= '1';
    layer3_outputs(2379) <= not(layer2_outputs(3388));
    layer3_outputs(2380) <= not(layer2_outputs(3607)) or (layer2_outputs(4875));
    layer3_outputs(2381) <= not((layer2_outputs(5302)) xor (layer2_outputs(6899)));
    layer3_outputs(2382) <= (layer2_outputs(6278)) and not (layer2_outputs(5695));
    layer3_outputs(2383) <= not(layer2_outputs(5740)) or (layer2_outputs(2452));
    layer3_outputs(2384) <= (layer2_outputs(2695)) and not (layer2_outputs(5182));
    layer3_outputs(2385) <= not(layer2_outputs(4637)) or (layer2_outputs(1854));
    layer3_outputs(2386) <= not((layer2_outputs(6392)) and (layer2_outputs(4434)));
    layer3_outputs(2387) <= not(layer2_outputs(1086));
    layer3_outputs(2388) <= (layer2_outputs(5257)) and not (layer2_outputs(1091));
    layer3_outputs(2389) <= (layer2_outputs(4240)) or (layer2_outputs(5238));
    layer3_outputs(2390) <= layer2_outputs(381);
    layer3_outputs(2391) <= layer2_outputs(207);
    layer3_outputs(2392) <= (layer2_outputs(7558)) or (layer2_outputs(6667));
    layer3_outputs(2393) <= (layer2_outputs(6430)) xor (layer2_outputs(7632));
    layer3_outputs(2394) <= layer2_outputs(4884);
    layer3_outputs(2395) <= layer2_outputs(813);
    layer3_outputs(2396) <= (layer2_outputs(83)) and not (layer2_outputs(3345));
    layer3_outputs(2397) <= (layer2_outputs(7506)) and not (layer2_outputs(2339));
    layer3_outputs(2398) <= layer2_outputs(1718);
    layer3_outputs(2399) <= not((layer2_outputs(7487)) or (layer2_outputs(4499)));
    layer3_outputs(2400) <= '1';
    layer3_outputs(2401) <= not((layer2_outputs(265)) and (layer2_outputs(5874)));
    layer3_outputs(2402) <= '0';
    layer3_outputs(2403) <= not(layer2_outputs(4054));
    layer3_outputs(2404) <= layer2_outputs(6411);
    layer3_outputs(2405) <= not(layer2_outputs(5020)) or (layer2_outputs(2674));
    layer3_outputs(2406) <= not(layer2_outputs(6953)) or (layer2_outputs(3778));
    layer3_outputs(2407) <= '1';
    layer3_outputs(2408) <= layer2_outputs(4014);
    layer3_outputs(2409) <= '0';
    layer3_outputs(2410) <= '0';
    layer3_outputs(2411) <= not(layer2_outputs(378)) or (layer2_outputs(6597));
    layer3_outputs(2412) <= not((layer2_outputs(4214)) and (layer2_outputs(7610)));
    layer3_outputs(2413) <= (layer2_outputs(7393)) and not (layer2_outputs(7243));
    layer3_outputs(2414) <= (layer2_outputs(6183)) and not (layer2_outputs(654));
    layer3_outputs(2415) <= not((layer2_outputs(2666)) or (layer2_outputs(7030)));
    layer3_outputs(2416) <= not(layer2_outputs(1513)) or (layer2_outputs(4247));
    layer3_outputs(2417) <= '0';
    layer3_outputs(2418) <= (layer2_outputs(557)) or (layer2_outputs(4515));
    layer3_outputs(2419) <= '1';
    layer3_outputs(2420) <= layer2_outputs(3990);
    layer3_outputs(2421) <= layer2_outputs(7410);
    layer3_outputs(2422) <= not(layer2_outputs(5573)) or (layer2_outputs(6888));
    layer3_outputs(2423) <= layer2_outputs(7576);
    layer3_outputs(2424) <= not(layer2_outputs(6368));
    layer3_outputs(2425) <= '0';
    layer3_outputs(2426) <= not(layer2_outputs(2624)) or (layer2_outputs(3832));
    layer3_outputs(2427) <= not((layer2_outputs(141)) or (layer2_outputs(1310)));
    layer3_outputs(2428) <= (layer2_outputs(408)) and (layer2_outputs(6821));
    layer3_outputs(2429) <= (layer2_outputs(2609)) xor (layer2_outputs(224));
    layer3_outputs(2430) <= (layer2_outputs(76)) and (layer2_outputs(1577));
    layer3_outputs(2431) <= not(layer2_outputs(1402));
    layer3_outputs(2432) <= layer2_outputs(4438);
    layer3_outputs(2433) <= not(layer2_outputs(952)) or (layer2_outputs(2789));
    layer3_outputs(2434) <= not(layer2_outputs(4073));
    layer3_outputs(2435) <= not(layer2_outputs(6612)) or (layer2_outputs(3072));
    layer3_outputs(2436) <= '0';
    layer3_outputs(2437) <= (layer2_outputs(1637)) and not (layer2_outputs(3236));
    layer3_outputs(2438) <= layer2_outputs(6454);
    layer3_outputs(2439) <= layer2_outputs(5922);
    layer3_outputs(2440) <= (layer2_outputs(40)) and (layer2_outputs(4521));
    layer3_outputs(2441) <= '1';
    layer3_outputs(2442) <= not(layer2_outputs(5635)) or (layer2_outputs(7480));
    layer3_outputs(2443) <= not(layer2_outputs(5571)) or (layer2_outputs(5262));
    layer3_outputs(2444) <= layer2_outputs(1656);
    layer3_outputs(2445) <= not(layer2_outputs(2119)) or (layer2_outputs(3027));
    layer3_outputs(2446) <= layer2_outputs(5909);
    layer3_outputs(2447) <= (layer2_outputs(1427)) and not (layer2_outputs(4947));
    layer3_outputs(2448) <= layer2_outputs(293);
    layer3_outputs(2449) <= not(layer2_outputs(3940));
    layer3_outputs(2450) <= '1';
    layer3_outputs(2451) <= '0';
    layer3_outputs(2452) <= not(layer2_outputs(7522)) or (layer2_outputs(4197));
    layer3_outputs(2453) <= (layer2_outputs(1294)) and not (layer2_outputs(4400));
    layer3_outputs(2454) <= layer2_outputs(2272);
    layer3_outputs(2455) <= not(layer2_outputs(3123)) or (layer2_outputs(796));
    layer3_outputs(2456) <= layer2_outputs(108);
    layer3_outputs(2457) <= (layer2_outputs(6848)) xor (layer2_outputs(1610));
    layer3_outputs(2458) <= not((layer2_outputs(809)) or (layer2_outputs(621)));
    layer3_outputs(2459) <= not(layer2_outputs(1701));
    layer3_outputs(2460) <= layer2_outputs(7264);
    layer3_outputs(2461) <= not(layer2_outputs(6280));
    layer3_outputs(2462) <= not(layer2_outputs(2330)) or (layer2_outputs(5528));
    layer3_outputs(2463) <= layer2_outputs(6402);
    layer3_outputs(2464) <= layer2_outputs(2151);
    layer3_outputs(2465) <= (layer2_outputs(3510)) or (layer2_outputs(805));
    layer3_outputs(2466) <= (layer2_outputs(3153)) and not (layer2_outputs(1054));
    layer3_outputs(2467) <= not((layer2_outputs(4260)) or (layer2_outputs(7180)));
    layer3_outputs(2468) <= '1';
    layer3_outputs(2469) <= (layer2_outputs(3223)) xor (layer2_outputs(4100));
    layer3_outputs(2470) <= not((layer2_outputs(6357)) and (layer2_outputs(6586)));
    layer3_outputs(2471) <= '0';
    layer3_outputs(2472) <= not((layer2_outputs(1040)) xor (layer2_outputs(479)));
    layer3_outputs(2473) <= (layer2_outputs(4679)) and (layer2_outputs(3210));
    layer3_outputs(2474) <= not((layer2_outputs(1571)) xor (layer2_outputs(6756)));
    layer3_outputs(2475) <= not(layer2_outputs(2830)) or (layer2_outputs(5349));
    layer3_outputs(2476) <= (layer2_outputs(4871)) and (layer2_outputs(947));
    layer3_outputs(2477) <= not((layer2_outputs(1462)) and (layer2_outputs(5963)));
    layer3_outputs(2478) <= not(layer2_outputs(6340));
    layer3_outputs(2479) <= layer2_outputs(203);
    layer3_outputs(2480) <= (layer2_outputs(3632)) or (layer2_outputs(1947));
    layer3_outputs(2481) <= (layer2_outputs(2307)) and (layer2_outputs(1908));
    layer3_outputs(2482) <= (layer2_outputs(4064)) and not (layer2_outputs(1581));
    layer3_outputs(2483) <= '0';
    layer3_outputs(2484) <= layer2_outputs(7200);
    layer3_outputs(2485) <= layer2_outputs(4145);
    layer3_outputs(2486) <= (layer2_outputs(126)) and not (layer2_outputs(1977));
    layer3_outputs(2487) <= '0';
    layer3_outputs(2488) <= not(layer2_outputs(1178));
    layer3_outputs(2489) <= layer2_outputs(6496);
    layer3_outputs(2490) <= not((layer2_outputs(5769)) xor (layer2_outputs(2389)));
    layer3_outputs(2491) <= (layer2_outputs(7149)) xor (layer2_outputs(4729));
    layer3_outputs(2492) <= not((layer2_outputs(4051)) and (layer2_outputs(2964)));
    layer3_outputs(2493) <= not(layer2_outputs(7263));
    layer3_outputs(2494) <= (layer2_outputs(283)) and not (layer2_outputs(977));
    layer3_outputs(2495) <= not((layer2_outputs(5687)) and (layer2_outputs(5249)));
    layer3_outputs(2496) <= (layer2_outputs(7046)) or (layer2_outputs(7314));
    layer3_outputs(2497) <= layer2_outputs(5970);
    layer3_outputs(2498) <= (layer2_outputs(3154)) and not (layer2_outputs(596));
    layer3_outputs(2499) <= layer2_outputs(3993);
    layer3_outputs(2500) <= not(layer2_outputs(6204)) or (layer2_outputs(938));
    layer3_outputs(2501) <= not(layer2_outputs(7318));
    layer3_outputs(2502) <= layer2_outputs(4459);
    layer3_outputs(2503) <= not(layer2_outputs(1682)) or (layer2_outputs(6176));
    layer3_outputs(2504) <= (layer2_outputs(5691)) and (layer2_outputs(596));
    layer3_outputs(2505) <= layer2_outputs(3772);
    layer3_outputs(2506) <= (layer2_outputs(5296)) or (layer2_outputs(5714));
    layer3_outputs(2507) <= (layer2_outputs(4101)) and not (layer2_outputs(4699));
    layer3_outputs(2508) <= '1';
    layer3_outputs(2509) <= not(layer2_outputs(1232));
    layer3_outputs(2510) <= layer2_outputs(6217);
    layer3_outputs(2511) <= '1';
    layer3_outputs(2512) <= not(layer2_outputs(3452));
    layer3_outputs(2513) <= layer2_outputs(6920);
    layer3_outputs(2514) <= not(layer2_outputs(7121)) or (layer2_outputs(4426));
    layer3_outputs(2515) <= not((layer2_outputs(4271)) and (layer2_outputs(2969)));
    layer3_outputs(2516) <= layer2_outputs(1879);
    layer3_outputs(2517) <= '0';
    layer3_outputs(2518) <= (layer2_outputs(4273)) and (layer2_outputs(6299));
    layer3_outputs(2519) <= layer2_outputs(4190);
    layer3_outputs(2520) <= layer2_outputs(3255);
    layer3_outputs(2521) <= (layer2_outputs(4536)) and not (layer2_outputs(6442));
    layer3_outputs(2522) <= (layer2_outputs(6808)) and (layer2_outputs(5470));
    layer3_outputs(2523) <= not((layer2_outputs(5003)) or (layer2_outputs(3325)));
    layer3_outputs(2524) <= not(layer2_outputs(3020));
    layer3_outputs(2525) <= not((layer2_outputs(735)) or (layer2_outputs(2604)));
    layer3_outputs(2526) <= not(layer2_outputs(428)) or (layer2_outputs(7098));
    layer3_outputs(2527) <= layer2_outputs(5673);
    layer3_outputs(2528) <= not(layer2_outputs(2503)) or (layer2_outputs(3128));
    layer3_outputs(2529) <= '1';
    layer3_outputs(2530) <= (layer2_outputs(3685)) and (layer2_outputs(4683));
    layer3_outputs(2531) <= (layer2_outputs(139)) and (layer2_outputs(1423));
    layer3_outputs(2532) <= not(layer2_outputs(6420)) or (layer2_outputs(5526));
    layer3_outputs(2533) <= not(layer2_outputs(5620)) or (layer2_outputs(5322));
    layer3_outputs(2534) <= not(layer2_outputs(4602)) or (layer2_outputs(7269));
    layer3_outputs(2535) <= layer2_outputs(2763);
    layer3_outputs(2536) <= not(layer2_outputs(3351)) or (layer2_outputs(2987));
    layer3_outputs(2537) <= (layer2_outputs(875)) and not (layer2_outputs(5560));
    layer3_outputs(2538) <= '1';
    layer3_outputs(2539) <= not((layer2_outputs(1635)) and (layer2_outputs(2330)));
    layer3_outputs(2540) <= '0';
    layer3_outputs(2541) <= (layer2_outputs(2261)) or (layer2_outputs(5255));
    layer3_outputs(2542) <= not((layer2_outputs(4443)) and (layer2_outputs(4700)));
    layer3_outputs(2543) <= not(layer2_outputs(2825)) or (layer2_outputs(3179));
    layer3_outputs(2544) <= (layer2_outputs(3129)) and (layer2_outputs(6486));
    layer3_outputs(2545) <= (layer2_outputs(3460)) and not (layer2_outputs(6104));
    layer3_outputs(2546) <= layer2_outputs(5158);
    layer3_outputs(2547) <= layer2_outputs(2484);
    layer3_outputs(2548) <= layer2_outputs(3280);
    layer3_outputs(2549) <= not(layer2_outputs(3826)) or (layer2_outputs(7583));
    layer3_outputs(2550) <= layer2_outputs(2593);
    layer3_outputs(2551) <= not(layer2_outputs(3798)) or (layer2_outputs(6414));
    layer3_outputs(2552) <= layer2_outputs(351);
    layer3_outputs(2553) <= (layer2_outputs(1424)) and (layer2_outputs(5058));
    layer3_outputs(2554) <= (layer2_outputs(1474)) or (layer2_outputs(4143));
    layer3_outputs(2555) <= layer2_outputs(7592);
    layer3_outputs(2556) <= not(layer2_outputs(4975)) or (layer2_outputs(3563));
    layer3_outputs(2557) <= not((layer2_outputs(2370)) and (layer2_outputs(7493)));
    layer3_outputs(2558) <= not(layer2_outputs(5613)) or (layer2_outputs(4876));
    layer3_outputs(2559) <= (layer2_outputs(2458)) and not (layer2_outputs(6183));
    layer3_outputs(2560) <= not(layer2_outputs(563));
    layer3_outputs(2561) <= layer2_outputs(5851);
    layer3_outputs(2562) <= layer2_outputs(6146);
    layer3_outputs(2563) <= not(layer2_outputs(7113));
    layer3_outputs(2564) <= not(layer2_outputs(4919));
    layer3_outputs(2565) <= layer2_outputs(3702);
    layer3_outputs(2566) <= (layer2_outputs(4680)) and not (layer2_outputs(3718));
    layer3_outputs(2567) <= not((layer2_outputs(2881)) and (layer2_outputs(312)));
    layer3_outputs(2568) <= (layer2_outputs(7499)) and not (layer2_outputs(4462));
    layer3_outputs(2569) <= not(layer2_outputs(3692));
    layer3_outputs(2570) <= not((layer2_outputs(2452)) or (layer2_outputs(1332)));
    layer3_outputs(2571) <= not(layer2_outputs(3930));
    layer3_outputs(2572) <= (layer2_outputs(3839)) or (layer2_outputs(3833));
    layer3_outputs(2573) <= not(layer2_outputs(1967));
    layer3_outputs(2574) <= not(layer2_outputs(2676)) or (layer2_outputs(7388));
    layer3_outputs(2575) <= '0';
    layer3_outputs(2576) <= not(layer2_outputs(4199));
    layer3_outputs(2577) <= layer2_outputs(7655);
    layer3_outputs(2578) <= layer2_outputs(5517);
    layer3_outputs(2579) <= (layer2_outputs(2153)) and not (layer2_outputs(5285));
    layer3_outputs(2580) <= not((layer2_outputs(2800)) and (layer2_outputs(6362)));
    layer3_outputs(2581) <= not(layer2_outputs(2472));
    layer3_outputs(2582) <= not(layer2_outputs(2797)) or (layer2_outputs(6112));
    layer3_outputs(2583) <= (layer2_outputs(6843)) or (layer2_outputs(3824));
    layer3_outputs(2584) <= layer2_outputs(7407);
    layer3_outputs(2585) <= not(layer2_outputs(6159));
    layer3_outputs(2586) <= '0';
    layer3_outputs(2587) <= layer2_outputs(6558);
    layer3_outputs(2588) <= '1';
    layer3_outputs(2589) <= (layer2_outputs(4169)) or (layer2_outputs(6701));
    layer3_outputs(2590) <= (layer2_outputs(4550)) or (layer2_outputs(425));
    layer3_outputs(2591) <= layer2_outputs(88);
    layer3_outputs(2592) <= not((layer2_outputs(7257)) xor (layer2_outputs(5743)));
    layer3_outputs(2593) <= not(layer2_outputs(2551)) or (layer2_outputs(7509));
    layer3_outputs(2594) <= not(layer2_outputs(4849));
    layer3_outputs(2595) <= not((layer2_outputs(6189)) xor (layer2_outputs(1268)));
    layer3_outputs(2596) <= not(layer2_outputs(6295)) or (layer2_outputs(4061));
    layer3_outputs(2597) <= (layer2_outputs(6471)) and not (layer2_outputs(5480));
    layer3_outputs(2598) <= (layer2_outputs(173)) and not (layer2_outputs(3304));
    layer3_outputs(2599) <= (layer2_outputs(1429)) and (layer2_outputs(7000));
    layer3_outputs(2600) <= not(layer2_outputs(7373));
    layer3_outputs(2601) <= not((layer2_outputs(3875)) or (layer2_outputs(90)));
    layer3_outputs(2602) <= (layer2_outputs(2723)) and (layer2_outputs(5098));
    layer3_outputs(2603) <= not(layer2_outputs(4988));
    layer3_outputs(2604) <= (layer2_outputs(740)) and not (layer2_outputs(5200));
    layer3_outputs(2605) <= layer2_outputs(1359);
    layer3_outputs(2606) <= not(layer2_outputs(3780)) or (layer2_outputs(1325));
    layer3_outputs(2607) <= not(layer2_outputs(1172));
    layer3_outputs(2608) <= layer2_outputs(1305);
    layer3_outputs(2609) <= not(layer2_outputs(1757)) or (layer2_outputs(2872));
    layer3_outputs(2610) <= layer2_outputs(5028);
    layer3_outputs(2611) <= not((layer2_outputs(2883)) or (layer2_outputs(218)));
    layer3_outputs(2612) <= '0';
    layer3_outputs(2613) <= '0';
    layer3_outputs(2614) <= not((layer2_outputs(441)) or (layer2_outputs(6980)));
    layer3_outputs(2615) <= not(layer2_outputs(7004));
    layer3_outputs(2616) <= layer2_outputs(2849);
    layer3_outputs(2617) <= (layer2_outputs(4776)) and (layer2_outputs(3118));
    layer3_outputs(2618) <= '1';
    layer3_outputs(2619) <= layer2_outputs(7443);
    layer3_outputs(2620) <= layer2_outputs(6799);
    layer3_outputs(2621) <= layer2_outputs(1393);
    layer3_outputs(2622) <= not(layer2_outputs(2857)) or (layer2_outputs(3207));
    layer3_outputs(2623) <= layer2_outputs(6001);
    layer3_outputs(2624) <= not(layer2_outputs(1390));
    layer3_outputs(2625) <= not(layer2_outputs(681));
    layer3_outputs(2626) <= not(layer2_outputs(5642)) or (layer2_outputs(5795));
    layer3_outputs(2627) <= not(layer2_outputs(2367));
    layer3_outputs(2628) <= (layer2_outputs(1457)) xor (layer2_outputs(4305));
    layer3_outputs(2629) <= not(layer2_outputs(5615)) or (layer2_outputs(3956));
    layer3_outputs(2630) <= (layer2_outputs(262)) and (layer2_outputs(2679));
    layer3_outputs(2631) <= not(layer2_outputs(7442));
    layer3_outputs(2632) <= not((layer2_outputs(958)) and (layer2_outputs(1902)));
    layer3_outputs(2633) <= '0';
    layer3_outputs(2634) <= not(layer2_outputs(5712));
    layer3_outputs(2635) <= (layer2_outputs(2058)) and not (layer2_outputs(2729));
    layer3_outputs(2636) <= (layer2_outputs(5345)) and (layer2_outputs(6997));
    layer3_outputs(2637) <= not(layer2_outputs(4914));
    layer3_outputs(2638) <= not(layer2_outputs(1467));
    layer3_outputs(2639) <= layer2_outputs(175);
    layer3_outputs(2640) <= not(layer2_outputs(7196));
    layer3_outputs(2641) <= not(layer2_outputs(3599)) or (layer2_outputs(3918));
    layer3_outputs(2642) <= layer2_outputs(7557);
    layer3_outputs(2643) <= (layer2_outputs(1105)) and not (layer2_outputs(3878));
    layer3_outputs(2644) <= '0';
    layer3_outputs(2645) <= layer2_outputs(2896);
    layer3_outputs(2646) <= not((layer2_outputs(1484)) and (layer2_outputs(6016)));
    layer3_outputs(2647) <= '0';
    layer3_outputs(2648) <= not((layer2_outputs(1863)) or (layer2_outputs(3367)));
    layer3_outputs(2649) <= (layer2_outputs(4808)) or (layer2_outputs(1177));
    layer3_outputs(2650) <= (layer2_outputs(4732)) and (layer2_outputs(6482));
    layer3_outputs(2651) <= (layer2_outputs(5206)) and not (layer2_outputs(935));
    layer3_outputs(2652) <= not((layer2_outputs(2217)) xor (layer2_outputs(1146)));
    layer3_outputs(2653) <= layer2_outputs(2451);
    layer3_outputs(2654) <= not((layer2_outputs(584)) and (layer2_outputs(2701)));
    layer3_outputs(2655) <= layer2_outputs(160);
    layer3_outputs(2656) <= not(layer2_outputs(5959));
    layer3_outputs(2657) <= not(layer2_outputs(2237));
    layer3_outputs(2658) <= not(layer2_outputs(4668));
    layer3_outputs(2659) <= layer2_outputs(1942);
    layer3_outputs(2660) <= not(layer2_outputs(2202)) or (layer2_outputs(1103));
    layer3_outputs(2661) <= '0';
    layer3_outputs(2662) <= not(layer2_outputs(3404));
    layer3_outputs(2663) <= layer2_outputs(3419);
    layer3_outputs(2664) <= not(layer2_outputs(2580));
    layer3_outputs(2665) <= (layer2_outputs(7332)) xor (layer2_outputs(5367));
    layer3_outputs(2666) <= (layer2_outputs(7221)) or (layer2_outputs(5168));
    layer3_outputs(2667) <= layer2_outputs(1983);
    layer3_outputs(2668) <= (layer2_outputs(5829)) and not (layer2_outputs(2792));
    layer3_outputs(2669) <= '0';
    layer3_outputs(2670) <= layer2_outputs(2913);
    layer3_outputs(2671) <= '1';
    layer3_outputs(2672) <= layer2_outputs(7434);
    layer3_outputs(2673) <= (layer2_outputs(624)) or (layer2_outputs(2513));
    layer3_outputs(2674) <= (layer2_outputs(3198)) and not (layer2_outputs(5247));
    layer3_outputs(2675) <= '1';
    layer3_outputs(2676) <= (layer2_outputs(5584)) and not (layer2_outputs(2404));
    layer3_outputs(2677) <= not(layer2_outputs(1566));
    layer3_outputs(2678) <= (layer2_outputs(7234)) and not (layer2_outputs(6154));
    layer3_outputs(2679) <= not(layer2_outputs(3065));
    layer3_outputs(2680) <= '0';
    layer3_outputs(2681) <= layer2_outputs(2650);
    layer3_outputs(2682) <= layer2_outputs(3469);
    layer3_outputs(2683) <= not(layer2_outputs(4088)) or (layer2_outputs(1669));
    layer3_outputs(2684) <= not(layer2_outputs(935)) or (layer2_outputs(2133));
    layer3_outputs(2685) <= not(layer2_outputs(1891)) or (layer2_outputs(4278));
    layer3_outputs(2686) <= '1';
    layer3_outputs(2687) <= '1';
    layer3_outputs(2688) <= (layer2_outputs(2095)) or (layer2_outputs(2958));
    layer3_outputs(2689) <= (layer2_outputs(5932)) or (layer2_outputs(3682));
    layer3_outputs(2690) <= layer2_outputs(3807);
    layer3_outputs(2691) <= layer2_outputs(1745);
    layer3_outputs(2692) <= not((layer2_outputs(2878)) and (layer2_outputs(7231)));
    layer3_outputs(2693) <= not(layer2_outputs(2388));
    layer3_outputs(2694) <= layer2_outputs(4358);
    layer3_outputs(2695) <= layer2_outputs(6790);
    layer3_outputs(2696) <= not(layer2_outputs(4385));
    layer3_outputs(2697) <= (layer2_outputs(3777)) or (layer2_outputs(256));
    layer3_outputs(2698) <= not(layer2_outputs(4518));
    layer3_outputs(2699) <= '1';
    layer3_outputs(2700) <= not((layer2_outputs(4991)) xor (layer2_outputs(2464)));
    layer3_outputs(2701) <= not(layer2_outputs(4788));
    layer3_outputs(2702) <= (layer2_outputs(381)) and not (layer2_outputs(3461));
    layer3_outputs(2703) <= not(layer2_outputs(6964));
    layer3_outputs(2704) <= not(layer2_outputs(164));
    layer3_outputs(2705) <= not((layer2_outputs(4707)) and (layer2_outputs(1677)));
    layer3_outputs(2706) <= layer2_outputs(1327);
    layer3_outputs(2707) <= '0';
    layer3_outputs(2708) <= not(layer2_outputs(4931));
    layer3_outputs(2709) <= layer2_outputs(2952);
    layer3_outputs(2710) <= (layer2_outputs(5511)) and not (layer2_outputs(4979));
    layer3_outputs(2711) <= (layer2_outputs(5295)) or (layer2_outputs(1706));
    layer3_outputs(2712) <= not(layer2_outputs(4941)) or (layer2_outputs(3030));
    layer3_outputs(2713) <= (layer2_outputs(3440)) or (layer2_outputs(1857));
    layer3_outputs(2714) <= (layer2_outputs(994)) or (layer2_outputs(3231));
    layer3_outputs(2715) <= (layer2_outputs(27)) xor (layer2_outputs(617));
    layer3_outputs(2716) <= layer2_outputs(6000);
    layer3_outputs(2717) <= (layer2_outputs(6015)) and not (layer2_outputs(3862));
    layer3_outputs(2718) <= not(layer2_outputs(6140)) or (layer2_outputs(1197));
    layer3_outputs(2719) <= layer2_outputs(598);
    layer3_outputs(2720) <= (layer2_outputs(682)) and not (layer2_outputs(4978));
    layer3_outputs(2721) <= layer2_outputs(3659);
    layer3_outputs(2722) <= not((layer2_outputs(2911)) and (layer2_outputs(96)));
    layer3_outputs(2723) <= not((layer2_outputs(6967)) or (layer2_outputs(704)));
    layer3_outputs(2724) <= not((layer2_outputs(4542)) or (layer2_outputs(6371)));
    layer3_outputs(2725) <= not((layer2_outputs(1649)) or (layer2_outputs(3329)));
    layer3_outputs(2726) <= (layer2_outputs(6644)) xor (layer2_outputs(4626));
    layer3_outputs(2727) <= not(layer2_outputs(1392));
    layer3_outputs(2728) <= '0';
    layer3_outputs(2729) <= not((layer2_outputs(7265)) and (layer2_outputs(5435)));
    layer3_outputs(2730) <= not(layer2_outputs(6180));
    layer3_outputs(2731) <= layer2_outputs(4076);
    layer3_outputs(2732) <= not(layer2_outputs(1849));
    layer3_outputs(2733) <= (layer2_outputs(5884)) and not (layer2_outputs(939));
    layer3_outputs(2734) <= (layer2_outputs(3725)) or (layer2_outputs(6751));
    layer3_outputs(2735) <= not(layer2_outputs(2141));
    layer3_outputs(2736) <= layer2_outputs(190);
    layer3_outputs(2737) <= (layer2_outputs(1336)) and not (layer2_outputs(1957));
    layer3_outputs(2738) <= not(layer2_outputs(3537)) or (layer2_outputs(1506));
    layer3_outputs(2739) <= (layer2_outputs(1468)) and not (layer2_outputs(6016));
    layer3_outputs(2740) <= (layer2_outputs(4089)) and not (layer2_outputs(3085));
    layer3_outputs(2741) <= not(layer2_outputs(6789));
    layer3_outputs(2742) <= not(layer2_outputs(3975));
    layer3_outputs(2743) <= not((layer2_outputs(4380)) and (layer2_outputs(1179)));
    layer3_outputs(2744) <= (layer2_outputs(7045)) and not (layer2_outputs(118));
    layer3_outputs(2745) <= not(layer2_outputs(4751));
    layer3_outputs(2746) <= layer2_outputs(278);
    layer3_outputs(2747) <= not((layer2_outputs(6492)) xor (layer2_outputs(6202)));
    layer3_outputs(2748) <= layer2_outputs(2421);
    layer3_outputs(2749) <= '0';
    layer3_outputs(2750) <= not(layer2_outputs(6429));
    layer3_outputs(2751) <= not((layer2_outputs(6913)) or (layer2_outputs(382)));
    layer3_outputs(2752) <= layer2_outputs(1124);
    layer3_outputs(2753) <= layer2_outputs(4468);
    layer3_outputs(2754) <= not(layer2_outputs(6512));
    layer3_outputs(2755) <= (layer2_outputs(1349)) and (layer2_outputs(2289));
    layer3_outputs(2756) <= layer2_outputs(1607);
    layer3_outputs(2757) <= layer2_outputs(3909);
    layer3_outputs(2758) <= not(layer2_outputs(972)) or (layer2_outputs(2089));
    layer3_outputs(2759) <= not(layer2_outputs(5655));
    layer3_outputs(2760) <= '0';
    layer3_outputs(2761) <= (layer2_outputs(1843)) and not (layer2_outputs(5798));
    layer3_outputs(2762) <= not(layer2_outputs(7304)) or (layer2_outputs(1187));
    layer3_outputs(2763) <= not((layer2_outputs(376)) and (layer2_outputs(622)));
    layer3_outputs(2764) <= not(layer2_outputs(924));
    layer3_outputs(2765) <= '1';
    layer3_outputs(2766) <= layer2_outputs(6396);
    layer3_outputs(2767) <= (layer2_outputs(7123)) and (layer2_outputs(2085));
    layer3_outputs(2768) <= not((layer2_outputs(1164)) and (layer2_outputs(6441)));
    layer3_outputs(2769) <= (layer2_outputs(3497)) or (layer2_outputs(5799));
    layer3_outputs(2770) <= layer2_outputs(2011);
    layer3_outputs(2771) <= layer2_outputs(3801);
    layer3_outputs(2772) <= (layer2_outputs(537)) and not (layer2_outputs(6119));
    layer3_outputs(2773) <= '1';
    layer3_outputs(2774) <= not(layer2_outputs(1355));
    layer3_outputs(2775) <= not((layer2_outputs(2739)) or (layer2_outputs(6179)));
    layer3_outputs(2776) <= not(layer2_outputs(3162)) or (layer2_outputs(5246));
    layer3_outputs(2777) <= (layer2_outputs(2161)) and not (layer2_outputs(6053));
    layer3_outputs(2778) <= not(layer2_outputs(4924));
    layer3_outputs(2779) <= not(layer2_outputs(4361));
    layer3_outputs(2780) <= '1';
    layer3_outputs(2781) <= '0';
    layer3_outputs(2782) <= layer2_outputs(3379);
    layer3_outputs(2783) <= layer2_outputs(5081);
    layer3_outputs(2784) <= (layer2_outputs(4981)) and (layer2_outputs(7647));
    layer3_outputs(2785) <= (layer2_outputs(5447)) and not (layer2_outputs(5294));
    layer3_outputs(2786) <= layer2_outputs(1852);
    layer3_outputs(2787) <= (layer2_outputs(1185)) and (layer2_outputs(1696));
    layer3_outputs(2788) <= (layer2_outputs(1011)) and not (layer2_outputs(3085));
    layer3_outputs(2789) <= '0';
    layer3_outputs(2790) <= layer2_outputs(2552);
    layer3_outputs(2791) <= (layer2_outputs(708)) and not (layer2_outputs(4658));
    layer3_outputs(2792) <= not((layer2_outputs(3534)) and (layer2_outputs(4161)));
    layer3_outputs(2793) <= layer2_outputs(2031);
    layer3_outputs(2794) <= layer2_outputs(4179);
    layer3_outputs(2795) <= not((layer2_outputs(964)) and (layer2_outputs(1229)));
    layer3_outputs(2796) <= not((layer2_outputs(6260)) and (layer2_outputs(7397)));
    layer3_outputs(2797) <= (layer2_outputs(7538)) and (layer2_outputs(6332));
    layer3_outputs(2798) <= not(layer2_outputs(3174)) or (layer2_outputs(3372));
    layer3_outputs(2799) <= '1';
    layer3_outputs(2800) <= (layer2_outputs(1168)) and not (layer2_outputs(397));
    layer3_outputs(2801) <= not(layer2_outputs(7203));
    layer3_outputs(2802) <= not(layer2_outputs(6064));
    layer3_outputs(2803) <= not(layer2_outputs(7575)) or (layer2_outputs(1880));
    layer3_outputs(2804) <= not(layer2_outputs(7495)) or (layer2_outputs(4292));
    layer3_outputs(2805) <= not((layer2_outputs(1759)) or (layer2_outputs(6210)));
    layer3_outputs(2806) <= not(layer2_outputs(1066)) or (layer2_outputs(1327));
    layer3_outputs(2807) <= layer2_outputs(6630);
    layer3_outputs(2808) <= not(layer2_outputs(5259));
    layer3_outputs(2809) <= layer2_outputs(4031);
    layer3_outputs(2810) <= (layer2_outputs(2783)) and (layer2_outputs(4940));
    layer3_outputs(2811) <= (layer2_outputs(4956)) xor (layer2_outputs(3106));
    layer3_outputs(2812) <= (layer2_outputs(3964)) and not (layer2_outputs(2874));
    layer3_outputs(2813) <= layer2_outputs(7135);
    layer3_outputs(2814) <= not(layer2_outputs(4954));
    layer3_outputs(2815) <= '0';
    layer3_outputs(2816) <= not(layer2_outputs(852));
    layer3_outputs(2817) <= (layer2_outputs(3122)) and not (layer2_outputs(3715));
    layer3_outputs(2818) <= (layer2_outputs(389)) and not (layer2_outputs(6796));
    layer3_outputs(2819) <= (layer2_outputs(2243)) and not (layer2_outputs(4244));
    layer3_outputs(2820) <= (layer2_outputs(925)) and (layer2_outputs(4526));
    layer3_outputs(2821) <= '1';
    layer3_outputs(2822) <= (layer2_outputs(2332)) and not (layer2_outputs(104));
    layer3_outputs(2823) <= not(layer2_outputs(7131)) or (layer2_outputs(4658));
    layer3_outputs(2824) <= layer2_outputs(965);
    layer3_outputs(2825) <= layer2_outputs(5822);
    layer3_outputs(2826) <= '0';
    layer3_outputs(2827) <= not(layer2_outputs(1684));
    layer3_outputs(2828) <= not((layer2_outputs(2945)) or (layer2_outputs(6387)));
    layer3_outputs(2829) <= (layer2_outputs(5652)) or (layer2_outputs(7113));
    layer3_outputs(2830) <= not(layer2_outputs(6238));
    layer3_outputs(2831) <= '1';
    layer3_outputs(2832) <= not(layer2_outputs(3337)) or (layer2_outputs(286));
    layer3_outputs(2833) <= not((layer2_outputs(7212)) or (layer2_outputs(5728)));
    layer3_outputs(2834) <= (layer2_outputs(4246)) and not (layer2_outputs(778));
    layer3_outputs(2835) <= '1';
    layer3_outputs(2836) <= (layer2_outputs(841)) and not (layer2_outputs(5572));
    layer3_outputs(2837) <= (layer2_outputs(3911)) or (layer2_outputs(6518));
    layer3_outputs(2838) <= layer2_outputs(2497);
    layer3_outputs(2839) <= not((layer2_outputs(1797)) or (layer2_outputs(2595)));
    layer3_outputs(2840) <= not((layer2_outputs(4347)) xor (layer2_outputs(338)));
    layer3_outputs(2841) <= (layer2_outputs(3074)) xor (layer2_outputs(5778));
    layer3_outputs(2842) <= not(layer2_outputs(2846));
    layer3_outputs(2843) <= not((layer2_outputs(5914)) and (layer2_outputs(5024)));
    layer3_outputs(2844) <= not(layer2_outputs(3095)) or (layer2_outputs(5303));
    layer3_outputs(2845) <= not(layer2_outputs(4364)) or (layer2_outputs(5366));
    layer3_outputs(2846) <= layer2_outputs(630);
    layer3_outputs(2847) <= not(layer2_outputs(3588));
    layer3_outputs(2848) <= not(layer2_outputs(6364));
    layer3_outputs(2849) <= layer2_outputs(6275);
    layer3_outputs(2850) <= layer2_outputs(6861);
    layer3_outputs(2851) <= (layer2_outputs(5858)) and not (layer2_outputs(1495));
    layer3_outputs(2852) <= (layer2_outputs(197)) or (layer2_outputs(6682));
    layer3_outputs(2853) <= layer2_outputs(2655);
    layer3_outputs(2854) <= '1';
    layer3_outputs(2855) <= not(layer2_outputs(2097)) or (layer2_outputs(2090));
    layer3_outputs(2856) <= not(layer2_outputs(3681)) or (layer2_outputs(419));
    layer3_outputs(2857) <= not((layer2_outputs(3013)) or (layer2_outputs(6853)));
    layer3_outputs(2858) <= not((layer2_outputs(2166)) xor (layer2_outputs(353)));
    layer3_outputs(2859) <= not((layer2_outputs(4300)) and (layer2_outputs(61)));
    layer3_outputs(2860) <= not((layer2_outputs(6365)) or (layer2_outputs(2766)));
    layer3_outputs(2861) <= layer2_outputs(1189);
    layer3_outputs(2862) <= not(layer2_outputs(3012)) or (layer2_outputs(91));
    layer3_outputs(2863) <= layer2_outputs(1606);
    layer3_outputs(2864) <= not((layer2_outputs(2336)) and (layer2_outputs(7219)));
    layer3_outputs(2865) <= not(layer2_outputs(3744)) or (layer2_outputs(485));
    layer3_outputs(2866) <= '1';
    layer3_outputs(2867) <= not((layer2_outputs(2189)) or (layer2_outputs(2479)));
    layer3_outputs(2868) <= not(layer2_outputs(726));
    layer3_outputs(2869) <= layer2_outputs(1601);
    layer3_outputs(2870) <= not(layer2_outputs(517)) or (layer2_outputs(2833));
    layer3_outputs(2871) <= not(layer2_outputs(5298));
    layer3_outputs(2872) <= not(layer2_outputs(3436));
    layer3_outputs(2873) <= (layer2_outputs(2147)) and (layer2_outputs(5519));
    layer3_outputs(2874) <= layer2_outputs(3056);
    layer3_outputs(2875) <= '0';
    layer3_outputs(2876) <= (layer2_outputs(7503)) and not (layer2_outputs(1897));
    layer3_outputs(2877) <= (layer2_outputs(5859)) and (layer2_outputs(1525));
    layer3_outputs(2878) <= not(layer2_outputs(4240));
    layer3_outputs(2879) <= not(layer2_outputs(3740));
    layer3_outputs(2880) <= (layer2_outputs(1868)) and not (layer2_outputs(6342));
    layer3_outputs(2881) <= layer2_outputs(7003);
    layer3_outputs(2882) <= not(layer2_outputs(6706)) or (layer2_outputs(4091));
    layer3_outputs(2883) <= layer2_outputs(3130);
    layer3_outputs(2884) <= not(layer2_outputs(3342));
    layer3_outputs(2885) <= not(layer2_outputs(4332));
    layer3_outputs(2886) <= not(layer2_outputs(4714));
    layer3_outputs(2887) <= not(layer2_outputs(7604));
    layer3_outputs(2888) <= (layer2_outputs(3319)) and not (layer2_outputs(5276));
    layer3_outputs(2889) <= not(layer2_outputs(6149)) or (layer2_outputs(6600));
    layer3_outputs(2890) <= '0';
    layer3_outputs(2891) <= not(layer2_outputs(1033)) or (layer2_outputs(6945));
    layer3_outputs(2892) <= not(layer2_outputs(4568));
    layer3_outputs(2893) <= '1';
    layer3_outputs(2894) <= '1';
    layer3_outputs(2895) <= not(layer2_outputs(929));
    layer3_outputs(2896) <= (layer2_outputs(6887)) and not (layer2_outputs(1702));
    layer3_outputs(2897) <= layer2_outputs(685);
    layer3_outputs(2898) <= layer2_outputs(4105);
    layer3_outputs(2899) <= not(layer2_outputs(170)) or (layer2_outputs(7307));
    layer3_outputs(2900) <= not(layer2_outputs(3423)) or (layer2_outputs(4183));
    layer3_outputs(2901) <= layer2_outputs(4377);
    layer3_outputs(2902) <= layer2_outputs(6879);
    layer3_outputs(2903) <= layer2_outputs(4451);
    layer3_outputs(2904) <= (layer2_outputs(4863)) or (layer2_outputs(6721));
    layer3_outputs(2905) <= layer2_outputs(5589);
    layer3_outputs(2906) <= '1';
    layer3_outputs(2907) <= not(layer2_outputs(4821)) or (layer2_outputs(2425));
    layer3_outputs(2908) <= '1';
    layer3_outputs(2909) <= (layer2_outputs(5491)) or (layer2_outputs(7370));
    layer3_outputs(2910) <= (layer2_outputs(2828)) and not (layer2_outputs(7566));
    layer3_outputs(2911) <= not((layer2_outputs(5051)) and (layer2_outputs(2077)));
    layer3_outputs(2912) <= (layer2_outputs(1079)) and not (layer2_outputs(2914));
    layer3_outputs(2913) <= (layer2_outputs(5265)) and (layer2_outputs(3026));
    layer3_outputs(2914) <= (layer2_outputs(7084)) or (layer2_outputs(2416));
    layer3_outputs(2915) <= not((layer2_outputs(5488)) or (layer2_outputs(5989)));
    layer3_outputs(2916) <= (layer2_outputs(593)) and (layer2_outputs(257));
    layer3_outputs(2917) <= not((layer2_outputs(5473)) or (layer2_outputs(2341)));
    layer3_outputs(2918) <= not(layer2_outputs(3059));
    layer3_outputs(2919) <= (layer2_outputs(334)) and not (layer2_outputs(485));
    layer3_outputs(2920) <= layer2_outputs(5714);
    layer3_outputs(2921) <= (layer2_outputs(4448)) or (layer2_outputs(2042));
    layer3_outputs(2922) <= not(layer2_outputs(7618));
    layer3_outputs(2923) <= layer2_outputs(240);
    layer3_outputs(2924) <= (layer2_outputs(4782)) and not (layer2_outputs(5612));
    layer3_outputs(2925) <= (layer2_outputs(1080)) and (layer2_outputs(477));
    layer3_outputs(2926) <= not((layer2_outputs(1241)) xor (layer2_outputs(4460)));
    layer3_outputs(2927) <= not((layer2_outputs(3821)) or (layer2_outputs(224)));
    layer3_outputs(2928) <= not((layer2_outputs(5221)) and (layer2_outputs(2150)));
    layer3_outputs(2929) <= not(layer2_outputs(2154));
    layer3_outputs(2930) <= layer2_outputs(6967);
    layer3_outputs(2931) <= not(layer2_outputs(2368));
    layer3_outputs(2932) <= not(layer2_outputs(6315));
    layer3_outputs(2933) <= (layer2_outputs(1618)) and not (layer2_outputs(1182));
    layer3_outputs(2934) <= (layer2_outputs(7030)) and (layer2_outputs(7193));
    layer3_outputs(2935) <= not(layer2_outputs(4933)) or (layer2_outputs(4541));
    layer3_outputs(2936) <= not(layer2_outputs(603)) or (layer2_outputs(3375));
    layer3_outputs(2937) <= (layer2_outputs(1307)) and not (layer2_outputs(3840));
    layer3_outputs(2938) <= (layer2_outputs(4412)) and not (layer2_outputs(3312));
    layer3_outputs(2939) <= not((layer2_outputs(452)) and (layer2_outputs(7308)));
    layer3_outputs(2940) <= not(layer2_outputs(5458)) or (layer2_outputs(3170));
    layer3_outputs(2941) <= '0';
    layer3_outputs(2942) <= not(layer2_outputs(1911));
    layer3_outputs(2943) <= (layer2_outputs(874)) and not (layer2_outputs(1324));
    layer3_outputs(2944) <= not((layer2_outputs(6174)) or (layer2_outputs(4908)));
    layer3_outputs(2945) <= (layer2_outputs(6865)) and not (layer2_outputs(1888));
    layer3_outputs(2946) <= layer2_outputs(7013);
    layer3_outputs(2947) <= not(layer2_outputs(7081)) or (layer2_outputs(4330));
    layer3_outputs(2948) <= not(layer2_outputs(4430));
    layer3_outputs(2949) <= '0';
    layer3_outputs(2950) <= '1';
    layer3_outputs(2951) <= (layer2_outputs(5671)) and not (layer2_outputs(1648));
    layer3_outputs(2952) <= '1';
    layer3_outputs(2953) <= not((layer2_outputs(5885)) and (layer2_outputs(3603)));
    layer3_outputs(2954) <= not(layer2_outputs(2760)) or (layer2_outputs(6));
    layer3_outputs(2955) <= '0';
    layer3_outputs(2956) <= not(layer2_outputs(49));
    layer3_outputs(2957) <= not((layer2_outputs(7678)) and (layer2_outputs(3642)));
    layer3_outputs(2958) <= not((layer2_outputs(6361)) and (layer2_outputs(4626)));
    layer3_outputs(2959) <= layer2_outputs(1135);
    layer3_outputs(2960) <= (layer2_outputs(3506)) and not (layer2_outputs(7587));
    layer3_outputs(2961) <= not(layer2_outputs(999)) or (layer2_outputs(7324));
    layer3_outputs(2962) <= not(layer2_outputs(4140)) or (layer2_outputs(1100));
    layer3_outputs(2963) <= not(layer2_outputs(7018));
    layer3_outputs(2964) <= (layer2_outputs(697)) and (layer2_outputs(5962));
    layer3_outputs(2965) <= layer2_outputs(2439);
    layer3_outputs(2966) <= (layer2_outputs(5563)) and not (layer2_outputs(7060));
    layer3_outputs(2967) <= not(layer2_outputs(3325));
    layer3_outputs(2968) <= (layer2_outputs(5872)) and (layer2_outputs(5120));
    layer3_outputs(2969) <= (layer2_outputs(7526)) or (layer2_outputs(657));
    layer3_outputs(2970) <= layer2_outputs(6545);
    layer3_outputs(2971) <= not(layer2_outputs(106));
    layer3_outputs(2972) <= layer2_outputs(3841);
    layer3_outputs(2973) <= layer2_outputs(6279);
    layer3_outputs(2974) <= layer2_outputs(3296);
    layer3_outputs(2975) <= (layer2_outputs(7237)) xor (layer2_outputs(5632));
    layer3_outputs(2976) <= not(layer2_outputs(1678)) or (layer2_outputs(5371));
    layer3_outputs(2977) <= (layer2_outputs(698)) or (layer2_outputs(7634));
    layer3_outputs(2978) <= not((layer2_outputs(2700)) and (layer2_outputs(1657)));
    layer3_outputs(2979) <= (layer2_outputs(6788)) or (layer2_outputs(6845));
    layer3_outputs(2980) <= layer2_outputs(4284);
    layer3_outputs(2981) <= '1';
    layer3_outputs(2982) <= '0';
    layer3_outputs(2983) <= not(layer2_outputs(3711));
    layer3_outputs(2984) <= not(layer2_outputs(3927)) or (layer2_outputs(2082));
    layer3_outputs(2985) <= layer2_outputs(186);
    layer3_outputs(2986) <= not(layer2_outputs(407));
    layer3_outputs(2987) <= not(layer2_outputs(1060));
    layer3_outputs(2988) <= not(layer2_outputs(6167)) or (layer2_outputs(3720));
    layer3_outputs(2989) <= (layer2_outputs(4101)) and not (layer2_outputs(7467));
    layer3_outputs(2990) <= not(layer2_outputs(3541));
    layer3_outputs(2991) <= (layer2_outputs(2027)) and not (layer2_outputs(7485));
    layer3_outputs(2992) <= (layer2_outputs(173)) and (layer2_outputs(5460));
    layer3_outputs(2993) <= not(layer2_outputs(3727));
    layer3_outputs(2994) <= (layer2_outputs(1794)) and (layer2_outputs(85));
    layer3_outputs(2995) <= not((layer2_outputs(5097)) xor (layer2_outputs(1192)));
    layer3_outputs(2996) <= not(layer2_outputs(7454));
    layer3_outputs(2997) <= (layer2_outputs(7340)) xor (layer2_outputs(2955));
    layer3_outputs(2998) <= not((layer2_outputs(7088)) or (layer2_outputs(6461)));
    layer3_outputs(2999) <= not(layer2_outputs(5538)) or (layer2_outputs(4221));
    layer3_outputs(3000) <= not(layer2_outputs(5063)) or (layer2_outputs(2753));
    layer3_outputs(3001) <= not((layer2_outputs(7183)) or (layer2_outputs(7518)));
    layer3_outputs(3002) <= not((layer2_outputs(484)) or (layer2_outputs(2507)));
    layer3_outputs(3003) <= layer2_outputs(928);
    layer3_outputs(3004) <= layer2_outputs(5794);
    layer3_outputs(3005) <= not((layer2_outputs(1939)) and (layer2_outputs(4389)));
    layer3_outputs(3006) <= not(layer2_outputs(3553));
    layer3_outputs(3007) <= not(layer2_outputs(7443));
    layer3_outputs(3008) <= '0';
    layer3_outputs(3009) <= not((layer2_outputs(6675)) and (layer2_outputs(455)));
    layer3_outputs(3010) <= not(layer2_outputs(3909));
    layer3_outputs(3011) <= not(layer2_outputs(3987));
    layer3_outputs(3012) <= layer2_outputs(7516);
    layer3_outputs(3013) <= (layer2_outputs(6269)) and not (layer2_outputs(5442));
    layer3_outputs(3014) <= (layer2_outputs(3278)) and (layer2_outputs(2157));
    layer3_outputs(3015) <= not((layer2_outputs(2223)) or (layer2_outputs(2901)));
    layer3_outputs(3016) <= not(layer2_outputs(5736)) or (layer2_outputs(4881));
    layer3_outputs(3017) <= not(layer2_outputs(4962));
    layer3_outputs(3018) <= not(layer2_outputs(1098));
    layer3_outputs(3019) <= '0';
    layer3_outputs(3020) <= not(layer2_outputs(288));
    layer3_outputs(3021) <= layer2_outputs(4910);
    layer3_outputs(3022) <= not(layer2_outputs(3545)) or (layer2_outputs(7671));
    layer3_outputs(3023) <= layer2_outputs(3474);
    layer3_outputs(3024) <= not(layer2_outputs(3943));
    layer3_outputs(3025) <= not(layer2_outputs(5210));
    layer3_outputs(3026) <= not(layer2_outputs(6633)) or (layer2_outputs(425));
    layer3_outputs(3027) <= (layer2_outputs(2136)) and (layer2_outputs(1777));
    layer3_outputs(3028) <= layer2_outputs(5761);
    layer3_outputs(3029) <= not(layer2_outputs(6737));
    layer3_outputs(3030) <= (layer2_outputs(216)) or (layer2_outputs(3617));
    layer3_outputs(3031) <= '0';
    layer3_outputs(3032) <= not((layer2_outputs(1452)) and (layer2_outputs(474)));
    layer3_outputs(3033) <= (layer2_outputs(2647)) xor (layer2_outputs(3062));
    layer3_outputs(3034) <= not(layer2_outputs(3795)) or (layer2_outputs(7152));
    layer3_outputs(3035) <= not(layer2_outputs(1018));
    layer3_outputs(3036) <= not((layer2_outputs(1379)) and (layer2_outputs(3593)));
    layer3_outputs(3037) <= (layer2_outputs(296)) and not (layer2_outputs(1755));
    layer3_outputs(3038) <= not(layer2_outputs(315));
    layer3_outputs(3039) <= not(layer2_outputs(3441));
    layer3_outputs(3040) <= (layer2_outputs(3676)) and (layer2_outputs(346));
    layer3_outputs(3041) <= (layer2_outputs(3151)) and not (layer2_outputs(6468));
    layer3_outputs(3042) <= not((layer2_outputs(2775)) and (layer2_outputs(2726)));
    layer3_outputs(3043) <= not((layer2_outputs(758)) or (layer2_outputs(5535)));
    layer3_outputs(3044) <= (layer2_outputs(3036)) and (layer2_outputs(7168));
    layer3_outputs(3045) <= (layer2_outputs(2533)) or (layer2_outputs(3493));
    layer3_outputs(3046) <= not(layer2_outputs(7233));
    layer3_outputs(3047) <= not((layer2_outputs(2984)) or (layer2_outputs(4682)));
    layer3_outputs(3048) <= not(layer2_outputs(7507)) or (layer2_outputs(317));
    layer3_outputs(3049) <= not((layer2_outputs(2408)) or (layer2_outputs(1227)));
    layer3_outputs(3050) <= not(layer2_outputs(1526));
    layer3_outputs(3051) <= (layer2_outputs(4098)) and (layer2_outputs(2999));
    layer3_outputs(3052) <= '0';
    layer3_outputs(3053) <= '1';
    layer3_outputs(3054) <= not(layer2_outputs(6582));
    layer3_outputs(3055) <= not(layer2_outputs(507));
    layer3_outputs(3056) <= not(layer2_outputs(5243));
    layer3_outputs(3057) <= layer2_outputs(2385);
    layer3_outputs(3058) <= not(layer2_outputs(2123)) or (layer2_outputs(5472));
    layer3_outputs(3059) <= (layer2_outputs(2911)) and (layer2_outputs(787));
    layer3_outputs(3060) <= (layer2_outputs(1272)) or (layer2_outputs(5980));
    layer3_outputs(3061) <= not(layer2_outputs(2910));
    layer3_outputs(3062) <= (layer2_outputs(7270)) or (layer2_outputs(1882));
    layer3_outputs(3063) <= '0';
    layer3_outputs(3064) <= layer2_outputs(204);
    layer3_outputs(3065) <= layer2_outputs(5284);
    layer3_outputs(3066) <= not((layer2_outputs(332)) or (layer2_outputs(3932)));
    layer3_outputs(3067) <= '1';
    layer3_outputs(3068) <= layer2_outputs(1188);
    layer3_outputs(3069) <= layer2_outputs(3884);
    layer3_outputs(3070) <= '0';
    layer3_outputs(3071) <= (layer2_outputs(646)) and (layer2_outputs(6627));
    layer3_outputs(3072) <= not((layer2_outputs(4831)) or (layer2_outputs(3712)));
    layer3_outputs(3073) <= not(layer2_outputs(3636));
    layer3_outputs(3074) <= not(layer2_outputs(3429));
    layer3_outputs(3075) <= not(layer2_outputs(78)) or (layer2_outputs(631));
    layer3_outputs(3076) <= (layer2_outputs(5376)) and not (layer2_outputs(4769));
    layer3_outputs(3077) <= not(layer2_outputs(5689));
    layer3_outputs(3078) <= (layer2_outputs(1577)) xor (layer2_outputs(4853));
    layer3_outputs(3079) <= not((layer2_outputs(2830)) and (layer2_outputs(4874)));
    layer3_outputs(3080) <= (layer2_outputs(782)) and not (layer2_outputs(801));
    layer3_outputs(3081) <= (layer2_outputs(5272)) or (layer2_outputs(4080));
    layer3_outputs(3082) <= (layer2_outputs(5900)) xor (layer2_outputs(5279));
    layer3_outputs(3083) <= (layer2_outputs(4508)) or (layer2_outputs(6556));
    layer3_outputs(3084) <= not(layer2_outputs(7377));
    layer3_outputs(3085) <= '0';
    layer3_outputs(3086) <= not((layer2_outputs(211)) or (layer2_outputs(1534)));
    layer3_outputs(3087) <= not((layer2_outputs(2127)) or (layer2_outputs(6664)));
    layer3_outputs(3088) <= '1';
    layer3_outputs(3089) <= '0';
    layer3_outputs(3090) <= '1';
    layer3_outputs(3091) <= not((layer2_outputs(1672)) xor (layer2_outputs(5901)));
    layer3_outputs(3092) <= not(layer2_outputs(1711)) or (layer2_outputs(1238));
    layer3_outputs(3093) <= (layer2_outputs(1124)) and not (layer2_outputs(7146));
    layer3_outputs(3094) <= not(layer2_outputs(476));
    layer3_outputs(3095) <= not(layer2_outputs(1139)) or (layer2_outputs(7028));
    layer3_outputs(3096) <= not(layer2_outputs(7191));
    layer3_outputs(3097) <= '0';
    layer3_outputs(3098) <= layer2_outputs(600);
    layer3_outputs(3099) <= (layer2_outputs(3393)) and (layer2_outputs(7306));
    layer3_outputs(3100) <= (layer2_outputs(5607)) and not (layer2_outputs(6544));
    layer3_outputs(3101) <= not((layer2_outputs(5507)) and (layer2_outputs(2822)));
    layer3_outputs(3102) <= not(layer2_outputs(3540)) or (layer2_outputs(7517));
    layer3_outputs(3103) <= not((layer2_outputs(2328)) and (layer2_outputs(1446)));
    layer3_outputs(3104) <= (layer2_outputs(6418)) xor (layer2_outputs(3904));
    layer3_outputs(3105) <= (layer2_outputs(3672)) and (layer2_outputs(5941));
    layer3_outputs(3106) <= (layer2_outputs(2725)) or (layer2_outputs(1061));
    layer3_outputs(3107) <= not((layer2_outputs(2123)) and (layer2_outputs(1841)));
    layer3_outputs(3108) <= layer2_outputs(7058);
    layer3_outputs(3109) <= not((layer2_outputs(3476)) and (layer2_outputs(304)));
    layer3_outputs(3110) <= not(layer2_outputs(6421)) or (layer2_outputs(4319));
    layer3_outputs(3111) <= (layer2_outputs(7104)) or (layer2_outputs(1564));
    layer3_outputs(3112) <= layer2_outputs(7342);
    layer3_outputs(3113) <= layer2_outputs(6206);
    layer3_outputs(3114) <= not(layer2_outputs(2019));
    layer3_outputs(3115) <= (layer2_outputs(2251)) and not (layer2_outputs(1487));
    layer3_outputs(3116) <= (layer2_outputs(6284)) or (layer2_outputs(6753));
    layer3_outputs(3117) <= not(layer2_outputs(3967));
    layer3_outputs(3118) <= (layer2_outputs(6113)) or (layer2_outputs(5174));
    layer3_outputs(3119) <= (layer2_outputs(5648)) and (layer2_outputs(7296));
    layer3_outputs(3120) <= (layer2_outputs(4880)) and (layer2_outputs(5924));
    layer3_outputs(3121) <= layer2_outputs(6404);
    layer3_outputs(3122) <= layer2_outputs(1407);
    layer3_outputs(3123) <= layer2_outputs(3134);
    layer3_outputs(3124) <= (layer2_outputs(3372)) or (layer2_outputs(7120));
    layer3_outputs(3125) <= '0';
    layer3_outputs(3126) <= layer2_outputs(3452);
    layer3_outputs(3127) <= not(layer2_outputs(2931)) or (layer2_outputs(2847));
    layer3_outputs(3128) <= not(layer2_outputs(634));
    layer3_outputs(3129) <= (layer2_outputs(6252)) or (layer2_outputs(4591));
    layer3_outputs(3130) <= '0';
    layer3_outputs(3131) <= layer2_outputs(4201);
    layer3_outputs(3132) <= not(layer2_outputs(594)) or (layer2_outputs(6759));
    layer3_outputs(3133) <= layer2_outputs(5828);
    layer3_outputs(3134) <= not(layer2_outputs(1789));
    layer3_outputs(3135) <= (layer2_outputs(744)) and not (layer2_outputs(1596));
    layer3_outputs(3136) <= not(layer2_outputs(5109));
    layer3_outputs(3137) <= layer2_outputs(1324);
    layer3_outputs(3138) <= not(layer2_outputs(3157));
    layer3_outputs(3139) <= not(layer2_outputs(3373));
    layer3_outputs(3140) <= (layer2_outputs(5080)) and not (layer2_outputs(2790));
    layer3_outputs(3141) <= not(layer2_outputs(4775));
    layer3_outputs(3142) <= not(layer2_outputs(6806));
    layer3_outputs(3143) <= not(layer2_outputs(6504));
    layer3_outputs(3144) <= (layer2_outputs(5556)) and not (layer2_outputs(7653));
    layer3_outputs(3145) <= '0';
    layer3_outputs(3146) <= (layer2_outputs(7340)) xor (layer2_outputs(3571));
    layer3_outputs(3147) <= (layer2_outputs(652)) and (layer2_outputs(2468));
    layer3_outputs(3148) <= layer2_outputs(3729);
    layer3_outputs(3149) <= (layer2_outputs(6234)) or (layer2_outputs(7305));
    layer3_outputs(3150) <= layer2_outputs(5476);
    layer3_outputs(3151) <= not(layer2_outputs(257)) or (layer2_outputs(5010));
    layer3_outputs(3152) <= (layer2_outputs(2592)) and (layer2_outputs(4340));
    layer3_outputs(3153) <= not(layer2_outputs(1568));
    layer3_outputs(3154) <= (layer2_outputs(261)) and not (layer2_outputs(6166));
    layer3_outputs(3155) <= '1';
    layer3_outputs(3156) <= (layer2_outputs(4961)) or (layer2_outputs(32));
    layer3_outputs(3157) <= layer2_outputs(5678);
    layer3_outputs(3158) <= not((layer2_outputs(6485)) and (layer2_outputs(2321)));
    layer3_outputs(3159) <= (layer2_outputs(1275)) and not (layer2_outputs(4578));
    layer3_outputs(3160) <= not(layer2_outputs(2205));
    layer3_outputs(3161) <= (layer2_outputs(6352)) or (layer2_outputs(4634));
    layer3_outputs(3162) <= not(layer2_outputs(4476));
    layer3_outputs(3163) <= layer2_outputs(3436);
    layer3_outputs(3164) <= '0';
    layer3_outputs(3165) <= not(layer2_outputs(640));
    layer3_outputs(3166) <= (layer2_outputs(3259)) or (layer2_outputs(5079));
    layer3_outputs(3167) <= not(layer2_outputs(60));
    layer3_outputs(3168) <= not(layer2_outputs(7061));
    layer3_outputs(3169) <= not(layer2_outputs(7228));
    layer3_outputs(3170) <= not((layer2_outputs(7116)) and (layer2_outputs(5818)));
    layer3_outputs(3171) <= layer2_outputs(1648);
    layer3_outputs(3172) <= layer2_outputs(412);
    layer3_outputs(3173) <= not(layer2_outputs(2154)) or (layer2_outputs(1511));
    layer3_outputs(3174) <= not((layer2_outputs(4341)) xor (layer2_outputs(807)));
    layer3_outputs(3175) <= layer2_outputs(1470);
    layer3_outputs(3176) <= layer2_outputs(6119);
    layer3_outputs(3177) <= layer2_outputs(3858);
    layer3_outputs(3178) <= (layer2_outputs(1222)) or (layer2_outputs(6859));
    layer3_outputs(3179) <= layer2_outputs(2402);
    layer3_outputs(3180) <= not(layer2_outputs(6293));
    layer3_outputs(3181) <= (layer2_outputs(2555)) and not (layer2_outputs(7190));
    layer3_outputs(3182) <= layer2_outputs(722);
    layer3_outputs(3183) <= not(layer2_outputs(33));
    layer3_outputs(3184) <= (layer2_outputs(223)) and not (layer2_outputs(1678));
    layer3_outputs(3185) <= not((layer2_outputs(4838)) and (layer2_outputs(2110)));
    layer3_outputs(3186) <= not(layer2_outputs(7273));
    layer3_outputs(3187) <= '0';
    layer3_outputs(3188) <= not(layer2_outputs(5682));
    layer3_outputs(3189) <= not((layer2_outputs(889)) or (layer2_outputs(3560)));
    layer3_outputs(3190) <= (layer2_outputs(2164)) and not (layer2_outputs(195));
    layer3_outputs(3191) <= not(layer2_outputs(1889)) or (layer2_outputs(1243));
    layer3_outputs(3192) <= not(layer2_outputs(7006)) or (layer2_outputs(4264));
    layer3_outputs(3193) <= (layer2_outputs(6884)) and not (layer2_outputs(7006));
    layer3_outputs(3194) <= not(layer2_outputs(1665));
    layer3_outputs(3195) <= '0';
    layer3_outputs(3196) <= '0';
    layer3_outputs(3197) <= not((layer2_outputs(4978)) or (layer2_outputs(1968)));
    layer3_outputs(3198) <= not(layer2_outputs(4617)) or (layer2_outputs(6127));
    layer3_outputs(3199) <= (layer2_outputs(1822)) and not (layer2_outputs(868));
    layer3_outputs(3200) <= not(layer2_outputs(2073));
    layer3_outputs(3201) <= '0';
    layer3_outputs(3202) <= not(layer2_outputs(7437));
    layer3_outputs(3203) <= layer2_outputs(4652);
    layer3_outputs(3204) <= not(layer2_outputs(5580)) or (layer2_outputs(3891));
    layer3_outputs(3205) <= not((layer2_outputs(1704)) or (layer2_outputs(4065)));
    layer3_outputs(3206) <= (layer2_outputs(4610)) and not (layer2_outputs(5388));
    layer3_outputs(3207) <= (layer2_outputs(1729)) and not (layer2_outputs(6769));
    layer3_outputs(3208) <= layer2_outputs(3985);
    layer3_outputs(3209) <= layer2_outputs(2297);
    layer3_outputs(3210) <= layer2_outputs(5007);
    layer3_outputs(3211) <= not(layer2_outputs(2121));
    layer3_outputs(3212) <= layer2_outputs(619);
    layer3_outputs(3213) <= not((layer2_outputs(6993)) or (layer2_outputs(5304)));
    layer3_outputs(3214) <= (layer2_outputs(6419)) or (layer2_outputs(6686));
    layer3_outputs(3215) <= layer2_outputs(6725);
    layer3_outputs(3216) <= (layer2_outputs(6881)) or (layer2_outputs(2403));
    layer3_outputs(3217) <= (layer2_outputs(4227)) or (layer2_outputs(5494));
    layer3_outputs(3218) <= not((layer2_outputs(2065)) xor (layer2_outputs(3716)));
    layer3_outputs(3219) <= '1';
    layer3_outputs(3220) <= not(layer2_outputs(4914)) or (layer2_outputs(3984));
    layer3_outputs(3221) <= not(layer2_outputs(3479));
    layer3_outputs(3222) <= not((layer2_outputs(6054)) or (layer2_outputs(5280)));
    layer3_outputs(3223) <= layer2_outputs(5322);
    layer3_outputs(3224) <= not(layer2_outputs(1258));
    layer3_outputs(3225) <= (layer2_outputs(3295)) and not (layer2_outputs(6663));
    layer3_outputs(3226) <= not(layer2_outputs(2345));
    layer3_outputs(3227) <= not(layer2_outputs(844));
    layer3_outputs(3228) <= not(layer2_outputs(1032)) or (layer2_outputs(5848));
    layer3_outputs(3229) <= not(layer2_outputs(6344)) or (layer2_outputs(4379));
    layer3_outputs(3230) <= (layer2_outputs(5019)) or (layer2_outputs(1451));
    layer3_outputs(3231) <= layer2_outputs(3652);
    layer3_outputs(3232) <= not(layer2_outputs(7358));
    layer3_outputs(3233) <= layer2_outputs(4370);
    layer3_outputs(3234) <= layer2_outputs(7);
    layer3_outputs(3235) <= not(layer2_outputs(7611));
    layer3_outputs(3236) <= layer2_outputs(7403);
    layer3_outputs(3237) <= (layer2_outputs(3448)) and (layer2_outputs(807));
    layer3_outputs(3238) <= (layer2_outputs(7361)) xor (layer2_outputs(7584));
    layer3_outputs(3239) <= layer2_outputs(855);
    layer3_outputs(3240) <= (layer2_outputs(660)) and not (layer2_outputs(5128));
    layer3_outputs(3241) <= layer2_outputs(6212);
    layer3_outputs(3242) <= (layer2_outputs(4209)) and not (layer2_outputs(5383));
    layer3_outputs(3243) <= not(layer2_outputs(4592));
    layer3_outputs(3244) <= (layer2_outputs(7252)) and not (layer2_outputs(4262));
    layer3_outputs(3245) <= not(layer2_outputs(3306));
    layer3_outputs(3246) <= not((layer2_outputs(3144)) xor (layer2_outputs(7095)));
    layer3_outputs(3247) <= (layer2_outputs(5375)) and not (layer2_outputs(65));
    layer3_outputs(3248) <= layer2_outputs(2991);
    layer3_outputs(3249) <= not(layer2_outputs(586)) or (layer2_outputs(2027));
    layer3_outputs(3250) <= '0';
    layer3_outputs(3251) <= '0';
    layer3_outputs(3252) <= '1';
    layer3_outputs(3253) <= not(layer2_outputs(6946));
    layer3_outputs(3254) <= layer2_outputs(4632);
    layer3_outputs(3255) <= layer2_outputs(402);
    layer3_outputs(3256) <= layer2_outputs(6631);
    layer3_outputs(3257) <= '0';
    layer3_outputs(3258) <= (layer2_outputs(3015)) and not (layer2_outputs(7338));
    layer3_outputs(3259) <= (layer2_outputs(1017)) and (layer2_outputs(7482));
    layer3_outputs(3260) <= (layer2_outputs(4439)) or (layer2_outputs(6923));
    layer3_outputs(3261) <= (layer2_outputs(59)) and not (layer2_outputs(1258));
    layer3_outputs(3262) <= '0';
    layer3_outputs(3263) <= not(layer2_outputs(1328));
    layer3_outputs(3264) <= (layer2_outputs(1059)) or (layer2_outputs(2199));
    layer3_outputs(3265) <= '0';
    layer3_outputs(3266) <= layer2_outputs(1399);
    layer3_outputs(3267) <= not((layer2_outputs(6412)) and (layer2_outputs(6223)));
    layer3_outputs(3268) <= (layer2_outputs(6296)) or (layer2_outputs(1940));
    layer3_outputs(3269) <= layer2_outputs(3358);
    layer3_outputs(3270) <= not(layer2_outputs(5408));
    layer3_outputs(3271) <= not(layer2_outputs(7672));
    layer3_outputs(3272) <= (layer2_outputs(3087)) or (layer2_outputs(2610));
    layer3_outputs(3273) <= (layer2_outputs(927)) and not (layer2_outputs(5048));
    layer3_outputs(3274) <= not((layer2_outputs(1961)) and (layer2_outputs(5257)));
    layer3_outputs(3275) <= (layer2_outputs(2886)) or (layer2_outputs(2603));
    layer3_outputs(3276) <= not((layer2_outputs(7409)) xor (layer2_outputs(2571)));
    layer3_outputs(3277) <= layer2_outputs(865);
    layer3_outputs(3278) <= not((layer2_outputs(525)) and (layer2_outputs(3584)));
    layer3_outputs(3279) <= (layer2_outputs(5587)) and (layer2_outputs(2253));
    layer3_outputs(3280) <= (layer2_outputs(771)) and not (layer2_outputs(7535));
    layer3_outputs(3281) <= '0';
    layer3_outputs(3282) <= not((layer2_outputs(4076)) and (layer2_outputs(6265)));
    layer3_outputs(3283) <= '0';
    layer3_outputs(3284) <= (layer2_outputs(4512)) or (layer2_outputs(6184));
    layer3_outputs(3285) <= not((layer2_outputs(5637)) and (layer2_outputs(7470)));
    layer3_outputs(3286) <= not(layer2_outputs(2143)) or (layer2_outputs(538));
    layer3_outputs(3287) <= not(layer2_outputs(4145));
    layer3_outputs(3288) <= (layer2_outputs(1530)) and (layer2_outputs(4445));
    layer3_outputs(3289) <= not(layer2_outputs(7085));
    layer3_outputs(3290) <= layer2_outputs(2501);
    layer3_outputs(3291) <= '0';
    layer3_outputs(3292) <= '0';
    layer3_outputs(3293) <= not(layer2_outputs(3666));
    layer3_outputs(3294) <= (layer2_outputs(7500)) and not (layer2_outputs(4365));
    layer3_outputs(3295) <= not(layer2_outputs(1005)) or (layer2_outputs(2175));
    layer3_outputs(3296) <= not(layer2_outputs(5245));
    layer3_outputs(3297) <= not(layer2_outputs(3836));
    layer3_outputs(3298) <= '1';
    layer3_outputs(3299) <= not((layer2_outputs(4864)) or (layer2_outputs(7198)));
    layer3_outputs(3300) <= '1';
    layer3_outputs(3301) <= not((layer2_outputs(6624)) and (layer2_outputs(2280)));
    layer3_outputs(3302) <= (layer2_outputs(3751)) and (layer2_outputs(606));
    layer3_outputs(3303) <= (layer2_outputs(6307)) and not (layer2_outputs(1581));
    layer3_outputs(3304) <= '0';
    layer3_outputs(3305) <= not(layer2_outputs(6211));
    layer3_outputs(3306) <= not((layer2_outputs(3341)) and (layer2_outputs(2859)));
    layer3_outputs(3307) <= not(layer2_outputs(6484)) or (layer2_outputs(5443));
    layer3_outputs(3308) <= not(layer2_outputs(916));
    layer3_outputs(3309) <= not(layer2_outputs(295));
    layer3_outputs(3310) <= not((layer2_outputs(4880)) xor (layer2_outputs(1982)));
    layer3_outputs(3311) <= not(layer2_outputs(6106));
    layer3_outputs(3312) <= not((layer2_outputs(3659)) and (layer2_outputs(2747)));
    layer3_outputs(3313) <= '1';
    layer3_outputs(3314) <= (layer2_outputs(5297)) and (layer2_outputs(4219));
    layer3_outputs(3315) <= layer2_outputs(6584);
    layer3_outputs(3316) <= (layer2_outputs(7195)) or (layer2_outputs(2686));
    layer3_outputs(3317) <= not(layer2_outputs(1482));
    layer3_outputs(3318) <= not(layer2_outputs(3385));
    layer3_outputs(3319) <= (layer2_outputs(6060)) and not (layer2_outputs(2649));
    layer3_outputs(3320) <= layer2_outputs(5017);
    layer3_outputs(3321) <= not(layer2_outputs(3344));
    layer3_outputs(3322) <= (layer2_outputs(1631)) and (layer2_outputs(2346));
    layer3_outputs(3323) <= '0';
    layer3_outputs(3324) <= not((layer2_outputs(3126)) and (layer2_outputs(1938)));
    layer3_outputs(3325) <= not((layer2_outputs(2098)) and (layer2_outputs(1036)));
    layer3_outputs(3326) <= (layer2_outputs(6432)) and (layer2_outputs(4551));
    layer3_outputs(3327) <= not(layer2_outputs(7432));
    layer3_outputs(3328) <= not((layer2_outputs(7277)) and (layer2_outputs(5737)));
    layer3_outputs(3329) <= not(layer2_outputs(2401));
    layer3_outputs(3330) <= layer2_outputs(264);
    layer3_outputs(3331) <= (layer2_outputs(2181)) and (layer2_outputs(2287));
    layer3_outputs(3332) <= layer2_outputs(6771);
    layer3_outputs(3333) <= (layer2_outputs(3948)) and not (layer2_outputs(1436));
    layer3_outputs(3334) <= not(layer2_outputs(5961)) or (layer2_outputs(4894));
    layer3_outputs(3335) <= layer2_outputs(6741);
    layer3_outputs(3336) <= (layer2_outputs(6460)) and not (layer2_outputs(1722));
    layer3_outputs(3337) <= not(layer2_outputs(5857));
    layer3_outputs(3338) <= layer2_outputs(3747);
    layer3_outputs(3339) <= (layer2_outputs(3884)) xor (layer2_outputs(6189));
    layer3_outputs(3340) <= not((layer2_outputs(1535)) xor (layer2_outputs(3846)));
    layer3_outputs(3341) <= layer2_outputs(3803);
    layer3_outputs(3342) <= '0';
    layer3_outputs(3343) <= layer2_outputs(5254);
    layer3_outputs(3344) <= layer2_outputs(894);
    layer3_outputs(3345) <= '1';
    layer3_outputs(3346) <= layer2_outputs(4504);
    layer3_outputs(3347) <= '1';
    layer3_outputs(3348) <= not(layer2_outputs(4177));
    layer3_outputs(3349) <= layer2_outputs(6013);
    layer3_outputs(3350) <= not(layer2_outputs(3939)) or (layer2_outputs(7429));
    layer3_outputs(3351) <= (layer2_outputs(3344)) and not (layer2_outputs(6190));
    layer3_outputs(3352) <= (layer2_outputs(2270)) or (layer2_outputs(6663));
    layer3_outputs(3353) <= layer2_outputs(6718);
    layer3_outputs(3354) <= (layer2_outputs(4681)) and (layer2_outputs(6638));
    layer3_outputs(3355) <= (layer2_outputs(1166)) and not (layer2_outputs(24));
    layer3_outputs(3356) <= layer2_outputs(1266);
    layer3_outputs(3357) <= (layer2_outputs(1751)) or (layer2_outputs(3131));
    layer3_outputs(3358) <= layer2_outputs(5510);
    layer3_outputs(3359) <= (layer2_outputs(7577)) and not (layer2_outputs(7240));
    layer3_outputs(3360) <= (layer2_outputs(7114)) and not (layer2_outputs(490));
    layer3_outputs(3361) <= layer2_outputs(6012);
    layer3_outputs(3362) <= not(layer2_outputs(4799)) or (layer2_outputs(475));
    layer3_outputs(3363) <= (layer2_outputs(1568)) and not (layer2_outputs(1206));
    layer3_outputs(3364) <= not(layer2_outputs(163)) or (layer2_outputs(6316));
    layer3_outputs(3365) <= layer2_outputs(434);
    layer3_outputs(3366) <= not(layer2_outputs(6001)) or (layer2_outputs(7636));
    layer3_outputs(3367) <= not(layer2_outputs(3341));
    layer3_outputs(3368) <= layer2_outputs(3166);
    layer3_outputs(3369) <= not((layer2_outputs(5152)) or (layer2_outputs(848)));
    layer3_outputs(3370) <= '0';
    layer3_outputs(3371) <= not(layer2_outputs(5885)) or (layer2_outputs(3185));
    layer3_outputs(3372) <= not(layer2_outputs(5280)) or (layer2_outputs(1510));
    layer3_outputs(3373) <= (layer2_outputs(2208)) and (layer2_outputs(6706));
    layer3_outputs(3374) <= '1';
    layer3_outputs(3375) <= not((layer2_outputs(6030)) and (layer2_outputs(972)));
    layer3_outputs(3376) <= not((layer2_outputs(6933)) xor (layer2_outputs(4747)));
    layer3_outputs(3377) <= not(layer2_outputs(1723));
    layer3_outputs(3378) <= '1';
    layer3_outputs(3379) <= '1';
    layer3_outputs(3380) <= not((layer2_outputs(1741)) or (layer2_outputs(3318)));
    layer3_outputs(3381) <= not(layer2_outputs(327));
    layer3_outputs(3382) <= (layer2_outputs(3456)) and not (layer2_outputs(787));
    layer3_outputs(3383) <= not((layer2_outputs(7600)) xor (layer2_outputs(1746)));
    layer3_outputs(3384) <= not((layer2_outputs(6138)) xor (layer2_outputs(4217)));
    layer3_outputs(3385) <= not(layer2_outputs(1351)) or (layer2_outputs(4036));
    layer3_outputs(3386) <= '0';
    layer3_outputs(3387) <= not(layer2_outputs(7209));
    layer3_outputs(3388) <= not(layer2_outputs(7419));
    layer3_outputs(3389) <= (layer2_outputs(4789)) and not (layer2_outputs(6289));
    layer3_outputs(3390) <= (layer2_outputs(4239)) and (layer2_outputs(6561));
    layer3_outputs(3391) <= not(layer2_outputs(4650));
    layer3_outputs(3392) <= (layer2_outputs(2292)) or (layer2_outputs(2768));
    layer3_outputs(3393) <= layer2_outputs(6825);
    layer3_outputs(3394) <= (layer2_outputs(1197)) and (layer2_outputs(1389));
    layer3_outputs(3395) <= '0';
    layer3_outputs(3396) <= not(layer2_outputs(2030)) or (layer2_outputs(5838));
    layer3_outputs(3397) <= not(layer2_outputs(4176)) or (layer2_outputs(1171));
    layer3_outputs(3398) <= not(layer2_outputs(2339));
    layer3_outputs(3399) <= (layer2_outputs(4485)) and (layer2_outputs(6060));
    layer3_outputs(3400) <= not(layer2_outputs(1972)) or (layer2_outputs(1242));
    layer3_outputs(3401) <= (layer2_outputs(1874)) and not (layer2_outputs(2384));
    layer3_outputs(3402) <= layer2_outputs(3597);
    layer3_outputs(3403) <= not((layer2_outputs(1021)) or (layer2_outputs(1970)));
    layer3_outputs(3404) <= not(layer2_outputs(5524));
    layer3_outputs(3405) <= '0';
    layer3_outputs(3406) <= '0';
    layer3_outputs(3407) <= '0';
    layer3_outputs(3408) <= not(layer2_outputs(2057));
    layer3_outputs(3409) <= layer2_outputs(2016);
    layer3_outputs(3410) <= not(layer2_outputs(2179)) or (layer2_outputs(1914));
    layer3_outputs(3411) <= not((layer2_outputs(815)) xor (layer2_outputs(4306)));
    layer3_outputs(3412) <= layer2_outputs(7054);
    layer3_outputs(3413) <= (layer2_outputs(5608)) or (layer2_outputs(6802));
    layer3_outputs(3414) <= layer2_outputs(7628);
    layer3_outputs(3415) <= not(layer2_outputs(6527));
    layer3_outputs(3416) <= not(layer2_outputs(689));
    layer3_outputs(3417) <= '0';
    layer3_outputs(3418) <= (layer2_outputs(842)) or (layer2_outputs(6718));
    layer3_outputs(3419) <= layer2_outputs(3581);
    layer3_outputs(3420) <= (layer2_outputs(966)) or (layer2_outputs(5464));
    layer3_outputs(3421) <= layer2_outputs(4045);
    layer3_outputs(3422) <= not(layer2_outputs(7075)) or (layer2_outputs(4809));
    layer3_outputs(3423) <= layer2_outputs(5763);
    layer3_outputs(3424) <= not(layer2_outputs(1038)) or (layer2_outputs(5653));
    layer3_outputs(3425) <= not(layer2_outputs(3131));
    layer3_outputs(3426) <= not(layer2_outputs(3158));
    layer3_outputs(3427) <= not((layer2_outputs(5518)) xor (layer2_outputs(7666)));
    layer3_outputs(3428) <= '1';
    layer3_outputs(3429) <= '0';
    layer3_outputs(3430) <= not(layer2_outputs(5254)) or (layer2_outputs(1592));
    layer3_outputs(3431) <= '1';
    layer3_outputs(3432) <= (layer2_outputs(1809)) or (layer2_outputs(7117));
    layer3_outputs(3433) <= (layer2_outputs(6407)) or (layer2_outputs(7216));
    layer3_outputs(3434) <= not(layer2_outputs(4543));
    layer3_outputs(3435) <= not((layer2_outputs(6787)) or (layer2_outputs(5825)));
    layer3_outputs(3436) <= '0';
    layer3_outputs(3437) <= layer2_outputs(2267);
    layer3_outputs(3438) <= not(layer2_outputs(699)) or (layer2_outputs(7203));
    layer3_outputs(3439) <= '1';
    layer3_outputs(3440) <= (layer2_outputs(4360)) and (layer2_outputs(1153));
    layer3_outputs(3441) <= not((layer2_outputs(6917)) xor (layer2_outputs(2700)));
    layer3_outputs(3442) <= not((layer2_outputs(7306)) or (layer2_outputs(6075)));
    layer3_outputs(3443) <= not(layer2_outputs(6615)) or (layer2_outputs(5423));
    layer3_outputs(3444) <= layer2_outputs(5315);
    layer3_outputs(3445) <= '1';
    layer3_outputs(3446) <= layer2_outputs(7436);
    layer3_outputs(3447) <= not(layer2_outputs(1426)) or (layer2_outputs(2128));
    layer3_outputs(3448) <= not(layer2_outputs(3611));
    layer3_outputs(3449) <= not((layer2_outputs(6781)) and (layer2_outputs(2585)));
    layer3_outputs(3450) <= '1';
    layer3_outputs(3451) <= not(layer2_outputs(6438));
    layer3_outputs(3452) <= not((layer2_outputs(2280)) and (layer2_outputs(881)));
    layer3_outputs(3453) <= not((layer2_outputs(1612)) and (layer2_outputs(372)));
    layer3_outputs(3454) <= not(layer2_outputs(2324));
    layer3_outputs(3455) <= layer2_outputs(1645);
    layer3_outputs(3456) <= not(layer2_outputs(4167));
    layer3_outputs(3457) <= (layer2_outputs(6128)) or (layer2_outputs(3307));
    layer3_outputs(3458) <= layer2_outputs(3930);
    layer3_outputs(3459) <= not((layer2_outputs(6969)) or (layer2_outputs(931)));
    layer3_outputs(3460) <= not((layer2_outputs(6755)) and (layer2_outputs(1146)));
    layer3_outputs(3461) <= not((layer2_outputs(264)) and (layer2_outputs(7023)));
    layer3_outputs(3462) <= not((layer2_outputs(4619)) or (layer2_outputs(3727)));
    layer3_outputs(3463) <= not(layer2_outputs(7295));
    layer3_outputs(3464) <= (layer2_outputs(7319)) and not (layer2_outputs(1212));
    layer3_outputs(3465) <= not((layer2_outputs(159)) or (layer2_outputs(1074)));
    layer3_outputs(3466) <= (layer2_outputs(7646)) and (layer2_outputs(1319));
    layer3_outputs(3467) <= (layer2_outputs(3551)) or (layer2_outputs(1673));
    layer3_outputs(3468) <= layer2_outputs(1207);
    layer3_outputs(3469) <= not(layer2_outputs(1271));
    layer3_outputs(3470) <= layer2_outputs(5338);
    layer3_outputs(3471) <= not((layer2_outputs(7546)) and (layer2_outputs(1073)));
    layer3_outputs(3472) <= (layer2_outputs(5086)) and not (layer2_outputs(3667));
    layer3_outputs(3473) <= '0';
    layer3_outputs(3474) <= not(layer2_outputs(3562));
    layer3_outputs(3475) <= (layer2_outputs(6584)) and not (layer2_outputs(199));
    layer3_outputs(3476) <= not(layer2_outputs(4819));
    layer3_outputs(3477) <= layer2_outputs(5537);
    layer3_outputs(3478) <= not(layer2_outputs(6088)) or (layer2_outputs(5499));
    layer3_outputs(3479) <= not(layer2_outputs(7403));
    layer3_outputs(3480) <= (layer2_outputs(2644)) and (layer2_outputs(4869));
    layer3_outputs(3481) <= (layer2_outputs(2311)) and not (layer2_outputs(217));
    layer3_outputs(3482) <= not(layer2_outputs(5507));
    layer3_outputs(3483) <= '1';
    layer3_outputs(3484) <= layer2_outputs(6330);
    layer3_outputs(3485) <= not((layer2_outputs(4291)) and (layer2_outputs(5699)));
    layer3_outputs(3486) <= not(layer2_outputs(5242)) or (layer2_outputs(1554));
    layer3_outputs(3487) <= not((layer2_outputs(1927)) or (layer2_outputs(4187)));
    layer3_outputs(3488) <= (layer2_outputs(1269)) and not (layer2_outputs(14));
    layer3_outputs(3489) <= not(layer2_outputs(1004));
    layer3_outputs(3490) <= layer2_outputs(793);
    layer3_outputs(3491) <= (layer2_outputs(1051)) or (layer2_outputs(2434));
    layer3_outputs(3492) <= layer2_outputs(6093);
    layer3_outputs(3493) <= '1';
    layer3_outputs(3494) <= '1';
    layer3_outputs(3495) <= not(layer2_outputs(3619));
    layer3_outputs(3496) <= not(layer2_outputs(3649));
    layer3_outputs(3497) <= '0';
    layer3_outputs(3498) <= not((layer2_outputs(5554)) or (layer2_outputs(4714)));
    layer3_outputs(3499) <= layer2_outputs(3347);
    layer3_outputs(3500) <= layer2_outputs(4630);
    layer3_outputs(3501) <= layer2_outputs(4436);
    layer3_outputs(3502) <= layer2_outputs(1833);
    layer3_outputs(3503) <= not(layer2_outputs(3409));
    layer3_outputs(3504) <= not(layer2_outputs(628));
    layer3_outputs(3505) <= (layer2_outputs(29)) and not (layer2_outputs(361));
    layer3_outputs(3506) <= '0';
    layer3_outputs(3507) <= not(layer2_outputs(864));
    layer3_outputs(3508) <= (layer2_outputs(554)) and (layer2_outputs(5785));
    layer3_outputs(3509) <= (layer2_outputs(5883)) and not (layer2_outputs(643));
    layer3_outputs(3510) <= layer2_outputs(7554);
    layer3_outputs(3511) <= not(layer2_outputs(1870));
    layer3_outputs(3512) <= not(layer2_outputs(421));
    layer3_outputs(3513) <= '1';
    layer3_outputs(3514) <= not(layer2_outputs(5366));
    layer3_outputs(3515) <= layer2_outputs(5575);
    layer3_outputs(3516) <= layer2_outputs(4125);
    layer3_outputs(3517) <= '0';
    layer3_outputs(3518) <= layer2_outputs(6872);
    layer3_outputs(3519) <= not(layer2_outputs(3033));
    layer3_outputs(3520) <= '0';
    layer3_outputs(3521) <= not(layer2_outputs(5513));
    layer3_outputs(3522) <= (layer2_outputs(3981)) and not (layer2_outputs(2144));
    layer3_outputs(3523) <= not(layer2_outputs(6607)) or (layer2_outputs(3896));
    layer3_outputs(3524) <= (layer2_outputs(6006)) and not (layer2_outputs(2012));
    layer3_outputs(3525) <= not(layer2_outputs(1988));
    layer3_outputs(3526) <= not(layer2_outputs(3810)) or (layer2_outputs(4256));
    layer3_outputs(3527) <= (layer2_outputs(384)) and (layer2_outputs(5111));
    layer3_outputs(3528) <= not(layer2_outputs(4074)) or (layer2_outputs(4544));
    layer3_outputs(3529) <= not((layer2_outputs(278)) or (layer2_outputs(2808)));
    layer3_outputs(3530) <= not(layer2_outputs(6641));
    layer3_outputs(3531) <= '0';
    layer3_outputs(3532) <= '1';
    layer3_outputs(3533) <= (layer2_outputs(1941)) and not (layer2_outputs(1376));
    layer3_outputs(3534) <= not(layer2_outputs(4412));
    layer3_outputs(3535) <= '0';
    layer3_outputs(3536) <= '0';
    layer3_outputs(3537) <= layer2_outputs(5170);
    layer3_outputs(3538) <= (layer2_outputs(358)) or (layer2_outputs(3611));
    layer3_outputs(3539) <= layer2_outputs(7363);
    layer3_outputs(3540) <= (layer2_outputs(5450)) and not (layer2_outputs(4383));
    layer3_outputs(3541) <= not(layer2_outputs(4487)) or (layer2_outputs(4271));
    layer3_outputs(3542) <= not(layer2_outputs(5540)) or (layer2_outputs(4877));
    layer3_outputs(3543) <= not(layer2_outputs(505)) or (layer2_outputs(6829));
    layer3_outputs(3544) <= not(layer2_outputs(5064)) or (layer2_outputs(5016));
    layer3_outputs(3545) <= (layer2_outputs(3066)) and not (layer2_outputs(1559));
    layer3_outputs(3546) <= not(layer2_outputs(1073)) or (layer2_outputs(2717));
    layer3_outputs(3547) <= (layer2_outputs(1003)) and not (layer2_outputs(1613));
    layer3_outputs(3548) <= (layer2_outputs(3628)) and not (layer2_outputs(202));
    layer3_outputs(3549) <= not((layer2_outputs(6390)) or (layer2_outputs(2556)));
    layer3_outputs(3550) <= (layer2_outputs(4509)) and (layer2_outputs(533));
    layer3_outputs(3551) <= (layer2_outputs(5068)) and not (layer2_outputs(446));
    layer3_outputs(3552) <= not(layer2_outputs(3282));
    layer3_outputs(3553) <= (layer2_outputs(3455)) and not (layer2_outputs(318));
    layer3_outputs(3554) <= not(layer2_outputs(4968)) or (layer2_outputs(1745));
    layer3_outputs(3555) <= not(layer2_outputs(6516));
    layer3_outputs(3556) <= layer2_outputs(5337);
    layer3_outputs(3557) <= not(layer2_outputs(1400));
    layer3_outputs(3558) <= (layer2_outputs(2305)) and not (layer2_outputs(943));
    layer3_outputs(3559) <= not((layer2_outputs(2904)) and (layer2_outputs(6503)));
    layer3_outputs(3560) <= not(layer2_outputs(773));
    layer3_outputs(3561) <= (layer2_outputs(5847)) or (layer2_outputs(320));
    layer3_outputs(3562) <= (layer2_outputs(309)) and not (layer2_outputs(7124));
    layer3_outputs(3563) <= not((layer2_outputs(1322)) xor (layer2_outputs(5063)));
    layer3_outputs(3564) <= (layer2_outputs(3753)) and not (layer2_outputs(3340));
    layer3_outputs(3565) <= (layer2_outputs(490)) and (layer2_outputs(3311));
    layer3_outputs(3566) <= '1';
    layer3_outputs(3567) <= '1';
    layer3_outputs(3568) <= (layer2_outputs(1020)) and (layer2_outputs(1206));
    layer3_outputs(3569) <= not(layer2_outputs(6446));
    layer3_outputs(3570) <= not(layer2_outputs(4896));
    layer3_outputs(3571) <= layer2_outputs(6271);
    layer3_outputs(3572) <= not(layer2_outputs(3508)) or (layer2_outputs(6089));
    layer3_outputs(3573) <= layer2_outputs(2868);
    layer3_outputs(3574) <= layer2_outputs(2855);
    layer3_outputs(3575) <= not(layer2_outputs(1495));
    layer3_outputs(3576) <= not((layer2_outputs(3671)) or (layer2_outputs(2798)));
    layer3_outputs(3577) <= (layer2_outputs(6804)) and (layer2_outputs(6020));
    layer3_outputs(3578) <= not(layer2_outputs(2347));
    layer3_outputs(3579) <= not((layer2_outputs(6635)) and (layer2_outputs(2209)));
    layer3_outputs(3580) <= not(layer2_outputs(335));
    layer3_outputs(3581) <= (layer2_outputs(5326)) xor (layer2_outputs(4003));
    layer3_outputs(3582) <= (layer2_outputs(671)) and not (layer2_outputs(6483));
    layer3_outputs(3583) <= not(layer2_outputs(506));
    layer3_outputs(3584) <= '1';
    layer3_outputs(3585) <= not((layer2_outputs(81)) or (layer2_outputs(3109)));
    layer3_outputs(3586) <= (layer2_outputs(653)) and not (layer2_outputs(3850));
    layer3_outputs(3587) <= not(layer2_outputs(7408)) or (layer2_outputs(5043));
    layer3_outputs(3588) <= '1';
    layer3_outputs(3589) <= not((layer2_outputs(400)) xor (layer2_outputs(42)));
    layer3_outputs(3590) <= not((layer2_outputs(4137)) and (layer2_outputs(1405)));
    layer3_outputs(3591) <= not(layer2_outputs(6339)) or (layer2_outputs(696));
    layer3_outputs(3592) <= not((layer2_outputs(140)) or (layer2_outputs(324)));
    layer3_outputs(3593) <= layer2_outputs(1152);
    layer3_outputs(3594) <= not(layer2_outputs(1712));
    layer3_outputs(3595) <= '1';
    layer3_outputs(3596) <= layer2_outputs(6232);
    layer3_outputs(3597) <= layer2_outputs(544);
    layer3_outputs(3598) <= layer2_outputs(6955);
    layer3_outputs(3599) <= not(layer2_outputs(5059));
    layer3_outputs(3600) <= layer2_outputs(6648);
    layer3_outputs(3601) <= (layer2_outputs(3183)) and not (layer2_outputs(3630));
    layer3_outputs(3602) <= (layer2_outputs(471)) and (layer2_outputs(2372));
    layer3_outputs(3603) <= layer2_outputs(7022);
    layer3_outputs(3604) <= not((layer2_outputs(3771)) and (layer2_outputs(6779)));
    layer3_outputs(3605) <= not(layer2_outputs(1210)) or (layer2_outputs(5385));
    layer3_outputs(3606) <= (layer2_outputs(636)) and (layer2_outputs(6297));
    layer3_outputs(3607) <= (layer2_outputs(6250)) xor (layer2_outputs(4639));
    layer3_outputs(3608) <= '0';
    layer3_outputs(3609) <= not(layer2_outputs(1214));
    layer3_outputs(3610) <= not(layer2_outputs(6086)) or (layer2_outputs(2067));
    layer3_outputs(3611) <= not((layer2_outputs(5999)) xor (layer2_outputs(5448)));
    layer3_outputs(3612) <= not(layer2_outputs(3877)) or (layer2_outputs(5));
    layer3_outputs(3613) <= (layer2_outputs(1660)) and (layer2_outputs(478));
    layer3_outputs(3614) <= not(layer2_outputs(4960));
    layer3_outputs(3615) <= '1';
    layer3_outputs(3616) <= layer2_outputs(315);
    layer3_outputs(3617) <= not((layer2_outputs(1963)) or (layer2_outputs(1478)));
    layer3_outputs(3618) <= layer2_outputs(5277);
    layer3_outputs(3619) <= layer2_outputs(6449);
    layer3_outputs(3620) <= (layer2_outputs(1224)) or (layer2_outputs(5053));
    layer3_outputs(3621) <= not(layer2_outputs(1315));
    layer3_outputs(3622) <= '0';
    layer3_outputs(3623) <= not(layer2_outputs(3520)) or (layer2_outputs(7436));
    layer3_outputs(3624) <= layer2_outputs(4694);
    layer3_outputs(3625) <= not((layer2_outputs(5915)) and (layer2_outputs(5710)));
    layer3_outputs(3626) <= not(layer2_outputs(4242)) or (layer2_outputs(5142));
    layer3_outputs(3627) <= (layer2_outputs(5867)) and not (layer2_outputs(6797));
    layer3_outputs(3628) <= not(layer2_outputs(723));
    layer3_outputs(3629) <= not(layer2_outputs(1));
    layer3_outputs(3630) <= '1';
    layer3_outputs(3631) <= not(layer2_outputs(6285));
    layer3_outputs(3632) <= layer2_outputs(4144);
    layer3_outputs(3633) <= layer2_outputs(3935);
    layer3_outputs(3634) <= not(layer2_outputs(5115)) or (layer2_outputs(4223));
    layer3_outputs(3635) <= '1';
    layer3_outputs(3636) <= '0';
    layer3_outputs(3637) <= layer2_outputs(2370);
    layer3_outputs(3638) <= (layer2_outputs(4540)) or (layer2_outputs(5217));
    layer3_outputs(3639) <= not(layer2_outputs(6834));
    layer3_outputs(3640) <= not(layer2_outputs(6251)) or (layer2_outputs(3763));
    layer3_outputs(3641) <= not(layer2_outputs(6205)) or (layer2_outputs(4438));
    layer3_outputs(3642) <= not(layer2_outputs(401));
    layer3_outputs(3643) <= '1';
    layer3_outputs(3644) <= '0';
    layer3_outputs(3645) <= not(layer2_outputs(6481)) or (layer2_outputs(241));
    layer3_outputs(3646) <= not(layer2_outputs(2505));
    layer3_outputs(3647) <= '0';
    layer3_outputs(3648) <= layer2_outputs(6549);
    layer3_outputs(3649) <= (layer2_outputs(4130)) and not (layer2_outputs(6225));
    layer3_outputs(3650) <= layer2_outputs(4790);
    layer3_outputs(3651) <= not(layer2_outputs(3291));
    layer3_outputs(3652) <= not(layer2_outputs(1447));
    layer3_outputs(3653) <= (layer2_outputs(3044)) and (layer2_outputs(5920));
    layer3_outputs(3654) <= not(layer2_outputs(4367));
    layer3_outputs(3655) <= (layer2_outputs(5070)) and not (layer2_outputs(146));
    layer3_outputs(3656) <= not((layer2_outputs(1440)) or (layer2_outputs(217)));
    layer3_outputs(3657) <= (layer2_outputs(4392)) or (layer2_outputs(4111));
    layer3_outputs(3658) <= not((layer2_outputs(7300)) and (layer2_outputs(165)));
    layer3_outputs(3659) <= not(layer2_outputs(5582));
    layer3_outputs(3660) <= '1';
    layer3_outputs(3661) <= layer2_outputs(4883);
    layer3_outputs(3662) <= not(layer2_outputs(4021)) or (layer2_outputs(4301));
    layer3_outputs(3663) <= not((layer2_outputs(16)) and (layer2_outputs(1691)));
    layer3_outputs(3664) <= not(layer2_outputs(887));
    layer3_outputs(3665) <= layer2_outputs(7011);
    layer3_outputs(3666) <= not(layer2_outputs(3209));
    layer3_outputs(3667) <= (layer2_outputs(5359)) xor (layer2_outputs(3036));
    layer3_outputs(3668) <= not(layer2_outputs(6832));
    layer3_outputs(3669) <= layer2_outputs(952);
    layer3_outputs(3670) <= not(layer2_outputs(754));
    layer3_outputs(3671) <= not(layer2_outputs(2774)) or (layer2_outputs(1398));
    layer3_outputs(3672) <= layer2_outputs(5150);
    layer3_outputs(3673) <= not(layer2_outputs(7121));
    layer3_outputs(3674) <= layer2_outputs(5809);
    layer3_outputs(3675) <= not(layer2_outputs(6366)) or (layer2_outputs(495));
    layer3_outputs(3676) <= (layer2_outputs(7280)) and not (layer2_outputs(3678));
    layer3_outputs(3677) <= (layer2_outputs(3292)) or (layer2_outputs(1252));
    layer3_outputs(3678) <= not((layer2_outputs(2369)) and (layer2_outputs(4192)));
    layer3_outputs(3679) <= not((layer2_outputs(3819)) and (layer2_outputs(4189)));
    layer3_outputs(3680) <= not(layer2_outputs(6587)) or (layer2_outputs(2947));
    layer3_outputs(3681) <= not(layer2_outputs(613));
    layer3_outputs(3682) <= layer2_outputs(2072);
    layer3_outputs(3683) <= layer2_outputs(5741);
    layer3_outputs(3684) <= not((layer2_outputs(2687)) or (layer2_outputs(1828)));
    layer3_outputs(3685) <= '0';
    layer3_outputs(3686) <= '1';
    layer3_outputs(3687) <= '0';
    layer3_outputs(3688) <= layer2_outputs(7386);
    layer3_outputs(3689) <= (layer2_outputs(6696)) and not (layer2_outputs(5072));
    layer3_outputs(3690) <= layer2_outputs(1433);
    layer3_outputs(3691) <= not(layer2_outputs(2871)) or (layer2_outputs(6907));
    layer3_outputs(3692) <= (layer2_outputs(2564)) and not (layer2_outputs(1663));
    layer3_outputs(3693) <= not(layer2_outputs(1506)) or (layer2_outputs(1390));
    layer3_outputs(3694) <= (layer2_outputs(3907)) or (layer2_outputs(3019));
    layer3_outputs(3695) <= layer2_outputs(6131);
    layer3_outputs(3696) <= not((layer2_outputs(3139)) xor (layer2_outputs(5763)));
    layer3_outputs(3697) <= not(layer2_outputs(4133));
    layer3_outputs(3698) <= layer2_outputs(4186);
    layer3_outputs(3699) <= not((layer2_outputs(1142)) and (layer2_outputs(6433)));
    layer3_outputs(3700) <= '1';
    layer3_outputs(3701) <= layer2_outputs(2745);
    layer3_outputs(3702) <= not(layer2_outputs(4359)) or (layer2_outputs(3060));
    layer3_outputs(3703) <= not((layer2_outputs(6454)) and (layer2_outputs(658)));
    layer3_outputs(3704) <= not(layer2_outputs(135));
    layer3_outputs(3705) <= not(layer2_outputs(4965));
    layer3_outputs(3706) <= not(layer2_outputs(2948)) or (layer2_outputs(4457));
    layer3_outputs(3707) <= '0';
    layer3_outputs(3708) <= not((layer2_outputs(7531)) or (layer2_outputs(4690)));
    layer3_outputs(3709) <= not(layer2_outputs(2222));
    layer3_outputs(3710) <= (layer2_outputs(4891)) or (layer2_outputs(5696));
    layer3_outputs(3711) <= (layer2_outputs(6142)) or (layer2_outputs(6122));
    layer3_outputs(3712) <= not((layer2_outputs(3044)) or (layer2_outputs(5457)));
    layer3_outputs(3713) <= (layer2_outputs(1494)) or (layer2_outputs(7110));
    layer3_outputs(3714) <= (layer2_outputs(7005)) and not (layer2_outputs(4980));
    layer3_outputs(3715) <= layer2_outputs(7648);
    layer3_outputs(3716) <= (layer2_outputs(6318)) and not (layer2_outputs(527));
    layer3_outputs(3717) <= not(layer2_outputs(2231)) or (layer2_outputs(3384));
    layer3_outputs(3718) <= not(layer2_outputs(4671)) or (layer2_outputs(5667));
    layer3_outputs(3719) <= '1';
    layer3_outputs(3720) <= not(layer2_outputs(3442)) or (layer2_outputs(5954));
    layer3_outputs(3721) <= (layer2_outputs(5267)) and not (layer2_outputs(1848));
    layer3_outputs(3722) <= not(layer2_outputs(1541));
    layer3_outputs(3723) <= not(layer2_outputs(5444)) or (layer2_outputs(4586));
    layer3_outputs(3724) <= (layer2_outputs(6847)) and not (layer2_outputs(3764));
    layer3_outputs(3725) <= not(layer2_outputs(4220));
    layer3_outputs(3726) <= not(layer2_outputs(1537)) or (layer2_outputs(802));
    layer3_outputs(3727) <= (layer2_outputs(1101)) and not (layer2_outputs(574));
    layer3_outputs(3728) <= (layer2_outputs(4302)) and not (layer2_outputs(3309));
    layer3_outputs(3729) <= not((layer2_outputs(1676)) or (layer2_outputs(7008)));
    layer3_outputs(3730) <= (layer2_outputs(6418)) xor (layer2_outputs(543));
    layer3_outputs(3731) <= not(layer2_outputs(4699)) or (layer2_outputs(6239));
    layer3_outputs(3732) <= not((layer2_outputs(2461)) and (layer2_outputs(7184)));
    layer3_outputs(3733) <= not((layer2_outputs(1382)) or (layer2_outputs(4813)));
    layer3_outputs(3734) <= not(layer2_outputs(2443));
    layer3_outputs(3735) <= layer2_outputs(575);
    layer3_outputs(3736) <= (layer2_outputs(6337)) and not (layer2_outputs(4517));
    layer3_outputs(3737) <= (layer2_outputs(3334)) and (layer2_outputs(2182));
    layer3_outputs(3738) <= (layer2_outputs(2036)) and not (layer2_outputs(6425));
    layer3_outputs(3739) <= not(layer2_outputs(4386)) or (layer2_outputs(2815));
    layer3_outputs(3740) <= (layer2_outputs(2180)) xor (layer2_outputs(2316));
    layer3_outputs(3741) <= (layer2_outputs(1890)) and not (layer2_outputs(1121));
    layer3_outputs(3742) <= (layer2_outputs(662)) and not (layer2_outputs(6069));
    layer3_outputs(3743) <= (layer2_outputs(469)) and not (layer2_outputs(1628));
    layer3_outputs(3744) <= (layer2_outputs(5142)) and not (layer2_outputs(3654));
    layer3_outputs(3745) <= (layer2_outputs(5701)) and (layer2_outputs(4068));
    layer3_outputs(3746) <= (layer2_outputs(2675)) and not (layer2_outputs(2137));
    layer3_outputs(3747) <= layer2_outputs(2923);
    layer3_outputs(3748) <= not(layer2_outputs(4866)) or (layer2_outputs(7024));
    layer3_outputs(3749) <= not((layer2_outputs(4948)) and (layer2_outputs(5137)));
    layer3_outputs(3750) <= layer2_outputs(6247);
    layer3_outputs(3751) <= not(layer2_outputs(6359));
    layer3_outputs(3752) <= not(layer2_outputs(6228));
    layer3_outputs(3753) <= (layer2_outputs(3269)) and (layer2_outputs(6055));
    layer3_outputs(3754) <= layer2_outputs(4644);
    layer3_outputs(3755) <= layer2_outputs(3160);
    layer3_outputs(3756) <= layer2_outputs(526);
    layer3_outputs(3757) <= '0';
    layer3_outputs(3758) <= (layer2_outputs(2173)) xor (layer2_outputs(1353));
    layer3_outputs(3759) <= (layer2_outputs(1498)) and not (layer2_outputs(1553));
    layer3_outputs(3760) <= (layer2_outputs(1786)) xor (layer2_outputs(739));
    layer3_outputs(3761) <= not(layer2_outputs(7192)) or (layer2_outputs(3289));
    layer3_outputs(3762) <= not((layer2_outputs(5179)) or (layer2_outputs(5310)));
    layer3_outputs(3763) <= layer2_outputs(1588);
    layer3_outputs(3764) <= not(layer2_outputs(1510)) or (layer2_outputs(4019));
    layer3_outputs(3765) <= not((layer2_outputs(728)) and (layer2_outputs(7052)));
    layer3_outputs(3766) <= not(layer2_outputs(5377));
    layer3_outputs(3767) <= not((layer2_outputs(942)) or (layer2_outputs(2391)));
    layer3_outputs(3768) <= layer2_outputs(521);
    layer3_outputs(3769) <= (layer2_outputs(5148)) and not (layer2_outputs(6937));
    layer3_outputs(3770) <= (layer2_outputs(6484)) or (layer2_outputs(2668));
    layer3_outputs(3771) <= layer2_outputs(232);
    layer3_outputs(3772) <= '0';
    layer3_outputs(3773) <= not(layer2_outputs(7244));
    layer3_outputs(3774) <= layer2_outputs(2801);
    layer3_outputs(3775) <= not(layer2_outputs(850));
    layer3_outputs(3776) <= layer2_outputs(140);
    layer3_outputs(3777) <= not(layer2_outputs(2466)) or (layer2_outputs(3573));
    layer3_outputs(3778) <= layer2_outputs(2546);
    layer3_outputs(3779) <= (layer2_outputs(2215)) or (layer2_outputs(3535));
    layer3_outputs(3780) <= (layer2_outputs(3134)) and not (layer2_outputs(5359));
    layer3_outputs(3781) <= layer2_outputs(7638);
    layer3_outputs(3782) <= (layer2_outputs(1231)) and not (layer2_outputs(3490));
    layer3_outputs(3783) <= not(layer2_outputs(53)) or (layer2_outputs(2640));
    layer3_outputs(3784) <= (layer2_outputs(3666)) and not (layer2_outputs(2862));
    layer3_outputs(3785) <= not((layer2_outputs(6576)) or (layer2_outputs(6143)));
    layer3_outputs(3786) <= not(layer2_outputs(3440)) or (layer2_outputs(6215));
    layer3_outputs(3787) <= not((layer2_outputs(2527)) and (layer2_outputs(3259)));
    layer3_outputs(3788) <= '0';
    layer3_outputs(3789) <= not(layer2_outputs(6619));
    layer3_outputs(3790) <= (layer2_outputs(4107)) and not (layer2_outputs(5562));
    layer3_outputs(3791) <= '0';
    layer3_outputs(3792) <= (layer2_outputs(2641)) and not (layer2_outputs(1452));
    layer3_outputs(3793) <= not(layer2_outputs(2919));
    layer3_outputs(3794) <= layer2_outputs(277);
    layer3_outputs(3795) <= not(layer2_outputs(6422)) or (layer2_outputs(1054));
    layer3_outputs(3796) <= (layer2_outputs(7233)) and not (layer2_outputs(4894));
    layer3_outputs(3797) <= not(layer2_outputs(3883));
    layer3_outputs(3798) <= layer2_outputs(7268);
    layer3_outputs(3799) <= '1';
    layer3_outputs(3800) <= not(layer2_outputs(6847));
    layer3_outputs(3801) <= layer2_outputs(6524);
    layer3_outputs(3802) <= (layer2_outputs(6907)) xor (layer2_outputs(6191));
    layer3_outputs(3803) <= layer2_outputs(2924);
    layer3_outputs(3804) <= (layer2_outputs(788)) and not (layer2_outputs(2748));
    layer3_outputs(3805) <= (layer2_outputs(3198)) and not (layer2_outputs(4053));
    layer3_outputs(3806) <= '0';
    layer3_outputs(3807) <= layer2_outputs(3169);
    layer3_outputs(3808) <= (layer2_outputs(3112)) and not (layer2_outputs(5278));
    layer3_outputs(3809) <= not(layer2_outputs(4989)) or (layer2_outputs(6911));
    layer3_outputs(3810) <= (layer2_outputs(3229)) and not (layer2_outputs(6389));
    layer3_outputs(3811) <= (layer2_outputs(3457)) or (layer2_outputs(403));
    layer3_outputs(3812) <= layer2_outputs(770);
    layer3_outputs(3813) <= layer2_outputs(2689);
    layer3_outputs(3814) <= layer2_outputs(514);
    layer3_outputs(3815) <= not(layer2_outputs(4529));
    layer3_outputs(3816) <= (layer2_outputs(6366)) and not (layer2_outputs(4641));
    layer3_outputs(3817) <= not((layer2_outputs(5606)) xor (layer2_outputs(868)));
    layer3_outputs(3818) <= (layer2_outputs(44)) and not (layer2_outputs(1805));
    layer3_outputs(3819) <= not((layer2_outputs(4290)) and (layer2_outputs(7160)));
    layer3_outputs(3820) <= (layer2_outputs(2683)) or (layer2_outputs(1339));
    layer3_outputs(3821) <= layer2_outputs(7312);
    layer3_outputs(3822) <= not(layer2_outputs(2010));
    layer3_outputs(3823) <= '1';
    layer3_outputs(3824) <= layer2_outputs(6649);
    layer3_outputs(3825) <= not(layer2_outputs(5803));
    layer3_outputs(3826) <= not(layer2_outputs(6291));
    layer3_outputs(3827) <= (layer2_outputs(6052)) or (layer2_outputs(2957));
    layer3_outputs(3828) <= (layer2_outputs(5796)) and not (layer2_outputs(5751));
    layer3_outputs(3829) <= not(layer2_outputs(921)) or (layer2_outputs(6186));
    layer3_outputs(3830) <= (layer2_outputs(509)) and not (layer2_outputs(1450));
    layer3_outputs(3831) <= '1';
    layer3_outputs(3832) <= '1';
    layer3_outputs(3833) <= not((layer2_outputs(2776)) xor (layer2_outputs(2160)));
    layer3_outputs(3834) <= not((layer2_outputs(1443)) xor (layer2_outputs(2296)));
    layer3_outputs(3835) <= (layer2_outputs(4388)) xor (layer2_outputs(4091));
    layer3_outputs(3836) <= '1';
    layer3_outputs(3837) <= not(layer2_outputs(5061)) or (layer2_outputs(4314));
    layer3_outputs(3838) <= not(layer2_outputs(642));
    layer3_outputs(3839) <= (layer2_outputs(5792)) or (layer2_outputs(7291));
    layer3_outputs(3840) <= not((layer2_outputs(1499)) or (layer2_outputs(21)));
    layer3_outputs(3841) <= not((layer2_outputs(5297)) and (layer2_outputs(1734)));
    layer3_outputs(3842) <= layer2_outputs(1812);
    layer3_outputs(3843) <= not(layer2_outputs(3380)) or (layer2_outputs(7666));
    layer3_outputs(3844) <= not(layer2_outputs(1872));
    layer3_outputs(3845) <= '1';
    layer3_outputs(3846) <= not(layer2_outputs(794)) or (layer2_outputs(2921));
    layer3_outputs(3847) <= not((layer2_outputs(2139)) xor (layer2_outputs(4635)));
    layer3_outputs(3848) <= not((layer2_outputs(114)) xor (layer2_outputs(4329)));
    layer3_outputs(3849) <= not(layer2_outputs(354));
    layer3_outputs(3850) <= (layer2_outputs(2746)) and not (layer2_outputs(3916));
    layer3_outputs(3851) <= (layer2_outputs(6455)) and not (layer2_outputs(5362));
    layer3_outputs(3852) <= not(layer2_outputs(4598));
    layer3_outputs(3853) <= layer2_outputs(6000);
    layer3_outputs(3854) <= layer2_outputs(6507);
    layer3_outputs(3855) <= (layer2_outputs(7614)) xor (layer2_outputs(5802));
    layer3_outputs(3856) <= layer2_outputs(3553);
    layer3_outputs(3857) <= (layer2_outputs(7070)) xor (layer2_outputs(5799));
    layer3_outputs(3858) <= not(layer2_outputs(174)) or (layer2_outputs(363));
    layer3_outputs(3859) <= (layer2_outputs(2143)) and not (layer2_outputs(2316));
    layer3_outputs(3860) <= not(layer2_outputs(575));
    layer3_outputs(3861) <= (layer2_outputs(227)) and (layer2_outputs(3680));
    layer3_outputs(3862) <= (layer2_outputs(6689)) and (layer2_outputs(1220));
    layer3_outputs(3863) <= '1';
    layer3_outputs(3864) <= layer2_outputs(4312);
    layer3_outputs(3865) <= not((layer2_outputs(3022)) and (layer2_outputs(252)));
    layer3_outputs(3866) <= not((layer2_outputs(6204)) or (layer2_outputs(566)));
    layer3_outputs(3867) <= not(layer2_outputs(274)) or (layer2_outputs(6975));
    layer3_outputs(3868) <= not(layer2_outputs(4049));
    layer3_outputs(3869) <= not((layer2_outputs(7576)) xor (layer2_outputs(5408)));
    layer3_outputs(3870) <= not(layer2_outputs(6643));
    layer3_outputs(3871) <= (layer2_outputs(2062)) and not (layer2_outputs(2053));
    layer3_outputs(3872) <= not((layer2_outputs(2267)) or (layer2_outputs(4245)));
    layer3_outputs(3873) <= not(layer2_outputs(4201)) or (layer2_outputs(3528));
    layer3_outputs(3874) <= not((layer2_outputs(7464)) and (layer2_outputs(5271)));
    layer3_outputs(3875) <= not(layer2_outputs(627));
    layer3_outputs(3876) <= not((layer2_outputs(1974)) and (layer2_outputs(7445)));
    layer3_outputs(3877) <= (layer2_outputs(4405)) or (layer2_outputs(1667));
    layer3_outputs(3878) <= layer2_outputs(2234);
    layer3_outputs(3879) <= (layer2_outputs(4769)) xor (layer2_outputs(2036));
    layer3_outputs(3880) <= not((layer2_outputs(2761)) or (layer2_outputs(5893)));
    layer3_outputs(3881) <= '0';
    layer3_outputs(3882) <= not((layer2_outputs(2702)) xor (layer2_outputs(4470)));
    layer3_outputs(3883) <= not(layer2_outputs(4631)) or (layer2_outputs(1320));
    layer3_outputs(3884) <= (layer2_outputs(4320)) and (layer2_outputs(3421));
    layer3_outputs(3885) <= (layer2_outputs(3389)) and (layer2_outputs(946));
    layer3_outputs(3886) <= layer2_outputs(6753);
    layer3_outputs(3887) <= '1';
    layer3_outputs(3888) <= (layer2_outputs(1079)) and not (layer2_outputs(429));
    layer3_outputs(3889) <= layer2_outputs(2463);
    layer3_outputs(3890) <= not(layer2_outputs(2807));
    layer3_outputs(3891) <= (layer2_outputs(6828)) and (layer2_outputs(883));
    layer3_outputs(3892) <= not((layer2_outputs(1960)) and (layer2_outputs(3883)));
    layer3_outputs(3893) <= not((layer2_outputs(616)) or (layer2_outputs(4928)));
    layer3_outputs(3894) <= '0';
    layer3_outputs(3895) <= '0';
    layer3_outputs(3896) <= '1';
    layer3_outputs(3897) <= not((layer2_outputs(3859)) or (layer2_outputs(6028)));
    layer3_outputs(3898) <= not((layer2_outputs(7543)) and (layer2_outputs(4739)));
    layer3_outputs(3899) <= (layer2_outputs(1082)) and not (layer2_outputs(6077));
    layer3_outputs(3900) <= not((layer2_outputs(4530)) or (layer2_outputs(700)));
    layer3_outputs(3901) <= not((layer2_outputs(4977)) and (layer2_outputs(2103)));
    layer3_outputs(3902) <= not((layer2_outputs(615)) or (layer2_outputs(91)));
    layer3_outputs(3903) <= '0';
    layer3_outputs(3904) <= layer2_outputs(2179);
    layer3_outputs(3905) <= layer2_outputs(551);
    layer3_outputs(3906) <= not(layer2_outputs(1475));
    layer3_outputs(3907) <= not(layer2_outputs(604));
    layer3_outputs(3908) <= not(layer2_outputs(5788)) or (layer2_outputs(2970));
    layer3_outputs(3909) <= not((layer2_outputs(1008)) or (layer2_outputs(7548)));
    layer3_outputs(3910) <= not(layer2_outputs(6123)) or (layer2_outputs(5592));
    layer3_outputs(3911) <= not(layer2_outputs(3335)) or (layer2_outputs(7375));
    layer3_outputs(3912) <= (layer2_outputs(1352)) and not (layer2_outputs(3459));
    layer3_outputs(3913) <= not(layer2_outputs(5369)) or (layer2_outputs(1575));
    layer3_outputs(3914) <= not(layer2_outputs(7128));
    layer3_outputs(3915) <= not(layer2_outputs(5325));
    layer3_outputs(3916) <= not(layer2_outputs(3842));
    layer3_outputs(3917) <= (layer2_outputs(2126)) and not (layer2_outputs(6602));
    layer3_outputs(3918) <= not(layer2_outputs(7482)) or (layer2_outputs(3766));
    layer3_outputs(3919) <= not((layer2_outputs(4109)) and (layer2_outputs(4195)));
    layer3_outputs(3920) <= not(layer2_outputs(606)) or (layer2_outputs(6038));
    layer3_outputs(3921) <= not((layer2_outputs(3447)) or (layer2_outputs(5068)));
    layer3_outputs(3922) <= not(layer2_outputs(7057));
    layer3_outputs(3923) <= not(layer2_outputs(1504));
    layer3_outputs(3924) <= not((layer2_outputs(3012)) and (layer2_outputs(511)));
    layer3_outputs(3925) <= (layer2_outputs(2596)) or (layer2_outputs(5774));
    layer3_outputs(3926) <= layer2_outputs(374);
    layer3_outputs(3927) <= (layer2_outputs(608)) xor (layer2_outputs(6943));
    layer3_outputs(3928) <= not((layer2_outputs(2117)) and (layer2_outputs(4686)));
    layer3_outputs(3929) <= layer2_outputs(6158);
    layer3_outputs(3930) <= (layer2_outputs(2782)) and not (layer2_outputs(1116));
    layer3_outputs(3931) <= (layer2_outputs(6308)) or (layer2_outputs(4966));
    layer3_outputs(3932) <= not(layer2_outputs(1922));
    layer3_outputs(3933) <= not(layer2_outputs(5685));
    layer3_outputs(3934) <= (layer2_outputs(2539)) or (layer2_outputs(1593));
    layer3_outputs(3935) <= layer2_outputs(1265);
    layer3_outputs(3936) <= layer2_outputs(1379);
    layer3_outputs(3937) <= not(layer2_outputs(3264));
    layer3_outputs(3938) <= (layer2_outputs(146)) and not (layer2_outputs(5948));
    layer3_outputs(3939) <= (layer2_outputs(6710)) and not (layer2_outputs(5561));
    layer3_outputs(3940) <= layer2_outputs(449);
    layer3_outputs(3941) <= not((layer2_outputs(5145)) and (layer2_outputs(1959)));
    layer3_outputs(3942) <= not((layer2_outputs(4764)) or (layer2_outputs(3099)));
    layer3_outputs(3943) <= (layer2_outputs(6520)) or (layer2_outputs(3955));
    layer3_outputs(3944) <= layer2_outputs(6137);
    layer3_outputs(3945) <= layer2_outputs(3547);
    layer3_outputs(3946) <= (layer2_outputs(1481)) and (layer2_outputs(3578));
    layer3_outputs(3947) <= (layer2_outputs(6738)) and not (layer2_outputs(4553));
    layer3_outputs(3948) <= not(layer2_outputs(3636));
    layer3_outputs(3949) <= not(layer2_outputs(4787));
    layer3_outputs(3950) <= not(layer2_outputs(929)) or (layer2_outputs(6100));
    layer3_outputs(3951) <= (layer2_outputs(4498)) and not (layer2_outputs(1314));
    layer3_outputs(3952) <= not(layer2_outputs(5405));
    layer3_outputs(3953) <= layer2_outputs(3622);
    layer3_outputs(3954) <= '1';
    layer3_outputs(3955) <= not(layer2_outputs(2489)) or (layer2_outputs(6182));
    layer3_outputs(3956) <= not((layer2_outputs(7239)) and (layer2_outputs(784)));
    layer3_outputs(3957) <= layer2_outputs(6937);
    layer3_outputs(3958) <= not((layer2_outputs(5648)) or (layer2_outputs(77)));
    layer3_outputs(3959) <= layer2_outputs(6995);
    layer3_outputs(3960) <= (layer2_outputs(5376)) and (layer2_outputs(5483));
    layer3_outputs(3961) <= (layer2_outputs(1776)) and not (layer2_outputs(6192));
    layer3_outputs(3962) <= not(layer2_outputs(3444)) or (layer2_outputs(3453));
    layer3_outputs(3963) <= not((layer2_outputs(1764)) and (layer2_outputs(7206)));
    layer3_outputs(3964) <= not((layer2_outputs(2825)) and (layer2_outputs(3951)));
    layer3_outputs(3965) <= '0';
    layer3_outputs(3966) <= (layer2_outputs(7096)) and not (layer2_outputs(7212));
    layer3_outputs(3967) <= layer2_outputs(4938);
    layer3_outputs(3968) <= layer2_outputs(5923);
    layer3_outputs(3969) <= '1';
    layer3_outputs(3970) <= (layer2_outputs(1040)) and (layer2_outputs(3544));
    layer3_outputs(3971) <= not(layer2_outputs(3395)) or (layer2_outputs(7160));
    layer3_outputs(3972) <= not(layer2_outputs(3985)) or (layer2_outputs(7303));
    layer3_outputs(3973) <= (layer2_outputs(5266)) and (layer2_outputs(2462));
    layer3_outputs(3974) <= '1';
    layer3_outputs(3975) <= layer2_outputs(7515);
    layer3_outputs(3976) <= (layer2_outputs(5833)) or (layer2_outputs(5898));
    layer3_outputs(3977) <= layer2_outputs(4657);
    layer3_outputs(3978) <= not((layer2_outputs(4339)) or (layer2_outputs(2715)));
    layer3_outputs(3979) <= (layer2_outputs(1161)) xor (layer2_outputs(1202));
    layer3_outputs(3980) <= (layer2_outputs(781)) xor (layer2_outputs(4623));
    layer3_outputs(3981) <= (layer2_outputs(3684)) and (layer2_outputs(5241));
    layer3_outputs(3982) <= not(layer2_outputs(6916));
    layer3_outputs(3983) <= layer2_outputs(2853);
    layer3_outputs(3984) <= layer2_outputs(5706);
    layer3_outputs(3985) <= (layer2_outputs(2404)) and (layer2_outputs(1986));
    layer3_outputs(3986) <= not(layer2_outputs(5621)) or (layer2_outputs(7230));
    layer3_outputs(3987) <= not((layer2_outputs(4480)) or (layer2_outputs(1988)));
    layer3_outputs(3988) <= not((layer2_outputs(6057)) or (layer2_outputs(917)));
    layer3_outputs(3989) <= not(layer2_outputs(4744));
    layer3_outputs(3990) <= not(layer2_outputs(2989)) or (layer2_outputs(882));
    layer3_outputs(3991) <= not(layer2_outputs(4486));
    layer3_outputs(3992) <= (layer2_outputs(5973)) or (layer2_outputs(7138));
    layer3_outputs(3993) <= layer2_outputs(6276);
    layer3_outputs(3994) <= (layer2_outputs(3286)) and not (layer2_outputs(6651));
    layer3_outputs(3995) <= (layer2_outputs(1562)) and (layer2_outputs(1053));
    layer3_outputs(3996) <= not((layer2_outputs(7440)) or (layer2_outputs(1907)));
    layer3_outputs(3997) <= (layer2_outputs(3557)) and not (layer2_outputs(328));
    layer3_outputs(3998) <= not((layer2_outputs(1809)) and (layer2_outputs(2059)));
    layer3_outputs(3999) <= layer2_outputs(2646);
    layer3_outputs(4000) <= not(layer2_outputs(4529));
    layer3_outputs(4001) <= not((layer2_outputs(2304)) and (layer2_outputs(7178)));
    layer3_outputs(4002) <= (layer2_outputs(5685)) and not (layer2_outputs(2482));
    layer3_outputs(4003) <= layer2_outputs(7050);
    layer3_outputs(4004) <= not((layer2_outputs(1599)) or (layer2_outputs(3417)));
    layer3_outputs(4005) <= not(layer2_outputs(5548)) or (layer2_outputs(3133));
    layer3_outputs(4006) <= layer2_outputs(6868);
    layer3_outputs(4007) <= (layer2_outputs(4423)) or (layer2_outputs(1507));
    layer3_outputs(4008) <= not(layer2_outputs(5324));
    layer3_outputs(4009) <= '0';
    layer3_outputs(4010) <= layer2_outputs(4901);
    layer3_outputs(4011) <= layer2_outputs(4048);
    layer3_outputs(4012) <= not((layer2_outputs(6704)) or (layer2_outputs(2512)));
    layer3_outputs(4013) <= (layer2_outputs(6625)) xor (layer2_outputs(1426));
    layer3_outputs(4014) <= not((layer2_outputs(859)) and (layer2_outputs(3898)));
    layer3_outputs(4015) <= not(layer2_outputs(2912));
    layer3_outputs(4016) <= not(layer2_outputs(3931));
    layer3_outputs(4017) <= not(layer2_outputs(6522));
    layer3_outputs(4018) <= not(layer2_outputs(4194)) or (layer2_outputs(3098));
    layer3_outputs(4019) <= layer2_outputs(386);
    layer3_outputs(4020) <= not(layer2_outputs(3093));
    layer3_outputs(4021) <= (layer2_outputs(1469)) xor (layer2_outputs(7422));
    layer3_outputs(4022) <= (layer2_outputs(6045)) or (layer2_outputs(432));
    layer3_outputs(4023) <= layer2_outputs(1238);
    layer3_outputs(4024) <= not(layer2_outputs(5845)) or (layer2_outputs(1914));
    layer3_outputs(4025) <= not(layer2_outputs(6800));
    layer3_outputs(4026) <= layer2_outputs(4673);
    layer3_outputs(4027) <= layer2_outputs(2453);
    layer3_outputs(4028) <= (layer2_outputs(1374)) and (layer2_outputs(6400));
    layer3_outputs(4029) <= not(layer2_outputs(2678)) or (layer2_outputs(5237));
    layer3_outputs(4030) <= not(layer2_outputs(845)) or (layer2_outputs(2429));
    layer3_outputs(4031) <= layer2_outputs(6722);
    layer3_outputs(4032) <= '1';
    layer3_outputs(4033) <= '0';
    layer3_outputs(4034) <= not((layer2_outputs(585)) xor (layer2_outputs(491)));
    layer3_outputs(4035) <= layer2_outputs(4065);
    layer3_outputs(4036) <= '0';
    layer3_outputs(4037) <= layer2_outputs(4937);
    layer3_outputs(4038) <= not((layer2_outputs(7274)) or (layer2_outputs(1951)));
    layer3_outputs(4039) <= '0';
    layer3_outputs(4040) <= (layer2_outputs(1203)) and not (layer2_outputs(2698));
    layer3_outputs(4041) <= (layer2_outputs(6879)) and not (layer2_outputs(2377));
    layer3_outputs(4042) <= layer2_outputs(198);
    layer3_outputs(4043) <= (layer2_outputs(5850)) xor (layer2_outputs(5581));
    layer3_outputs(4044) <= (layer2_outputs(6083)) and (layer2_outputs(6962));
    layer3_outputs(4045) <= layer2_outputs(6801);
    layer3_outputs(4046) <= (layer2_outputs(6381)) and not (layer2_outputs(808));
    layer3_outputs(4047) <= (layer2_outputs(1997)) xor (layer2_outputs(1300));
    layer3_outputs(4048) <= (layer2_outputs(6727)) or (layer2_outputs(2771));
    layer3_outputs(4049) <= not(layer2_outputs(4873)) or (layer2_outputs(2287));
    layer3_outputs(4050) <= not(layer2_outputs(3677)) or (layer2_outputs(6476));
    layer3_outputs(4051) <= not(layer2_outputs(6759));
    layer3_outputs(4052) <= (layer2_outputs(6294)) and not (layer2_outputs(1421));
    layer3_outputs(4053) <= not(layer2_outputs(4890));
    layer3_outputs(4054) <= not((layer2_outputs(1929)) and (layer2_outputs(5416)));
    layer3_outputs(4055) <= (layer2_outputs(5581)) or (layer2_outputs(3697));
    layer3_outputs(4056) <= (layer2_outputs(5198)) and not (layer2_outputs(6985));
    layer3_outputs(4057) <= not(layer2_outputs(6434));
    layer3_outputs(4058) <= (layer2_outputs(4288)) and (layer2_outputs(2046));
    layer3_outputs(4059) <= (layer2_outputs(6300)) and not (layer2_outputs(5166));
    layer3_outputs(4060) <= not(layer2_outputs(1771));
    layer3_outputs(4061) <= (layer2_outputs(1741)) or (layer2_outputs(7427));
    layer3_outputs(4062) <= (layer2_outputs(7495)) and (layer2_outputs(6218));
    layer3_outputs(4063) <= not((layer2_outputs(3360)) and (layer2_outputs(5352)));
    layer3_outputs(4064) <= (layer2_outputs(5719)) and (layer2_outputs(1106));
    layer3_outputs(4065) <= layer2_outputs(4737);
    layer3_outputs(4066) <= layer2_outputs(1020);
    layer3_outputs(4067) <= '1';
    layer3_outputs(4068) <= (layer2_outputs(2823)) and not (layer2_outputs(4578));
    layer3_outputs(4069) <= not((layer2_outputs(6752)) xor (layer2_outputs(6832)));
    layer3_outputs(4070) <= not(layer2_outputs(4771)) or (layer2_outputs(7015));
    layer3_outputs(4071) <= (layer2_outputs(6614)) and not (layer2_outputs(821));
    layer3_outputs(4072) <= layer2_outputs(1920);
    layer3_outputs(4073) <= '0';
    layer3_outputs(4074) <= not(layer2_outputs(5548)) or (layer2_outputs(6808));
    layer3_outputs(4075) <= not(layer2_outputs(5535)) or (layer2_outputs(5025));
    layer3_outputs(4076) <= not(layer2_outputs(886)) or (layer2_outputs(6020));
    layer3_outputs(4077) <= not((layer2_outputs(5349)) or (layer2_outputs(5819)));
    layer3_outputs(4078) <= not(layer2_outputs(846)) or (layer2_outputs(6475));
    layer3_outputs(4079) <= not(layer2_outputs(7567));
    layer3_outputs(4080) <= layer2_outputs(6099);
    layer3_outputs(4081) <= layer2_outputs(6861);
    layer3_outputs(4082) <= not(layer2_outputs(1388));
    layer3_outputs(4083) <= not((layer2_outputs(5026)) xor (layer2_outputs(6783)));
    layer3_outputs(4084) <= (layer2_outputs(255)) or (layer2_outputs(839));
    layer3_outputs(4085) <= not((layer2_outputs(6115)) xor (layer2_outputs(5075)));
    layer3_outputs(4086) <= not(layer2_outputs(337));
    layer3_outputs(4087) <= not((layer2_outputs(973)) and (layer2_outputs(6883)));
    layer3_outputs(4088) <= (layer2_outputs(184)) or (layer2_outputs(2046));
    layer3_outputs(4089) <= layer2_outputs(7356);
    layer3_outputs(4090) <= (layer2_outputs(4027)) and not (layer2_outputs(6166));
    layer3_outputs(4091) <= (layer2_outputs(6466)) and not (layer2_outputs(786));
    layer3_outputs(4092) <= (layer2_outputs(3211)) or (layer2_outputs(4311));
    layer3_outputs(4093) <= layer2_outputs(5082);
    layer3_outputs(4094) <= layer2_outputs(2792);
    layer3_outputs(4095) <= layer2_outputs(4921);
    layer3_outputs(4096) <= not((layer2_outputs(3057)) xor (layer2_outputs(4655)));
    layer3_outputs(4097) <= layer2_outputs(2159);
    layer3_outputs(4098) <= (layer2_outputs(3882)) or (layer2_outputs(7188));
    layer3_outputs(4099) <= '0';
    layer3_outputs(4100) <= not(layer2_outputs(3269));
    layer3_outputs(4101) <= '1';
    layer3_outputs(4102) <= '0';
    layer3_outputs(4103) <= not((layer2_outputs(7639)) and (layer2_outputs(4616)));
    layer3_outputs(4104) <= (layer2_outputs(1276)) and not (layer2_outputs(2654));
    layer3_outputs(4105) <= not((layer2_outputs(5654)) or (layer2_outputs(4556)));
    layer3_outputs(4106) <= (layer2_outputs(2796)) or (layer2_outputs(4461));
    layer3_outputs(4107) <= (layer2_outputs(4163)) or (layer2_outputs(2253));
    layer3_outputs(4108) <= not(layer2_outputs(6537)) or (layer2_outputs(982));
    layer3_outputs(4109) <= not(layer2_outputs(1273)) or (layer2_outputs(2850));
    layer3_outputs(4110) <= layer2_outputs(7004);
    layer3_outputs(4111) <= not((layer2_outputs(1270)) or (layer2_outputs(2759)));
    layer3_outputs(4112) <= not(layer2_outputs(5760));
    layer3_outputs(4113) <= not(layer2_outputs(5652));
    layer3_outputs(4114) <= not((layer2_outputs(4732)) or (layer2_outputs(7276)));
    layer3_outputs(4115) <= (layer2_outputs(5887)) xor (layer2_outputs(5999));
    layer3_outputs(4116) <= not(layer2_outputs(1646));
    layer3_outputs(4117) <= layer2_outputs(2795);
    layer3_outputs(4118) <= not((layer2_outputs(6932)) or (layer2_outputs(3128)));
    layer3_outputs(4119) <= layer2_outputs(1245);
    layer3_outputs(4120) <= not(layer2_outputs(2672));
    layer3_outputs(4121) <= '1';
    layer3_outputs(4122) <= layer2_outputs(5387);
    layer3_outputs(4123) <= '0';
    layer3_outputs(4124) <= (layer2_outputs(2198)) and (layer2_outputs(7110));
    layer3_outputs(4125) <= not(layer2_outputs(4260));
    layer3_outputs(4126) <= (layer2_outputs(4705)) and not (layer2_outputs(831));
    layer3_outputs(4127) <= layer2_outputs(103);
    layer3_outputs(4128) <= not(layer2_outputs(221));
    layer3_outputs(4129) <= not((layer2_outputs(3812)) and (layer2_outputs(2667)));
    layer3_outputs(4130) <= not(layer2_outputs(266));
    layer3_outputs(4131) <= layer2_outputs(6870);
    layer3_outputs(4132) <= layer2_outputs(7478);
    layer3_outputs(4133) <= '1';
    layer3_outputs(4134) <= (layer2_outputs(5461)) or (layer2_outputs(5998));
    layer3_outputs(4135) <= not((layer2_outputs(468)) or (layer2_outputs(4918)));
    layer3_outputs(4136) <= '0';
    layer3_outputs(4137) <= (layer2_outputs(7491)) and not (layer2_outputs(3073));
    layer3_outputs(4138) <= (layer2_outputs(2008)) and (layer2_outputs(2399));
    layer3_outputs(4139) <= not(layer2_outputs(4904));
    layer3_outputs(4140) <= (layer2_outputs(1181)) or (layer2_outputs(1787));
    layer3_outputs(4141) <= not((layer2_outputs(4276)) and (layer2_outputs(907)));
    layer3_outputs(4142) <= layer2_outputs(6719);
    layer3_outputs(4143) <= not(layer2_outputs(7294));
    layer3_outputs(4144) <= (layer2_outputs(3902)) and not (layer2_outputs(6222));
    layer3_outputs(4145) <= layer2_outputs(637);
    layer3_outputs(4146) <= '1';
    layer3_outputs(4147) <= not(layer2_outputs(6908));
    layer3_outputs(4148) <= (layer2_outputs(75)) xor (layer2_outputs(4251));
    layer3_outputs(4149) <= not((layer2_outputs(6699)) and (layer2_outputs(3213)));
    layer3_outputs(4150) <= not(layer2_outputs(3441)) or (layer2_outputs(3970));
    layer3_outputs(4151) <= not((layer2_outputs(4876)) and (layer2_outputs(5552)));
    layer3_outputs(4152) <= not(layer2_outputs(5009)) or (layer2_outputs(231));
    layer3_outputs(4153) <= not((layer2_outputs(7034)) or (layer2_outputs(1825)));
    layer3_outputs(4154) <= not(layer2_outputs(2326));
    layer3_outputs(4155) <= not((layer2_outputs(1198)) and (layer2_outputs(5382)));
    layer3_outputs(4156) <= '0';
    layer3_outputs(4157) <= layer2_outputs(2269);
    layer3_outputs(4158) <= layer2_outputs(638);
    layer3_outputs(4159) <= layer2_outputs(7172);
    layer3_outputs(4160) <= not(layer2_outputs(6543));
    layer3_outputs(4161) <= (layer2_outputs(4)) and not (layer2_outputs(5837));
    layer3_outputs(4162) <= not((layer2_outputs(1618)) and (layer2_outputs(6310)));
    layer3_outputs(4163) <= not((layer2_outputs(665)) or (layer2_outputs(5100)));
    layer3_outputs(4164) <= (layer2_outputs(3886)) or (layer2_outputs(4114));
    layer3_outputs(4165) <= not((layer2_outputs(1807)) and (layer2_outputs(6213)));
    layer3_outputs(4166) <= '0';
    layer3_outputs(4167) <= (layer2_outputs(1458)) and not (layer2_outputs(7313));
    layer3_outputs(4168) <= (layer2_outputs(175)) and not (layer2_outputs(5281));
    layer3_outputs(4169) <= '1';
    layer3_outputs(4170) <= '1';
    layer3_outputs(4171) <= (layer2_outputs(3676)) and not (layer2_outputs(2769));
    layer3_outputs(4172) <= not((layer2_outputs(6009)) and (layer2_outputs(1900)));
    layer3_outputs(4173) <= (layer2_outputs(5094)) xor (layer2_outputs(921));
    layer3_outputs(4174) <= (layer2_outputs(2937)) xor (layer2_outputs(2565));
    layer3_outputs(4175) <= not((layer2_outputs(1599)) or (layer2_outputs(1877)));
    layer3_outputs(4176) <= not(layer2_outputs(5106));
    layer3_outputs(4177) <= not(layer2_outputs(3179)) or (layer2_outputs(5684));
    layer3_outputs(4178) <= not(layer2_outputs(3945)) or (layer2_outputs(2098));
    layer3_outputs(4179) <= not(layer2_outputs(3472)) or (layer2_outputs(5856));
    layer3_outputs(4180) <= not(layer2_outputs(6145));
    layer3_outputs(4181) <= (layer2_outputs(2304)) or (layer2_outputs(815));
    layer3_outputs(4182) <= not(layer2_outputs(1382));
    layer3_outputs(4183) <= '1';
    layer3_outputs(4184) <= '0';
    layer3_outputs(4185) <= not((layer2_outputs(3275)) and (layer2_outputs(1957)));
    layer3_outputs(4186) <= not(layer2_outputs(478));
    layer3_outputs(4187) <= not((layer2_outputs(5092)) and (layer2_outputs(7136)));
    layer3_outputs(4188) <= not((layer2_outputs(2633)) or (layer2_outputs(5358)));
    layer3_outputs(4189) <= '1';
    layer3_outputs(4190) <= not((layer2_outputs(3094)) or (layer2_outputs(3873)));
    layer3_outputs(4191) <= not(layer2_outputs(4495));
    layer3_outputs(4192) <= not(layer2_outputs(2978));
    layer3_outputs(4193) <= (layer2_outputs(3518)) or (layer2_outputs(4238));
    layer3_outputs(4194) <= not(layer2_outputs(7278));
    layer3_outputs(4195) <= layer2_outputs(2344);
    layer3_outputs(4196) <= (layer2_outputs(6966)) and not (layer2_outputs(7446));
    layer3_outputs(4197) <= layer2_outputs(4326);
    layer3_outputs(4198) <= not(layer2_outputs(3374)) or (layer2_outputs(7213));
    layer3_outputs(4199) <= not(layer2_outputs(2639));
    layer3_outputs(4200) <= not((layer2_outputs(1765)) or (layer2_outputs(6752)));
    layer3_outputs(4201) <= not(layer2_outputs(4336));
    layer3_outputs(4202) <= layer2_outputs(4583);
    layer3_outputs(4203) <= (layer2_outputs(3919)) and not (layer2_outputs(691));
    layer3_outputs(4204) <= not(layer2_outputs(450)) or (layer2_outputs(2383));
    layer3_outputs(4205) <= not((layer2_outputs(2335)) or (layer2_outputs(719)));
    layer3_outputs(4206) <= layer2_outputs(4797);
    layer3_outputs(4207) <= not(layer2_outputs(887));
    layer3_outputs(4208) <= layer2_outputs(292);
    layer3_outputs(4209) <= not(layer2_outputs(5038)) or (layer2_outputs(7100));
    layer3_outputs(4210) <= not(layer2_outputs(3115)) or (layer2_outputs(4613));
    layer3_outputs(4211) <= layer2_outputs(6927);
    layer3_outputs(4212) <= '0';
    layer3_outputs(4213) <= not((layer2_outputs(3834)) or (layer2_outputs(145)));
    layer3_outputs(4214) <= '1';
    layer3_outputs(4215) <= not(layer2_outputs(2491));
    layer3_outputs(4216) <= (layer2_outputs(2605)) and not (layer2_outputs(5078));
    layer3_outputs(4217) <= not(layer2_outputs(3033));
    layer3_outputs(4218) <= (layer2_outputs(376)) and not (layer2_outputs(340));
    layer3_outputs(4219) <= '0';
    layer3_outputs(4220) <= not(layer2_outputs(2720)) or (layer2_outputs(6645));
    layer3_outputs(4221) <= layer2_outputs(3357);
    layer3_outputs(4222) <= (layer2_outputs(6612)) and (layer2_outputs(360));
    layer3_outputs(4223) <= not((layer2_outputs(2607)) or (layer2_outputs(298)));
    layer3_outputs(4224) <= (layer2_outputs(2160)) and not (layer2_outputs(4785));
    layer3_outputs(4225) <= '1';
    layer3_outputs(4226) <= layer2_outputs(4467);
    layer3_outputs(4227) <= (layer2_outputs(7477)) or (layer2_outputs(5702));
    layer3_outputs(4228) <= (layer2_outputs(0)) and (layer2_outputs(5776));
    layer3_outputs(4229) <= layer2_outputs(7067);
    layer3_outputs(4230) <= (layer2_outputs(1705)) and not (layer2_outputs(6226));
    layer3_outputs(4231) <= not(layer2_outputs(2066));
    layer3_outputs(4232) <= (layer2_outputs(6150)) or (layer2_outputs(5694));
    layer3_outputs(4233) <= (layer2_outputs(1699)) and (layer2_outputs(2308));
    layer3_outputs(4234) <= (layer2_outputs(5732)) xor (layer2_outputs(1910));
    layer3_outputs(4235) <= not(layer2_outputs(1940)) or (layer2_outputs(1966));
    layer3_outputs(4236) <= not((layer2_outputs(2416)) and (layer2_outputs(3119)));
    layer3_outputs(4237) <= layer2_outputs(150);
    layer3_outputs(4238) <= layer2_outputs(717);
    layer3_outputs(4239) <= layer2_outputs(1846);
    layer3_outputs(4240) <= layer2_outputs(5397);
    layer3_outputs(4241) <= (layer2_outputs(1397)) xor (layer2_outputs(93));
    layer3_outputs(4242) <= '1';
    layer3_outputs(4243) <= '1';
    layer3_outputs(4244) <= layer2_outputs(7244);
    layer3_outputs(4245) <= layer2_outputs(5616);
    layer3_outputs(4246) <= (layer2_outputs(5334)) and (layer2_outputs(4665));
    layer3_outputs(4247) <= not(layer2_outputs(6774));
    layer3_outputs(4248) <= layer2_outputs(4424);
    layer3_outputs(4249) <= not(layer2_outputs(6093)) or (layer2_outputs(3600));
    layer3_outputs(4250) <= (layer2_outputs(4211)) or (layer2_outputs(1070));
    layer3_outputs(4251) <= layer2_outputs(4907);
    layer3_outputs(4252) <= '0';
    layer3_outputs(4253) <= layer2_outputs(4396);
    layer3_outputs(4254) <= (layer2_outputs(6609)) and (layer2_outputs(4234));
    layer3_outputs(4255) <= (layer2_outputs(4960)) and (layer2_outputs(5492));
    layer3_outputs(4256) <= (layer2_outputs(3853)) and not (layer2_outputs(5301));
    layer3_outputs(4257) <= not(layer2_outputs(2));
    layer3_outputs(4258) <= '1';
    layer3_outputs(4259) <= layer2_outputs(4588);
    layer3_outputs(4260) <= layer2_outputs(1096);
    layer3_outputs(4261) <= layer2_outputs(4860);
    layer3_outputs(4262) <= not((layer2_outputs(7398)) or (layer2_outputs(7578)));
    layer3_outputs(4263) <= not((layer2_outputs(1941)) or (layer2_outputs(6439)));
    layer3_outputs(4264) <= layer2_outputs(7220);
    layer3_outputs(4265) <= (layer2_outputs(4475)) and not (layer2_outputs(3865));
    layer3_outputs(4266) <= not(layer2_outputs(5675));
    layer3_outputs(4267) <= (layer2_outputs(5554)) and (layer2_outputs(4811));
    layer3_outputs(4268) <= '1';
    layer3_outputs(4269) <= (layer2_outputs(5405)) and not (layer2_outputs(2026));
    layer3_outputs(4270) <= (layer2_outputs(5006)) and (layer2_outputs(6755));
    layer3_outputs(4271) <= '1';
    layer3_outputs(4272) <= not(layer2_outputs(5041));
    layer3_outputs(4273) <= not(layer2_outputs(4624));
    layer3_outputs(4274) <= not(layer2_outputs(5591));
    layer3_outputs(4275) <= '0';
    layer3_outputs(4276) <= layer2_outputs(4911);
    layer3_outputs(4277) <= layer2_outputs(5159);
    layer3_outputs(4278) <= (layer2_outputs(6894)) and (layer2_outputs(2934));
    layer3_outputs(4279) <= layer2_outputs(6827);
    layer3_outputs(4280) <= (layer2_outputs(7609)) and not (layer2_outputs(3443));
    layer3_outputs(4281) <= (layer2_outputs(1396)) or (layer2_outputs(7670));
    layer3_outputs(4282) <= '1';
    layer3_outputs(4283) <= not((layer2_outputs(2875)) xor (layer2_outputs(1989)));
    layer3_outputs(4284) <= not(layer2_outputs(3730));
    layer3_outputs(4285) <= not(layer2_outputs(4589)) or (layer2_outputs(2418));
    layer3_outputs(4286) <= not(layer2_outputs(7587)) or (layer2_outputs(7125));
    layer3_outputs(4287) <= not(layer2_outputs(7538)) or (layer2_outputs(1619));
    layer3_outputs(4288) <= layer2_outputs(5429);
    layer3_outputs(4289) <= (layer2_outputs(7132)) and not (layer2_outputs(4958));
    layer3_outputs(4290) <= layer2_outputs(5318);
    layer3_outputs(4291) <= not(layer2_outputs(5268));
    layer3_outputs(4292) <= (layer2_outputs(4927)) and (layer2_outputs(2508));
    layer3_outputs(4293) <= not(layer2_outputs(2939));
    layer3_outputs(4294) <= not(layer2_outputs(899));
    layer3_outputs(4295) <= not(layer2_outputs(3388)) or (layer2_outputs(5601));
    layer3_outputs(4296) <= (layer2_outputs(6505)) and not (layer2_outputs(6096));
    layer3_outputs(4297) <= layer2_outputs(2147);
    layer3_outputs(4298) <= layer2_outputs(5643);
    layer3_outputs(4299) <= not(layer2_outputs(2541));
    layer3_outputs(4300) <= layer2_outputs(4567);
    layer3_outputs(4301) <= (layer2_outputs(5110)) or (layer2_outputs(1128));
    layer3_outputs(4302) <= (layer2_outputs(781)) and not (layer2_outputs(1157));
    layer3_outputs(4303) <= (layer2_outputs(531)) and not (layer2_outputs(2574));
    layer3_outputs(4304) <= '0';
    layer3_outputs(4305) <= '0';
    layer3_outputs(4306) <= (layer2_outputs(2890)) and not (layer2_outputs(1779));
    layer3_outputs(4307) <= layer2_outputs(6916);
    layer3_outputs(4308) <= not((layer2_outputs(6169)) xor (layer2_outputs(7492)));
    layer3_outputs(4309) <= not(layer2_outputs(5794)) or (layer2_outputs(4735));
    layer3_outputs(4310) <= (layer2_outputs(2795)) or (layer2_outputs(5446));
    layer3_outputs(4311) <= not(layer2_outputs(685));
    layer3_outputs(4312) <= not(layer2_outputs(1009)) or (layer2_outputs(1309));
    layer3_outputs(4313) <= not(layer2_outputs(7514));
    layer3_outputs(4314) <= not((layer2_outputs(6790)) and (layer2_outputs(4272)));
    layer3_outputs(4315) <= (layer2_outputs(1990)) or (layer2_outputs(7658));
    layer3_outputs(4316) <= not(layer2_outputs(1156));
    layer3_outputs(4317) <= '0';
    layer3_outputs(4318) <= not((layer2_outputs(2599)) xor (layer2_outputs(1437)));
    layer3_outputs(4319) <= (layer2_outputs(2303)) and not (layer2_outputs(6817));
    layer3_outputs(4320) <= not(layer2_outputs(3349));
    layer3_outputs(4321) <= not((layer2_outputs(3092)) and (layer2_outputs(902)));
    layer3_outputs(4322) <= (layer2_outputs(4342)) and not (layer2_outputs(7427));
    layer3_outputs(4323) <= not(layer2_outputs(6760));
    layer3_outputs(4324) <= not(layer2_outputs(6669)) or (layer2_outputs(7461));
    layer3_outputs(4325) <= not(layer2_outputs(2894)) or (layer2_outputs(1766));
    layer3_outputs(4326) <= not((layer2_outputs(4516)) xor (layer2_outputs(2023)));
    layer3_outputs(4327) <= not((layer2_outputs(431)) and (layer2_outputs(4289)));
    layer3_outputs(4328) <= not(layer2_outputs(7633));
    layer3_outputs(4329) <= '1';
    layer3_outputs(4330) <= (layer2_outputs(6473)) and not (layer2_outputs(6009));
    layer3_outputs(4331) <= layer2_outputs(240);
    layer3_outputs(4332) <= layer2_outputs(6237);
    layer3_outputs(4333) <= (layer2_outputs(1357)) and not (layer2_outputs(416));
    layer3_outputs(4334) <= not(layer2_outputs(5201));
    layer3_outputs(4335) <= layer2_outputs(5756);
    layer3_outputs(4336) <= not(layer2_outputs(2641));
    layer3_outputs(4337) <= layer2_outputs(6067);
    layer3_outputs(4338) <= (layer2_outputs(4001)) and not (layer2_outputs(3617));
    layer3_outputs(4339) <= not(layer2_outputs(2992)) or (layer2_outputs(1384));
    layer3_outputs(4340) <= (layer2_outputs(4122)) and not (layer2_outputs(1816));
    layer3_outputs(4341) <= not(layer2_outputs(4900));
    layer3_outputs(4342) <= layer2_outputs(4437);
    layer3_outputs(4343) <= not((layer2_outputs(3530)) or (layer2_outputs(5413)));
    layer3_outputs(4344) <= not((layer2_outputs(4758)) and (layer2_outputs(5347)));
    layer3_outputs(4345) <= not(layer2_outputs(7488));
    layer3_outputs(4346) <= not((layer2_outputs(6910)) and (layer2_outputs(3047)));
    layer3_outputs(4347) <= not(layer2_outputs(2952));
    layer3_outputs(4348) <= (layer2_outputs(5262)) and not (layer2_outputs(2009));
    layer3_outputs(4349) <= not(layer2_outputs(38));
    layer3_outputs(4350) <= not(layer2_outputs(3669));
    layer3_outputs(4351) <= layer2_outputs(675);
    layer3_outputs(4352) <= (layer2_outputs(7383)) and (layer2_outputs(651));
    layer3_outputs(4353) <= '1';
    layer3_outputs(4354) <= layer2_outputs(1092);
    layer3_outputs(4355) <= layer2_outputs(2710);
    layer3_outputs(4356) <= (layer2_outputs(6676)) and not (layer2_outputs(4335));
    layer3_outputs(4357) <= (layer2_outputs(5952)) or (layer2_outputs(2872));
    layer3_outputs(4358) <= (layer2_outputs(4834)) and not (layer2_outputs(7545));
    layer3_outputs(4359) <= not(layer2_outputs(5230));
    layer3_outputs(4360) <= layer2_outputs(7162);
    layer3_outputs(4361) <= layer2_outputs(4897);
    layer3_outputs(4362) <= (layer2_outputs(7535)) and not (layer2_outputs(2540));
    layer3_outputs(4363) <= not(layer2_outputs(281)) or (layer2_outputs(1011));
    layer3_outputs(4364) <= (layer2_outputs(704)) or (layer2_outputs(2354));
    layer3_outputs(4365) <= layer2_outputs(1558);
    layer3_outputs(4366) <= '1';
    layer3_outputs(4367) <= layer2_outputs(2941);
    layer3_outputs(4368) <= '0';
    layer3_outputs(4369) <= not(layer2_outputs(4252));
    layer3_outputs(4370) <= layer2_outputs(5591);
    layer3_outputs(4371) <= layer2_outputs(2576);
    layer3_outputs(4372) <= (layer2_outputs(4615)) and not (layer2_outputs(1810));
    layer3_outputs(4373) <= (layer2_outputs(2793)) and not (layer2_outputs(2060));
    layer3_outputs(4374) <= '1';
    layer3_outputs(4375) <= not((layer2_outputs(962)) or (layer2_outputs(279)));
    layer3_outputs(4376) <= (layer2_outputs(6542)) or (layer2_outputs(2750));
    layer3_outputs(4377) <= layer2_outputs(6791);
    layer3_outputs(4378) <= not(layer2_outputs(1408));
    layer3_outputs(4379) <= not((layer2_outputs(1055)) and (layer2_outputs(3293)));
    layer3_outputs(4380) <= not(layer2_outputs(4648)) or (layer2_outputs(3434));
    layer3_outputs(4381) <= layer2_outputs(6560);
    layer3_outputs(4382) <= not((layer2_outputs(4079)) and (layer2_outputs(1367)));
    layer3_outputs(4383) <= not(layer2_outputs(1964));
    layer3_outputs(4384) <= not(layer2_outputs(2266)) or (layer2_outputs(4369));
    layer3_outputs(4385) <= not(layer2_outputs(5579));
    layer3_outputs(4386) <= not(layer2_outputs(6393)) or (layer2_outputs(1780));
    layer3_outputs(4387) <= (layer2_outputs(5515)) and not (layer2_outputs(3310));
    layer3_outputs(4388) <= not((layer2_outputs(5363)) xor (layer2_outputs(2955)));
    layer3_outputs(4389) <= layer2_outputs(633);
    layer3_outputs(4390) <= (layer2_outputs(1355)) and not (layer2_outputs(4222));
    layer3_outputs(4391) <= not(layer2_outputs(92));
    layer3_outputs(4392) <= '0';
    layer3_outputs(4393) <= layer2_outputs(5154);
    layer3_outputs(4394) <= not((layer2_outputs(4351)) and (layer2_outputs(7298)));
    layer3_outputs(4395) <= layer2_outputs(1569);
    layer3_outputs(4396) <= not(layer2_outputs(5027)) or (layer2_outputs(5560));
    layer3_outputs(4397) <= (layer2_outputs(7112)) xor (layer2_outputs(6772));
    layer3_outputs(4398) <= (layer2_outputs(5539)) and not (layer2_outputs(7137));
    layer3_outputs(4399) <= layer2_outputs(1088);
    layer3_outputs(4400) <= not(layer2_outputs(5555));
    layer3_outputs(4401) <= '0';
    layer3_outputs(4402) <= not(layer2_outputs(2353));
    layer3_outputs(4403) <= not(layer2_outputs(6173));
    layer3_outputs(4404) <= (layer2_outputs(5085)) and (layer2_outputs(6100));
    layer3_outputs(4405) <= not(layer2_outputs(6948));
    layer3_outputs(4406) <= not(layer2_outputs(2996));
    layer3_outputs(4407) <= not(layer2_outputs(2561)) or (layer2_outputs(2017));
    layer3_outputs(4408) <= not(layer2_outputs(5815));
    layer3_outputs(4409) <= not(layer2_outputs(2364));
    layer3_outputs(4410) <= not(layer2_outputs(6841));
    layer3_outputs(4411) <= (layer2_outputs(2035)) or (layer2_outputs(860));
    layer3_outputs(4412) <= not(layer2_outputs(4657));
    layer3_outputs(4413) <= layer2_outputs(4998);
    layer3_outputs(4414) <= not(layer2_outputs(1093)) or (layer2_outputs(4672));
    layer3_outputs(4415) <= (layer2_outputs(4115)) and (layer2_outputs(1530));
    layer3_outputs(4416) <= layer2_outputs(915);
    layer3_outputs(4417) <= (layer2_outputs(5189)) and not (layer2_outputs(7449));
    layer3_outputs(4418) <= not((layer2_outputs(561)) or (layer2_outputs(4859)));
    layer3_outputs(4419) <= layer2_outputs(3759);
    layer3_outputs(4420) <= not((layer2_outputs(4369)) and (layer2_outputs(1192)));
    layer3_outputs(4421) <= not(layer2_outputs(3463));
    layer3_outputs(4422) <= not(layer2_outputs(7583)) or (layer2_outputs(5352));
    layer3_outputs(4423) <= not(layer2_outputs(7320));
    layer3_outputs(4424) <= '1';
    layer3_outputs(4425) <= not((layer2_outputs(2095)) or (layer2_outputs(1584)));
    layer3_outputs(4426) <= layer2_outputs(2929);
    layer3_outputs(4427) <= layer2_outputs(4149);
    layer3_outputs(4428) <= not(layer2_outputs(5596));
    layer3_outputs(4429) <= not((layer2_outputs(6329)) and (layer2_outputs(4264)));
    layer3_outputs(4430) <= (layer2_outputs(6126)) or (layer2_outputs(7603));
    layer3_outputs(4431) <= not(layer2_outputs(1301)) or (layer2_outputs(959));
    layer3_outputs(4432) <= not(layer2_outputs(6467));
    layer3_outputs(4433) <= not(layer2_outputs(6677)) or (layer2_outputs(46));
    layer3_outputs(4434) <= layer2_outputs(4806);
    layer3_outputs(4435) <= (layer2_outputs(1304)) and not (layer2_outputs(7520));
    layer3_outputs(4436) <= not(layer2_outputs(5527)) or (layer2_outputs(4620));
    layer3_outputs(4437) <= not((layer2_outputs(7262)) or (layer2_outputs(743)));
    layer3_outputs(4438) <= layer2_outputs(4159);
    layer3_outputs(4439) <= layer2_outputs(2755);
    layer3_outputs(4440) <= (layer2_outputs(2494)) and (layer2_outputs(3504));
    layer3_outputs(4441) <= not(layer2_outputs(7140));
    layer3_outputs(4442) <= (layer2_outputs(2140)) or (layer2_outputs(4774));
    layer3_outputs(4443) <= layer2_outputs(1286);
    layer3_outputs(4444) <= layer2_outputs(1318);
    layer3_outputs(4445) <= '0';
    layer3_outputs(4446) <= layer2_outputs(2121);
    layer3_outputs(4447) <= not(layer2_outputs(7391));
    layer3_outputs(4448) <= (layer2_outputs(7515)) and not (layer2_outputs(7073));
    layer3_outputs(4449) <= not((layer2_outputs(6124)) xor (layer2_outputs(6616)));
    layer3_outputs(4450) <= not(layer2_outputs(7637));
    layer3_outputs(4451) <= not(layer2_outputs(1735)) or (layer2_outputs(271));
    layer3_outputs(4452) <= not(layer2_outputs(7457));
    layer3_outputs(4453) <= not(layer2_outputs(1822)) or (layer2_outputs(4621));
    layer3_outputs(4454) <= not(layer2_outputs(1414));
    layer3_outputs(4455) <= layer2_outputs(2279);
    layer3_outputs(4456) <= (layer2_outputs(777)) and (layer2_outputs(6024));
    layer3_outputs(4457) <= not(layer2_outputs(249));
    layer3_outputs(4458) <= not(layer2_outputs(4064));
    layer3_outputs(4459) <= layer2_outputs(5661);
    layer3_outputs(4460) <= not(layer2_outputs(7202));
    layer3_outputs(4461) <= (layer2_outputs(7036)) or (layer2_outputs(3835));
    layer3_outputs(4462) <= '0';
    layer3_outputs(4463) <= not((layer2_outputs(1441)) xor (layer2_outputs(6810)));
    layer3_outputs(4464) <= not(layer2_outputs(2014));
    layer3_outputs(4465) <= layer2_outputs(2827);
    layer3_outputs(4466) <= '0';
    layer3_outputs(4467) <= not((layer2_outputs(3304)) and (layer2_outputs(1031)));
    layer3_outputs(4468) <= (layer2_outputs(7090)) and not (layer2_outputs(5118));
    layer3_outputs(4469) <= not(layer2_outputs(2729));
    layer3_outputs(4470) <= not((layer2_outputs(7326)) and (layer2_outputs(2493)));
    layer3_outputs(4471) <= not(layer2_outputs(151));
    layer3_outputs(4472) <= '1';
    layer3_outputs(4473) <= '1';
    layer3_outputs(4474) <= '0';
    layer3_outputs(4475) <= not(layer2_outputs(302));
    layer3_outputs(4476) <= layer2_outputs(3402);
    layer3_outputs(4477) <= (layer2_outputs(1047)) and not (layer2_outputs(1664));
    layer3_outputs(4478) <= (layer2_outputs(548)) or (layer2_outputs(6102));
    layer3_outputs(4479) <= not((layer2_outputs(1815)) or (layer2_outputs(68)));
    layer3_outputs(4480) <= layer2_outputs(4413);
    layer3_outputs(4481) <= (layer2_outputs(7257)) and (layer2_outputs(3784));
    layer3_outputs(4482) <= not(layer2_outputs(2310));
    layer3_outputs(4483) <= not(layer2_outputs(512));
    layer3_outputs(4484) <= '0';
    layer3_outputs(4485) <= layer2_outputs(5222);
    layer3_outputs(4486) <= (layer2_outputs(1820)) and not (layer2_outputs(7207));
    layer3_outputs(4487) <= (layer2_outputs(7025)) and (layer2_outputs(1669));
    layer3_outputs(4488) <= not(layer2_outputs(284));
    layer3_outputs(4489) <= (layer2_outputs(2442)) and (layer2_outputs(4072));
    layer3_outputs(4490) <= (layer2_outputs(5713)) or (layer2_outputs(676));
    layer3_outputs(4491) <= layer2_outputs(3422);
    layer3_outputs(4492) <= (layer2_outputs(5677)) and (layer2_outputs(3410));
    layer3_outputs(4493) <= not(layer2_outputs(4779)) or (layer2_outputs(1563));
    layer3_outputs(4494) <= '0';
    layer3_outputs(4495) <= (layer2_outputs(6593)) or (layer2_outputs(5566));
    layer3_outputs(4496) <= (layer2_outputs(5479)) or (layer2_outputs(1297));
    layer3_outputs(4497) <= layer2_outputs(6553);
    layer3_outputs(4498) <= (layer2_outputs(4414)) and not (layer2_outputs(995));
    layer3_outputs(4499) <= '1';
    layer3_outputs(4500) <= '0';
    layer3_outputs(4501) <= (layer2_outputs(4417)) and (layer2_outputs(5919));
    layer3_outputs(4502) <= layer2_outputs(6247);
    layer3_outputs(4503) <= (layer2_outputs(3055)) or (layer2_outputs(46));
    layer3_outputs(4504) <= (layer2_outputs(2724)) and not (layer2_outputs(7014));
    layer3_outputs(4505) <= not(layer2_outputs(6579));
    layer3_outputs(4506) <= not(layer2_outputs(7597)) or (layer2_outputs(4042));
    layer3_outputs(4507) <= not((layer2_outputs(6026)) or (layer2_outputs(635)));
    layer3_outputs(4508) <= not(layer2_outputs(470));
    layer3_outputs(4509) <= (layer2_outputs(2119)) and (layer2_outputs(3754));
    layer3_outputs(4510) <= layer2_outputs(6656);
    layer3_outputs(4511) <= not(layer2_outputs(2548)) or (layer2_outputs(729));
    layer3_outputs(4512) <= not((layer2_outputs(2509)) and (layer2_outputs(1663)));
    layer3_outputs(4513) <= not(layer2_outputs(3270));
    layer3_outputs(4514) <= '0';
    layer3_outputs(4515) <= not(layer2_outputs(238)) or (layer2_outputs(7011));
    layer3_outputs(4516) <= not(layer2_outputs(2511)) or (layer2_outputs(1418));
    layer3_outputs(4517) <= (layer2_outputs(6740)) or (layer2_outputs(6729));
    layer3_outputs(4518) <= (layer2_outputs(6764)) or (layer2_outputs(6745));
    layer3_outputs(4519) <= layer2_outputs(1919);
    layer3_outputs(4520) <= not(layer2_outputs(6227));
    layer3_outputs(4521) <= (layer2_outputs(2477)) or (layer2_outputs(2108));
    layer3_outputs(4522) <= not(layer2_outputs(5018)) or (layer2_outputs(538));
    layer3_outputs(4523) <= (layer2_outputs(2309)) and not (layer2_outputs(3007));
    layer3_outputs(4524) <= layer2_outputs(6483);
    layer3_outputs(4525) <= (layer2_outputs(7300)) and (layer2_outputs(5995));
    layer3_outputs(4526) <= layer2_outputs(5215);
    layer3_outputs(4527) <= layer2_outputs(2396);
    layer3_outputs(4528) <= layer2_outputs(4207);
    layer3_outputs(4529) <= (layer2_outputs(2586)) and not (layer2_outputs(5629));
    layer3_outputs(4530) <= not(layer2_outputs(6715));
    layer3_outputs(4531) <= layer2_outputs(7270);
    layer3_outputs(4532) <= layer2_outputs(1998);
    layer3_outputs(4533) <= not(layer2_outputs(6828)) or (layer2_outputs(5172));
    layer3_outputs(4534) <= layer2_outputs(5196);
    layer3_outputs(4535) <= not(layer2_outputs(4442));
    layer3_outputs(4536) <= layer2_outputs(1930);
    layer3_outputs(4537) <= (layer2_outputs(7174)) and (layer2_outputs(5234));
    layer3_outputs(4538) <= not(layer2_outputs(2437));
    layer3_outputs(4539) <= layer2_outputs(3974);
    layer3_outputs(4540) <= (layer2_outputs(7230)) and (layer2_outputs(7532));
    layer3_outputs(4541) <= not(layer2_outputs(757)) or (layer2_outputs(3376));
    layer3_outputs(4542) <= not((layer2_outputs(4675)) and (layer2_outputs(2943)));
    layer3_outputs(4543) <= '1';
    layer3_outputs(4544) <= (layer2_outputs(2020)) and (layer2_outputs(1465));
    layer3_outputs(4545) <= layer2_outputs(28);
    layer3_outputs(4546) <= not((layer2_outputs(3472)) or (layer2_outputs(4267)));
    layer3_outputs(4547) <= layer2_outputs(5261);
    layer3_outputs(4548) <= not(layer2_outputs(1854)) or (layer2_outputs(7497));
    layer3_outputs(4549) <= (layer2_outputs(6149)) and (layer2_outputs(463));
    layer3_outputs(4550) <= (layer2_outputs(4359)) and not (layer2_outputs(6368));
    layer3_outputs(4551) <= not(layer2_outputs(6156));
    layer3_outputs(4552) <= not(layer2_outputs(6819)) or (layer2_outputs(4080));
    layer3_outputs(4553) <= not(layer2_outputs(6465));
    layer3_outputs(4554) <= (layer2_outputs(2567)) and not (layer2_outputs(1989));
    layer3_outputs(4555) <= not((layer2_outputs(2410)) or (layer2_outputs(7525)));
    layer3_outputs(4556) <= (layer2_outputs(1992)) and (layer2_outputs(1281));
    layer3_outputs(4557) <= '1';
    layer3_outputs(4558) <= layer2_outputs(5204);
    layer3_outputs(4559) <= layer2_outputs(6900);
    layer3_outputs(4560) <= (layer2_outputs(6079)) and not (layer2_outputs(4061));
    layer3_outputs(4561) <= layer2_outputs(366);
    layer3_outputs(4562) <= layer2_outputs(500);
    layer3_outputs(4563) <= '0';
    layer3_outputs(4564) <= '0';
    layer3_outputs(4565) <= layer2_outputs(5986);
    layer3_outputs(4566) <= not((layer2_outputs(3214)) or (layer2_outputs(2864)));
    layer3_outputs(4567) <= not((layer2_outputs(3178)) or (layer2_outputs(5087)));
    layer3_outputs(4568) <= (layer2_outputs(818)) and (layer2_outputs(1950));
    layer3_outputs(4569) <= not(layer2_outputs(2606));
    layer3_outputs(4570) <= (layer2_outputs(3794)) xor (layer2_outputs(1486));
    layer3_outputs(4571) <= layer2_outputs(2334);
    layer3_outputs(4572) <= not(layer2_outputs(3109)) or (layer2_outputs(3299));
    layer3_outputs(4573) <= not(layer2_outputs(2949));
    layer3_outputs(4574) <= not((layer2_outputs(1194)) or (layer2_outputs(4519)));
    layer3_outputs(4575) <= not(layer2_outputs(5357));
    layer3_outputs(4576) <= layer2_outputs(6159);
    layer3_outputs(4577) <= (layer2_outputs(3657)) and not (layer2_outputs(2254));
    layer3_outputs(4578) <= '0';
    layer3_outputs(4579) <= not(layer2_outputs(95));
    layer3_outputs(4580) <= not(layer2_outputs(3164));
    layer3_outputs(4581) <= '0';
    layer3_outputs(4582) <= (layer2_outputs(3917)) and not (layer2_outputs(2839));
    layer3_outputs(4583) <= (layer2_outputs(5463)) and not (layer2_outputs(2273));
    layer3_outputs(4584) <= (layer2_outputs(6862)) or (layer2_outputs(5706));
    layer3_outputs(4585) <= layer2_outputs(5804);
    layer3_outputs(4586) <= layer2_outputs(7537);
    layer3_outputs(4587) <= not((layer2_outputs(6102)) and (layer2_outputs(7049)));
    layer3_outputs(4588) <= layer2_outputs(3906);
    layer3_outputs(4589) <= not((layer2_outputs(1902)) and (layer2_outputs(2363)));
    layer3_outputs(4590) <= '1';
    layer3_outputs(4591) <= (layer2_outputs(4368)) and not (layer2_outputs(5759));
    layer3_outputs(4592) <= not(layer2_outputs(4835)) or (layer2_outputs(6378));
    layer3_outputs(4593) <= not(layer2_outputs(2478));
    layer3_outputs(4594) <= not(layer2_outputs(1065)) or (layer2_outputs(2828));
    layer3_outputs(4595) <= layer2_outputs(6683);
    layer3_outputs(4596) <= not(layer2_outputs(3808)) or (layer2_outputs(5980));
    layer3_outputs(4597) <= not(layer2_outputs(40)) or (layer2_outputs(4756));
    layer3_outputs(4598) <= layer2_outputs(724);
    layer3_outputs(4599) <= not(layer2_outputs(5371)) or (layer2_outputs(2190));
    layer3_outputs(4600) <= layer2_outputs(532);
    layer3_outputs(4601) <= (layer2_outputs(3264)) xor (layer2_outputs(6502));
    layer3_outputs(4602) <= (layer2_outputs(3267)) or (layer2_outputs(5967));
    layer3_outputs(4603) <= not(layer2_outputs(4355)) or (layer2_outputs(6766));
    layer3_outputs(4604) <= layer2_outputs(6625);
    layer3_outputs(4605) <= layer2_outputs(572);
    layer3_outputs(4606) <= layer2_outputs(5628);
    layer3_outputs(4607) <= not(layer2_outputs(5862));
    layer3_outputs(4608) <= layer2_outputs(1818);
    layer3_outputs(4609) <= (layer2_outputs(3924)) and not (layer2_outputs(6958));
    layer3_outputs(4610) <= layer2_outputs(3247);
    layer3_outputs(4611) <= '1';
    layer3_outputs(4612) <= '1';
    layer3_outputs(4613) <= (layer2_outputs(1850)) and not (layer2_outputs(226));
    layer3_outputs(4614) <= layer2_outputs(1862);
    layer3_outputs(4615) <= not(layer2_outputs(4376)) or (layer2_outputs(1675));
    layer3_outputs(4616) <= layer2_outputs(5982);
    layer3_outputs(4617) <= layer2_outputs(2419);
    layer3_outputs(4618) <= layer2_outputs(4953);
    layer3_outputs(4619) <= not((layer2_outputs(4442)) or (layer2_outputs(636)));
    layer3_outputs(4620) <= layer2_outputs(2924);
    layer3_outputs(4621) <= '1';
    layer3_outputs(4622) <= (layer2_outputs(3759)) and not (layer2_outputs(911));
    layer3_outputs(4623) <= (layer2_outputs(1026)) and (layer2_outputs(2968));
    layer3_outputs(4624) <= '0';
    layer3_outputs(4625) <= (layer2_outputs(737)) and not (layer2_outputs(5054));
    layer3_outputs(4626) <= '1';
    layer3_outputs(4627) <= layer2_outputs(6807);
    layer3_outputs(4628) <= '1';
    layer3_outputs(4629) <= not(layer2_outputs(2759)) or (layer2_outputs(2856));
    layer3_outputs(4630) <= '1';
    layer3_outputs(4631) <= not(layer2_outputs(5163));
    layer3_outputs(4632) <= (layer2_outputs(5129)) and not (layer2_outputs(7669));
    layer3_outputs(4633) <= not((layer2_outputs(7565)) and (layer2_outputs(923)));
    layer3_outputs(4634) <= not((layer2_outputs(4136)) or (layer2_outputs(1284)));
    layer3_outputs(4635) <= (layer2_outputs(1449)) or (layer2_outputs(3346));
    layer3_outputs(4636) <= not((layer2_outputs(6867)) or (layer2_outputs(111)));
    layer3_outputs(4637) <= not(layer2_outputs(4020));
    layer3_outputs(4638) <= not((layer2_outputs(3624)) or (layer2_outputs(495)));
    layer3_outputs(4639) <= layer2_outputs(2078);
    layer3_outputs(4640) <= (layer2_outputs(1640)) or (layer2_outputs(7580));
    layer3_outputs(4641) <= not(layer2_outputs(18));
    layer3_outputs(4642) <= not(layer2_outputs(3743));
    layer3_outputs(4643) <= (layer2_outputs(3115)) and not (layer2_outputs(458));
    layer3_outputs(4644) <= layer2_outputs(513);
    layer3_outputs(4645) <= not(layer2_outputs(6377));
    layer3_outputs(4646) <= not(layer2_outputs(6408));
    layer3_outputs(4647) <= (layer2_outputs(7246)) and not (layer2_outputs(6960));
    layer3_outputs(4648) <= layer2_outputs(5250);
    layer3_outputs(4649) <= (layer2_outputs(6130)) and (layer2_outputs(212));
    layer3_outputs(4650) <= (layer2_outputs(7021)) and not (layer2_outputs(4584));
    layer3_outputs(4651) <= not(layer2_outputs(2494));
    layer3_outputs(4652) <= not(layer2_outputs(3520));
    layer3_outputs(4653) <= not(layer2_outputs(4677));
    layer3_outputs(4654) <= not((layer2_outputs(3864)) or (layer2_outputs(343)));
    layer3_outputs(4655) <= layer2_outputs(6434);
    layer3_outputs(4656) <= '0';
    layer3_outputs(4657) <= '1';
    layer3_outputs(4658) <= not(layer2_outputs(4912));
    layer3_outputs(4659) <= not((layer2_outputs(3291)) and (layer2_outputs(6682)));
    layer3_outputs(4660) <= not((layer2_outputs(6383)) or (layer2_outputs(4265)));
    layer3_outputs(4661) <= '1';
    layer3_outputs(4662) <= '1';
    layer3_outputs(4663) <= not(layer2_outputs(3090));
    layer3_outputs(4664) <= (layer2_outputs(7563)) or (layer2_outputs(5453));
    layer3_outputs(4665) <= not(layer2_outputs(7378)) or (layer2_outputs(5190));
    layer3_outputs(4666) <= not(layer2_outputs(2744));
    layer3_outputs(4667) <= (layer2_outputs(1921)) and not (layer2_outputs(6248));
    layer3_outputs(4668) <= not(layer2_outputs(2337));
    layer3_outputs(4669) <= (layer2_outputs(1769)) xor (layer2_outputs(4953));
    layer3_outputs(4670) <= (layer2_outputs(4762)) or (layer2_outputs(978));
    layer3_outputs(4671) <= (layer2_outputs(7402)) xor (layer2_outputs(1688));
    layer3_outputs(4672) <= layer2_outputs(3071);
    layer3_outputs(4673) <= not(layer2_outputs(863));
    layer3_outputs(4674) <= '0';
    layer3_outputs(4675) <= layer2_outputs(4401);
    layer3_outputs(4676) <= not(layer2_outputs(5713));
    layer3_outputs(4677) <= not(layer2_outputs(2241)) or (layer2_outputs(1710));
    layer3_outputs(4678) <= not(layer2_outputs(709));
    layer3_outputs(4679) <= not(layer2_outputs(4071)) or (layer2_outputs(227));
    layer3_outputs(4680) <= not(layer2_outputs(611));
    layer3_outputs(4681) <= not((layer2_outputs(6284)) or (layer2_outputs(4116)));
    layer3_outputs(4682) <= layer2_outputs(4952);
    layer3_outputs(4683) <= (layer2_outputs(6565)) xor (layer2_outputs(6574));
    layer3_outputs(4684) <= layer2_outputs(6495);
    layer3_outputs(4685) <= not(layer2_outputs(7387));
    layer3_outputs(4686) <= layer2_outputs(2016);
    layer3_outputs(4687) <= (layer2_outputs(3708)) or (layer2_outputs(3984));
    layer3_outputs(4688) <= (layer2_outputs(2914)) and not (layer2_outputs(7553));
    layer3_outputs(4689) <= '1';
    layer3_outputs(4690) <= not(layer2_outputs(1792));
    layer3_outputs(4691) <= not(layer2_outputs(7575));
    layer3_outputs(4692) <= not((layer2_outputs(541)) xor (layer2_outputs(6107)));
    layer3_outputs(4693) <= (layer2_outputs(4184)) and not (layer2_outputs(7153));
    layer3_outputs(4694) <= (layer2_outputs(79)) and (layer2_outputs(625));
    layer3_outputs(4695) <= not(layer2_outputs(6035));
    layer3_outputs(4696) <= (layer2_outputs(5888)) or (layer2_outputs(7165));
    layer3_outputs(4697) <= not(layer2_outputs(895));
    layer3_outputs(4698) <= '1';
    layer3_outputs(4699) <= (layer2_outputs(5801)) and (layer2_outputs(268));
    layer3_outputs(4700) <= (layer2_outputs(5343)) and not (layer2_outputs(6));
    layer3_outputs(4701) <= layer2_outputs(7155);
    layer3_outputs(4702) <= (layer2_outputs(804)) and not (layer2_outputs(5515));
    layer3_outputs(4703) <= not(layer2_outputs(4284));
    layer3_outputs(4704) <= not(layer2_outputs(7581));
    layer3_outputs(4705) <= layer2_outputs(3487);
    layer3_outputs(4706) <= (layer2_outputs(6734)) and (layer2_outputs(377));
    layer3_outputs(4707) <= (layer2_outputs(667)) and not (layer2_outputs(828));
    layer3_outputs(4708) <= not((layer2_outputs(3618)) or (layer2_outputs(1348)));
    layer3_outputs(4709) <= '1';
    layer3_outputs(4710) <= layer2_outputs(4862);
    layer3_outputs(4711) <= layer2_outputs(3937);
    layer3_outputs(4712) <= layer2_outputs(1810);
    layer3_outputs(4713) <= layer2_outputs(4103);
    layer3_outputs(4714) <= layer2_outputs(4972);
    layer3_outputs(4715) <= '1';
    layer3_outputs(4716) <= layer2_outputs(5033);
    layer3_outputs(4717) <= not((layer2_outputs(6113)) or (layer2_outputs(6063)));
    layer3_outputs(4718) <= (layer2_outputs(981)) and (layer2_outputs(6398));
    layer3_outputs(4719) <= not(layer2_outputs(3678)) or (layer2_outputs(7039));
    layer3_outputs(4720) <= '1';
    layer3_outputs(4721) <= layer2_outputs(975);
    layer3_outputs(4722) <= '1';
    layer3_outputs(4723) <= not(layer2_outputs(4998));
    layer3_outputs(4724) <= '1';
    layer3_outputs(4725) <= not((layer2_outputs(5603)) or (layer2_outputs(7053)));
    layer3_outputs(4726) <= (layer2_outputs(7605)) and not (layer2_outputs(2966));
    layer3_outputs(4727) <= '0';
    layer3_outputs(4728) <= not(layer2_outputs(6608)) or (layer2_outputs(2764));
    layer3_outputs(4729) <= not((layer2_outputs(6139)) or (layer2_outputs(3100)));
    layer3_outputs(4730) <= layer2_outputs(6703);
    layer3_outputs(4731) <= (layer2_outputs(3718)) and (layer2_outputs(3998));
    layer3_outputs(4732) <= not(layer2_outputs(4569));
    layer3_outputs(4733) <= not(layer2_outputs(6035));
    layer3_outputs(4734) <= layer2_outputs(2387);
    layer3_outputs(4735) <= not(layer2_outputs(683));
    layer3_outputs(4736) <= (layer2_outputs(5090)) and not (layer2_outputs(6714));
    layer3_outputs(4737) <= '1';
    layer3_outputs(4738) <= not((layer2_outputs(7285)) and (layer2_outputs(2977)));
    layer3_outputs(4739) <= not(layer2_outputs(5444)) or (layer2_outputs(6103));
    layer3_outputs(4740) <= not(layer2_outputs(2507));
    layer3_outputs(4741) <= (layer2_outputs(4632)) and not (layer2_outputs(2481));
    layer3_outputs(4742) <= '1';
    layer3_outputs(4743) <= layer2_outputs(2716);
    layer3_outputs(4744) <= layer2_outputs(4346);
    layer3_outputs(4745) <= layer2_outputs(4084);
    layer3_outputs(4746) <= not(layer2_outputs(1628));
    layer3_outputs(4747) <= layer2_outputs(4721);
    layer3_outputs(4748) <= not((layer2_outputs(909)) or (layer2_outputs(1813)));
    layer3_outputs(4749) <= layer2_outputs(522);
    layer3_outputs(4750) <= (layer2_outputs(5938)) and not (layer2_outputs(3863));
    layer3_outputs(4751) <= not(layer2_outputs(6933)) or (layer2_outputs(1025));
    layer3_outputs(4752) <= '1';
    layer3_outputs(4753) <= not((layer2_outputs(1882)) or (layer2_outputs(4129)));
    layer3_outputs(4754) <= (layer2_outputs(4097)) and (layer2_outputs(1656));
    layer3_outputs(4755) <= (layer2_outputs(2381)) or (layer2_outputs(6639));
    layer3_outputs(4756) <= not((layer2_outputs(5470)) or (layer2_outputs(6472)));
    layer3_outputs(4757) <= layer2_outputs(5894);
    layer3_outputs(4758) <= (layer2_outputs(1954)) and not (layer2_outputs(6158));
    layer3_outputs(4759) <= (layer2_outputs(5232)) and not (layer2_outputs(2322));
    layer3_outputs(4760) <= (layer2_outputs(2740)) and not (layer2_outputs(3584));
    layer3_outputs(4761) <= not(layer2_outputs(3495));
    layer3_outputs(4762) <= layer2_outputs(280);
    layer3_outputs(4763) <= (layer2_outputs(1025)) and not (layer2_outputs(4293));
    layer3_outputs(4764) <= (layer2_outputs(3375)) and not (layer2_outputs(752));
    layer3_outputs(4765) <= '0';
    layer3_outputs(4766) <= '1';
    layer3_outputs(4767) <= (layer2_outputs(2106)) and not (layer2_outputs(4477));
    layer3_outputs(4768) <= not(layer2_outputs(4486));
    layer3_outputs(4769) <= layer2_outputs(3687);
    layer3_outputs(4770) <= not((layer2_outputs(1866)) or (layer2_outputs(2731)));
    layer3_outputs(4771) <= layer2_outputs(1282);
    layer3_outputs(4772) <= layer2_outputs(2257);
    layer3_outputs(4773) <= '0';
    layer3_outputs(4774) <= layer2_outputs(2195);
    layer3_outputs(4775) <= not((layer2_outputs(1832)) and (layer2_outputs(7656)));
    layer3_outputs(4776) <= not(layer2_outputs(6572));
    layer3_outputs(4777) <= (layer2_outputs(2591)) or (layer2_outputs(791));
    layer3_outputs(4778) <= '1';
    layer3_outputs(4779) <= (layer2_outputs(354)) and not (layer2_outputs(4130));
    layer3_outputs(4780) <= not((layer2_outputs(745)) and (layer2_outputs(4131)));
    layer3_outputs(4781) <= layer2_outputs(5329);
    layer3_outputs(4782) <= not(layer2_outputs(6010));
    layer3_outputs(4783) <= (layer2_outputs(5232)) or (layer2_outputs(1798));
    layer3_outputs(4784) <= '1';
    layer3_outputs(4785) <= not(layer2_outputs(4909));
    layer3_outputs(4786) <= (layer2_outputs(3608)) and not (layer2_outputs(2880));
    layer3_outputs(4787) <= layer2_outputs(3530);
    layer3_outputs(4788) <= layer2_outputs(491);
    layer3_outputs(4789) <= not((layer2_outputs(4606)) and (layer2_outputs(2529)));
    layer3_outputs(4790) <= layer2_outputs(2763);
    layer3_outputs(4791) <= not((layer2_outputs(5431)) and (layer2_outputs(3558)));
    layer3_outputs(4792) <= not(layer2_outputs(2859));
    layer3_outputs(4793) <= not((layer2_outputs(6631)) and (layer2_outputs(1101)));
    layer3_outputs(4794) <= not(layer2_outputs(3416));
    layer3_outputs(4795) <= (layer2_outputs(5810)) and not (layer2_outputs(2165));
    layer3_outputs(4796) <= (layer2_outputs(6261)) and not (layer2_outputs(6602));
    layer3_outputs(4797) <= layer2_outputs(945);
    layer3_outputs(4798) <= layer2_outputs(4659);
    layer3_outputs(4799) <= layer2_outputs(3679);
    layer3_outputs(4800) <= not(layer2_outputs(7330));
    layer3_outputs(4801) <= not(layer2_outputs(2156));
    layer3_outputs(4802) <= (layer2_outputs(1623)) and (layer2_outputs(6287));
    layer3_outputs(4803) <= (layer2_outputs(6447)) and (layer2_outputs(4830));
    layer3_outputs(4804) <= not(layer2_outputs(1615));
    layer3_outputs(4805) <= layer2_outputs(2868);
    layer3_outputs(4806) <= layer2_outputs(1872);
    layer3_outputs(4807) <= '1';
    layer3_outputs(4808) <= layer2_outputs(1527);
    layer3_outputs(4809) <= layer2_outputs(1875);
    layer3_outputs(4810) <= (layer2_outputs(2054)) and (layer2_outputs(3867));
    layer3_outputs(4811) <= not(layer2_outputs(2953));
    layer3_outputs(4812) <= not(layer2_outputs(6445));
    layer3_outputs(4813) <= not((layer2_outputs(7322)) or (layer2_outputs(1137)));
    layer3_outputs(4814) <= not(layer2_outputs(5830));
    layer3_outputs(4815) <= '1';
    layer3_outputs(4816) <= not(layer2_outputs(6085));
    layer3_outputs(4817) <= not((layer2_outputs(7410)) or (layer2_outputs(1301)));
    layer3_outputs(4818) <= not(layer2_outputs(4283)) or (layer2_outputs(2285));
    layer3_outputs(4819) <= '1';
    layer3_outputs(4820) <= not(layer2_outputs(5618));
    layer3_outputs(4821) <= (layer2_outputs(390)) and not (layer2_outputs(1772));
    layer3_outputs(4822) <= (layer2_outputs(7463)) or (layer2_outputs(4490));
    layer3_outputs(4823) <= (layer2_outputs(382)) or (layer2_outputs(1706));
    layer3_outputs(4824) <= layer2_outputs(4429);
    layer3_outputs(4825) <= not(layer2_outputs(3698));
    layer3_outputs(4826) <= not((layer2_outputs(2744)) and (layer2_outputs(1889)));
    layer3_outputs(4827) <= not(layer2_outputs(2504)) or (layer2_outputs(2185));
    layer3_outputs(4828) <= layer2_outputs(2582);
    layer3_outputs(4829) <= not(layer2_outputs(84));
    layer3_outputs(4830) <= not(layer2_outputs(6478));
    layer3_outputs(4831) <= (layer2_outputs(4843)) and not (layer2_outputs(1231));
    layer3_outputs(4832) <= not((layer2_outputs(7107)) or (layer2_outputs(4738)));
    layer3_outputs(4833) <= not((layer2_outputs(1778)) or (layer2_outputs(383)));
    layer3_outputs(4834) <= layer2_outputs(7579);
    layer3_outputs(4835) <= layer2_outputs(2293);
    layer3_outputs(4836) <= not(layer2_outputs(7127)) or (layer2_outputs(1632));
    layer3_outputs(4837) <= '0';
    layer3_outputs(4838) <= '0';
    layer3_outputs(4839) <= '0';
    layer3_outputs(4840) <= layer2_outputs(4160);
    layer3_outputs(4841) <= not(layer2_outputs(5818)) or (layer2_outputs(2919));
    layer3_outputs(4842) <= not(layer2_outputs(251));
    layer3_outputs(4843) <= not(layer2_outputs(1286)) or (layer2_outputs(2456));
    layer3_outputs(4844) <= (layer2_outputs(6074)) and not (layer2_outputs(3773));
    layer3_outputs(4845) <= '1';
    layer3_outputs(4846) <= not(layer2_outputs(5546)) or (layer2_outputs(2428));
    layer3_outputs(4847) <= (layer2_outputs(2969)) and not (layer2_outputs(4338));
    layer3_outputs(4848) <= (layer2_outputs(2172)) and (layer2_outputs(4760));
    layer3_outputs(4849) <= not(layer2_outputs(5344));
    layer3_outputs(4850) <= (layer2_outputs(5660)) or (layer2_outputs(4937));
    layer3_outputs(4851) <= not(layer2_outputs(7327)) or (layer2_outputs(2470));
    layer3_outputs(4852) <= (layer2_outputs(988)) and (layer2_outputs(592));
    layer3_outputs(4853) <= (layer2_outputs(2341)) and (layer2_outputs(7187));
    layer3_outputs(4854) <= layer2_outputs(3647);
    layer3_outputs(4855) <= not(layer2_outputs(2003));
    layer3_outputs(4856) <= (layer2_outputs(867)) and not (layer2_outputs(2029));
    layer3_outputs(4857) <= (layer2_outputs(3511)) and not (layer2_outputs(1400));
    layer3_outputs(4858) <= '1';
    layer3_outputs(4859) <= (layer2_outputs(3302)) and (layer2_outputs(7062));
    layer3_outputs(4860) <= not((layer2_outputs(5725)) xor (layer2_outputs(7038)));
    layer3_outputs(4861) <= not((layer2_outputs(6944)) and (layer2_outputs(541)));
    layer3_outputs(4862) <= layer2_outputs(369);
    layer3_outputs(4863) <= (layer2_outputs(5319)) and not (layer2_outputs(2629));
    layer3_outputs(4864) <= not(layer2_outputs(3117));
    layer3_outputs(4865) <= (layer2_outputs(6477)) or (layer2_outputs(1534));
    layer3_outputs(4866) <= layer2_outputs(7445);
    layer3_outputs(4867) <= (layer2_outputs(7184)) and (layer2_outputs(5735));
    layer3_outputs(4868) <= layer2_outputs(2234);
    layer3_outputs(4869) <= '0';
    layer3_outputs(4870) <= not(layer2_outputs(7109)) or (layer2_outputs(4157));
    layer3_outputs(4871) <= not(layer2_outputs(2040)) or (layer2_outputs(566));
    layer3_outputs(4872) <= (layer2_outputs(4196)) and (layer2_outputs(5034));
    layer3_outputs(4873) <= not(layer2_outputs(3623));
    layer3_outputs(4874) <= (layer2_outputs(3050)) and not (layer2_outputs(7572));
    layer3_outputs(4875) <= not(layer2_outputs(2340));
    layer3_outputs(4876) <= not(layer2_outputs(2829));
    layer3_outputs(4877) <= '0';
    layer3_outputs(4878) <= (layer2_outputs(5570)) or (layer2_outputs(6629));
    layer3_outputs(4879) <= '1';
    layer3_outputs(4880) <= (layer2_outputs(329)) and not (layer2_outputs(3731));
    layer3_outputs(4881) <= layer2_outputs(3552);
    layer3_outputs(4882) <= layer2_outputs(30);
    layer3_outputs(4883) <= (layer2_outputs(4807)) and not (layer2_outputs(1532));
    layer3_outputs(4884) <= layer2_outputs(5523);
    layer3_outputs(4885) <= '0';
    layer3_outputs(4886) <= '1';
    layer3_outputs(4887) <= not(layer2_outputs(2779));
    layer3_outputs(4888) <= '1';
    layer3_outputs(4889) <= layer2_outputs(2196);
    layer3_outputs(4890) <= (layer2_outputs(5749)) and not (layer2_outputs(2966));
    layer3_outputs(4891) <= layer2_outputs(4811);
    layer3_outputs(4892) <= layer2_outputs(3276);
    layer3_outputs(4893) <= '0';
    layer3_outputs(4894) <= not((layer2_outputs(2928)) or (layer2_outputs(6254)));
    layer3_outputs(4895) <= not(layer2_outputs(1539));
    layer3_outputs(4896) <= (layer2_outputs(1122)) and (layer2_outputs(1525));
    layer3_outputs(4897) <= (layer2_outputs(4942)) xor (layer2_outputs(6498));
    layer3_outputs(4898) <= not((layer2_outputs(6589)) xor (layer2_outputs(3380)));
    layer3_outputs(4899) <= layer2_outputs(6131);
    layer3_outputs(4900) <= not(layer2_outputs(2210));
    layer3_outputs(4901) <= layer2_outputs(786);
    layer3_outputs(4902) <= not(layer2_outputs(6351));
    layer3_outputs(4903) <= layer2_outputs(5155);
    layer3_outputs(4904) <= not(layer2_outputs(2218));
    layer3_outputs(4905) <= layer2_outputs(7424);
    layer3_outputs(4906) <= '0';
    layer3_outputs(4907) <= not(layer2_outputs(318)) or (layer2_outputs(2888));
    layer3_outputs(4908) <= (layer2_outputs(2693)) or (layer2_outputs(2811));
    layer3_outputs(4909) <= layer2_outputs(6547);
    layer3_outputs(4910) <= not(layer2_outputs(3365));
    layer3_outputs(4911) <= '1';
    layer3_outputs(4912) <= not(layer2_outputs(4758));
    layer3_outputs(4913) <= not(layer2_outputs(473));
    layer3_outputs(4914) <= '1';
    layer3_outputs(4915) <= (layer2_outputs(4360)) and not (layer2_outputs(2314));
    layer3_outputs(4916) <= not((layer2_outputs(4150)) or (layer2_outputs(5541)));
    layer3_outputs(4917) <= layer2_outputs(1566);
    layer3_outputs(4918) <= not(layer2_outputs(3078));
    layer3_outputs(4919) <= not((layer2_outputs(6919)) or (layer2_outputs(5870)));
    layer3_outputs(4920) <= (layer2_outputs(5145)) and (layer2_outputs(7337));
    layer3_outputs(4921) <= not(layer2_outputs(5764));
    layer3_outputs(4922) <= layer2_outputs(1837);
    layer3_outputs(4923) <= '1';
    layer3_outputs(4924) <= '1';
    layer3_outputs(4925) <= '0';
    layer3_outputs(4926) <= (layer2_outputs(1489)) and not (layer2_outputs(3127));
    layer3_outputs(4927) <= not((layer2_outputs(5792)) or (layer2_outputs(3798)));
    layer3_outputs(4928) <= not(layer2_outputs(4883));
    layer3_outputs(4929) <= (layer2_outputs(4831)) and not (layer2_outputs(2519));
    layer3_outputs(4930) <= not((layer2_outputs(664)) and (layer2_outputs(5023)));
    layer3_outputs(4931) <= not(layer2_outputs(7037)) or (layer2_outputs(414));
    layer3_outputs(4932) <= (layer2_outputs(4881)) and not (layer2_outputs(569));
    layer3_outputs(4933) <= not(layer2_outputs(5323)) or (layer2_outputs(4166));
    layer3_outputs(4934) <= layer2_outputs(6772);
    layer3_outputs(4935) <= (layer2_outputs(6129)) and not (layer2_outputs(4854));
    layer3_outputs(4936) <= (layer2_outputs(1984)) and not (layer2_outputs(5723));
    layer3_outputs(4937) <= (layer2_outputs(1951)) xor (layer2_outputs(4877));
    layer3_outputs(4938) <= (layer2_outputs(4112)) and not (layer2_outputs(3280));
    layer3_outputs(4939) <= (layer2_outputs(4562)) or (layer2_outputs(2178));
    layer3_outputs(4940) <= not((layer2_outputs(6322)) xor (layer2_outputs(7152)));
    layer3_outputs(4941) <= (layer2_outputs(5229)) and (layer2_outputs(5739));
    layer3_outputs(4942) <= layer2_outputs(6938);
    layer3_outputs(4943) <= not(layer2_outputs(5081));
    layer3_outputs(4944) <= '1';
    layer3_outputs(4945) <= (layer2_outputs(5656)) or (layer2_outputs(2459));
    layer3_outputs(4946) <= '1';
    layer3_outputs(4947) <= '0';
    layer3_outputs(4948) <= not(layer2_outputs(548)) or (layer2_outputs(4398));
    layer3_outputs(4949) <= layer2_outputs(1350);
    layer3_outputs(4950) <= layer2_outputs(7601);
    layer3_outputs(4951) <= not(layer2_outputs(408));
    layer3_outputs(4952) <= '1';
    layer3_outputs(4953) <= (layer2_outputs(5387)) xor (layer2_outputs(472));
    layer3_outputs(4954) <= not(layer2_outputs(7620));
    layer3_outputs(4955) <= not(layer2_outputs(3069));
    layer3_outputs(4956) <= (layer2_outputs(1414)) and (layer2_outputs(6161));
    layer3_outputs(4957) <= (layer2_outputs(4560)) and not (layer2_outputs(545));
    layer3_outputs(4958) <= not(layer2_outputs(629));
    layer3_outputs(4959) <= not(layer2_outputs(3681));
    layer3_outputs(4960) <= (layer2_outputs(5791)) and not (layer2_outputs(4755));
    layer3_outputs(4961) <= not((layer2_outputs(2669)) and (layer2_outputs(1557)));
    layer3_outputs(4962) <= layer2_outputs(7360);
    layer3_outputs(4963) <= (layer2_outputs(6118)) and not (layer2_outputs(3023));
    layer3_outputs(4964) <= not(layer2_outputs(1785));
    layer3_outputs(4965) <= (layer2_outputs(4977)) and (layer2_outputs(2264));
    layer3_outputs(4966) <= not(layer2_outputs(292));
    layer3_outputs(4967) <= not(layer2_outputs(6578));
    layer3_outputs(4968) <= (layer2_outputs(5090)) and not (layer2_outputs(437));
    layer3_outputs(4969) <= not(layer2_outputs(385)) or (layer2_outputs(2477));
    layer3_outputs(4970) <= (layer2_outputs(489)) and not (layer2_outputs(4921));
    layer3_outputs(4971) <= not(layer2_outputs(2114)) or (layer2_outputs(847));
    layer3_outputs(4972) <= not((layer2_outputs(75)) or (layer2_outputs(1108)));
    layer3_outputs(4973) <= not(layer2_outputs(1824));
    layer3_outputs(4974) <= '0';
    layer3_outputs(4975) <= not(layer2_outputs(4557));
    layer3_outputs(4976) <= not(layer2_outputs(4909)) or (layer2_outputs(6292));
    layer3_outputs(4977) <= (layer2_outputs(1240)) and not (layer2_outputs(5381));
    layer3_outputs(4978) <= layer2_outputs(7585);
    layer3_outputs(4979) <= not(layer2_outputs(134)) or (layer2_outputs(623));
    layer3_outputs(4980) <= layer2_outputs(6091);
    layer3_outputs(4981) <= layer2_outputs(1589);
    layer3_outputs(4982) <= '1';
    layer3_outputs(4983) <= not(layer2_outputs(5290));
    layer3_outputs(4984) <= not(layer2_outputs(4761)) or (layer2_outputs(423));
    layer3_outputs(4985) <= (layer2_outputs(6532)) or (layer2_outputs(4212));
    layer3_outputs(4986) <= not((layer2_outputs(7599)) xor (layer2_outputs(6869)));
    layer3_outputs(4987) <= not(layer2_outputs(215));
    layer3_outputs(4988) <= not((layer2_outputs(7529)) or (layer2_outputs(6236)));
    layer3_outputs(4989) <= layer2_outputs(58);
    layer3_outputs(4990) <= (layer2_outputs(1700)) and (layer2_outputs(2713));
    layer3_outputs(4991) <= not(layer2_outputs(7519));
    layer3_outputs(4992) <= '0';
    layer3_outputs(4993) <= (layer2_outputs(4204)) and not (layer2_outputs(7670));
    layer3_outputs(4994) <= layer2_outputs(4333);
    layer3_outputs(4995) <= (layer2_outputs(4279)) and not (layer2_outputs(469));
    layer3_outputs(4996) <= not((layer2_outputs(3887)) and (layer2_outputs(3383)));
    layer3_outputs(4997) <= not(layer2_outputs(196));
    layer3_outputs(4998) <= (layer2_outputs(1750)) and not (layer2_outputs(368));
    layer3_outputs(4999) <= not((layer2_outputs(3925)) and (layer2_outputs(668)));
    layer3_outputs(5000) <= layer2_outputs(7633);
    layer3_outputs(5001) <= not(layer2_outputs(5379));
    layer3_outputs(5002) <= '0';
    layer3_outputs(5003) <= (layer2_outputs(1253)) or (layer2_outputs(3958));
    layer3_outputs(5004) <= (layer2_outputs(1871)) and (layer2_outputs(3322));
    layer3_outputs(5005) <= not((layer2_outputs(1642)) and (layer2_outputs(3846)));
    layer3_outputs(5006) <= (layer2_outputs(5984)) and not (layer2_outputs(1250));
    layer3_outputs(5007) <= not(layer2_outputs(7438));
    layer3_outputs(5008) <= layer2_outputs(5273);
    layer3_outputs(5009) <= not(layer2_outputs(2451)) or (layer2_outputs(6617));
    layer3_outputs(5010) <= not((layer2_outputs(6526)) xor (layer2_outputs(4608)));
    layer3_outputs(5011) <= '0';
    layer3_outputs(5012) <= not(layer2_outputs(5021));
    layer3_outputs(5013) <= layer2_outputs(5604);
    layer3_outputs(5014) <= not(layer2_outputs(4587));
    layer3_outputs(5015) <= not(layer2_outputs(2656)) or (layer2_outputs(7298));
    layer3_outputs(5016) <= not((layer2_outputs(1687)) and (layer2_outputs(3950)));
    layer3_outputs(5017) <= '0';
    layer3_outputs(5018) <= not(layer2_outputs(1031)) or (layer2_outputs(4552));
    layer3_outputs(5019) <= (layer2_outputs(5860)) xor (layer2_outputs(3412));
    layer3_outputs(5020) <= layer2_outputs(2712);
    layer3_outputs(5021) <= layer2_outputs(3199);
    layer3_outputs(5022) <= not(layer2_outputs(6492)) or (layer2_outputs(6766));
    layer3_outputs(5023) <= not((layer2_outputs(2601)) or (layer2_outputs(1571)));
    layer3_outputs(5024) <= '0';
    layer3_outputs(5025) <= layer2_outputs(4225);
    layer3_outputs(5026) <= layer2_outputs(6208);
    layer3_outputs(5027) <= not(layer2_outputs(2430)) or (layer2_outputs(884));
    layer3_outputs(5028) <= not(layer2_outputs(783)) or (layer2_outputs(1027));
    layer3_outputs(5029) <= not((layer2_outputs(2628)) or (layer2_outputs(7070)));
    layer3_outputs(5030) <= not(layer2_outputs(7157));
    layer3_outputs(5031) <= not(layer2_outputs(5910));
    layer3_outputs(5032) <= layer2_outputs(2375);
    layer3_outputs(5033) <= (layer2_outputs(4283)) xor (layer2_outputs(4494));
    layer3_outputs(5034) <= layer2_outputs(5158);
    layer3_outputs(5035) <= '1';
    layer3_outputs(5036) <= (layer2_outputs(3907)) and not (layer2_outputs(5506));
    layer3_outputs(5037) <= layer2_outputs(4983);
    layer3_outputs(5038) <= not((layer2_outputs(5704)) xor (layer2_outputs(2385)));
    layer3_outputs(5039) <= (layer2_outputs(2602)) and not (layer2_outputs(1895));
    layer3_outputs(5040) <= not((layer2_outputs(1702)) and (layer2_outputs(1523)));
    layer3_outputs(5041) <= layer2_outputs(7400);
    layer3_outputs(5042) <= layer2_outputs(1837);
    layer3_outputs(5043) <= (layer2_outputs(1093)) and not (layer2_outputs(137));
    layer3_outputs(5044) <= not(layer2_outputs(7476)) or (layer2_outputs(2544));
    layer3_outputs(5045) <= not(layer2_outputs(4873));
    layer3_outputs(5046) <= not((layer2_outputs(6757)) or (layer2_outputs(998)));
    layer3_outputs(5047) <= (layer2_outputs(2622)) or (layer2_outputs(2834));
    layer3_outputs(5048) <= not(layer2_outputs(3978));
    layer3_outputs(5049) <= (layer2_outputs(1342)) and not (layer2_outputs(6860));
    layer3_outputs(5050) <= not(layer2_outputs(789));
    layer3_outputs(5051) <= not((layer2_outputs(1277)) and (layer2_outputs(2191)));
    layer3_outputs(5052) <= not(layer2_outputs(7171));
    layer3_outputs(5053) <= not((layer2_outputs(5343)) or (layer2_outputs(6257)));
    layer3_outputs(5054) <= layer2_outputs(2255);
    layer3_outputs(5055) <= not((layer2_outputs(7119)) and (layer2_outputs(5942)));
    layer3_outputs(5056) <= '1';
    layer3_outputs(5057) <= (layer2_outputs(1658)) and (layer2_outputs(5239));
    layer3_outputs(5058) <= not(layer2_outputs(1574));
    layer3_outputs(5059) <= '0';
    layer3_outputs(5060) <= (layer2_outputs(5315)) and (layer2_outputs(5195));
    layer3_outputs(5061) <= '1';
    layer3_outputs(5062) <= (layer2_outputs(6501)) or (layer2_outputs(1368));
    layer3_outputs(5063) <= layer2_outputs(4799);
    layer3_outputs(5064) <= '1';
    layer3_outputs(5065) <= not((layer2_outputs(1603)) and (layer2_outputs(5866)));
    layer3_outputs(5066) <= not(layer2_outputs(6353)) or (layer2_outputs(7112));
    layer3_outputs(5067) <= '1';
    layer3_outputs(5068) <= not(layer2_outputs(4458)) or (layer2_outputs(4047));
    layer3_outputs(5069) <= (layer2_outputs(6304)) and not (layer2_outputs(5680));
    layer3_outputs(5070) <= layer2_outputs(2241);
    layer3_outputs(5071) <= '0';
    layer3_outputs(5072) <= (layer2_outputs(714)) and not (layer2_outputs(3462));
    layer3_outputs(5073) <= '1';
    layer3_outputs(5074) <= (layer2_outputs(3802)) xor (layer2_outputs(280));
    layer3_outputs(5075) <= (layer2_outputs(3058)) and (layer2_outputs(5512));
    layer3_outputs(5076) <= not((layer2_outputs(6686)) xor (layer2_outputs(5828)));
    layer3_outputs(5077) <= '1';
    layer3_outputs(5078) <= (layer2_outputs(7117)) xor (layer2_outputs(1285));
    layer3_outputs(5079) <= layer2_outputs(1873);
    layer3_outputs(5080) <= (layer2_outputs(3650)) and not (layer2_outputs(6209));
    layer3_outputs(5081) <= layer2_outputs(3212);
    layer3_outputs(5082) <= layer2_outputs(1876);
    layer3_outputs(5083) <= not(layer2_outputs(1916));
    layer3_outputs(5084) <= not(layer2_outputs(466));
    layer3_outputs(5085) <= (layer2_outputs(2129)) xor (layer2_outputs(2547));
    layer3_outputs(5086) <= (layer2_outputs(4478)) and (layer2_outputs(2274));
    layer3_outputs(5087) <= not(layer2_outputs(161)) or (layer2_outputs(518));
    layer3_outputs(5088) <= layer2_outputs(1527);
    layer3_outputs(5089) <= (layer2_outputs(1050)) or (layer2_outputs(7665));
    layer3_outputs(5090) <= not(layer2_outputs(3882)) or (layer2_outputs(2756));
    layer3_outputs(5091) <= not(layer2_outputs(7288));
    layer3_outputs(5092) <= not(layer2_outputs(5272)) or (layer2_outputs(4429));
    layer3_outputs(5093) <= not(layer2_outputs(2632)) or (layer2_outputs(2064));
    layer3_outputs(5094) <= '1';
    layer3_outputs(5095) <= layer2_outputs(5772);
    layer3_outputs(5096) <= layer2_outputs(316);
    layer3_outputs(5097) <= not((layer2_outputs(559)) and (layer2_outputs(5863)));
    layer3_outputs(5098) <= not(layer2_outputs(7662));
    layer3_outputs(5099) <= '0';
    layer3_outputs(5100) <= not((layer2_outputs(5940)) xor (layer2_outputs(1039)));
    layer3_outputs(5101) <= not(layer2_outputs(6135));
    layer3_outputs(5102) <= not((layer2_outputs(3901)) or (layer2_outputs(3791)));
    layer3_outputs(5103) <= layer2_outputs(1586);
    layer3_outputs(5104) <= not(layer2_outputs(6487));
    layer3_outputs(5105) <= '1';
    layer3_outputs(5106) <= '0';
    layer3_outputs(5107) <= not((layer2_outputs(5841)) or (layer2_outputs(3410)));
    layer3_outputs(5108) <= '1';
    layer3_outputs(5109) <= (layer2_outputs(571)) and not (layer2_outputs(2455));
    layer3_outputs(5110) <= (layer2_outputs(1112)) and not (layer2_outputs(888));
    layer3_outputs(5111) <= not(layer2_outputs(4034));
    layer3_outputs(5112) <= '0';
    layer3_outputs(5113) <= not(layer2_outputs(7626)) or (layer2_outputs(1058));
    layer3_outputs(5114) <= layer2_outputs(1555);
    layer3_outputs(5115) <= '1';
    layer3_outputs(5116) <= not(layer2_outputs(1175)) or (layer2_outputs(5037));
    layer3_outputs(5117) <= layer2_outputs(510);
    layer3_outputs(5118) <= (layer2_outputs(7444)) and not (layer2_outputs(2427));
    layer3_outputs(5119) <= (layer2_outputs(4690)) or (layer2_outputs(3760));
    layer3_outputs(5120) <= (layer2_outputs(7421)) and (layer2_outputs(3362));
    layer3_outputs(5121) <= layer2_outputs(4579);
    layer3_outputs(5122) <= (layer2_outputs(2443)) and not (layer2_outputs(2014));
    layer3_outputs(5123) <= not(layer2_outputs(1198)) or (layer2_outputs(5160));
    layer3_outputs(5124) <= not(layer2_outputs(6715));
    layer3_outputs(5125) <= not((layer2_outputs(1817)) and (layer2_outputs(2962)));
    layer3_outputs(5126) <= layer2_outputs(3333);
    layer3_outputs(5127) <= (layer2_outputs(71)) and (layer2_outputs(1508));
    layer3_outputs(5128) <= '1';
    layer3_outputs(5129) <= (layer2_outputs(7669)) and not (layer2_outputs(5095));
    layer3_outputs(5130) <= not(layer2_outputs(6144)) or (layer2_outputs(7019));
    layer3_outputs(5131) <= not((layer2_outputs(4617)) or (layer2_outputs(4801)));
    layer3_outputs(5132) <= layer2_outputs(1127);
    layer3_outputs(5133) <= not(layer2_outputs(1858));
    layer3_outputs(5134) <= not(layer2_outputs(2276)) or (layer2_outputs(3529));
    layer3_outputs(5135) <= not((layer2_outputs(1365)) and (layer2_outputs(1666)));
    layer3_outputs(5136) <= not(layer2_outputs(6681)) or (layer2_outputs(2976));
    layer3_outputs(5137) <= not(layer2_outputs(5872));
    layer3_outputs(5138) <= '0';
    layer3_outputs(5139) <= layer2_outputs(2992);
    layer3_outputs(5140) <= layer2_outputs(8);
    layer3_outputs(5141) <= '1';
    layer3_outputs(5142) <= (layer2_outputs(730)) and not (layer2_outputs(7382));
    layer3_outputs(5143) <= not(layer2_outputs(5252));
    layer3_outputs(5144) <= (layer2_outputs(6805)) and not (layer2_outputs(3889));
    layer3_outputs(5145) <= not(layer2_outputs(5508));
    layer3_outputs(5146) <= '1';
    layer3_outputs(5147) <= layer2_outputs(2207);
    layer3_outputs(5148) <= not(layer2_outputs(2094)) or (layer2_outputs(4142));
    layer3_outputs(5149) <= layer2_outputs(3521);
    layer3_outputs(5150) <= (layer2_outputs(677)) xor (layer2_outputs(5543));
    layer3_outputs(5151) <= '0';
    layer3_outputs(5152) <= not((layer2_outputs(3602)) and (layer2_outputs(4747)));
    layer3_outputs(5153) <= (layer2_outputs(2762)) and (layer2_outputs(4957));
    layer3_outputs(5154) <= not(layer2_outputs(377)) or (layer2_outputs(6884));
    layer3_outputs(5155) <= not(layer2_outputs(2479)) or (layer2_outputs(4737));
    layer3_outputs(5156) <= (layer2_outputs(5121)) or (layer2_outputs(6173));
    layer3_outputs(5157) <= not((layer2_outputs(5388)) xor (layer2_outputs(957)));
    layer3_outputs(5158) <= not(layer2_outputs(1799));
    layer3_outputs(5159) <= not(layer2_outputs(7122)) or (layer2_outputs(694));
    layer3_outputs(5160) <= layer2_outputs(1926);
    layer3_outputs(5161) <= (layer2_outputs(6048)) and not (layer2_outputs(5373));
    layer3_outputs(5162) <= '1';
    layer3_outputs(5163) <= not((layer2_outputs(5042)) and (layer2_outputs(5917)));
    layer3_outputs(5164) <= not(layer2_outputs(1453));
    layer3_outputs(5165) <= (layer2_outputs(7543)) and not (layer2_outputs(3876));
    layer3_outputs(5166) <= not(layer2_outputs(3843));
    layer3_outputs(5167) <= (layer2_outputs(953)) and (layer2_outputs(5263));
    layer3_outputs(5168) <= not(layer2_outputs(448));
    layer3_outputs(5169) <= not((layer2_outputs(6599)) or (layer2_outputs(1794)));
    layer3_outputs(5170) <= '0';
    layer3_outputs(5171) <= not(layer2_outputs(1946));
    layer3_outputs(5172) <= '0';
    layer3_outputs(5173) <= layer2_outputs(3403);
    layer3_outputs(5174) <= (layer2_outputs(4033)) and not (layer2_outputs(6069));
    layer3_outputs(5175) <= '1';
    layer3_outputs(5176) <= not(layer2_outputs(4204)) or (layer2_outputs(2965));
    layer3_outputs(5177) <= not(layer2_outputs(5769)) or (layer2_outputs(4108));
    layer3_outputs(5178) <= not(layer2_outputs(3)) or (layer2_outputs(4236));
    layer3_outputs(5179) <= not(layer2_outputs(5209));
    layer3_outputs(5180) <= not(layer2_outputs(1133)) or (layer2_outputs(774));
    layer3_outputs(5181) <= not((layer2_outputs(6978)) and (layer2_outputs(6256)));
    layer3_outputs(5182) <= '1';
    layer3_outputs(5183) <= not(layer2_outputs(7012));
    layer3_outputs(5184) <= not(layer2_outputs(4691));
    layer3_outputs(5185) <= '0';
    layer3_outputs(5186) <= (layer2_outputs(861)) or (layer2_outputs(1765));
    layer3_outputs(5187) <= layer2_outputs(3941);
    layer3_outputs(5188) <= layer2_outputs(6397);
    layer3_outputs(5189) <= not(layer2_outputs(2470)) or (layer2_outputs(1594));
    layer3_outputs(5190) <= not((layer2_outputs(2959)) or (layer2_outputs(1641)));
    layer3_outputs(5191) <= layer2_outputs(1879);
    layer3_outputs(5192) <= not((layer2_outputs(6795)) and (layer2_outputs(1729)));
    layer3_outputs(5193) <= (layer2_outputs(4537)) and (layer2_outputs(4195));
    layer3_outputs(5194) <= layer2_outputs(1763);
    layer3_outputs(5195) <= (layer2_outputs(1659)) and not (layer2_outputs(5039));
    layer3_outputs(5196) <= (layer2_outputs(3653)) and not (layer2_outputs(143));
    layer3_outputs(5197) <= not((layer2_outputs(7123)) xor (layer2_outputs(1087)));
    layer3_outputs(5198) <= layer2_outputs(7082);
    layer3_outputs(5199) <= '1';
    layer3_outputs(5200) <= not(layer2_outputs(1001));
    layer3_outputs(5201) <= layer2_outputs(3964);
    layer3_outputs(5202) <= '1';
    layer3_outputs(5203) <= not(layer2_outputs(3980));
    layer3_outputs(5204) <= not((layer2_outputs(5790)) and (layer2_outputs(4973)));
    layer3_outputs(5205) <= layer2_outputs(7267);
    layer3_outputs(5206) <= not(layer2_outputs(4741));
    layer3_outputs(5207) <= not(layer2_outputs(165));
    layer3_outputs(5208) <= not((layer2_outputs(2067)) or (layer2_outputs(4012)));
    layer3_outputs(5209) <= not((layer2_outputs(179)) or (layer2_outputs(6764)));
    layer3_outputs(5210) <= not(layer2_outputs(4043));
    layer3_outputs(5211) <= (layer2_outputs(2490)) and not (layer2_outputs(1165));
    layer3_outputs(5212) <= (layer2_outputs(2293)) or (layer2_outputs(1074));
    layer3_outputs(5213) <= not(layer2_outputs(2620)) or (layer2_outputs(1505));
    layer3_outputs(5214) <= '0';
    layer3_outputs(5215) <= not(layer2_outputs(6485));
    layer3_outputs(5216) <= (layer2_outputs(494)) and not (layer2_outputs(2645));
    layer3_outputs(5217) <= (layer2_outputs(908)) and (layer2_outputs(5899));
    layer3_outputs(5218) <= layer2_outputs(2456);
    layer3_outputs(5219) <= layer2_outputs(4372);
    layer3_outputs(5220) <= layer2_outputs(4095);
    layer3_outputs(5221) <= layer2_outputs(2552);
    layer3_outputs(5222) <= (layer2_outputs(2566)) and (layer2_outputs(5269));
    layer3_outputs(5223) <= not(layer2_outputs(6803));
    layer3_outputs(5224) <= not(layer2_outputs(6022));
    layer3_outputs(5225) <= not(layer2_outputs(1994)) or (layer2_outputs(3176));
    layer3_outputs(5226) <= (layer2_outputs(5413)) or (layer2_outputs(5609));
    layer3_outputs(5227) <= (layer2_outputs(7042)) or (layer2_outputs(1322));
    layer3_outputs(5228) <= not(layer2_outputs(2815));
    layer3_outputs(5229) <= layer2_outputs(2848);
    layer3_outputs(5230) <= not(layer2_outputs(1880)) or (layer2_outputs(7454));
    layer3_outputs(5231) <= (layer2_outputs(2444)) and not (layer2_outputs(1183));
    layer3_outputs(5232) <= (layer2_outputs(5638)) and not (layer2_outputs(7600));
    layer3_outputs(5233) <= not(layer2_outputs(2600)) or (layer2_outputs(6775));
    layer3_outputs(5234) <= '0';
    layer3_outputs(5235) <= not(layer2_outputs(1717)) or (layer2_outputs(3707));
    layer3_outputs(5236) <= layer2_outputs(6444);
    layer3_outputs(5237) <= (layer2_outputs(1770)) or (layer2_outputs(1429));
    layer3_outputs(5238) <= not(layer2_outputs(2318)) or (layer2_outputs(1342));
    layer3_outputs(5239) <= not(layer2_outputs(4676));
    layer3_outputs(5240) <= not((layer2_outputs(6914)) and (layer2_outputs(1557)));
    layer3_outputs(5241) <= layer2_outputs(2654);
    layer3_outputs(5242) <= layer2_outputs(655);
    layer3_outputs(5243) <= (layer2_outputs(3911)) and not (layer2_outputs(7086));
    layer3_outputs(5244) <= not(layer2_outputs(4473));
    layer3_outputs(5245) <= '1';
    layer3_outputs(5246) <= '1';
    layer3_outputs(5247) <= '1';
    layer3_outputs(5248) <= (layer2_outputs(4600)) or (layer2_outputs(5313));
    layer3_outputs(5249) <= not(layer2_outputs(7492));
    layer3_outputs(5250) <= not(layer2_outputs(7265));
    layer3_outputs(5251) <= not((layer2_outputs(536)) and (layer2_outputs(4358)));
    layer3_outputs(5252) <= not(layer2_outputs(664)) or (layer2_outputs(6427));
    layer3_outputs(5253) <= not(layer2_outputs(4739));
    layer3_outputs(5254) <= (layer2_outputs(202)) and not (layer2_outputs(3250));
    layer3_outputs(5255) <= not(layer2_outputs(6451)) or (layer2_outputs(2220));
    layer3_outputs(5256) <= '0';
    layer3_outputs(5257) <= '0';
    layer3_outputs(5258) <= (layer2_outputs(7540)) and not (layer2_outputs(5733));
    layer3_outputs(5259) <= '1';
    layer3_outputs(5260) <= not(layer2_outputs(5456));
    layer3_outputs(5261) <= not(layer2_outputs(7430));
    layer3_outputs(5262) <= (layer2_outputs(6777)) and not (layer2_outputs(7389));
    layer3_outputs(5263) <= not(layer2_outputs(2245));
    layer3_outputs(5264) <= (layer2_outputs(741)) and not (layer2_outputs(2076));
    layer3_outputs(5265) <= layer2_outputs(2383);
    layer3_outputs(5266) <= not(layer2_outputs(5559)) or (layer2_outputs(4203));
    layer3_outputs(5267) <= not(layer2_outputs(2909));
    layer3_outputs(5268) <= '0';
    layer3_outputs(5269) <= layer2_outputs(4354);
    layer3_outputs(5270) <= not((layer2_outputs(7022)) or (layer2_outputs(4888)));
    layer3_outputs(5271) <= layer2_outputs(3596);
    layer3_outputs(5272) <= '1';
    layer3_outputs(5273) <= not(layer2_outputs(3045));
    layer3_outputs(5274) <= layer2_outputs(1432);
    layer3_outputs(5275) <= '0';
    layer3_outputs(5276) <= layer2_outputs(48);
    layer3_outputs(5277) <= layer2_outputs(5270);
    layer3_outputs(5278) <= (layer2_outputs(5695)) and not (layer2_outputs(4885));
    layer3_outputs(5279) <= not((layer2_outputs(3732)) or (layer2_outputs(6862)));
    layer3_outputs(5280) <= '0';
    layer3_outputs(5281) <= not((layer2_outputs(7057)) and (layer2_outputs(301)));
    layer3_outputs(5282) <= not((layer2_outputs(3275)) or (layer2_outputs(618)));
    layer3_outputs(5283) <= (layer2_outputs(2559)) and (layer2_outputs(6262));
    layer3_outputs(5284) <= (layer2_outputs(2193)) or (layer2_outputs(2674));
    layer3_outputs(5285) <= not(layer2_outputs(4334));
    layer3_outputs(5286) <= (layer2_outputs(2600)) and not (layer2_outputs(3626));
    layer3_outputs(5287) <= '0';
    layer3_outputs(5288) <= not(layer2_outputs(5747));
    layer3_outputs(5289) <= (layer2_outputs(3059)) and (layer2_outputs(2247));
    layer3_outputs(5290) <= (layer2_outputs(6835)) and not (layer2_outputs(2954));
    layer3_outputs(5291) <= (layer2_outputs(6587)) and not (layer2_outputs(4833));
    layer3_outputs(5292) <= '1';
    layer3_outputs(5293) <= '1';
    layer3_outputs(5294) <= not((layer2_outputs(4067)) or (layer2_outputs(251)));
    layer3_outputs(5295) <= (layer2_outputs(560)) and (layer2_outputs(708));
    layer3_outputs(5296) <= not((layer2_outputs(3805)) or (layer2_outputs(7133)));
    layer3_outputs(5297) <= not((layer2_outputs(2979)) and (layer2_outputs(3854)));
    layer3_outputs(5298) <= (layer2_outputs(822)) and not (layer2_outputs(4376));
    layer3_outputs(5299) <= layer2_outputs(3713);
    layer3_outputs(5300) <= '1';
    layer3_outputs(5301) <= layer2_outputs(6739);
    layer3_outputs(5302) <= layer2_outputs(2457);
    layer3_outputs(5303) <= layer2_outputs(269);
    layer3_outputs(5304) <= not(layer2_outputs(5015)) or (layer2_outputs(522));
    layer3_outputs(5305) <= layer2_outputs(3140);
    layer3_outputs(5306) <= layer2_outputs(6582);
    layer3_outputs(5307) <= (layer2_outputs(7598)) and (layer2_outputs(2381));
    layer3_outputs(5308) <= not(layer2_outputs(6280));
    layer3_outputs(5309) <= (layer2_outputs(4224)) and not (layer2_outputs(7102));
    layer3_outputs(5310) <= not((layer2_outputs(3366)) and (layer2_outputs(6737)));
    layer3_outputs(5311) <= not((layer2_outputs(2487)) and (layer2_outputs(2275)));
    layer3_outputs(5312) <= layer2_outputs(5624);
    layer3_outputs(5313) <= '1';
    layer3_outputs(5314) <= layer2_outputs(718);
    layer3_outputs(5315) <= not(layer2_outputs(3869));
    layer3_outputs(5316) <= not(layer2_outputs(3809));
    layer3_outputs(5317) <= (layer2_outputs(720)) and not (layer2_outputs(5985));
    layer3_outputs(5318) <= not((layer2_outputs(3005)) and (layer2_outputs(3823)));
    layer3_outputs(5319) <= (layer2_outputs(3988)) and not (layer2_outputs(7243));
    layer3_outputs(5320) <= layer2_outputs(2896);
    layer3_outputs(5321) <= layer2_outputs(7418);
    layer3_outputs(5322) <= not((layer2_outputs(4452)) xor (layer2_outputs(3253)));
    layer3_outputs(5323) <= (layer2_outputs(4601)) and (layer2_outputs(3910));
    layer3_outputs(5324) <= not(layer2_outputs(3116));
    layer3_outputs(5325) <= not(layer2_outputs(3832));
    layer3_outputs(5326) <= '1';
    layer3_outputs(5327) <= (layer2_outputs(6798)) or (layer2_outputs(5147));
    layer3_outputs(5328) <= not((layer2_outputs(2058)) or (layer2_outputs(5235)));
    layer3_outputs(5329) <= '0';
    layer3_outputs(5330) <= not(layer2_outputs(3982));
    layer3_outputs(5331) <= layer2_outputs(1662);
    layer3_outputs(5332) <= '0';
    layer3_outputs(5333) <= (layer2_outputs(2542)) and (layer2_outputs(6054));
    layer3_outputs(5334) <= '1';
    layer3_outputs(5335) <= layer2_outputs(6662);
    layer3_outputs(5336) <= (layer2_outputs(2778)) and (layer2_outputs(6639));
    layer3_outputs(5337) <= '1';
    layer3_outputs(5338) <= not(layer2_outputs(1617));
    layer3_outputs(5339) <= not((layer2_outputs(1570)) or (layer2_outputs(4585)));
    layer3_outputs(5340) <= layer2_outputs(1007);
    layer3_outputs(5341) <= layer2_outputs(5011);
    layer3_outputs(5342) <= (layer2_outputs(2284)) or (layer2_outputs(5933));
    layer3_outputs(5343) <= not(layer2_outputs(7310));
    layer3_outputs(5344) <= (layer2_outputs(3155)) or (layer2_outputs(5383));
    layer3_outputs(5345) <= not(layer2_outputs(4504)) or (layer2_outputs(679));
    layer3_outputs(5346) <= layer2_outputs(721);
    layer3_outputs(5347) <= not((layer2_outputs(1489)) and (layer2_outputs(101)));
    layer3_outputs(5348) <= '0';
    layer3_outputs(5349) <= not(layer2_outputs(854));
    layer3_outputs(5350) <= not(layer2_outputs(5707));
    layer3_outputs(5351) <= not(layer2_outputs(2040));
    layer3_outputs(5352) <= layer2_outputs(6561);
    layer3_outputs(5353) <= not((layer2_outputs(3055)) or (layer2_outputs(6653)));
    layer3_outputs(5354) <= not(layer2_outputs(4366)) or (layer2_outputs(113));
    layer3_outputs(5355) <= not(layer2_outputs(1022));
    layer3_outputs(5356) <= not(layer2_outputs(2362));
    layer3_outputs(5357) <= not(layer2_outputs(1386)) or (layer2_outputs(5521));
    layer3_outputs(5358) <= (layer2_outputs(2812)) and not (layer2_outputs(797));
    layer3_outputs(5359) <= '1';
    layer3_outputs(5360) <= not(layer2_outputs(965));
    layer3_outputs(5361) <= layer2_outputs(6459);
    layer3_outputs(5362) <= not(layer2_outputs(6116)) or (layer2_outputs(6591));
    layer3_outputs(5363) <= (layer2_outputs(5445)) and not (layer2_outputs(325));
    layer3_outputs(5364) <= not((layer2_outputs(4353)) or (layer2_outputs(7659)));
    layer3_outputs(5365) <= layer2_outputs(1244);
    layer3_outputs(5366) <= (layer2_outputs(1053)) or (layer2_outputs(6076));
    layer3_outputs(5367) <= (layer2_outputs(3897)) and not (layer2_outputs(2538));
    layer3_outputs(5368) <= not(layer2_outputs(4829));
    layer3_outputs(5369) <= not((layer2_outputs(7634)) xor (layer2_outputs(6595)));
    layer3_outputs(5370) <= not(layer2_outputs(6526));
    layer3_outputs(5371) <= not(layer2_outputs(1344));
    layer3_outputs(5372) <= (layer2_outputs(87)) and not (layer2_outputs(2356));
    layer3_outputs(5373) <= not(layer2_outputs(6513)) or (layer2_outputs(1217));
    layer3_outputs(5374) <= '1';
    layer3_outputs(5375) <= (layer2_outputs(6059)) or (layer2_outputs(86));
    layer3_outputs(5376) <= layer2_outputs(6936);
    layer3_outputs(5377) <= not(layer2_outputs(1607)) or (layer2_outputs(5600));
    layer3_outputs(5378) <= (layer2_outputs(7027)) and not (layer2_outputs(3848));
    layer3_outputs(5379) <= layer2_outputs(5424);
    layer3_outputs(5380) <= not(layer2_outputs(5134)) or (layer2_outputs(2136));
    layer3_outputs(5381) <= not(layer2_outputs(82)) or (layer2_outputs(5180));
    layer3_outputs(5382) <= not((layer2_outputs(6433)) and (layer2_outputs(2300)));
    layer3_outputs(5383) <= (layer2_outputs(3733)) or (layer2_outputs(7158));
    layer3_outputs(5384) <= not((layer2_outputs(7497)) or (layer2_outputs(3607)));
    layer3_outputs(5385) <= (layer2_outputs(2960)) or (layer2_outputs(5014));
    layer3_outputs(5386) <= not(layer2_outputs(2089));
    layer3_outputs(5387) <= layer2_outputs(3663);
    layer3_outputs(5388) <= not(layer2_outputs(2627)) or (layer2_outputs(413));
    layer3_outputs(5389) <= not((layer2_outputs(6586)) or (layer2_outputs(3298)));
    layer3_outputs(5390) <= not(layer2_outputs(7524)) or (layer2_outputs(6106));
    layer3_outputs(5391) <= (layer2_outputs(5707)) and (layer2_outputs(5306));
    layer3_outputs(5392) <= layer2_outputs(2052);
    layer3_outputs(5393) <= '1';
    layer3_outputs(5394) <= layer2_outputs(6214);
    layer3_outputs(5395) <= layer2_outputs(7330);
    layer3_outputs(5396) <= not((layer2_outputs(3885)) or (layer2_outputs(5645)));
    layer3_outputs(5397) <= (layer2_outputs(6818)) or (layer2_outputs(692));
    layer3_outputs(5398) <= not(layer2_outputs(862));
    layer3_outputs(5399) <= '0';
    layer3_outputs(5400) <= (layer2_outputs(610)) xor (layer2_outputs(1936));
    layer3_outputs(5401) <= (layer2_outputs(7019)) or (layer2_outputs(6895));
    layer3_outputs(5402) <= layer2_outputs(5747);
    layer3_outputs(5403) <= not(layer2_outputs(971)) or (layer2_outputs(4524));
    layer3_outputs(5404) <= (layer2_outputs(1878)) and not (layer2_outputs(784));
    layer3_outputs(5405) <= layer2_outputs(1378);
    layer3_outputs(5406) <= layer2_outputs(3271);
    layer3_outputs(5407) <= (layer2_outputs(5117)) or (layer2_outputs(100));
    layer3_outputs(5408) <= layer2_outputs(112);
    layer3_outputs(5409) <= not(layer2_outputs(5030));
    layer3_outputs(5410) <= (layer2_outputs(5718)) xor (layer2_outputs(2232));
    layer3_outputs(5411) <= layer2_outputs(3525);
    layer3_outputs(5412) <= not(layer2_outputs(5553)) or (layer2_outputs(3278));
    layer3_outputs(5413) <= not((layer2_outputs(83)) and (layer2_outputs(5969)));
    layer3_outputs(5414) <= layer2_outputs(5595);
    layer3_outputs(5415) <= '0';
    layer3_outputs(5416) <= not(layer2_outputs(1727));
    layer3_outputs(5417) <= not(layer2_outputs(572));
    layer3_outputs(5418) <= '1';
    layer3_outputs(5419) <= (layer2_outputs(885)) and not (layer2_outputs(7617));
    layer3_outputs(5420) <= not((layer2_outputs(1120)) and (layer2_outputs(7016)));
    layer3_outputs(5421) <= (layer2_outputs(4217)) xor (layer2_outputs(1098));
    layer3_outputs(5422) <= not(layer2_outputs(2806));
    layer3_outputs(5423) <= '1';
    layer3_outputs(5424) <= not(layer2_outputs(3585)) or (layer2_outputs(4599));
    layer3_outputs(5425) <= not(layer2_outputs(5598)) or (layer2_outputs(7099));
    layer3_outputs(5426) <= not(layer2_outputs(6070));
    layer3_outputs(5427) <= (layer2_outputs(3833)) and not (layer2_outputs(2769));
    layer3_outputs(5428) <= (layer2_outputs(245)) and (layer2_outputs(3518));
    layer3_outputs(5429) <= not(layer2_outputs(580)) or (layer2_outputs(5177));
    layer3_outputs(5430) <= (layer2_outputs(6380)) or (layer2_outputs(3881));
    layer3_outputs(5431) <= not((layer2_outputs(897)) and (layer2_outputs(741)));
    layer3_outputs(5432) <= not(layer2_outputs(1621));
    layer3_outputs(5433) <= (layer2_outputs(7156)) or (layer2_outputs(4524));
    layer3_outputs(5434) <= not(layer2_outputs(4363)) or (layer2_outputs(7115));
    layer3_outputs(5435) <= (layer2_outputs(5486)) and not (layer2_outputs(5156));
    layer3_outputs(5436) <= layer2_outputs(1913);
    layer3_outputs(5437) <= '0';
    layer3_outputs(5438) <= not(layer2_outputs(3303));
    layer3_outputs(5439) <= not(layer2_outputs(6952));
    layer3_outputs(5440) <= not(layer2_outputs(2364));
    layer3_outputs(5441) <= '0';
    layer3_outputs(5442) <= not((layer2_outputs(5414)) and (layer2_outputs(720)));
    layer3_outputs(5443) <= layer2_outputs(1767);
    layer3_outputs(5444) <= (layer2_outputs(6378)) xor (layer2_outputs(6347));
    layer3_outputs(5445) <= (layer2_outputs(2229)) and (layer2_outputs(1720));
    layer3_outputs(5446) <= '0';
    layer3_outputs(5447) <= (layer2_outputs(7320)) and (layer2_outputs(6323));
    layer3_outputs(5448) <= not(layer2_outputs(6250));
    layer3_outputs(5449) <= not(layer2_outputs(7322));
    layer3_outputs(5450) <= not(layer2_outputs(6438)) or (layer2_outputs(4719));
    layer3_outputs(5451) <= not(layer2_outputs(5282)) or (layer2_outputs(3581));
    layer3_outputs(5452) <= not((layer2_outputs(1209)) or (layer2_outputs(2078)));
    layer3_outputs(5453) <= layer2_outputs(4667);
    layer3_outputs(5454) <= (layer2_outputs(6493)) and not (layer2_outputs(2313));
    layer3_outputs(5455) <= (layer2_outputs(5536)) and not (layer2_outputs(4104));
    layer3_outputs(5456) <= not(layer2_outputs(5229)) or (layer2_outputs(4576));
    layer3_outputs(5457) <= not(layer2_outputs(6185));
    layer3_outputs(5458) <= layer2_outputs(2433);
    layer3_outputs(5459) <= not((layer2_outputs(1796)) and (layer2_outputs(5855)));
    layer3_outputs(5460) <= layer2_outputs(3706);
    layer3_outputs(5461) <= not((layer2_outputs(5088)) or (layer2_outputs(1578)));
    layer3_outputs(5462) <= '1';
    layer3_outputs(5463) <= (layer2_outputs(4291)) and not (layer2_outputs(4472));
    layer3_outputs(5464) <= not(layer2_outputs(1881));
    layer3_outputs(5465) <= not((layer2_outputs(6090)) xor (layer2_outputs(2550)));
    layer3_outputs(5466) <= not(layer2_outputs(3634));
    layer3_outputs(5467) <= (layer2_outputs(6140)) or (layer2_outputs(2551));
    layer3_outputs(5468) <= layer2_outputs(2538);
    layer3_outputs(5469) <= '1';
    layer3_outputs(5470) <= not(layer2_outputs(2774));
    layer3_outputs(5471) <= not(layer2_outputs(4670)) or (layer2_outputs(3531));
    layer3_outputs(5472) <= not(layer2_outputs(1839)) or (layer2_outputs(7141));
    layer3_outputs(5473) <= not((layer2_outputs(2690)) and (layer2_outputs(5009)));
    layer3_outputs(5474) <= (layer2_outputs(1491)) or (layer2_outputs(3338));
    layer3_outputs(5475) <= (layer2_outputs(4496)) and not (layer2_outputs(4730));
    layer3_outputs(5476) <= (layer2_outputs(7292)) and (layer2_outputs(3590));
    layer3_outputs(5477) <= not(layer2_outputs(2765));
    layer3_outputs(5478) <= layer2_outputs(2820);
    layer3_outputs(5479) <= (layer2_outputs(4365)) and (layer2_outputs(6394));
    layer3_outputs(5480) <= not(layer2_outputs(1597));
    layer3_outputs(5481) <= (layer2_outputs(3516)) and not (layer2_outputs(6548));
    layer3_outputs(5482) <= not(layer2_outputs(2406));
    layer3_outputs(5483) <= not(layer2_outputs(1942));
    layer3_outputs(5484) <= layer2_outputs(4326);
    layer3_outputs(5485) <= not(layer2_outputs(445)) or (layer2_outputs(3776));
    layer3_outputs(5486) <= '1';
    layer3_outputs(5487) <= not(layer2_outputs(4711));
    layer3_outputs(5488) <= '1';
    layer3_outputs(5489) <= layer2_outputs(1664);
    layer3_outputs(5490) <= not((layer2_outputs(6707)) xor (layer2_outputs(1830)));
    layer3_outputs(5491) <= (layer2_outputs(4748)) and not (layer2_outputs(4678));
    layer3_outputs(5492) <= not(layer2_outputs(3905));
    layer3_outputs(5493) <= (layer2_outputs(7560)) or (layer2_outputs(6991));
    layer3_outputs(5494) <= not((layer2_outputs(4060)) or (layer2_outputs(3507)));
    layer3_outputs(5495) <= (layer2_outputs(3435)) and (layer2_outputs(3595));
    layer3_outputs(5496) <= (layer2_outputs(3272)) or (layer2_outputs(3276));
    layer3_outputs(5497) <= (layer2_outputs(4729)) and (layer2_outputs(2007));
    layer3_outputs(5498) <= (layer2_outputs(5765)) or (layer2_outputs(1049));
    layer3_outputs(5499) <= not(layer2_outputs(237));
    layer3_outputs(5500) <= (layer2_outputs(7625)) and not (layer2_outputs(6050));
    layer3_outputs(5501) <= not(layer2_outputs(6091)) or (layer2_outputs(6428));
    layer3_outputs(5502) <= not(layer2_outputs(6194)) or (layer2_outputs(5292));
    layer3_outputs(5503) <= (layer2_outputs(2711)) and not (layer2_outputs(177));
    layer3_outputs(5504) <= not(layer2_outputs(5433)) or (layer2_outputs(1565));
    layer3_outputs(5505) <= not(layer2_outputs(2091));
    layer3_outputs(5506) <= not(layer2_outputs(2162)) or (layer2_outputs(6603));
    layer3_outputs(5507) <= layer2_outputs(556);
    layer3_outputs(5508) <= (layer2_outputs(5133)) and not (layer2_outputs(361));
    layer3_outputs(5509) <= layer2_outputs(6746);
    layer3_outputs(5510) <= not((layer2_outputs(4092)) or (layer2_outputs(5753)));
    layer3_outputs(5511) <= not((layer2_outputs(7044)) and (layer2_outputs(4353)));
    layer3_outputs(5512) <= not(layer2_outputs(3418));
    layer3_outputs(5513) <= layer2_outputs(7516);
    layer3_outputs(5514) <= '0';
    layer3_outputs(5515) <= not((layer2_outputs(6839)) or (layer2_outputs(2374)));
    layer3_outputs(5516) <= not((layer2_outputs(687)) xor (layer2_outputs(2379)));
    layer3_outputs(5517) <= (layer2_outputs(6821)) and (layer2_outputs(5409));
    layer3_outputs(5518) <= not((layer2_outputs(2723)) or (layer2_outputs(6697)));
    layer3_outputs(5519) <= layer2_outputs(534);
    layer3_outputs(5520) <= not((layer2_outputs(5000)) or (layer2_outputs(4731)));
    layer3_outputs(5521) <= '1';
    layer3_outputs(5522) <= '1';
    layer3_outputs(5523) <= not(layer2_outputs(6691)) or (layer2_outputs(3755));
    layer3_outputs(5524) <= not((layer2_outputs(3738)) or (layer2_outputs(4772)));
    layer3_outputs(5525) <= '1';
    layer3_outputs(5526) <= layer2_outputs(2556);
    layer3_outputs(5527) <= (layer2_outputs(2854)) xor (layer2_outputs(4797));
    layer3_outputs(5528) <= not(layer2_outputs(194));
    layer3_outputs(5529) <= (layer2_outputs(543)) or (layer2_outputs(367));
    layer3_outputs(5530) <= '1';
    layer3_outputs(5531) <= not(layer2_outputs(6036)) or (layer2_outputs(1929));
    layer3_outputs(5532) <= (layer2_outputs(2288)) and not (layer2_outputs(3855));
    layer3_outputs(5533) <= '0';
    layer3_outputs(5534) <= not(layer2_outputs(2716));
    layer3_outputs(5535) <= (layer2_outputs(6206)) or (layer2_outputs(1373));
    layer3_outputs(5536) <= not(layer2_outputs(5144));
    layer3_outputs(5537) <= layer2_outputs(115);
    layer3_outputs(5538) <= layer2_outputs(2718);
    layer3_outputs(5539) <= not((layer2_outputs(6169)) and (layer2_outputs(7275)));
    layer3_outputs(5540) <= not((layer2_outputs(6198)) or (layer2_outputs(5126)));
    layer3_outputs(5541) <= not((layer2_outputs(4554)) or (layer2_outputs(3621)));
    layer3_outputs(5542) <= not(layer2_outputs(6674)) or (layer2_outputs(394));
    layer3_outputs(5543) <= (layer2_outputs(4661)) and (layer2_outputs(3707));
    layer3_outputs(5544) <= layer2_outputs(3816);
    layer3_outputs(5545) <= not(layer2_outputs(6344));
    layer3_outputs(5546) <= layer2_outputs(3916);
    layer3_outputs(5547) <= layer2_outputs(4170);
    layer3_outputs(5548) <= not(layer2_outputs(295));
    layer3_outputs(5549) <= '1';
    layer3_outputs(5550) <= not(layer2_outputs(6650));
    layer3_outputs(5551) <= not((layer2_outputs(4440)) xor (layer2_outputs(4448)));
    layer3_outputs(5552) <= not((layer2_outputs(4384)) or (layer2_outputs(5211)));
    layer3_outputs(5553) <= (layer2_outputs(2508)) or (layer2_outputs(4209));
    layer3_outputs(5554) <= (layer2_outputs(7147)) and not (layer2_outputs(1195));
    layer3_outputs(5555) <= '0';
    layer3_outputs(5556) <= (layer2_outputs(5309)) and (layer2_outputs(2170));
    layer3_outputs(5557) <= not((layer2_outputs(7635)) and (layer2_outputs(6690)));
    layer3_outputs(5558) <= not(layer2_outputs(7450));
    layer3_outputs(5559) <= not(layer2_outputs(7167)) or (layer2_outputs(6745));
    layer3_outputs(5560) <= not(layer2_outputs(5061));
    layer3_outputs(5561) <= not(layer2_outputs(6233));
    layer3_outputs(5562) <= not((layer2_outputs(5813)) and (layer2_outputs(6852)));
    layer3_outputs(5563) <= (layer2_outputs(5639)) xor (layer2_outputs(3132));
    layer3_outputs(5564) <= not(layer2_outputs(4385)) or (layer2_outputs(5056));
    layer3_outputs(5565) <= (layer2_outputs(1455)) or (layer2_outputs(3633));
    layer3_outputs(5566) <= not(layer2_outputs(150));
    layer3_outputs(5567) <= '0';
    layer3_outputs(5568) <= (layer2_outputs(3238)) and not (layer2_outputs(6918));
    layer3_outputs(5569) <= not((layer2_outputs(7139)) or (layer2_outputs(5122)));
    layer3_outputs(5570) <= layer2_outputs(5978);
    layer3_outputs(5571) <= not((layer2_outputs(5102)) and (layer2_outputs(2096)));
    layer3_outputs(5572) <= not((layer2_outputs(7279)) and (layer2_outputs(4805)));
    layer3_outputs(5573) <= not(layer2_outputs(1841)) or (layer2_outputs(3184));
    layer3_outputs(5574) <= not(layer2_outputs(1819));
    layer3_outputs(5575) <= (layer2_outputs(6246)) and (layer2_outputs(5834));
    layer3_outputs(5576) <= (layer2_outputs(6479)) and not (layer2_outputs(3272));
    layer3_outputs(5577) <= not(layer2_outputs(99));
    layer3_outputs(5578) <= '1';
    layer3_outputs(5579) <= not(layer2_outputs(5259));
    layer3_outputs(5580) <= (layer2_outputs(5906)) or (layer2_outputs(5834));
    layer3_outputs(5581) <= (layer2_outputs(1717)) and not (layer2_outputs(4784));
    layer3_outputs(5582) <= not((layer2_outputs(1235)) or (layer2_outputs(519)));
    layer3_outputs(5583) <= (layer2_outputs(3445)) xor (layer2_outputs(5023));
    layer3_outputs(5584) <= '1';
    layer3_outputs(5585) <= not(layer2_outputs(3540));
    layer3_outputs(5586) <= not(layer2_outputs(3437)) or (layer2_outputs(1436));
    layer3_outputs(5587) <= not((layer2_outputs(4287)) or (layer2_outputs(607)));
    layer3_outputs(5588) <= not(layer2_outputs(2691)) or (layer2_outputs(4638));
    layer3_outputs(5589) <= '1';
    layer3_outputs(5590) <= not((layer2_outputs(4507)) and (layer2_outputs(325)));
    layer3_outputs(5591) <= (layer2_outputs(3322)) and not (layer2_outputs(4706));
    layer3_outputs(5592) <= not(layer2_outputs(5209)) or (layer2_outputs(6583));
    layer3_outputs(5593) <= (layer2_outputs(4587)) and (layer2_outputs(1617));
    layer3_outputs(5594) <= not((layer2_outputs(6068)) or (layer2_outputs(1835)));
    layer3_outputs(5595) <= not((layer2_outputs(2114)) and (layer2_outputs(1307)));
    layer3_outputs(5596) <= (layer2_outputs(3171)) and not (layer2_outputs(5256));
    layer3_outputs(5597) <= layer2_outputs(6892);
    layer3_outputs(5598) <= not(layer2_outputs(4912));
    layer3_outputs(5599) <= '0';
    layer3_outputs(5600) <= not((layer2_outputs(299)) and (layer2_outputs(1493)));
    layer3_outputs(5601) <= '1';
    layer3_outputs(5602) <= '0';
    layer3_outputs(5603) <= not(layer2_outputs(429)) or (layer2_outputs(1920));
    layer3_outputs(5604) <= '0';
    layer3_outputs(5605) <= not((layer2_outputs(4815)) and (layer2_outputs(2362)));
    layer3_outputs(5606) <= '1';
    layer3_outputs(5607) <= (layer2_outputs(1109)) or (layer2_outputs(2684));
    layer3_outputs(5608) <= '0';
    layer3_outputs(5609) <= layer2_outputs(621);
    layer3_outputs(5610) <= layer2_outputs(2787);
    layer3_outputs(5611) <= '1';
    layer3_outputs(5612) <= layer2_outputs(3942);
    layer3_outputs(5613) <= layer2_outputs(4410);
    layer3_outputs(5614) <= not((layer2_outputs(2510)) and (layer2_outputs(58)));
    layer3_outputs(5615) <= not(layer2_outputs(4814)) or (layer2_outputs(4996));
    layer3_outputs(5616) <= not(layer2_outputs(3503)) or (layer2_outputs(3668));
    layer3_outputs(5617) <= layer2_outputs(2243);
    layer3_outputs(5618) <= not(layer2_outputs(7119)) or (layer2_outputs(7439));
    layer3_outputs(5619) <= layer2_outputs(558);
    layer3_outputs(5620) <= not(layer2_outputs(3763)) or (layer2_outputs(5723));
    layer3_outputs(5621) <= not((layer2_outputs(4844)) or (layer2_outputs(147)));
    layer3_outputs(5622) <= not(layer2_outputs(70));
    layer3_outputs(5623) <= not(layer2_outputs(3107));
    layer3_outputs(5624) <= layer2_outputs(973);
    layer3_outputs(5625) <= (layer2_outputs(2987)) xor (layer2_outputs(3837));
    layer3_outputs(5626) <= not((layer2_outputs(876)) or (layer2_outputs(296)));
    layer3_outputs(5627) <= '0';
    layer3_outputs(5628) <= layer2_outputs(6231);
    layer3_outputs(5629) <= layer2_outputs(1422);
    layer3_outputs(5630) <= layer2_outputs(1560);
    layer3_outputs(5631) <= layer2_outputs(3783);
    layer3_outputs(5632) <= (layer2_outputs(5283)) or (layer2_outputs(3961));
    layer3_outputs(5633) <= (layer2_outputs(2029)) or (layer2_outputs(4123));
    layer3_outputs(5634) <= '1';
    layer3_outputs(5635) <= layer2_outputs(5742);
    layer3_outputs(5636) <= (layer2_outputs(4015)) or (layer2_outputs(6032));
    layer3_outputs(5637) <= (layer2_outputs(1370)) or (layer2_outputs(1739));
    layer3_outputs(5638) <= not(layer2_outputs(7511)) or (layer2_outputs(2361));
    layer3_outputs(5639) <= not(layer2_outputs(3735));
    layer3_outputs(5640) <= (layer2_outputs(814)) and (layer2_outputs(7302));
    layer3_outputs(5641) <= layer2_outputs(5843);
    layer3_outputs(5642) <= (layer2_outputs(595)) xor (layer2_outputs(6148));
    layer3_outputs(5643) <= layer2_outputs(3132);
    layer3_outputs(5644) <= (layer2_outputs(7229)) or (layer2_outputs(3826));
    layer3_outputs(5645) <= not(layer2_outputs(2474)) or (layer2_outputs(5807));
    layer3_outputs(5646) <= (layer2_outputs(2581)) or (layer2_outputs(6041));
    layer3_outputs(5647) <= layer2_outputs(3512);
    layer3_outputs(5648) <= not(layer2_outputs(6421));
    layer3_outputs(5649) <= (layer2_outputs(1331)) and not (layer2_outputs(5202));
    layer3_outputs(5650) <= (layer2_outputs(6181)) and not (layer2_outputs(5004));
    layer3_outputs(5651) <= not(layer2_outputs(760)) or (layer2_outputs(5895));
    layer3_outputs(5652) <= (layer2_outputs(1781)) and (layer2_outputs(4372));
    layer3_outputs(5653) <= (layer2_outputs(6890)) and not (layer2_outputs(6287));
    layer3_outputs(5654) <= (layer2_outputs(6101)) and (layer2_outputs(3992));
    layer3_outputs(5655) <= layer2_outputs(3323);
    layer3_outputs(5656) <= (layer2_outputs(5407)) or (layer2_outputs(4466));
    layer3_outputs(5657) <= (layer2_outputs(156)) and not (layer2_outputs(5853));
    layer3_outputs(5658) <= layer2_outputs(4281);
    layer3_outputs(5659) <= layer2_outputs(6540);
    layer3_outputs(5660) <= layer2_outputs(6256);
    layer3_outputs(5661) <= '0';
    layer3_outputs(5662) <= '0';
    layer3_outputs(5663) <= not((layer2_outputs(2520)) and (layer2_outputs(5926)));
    layer3_outputs(5664) <= layer2_outputs(7601);
    layer3_outputs(5665) <= '0';
    layer3_outputs(5666) <= (layer2_outputs(3903)) and (layer2_outputs(5442));
    layer3_outputs(5667) <= (layer2_outputs(5983)) xor (layer2_outputs(2575));
    layer3_outputs(5668) <= layer2_outputs(417);
    layer3_outputs(5669) <= not((layer2_outputs(4070)) or (layer2_outputs(5653)));
    layer3_outputs(5670) <= layer2_outputs(5869);
    layer3_outputs(5671) <= layer2_outputs(842);
    layer3_outputs(5672) <= not(layer2_outputs(3691)) or (layer2_outputs(5047));
    layer3_outputs(5673) <= (layer2_outputs(1412)) and (layer2_outputs(3995));
    layer3_outputs(5674) <= '0';
    layer3_outputs(5675) <= not(layer2_outputs(7494));
    layer3_outputs(5676) <= not((layer2_outputs(4317)) or (layer2_outputs(2008)));
    layer3_outputs(5677) <= '0';
    layer3_outputs(5678) <= layer2_outputs(844);
    layer3_outputs(5679) <= layer2_outputs(5748);
    layer3_outputs(5680) <= not(layer2_outputs(5270));
    layer3_outputs(5681) <= '0';
    layer3_outputs(5682) <= '1';
    layer3_outputs(5683) <= not((layer2_outputs(6681)) or (layer2_outputs(5867)));
    layer3_outputs(5684) <= not(layer2_outputs(3474)) or (layer2_outputs(3959));
    layer3_outputs(5685) <= not(layer2_outputs(6476)) or (layer2_outputs(2336));
    layer3_outputs(5686) <= '1';
    layer3_outputs(5687) <= not((layer2_outputs(3561)) and (layer2_outputs(1269)));
    layer3_outputs(5688) <= (layer2_outputs(1842)) and not (layer2_outputs(1614));
    layer3_outputs(5689) <= layer2_outputs(5195);
    layer3_outputs(5690) <= layer2_outputs(3710);
    layer3_outputs(5691) <= not(layer2_outputs(3359)) or (layer2_outputs(4502));
    layer3_outputs(5692) <= (layer2_outputs(6121)) and not (layer2_outputs(7488));
    layer3_outputs(5693) <= (layer2_outputs(3203)) and not (layer2_outputs(3831));
    layer3_outputs(5694) <= not(layer2_outputs(6607));
    layer3_outputs(5695) <= not(layer2_outputs(930));
    layer3_outputs(5696) <= layer2_outputs(6423);
    layer3_outputs(5697) <= (layer2_outputs(4030)) and (layer2_outputs(7266));
    layer3_outputs(5698) <= not(layer2_outputs(3227));
    layer3_outputs(5699) <= not(layer2_outputs(1134)) or (layer2_outputs(926));
    layer3_outputs(5700) <= not(layer2_outputs(5300));
    layer3_outputs(5701) <= layer2_outputs(7209);
    layer3_outputs(5702) <= not(layer2_outputs(5478)) or (layer2_outputs(7677));
    layer3_outputs(5703) <= (layer2_outputs(4089)) and (layer2_outputs(5329));
    layer3_outputs(5704) <= not(layer2_outputs(4010));
    layer3_outputs(5705) <= (layer2_outputs(3407)) and not (layer2_outputs(2844));
    layer3_outputs(5706) <= not((layer2_outputs(3078)) or (layer2_outputs(1253)));
    layer3_outputs(5707) <= (layer2_outputs(567)) and (layer2_outputs(6167));
    layer3_outputs(5708) <= (layer2_outputs(6219)) and not (layer2_outputs(6178));
    layer3_outputs(5709) <= not(layer2_outputs(6660)) or (layer2_outputs(3310));
    layer3_outputs(5710) <= not(layer2_outputs(5330)) or (layer2_outputs(3086));
    layer3_outputs(5711) <= not(layer2_outputs(2675));
    layer3_outputs(5712) <= not((layer2_outputs(5031)) and (layer2_outputs(5805)));
    layer3_outputs(5713) <= layer2_outputs(5105);
    layer3_outputs(5714) <= (layer2_outputs(15)) and not (layer2_outputs(4425));
    layer3_outputs(5715) <= (layer2_outputs(1591)) and (layer2_outputs(36));
    layer3_outputs(5716) <= (layer2_outputs(4749)) xor (layer2_outputs(6778));
    layer3_outputs(5717) <= not(layer2_outputs(1541));
    layer3_outputs(5718) <= not(layer2_outputs(1377));
    layer3_outputs(5719) <= layer2_outputs(6912);
    layer3_outputs(5720) <= '1';
    layer3_outputs(5721) <= layer2_outputs(6337);
    layer3_outputs(5722) <= not(layer2_outputs(6763));
    layer3_outputs(5723) <= not(layer2_outputs(4922));
    layer3_outputs(5724) <= not(layer2_outputs(7331)) or (layer2_outputs(2225));
    layer3_outputs(5725) <= layer2_outputs(447);
    layer3_outputs(5726) <= not((layer2_outputs(3565)) xor (layer2_outputs(3957)));
    layer3_outputs(5727) <= not(layer2_outputs(618)) or (layer2_outputs(7582));
    layer3_outputs(5728) <= (layer2_outputs(4545)) and not (layer2_outputs(562));
    layer3_outputs(5729) <= not(layer2_outputs(881)) or (layer2_outputs(1141));
    layer3_outputs(5730) <= not(layer2_outputs(7536));
    layer3_outputs(5731) <= (layer2_outputs(582)) and not (layer2_outputs(3030));
    layer3_outputs(5732) <= layer2_outputs(6961);
    layer3_outputs(5733) <= not((layer2_outputs(987)) or (layer2_outputs(4368)));
    layer3_outputs(5734) <= not(layer2_outputs(3394));
    layer3_outputs(5735) <= layer2_outputs(3386);
    layer3_outputs(5736) <= (layer2_outputs(2545)) and not (layer2_outputs(3842));
    layer3_outputs(5737) <= '0';
    layer3_outputs(5738) <= '0';
    layer3_outputs(5739) <= (layer2_outputs(5412)) and not (layer2_outputs(2094));
    layer3_outputs(5740) <= not((layer2_outputs(5960)) or (layer2_outputs(4424)));
    layer3_outputs(5741) <= layer2_outputs(6826);
    layer3_outputs(5742) <= (layer2_outputs(3719)) and not (layer2_outputs(136));
    layer3_outputs(5743) <= (layer2_outputs(1199)) and not (layer2_outputs(6215));
    layer3_outputs(5744) <= not(layer2_outputs(6982)) or (layer2_outputs(7570));
    layer3_outputs(5745) <= not(layer2_outputs(170));
    layer3_outputs(5746) <= layer2_outputs(275);
    layer3_outputs(5747) <= (layer2_outputs(2898)) and not (layer2_outputs(3080));
    layer3_outputs(5748) <= not(layer2_outputs(4954));
    layer3_outputs(5749) <= '1';
    layer3_outputs(5750) <= not((layer2_outputs(628)) and (layer2_outputs(7054)));
    layer3_outputs(5751) <= layer2_outputs(504);
    layer3_outputs(5752) <= not(layer2_outputs(5787));
    layer3_outputs(5753) <= not(layer2_outputs(6929)) or (layer2_outputs(3723));
    layer3_outputs(5754) <= (layer2_outputs(7542)) and not (layer2_outputs(1830));
    layer3_outputs(5755) <= (layer2_outputs(2733)) or (layer2_outputs(6620));
    layer3_outputs(5756) <= (layer2_outputs(5561)) xor (layer2_outputs(1733));
    layer3_outputs(5757) <= not((layer2_outputs(3358)) or (layer2_outputs(1616)));
    layer3_outputs(5758) <= not((layer2_outputs(6505)) or (layer2_outputs(2471)));
    layer3_outputs(5759) <= '0';
    layer3_outputs(5760) <= (layer2_outputs(4422)) and not (layer2_outputs(3350));
    layer3_outputs(5761) <= '1';
    layer3_outputs(5762) <= not(layer2_outputs(6875));
    layer3_outputs(5763) <= not(layer2_outputs(993));
    layer3_outputs(5764) <= not(layer2_outputs(4759)) or (layer2_outputs(6895));
    layer3_outputs(5765) <= not(layer2_outputs(3245));
    layer3_outputs(5766) <= (layer2_outputs(3254)) or (layer2_outputs(3432));
    layer3_outputs(5767) <= layer2_outputs(6840);
    layer3_outputs(5768) <= (layer2_outputs(2546)) or (layer2_outputs(2201));
    layer3_outputs(5769) <= not(layer2_outputs(5108));
    layer3_outputs(5770) <= (layer2_outputs(4234)) and (layer2_outputs(1423));
    layer3_outputs(5771) <= (layer2_outputs(15)) and not (layer2_outputs(1507));
    layer3_outputs(5772) <= not(layer2_outputs(1102)) or (layer2_outputs(6332));
    layer3_outputs(5773) <= (layer2_outputs(3144)) and (layer2_outputs(4572));
    layer3_outputs(5774) <= not(layer2_outputs(4565));
    layer3_outputs(5775) <= (layer2_outputs(3570)) xor (layer2_outputs(4506));
    layer3_outputs(5776) <= not(layer2_outputs(2616));
    layer3_outputs(5777) <= not((layer2_outputs(4534)) or (layer2_outputs(2145)));
    layer3_outputs(5778) <= (layer2_outputs(7283)) and (layer2_outputs(3601));
    layer3_outputs(5779) <= not(layer2_outputs(7597));
    layer3_outputs(5780) <= (layer2_outputs(4052)) and not (layer2_outputs(2532));
    layer3_outputs(5781) <= layer2_outputs(1218);
    layer3_outputs(5782) <= not((layer2_outputs(4696)) and (layer2_outputs(4082)));
    layer3_outputs(5783) <= layer2_outputs(4938);
    layer3_outputs(5784) <= '1';
    layer3_outputs(5785) <= layer2_outputs(3574);
    layer3_outputs(5786) <= not((layer2_outputs(1223)) or (layer2_outputs(25)));
    layer3_outputs(5787) <= not((layer2_outputs(6909)) and (layer2_outputs(2523)));
    layer3_outputs(5788) <= layer2_outputs(7643);
    layer3_outputs(5789) <= not(layer2_outputs(4630));
    layer3_outputs(5790) <= not(layer2_outputs(5342));
    layer3_outputs(5791) <= (layer2_outputs(479)) and not (layer2_outputs(3041));
    layer3_outputs(5792) <= '1';
    layer3_outputs(5793) <= (layer2_outputs(3647)) or (layer2_outputs(371));
    layer3_outputs(5794) <= (layer2_outputs(5704)) and not (layer2_outputs(7667));
    layer3_outputs(5795) <= (layer2_outputs(1368)) and not (layer2_outputs(4407));
    layer3_outputs(5796) <= '0';
    layer3_outputs(5797) <= layer2_outputs(1077);
    layer3_outputs(5798) <= not(layer2_outputs(6685));
    layer3_outputs(5799) <= (layer2_outputs(2525)) or (layer2_outputs(693));
    layer3_outputs(5800) <= (layer2_outputs(35)) xor (layer2_outputs(5409));
    layer3_outputs(5801) <= layer2_outputs(4624);
    layer3_outputs(5802) <= layer2_outputs(4085);
    layer3_outputs(5803) <= layer2_outputs(5311);
    layer3_outputs(5804) <= not(layer2_outputs(7676));
    layer3_outputs(5805) <= not(layer2_outputs(3009)) or (layer2_outputs(670));
    layer3_outputs(5806) <= (layer2_outputs(3637)) xor (layer2_outputs(2544));
    layer3_outputs(5807) <= layer2_outputs(7479);
    layer3_outputs(5808) <= not((layer2_outputs(5699)) or (layer2_outputs(6386)));
    layer3_outputs(5809) <= not((layer2_outputs(6391)) or (layer2_outputs(4556)));
    layer3_outputs(5810) <= layer2_outputs(6456);
    layer3_outputs(5811) <= not(layer2_outputs(7463));
    layer3_outputs(5812) <= (layer2_outputs(4445)) and not (layer2_outputs(2681));
    layer3_outputs(5813) <= layer2_outputs(6566);
    layer3_outputs(5814) <= not(layer2_outputs(1533));
    layer3_outputs(5815) <= layer2_outputs(145);
    layer3_outputs(5816) <= (layer2_outputs(6351)) or (layer2_outputs(6547));
    layer3_outputs(5817) <= not((layer2_outputs(7311)) and (layer2_outputs(5456)));
    layer3_outputs(5818) <= not(layer2_outputs(1500)) or (layer2_outputs(4296));
    layer3_outputs(5819) <= layer2_outputs(4902);
    layer3_outputs(5820) <= not(layer2_outputs(6537)) or (layer2_outputs(6994));
    layer3_outputs(5821) <= layer2_outputs(3760);
    layer3_outputs(5822) <= not(layer2_outputs(2398)) or (layer2_outputs(1064));
    layer3_outputs(5823) <= not(layer2_outputs(1725)) or (layer2_outputs(2060));
    layer3_outputs(5824) <= not((layer2_outputs(7135)) and (layer2_outputs(3279)));
    layer3_outputs(5825) <= '0';
    layer3_outputs(5826) <= (layer2_outputs(5790)) and (layer2_outputs(825));
    layer3_outputs(5827) <= not(layer2_outputs(5468));
    layer3_outputs(5828) <= layer2_outputs(6399);
    layer3_outputs(5829) <= layer2_outputs(2337);
    layer3_outputs(5830) <= layer2_outputs(6019);
    layer3_outputs(5831) <= (layer2_outputs(2355)) and not (layer2_outputs(1932));
    layer3_outputs(5832) <= not(layer2_outputs(6873));
    layer3_outputs(5833) <= layer2_outputs(2809);
    layer3_outputs(5834) <= (layer2_outputs(1233)) and not (layer2_outputs(499));
    layer3_outputs(5835) <= not((layer2_outputs(2886)) or (layer2_outputs(2176)));
    layer3_outputs(5836) <= layer2_outputs(956);
    layer3_outputs(5837) <= (layer2_outputs(176)) and not (layer2_outputs(1395));
    layer3_outputs(5838) <= not(layer2_outputs(2557)) or (layer2_outputs(7385));
    layer3_outputs(5839) <= '0';
    layer3_outputs(5840) <= (layer2_outputs(858)) and (layer2_outputs(4868));
    layer3_outputs(5841) <= not(layer2_outputs(424));
    layer3_outputs(5842) <= not(layer2_outputs(1310));
    layer3_outputs(5843) <= not(layer2_outputs(1570));
    layer3_outputs(5844) <= (layer2_outputs(6961)) and not (layer2_outputs(2050));
    layer3_outputs(5845) <= (layer2_outputs(460)) or (layer2_outputs(5676));
    layer3_outputs(5846) <= (layer2_outputs(233)) and not (layer2_outputs(6108));
    layer3_outputs(5847) <= '1';
    layer3_outputs(5848) <= (layer2_outputs(6541)) and (layer2_outputs(4664));
    layer3_outputs(5849) <= layer2_outputs(119);
    layer3_outputs(5850) <= not((layer2_outputs(962)) or (layer2_outputs(2558)));
    layer3_outputs(5851) <= (layer2_outputs(5693)) and (layer2_outputs(4817));
    layer3_outputs(5852) <= (layer2_outputs(7421)) xor (layer2_outputs(6514));
    layer3_outputs(5853) <= not(layer2_outputs(5477));
    layer3_outputs(5854) <= not(layer2_outputs(7348));
    layer3_outputs(5855) <= '1';
    layer3_outputs(5856) <= (layer2_outputs(510)) or (layer2_outputs(5989));
    layer3_outputs(5857) <= (layer2_outputs(3627)) and (layer2_outputs(7638));
    layer3_outputs(5858) <= not(layer2_outputs(2487)) or (layer2_outputs(4810));
    layer3_outputs(5859) <= not((layer2_outputs(1356)) and (layer2_outputs(6355)));
    layer3_outputs(5860) <= (layer2_outputs(4642)) and not (layer2_outputs(7512));
    layer3_outputs(5861) <= (layer2_outputs(3195)) and not (layer2_outputs(1520));
    layer3_outputs(5862) <= not((layer2_outputs(7431)) and (layer2_outputs(1144)));
    layer3_outputs(5863) <= (layer2_outputs(5812)) and (layer2_outputs(2683));
    layer3_outputs(5864) <= layer2_outputs(23);
    layer3_outputs(5865) <= not((layer2_outputs(6826)) xor (layer2_outputs(4066)));
    layer3_outputs(5866) <= '0';
    layer3_outputs(5867) <= not((layer2_outputs(6678)) or (layer2_outputs(3976)));
    layer3_outputs(5868) <= layer2_outputs(241);
    layer3_outputs(5869) <= '1';
    layer3_outputs(5870) <= (layer2_outputs(5730)) and not (layer2_outputs(4772));
    layer3_outputs(5871) <= not(layer2_outputs(1160));
    layer3_outputs(5872) <= not((layer2_outputs(5153)) and (layer2_outputs(3081)));
    layer3_outputs(5873) <= '0';
    layer3_outputs(5874) <= not((layer2_outputs(6338)) xor (layer2_outputs(6313)));
    layer3_outputs(5875) <= not((layer2_outputs(5336)) or (layer2_outputs(6912)));
    layer3_outputs(5876) <= not(layer2_outputs(3887));
    layer3_outputs(5877) <= (layer2_outputs(259)) or (layer2_outputs(5847));
    layer3_outputs(5878) <= (layer2_outputs(1144)) xor (layer2_outputs(693));
    layer3_outputs(5879) <= not(layer2_outputs(6673));
    layer3_outputs(5880) <= (layer2_outputs(3136)) and not (layer2_outputs(5127));
    layer3_outputs(5881) <= (layer2_outputs(6162)) and (layer2_outputs(4178));
    layer3_outputs(5882) <= not(layer2_outputs(882));
    layer3_outputs(5883) <= (layer2_outputs(1543)) and not (layer2_outputs(3051));
    layer3_outputs(5884) <= layer2_outputs(4223);
    layer3_outputs(5885) <= (layer2_outputs(5012)) xor (layer2_outputs(4599));
    layer3_outputs(5886) <= layer2_outputs(6497);
    layer3_outputs(5887) <= (layer2_outputs(5124)) and (layer2_outputs(7282));
    layer3_outputs(5888) <= not(layer2_outputs(3091)) or (layer2_outputs(7472));
    layer3_outputs(5889) <= not(layer2_outputs(6360));
    layer3_outputs(5890) <= not((layer2_outputs(3587)) and (layer2_outputs(3941)));
    layer3_outputs(5891) <= '0';
    layer3_outputs(5892) <= layer2_outputs(6361);
    layer3_outputs(5893) <= (layer2_outputs(1595)) or (layer2_outputs(5054));
    layer3_outputs(5894) <= not(layer2_outputs(5225));
    layer3_outputs(5895) <= not(layer2_outputs(1482));
    layer3_outputs(5896) <= not(layer2_outputs(1945));
    layer3_outputs(5897) <= (layer2_outputs(2801)) or (layer2_outputs(5454));
    layer3_outputs(5898) <= not((layer2_outputs(6228)) or (layer2_outputs(7010)));
    layer3_outputs(5899) <= (layer2_outputs(1531)) and (layer2_outputs(4110));
    layer3_outputs(5900) <= not((layer2_outputs(5044)) or (layer2_outputs(5977)));
    layer3_outputs(5901) <= (layer2_outputs(5293)) or (layer2_outputs(1749));
    layer3_outputs(5902) <= not((layer2_outputs(6806)) or (layer2_outputs(6241)));
    layer3_outputs(5903) <= layer2_outputs(5679);
    layer3_outputs(5904) <= not((layer2_outputs(721)) and (layer2_outputs(5553)));
    layer3_outputs(5905) <= not(layer2_outputs(907)) or (layer2_outputs(7205));
    layer3_outputs(5906) <= not(layer2_outputs(6833)) or (layer2_outputs(5928));
    layer3_outputs(5907) <= (layer2_outputs(3163)) or (layer2_outputs(5164));
    layer3_outputs(5908) <= not((layer2_outputs(3996)) xor (layer2_outputs(7411)));
    layer3_outputs(5909) <= layer2_outputs(467);
    layer3_outputs(5910) <= '1';
    layer3_outputs(5911) <= not((layer2_outputs(6130)) or (layer2_outputs(3934)));
    layer3_outputs(5912) <= not(layer2_outputs(3628));
    layer3_outputs(5913) <= (layer2_outputs(1147)) and (layer2_outputs(4142));
    layer3_outputs(5914) <= not(layer2_outputs(149));
    layer3_outputs(5915) <= layer2_outputs(220);
    layer3_outputs(5916) <= not(layer2_outputs(49));
    layer3_outputs(5917) <= layer2_outputs(1621);
    layer3_outputs(5918) <= (layer2_outputs(4997)) or (layer2_outputs(5720));
    layer3_outputs(5919) <= not(layer2_outputs(4716)) or (layer2_outputs(4032));
    layer3_outputs(5920) <= not(layer2_outputs(3936)) or (layer2_outputs(3631));
    layer3_outputs(5921) <= (layer2_outputs(5339)) and not (layer2_outputs(2203));
    layer3_outputs(5922) <= (layer2_outputs(4000)) and not (layer2_outputs(2979));
    layer3_outputs(5923) <= (layer2_outputs(1466)) and not (layer2_outputs(1008));
    layer3_outputs(5924) <= layer2_outputs(103);
    layer3_outputs(5925) <= (layer2_outputs(1895)) and not (layer2_outputs(6732));
    layer3_outputs(5926) <= not(layer2_outputs(4131));
    layer3_outputs(5927) <= layer2_outputs(5877);
    layer3_outputs(5928) <= (layer2_outputs(4392)) xor (layer2_outputs(3921));
    layer3_outputs(5929) <= layer2_outputs(3567);
    layer3_outputs(5930) <= not(layer2_outputs(4477));
    layer3_outputs(5931) <= (layer2_outputs(3233)) and (layer2_outputs(4463));
    layer3_outputs(5932) <= layer2_outputs(155);
    layer3_outputs(5933) <= (layer2_outputs(6618)) and (layer2_outputs(5267));
    layer3_outputs(5934) <= not(layer2_outputs(2005));
    layer3_outputs(5935) <= not(layer2_outputs(6947)) or (layer2_outputs(6936));
    layer3_outputs(5936) <= not(layer2_outputs(748)) or (layer2_outputs(1029));
    layer3_outputs(5937) <= layer2_outputs(4289);
    layer3_outputs(5938) <= layer2_outputs(5991);
    layer3_outputs(5939) <= (layer2_outputs(5645)) or (layer2_outputs(133));
    layer3_outputs(5940) <= not(layer2_outputs(431));
    layer3_outputs(5941) <= '1';
    layer3_outputs(5942) <= not(layer2_outputs(1467));
    layer3_outputs(5943) <= '1';
    layer3_outputs(5944) <= (layer2_outputs(7458)) or (layer2_outputs(4343));
    layer3_outputs(5945) <= not(layer2_outputs(6500));
    layer3_outputs(5946) <= not((layer2_outputs(866)) xor (layer2_outputs(507)));
    layer3_outputs(5947) <= (layer2_outputs(4038)) and (layer2_outputs(5392));
    layer3_outputs(5948) <= layer2_outputs(418);
    layer3_outputs(5949) <= '1';
    layer3_outputs(5950) <= not((layer2_outputs(5726)) and (layer2_outputs(1883)));
    layer3_outputs(5951) <= not(layer2_outputs(333)) or (layer2_outputs(3415));
    layer3_outputs(5952) <= not((layer2_outputs(2015)) and (layer2_outputs(6983)));
    layer3_outputs(5953) <= '1';
    layer3_outputs(5954) <= not(layer2_outputs(3456));
    layer3_outputs(5955) <= layer2_outputs(3156);
    layer3_outputs(5956) <= layer2_outputs(1755);
    layer3_outputs(5957) <= not(layer2_outputs(5151)) or (layer2_outputs(5328));
    layer3_outputs(5958) <= not(layer2_outputs(1417)) or (layer2_outputs(1099));
    layer3_outputs(5959) <= layer2_outputs(3205);
    layer3_outputs(5960) <= (layer2_outputs(2066)) or (layer2_outputs(7654));
    layer3_outputs(5961) <= (layer2_outputs(1204)) and (layer2_outputs(6992));
    layer3_outputs(5962) <= not(layer2_outputs(4770));
    layer3_outputs(5963) <= not(layer2_outputs(1660)) or (layer2_outputs(6858));
    layer3_outputs(5964) <= layer2_outputs(1933);
    layer3_outputs(5965) <= not(layer2_outputs(1138));
    layer3_outputs(5966) <= (layer2_outputs(6379)) and not (layer2_outputs(2218));
    layer3_outputs(5967) <= not((layer2_outputs(5871)) and (layer2_outputs(3825)));
    layer3_outputs(5968) <= not(layer2_outputs(5654));
    layer3_outputs(5969) <= layer2_outputs(1640);
    layer3_outputs(5970) <= not(layer2_outputs(7674)) or (layer2_outputs(4505));
    layer3_outputs(5971) <= not(layer2_outputs(5964));
    layer3_outputs(5972) <= (layer2_outputs(4491)) and (layer2_outputs(2035));
    layer3_outputs(5973) <= '0';
    layer3_outputs(5974) <= not(layer2_outputs(4018)) or (layer2_outputs(2155));
    layer3_outputs(5975) <= not((layer2_outputs(2836)) xor (layer2_outputs(4594)));
    layer3_outputs(5976) <= layer2_outputs(3703);
    layer3_outputs(5977) <= layer2_outputs(4951);
    layer3_outputs(5978) <= not((layer2_outputs(4151)) or (layer2_outputs(3465)));
    layer3_outputs(5979) <= layer2_outputs(2463);
    layer3_outputs(5980) <= layer2_outputs(2537);
    layer3_outputs(5981) <= not(layer2_outputs(659));
    layer3_outputs(5982) <= (layer2_outputs(3068)) and not (layer2_outputs(2021));
    layer3_outputs(5983) <= not(layer2_outputs(877));
    layer3_outputs(5984) <= not(layer2_outputs(6521));
    layer3_outputs(5985) <= (layer2_outputs(3313)) xor (layer2_outputs(5833));
    layer3_outputs(5986) <= not(layer2_outputs(4985));
    layer3_outputs(5987) <= not((layer2_outputs(589)) or (layer2_outputs(840)));
    layer3_outputs(5988) <= layer2_outputs(5451);
    layer3_outputs(5989) <= not(layer2_outputs(1190)) or (layer2_outputs(4622));
    layer3_outputs(5990) <= (layer2_outputs(1476)) and (layer2_outputs(3362));
    layer3_outputs(5991) <= layer2_outputs(5207);
    layer3_outputs(5992) <= '0';
    layer3_outputs(5993) <= not((layer2_outputs(36)) or (layer2_outputs(4408)));
    layer3_outputs(5994) <= not(layer2_outputs(6335));
    layer3_outputs(5995) <= layer2_outputs(5047);
    layer3_outputs(5996) <= (layer2_outputs(3592)) and not (layer2_outputs(5934));
    layer3_outputs(5997) <= (layer2_outputs(1048)) or (layer2_outputs(6288));
    layer3_outputs(5998) <= layer2_outputs(2594);
    layer3_outputs(5999) <= '1';
    layer3_outputs(6000) <= (layer2_outputs(6445)) or (layer2_outputs(768));
    layer3_outputs(6001) <= (layer2_outputs(4764)) and not (layer2_outputs(2915));
    layer3_outputs(6002) <= not(layer2_outputs(10)) or (layer2_outputs(6550));
    layer3_outputs(6003) <= layer2_outputs(768);
    layer3_outputs(6004) <= layer2_outputs(3195);
    layer3_outputs(6005) <= '0';
    layer3_outputs(6006) <= (layer2_outputs(2597)) and (layer2_outputs(3428));
    layer3_outputs(6007) <= (layer2_outputs(1439)) or (layer2_outputs(1801));
    layer3_outputs(6008) <= not(layer2_outputs(1176)) or (layer2_outputs(1165));
    layer3_outputs(6009) <= not(layer2_outputs(525));
    layer3_outputs(6010) <= layer2_outputs(4173);
    layer3_outputs(6011) <= (layer2_outputs(7066)) and (layer2_outputs(570));
    layer3_outputs(6012) <= not((layer2_outputs(7000)) or (layer2_outputs(5903)));
    layer3_outputs(6013) <= (layer2_outputs(5374)) and not (layer2_outputs(1761));
    layer3_outputs(6014) <= not(layer2_outputs(1635));
    layer3_outputs(6015) <= not(layer2_outputs(4735)) or (layer2_outputs(779));
    layer3_outputs(6016) <= not(layer2_outputs(6342));
    layer3_outputs(6017) <= layer2_outputs(2189);
    layer3_outputs(6018) <= not((layer2_outputs(2378)) xor (layer2_outputs(180)));
    layer3_outputs(6019) <= layer2_outputs(1547);
    layer3_outputs(6020) <= layer2_outputs(7661);
    layer3_outputs(6021) <= not((layer2_outputs(7473)) and (layer2_outputs(6553)));
    layer3_outputs(6022) <= '0';
    layer3_outputs(6023) <= (layer2_outputs(1127)) or (layer2_outputs(674));
    layer3_outputs(6024) <= not(layer2_outputs(1107));
    layer3_outputs(6025) <= (layer2_outputs(6823)) and not (layer2_outputs(1257));
    layer3_outputs(6026) <= (layer2_outputs(7201)) and (layer2_outputs(4590));
    layer3_outputs(6027) <= '0';
    layer3_outputs(6028) <= not(layer2_outputs(7624));
    layer3_outputs(6029) <= '0';
    layer3_outputs(6030) <= layer2_outputs(7664);
    layer3_outputs(6031) <= not(layer2_outputs(7061)) or (layer2_outputs(1522));
    layer3_outputs(6032) <= not((layer2_outputs(7655)) or (layer2_outputs(2994)));
    layer3_outputs(6033) <= layer2_outputs(5583);
    layer3_outputs(6034) <= not(layer2_outputs(3398)) or (layer2_outputs(2583));
    layer3_outputs(6035) <= layer2_outputs(6397);
    layer3_outputs(6036) <= layer2_outputs(4138);
    layer3_outputs(6037) <= not(layer2_outputs(304)) or (layer2_outputs(5902));
    layer3_outputs(6038) <= not(layer2_outputs(6783));
    layer3_outputs(6039) <= not((layer2_outputs(7103)) and (layer2_outputs(1945)));
    layer3_outputs(6040) <= (layer2_outputs(3450)) xor (layer2_outputs(6784));
    layer3_outputs(6041) <= layer2_outputs(5008);
    layer3_outputs(6042) <= (layer2_outputs(2845)) or (layer2_outputs(6846));
    layer3_outputs(6043) <= not(layer2_outputs(3779)) or (layer2_outputs(6609));
    layer3_outputs(6044) <= layer2_outputs(6117);
    layer3_outputs(6045) <= '1';
    layer3_outputs(6046) <= layer2_outputs(3049);
    layer3_outputs(6047) <= not((layer2_outputs(7572)) or (layer2_outputs(3182)));
    layer3_outputs(6048) <= (layer2_outputs(6365)) and not (layer2_outputs(5931));
    layer3_outputs(6049) <= not((layer2_outputs(5438)) and (layer2_outputs(4581)));
    layer3_outputs(6050) <= (layer2_outputs(7462)) and not (layer2_outputs(5216));
    layer3_outputs(6051) <= not((layer2_outputs(4246)) or (layer2_outputs(7531)));
    layer3_outputs(6052) <= '1';
    layer3_outputs(6053) <= not(layer2_outputs(1213)) or (layer2_outputs(7413));
    layer3_outputs(6054) <= '0';
    layer3_outputs(6055) <= layer2_outputs(831);
    layer3_outputs(6056) <= '1';
    layer3_outputs(6057) <= '0';
    layer3_outputs(6058) <= not((layer2_outputs(1791)) and (layer2_outputs(2166)));
    layer3_outputs(6059) <= not((layer2_outputs(7665)) or (layer2_outputs(5128)));
    layer3_outputs(6060) <= not(layer2_outputs(2962)) or (layer2_outputs(2055));
    layer3_outputs(6061) <= (layer2_outputs(3739)) or (layer2_outputs(1894));
    layer3_outputs(6062) <= not(layer2_outputs(6611));
    layer3_outputs(6063) <= '0';
    layer3_outputs(6064) <= not(layer2_outputs(6515)) or (layer2_outputs(2269));
    layer3_outputs(6065) <= '0';
    layer3_outputs(6066) <= not(layer2_outputs(4427));
    layer3_outputs(6067) <= (layer2_outputs(2515)) or (layer2_outputs(1539));
    layer3_outputs(6068) <= layer2_outputs(5477);
    layer3_outputs(6069) <= '0';
    layer3_outputs(6070) <= not(layer2_outputs(290));
    layer3_outputs(6071) <= not((layer2_outputs(4627)) and (layer2_outputs(1014)));
    layer3_outputs(6072) <= (layer2_outputs(6965)) and not (layer2_outputs(5484));
    layer3_outputs(6073) <= not(layer2_outputs(6037)) or (layer2_outputs(3167));
    layer3_outputs(6074) <= not(layer2_outputs(2122));
    layer3_outputs(6075) <= '1';
    layer3_outputs(6076) <= not(layer2_outputs(426));
    layer3_outputs(6077) <= not(layer2_outputs(3582)) or (layer2_outputs(3204));
    layer3_outputs(6078) <= layer2_outputs(3218);
    layer3_outputs(6079) <= not(layer2_outputs(6193)) or (layer2_outputs(3338));
    layer3_outputs(6080) <= layer2_outputs(6066);
    layer3_outputs(6081) <= (layer2_outputs(1236)) and not (layer2_outputs(4173));
    layer3_outputs(6082) <= (layer2_outputs(5599)) or (layer2_outputs(183));
    layer3_outputs(6083) <= not(layer2_outputs(6905));
    layer3_outputs(6084) <= '0';
    layer3_outputs(6085) <= layer2_outputs(1063);
    layer3_outputs(6086) <= (layer2_outputs(22)) and not (layer2_outputs(2617));
    layer3_outputs(6087) <= not((layer2_outputs(5122)) or (layer2_outputs(3102)));
    layer3_outputs(6088) <= '1';
    layer3_outputs(6089) <= not((layer2_outputs(2003)) or (layer2_outputs(3999)));
    layer3_outputs(6090) <= (layer2_outputs(7001)) and not (layer2_outputs(1770));
    layer3_outputs(6091) <= (layer2_outputs(236)) and not (layer2_outputs(703));
    layer3_outputs(6092) <= not(layer2_outputs(3426));
    layer3_outputs(6093) <= '1';
    layer3_outputs(6094) <= '0';
    layer3_outputs(6095) <= (layer2_outputs(7629)) or (layer2_outputs(6121));
    layer3_outputs(6096) <= not(layer2_outputs(3569));
    layer3_outputs(6097) <= not(layer2_outputs(5168));
    layer3_outputs(6098) <= layer2_outputs(3121);
    layer3_outputs(6099) <= not(layer2_outputs(5615));
    layer3_outputs(6100) <= layer2_outputs(168);
    layer3_outputs(6101) <= (layer2_outputs(3260)) and not (layer2_outputs(3025));
    layer3_outputs(6102) <= not(layer2_outputs(5171)) or (layer2_outputs(5191));
    layer3_outputs(6103) <= not(layer2_outputs(6581)) or (layer2_outputs(4381));
    layer3_outputs(6104) <= not(layer2_outputs(5665));
    layer3_outputs(6105) <= layer2_outputs(7086);
    layer3_outputs(6106) <= (layer2_outputs(2618)) and not (layer2_outputs(4362));
    layer3_outputs(6107) <= '1';
    layer3_outputs(6108) <= not(layer2_outputs(4522));
    layer3_outputs(6109) <= not((layer2_outputs(1215)) xor (layer2_outputs(1997)));
    layer3_outputs(6110) <= (layer2_outputs(391)) and (layer2_outputs(4310));
    layer3_outputs(6111) <= (layer2_outputs(2582)) and (layer2_outputs(727));
    layer3_outputs(6112) <= not(layer2_outputs(4964));
    layer3_outputs(6113) <= layer2_outputs(7566);
    layer3_outputs(6114) <= not((layer2_outputs(6866)) or (layer2_outputs(5625)));
    layer3_outputs(6115) <= '1';
    layer3_outputs(6116) <= layer2_outputs(3808);
    layer3_outputs(6117) <= (layer2_outputs(795)) and not (layer2_outputs(4496));
    layer3_outputs(6118) <= layer2_outputs(7164);
    layer3_outputs(6119) <= '1';
    layer3_outputs(6120) <= '0';
    layer3_outputs(6121) <= '0';
    layer3_outputs(6122) <= not(layer2_outputs(2771));
    layer3_outputs(6123) <= (layer2_outputs(780)) and not (layer2_outputs(3946));
    layer3_outputs(6124) <= (layer2_outputs(7409)) and not (layer2_outputs(2642));
    layer3_outputs(6125) <= not((layer2_outputs(4404)) or (layer2_outputs(468)));
    layer3_outputs(6126) <= not(layer2_outputs(5163));
    layer3_outputs(6127) <= (layer2_outputs(5417)) or (layer2_outputs(738));
    layer3_outputs(6128) <= not(layer2_outputs(341));
    layer3_outputs(6129) <= not(layer2_outputs(2319)) or (layer2_outputs(1748));
    layer3_outputs(6130) <= (layer2_outputs(1917)) and not (layer2_outputs(3872));
    layer3_outputs(6131) <= not(layer2_outputs(6465)) or (layer2_outputs(5974));
    layer3_outputs(6132) <= not(layer2_outputs(2767)) or (layer2_outputs(5865));
    layer3_outputs(6133) <= not(layer2_outputs(3204)) or (layer2_outputs(2355));
    layer3_outputs(6134) <= layer2_outputs(1150);
    layer3_outputs(6135) <= layer2_outputs(2520);
    layer3_outputs(6136) <= not(layer2_outputs(5530)) or (layer2_outputs(4870));
    layer3_outputs(6137) <= '0';
    layer3_outputs(6138) <= not(layer2_outputs(1438));
    layer3_outputs(6139) <= layer2_outputs(2985);
    layer3_outputs(6140) <= not((layer2_outputs(64)) or (layer2_outputs(4717)));
    layer3_outputs(6141) <= layer2_outputs(2275);
    layer3_outputs(6142) <= not((layer2_outputs(4670)) or (layer2_outputs(7334)));
    layer3_outputs(6143) <= (layer2_outputs(3787)) or (layer2_outputs(4044));
    layer3_outputs(6144) <= '0';
    layer3_outputs(6145) <= layer2_outputs(3031);
    layer3_outputs(6146) <= not((layer2_outputs(2506)) xor (layer2_outputs(6479)));
    layer3_outputs(6147) <= layer2_outputs(6613);
    layer3_outputs(6148) <= (layer2_outputs(1287)) or (layer2_outputs(1857));
    layer3_outputs(6149) <= not(layer2_outputs(6348)) or (layer2_outputs(2013));
    layer3_outputs(6150) <= (layer2_outputs(6558)) and not (layer2_outputs(2064));
    layer3_outputs(6151) <= (layer2_outputs(763)) and not (layer2_outputs(1180));
    layer3_outputs(6152) <= not(layer2_outputs(5498)) or (layer2_outputs(4032));
    layer3_outputs(6153) <= '0';
    layer3_outputs(6154) <= layer2_outputs(612);
    layer3_outputs(6155) <= (layer2_outputs(860)) and not (layer2_outputs(2140));
    layer3_outputs(6156) <= not((layer2_outputs(5766)) and (layer2_outputs(2710)));
    layer3_outputs(6157) <= not(layer2_outputs(6214)) or (layer2_outputs(6927));
    layer3_outputs(6158) <= not((layer2_outputs(301)) and (layer2_outputs(718)));
    layer3_outputs(6159) <= not(layer2_outputs(7042));
    layer3_outputs(6160) <= not((layer2_outputs(578)) and (layer2_outputs(5997)));
    layer3_outputs(6161) <= not(layer2_outputs(7594));
    layer3_outputs(6162) <= '1';
    layer3_outputs(6163) <= not(layer2_outputs(7064)) or (layer2_outputs(4548));
    layer3_outputs(6164) <= not((layer2_outputs(5130)) or (layer2_outputs(4301)));
    layer3_outputs(6165) <= layer2_outputs(2070);
    layer3_outputs(6166) <= '1';
    layer3_outputs(6167) <= (layer2_outputs(5768)) and (layer2_outputs(6784));
    layer3_outputs(6168) <= (layer2_outputs(4687)) and not (layer2_outputs(7115));
    layer3_outputs(6169) <= '0';
    layer3_outputs(6170) <= not(layer2_outputs(2778)) or (layer2_outputs(837));
    layer3_outputs(6171) <= not(layer2_outputs(564)) or (layer2_outputs(12));
    layer3_outputs(6172) <= not(layer2_outputs(5164)) or (layer2_outputs(7357));
    layer3_outputs(6173) <= (layer2_outputs(1720)) and (layer2_outputs(705));
    layer3_outputs(6174) <= layer2_outputs(6043);
    layer3_outputs(6175) <= (layer2_outputs(823)) and not (layer2_outputs(2459));
    layer3_outputs(6176) <= (layer2_outputs(593)) and not (layer2_outputs(3083));
    layer3_outputs(6177) <= not((layer2_outputs(6814)) xor (layer2_outputs(5212)));
    layer3_outputs(6178) <= (layer2_outputs(4859)) and (layer2_outputs(255));
    layer3_outputs(6179) <= not(layer2_outputs(2611));
    layer3_outputs(6180) <= '0';
    layer3_outputs(6181) <= not((layer2_outputs(2695)) or (layer2_outputs(6293)));
    layer3_outputs(6182) <= not(layer2_outputs(2963)) or (layer2_outputs(5076));
    layer3_outputs(6183) <= '1';
    layer3_outputs(6184) <= (layer2_outputs(5137)) and not (layer2_outputs(3116));
    layer3_outputs(6185) <= not((layer2_outputs(810)) or (layer2_outputs(289)));
    layer3_outputs(6186) <= layer2_outputs(6232);
    layer3_outputs(6187) <= layer2_outputs(452);
    layer3_outputs(6188) <= not(layer2_outputs(527));
    layer3_outputs(6189) <= (layer2_outputs(6666)) or (layer2_outputs(7032));
    layer3_outputs(6190) <= not(layer2_outputs(313));
    layer3_outputs(6191) <= layer2_outputs(2116);
    layer3_outputs(6192) <= (layer2_outputs(5055)) xor (layer2_outputs(5726));
    layer3_outputs(6193) <= (layer2_outputs(6271)) xor (layer2_outputs(164));
    layer3_outputs(6194) <= not((layer2_outputs(2208)) or (layer2_outputs(6588)));
    layer3_outputs(6195) <= (layer2_outputs(2386)) and not (layer2_outputs(1041));
    layer3_outputs(6196) <= (layer2_outputs(1033)) and not (layer2_outputs(1394));
    layer3_outputs(6197) <= '1';
    layer3_outputs(6198) <= (layer2_outputs(7002)) and not (layer2_outputs(4959));
    layer3_outputs(6199) <= layer2_outputs(178);
    layer3_outputs(6200) <= (layer2_outputs(7350)) xor (layer2_outputs(604));
    layer3_outputs(6201) <= not(layer2_outputs(6562)) or (layer2_outputs(6798));
    layer3_outputs(6202) <= not(layer2_outputs(6516));
    layer3_outputs(6203) <= not(layer2_outputs(2371));
    layer3_outputs(6204) <= '0';
    layer3_outputs(6205) <= (layer2_outputs(4019)) and not (layer2_outputs(6136));
    layer3_outputs(6206) <= (layer2_outputs(3038)) or (layer2_outputs(4525));
    layer3_outputs(6207) <= not((layer2_outputs(2965)) and (layer2_outputs(2885)));
    layer3_outputs(6208) <= (layer2_outputs(5518)) and (layer2_outputs(1363));
    layer3_outputs(6209) <= not(layer2_outputs(2596)) or (layer2_outputs(2303));
    layer3_outputs(6210) <= layer2_outputs(2977);
    layer3_outputs(6211) <= not(layer2_outputs(4563));
    layer3_outputs(6212) <= '0';
    layer3_outputs(6213) <= not(layer2_outputs(3954)) or (layer2_outputs(964));
    layer3_outputs(6214) <= not((layer2_outputs(7673)) and (layer2_outputs(447)));
    layer3_outputs(6215) <= not((layer2_outputs(5708)) and (layer2_outputs(3773)));
    layer3_outputs(6216) <= not((layer2_outputs(1203)) and (layer2_outputs(4120)));
    layer3_outputs(6217) <= not(layer2_outputs(3768)) or (layer2_outputs(152));
    layer3_outputs(6218) <= layer2_outputs(2664);
    layer3_outputs(6219) <= not(layer2_outputs(2338));
    layer3_outputs(6220) <= (layer2_outputs(4293)) and (layer2_outputs(64));
    layer3_outputs(6221) <= not((layer2_outputs(5266)) and (layer2_outputs(2115)));
    layer3_outputs(6222) <= (layer2_outputs(2038)) xor (layer2_outputs(350));
    layer3_outputs(6223) <= '1';
    layer3_outputs(6224) <= (layer2_outputs(4723)) or (layer2_outputs(5881));
    layer3_outputs(6225) <= not((layer2_outputs(5231)) xor (layer2_outputs(6989)));
    layer3_outputs(6226) <= not((layer2_outputs(4266)) or (layer2_outputs(1726)));
    layer3_outputs(6227) <= not((layer2_outputs(6652)) and (layer2_outputs(4377)));
    layer3_outputs(6228) <= not(layer2_outputs(7468));
    layer3_outputs(6229) <= not(layer2_outputs(936));
    layer3_outputs(6230) <= layer2_outputs(3206);
    layer3_outputs(6231) <= not((layer2_outputs(2184)) and (layer2_outputs(3789)));
    layer3_outputs(6232) <= not(layer2_outputs(4844));
    layer3_outputs(6233) <= layer2_outputs(3728);
    layer3_outputs(6234) <= not(layer2_outputs(5514)) or (layer2_outputs(5289));
    layer3_outputs(6235) <= not(layer2_outputs(480));
    layer3_outputs(6236) <= not(layer2_outputs(4297));
    layer3_outputs(6237) <= not((layer2_outputs(5797)) or (layer2_outputs(4559)));
    layer3_outputs(6238) <= '0';
    layer3_outputs(6239) <= not(layer2_outputs(4999));
    layer3_outputs(6240) <= (layer2_outputs(423)) and (layer2_outputs(7479));
    layer3_outputs(6241) <= (layer2_outputs(4436)) or (layer2_outputs(481));
    layer3_outputs(6242) <= layer2_outputs(601);
    layer3_outputs(6243) <= layer2_outputs(2870);
    layer3_outputs(6244) <= '0';
    layer3_outputs(6245) <= '0';
    layer3_outputs(6246) <= not((layer2_outputs(6315)) and (layer2_outputs(4579)));
    layer3_outputs(6247) <= not((layer2_outputs(4945)) and (layer2_outputs(4005)));
    layer3_outputs(6248) <= layer2_outputs(2177);
    layer3_outputs(6249) <= not(layer2_outputs(477)) or (layer2_outputs(4208));
    layer3_outputs(6250) <= not(layer2_outputs(1922));
    layer3_outputs(6251) <= (layer2_outputs(2445)) or (layer2_outputs(5750));
    layer3_outputs(6252) <= '1';
    layer3_outputs(6253) <= not(layer2_outputs(3320));
    layer3_outputs(6254) <= (layer2_outputs(2703)) xor (layer2_outputs(7647));
    layer3_outputs(6255) <= '0';
    layer3_outputs(6256) <= not(layer2_outputs(1792));
    layer3_outputs(6257) <= not(layer2_outputs(3788)) or (layer2_outputs(7619));
    layer3_outputs(6258) <= (layer2_outputs(61)) and not (layer2_outputs(3192));
    layer3_outputs(6259) <= (layer2_outputs(2789)) and (layer2_outputs(4361));
    layer3_outputs(6260) <= not((layer2_outputs(6363)) or (layer2_outputs(6269)));
    layer3_outputs(6261) <= '0';
    layer3_outputs(6262) <= (layer2_outputs(7275)) or (layer2_outputs(4965));
    layer3_outputs(6263) <= not(layer2_outputs(7185));
    layer3_outputs(6264) <= not(layer2_outputs(3151)) or (layer2_outputs(5382));
    layer3_outputs(6265) <= layer2_outputs(1361);
    layer3_outputs(6266) <= not((layer2_outputs(1545)) or (layer2_outputs(3614)));
    layer3_outputs(6267) <= not(layer2_outputs(130)) or (layer2_outputs(2699));
    layer3_outputs(6268) <= not((layer2_outputs(515)) xor (layer2_outputs(1083)));
    layer3_outputs(6269) <= layer2_outputs(2558);
    layer3_outputs(6270) <= not(layer2_outputs(7362)) or (layer2_outputs(1262));
    layer3_outputs(6271) <= '0';
    layer3_outputs(6272) <= not(layer2_outputs(3412));
    layer3_outputs(6273) <= (layer2_outputs(5019)) and (layer2_outputs(5529));
    layer3_outputs(6274) <= not((layer2_outputs(5831)) and (layer2_outputs(1808)));
    layer3_outputs(6275) <= layer2_outputs(422);
    layer3_outputs(6276) <= '0';
    layer3_outputs(6277) <= not(layer2_outputs(498));
    layer3_outputs(6278) <= not((layer2_outputs(6926)) and (layer2_outputs(3063)));
    layer3_outputs(6279) <= layer2_outputs(661);
    layer3_outputs(6280) <= layer2_outputs(5635);
    layer3_outputs(6281) <= (layer2_outputs(1290)) and not (layer2_outputs(2082));
    layer3_outputs(6282) <= layer2_outputs(4560);
    layer3_outputs(6283) <= layer2_outputs(5355);
    layer3_outputs(6284) <= (layer2_outputs(3177)) and not (layer2_outputs(3837));
    layer3_outputs(6285) <= '0';
    layer3_outputs(6286) <= layer2_outputs(4050);
    layer3_outputs(6287) <= not((layer2_outputs(1713)) and (layer2_outputs(7111)));
    layer3_outputs(6288) <= not(layer2_outputs(5510));
    layer3_outputs(6289) <= not(layer2_outputs(3337));
    layer3_outputs(6290) <= '0';
    layer3_outputs(6291) <= not((layer2_outputs(3938)) or (layer2_outputs(4303)));
    layer3_outputs(6292) <= (layer2_outputs(2543)) and (layer2_outputs(2686));
    layer3_outputs(6293) <= layer2_outputs(6463);
    layer3_outputs(6294) <= not(layer2_outputs(3004));
    layer3_outputs(6295) <= not((layer2_outputs(2365)) and (layer2_outputs(1836)));
    layer3_outputs(6296) <= layer2_outputs(2927);
    layer3_outputs(6297) <= layer2_outputs(1434);
    layer3_outputs(6298) <= layer2_outputs(6991);
    layer3_outputs(6299) <= not((layer2_outputs(1695)) xor (layer2_outputs(4708)));
    layer3_outputs(6300) <= layer2_outputs(1346);
    layer3_outputs(6301) <= (layer2_outputs(3937)) and not (layer2_outputs(4057));
    layer3_outputs(6302) <= not(layer2_outputs(1473)) or (layer2_outputs(1666));
    layer3_outputs(6303) <= layer2_outputs(2358);
    layer3_outputs(6304) <= not(layer2_outputs(6528));
    layer3_outputs(6305) <= not(layer2_outputs(523));
    layer3_outputs(6306) <= not(layer2_outputs(4990));
    layer3_outputs(6307) <= layer2_outputs(3669);
    layer3_outputs(6308) <= not(layer2_outputs(7089));
    layer3_outputs(6309) <= not(layer2_outputs(550));
    layer3_outputs(6310) <= not(layer2_outputs(395));
    layer3_outputs(6311) <= not(layer2_outputs(4460));
    layer3_outputs(6312) <= (layer2_outputs(2980)) and not (layer2_outputs(6385));
    layer3_outputs(6313) <= not(layer2_outputs(6440));
    layer3_outputs(6314) <= not(layer2_outputs(3471));
    layer3_outputs(6315) <= not((layer2_outputs(639)) or (layer2_outputs(5318)));
    layer3_outputs(6316) <= not((layer2_outputs(3988)) xor (layer2_outputs(1751)));
    layer3_outputs(6317) <= layer2_outputs(4853);
    layer3_outputs(6318) <= not(layer2_outputs(4744)) or (layer2_outputs(582));
    layer3_outputs(6319) <= '0';
    layer3_outputs(6320) <= layer2_outputs(4589);
    layer3_outputs(6321) <= not(layer2_outputs(3656));
    layer3_outputs(6322) <= not((layer2_outputs(5525)) or (layer2_outputs(7260)));
    layer3_outputs(6323) <= not((layer2_outputs(1975)) xor (layer2_outputs(4983)));
    layer3_outputs(6324) <= not(layer2_outputs(1421)) or (layer2_outputs(1123));
    layer3_outputs(6325) <= not((layer2_outputs(117)) or (layer2_outputs(156)));
    layer3_outputs(6326) <= layer2_outputs(5141);
    layer3_outputs(6327) <= not((layer2_outputs(4503)) and (layer2_outputs(6462)));
    layer3_outputs(6328) <= layer2_outputs(2572);
    layer3_outputs(6329) <= not((layer2_outputs(3980)) and (layer2_outputs(4822)));
    layer3_outputs(6330) <= not(layer2_outputs(1826));
    layer3_outputs(6331) <= not(layer2_outputs(1108)) or (layer2_outputs(5661));
    layer3_outputs(6332) <= not(layer2_outputs(7594)) or (layer2_outputs(2056));
    layer3_outputs(6333) <= (layer2_outputs(6668)) and not (layer2_outputs(6132));
    layer3_outputs(6334) <= not((layer2_outputs(1573)) and (layer2_outputs(277)));
    layer3_outputs(6335) <= not(layer2_outputs(5534));
    layer3_outputs(6336) <= '1';
    layer3_outputs(6337) <= layer2_outputs(4409);
    layer3_outputs(6338) <= not(layer2_outputs(1404));
    layer3_outputs(6339) <= '0';
    layer3_outputs(6340) <= not(layer2_outputs(5672)) or (layer2_outputs(3947));
    layer3_outputs(6341) <= not((layer2_outputs(30)) and (layer2_outputs(750)));
    layer3_outputs(6342) <= layer2_outputs(5590);
    layer3_outputs(6343) <= (layer2_outputs(102)) and not (layer2_outputs(884));
    layer3_outputs(6344) <= not(layer2_outputs(6003));
    layer3_outputs(6345) <= not(layer2_outputs(2103)) or (layer2_outputs(871));
    layer3_outputs(6346) <= not((layer2_outputs(7628)) or (layer2_outputs(8)));
    layer3_outputs(6347) <= (layer2_outputs(456)) or (layer2_outputs(6683));
    layer3_outputs(6348) <= not((layer2_outputs(610)) and (layer2_outputs(2516)));
    layer3_outputs(6349) <= not(layer2_outputs(4153));
    layer3_outputs(6350) <= (layer2_outputs(3632)) or (layer2_outputs(5889));
    layer3_outputs(6351) <= not((layer2_outputs(6636)) or (layer2_outputs(2877)));
    layer3_outputs(6352) <= (layer2_outputs(3509)) and not (layer2_outputs(6295));
    layer3_outputs(6353) <= not(layer2_outputs(2783));
    layer3_outputs(6354) <= layer2_outputs(6245);
    layer3_outputs(6355) <= (layer2_outputs(4152)) or (layer2_outputs(3519));
    layer3_outputs(6356) <= not((layer2_outputs(4155)) and (layer2_outputs(4268)));
    layer3_outputs(6357) <= not((layer2_outputs(4162)) xor (layer2_outputs(912)));
    layer3_outputs(6358) <= (layer2_outputs(1028)) and not (layer2_outputs(2158));
    layer3_outputs(6359) <= not((layer2_outputs(2049)) or (layer2_outputs(2913)));
    layer3_outputs(6360) <= not(layer2_outputs(4167)) or (layer2_outputs(1928));
    layer3_outputs(6361) <= not(layer2_outputs(3573));
    layer3_outputs(6362) <= not((layer2_outputs(7142)) and (layer2_outputs(3655)));
    layer3_outputs(6363) <= '0';
    layer3_outputs(6364) <= layer2_outputs(3052);
    layer3_outputs(6365) <= not((layer2_outputs(4553)) or (layer2_outputs(2467)));
    layer3_outputs(6366) <= layer2_outputs(1281);
    layer3_outputs(6367) <= '1';
    layer3_outputs(6368) <= '1';
    layer3_outputs(6369) <= '1';
    layer3_outputs(6370) <= not(layer2_outputs(4022)) or (layer2_outputs(128));
    layer3_outputs(6371) <= not((layer2_outputs(5881)) or (layer2_outputs(7038)));
    layer3_outputs(6372) <= (layer2_outputs(7335)) and not (layer2_outputs(3892));
    layer3_outputs(6373) <= layer2_outputs(3757);
    layer3_outputs(6374) <= not((layer2_outputs(88)) or (layer2_outputs(1318)));
    layer3_outputs(6375) <= layer2_outputs(3390);
    layer3_outputs(6376) <= layer2_outputs(80);
    layer3_outputs(6377) <= not(layer2_outputs(1072));
    layer3_outputs(6378) <= not((layer2_outputs(3017)) and (layer2_outputs(3643)));
    layer3_outputs(6379) <= layer2_outputs(1459);
    layer3_outputs(6380) <= layer2_outputs(6086);
    layer3_outputs(6381) <= (layer2_outputs(2865)) and not (layer2_outputs(6266));
    layer3_outputs(6382) <= not(layer2_outputs(273));
    layer3_outputs(6383) <= (layer2_outputs(4079)) or (layer2_outputs(6413));
    layer3_outputs(6384) <= (layer2_outputs(5282)) and not (layer2_outputs(1903));
    layer3_outputs(6385) <= layer2_outputs(5454);
    layer3_outputs(6386) <= (layer2_outputs(5544)) and not (layer2_outputs(1375));
    layer3_outputs(6387) <= not(layer2_outputs(6598));
    layer3_outputs(6388) <= not((layer2_outputs(5031)) xor (layer2_outputs(513)));
    layer3_outputs(6389) <= not(layer2_outputs(6412));
    layer3_outputs(6390) <= not((layer2_outputs(6146)) or (layer2_outputs(812)));
    layer3_outputs(6391) <= not(layer2_outputs(7653));
    layer3_outputs(6392) <= not(layer2_outputs(7533));
    layer3_outputs(6393) <= not(layer2_outputs(5103));
    layer3_outputs(6394) <= layer2_outputs(3468);
    layer3_outputs(6395) <= (layer2_outputs(7613)) and not (layer2_outputs(6744));
    layer3_outputs(6396) <= not(layer2_outputs(7001));
    layer3_outputs(6397) <= (layer2_outputs(3193)) and (layer2_outputs(4085));
    layer3_outputs(6398) <= not((layer2_outputs(247)) and (layer2_outputs(6567)));
    layer3_outputs(6399) <= (layer2_outputs(6224)) and not (layer2_outputs(2436));
    layer3_outputs(6400) <= (layer2_outputs(5406)) and not (layer2_outputs(7449));
    layer3_outputs(6401) <= layer2_outputs(2900);
    layer3_outputs(6402) <= not((layer2_outputs(1230)) and (layer2_outputs(5773)));
    layer3_outputs(6403) <= not((layer2_outputs(7610)) and (layer2_outputs(5394)));
    layer3_outputs(6404) <= (layer2_outputs(6336)) and not (layer2_outputs(489));
    layer3_outputs(6405) <= not(layer2_outputs(2420));
    layer3_outputs(6406) <= '0';
    layer3_outputs(6407) <= not(layer2_outputs(4976));
    layer3_outputs(6408) <= not(layer2_outputs(2376));
    layer3_outputs(6409) <= layer2_outputs(6473);
    layer3_outputs(6410) <= layer2_outputs(41);
    layer3_outputs(6411) <= layer2_outputs(270);
    layer3_outputs(6412) <= (layer2_outputs(5722)) and not (layer2_outputs(4644));
    layer3_outputs(6413) <= '1';
    layer3_outputs(6414) <= (layer2_outputs(6191)) and not (layer2_outputs(6450));
    layer3_outputs(6415) <= layer2_outputs(4328);
    layer3_outputs(6416) <= (layer2_outputs(4738)) and not (layer2_outputs(3847));
    layer3_outputs(6417) <= not(layer2_outputs(5859));
    layer3_outputs(6418) <= layer2_outputs(5457);
    layer3_outputs(6419) <= not(layer2_outputs(5500));
    layer3_outputs(6420) <= not(layer2_outputs(3969)) or (layer2_outputs(7227));
    layer3_outputs(6421) <= (layer2_outputs(1104)) or (layer2_outputs(5420));
    layer3_outputs(6422) <= not((layer2_outputs(6728)) or (layer2_outputs(1330)));
    layer3_outputs(6423) <= layer2_outputs(7418);
    layer3_outputs(6424) <= layer2_outputs(6312);
    layer3_outputs(6425) <= not(layer2_outputs(2645));
    layer3_outputs(6426) <= (layer2_outputs(3812)) and not (layer2_outputs(3700));
    layer3_outputs(6427) <= not((layer2_outputs(1876)) or (layer2_outputs(1410)));
    layer3_outputs(6428) <= layer2_outputs(1579);
    layer3_outputs(6429) <= not(layer2_outputs(149)) or (layer2_outputs(2112));
    layer3_outputs(6430) <= not((layer2_outputs(5317)) and (layer2_outputs(7087)));
    layer3_outputs(6431) <= not(layer2_outputs(4250));
    layer3_outputs(6432) <= not(layer2_outputs(4023));
    layer3_outputs(6433) <= (layer2_outputs(80)) and (layer2_outputs(1556));
    layer3_outputs(6434) <= not(layer2_outputs(4484));
    layer3_outputs(6435) <= not(layer2_outputs(4943)) or (layer2_outputs(7663));
    layer3_outputs(6436) <= '0';
    layer3_outputs(6437) <= not((layer2_outputs(7130)) and (layer2_outputs(2731)));
    layer3_outputs(6438) <= (layer2_outputs(4090)) and (layer2_outputs(5312));
    layer3_outputs(6439) <= layer2_outputs(688);
    layer3_outputs(6440) <= layer2_outputs(2954);
    layer3_outputs(6441) <= not(layer2_outputs(803)) or (layer2_outputs(7549));
    layer3_outputs(6442) <= (layer2_outputs(1153)) and not (layer2_outputs(3521));
    layer3_outputs(6443) <= not((layer2_outputs(342)) xor (layer2_outputs(6950)));
    layer3_outputs(6444) <= not((layer2_outputs(5269)) xor (layer2_outputs(2640)));
    layer3_outputs(6445) <= layer2_outputs(5199);
    layer3_outputs(6446) <= (layer2_outputs(7189)) and not (layer2_outputs(1438));
    layer3_outputs(6447) <= not(layer2_outputs(3621));
    layer3_outputs(6448) <= not(layer2_outputs(740));
    layer3_outputs(6449) <= (layer2_outputs(5154)) or (layer2_outputs(4702));
    layer3_outputs(6450) <= not(layer2_outputs(5268));
    layer3_outputs(6451) <= not(layer2_outputs(5937));
    layer3_outputs(6452) <= layer2_outputs(2660);
    layer3_outputs(6453) <= not((layer2_outputs(5325)) and (layer2_outputs(2022)));
    layer3_outputs(6454) <= not(layer2_outputs(5849));
    layer3_outputs(6455) <= (layer2_outputs(1085)) and not (layer2_outputs(4345));
    layer3_outputs(6456) <= not(layer2_outputs(1907));
    layer3_outputs(6457) <= not(layer2_outputs(2903));
    layer3_outputs(6458) <= not((layer2_outputs(4763)) and (layer2_outputs(5734)));
    layer3_outputs(6459) <= not((layer2_outputs(7161)) or (layer2_outputs(1041)));
    layer3_outputs(6460) <= layer2_outputs(2159);
    layer3_outputs(6461) <= not((layer2_outputs(3856)) xor (layer2_outputs(2490)));
    layer3_outputs(6462) <= not(layer2_outputs(6040));
    layer3_outputs(6463) <= not(layer2_outputs(3453));
    layer3_outputs(6464) <= not(layer2_outputs(5378));
    layer3_outputs(6465) <= (layer2_outputs(7650)) and not (layer2_outputs(2485));
    layer3_outputs(6466) <= (layer2_outputs(4099)) xor (layer2_outputs(969));
    layer3_outputs(6467) <= (layer2_outputs(5498)) and not (layer2_outputs(2737));
    layer3_outputs(6468) <= '0';
    layer3_outputs(6469) <= not(layer2_outputs(1472)) or (layer2_outputs(2448));
    layer3_outputs(6470) <= not(layer2_outputs(2953));
    layer3_outputs(6471) <= (layer2_outputs(7604)) xor (layer2_outputs(7519));
    layer3_outputs(6472) <= not(layer2_outputs(2555));
    layer3_outputs(6473) <= not(layer2_outputs(6929)) or (layer2_outputs(4669));
    layer3_outputs(6474) <= layer2_outputs(1626);
    layer3_outputs(6475) <= (layer2_outputs(2934)) and (layer2_outputs(6904));
    layer3_outputs(6476) <= '1';
    layer3_outputs(6477) <= (layer2_outputs(1867)) and not (layer2_outputs(7392));
    layer3_outputs(6478) <= '0';
    layer3_outputs(6479) <= not(layer2_outputs(1007)) or (layer2_outputs(5074));
    layer3_outputs(6480) <= not(layer2_outputs(865)) or (layer2_outputs(7366));
    layer3_outputs(6481) <= not(layer2_outputs(7020));
    layer3_outputs(6482) <= not(layer2_outputs(5491));
    layer3_outputs(6483) <= not(layer2_outputs(4733)) or (layer2_outputs(6986));
    layer3_outputs(6484) <= not((layer2_outputs(7208)) or (layer2_outputs(953)));
    layer3_outputs(6485) <= (layer2_outputs(5725)) and not (layer2_outputs(6693));
    layer3_outputs(6486) <= '1';
    layer3_outputs(6487) <= not((layer2_outputs(553)) and (layer2_outputs(5451)));
    layer3_outputs(6488) <= layer2_outputs(4904);
    layer3_outputs(6489) <= not(layer2_outputs(3810));
    layer3_outputs(6490) <= layer2_outputs(2936);
    layer3_outputs(6491) <= layer2_outputs(93);
    layer3_outputs(6492) <= not(layer2_outputs(6559)) or (layer2_outputs(6073));
    layer3_outputs(6493) <= not(layer2_outputs(4879));
    layer3_outputs(6494) <= (layer2_outputs(1158)) and not (layer2_outputs(5233));
    layer3_outputs(6495) <= not(layer2_outputs(1781));
    layer3_outputs(6496) <= not(layer2_outputs(1600)) or (layer2_outputs(7379));
    layer3_outputs(6497) <= (layer2_outputs(7190)) and not (layer2_outputs(1398));
    layer3_outputs(6498) <= not((layer2_outputs(6843)) or (layer2_outputs(1844)));
    layer3_outputs(6499) <= not(layer2_outputs(5879));
    layer3_outputs(6500) <= (layer2_outputs(5425)) and not (layer2_outputs(3811));
    layer3_outputs(6501) <= not(layer2_outputs(3336));
    layer3_outputs(6502) <= not(layer2_outputs(1378)) or (layer2_outputs(160));
    layer3_outputs(6503) <= (layer2_outputs(1771)) xor (layer2_outputs(2197));
    layer3_outputs(6504) <= '1';
    layer3_outputs(6505) <= (layer2_outputs(2361)) and (layer2_outputs(7245));
    layer3_outputs(6506) <= (layer2_outputs(7308)) or (layer2_outputs(6935));
    layer3_outputs(6507) <= not(layer2_outputs(6777));
    layer3_outputs(6508) <= not((layer2_outputs(6592)) and (layer2_outputs(3451)));
    layer3_outputs(6509) <= (layer2_outputs(2032)) and not (layer2_outputs(1795));
    layer3_outputs(6510) <= layer2_outputs(4935);
    layer3_outputs(6511) <= not(layer2_outputs(1213)) or (layer2_outputs(4945));
    layer3_outputs(6512) <= '1';
    layer3_outputs(6513) <= (layer2_outputs(3629)) and not (layer2_outputs(988));
    layer3_outputs(6514) <= (layer2_outputs(5597)) or (layer2_outputs(6824));
    layer3_outputs(6515) <= (layer2_outputs(7013)) or (layer2_outputs(6677));
    layer3_outputs(6516) <= not(layer2_outputs(6480));
    layer3_outputs(6517) <= not(layer2_outputs(4514)) or (layer2_outputs(5141));
    layer3_outputs(6518) <= not((layer2_outputs(6942)) and (layer2_outputs(5338)));
    layer3_outputs(6519) <= '0';
    layer3_outputs(6520) <= not(layer2_outputs(2813)) or (layer2_outputs(599));
    layer3_outputs(6521) <= layer2_outputs(6906);
    layer3_outputs(6522) <= not(layer2_outputs(4903)) or (layer2_outputs(1775));
    layer3_outputs(6523) <= not(layer2_outputs(939));
    layer3_outputs(6524) <= layer2_outputs(2409);
    layer3_outputs(6525) <= (layer2_outputs(4992)) and (layer2_outputs(187));
    layer3_outputs(6526) <= '0';
    layer3_outputs(6527) <= (layer2_outputs(2858)) or (layer2_outputs(95));
    layer3_outputs(6528) <= (layer2_outputs(3651)) and (layer2_outputs(3566));
    layer3_outputs(6529) <= '1';
    layer3_outputs(6530) <= (layer2_outputs(7371)) or (layer2_outputs(5307));
    layer3_outputs(6531) <= not((layer2_outputs(1707)) or (layer2_outputs(609)));
    layer3_outputs(6532) <= not(layer2_outputs(2829));
    layer3_outputs(6533) <= layer2_outputs(1553);
    layer3_outputs(6534) <= layer2_outputs(5437);
    layer3_outputs(6535) <= not(layer2_outputs(4595)) or (layer2_outputs(5455));
    layer3_outputs(6536) <= not(layer2_outputs(7364)) or (layer2_outputs(6027));
    layer3_outputs(6537) <= (layer2_outputs(4492)) and not (layer2_outputs(171));
    layer3_outputs(6538) <= '1';
    layer3_outputs(6539) <= layer2_outputs(6262);
    layer3_outputs(6540) <= (layer2_outputs(5966)) and not (layer2_outputs(4918));
    layer3_outputs(6541) <= (layer2_outputs(3079)) and (layer2_outputs(6857));
    layer3_outputs(6542) <= (layer2_outputs(4386)) and (layer2_outputs(3866));
    layer3_outputs(6543) <= not(layer2_outputs(3755));
    layer3_outputs(6544) <= not((layer2_outputs(2736)) and (layer2_outputs(5215)));
    layer3_outputs(6545) <= layer2_outputs(2951);
    layer3_outputs(6546) <= layer2_outputs(4532);
    layer3_outputs(6547) <= (layer2_outputs(10)) and not (layer2_outputs(2489));
    layer3_outputs(6548) <= not((layer2_outputs(2810)) or (layer2_outputs(2249)));
    layer3_outputs(6549) <= layer2_outputs(116);
    layer3_outputs(6550) <= '1';
    layer3_outputs(6551) <= not((layer2_outputs(2131)) or (layer2_outputs(2333)));
    layer3_outputs(6552) <= not((layer2_outputs(5669)) or (layer2_outputs(2277)));
    layer3_outputs(6553) <= '1';
    layer3_outputs(6554) <= '0';
    layer3_outputs(6555) <= '1';
    layer3_outputs(6556) <= not(layer2_outputs(6199)) or (layer2_outputs(2513));
    layer3_outputs(6557) <= (layer2_outputs(123)) or (layer2_outputs(5971));
    layer3_outputs(6558) <= (layer2_outputs(2183)) and not (layer2_outputs(5401));
    layer3_outputs(6559) <= not(layer2_outputs(9));
    layer3_outputs(6560) <= not((layer2_outputs(7018)) and (layer2_outputs(6503)));
    layer3_outputs(6561) <= layer2_outputs(3762);
    layer3_outputs(6562) <= (layer2_outputs(3682)) and not (layer2_outputs(2092));
    layer3_outputs(6563) <= not(layer2_outputs(2844)) or (layer2_outputs(2360));
    layer3_outputs(6564) <= (layer2_outputs(4842)) and (layer2_outputs(3935));
    layer3_outputs(6565) <= '0';
    layer3_outputs(6566) <= not(layer2_outputs(5521)) or (layer2_outputs(4841));
    layer3_outputs(6567) <= (layer2_outputs(5495)) and not (layer2_outputs(5227));
    layer3_outputs(6568) <= '0';
    layer3_outputs(6569) <= '1';
    layer3_outputs(6570) <= layer2_outputs(2777);
    layer3_outputs(6571) <= not(layer2_outputs(3254));
    layer3_outputs(6572) <= (layer2_outputs(5180)) and not (layer2_outputs(5281));
    layer3_outputs(6573) <= not(layer2_outputs(822));
    layer3_outputs(6574) <= not(layer2_outputs(3438)) or (layer2_outputs(6692));
    layer3_outputs(6575) <= not((layer2_outputs(7092)) and (layer2_outputs(1219)));
    layer3_outputs(6576) <= not(layer2_outputs(5183)) or (layer2_outputs(4308));
    layer3_outputs(6577) <= (layer2_outputs(4910)) or (layer2_outputs(7364));
    layer3_outputs(6578) <= not(layer2_outputs(2897));
    layer3_outputs(6579) <= layer2_outputs(1221);
    layer3_outputs(6580) <= not(layer2_outputs(1425));
    layer3_outputs(6581) <= layer2_outputs(1445);
    layer3_outputs(6582) <= not((layer2_outputs(6878)) or (layer2_outputs(2618)));
    layer3_outputs(6583) <= (layer2_outputs(6063)) and not (layer2_outputs(2814));
    layer3_outputs(6584) <= layer2_outputs(6283);
    layer3_outputs(6585) <= not(layer2_outputs(5233));
    layer3_outputs(6586) <= (layer2_outputs(4722)) xor (layer2_outputs(3315));
    layer3_outputs(6587) <= (layer2_outputs(4536)) and not (layer2_outputs(3890));
    layer3_outputs(6588) <= (layer2_outputs(1788)) and (layer2_outputs(2988));
    layer3_outputs(6589) <= not(layer2_outputs(6624));
    layer3_outputs(6590) <= '1';
    layer3_outputs(6591) <= not(layer2_outputs(6321));
    layer3_outputs(6592) <= '1';
    layer3_outputs(6593) <= (layer2_outputs(1881)) or (layer2_outputs(5559));
    layer3_outputs(6594) <= layer2_outputs(3496);
    layer3_outputs(6595) <= (layer2_outputs(421)) or (layer2_outputs(4651));
    layer3_outputs(6596) <= (layer2_outputs(3466)) or (layer2_outputs(1360));
    layer3_outputs(6597) <= not((layer2_outputs(6338)) or (layer2_outputs(248)));
    layer3_outputs(6598) <= (layer2_outputs(2785)) and not (layer2_outputs(5086));
    layer3_outputs(6599) <= (layer2_outputs(5516)) xor (layer2_outputs(6490));
    layer3_outputs(6600) <= not(layer2_outputs(6863)) or (layer2_outputs(60));
    layer3_outputs(6601) <= '0';
    layer3_outputs(6602) <= (layer2_outputs(2517)) and (layer2_outputs(3346));
    layer3_outputs(6603) <= not((layer2_outputs(6047)) and (layer2_outputs(2707)));
    layer3_outputs(6604) <= not((layer2_outputs(2213)) or (layer2_outputs(3125)));
    layer3_outputs(6605) <= '1';
    layer3_outputs(6606) <= not(layer2_outputs(2187));
    layer3_outputs(6607) <= not(layer2_outputs(1420));
    layer3_outputs(6608) <= (layer2_outputs(7398)) and (layer2_outputs(6304));
    layer3_outputs(6609) <= not(layer2_outputs(5969)) or (layer2_outputs(5576));
    layer3_outputs(6610) <= layer2_outputs(3357);
    layer3_outputs(6611) <= not(layer2_outputs(6642));
    layer3_outputs(6612) <= not(layer2_outputs(5832)) or (layer2_outputs(3041));
    layer3_outputs(6613) <= layer2_outputs(6581);
    layer3_outputs(6614) <= '0';
    layer3_outputs(6615) <= (layer2_outputs(4786)) and (layer2_outputs(857));
    layer3_outputs(6616) <= not(layer2_outputs(7155));
    layer3_outputs(6617) <= not(layer2_outputs(6018)) or (layer2_outputs(7315));
    layer3_outputs(6618) <= not(layer2_outputs(6732));
    layer3_outputs(6619) <= not(layer2_outputs(3005));
    layer3_outputs(6620) <= not(layer2_outputs(1593));
    layer3_outputs(6621) <= '0';
    layer3_outputs(6622) <= '1';
    layer3_outputs(6623) <= (layer2_outputs(5857)) and (layer2_outputs(5161));
    layer3_outputs(6624) <= not((layer2_outputs(5165)) and (layer2_outputs(5046)));
    layer3_outputs(6625) <= '0';
    layer3_outputs(6626) <= not(layer2_outputs(6734));
    layer3_outputs(6627) <= (layer2_outputs(2599)) and (layer2_outputs(2407));
    layer3_outputs(6628) <= (layer2_outputs(2800)) or (layer2_outputs(4781));
    layer3_outputs(6629) <= not((layer2_outputs(2051)) or (layer2_outputs(7266)));
    layer3_outputs(6630) <= layer2_outputs(5205);
    layer3_outputs(6631) <= (layer2_outputs(5882)) and not (layer2_outputs(43));
    layer3_outputs(6632) <= (layer2_outputs(3191)) and not (layer2_outputs(2200));
    layer3_outputs(6633) <= not((layer2_outputs(1263)) and (layer2_outputs(5923)));
    layer3_outputs(6634) <= layer2_outputs(4399);
    layer3_outputs(6635) <= layer2_outputs(87);
    layer3_outputs(6636) <= not((layer2_outputs(736)) and (layer2_outputs(519)));
    layer3_outputs(6637) <= (layer2_outputs(1965)) and (layer2_outputs(7186));
    layer3_outputs(6638) <= (layer2_outputs(2720)) and (layer2_outputs(47));
    layer3_outputs(6639) <= not(layer2_outputs(6773)) or (layer2_outputs(713));
    layer3_outputs(6640) <= (layer2_outputs(2312)) and not (layer2_outputs(800));
    layer3_outputs(6641) <= '0';
    layer3_outputs(6642) <= (layer2_outputs(1042)) and (layer2_outputs(7084));
    layer3_outputs(6643) <= not((layer2_outputs(3342)) or (layer2_outputs(3775)));
    layer3_outputs(6644) <= (layer2_outputs(6101)) or (layer2_outputs(5631));
    layer3_outputs(6645) <= not((layer2_outputs(3221)) or (layer2_outputs(2784)));
    layer3_outputs(6646) <= '1';
    layer3_outputs(6647) <= (layer2_outputs(820)) and not (layer2_outputs(4016));
    layer3_outputs(6648) <= not(layer2_outputs(1586));
    layer3_outputs(6649) <= (layer2_outputs(6749)) or (layer2_outputs(3433));
    layer3_outputs(6650) <= layer2_outputs(4631);
    layer3_outputs(6651) <= layer2_outputs(6531);
    layer3_outputs(6652) <= (layer2_outputs(3953)) and not (layer2_outputs(1064));
    layer3_outputs(6653) <= layer2_outputs(4988);
    layer3_outputs(6654) <= not(layer2_outputs(2526));
    layer3_outputs(6655) <= not(layer2_outputs(7258)) or (layer2_outputs(1160));
    layer3_outputs(6656) <= not(layer2_outputs(3594));
    layer3_outputs(6657) <= (layer2_outputs(3354)) and not (layer2_outputs(624));
    layer3_outputs(6658) <= not((layer2_outputs(5831)) or (layer2_outputs(308)));
    layer3_outputs(6659) <= (layer2_outputs(7037)) and not (layer2_outputs(4695));
    layer3_outputs(6660) <= '1';
    layer3_outputs(6661) <= layer2_outputs(1090);
    layer3_outputs(6662) <= not((layer2_outputs(6185)) and (layer2_outputs(3267)));
    layer3_outputs(6663) <= not((layer2_outputs(5762)) or (layer2_outputs(2799)));
    layer3_outputs(6664) <= not(layer2_outputs(5840));
    layer3_outputs(6665) <= layer2_outputs(3114);
    layer3_outputs(6666) <= layer2_outputs(3315);
    layer3_outputs(6667) <= not(layer2_outputs(3273));
    layer3_outputs(6668) <= not(layer2_outputs(970)) or (layer2_outputs(5966));
    layer3_outputs(6669) <= (layer2_outputs(5873)) or (layer2_outputs(2705));
    layer3_outputs(6670) <= (layer2_outputs(4825)) and (layer2_outputs(5686));
    layer3_outputs(6671) <= not(layer2_outputs(6050));
    layer3_outputs(6672) <= (layer2_outputs(2658)) and not (layer2_outputs(1677));
    layer3_outputs(6673) <= not(layer2_outputs(3874));
    layer3_outputs(6674) <= (layer2_outputs(1249)) and (layer2_outputs(5748));
    layer3_outputs(6675) <= not(layer2_outputs(6842));
    layer3_outputs(6676) <= not((layer2_outputs(3467)) and (layer2_outputs(3840)));
    layer3_outputs(6677) <= not(layer2_outputs(3631)) or (layer2_outputs(4278));
    layer3_outputs(6678) <= layer2_outputs(4227);
    layer3_outputs(6679) <= not(layer2_outputs(4025)) or (layer2_outputs(5753));
    layer3_outputs(6680) <= (layer2_outputs(230)) and (layer2_outputs(5817));
    layer3_outputs(6681) <= layer2_outputs(5659);
    layer3_outputs(6682) <= not(layer2_outputs(1035));
    layer3_outputs(6683) <= (layer2_outputs(6758)) xor (layer2_outputs(7613));
    layer3_outputs(6684) <= (layer2_outputs(5487)) and not (layer2_outputs(6692));
    layer3_outputs(6685) <= not(layer2_outputs(4970));
    layer3_outputs(6686) <= layer2_outputs(7085);
    layer3_outputs(6687) <= layer2_outputs(2843);
    layer3_outputs(6688) <= not(layer2_outputs(3274)) or (layer2_outputs(1517));
    layer3_outputs(6689) <= layer2_outputs(1582);
    layer3_outputs(6690) <= layer2_outputs(285);
    layer3_outputs(6691) <= not(layer2_outputs(700));
    layer3_outputs(6692) <= '1';
    layer3_outputs(6693) <= not(layer2_outputs(443));
    layer3_outputs(6694) <= (layer2_outputs(4115)) and not (layer2_outputs(4605));
    layer3_outputs(6695) <= '0';
    layer3_outputs(6696) <= (layer2_outputs(2408)) and not (layer2_outputs(5117));
    layer3_outputs(6697) <= (layer2_outputs(6594)) or (layer2_outputs(1522));
    layer3_outputs(6698) <= not(layer2_outputs(5177));
    layer3_outputs(6699) <= not(layer2_outputs(3414)) or (layer2_outputs(619));
    layer3_outputs(6700) <= layer2_outputs(3353);
    layer3_outputs(6701) <= (layer2_outputs(7034)) and (layer2_outputs(7046));
    layer3_outputs(6702) <= '1';
    layer3_outputs(6703) <= not(layer2_outputs(2803)) or (layer2_outputs(233));
    layer3_outputs(6704) <= layer2_outputs(86);
    layer3_outputs(6705) <= '1';
    layer3_outputs(6706) <= (layer2_outputs(2730)) and (layer2_outputs(4790));
    layer3_outputs(6707) <= not((layer2_outputs(773)) or (layer2_outputs(2048)));
    layer3_outputs(6708) <= layer2_outputs(6842);
    layer3_outputs(6709) <= not(layer2_outputs(4118));
    layer3_outputs(6710) <= not(layer2_outputs(4003));
    layer3_outputs(6711) <= '0';
    layer3_outputs(6712) <= (layer2_outputs(6540)) and (layer2_outputs(5585));
    layer3_outputs(6713) <= '0';
    layer3_outputs(6714) <= not(layer2_outputs(3868));
    layer3_outputs(6715) <= not((layer2_outputs(2743)) or (layer2_outputs(4786)));
    layer3_outputs(6716) <= layer2_outputs(4618);
    layer3_outputs(6717) <= '0';
    layer3_outputs(6718) <= not((layer2_outputs(2375)) or (layer2_outputs(2926)));
    layer3_outputs(6719) <= (layer2_outputs(5185)) or (layer2_outputs(7569));
    layer3_outputs(6720) <= layer2_outputs(5321);
    layer3_outputs(6721) <= '1';
    layer3_outputs(6722) <= not((layer2_outputs(6552)) or (layer2_outputs(2651)));
    layer3_outputs(6723) <= '0';
    layer3_outputs(6724) <= '0';
    layer3_outputs(6725) <= '1';
    layer3_outputs(6726) <= layer2_outputs(6698);
    layer3_outputs(6727) <= not(layer2_outputs(5772));
    layer3_outputs(6728) <= not(layer2_outputs(158));
    layer3_outputs(6729) <= '1';
    layer3_outputs(6730) <= not(layer2_outputs(2044));
    layer3_outputs(6731) <= layer2_outputs(5781);
    layer3_outputs(6732) <= layer2_outputs(6217);
    layer3_outputs(6733) <= layer2_outputs(1629);
    layer3_outputs(6734) <= not(layer2_outputs(6314)) or (layer2_outputs(3378));
    layer3_outputs(6735) <= not((layer2_outputs(1956)) or (layer2_outputs(4950)));
    layer3_outputs(6736) <= not(layer2_outputs(1512));
    layer3_outputs(6737) <= not(layer2_outputs(6941)) or (layer2_outputs(895));
    layer3_outputs(6738) <= not((layer2_outputs(4989)) and (layer2_outputs(6327)));
    layer3_outputs(6739) <= not(layer2_outputs(4029));
    layer3_outputs(6740) <= (layer2_outputs(1086)) and (layer2_outputs(4146));
    layer3_outputs(6741) <= not(layer2_outputs(1009)) or (layer2_outputs(2773));
    layer3_outputs(6742) <= not((layer2_outputs(5737)) and (layer2_outputs(2502)));
    layer3_outputs(6743) <= layer2_outputs(2285);
    layer3_outputs(6744) <= (layer2_outputs(252)) and not (layer2_outputs(3580));
    layer3_outputs(6745) <= (layer2_outputs(1734)) and not (layer2_outputs(2126));
    layer3_outputs(6746) <= layer2_outputs(7435);
    layer3_outputs(6747) <= layer2_outputs(6595);
    layer3_outputs(6748) <= '1';
    layer3_outputs(6749) <= not(layer2_outputs(981)) or (layer2_outputs(6023));
    layer3_outputs(6750) <= (layer2_outputs(1249)) or (layer2_outputs(6636));
    layer3_outputs(6751) <= (layer2_outputs(7499)) or (layer2_outputs(2833));
    layer3_outputs(6752) <= not((layer2_outputs(5784)) or (layer2_outputs(3831)));
    layer3_outputs(6753) <= not(layer2_outputs(380));
    layer3_outputs(6754) <= layer2_outputs(1279);
    layer3_outputs(6755) <= (layer2_outputs(3052)) and (layer2_outputs(674));
    layer3_outputs(6756) <= not(layer2_outputs(4348));
    layer3_outputs(6757) <= not(layer2_outputs(6403));
    layer3_outputs(6758) <= not((layer2_outputs(4848)) or (layer2_outputs(2006)));
    layer3_outputs(6759) <= (layer2_outputs(3306)) and not (layer2_outputs(7595));
    layer3_outputs(6760) <= (layer2_outputs(6954)) xor (layer2_outputs(2714));
    layer3_outputs(6761) <= not(layer2_outputs(2334));
    layer3_outputs(6762) <= not(layer2_outputs(6325));
    layer3_outputs(6763) <= (layer2_outputs(5428)) or (layer2_outputs(2613));
    layer3_outputs(6764) <= not((layer2_outputs(4181)) or (layer2_outputs(1935)));
    layer3_outputs(6765) <= layer2_outputs(7459);
    layer3_outputs(6766) <= (layer2_outputs(7147)) and not (layer2_outputs(3345));
    layer3_outputs(6767) <= not(layer2_outputs(461)) or (layer2_outputs(2584));
    layer3_outputs(6768) <= layer2_outputs(5832);
    layer3_outputs(6769) <= not(layer2_outputs(5449)) or (layer2_outputs(3736));
    layer3_outputs(6770) <= '0';
    layer3_outputs(6771) <= not((layer2_outputs(5495)) xor (layer2_outputs(7565)));
    layer3_outputs(6772) <= (layer2_outputs(4791)) and not (layer2_outputs(7329));
    layer3_outputs(6773) <= not((layer2_outputs(6511)) and (layer2_outputs(6472)));
    layer3_outputs(6774) <= layer2_outputs(4602);
    layer3_outputs(6775) <= '0';
    layer3_outputs(6776) <= layer2_outputs(7618);
    layer3_outputs(6777) <= not((layer2_outputs(4544)) and (layer2_outputs(5976)));
    layer3_outputs(6778) <= (layer2_outputs(7483)) or (layer2_outputs(3149));
    layer3_outputs(6779) <= '1';
    layer3_outputs(6780) <= layer2_outputs(2146);
    layer3_outputs(6781) <= layer2_outputs(5011);
    layer3_outputs(6782) <= not(layer2_outputs(1630));
    layer3_outputs(6783) <= layer2_outputs(2605);
    layer3_outputs(6784) <= (layer2_outputs(5729)) or (layer2_outputs(5578));
    layer3_outputs(6785) <= '0';
    layer3_outputs(6786) <= (layer2_outputs(6220)) and not (layer2_outputs(7217));
    layer3_outputs(6787) <= not((layer2_outputs(6998)) and (layer2_outputs(4701)));
    layer3_outputs(6788) <= not((layer2_outputs(6299)) and (layer2_outputs(4455)));
    layer3_outputs(6789) <= layer2_outputs(3800);
    layer3_outputs(6790) <= not((layer2_outputs(1798)) and (layer2_outputs(1756)));
    layer3_outputs(6791) <= not(layer2_outputs(4979)) or (layer2_outputs(1173));
    layer3_outputs(6792) <= layer2_outputs(5526);
    layer3_outputs(6793) <= not(layer2_outputs(6990));
    layer3_outputs(6794) <= not(layer2_outputs(3217));
    layer3_outputs(6795) <= not(layer2_outputs(7622));
    layer3_outputs(6796) <= '1';
    layer3_outputs(6797) <= '0';
    layer3_outputs(6798) <= not((layer2_outputs(709)) or (layer2_outputs(2592)));
    layer3_outputs(6799) <= not(layer2_outputs(1719));
    layer3_outputs(6800) <= (layer2_outputs(78)) or (layer2_outputs(3699));
    layer3_outputs(6801) <= (layer2_outputs(2214)) and not (layer2_outputs(711));
    layer3_outputs(6802) <= layer2_outputs(3100);
    layer3_outputs(6803) <= not(layer2_outputs(442)) or (layer2_outputs(762));
    layer3_outputs(6804) <= layer2_outputs(348);
    layer3_outputs(6805) <= not(layer2_outputs(355));
    layer3_outputs(6806) <= '0';
    layer3_outputs(6807) <= not(layer2_outputs(726));
    layer3_outputs(6808) <= '0';
    layer3_outputs(6809) <= not(layer2_outputs(488));
    layer3_outputs(6810) <= (layer2_outputs(3541)) xor (layer2_outputs(2134));
    layer3_outputs(6811) <= not(layer2_outputs(4855)) or (layer2_outputs(6382));
    layer3_outputs(6812) <= not(layer2_outputs(4564)) or (layer2_outputs(2895));
    layer3_outputs(6813) <= layer2_outputs(2081);
    layer3_outputs(6814) <= not(layer2_outputs(6229)) or (layer2_outputs(6901));
    layer3_outputs(6815) <= not((layer2_outputs(6660)) and (layer2_outputs(4838)));
    layer3_outputs(6816) <= (layer2_outputs(1148)) and not (layer2_outputs(7223));
    layer3_outputs(6817) <= '0';
    layer3_outputs(6818) <= (layer2_outputs(6085)) and (layer2_outputs(4189));
    layer3_outputs(6819) <= not(layer2_outputs(363)) or (layer2_outputs(6079));
    layer3_outputs(6820) <= not(layer2_outputs(3591));
    layer3_outputs(6821) <= layer2_outputs(2328);
    layer3_outputs(6822) <= not(layer2_outputs(1820)) or (layer2_outputs(411));
    layer3_outputs(6823) <= '1';
    layer3_outputs(6824) <= (layer2_outputs(1625)) and (layer2_outputs(2047));
    layer3_outputs(6825) <= layer2_outputs(2781);
    layer3_outputs(6826) <= (layer2_outputs(5606)) and not (layer2_outputs(6355));
    layer3_outputs(6827) <= layer2_outputs(6494);
    layer3_outputs(6828) <= not(layer2_outputs(623));
    layer3_outputs(6829) <= layer2_outputs(5886);
    layer3_outputs(6830) <= layer2_outputs(1859);
    layer3_outputs(6831) <= layer2_outputs(6867);
    layer3_outputs(6832) <= not((layer2_outputs(89)) xor (layer2_outputs(4338)));
    layer3_outputs(6833) <= not(layer2_outputs(5766));
    layer3_outputs(6834) <= (layer2_outputs(5927)) and not (layer2_outputs(6370));
    layer3_outputs(6835) <= not(layer2_outputs(2449));
    layer3_outputs(6836) <= not((layer2_outputs(3444)) and (layer2_outputs(5537)));
    layer3_outputs(6837) <= not(layer2_outputs(3086));
    layer3_outputs(6838) <= not(layer2_outputs(6713));
    layer3_outputs(6839) <= not((layer2_outputs(6104)) and (layer2_outputs(1444)));
    layer3_outputs(6840) <= not(layer2_outputs(1611));
    layer3_outputs(6841) <= not(layer2_outputs(362)) or (layer2_outputs(4546));
    layer3_outputs(6842) <= (layer2_outputs(1119)) and not (layer2_outputs(1610));
    layer3_outputs(6843) <= '0';
    layer3_outputs(6844) <= not(layer2_outputs(1875));
    layer3_outputs(6845) <= '0';
    layer3_outputs(6846) <= (layer2_outputs(7667)) and not (layer2_outputs(2821));
    layer3_outputs(6847) <= layer2_outputs(2186);
    layer3_outputs(6848) <= not(layer2_outputs(2978));
    layer3_outputs(6849) <= not((layer2_outputs(5070)) and (layer2_outputs(4712)));
    layer3_outputs(6850) <= (layer2_outputs(6841)) and not (layer2_outputs(6386));
    layer3_outputs(6851) <= not(layer2_outputs(427)) or (layer2_outputs(829));
    layer3_outputs(6852) <= not(layer2_outputs(6325));
    layer3_outputs(6853) <= '1';
    layer3_outputs(6854) <= layer2_outputs(6300);
    layer3_outputs(6855) <= (layer2_outputs(3978)) and not (layer2_outputs(4484));
    layer3_outputs(6856) <= layer2_outputs(6046);
    layer3_outputs(6857) <= not((layer2_outputs(497)) xor (layer2_outputs(5639)));
    layer3_outputs(6858) <= (layer2_outputs(3303)) and not (layer2_outputs(3992));
    layer3_outputs(6859) <= not(layer2_outputs(3813)) or (layer2_outputs(3920));
    layer3_outputs(6860) <= layer2_outputs(5959);
    layer3_outputs(6861) <= layer2_outputs(3648);
    layer3_outputs(6862) <= layer2_outputs(2839);
    layer3_outputs(6863) <= not(layer2_outputs(2597)) or (layer2_outputs(3450));
    layer3_outputs(6864) <= layer2_outputs(2246);
    layer3_outputs(6865) <= layer2_outputs(2831);
    layer3_outputs(6866) <= not((layer2_outputs(7612)) or (layer2_outputs(5544)));
    layer3_outputs(6867) <= not(layer2_outputs(4845)) or (layer2_outputs(6474));
    layer3_outputs(6868) <= not(layer2_outputs(3143)) or (layer2_outputs(3273));
    layer3_outputs(6869) <= (layer2_outputs(3526)) and not (layer2_outputs(4453));
    layer3_outputs(6870) <= (layer2_outputs(3784)) and not (layer2_outputs(1848));
    layer3_outputs(6871) <= not((layer2_outputs(5132)) or (layer2_outputs(7369)));
    layer3_outputs(6872) <= layer2_outputs(1730);
    layer3_outputs(6873) <= '0';
    layer3_outputs(6874) <= (layer2_outputs(5326)) xor (layer2_outputs(6242));
    layer3_outputs(6875) <= not(layer2_outputs(645));
    layer3_outputs(6876) <= layer2_outputs(2559);
    layer3_outputs(6877) <= layer2_outputs(695);
    layer3_outputs(6878) <= (layer2_outputs(2118)) and not (layer2_outputs(4171));
    layer3_outputs(6879) <= '0';
    layer3_outputs(6880) <= not(layer2_outputs(5139)) or (layer2_outputs(238));
    layer3_outputs(6881) <= not(layer2_outputs(4845));
    layer3_outputs(6882) <= (layer2_outputs(6122)) and not (layer2_outputs(7489));
    layer3_outputs(6883) <= (layer2_outputs(727)) and (layer2_outputs(6331));
    layer3_outputs(6884) <= not(layer2_outputs(2240));
    layer3_outputs(6885) <= not((layer2_outputs(1305)) xor (layer2_outputs(5027)));
    layer3_outputs(6886) <= not(layer2_outputs(6006));
    layer3_outputs(6887) <= (layer2_outputs(7474)) and not (layer2_outputs(5675));
    layer3_outputs(6888) <= not(layer2_outputs(5632));
    layer3_outputs(6889) <= (layer2_outputs(6981)) and not (layer2_outputs(1950));
    layer3_outputs(6890) <= layer2_outputs(4612);
    layer3_outputs(6891) <= not(layer2_outputs(2677));
    layer3_outputs(6892) <= not(layer2_outputs(530));
    layer3_outputs(6893) <= not(layer2_outputs(5918));
    layer3_outputs(6894) <= not(layer2_outputs(5077));
    layer3_outputs(6895) <= (layer2_outputs(6740)) and (layer2_outputs(7578));
    layer3_outputs(6896) <= not(layer2_outputs(3146));
    layer3_outputs(6897) <= (layer2_outputs(4214)) or (layer2_outputs(5422));
    layer3_outputs(6898) <= not(layer2_outputs(5301));
    layer3_outputs(6899) <= (layer2_outputs(7164)) and not (layer2_outputs(5156));
    layer3_outputs(6900) <= (layer2_outputs(3505)) and not (layer2_outputs(2877));
    layer3_outputs(6901) <= '0';
    layer3_outputs(6902) <= (layer2_outputs(3561)) and (layer2_outputs(1149));
    layer3_outputs(6903) <= layer2_outputs(6853);
    layer3_outputs(6904) <= not((layer2_outputs(3426)) and (layer2_outputs(6510)));
    layer3_outputs(6905) <= '0';
    layer3_outputs(6906) <= (layer2_outputs(4337)) and not (layer2_outputs(5344));
    layer3_outputs(6907) <= (layer2_outputs(697)) or (layer2_outputs(2097));
    layer3_outputs(6908) <= not((layer2_outputs(6856)) and (layer2_outputs(4255)));
    layer3_outputs(6909) <= layer2_outputs(1182);
    layer3_outputs(6910) <= layer2_outputs(6793);
    layer3_outputs(6911) <= layer2_outputs(6628);
    layer3_outputs(6912) <= (layer2_outputs(547)) and not (layer2_outputs(869));
    layer3_outputs(6913) <= not(layer2_outputs(1260)) or (layer2_outputs(5173));
    layer3_outputs(6914) <= not((layer2_outputs(1952)) and (layer2_outputs(2017)));
    layer3_outputs(6915) <= not(layer2_outputs(5863)) or (layer2_outputs(5097));
    layer3_outputs(6916) <= '0';
    layer3_outputs(6917) <= '0';
    layer3_outputs(6918) <= not(layer2_outputs(3024)) or (layer2_outputs(6679));
    layer3_outputs(6919) <= not((layer2_outputs(1754)) xor (layer2_outputs(2301)));
    layer3_outputs(6920) <= layer2_outputs(2719);
    layer3_outputs(6921) <= not((layer2_outputs(5957)) or (layer2_outputs(1211)));
    layer3_outputs(6922) <= not(layer2_outputs(7199));
    layer3_outputs(6923) <= not(layer2_outputs(931));
    layer3_outputs(6924) <= (layer2_outputs(4555)) or (layer2_outputs(3040));
    layer3_outputs(6925) <= layer2_outputs(3073);
    layer3_outputs(6926) <= not(layer2_outputs(4094));
    layer3_outputs(6927) <= '1';
    layer3_outputs(6928) <= not(layer2_outputs(2326)) or (layer2_outputs(4016));
    layer3_outputs(6929) <= not(layer2_outputs(3208)) or (layer2_outputs(386));
    layer3_outputs(6930) <= (layer2_outputs(2439)) or (layer2_outputs(7579));
    layer3_outputs(6931) <= (layer2_outputs(3409)) or (layer2_outputs(7309));
    layer3_outputs(6932) <= (layer2_outputs(4300)) and not (layer2_outputs(3457));
    layer3_outputs(6933) <= not((layer2_outputs(5230)) and (layer2_outputs(775)));
    layer3_outputs(6934) <= (layer2_outputs(1062)) or (layer2_outputs(6478));
    layer3_outputs(6935) <= layer2_outputs(1425);
    layer3_outputs(6936) <= not((layer2_outputs(1265)) and (layer2_outputs(746)));
    layer3_outputs(6937) <= (layer2_outputs(1679)) or (layer2_outputs(1448));
    layer3_outputs(6938) <= (layer2_outputs(499)) and (layer2_outputs(6353));
    layer3_outputs(6939) <= (layer2_outputs(2725)) and not (layer2_outputs(444));
    layer3_outputs(6940) <= (layer2_outputs(2422)) and not (layer2_outputs(7602));
    layer3_outputs(6941) <= not((layer2_outputs(6707)) and (layer2_outputs(4456)));
    layer3_outputs(6942) <= not(layer2_outputs(6902));
    layer3_outputs(6943) <= not(layer2_outputs(4488));
    layer3_outputs(6944) <= (layer2_outputs(1917)) or (layer2_outputs(3529));
    layer3_outputs(6945) <= not(layer2_outputs(2486)) or (layer2_outputs(3547));
    layer3_outputs(6946) <= '1';
    layer3_outputs(6947) <= '1';
    layer3_outputs(6948) <= not(layer2_outputs(1793)) or (layer2_outputs(6401));
    layer3_outputs(6949) <= layer2_outputs(1497);
    layer3_outputs(6950) <= not(layer2_outputs(466)) or (layer2_outputs(1492));
    layer3_outputs(6951) <= (layer2_outputs(3963)) xor (layer2_outputs(5680));
    layer3_outputs(6952) <= not(layer2_outputs(1670)) or (layer2_outputs(3239));
    layer3_outputs(6953) <= not(layer2_outputs(5996));
    layer3_outputs(6954) <= (layer2_outputs(6462)) xor (layer2_outputs(6081));
    layer3_outputs(6955) <= (layer2_outputs(4302)) or (layer2_outputs(6563));
    layer3_outputs(6956) <= '1';
    layer3_outputs(6957) <= not(layer2_outputs(5219));
    layer3_outputs(6958) <= layer2_outputs(1646);
    layer3_outputs(6959) <= (layer2_outputs(3566)) and not (layer2_outputs(611));
    layer3_outputs(6960) <= (layer2_outputs(3420)) and not (layer2_outputs(7447));
    layer3_outputs(6961) <= layer2_outputs(898);
    layer3_outputs(6962) <= not(layer2_outputs(864));
    layer3_outputs(6963) <= not((layer2_outputs(1239)) xor (layer2_outputs(6996)));
    layer3_outputs(6964) <= layer2_outputs(3480);
    layer3_outputs(6965) <= layer2_outputs(124);
    layer3_outputs(6966) <= layer2_outputs(7629);
    layer3_outputs(6967) <= not(layer2_outputs(7557));
    layer3_outputs(6968) <= not((layer2_outputs(6954)) and (layer2_outputs(4106)));
    layer3_outputs(6969) <= not((layer2_outputs(4777)) or (layer2_outputs(5587)));
    layer3_outputs(6970) <= not(layer2_outputs(4004));
    layer3_outputs(6971) <= (layer2_outputs(4971)) and (layer2_outputs(2657));
    layer3_outputs(6972) <= '1';
    layer3_outputs(6973) <= (layer2_outputs(2692)) and not (layer2_outputs(2242));
    layer3_outputs(6974) <= (layer2_outputs(4251)) and not (layer2_outputs(3212));
    layer3_outputs(6975) <= (layer2_outputs(7534)) or (layer2_outputs(1456));
    layer3_outputs(6976) <= (layer2_outputs(4588)) and not (layer2_outputs(5712));
    layer3_outputs(6977) <= not(layer2_outputs(1058));
    layer3_outputs(6978) <= layer2_outputs(6940);
    layer3_outputs(6979) <= (layer2_outputs(3494)) and not (layer2_outputs(7404));
    layer3_outputs(6980) <= '1';
    layer3_outputs(6981) <= layer2_outputs(549);
    layer3_outputs(6982) <= not(layer2_outputs(6809)) or (layer2_outputs(6343));
    layer3_outputs(6983) <= (layer2_outputs(6111)) and not (layer2_outputs(4165));
    layer3_outputs(6984) <= (layer2_outputs(3465)) or (layer2_outputs(7395));
    layer3_outputs(6985) <= '0';
    layer3_outputs(6986) <= '0';
    layer3_outputs(6987) <= layer2_outputs(2482);
    layer3_outputs(6988) <= layer2_outputs(3956);
    layer3_outputs(6989) <= layer2_outputs(940);
    layer3_outputs(6990) <= not(layer2_outputs(3861)) or (layer2_outputs(1703));
    layer3_outputs(6991) <= not(layer2_outputs(4241)) or (layer2_outputs(1680));
    layer3_outputs(6992) <= not((layer2_outputs(3286)) and (layer2_outputs(1137)));
    layer3_outputs(6993) <= not(layer2_outputs(5874)) or (layer2_outputs(2146));
    layer3_outputs(6994) <= '1';
    layer3_outputs(6995) <= layer2_outputs(3446);
    layer3_outputs(6996) <= not(layer2_outputs(1471)) or (layer2_outputs(2865));
    layer3_outputs(6997) <= not(layer2_outputs(6200)) or (layer2_outputs(5981));
    layer3_outputs(6998) <= not(layer2_outputs(6200));
    layer3_outputs(6999) <= not(layer2_outputs(600));
    layer3_outputs(7000) <= '0';
    layer3_outputs(7001) <= '1';
    layer3_outputs(7002) <= not((layer2_outputs(5174)) or (layer2_outputs(4713)));
    layer3_outputs(7003) <= layer2_outputs(4313);
    layer3_outputs(7004) <= (layer2_outputs(528)) and (layer2_outputs(3221));
    layer3_outputs(7005) <= not((layer2_outputs(6731)) or (layer2_outputs(94)));
    layer3_outputs(7006) <= not(layer2_outputs(7417)) or (layer2_outputs(2216));
    layer3_outputs(7007) <= not(layer2_outputs(4371));
    layer3_outputs(7008) <= not((layer2_outputs(4974)) or (layer2_outputs(879)));
    layer3_outputs(7009) <= not(layer2_outputs(2051)) or (layer2_outputs(762));
    layer3_outputs(7010) <= not(layer2_outputs(7012));
    layer3_outputs(7011) <= (layer2_outputs(4824)) and not (layer2_outputs(6517));
    layer3_outputs(7012) <= '1';
    layer3_outputs(7013) <= (layer2_outputs(5088)) and (layer2_outputs(4576));
    layer3_outputs(7014) <= (layer2_outputs(1858)) and (layer2_outputs(2577));
    layer3_outputs(7015) <= not((layer2_outputs(6367)) xor (layer2_outputs(345)));
    layer3_outputs(7016) <= not((layer2_outputs(4425)) or (layer2_outputs(1268)));
    layer3_outputs(7017) <= (layer2_outputs(3726)) and not (layer2_outputs(616));
    layer3_outputs(7018) <= layer2_outputs(3712);
    layer3_outputs(7019) <= not(layer2_outputs(214)) or (layer2_outputs(4792));
    layer3_outputs(7020) <= '0';
    layer3_outputs(7021) <= (layer2_outputs(2193)) and not (layer2_outputs(4123));
    layer3_outputs(7022) <= '1';
    layer3_outputs(7023) <= layer2_outputs(4967);
    layer3_outputs(7024) <= not(layer2_outputs(5927)) or (layer2_outputs(5037));
    layer3_outputs(7025) <= not((layer2_outputs(5956)) and (layer2_outputs(200)));
    layer3_outputs(7026) <= not(layer2_outputs(4164));
    layer3_outputs(7027) <= (layer2_outputs(6328)) xor (layer2_outputs(1629));
    layer3_outputs(7028) <= not(layer2_outputs(5711)) or (layer2_outputs(5101));
    layer3_outputs(7029) <= not((layer2_outputs(5427)) and (layer2_outputs(3989)));
    layer3_outputs(7030) <= '1';
    layer3_outputs(7031) <= not((layer2_outputs(3373)) or (layer2_outputs(5767)));
    layer3_outputs(7032) <= not((layer2_outputs(5605)) or (layer2_outputs(3282)));
    layer3_outputs(7033) <= layer2_outputs(3635);
    layer3_outputs(7034) <= not((layer2_outputs(7040)) and (layer2_outputs(1946)));
    layer3_outputs(7035) <= (layer2_outputs(2997)) xor (layer2_outputs(248));
    layer3_outputs(7036) <= not(layer2_outputs(3045)) or (layer2_outputs(3743));
    layer3_outputs(7037) <= not((layer2_outputs(3026)) and (layer2_outputs(7571)));
    layer3_outputs(7038) <= (layer2_outputs(6850)) and (layer2_outputs(275));
    layer3_outputs(7039) <= not(layer2_outputs(4298)) or (layer2_outputs(1993));
    layer3_outputs(7040) <= (layer2_outputs(4239)) and not (layer2_outputs(712));
    layer3_outputs(7041) <= layer2_outputs(7150);
    layer3_outputs(7042) <= '1';
    layer3_outputs(7043) <= not(layer2_outputs(970)) or (layer2_outputs(1619));
    layer3_outputs(7044) <= (layer2_outputs(4650)) or (layer2_outputs(1963));
    layer3_outputs(7045) <= (layer2_outputs(5826)) and not (layer2_outputs(7662));
    layer3_outputs(7046) <= '0';
    layer3_outputs(7047) <= not(layer2_outputs(7586));
    layer3_outputs(7048) <= layer2_outputs(4062);
    layer3_outputs(7049) <= not(layer2_outputs(1076));
    layer3_outputs(7050) <= (layer2_outputs(3473)) and (layer2_outputs(7414));
    layer3_outputs(7051) <= layer2_outputs(1969);
    layer3_outputs(7052) <= not(layer2_outputs(1488));
    layer3_outputs(7053) <= (layer2_outputs(1015)) and not (layer2_outputs(5973));
    layer3_outputs(7054) <= layer2_outputs(3796);
    layer3_outputs(7055) <= not(layer2_outputs(7175)) or (layer2_outputs(4295));
    layer3_outputs(7056) <= layer2_outputs(6915);
    layer3_outputs(7057) <= '1';
    layer3_outputs(7058) <= not(layer2_outputs(4467));
    layer3_outputs(7059) <= layer2_outputs(7256);
    layer3_outputs(7060) <= (layer2_outputs(2329)) and (layer2_outputs(5905));
    layer3_outputs(7061) <= layer2_outputs(3243);
    layer3_outputs(7062) <= not(layer2_outputs(2711)) or (layer2_outputs(6523));
    layer3_outputs(7063) <= not(layer2_outputs(5633));
    layer3_outputs(7064) <= layer2_outputs(6494);
    layer3_outputs(7065) <= layer2_outputs(1811);
    layer3_outputs(7066) <= (layer2_outputs(7314)) and not (layer2_outputs(3804));
    layer3_outputs(7067) <= layer2_outputs(7607);
    layer3_outputs(7068) <= not(layer2_outputs(4681));
    layer3_outputs(7069) <= (layer2_outputs(3696)) and (layer2_outputs(66));
    layer3_outputs(7070) <= not(layer2_outputs(3562));
    layer3_outputs(7071) <= not((layer2_outputs(3495)) or (layer2_outputs(2438)));
    layer3_outputs(7072) <= not((layer2_outputs(6813)) and (layer2_outputs(113)));
    layer3_outputs(7073) <= not((layer2_outputs(7254)) and (layer2_outputs(2142)));
    layer3_outputs(7074) <= layer2_outputs(1114);
    layer3_outputs(7075) <= (layer2_outputs(4348)) and (layer2_outputs(3888));
    layer3_outputs(7076) <= not(layer2_outputs(6341)) or (layer2_outputs(5568));
    layer3_outputs(7077) <= '1';
    layer3_outputs(7078) <= not(layer2_outputs(5536));
    layer3_outputs(7079) <= not(layer2_outputs(6972)) or (layer2_outputs(1374));
    layer3_outputs(7080) <= layer2_outputs(3546);
    layer3_outputs(7081) <= not(layer2_outputs(7675));
    layer3_outputs(7082) <= not((layer2_outputs(3071)) and (layer2_outputs(6193)));
    layer3_outputs(7083) <= '1';
    layer3_outputs(7084) <= (layer2_outputs(1316)) and not (layer2_outputs(6970));
    layer3_outputs(7085) <= not(layer2_outputs(143));
    layer3_outputs(7086) <= layer2_outputs(6259);
    layer3_outputs(7087) <= not((layer2_outputs(3213)) xor (layer2_outputs(1317)));
    layer3_outputs(7088) <= '1';
    layer3_outputs(7089) <= not(layer2_outputs(6427)) or (layer2_outputs(6490));
    layer3_outputs(7090) <= not(layer2_outputs(7226));
    layer3_outputs(7091) <= not(layer2_outputs(1932));
    layer3_outputs(7092) <= (layer2_outputs(4443)) and (layer2_outputs(2958));
    layer3_outputs(7093) <= not(layer2_outputs(5130));
    layer3_outputs(7094) <= (layer2_outputs(4792)) and (layer2_outputs(4168));
    layer3_outputs(7095) <= layer2_outputs(3830);
    layer3_outputs(7096) <= (layer2_outputs(4506)) and (layer2_outputs(5146));
    layer3_outputs(7097) <= '1';
    layer3_outputs(7098) <= '0';
    layer3_outputs(7099) <= not(layer2_outputs(5791));
    layer3_outputs(7100) <= not(layer2_outputs(7649));
    layer3_outputs(7101) <= layer2_outputs(2473);
    layer3_outputs(7102) <= not((layer2_outputs(7224)) or (layer2_outputs(4733)));
    layer3_outputs(7103) <= not((layer2_outputs(6155)) or (layer2_outputs(2465)));
    layer3_outputs(7104) <= layer2_outputs(1948);
    layer3_outputs(7105) <= layer2_outputs(2053);
    layer3_outputs(7106) <= not((layer2_outputs(2726)) or (layer2_outputs(4354)));
    layer3_outputs(7107) <= layer2_outputs(1243);
    layer3_outputs(7108) <= not(layer2_outputs(1473)) or (layer2_outputs(4558));
    layer3_outputs(7109) <= '1';
    layer3_outputs(7110) <= layer2_outputs(3196);
    layer3_outputs(7111) <= not((layer2_outputs(6723)) or (layer2_outputs(1847)));
    layer3_outputs(7112) <= not(layer2_outputs(4776));
    layer3_outputs(7113) <= '0';
    layer3_outputs(7114) <= layer2_outputs(4153);
    layer3_outputs(7115) <= '0';
    layer3_outputs(7116) <= layer2_outputs(4294);
    layer3_outputs(7117) <= (layer2_outputs(5895)) and not (layer2_outputs(97));
    layer3_outputs(7118) <= not(layer2_outputs(1634));
    layer3_outputs(7119) <= not(layer2_outputs(4350)) or (layer2_outputs(7603));
    layer3_outputs(7120) <= not((layer2_outputs(7271)) and (layer2_outputs(5705)));
    layer3_outputs(7121) <= not((layer2_outputs(6804)) xor (layer2_outputs(2449)));
    layer3_outputs(7122) <= layer2_outputs(3314);
    layer3_outputs(7123) <= layer2_outputs(99);
    layer3_outputs(7124) <= (layer2_outputs(5672)) and (layer2_outputs(1994));
    layer3_outputs(7125) <= not((layer2_outputs(4594)) and (layer2_outputs(4523)));
    layer3_outputs(7126) <= (layer2_outputs(573)) or (layer2_outputs(1925));
    layer3_outputs(7127) <= '1';
    layer3_outputs(7128) <= not((layer2_outputs(4943)) or (layer2_outputs(7354)));
    layer3_outputs(7129) <= layer2_outputs(1430);
    layer3_outputs(7130) <= (layer2_outputs(5892)) and not (layer2_outputs(6411));
    layer3_outputs(7131) <= '1';
    layer3_outputs(7132) <= not(layer2_outputs(4662)) or (layer2_outputs(3815));
    layer3_outputs(7133) <= (layer2_outputs(2184)) and not (layer2_outputs(2880));
    layer3_outputs(7134) <= not(layer2_outputs(1081)) or (layer2_outputs(2260));
    layer3_outputs(7135) <= layer2_outputs(5949);
    layer3_outputs(7136) <= not((layer2_outputs(5289)) and (layer2_outputs(2648)));
    layer3_outputs(7137) <= not(layer2_outputs(3035)) or (layer2_outputs(2297));
    layer3_outputs(7138) <= '0';
    layer3_outputs(7139) <= (layer2_outputs(3619)) or (layer2_outputs(5669));
    layer3_outputs(7140) <= '0';
    layer3_outputs(7141) <= not((layer2_outputs(226)) and (layer2_outputs(5997)));
    layer3_outputs(7142) <= not((layer2_outputs(6994)) or (layer2_outputs(4509)));
    layer3_outputs(7143) <= not(layer2_outputs(3308));
    layer3_outputs(7144) <= (layer2_outputs(5558)) and not (layer2_outputs(6364));
    layer3_outputs(7145) <= not((layer2_outputs(1190)) xor (layer2_outputs(1177)));
    layer3_outputs(7146) <= (layer2_outputs(5350)) and not (layer2_outputs(108));
    layer3_outputs(7147) <= not(layer2_outputs(2074));
    layer3_outputs(7148) <= (layer2_outputs(2545)) and not (layer2_outputs(5469));
    layer3_outputs(7149) <= '0';
    layer3_outputs(7150) <= not(layer2_outputs(3934)) or (layer2_outputs(5622));
    layer3_outputs(7151) <= (layer2_outputs(4930)) or (layer2_outputs(6964));
    layer3_outputs(7152) <= not(layer2_outputs(3425));
    layer3_outputs(7153) <= not(layer2_outputs(876)) or (layer2_outputs(5190));
    layer3_outputs(7154) <= not((layer2_outputs(1991)) or (layer2_outputs(1215)));
    layer3_outputs(7155) <= not(layer2_outputs(3652));
    layer3_outputs(7156) <= not((layer2_outputs(2255)) and (layer2_outputs(2983)));
    layer3_outputs(7157) <= not((layer2_outputs(3454)) and (layer2_outputs(3091)));
    layer3_outputs(7158) <= not(layer2_outputs(1561)) or (layer2_outputs(4604));
    layer3_outputs(7159) <= (layer2_outputs(242)) and (layer2_outputs(7063));
    layer3_outputs(7160) <= not(layer2_outputs(7460)) or (layer2_outputs(5935));
    layer3_outputs(7161) <= not(layer2_outputs(1479)) or (layer2_outputs(1821));
    layer3_outputs(7162) <= layer2_outputs(3161);
    layer3_outputs(7163) <= (layer2_outputs(109)) and (layer2_outputs(7352));
    layer3_outputs(7164) <= layer2_outputs(3706);
    layer3_outputs(7165) <= not(layer2_outputs(4489));
    layer3_outputs(7166) <= '0';
    layer3_outputs(7167) <= (layer2_outputs(2788)) xor (layer2_outputs(5752));
    layer3_outputs(7168) <= layer2_outputs(6504);
    layer3_outputs(7169) <= '0';
    layer3_outputs(7170) <= (layer2_outputs(1272)) or (layer2_outputs(5887));
    layer3_outputs(7171) <= not(layer2_outputs(3640));
    layer3_outputs(7172) <= not((layer2_outputs(808)) and (layer2_outputs(5642)));
    layer3_outputs(7173) <= not((layer2_outputs(3946)) and (layer2_outputs(2226)));
    layer3_outputs(7174) <= not(layer2_outputs(6851));
    layer3_outputs(7175) <= not(layer2_outputs(2256));
    layer3_outputs(7176) <= layer2_outputs(3522);
    layer3_outputs(7177) <= not(layer2_outputs(1783));
    layer3_outputs(7178) <= not((layer2_outputs(684)) or (layer2_outputs(7352)));
    layer3_outputs(7179) <= not(layer2_outputs(7509));
    layer3_outputs(7180) <= (layer2_outputs(5519)) and not (layer2_outputs(1838));
    layer3_outputs(7181) <= not((layer2_outputs(6979)) or (layer2_outputs(5789)));
    layer3_outputs(7182) <= (layer2_outputs(1584)) xor (layer2_outputs(242));
    layer3_outputs(7183) <= (layer2_outputs(4952)) and (layer2_outputs(5870));
    layer3_outputs(7184) <= layer2_outputs(167);
    layer3_outputs(7185) <= not(layer2_outputs(1067));
    layer3_outputs(7186) <= not((layer2_outputs(5131)) and (layer2_outputs(739)));
    layer3_outputs(7187) <= (layer2_outputs(253)) and (layer2_outputs(6952));
    layer3_outputs(7188) <= not((layer2_outputs(2351)) or (layer2_outputs(6470)));
    layer3_outputs(7189) <= (layer2_outputs(5949)) and (layer2_outputs(1681));
    layer3_outputs(7190) <= not(layer2_outputs(2915)) or (layer2_outputs(2923));
    layer3_outputs(7191) <= layer2_outputs(4852);
    layer3_outputs(7192) <= not(layer2_outputs(6005));
    layer3_outputs(7193) <= layer2_outputs(5324);
    layer3_outputs(7194) <= '0';
    layer3_outputs(7195) <= (layer2_outputs(3321)) xor (layer2_outputs(5611));
    layer3_outputs(7196) <= layer2_outputs(1740);
    layer3_outputs(7197) <= layer2_outputs(3147);
    layer3_outputs(7198) <= (layer2_outputs(6560)) and not (layer2_outputs(5904));
    layer3_outputs(7199) <= layer2_outputs(6942);
    layer3_outputs(7200) <= not(layer2_outputs(969));
    layer3_outputs(7201) <= not(layer2_outputs(2331));
    layer3_outputs(7202) <= layer2_outputs(871);
    layer3_outputs(7203) <= not(layer2_outputs(2198));
    layer3_outputs(7204) <= '1';
    layer3_outputs(7205) <= not((layer2_outputs(1299)) or (layer2_outputs(2653)));
    layer3_outputs(7206) <= not(layer2_outputs(2433));
    layer3_outputs(7207) <= (layer2_outputs(1331)) or (layer2_outputs(237));
    layer3_outputs(7208) <= not((layer2_outputs(2152)) and (layer2_outputs(4879)));
    layer3_outputs(7209) <= (layer2_outputs(157)) and not (layer2_outputs(7355));
    layer3_outputs(7210) <= (layer2_outputs(7630)) and not (layer2_outputs(1674));
    layer3_outputs(7211) <= layer2_outputs(1649);
    layer3_outputs(7212) <= (layer2_outputs(1325)) xor (layer2_outputs(5149));
    layer3_outputs(7213) <= layer2_outputs(1259);
    layer3_outputs(7214) <= layer2_outputs(2570);
    layer3_outputs(7215) <= '0';
    layer3_outputs(7216) <= not(layer2_outputs(1387));
    layer3_outputs(7217) <= not(layer2_outputs(2188));
    layer3_outputs(7218) <= layer2_outputs(4511);
    layer3_outputs(7219) <= not(layer2_outputs(294)) or (layer2_outputs(5056));
    layer3_outputs(7220) <= not(layer2_outputs(3065));
    layer3_outputs(7221) <= (layer2_outputs(57)) and (layer2_outputs(4722));
    layer3_outputs(7222) <= not((layer2_outputs(2384)) or (layer2_outputs(2473)));
    layer3_outputs(7223) <= not(layer2_outputs(3124));
    layer3_outputs(7224) <= '0';
    layer3_outputs(7225) <= not(layer2_outputs(3197)) or (layer2_outputs(4205));
    layer3_outputs(7226) <= layer2_outputs(3785);
    layer3_outputs(7227) <= not(layer2_outputs(7381));
    layer3_outputs(7228) <= not((layer2_outputs(6579)) and (layer2_outputs(3249)));
    layer3_outputs(7229) <= (layer2_outputs(529)) and not (layer2_outputs(2290));
    layer3_outputs(7230) <= not(layer2_outputs(4413));
    layer3_outputs(7231) <= (layer2_outputs(2028)) and not (layer2_outputs(677));
    layer3_outputs(7232) <= not(layer2_outputs(2306));
    layer3_outputs(7233) <= layer2_outputs(3698);
    layer3_outputs(7234) <= not(layer2_outputs(4511)) or (layer2_outputs(393));
    layer3_outputs(7235) <= not(layer2_outputs(6053));
    layer3_outputs(7236) <= (layer2_outputs(243)) and not (layer2_outputs(2333));
    layer3_outputs(7237) <= not(layer2_outputs(901)) or (layer2_outputs(6125));
    layer3_outputs(7238) <= not(layer2_outputs(6797)) or (layer2_outputs(2691));
    layer3_outputs(7239) <= layer2_outputs(4082);
    layer3_outputs(7240) <= not((layer2_outputs(1756)) xor (layer2_outputs(5398)));
    layer3_outputs(7241) <= (layer2_outputs(6536)) and (layer2_outputs(3219));
    layer3_outputs(7242) <= (layer2_outputs(2264)) and not (layer2_outputs(3572));
    layer3_outputs(7243) <= not(layer2_outputs(365)) or (layer2_outputs(731));
    layer3_outputs(7244) <= (layer2_outputs(6873)) and not (layer2_outputs(7526));
    layer3_outputs(7245) <= (layer2_outputs(7214)) and not (layer2_outputs(2423));
    layer3_outputs(7246) <= (layer2_outputs(794)) xor (layer2_outputs(7192));
    layer3_outputs(7247) <= not((layer2_outputs(1731)) and (layer2_outputs(7101)));
    layer3_outputs(7248) <= not(layer2_outputs(1159)) or (layer2_outputs(3105));
    layer3_outputs(7249) <= layer2_outputs(7157);
    layer3_outputs(7250) <= layer2_outputs(2351);
    layer3_outputs(7251) <= layer2_outputs(6711);
    layer3_outputs(7252) <= (layer2_outputs(6710)) and not (layer2_outputs(1366));
    layer3_outputs(7253) <= not((layer2_outputs(198)) or (layer2_outputs(7606)));
    layer3_outputs(7254) <= not(layer2_outputs(2751));
    layer3_outputs(7255) <= not(layer2_outputs(4850)) or (layer2_outputs(7596));
    layer3_outputs(7256) <= not(layer2_outputs(2917));
    layer3_outputs(7257) <= not(layer2_outputs(2852));
    layer3_outputs(7258) <= layer2_outputs(4577);
    layer3_outputs(7259) <= not((layer2_outputs(1319)) and (layer2_outputs(6237)));
    layer3_outputs(7260) <= not((layer2_outputs(7423)) and (layer2_outputs(2918)));
    layer3_outputs(7261) <= layer2_outputs(228);
    layer3_outputs(7262) <= layer2_outputs(1538);
    layer3_outputs(7263) <= (layer2_outputs(5360)) or (layer2_outputs(626));
    layer3_outputs(7264) <= (layer2_outputs(6499)) xor (layer2_outputs(5138));
    layer3_outputs(7265) <= layer2_outputs(5854);
    layer3_outputs(7266) <= layer2_outputs(1252);
    layer3_outputs(7267) <= not(layer2_outputs(3648));
    layer3_outputs(7268) <= not((layer2_outputs(7635)) or (layer2_outputs(1381)));
    layer3_outputs(7269) <= not(layer2_outputs(4049));
    layer3_outputs(7270) <= not((layer2_outputs(6673)) and (layer2_outputs(7556)));
    layer3_outputs(7271) <= not(layer2_outputs(3771));
    layer3_outputs(7272) <= not(layer2_outputs(7200));
    layer3_outputs(7273) <= not((layer2_outputs(3459)) xor (layer2_outputs(350)));
    layer3_outputs(7274) <= not((layer2_outputs(3722)) and (layer2_outputs(4435)));
    layer3_outputs(7275) <= (layer2_outputs(6695)) or (layer2_outputs(6703));
    layer3_outputs(7276) <= '0';
    layer3_outputs(7277) <= not(layer2_outputs(1045));
    layer3_outputs(7278) <= not(layer2_outputs(7384)) or (layer2_outputs(4057));
    layer3_outputs(7279) <= not((layer2_outputs(1478)) or (layer2_outputs(5182)));
    layer3_outputs(7280) <= '1';
    layer3_outputs(7281) <= (layer2_outputs(5092)) and (layer2_outputs(6576));
    layer3_outputs(7282) <= not(layer2_outputs(4856));
    layer3_outputs(7283) <= layer2_outputs(4352);
    layer3_outputs(7284) <= not((layer2_outputs(7242)) and (layer2_outputs(6460)));
    layer3_outputs(7285) <= not(layer2_outputs(2201)) or (layer2_outputs(6373));
    layer3_outputs(7286) <= (layer2_outputs(3401)) and not (layer2_outputs(6877));
    layer3_outputs(7287) <= not(layer2_outputs(2998)) or (layer2_outputs(6168));
    layer3_outputs(7288) <= not(layer2_outputs(545));
    layer3_outputs(7289) <= (layer2_outputs(483)) or (layer2_outputs(4018));
    layer3_outputs(7290) <= '0';
    layer3_outputs(7291) <= (layer2_outputs(5940)) and not (layer2_outputs(5205));
    layer3_outputs(7292) <= (layer2_outputs(2808)) or (layer2_outputs(4011));
    layer3_outputs(7293) <= not((layer2_outputs(5651)) and (layer2_outputs(3901)));
    layer3_outputs(7294) <= not(layer2_outputs(1747));
    layer3_outputs(7295) <= not(layer2_outputs(2883)) or (layer2_outputs(5140));
    layer3_outputs(7296) <= not(layer2_outputs(4474));
    layer3_outputs(7297) <= layer2_outputs(5743);
    layer3_outputs(7298) <= (layer2_outputs(5952)) or (layer2_outputs(7077));
    layer3_outputs(7299) <= not((layer2_outputs(5821)) or (layer2_outputs(2469)));
    layer3_outputs(7300) <= not((layer2_outputs(5351)) or (layer2_outputs(5852)));
    layer3_outputs(7301) <= (layer2_outputs(4646)) xor (layer2_outputs(6539));
    layer3_outputs(7302) <= '0';
    layer3_outputs(7303) <= layer2_outputs(733);
    layer3_outputs(7304) <= '1';
    layer3_outputs(7305) <= not(layer2_outputs(4014));
    layer3_outputs(7306) <= not(layer2_outputs(2350));
    layer3_outputs(7307) <= not(layer2_outputs(1667));
    layer3_outputs(7308) <= (layer2_outputs(2083)) and not (layer2_outputs(1981));
    layer3_outputs(7309) <= layer2_outputs(7529);
    layer3_outputs(7310) <= not(layer2_outputs(1169));
    layer3_outputs(7311) <= (layer2_outputs(6437)) xor (layer2_outputs(5402));
    layer3_outputs(7312) <= (layer2_outputs(4836)) and not (layer2_outputs(6044));
    layer3_outputs(7313) <= not(layer2_outputs(7512));
    layer3_outputs(7314) <= '0';
    layer3_outputs(7315) <= layer2_outputs(2533);
    layer3_outputs(7316) <= (layer2_outputs(5715)) and not (layer2_outputs(7074));
    layer3_outputs(7317) <= not((layer2_outputs(7415)) and (layer2_outputs(5889)));
    layer3_outputs(7318) <= (layer2_outputs(4987)) and not (layer2_outputs(2191));
    layer3_outputs(7319) <= (layer2_outputs(1704)) and (layer2_outputs(3793));
    layer3_outputs(7320) <= '1';
    layer3_outputs(7321) <= not(layer2_outputs(1085));
    layer3_outputs(7322) <= (layer2_outputs(5087)) and (layer2_outputs(7486));
    layer3_outputs(7323) <= not(layer2_outputs(5728));
    layer3_outputs(7324) <= layer2_outputs(2822);
    layer3_outputs(7325) <= (layer2_outputs(2079)) or (layer2_outputs(6028));
    layer3_outputs(7326) <= (layer2_outputs(5720)) or (layer2_outputs(2168));
    layer3_outputs(7327) <= not(layer2_outputs(3014));
    layer3_outputs(7328) <= layer2_outputs(3394);
    layer3_outputs(7329) <= layer2_outputs(892);
    layer3_outputs(7330) <= '1';
    layer3_outputs(7331) <= layer2_outputs(7592);
    layer3_outputs(7332) <= layer2_outputs(1471);
    layer3_outputs(7333) <= not(layer2_outputs(4803));
    layer3_outputs(7334) <= layer2_outputs(2621);
    layer3_outputs(7335) <= not(layer2_outputs(6844));
    layer3_outputs(7336) <= not(layer2_outputs(4533)) or (layer2_outputs(6407));
    layer3_outputs(7337) <= '1';
    layer3_outputs(7338) <= layer2_outputs(1481);
    layer3_outputs(7339) <= not(layer2_outputs(1823));
    layer3_outputs(7340) <= (layer2_outputs(4402)) and not (layer2_outputs(1740));
    layer3_outputs(7341) <= not((layer2_outputs(69)) and (layer2_outputs(67)));
    layer3_outputs(7342) <= layer2_outputs(7065);
    layer3_outputs(7343) <= not((layer2_outputs(3602)) and (layer2_outputs(3845)));
    layer3_outputs(7344) <= not(layer2_outputs(6046));
    layer3_outputs(7345) <= not(layer2_outputs(6733)) or (layer2_outputs(1652));
    layer3_outputs(7346) <= '1';
    layer3_outputs(7347) <= not((layer2_outputs(6781)) and (layer2_outputs(1444)));
    layer3_outputs(7348) <= not(layer2_outputs(1126));
    layer3_outputs(7349) <= not(layer2_outputs(2050));
    layer3_outputs(7350) <= not(layer2_outputs(5250));
    layer3_outputs(7351) <= not(layer2_outputs(793));
    layer3_outputs(7352) <= not((layer2_outputs(2516)) and (layer2_outputs(5835)));
    layer3_outputs(7353) <= not(layer2_outputs(6573));
    layer3_outputs(7354) <= not((layer2_outputs(6871)) and (layer2_outputs(3856)));
    layer3_outputs(7355) <= not((layer2_outputs(4898)) and (layer2_outputs(6859)));
    layer3_outputs(7356) <= not((layer2_outputs(1218)) and (layer2_outputs(5126)));
    layer3_outputs(7357) <= not(layer2_outputs(218));
    layer3_outputs(7358) <= (layer2_outputs(5487)) and not (layer2_outputs(4397));
    layer3_outputs(7359) <= layer2_outputs(832);
    layer3_outputs(7360) <= layer2_outputs(7332);
    layer3_outputs(7361) <= not((layer2_outputs(2142)) or (layer2_outputs(3032)));
    layer3_outputs(7362) <= layer2_outputs(885);
    layer3_outputs(7363) <= (layer2_outputs(6281)) and not (layer2_outputs(612));
    layer3_outputs(7364) <= layer2_outputs(1477);
    layer3_outputs(7365) <= not(layer2_outputs(7029));
    layer3_outputs(7366) <= not((layer2_outputs(4746)) and (layer2_outputs(757)));
    layer3_outputs(7367) <= (layer2_outputs(5298)) or (layer2_outputs(3770));
    layer3_outputs(7368) <= not(layer2_outputs(6987)) or (layer2_outputs(6699));
    layer3_outputs(7369) <= '1';
    layer3_outputs(7370) <= '0';
    layer3_outputs(7371) <= not((layer2_outputs(5305)) and (layer2_outputs(4164)));
    layer3_outputs(7372) <= layer2_outputs(1299);
    layer3_outputs(7373) <= not((layer2_outputs(4312)) xor (layer2_outputs(1446)));
    layer3_outputs(7374) <= (layer2_outputs(6209)) and not (layer2_outputs(1004));
    layer3_outputs(7375) <= not(layer2_outputs(1947)) or (layer2_outputs(7240));
    layer3_outputs(7376) <= not(layer2_outputs(3504));
    layer3_outputs(7377) <= layer2_outputs(4725);
    layer3_outputs(7378) <= not(layer2_outputs(1185)) or (layer2_outputs(4497));
    layer3_outputs(7379) <= (layer2_outputs(2717)) or (layer2_outputs(4596));
    layer3_outputs(7380) <= (layer2_outputs(3230)) and (layer2_outputs(4017));
    layer3_outputs(7381) <= '0';
    layer3_outputs(7382) <= not(layer2_outputs(765));
    layer3_outputs(7383) <= (layer2_outputs(6493)) and not (layer2_outputs(4206));
    layer3_outputs(7384) <= layer2_outputs(5836);
    layer3_outputs(7385) <= not(layer2_outputs(5657));
    layer3_outputs(7386) <= (layer2_outputs(3560)) and (layer2_outputs(4975));
    layer3_outputs(7387) <= '0';
    layer3_outputs(7388) <= not((layer2_outputs(5368)) or (layer2_outputs(4037)));
    layer3_outputs(7389) <= not((layer2_outputs(2647)) and (layer2_outputs(4015)));
    layer3_outputs(7390) <= not(layer2_outputs(6816));
    layer3_outputs(7391) <= '1';
    layer3_outputs(7392) <= not(layer2_outputs(3965));
    layer3_outputs(7393) <= '0';
    layer3_outputs(7394) <= layer2_outputs(2194);
    layer3_outputs(7395) <= (layer2_outputs(1350)) and not (layer2_outputs(4878));
    layer3_outputs(7396) <= not((layer2_outputs(6018)) xor (layer2_outputs(2930)));
    layer3_outputs(7397) <= layer2_outputs(2080);
    layer3_outputs(7398) <= (layer2_outputs(5754)) or (layer2_outputs(3400));
    layer3_outputs(7399) <= not(layer2_outputs(7167));
    layer3_outputs(7400) <= '1';
    layer3_outputs(7401) <= not(layer2_outputs(7657)) or (layer2_outputs(472));
    layer3_outputs(7402) <= (layer2_outputs(3466)) and not (layer2_outputs(5132));
    layer3_outputs(7403) <= (layer2_outputs(4766)) or (layer2_outputs(5410));
    layer3_outputs(7404) <= layer2_outputs(4024);
    layer3_outputs(7405) <= '0';
    layer3_outputs(7406) <= not(layer2_outputs(5014)) or (layer2_outputs(493));
    layer3_outputs(7407) <= not(layer2_outputs(626)) or (layer2_outputs(1219));
    layer3_outputs(7408) <= not(layer2_outputs(3792)) or (layer2_outputs(3630));
    layer3_outputs(7409) <= layer2_outputs(6017);
    layer3_outputs(7410) <= (layer2_outputs(3494)) and (layer2_outputs(3485));
    layer3_outputs(7411) <= not(layer2_outputs(5279));
    layer3_outputs(7412) <= not(layer2_outputs(5823));
    layer3_outputs(7413) <= layer2_outputs(4902);
    layer3_outputs(7414) <= layer2_outputs(7625);
    layer3_outputs(7415) <= not((layer2_outputs(1580)) or (layer2_outputs(5876)));
    layer3_outputs(7416) <= layer2_outputs(5300);
    layer3_outputs(7417) <= not(layer2_outputs(3169));
    layer3_outputs(7418) <= (layer2_outputs(5656)) or (layer2_outputs(591));
    layer3_outputs(7419) <= not(layer2_outputs(3429));
    layer3_outputs(7420) <= not(layer2_outputs(1081));
    layer3_outputs(7421) <= '0';
    layer3_outputs(7422) <= (layer2_outputs(3569)) and (layer2_outputs(4395));
    layer3_outputs(7423) <= not(layer2_outputs(1763)) or (layer2_outputs(1587));
    layer3_outputs(7424) <= '0';
    layer3_outputs(7425) <= (layer2_outputs(2088)) and (layer2_outputs(960));
    layer3_outputs(7426) <= '1';
    layer3_outputs(7427) <= not(layer2_outputs(101)) or (layer2_outputs(6575));
    layer3_outputs(7428) <= layer2_outputs(1460);
    layer3_outputs(7429) <= not((layer2_outputs(3309)) xor (layer2_outputs(6980)));
    layer3_outputs(7430) <= (layer2_outputs(5240)) or (layer2_outputs(4040));
    layer3_outputs(7431) <= not((layer2_outputs(3509)) and (layer2_outputs(2803)));
    layer3_outputs(7432) <= not(layer2_outputs(6171));
    layer3_outputs(7433) <= layer2_outputs(3598);
    layer3_outputs(7434) <= '0';
    layer3_outputs(7435) <= not(layer2_outputs(4489));
    layer3_outputs(7436) <= (layer2_outputs(7471)) or (layer2_outputs(1110));
    layer3_outputs(7437) <= '0';
    layer3_outputs(7438) <= layer2_outputs(3608);
    layer3_outputs(7439) <= (layer2_outputs(4990)) and not (layer2_outputs(463));
    layer3_outputs(7440) <= (layer2_outputs(7541)) and (layer2_outputs(1225));
    layer3_outputs(7441) <= layer2_outputs(4531);
    layer3_outputs(7442) <= not(layer2_outputs(4229));
    layer3_outputs(7443) <= layer2_outputs(3908);
    layer3_outputs(7444) <= not(layer2_outputs(6123)) or (layer2_outputs(1899));
    layer3_outputs(7445) <= layer2_outputs(631);
    layer3_outputs(7446) <= not(layer2_outputs(531)) or (layer2_outputs(5153));
    layer3_outputs(7447) <= not(layer2_outputs(516));
    layer3_outputs(7448) <= not(layer2_outputs(1019));
    layer3_outputs(7449) <= (layer2_outputs(7026)) and (layer2_outputs(6882));
    layer3_outputs(7450) <= not((layer2_outputs(1376)) and (layer2_outputs(5355)));
    layer3_outputs(7451) <= not((layer2_outputs(1961)) or (layer2_outputs(390)));
    layer3_outputs(7452) <= not(layer2_outputs(1051));
    layer3_outputs(7453) <= not(layer2_outputs(2842));
    layer3_outputs(7454) <= not(layer2_outputs(6141));
    layer3_outputs(7455) <= (layer2_outputs(4474)) and not (layer2_outputs(2061));
    layer3_outputs(7456) <= not(layer2_outputs(3374)) or (layer2_outputs(5771));
    layer3_outputs(7457) <= not(layer2_outputs(6409));
    layer3_outputs(7458) <= not(layer2_outputs(5897));
    layer3_outputs(7459) <= (layer2_outputs(2181)) and not (layer2_outputs(6109));
    layer3_outputs(7460) <= not((layer2_outputs(5213)) or (layer2_outputs(1634)));
    layer3_outputs(7461) <= not(layer2_outputs(6186));
    layer3_outputs(7462) <= not(layer2_outputs(4432)) or (layer2_outputs(4539));
    layer3_outputs(7463) <= layer2_outputs(5015);
    layer3_outputs(7464) <= not((layer2_outputs(3263)) and (layer2_outputs(2930)));
    layer3_outputs(7465) <= (layer2_outputs(6078)) and not (layer2_outputs(1180));
    layer3_outputs(7466) <= not((layer2_outputs(2205)) or (layer2_outputs(142)));
    layer3_outputs(7467) <= (layer2_outputs(3915)) or (layer2_outputs(5245));
    layer3_outputs(7468) <= '1';
    layer3_outputs(7469) <= (layer2_outputs(5183)) xor (layer2_outputs(1099));
    layer3_outputs(7470) <= (layer2_outputs(2869)) and not (layer2_outputs(276));
    layer3_outputs(7471) <= layer2_outputs(488);
    layer3_outputs(7472) <= '0';
    layer3_outputs(7473) <= layer2_outputs(6708);
    layer3_outputs(7474) <= not(layer2_outputs(5731));
    layer3_outputs(7475) <= layer2_outputs(4190);
    layer3_outputs(7476) <= layer2_outputs(3133);
    layer3_outputs(7477) <= (layer2_outputs(7548)) and (layer2_outputs(535));
    layer3_outputs(7478) <= not(layer2_outputs(393));
    layer3_outputs(7479) <= (layer2_outputs(1871)) or (layer2_outputs(7211));
    layer3_outputs(7480) <= (layer2_outputs(1680)) or (layer2_outputs(4433));
    layer3_outputs(7481) <= '0';
    layer3_outputs(7482) <= '1';
    layer3_outputs(7483) <= (layer2_outputs(6289)) or (layer2_outputs(2623));
    layer3_outputs(7484) <= not(layer2_outputs(2504));
    layer3_outputs(7485) <= '1';
    layer3_outputs(7486) <= not((layer2_outputs(3806)) or (layer2_outputs(7007)));
    layer3_outputs(7487) <= not((layer2_outputs(997)) and (layer2_outputs(326)));
    layer3_outputs(7488) <= not(layer2_outputs(2062));
    layer3_outputs(7489) <= not(layer2_outputs(5287));
    layer3_outputs(7490) <= (layer2_outputs(117)) and not (layer2_outputs(3140));
    layer3_outputs(7491) <= not(layer2_outputs(6333));
    layer3_outputs(7492) <= (layer2_outputs(4584)) and (layer2_outputs(6551));
    layer3_outputs(7493) <= not(layer2_outputs(5502));
    layer3_outputs(7494) <= '1';
    layer3_outputs(7495) <= not(layer2_outputs(5226)) or (layer2_outputs(7540));
    layer3_outputs(7496) <= layer2_outputs(1681);
    layer3_outputs(7497) <= (layer2_outputs(5588)) and not (layer2_outputs(850));
    layer3_outputs(7498) <= not(layer2_outputs(2291)) or (layer2_outputs(4916));
    layer3_outputs(7499) <= not((layer2_outputs(6812)) and (layer2_outputs(7642)));
    layer3_outputs(7500) <= (layer2_outputs(2421)) or (layer2_outputs(6831));
    layer3_outputs(7501) <= (layer2_outputs(3714)) or (layer2_outputs(1371));
    layer3_outputs(7502) <= '1';
    layer3_outputs(7503) <= not(layer2_outputs(2011)) or (layer2_outputs(2742));
    layer3_outputs(7504) <= not(layer2_outputs(358));
    layer3_outputs(7505) <= layer2_outputs(7478);
    layer3_outputs(7506) <= '1';
    layer3_outputs(7507) <= layer2_outputs(4718);
    layer3_outputs(7508) <= '0';
    layer3_outputs(7509) <= '0';
    layer3_outputs(7510) <= not(layer2_outputs(7088));
    layer3_outputs(7511) <= not(layer2_outputs(2022)) or (layer2_outputs(4942));
    layer3_outputs(7512) <= layer2_outputs(3728);
    layer3_outputs(7513) <= (layer2_outputs(5340)) and not (layer2_outputs(3533));
    layer3_outputs(7514) <= not(layer2_outputs(1278));
    layer3_outputs(7515) <= (layer2_outputs(2004)) or (layer2_outputs(3725));
    layer3_outputs(7516) <= not(layer2_outputs(3871)) or (layer2_outputs(949));
    layer3_outputs(7517) <= (layer2_outputs(2927)) and not (layer2_outputs(5929));
    layer3_outputs(7518) <= layer2_outputs(5715);
    layer3_outputs(7519) <= '1';
    layer3_outputs(7520) <= '0';
    layer3_outputs(7521) <= (layer2_outputs(2863)) and not (layer2_outputs(7562));
    layer3_outputs(7522) <= not(layer2_outputs(714)) or (layer2_outputs(5089));
    layer3_outputs(7523) <= not((layer2_outputs(2414)) and (layer2_outputs(5012)));
    layer3_outputs(7524) <= (layer2_outputs(7028)) and (layer2_outputs(6743));
    layer3_outputs(7525) <= (layer2_outputs(2791)) or (layer2_outputs(6725));
    layer3_outputs(7526) <= layer2_outputs(454);
    layer3_outputs(7527) <= not((layer2_outputs(3245)) and (layer2_outputs(7264)));
    layer3_outputs(7528) <= (layer2_outputs(5377)) and not (layer2_outputs(7343));
    layer3_outputs(7529) <= not((layer2_outputs(6334)) and (layer2_outputs(4708)));
    layer3_outputs(7530) <= not(layer2_outputs(827));
    layer3_outputs(7531) <= layer2_outputs(3279);
    layer3_outputs(7532) <= layer2_outputs(7376);
    layer3_outputs(7533) <= (layer2_outputs(5171)) and not (layer2_outputs(1518));
    layer3_outputs(7534) <= layer2_outputs(4378);
    layer3_outputs(7535) <= (layer2_outputs(7331)) and not (layer2_outputs(5595));
    layer3_outputs(7536) <= not(layer2_outputs(7372));
    layer3_outputs(7537) <= not(layer2_outputs(6680));
    layer3_outputs(7538) <= layer2_outputs(1697);
    layer3_outputs(7539) <= not((layer2_outputs(750)) xor (layer2_outputs(2818)));
    layer3_outputs(7540) <= not(layer2_outputs(4851));
    layer3_outputs(7541) <= not((layer2_outputs(6651)) and (layer2_outputs(6830)));
    layer3_outputs(7542) <= not((layer2_outputs(4418)) and (layer2_outputs(2124)));
    layer3_outputs(7543) <= (layer2_outputs(2475)) and not (layer2_outputs(3970));
    layer3_outputs(7544) <= layer2_outputs(4147);
    layer3_outputs(7545) <= not((layer2_outputs(2135)) xor (layer2_outputs(4184)));
    layer3_outputs(7546) <= not(layer2_outputs(1143));
    layer3_outputs(7547) <= (layer2_outputs(4121)) and not (layer2_outputs(3226));
    layer3_outputs(7548) <= (layer2_outputs(110)) and (layer2_outputs(1296));
    layer3_outputs(7549) <= layer2_outputs(3194);
    layer3_outputs(7550) <= layer2_outputs(7573);
    layer3_outputs(7551) <= '1';
    layer3_outputs(7552) <= not(layer2_outputs(2739));
    layer3_outputs(7553) <= layer2_outputs(2610);
    layer3_outputs(7554) <= (layer2_outputs(7346)) and not (layer2_outputs(2562));
    layer3_outputs(7555) <= not((layer2_outputs(3701)) and (layer2_outputs(4804)));
    layer3_outputs(7556) <= (layer2_outputs(4230)) xor (layer2_outputs(1000));
    layer3_outputs(7557) <= '0';
    layer3_outputs(7558) <= not(layer2_outputs(6628)) or (layer2_outputs(5436));
    layer3_outputs(7559) <= layer2_outputs(7621);
    layer3_outputs(7560) <= (layer2_outputs(3522)) and not (layer2_outputs(4122));
    layer3_outputs(7561) <= not(layer2_outputs(365)) or (layer2_outputs(779));
    layer3_outputs(7562) <= (layer2_outputs(6971)) or (layer2_outputs(7458));
    layer3_outputs(7563) <= (layer2_outputs(1220)) and (layer2_outputs(3178));
    layer3_outputs(7564) <= '1';
    layer3_outputs(7565) <= (layer2_outputs(1113)) and (layer2_outputs(7295));
    layer3_outputs(7566) <= (layer2_outputs(5330)) or (layer2_outputs(5869));
    layer3_outputs(7567) <= not(layer2_outputs(2832));
    layer3_outputs(7568) <= (layer2_outputs(4419)) and not (layer2_outputs(6617));
    layer3_outputs(7569) <= not((layer2_outputs(7175)) or (layer2_outputs(753)));
    layer3_outputs(7570) <= not(layer2_outputs(1029));
    layer3_outputs(7571) <= layer2_outputs(3872);
    layer3_outputs(7572) <= layer2_outputs(1788);
    layer3_outputs(7573) <= (layer2_outputs(1655)) and (layer2_outputs(1427));
    layer3_outputs(7574) <= not(layer2_outputs(975));
    layer3_outputs(7575) <= not(layer2_outputs(2353));
    layer3_outputs(7576) <= (layer2_outputs(2213)) and not (layer2_outputs(2366));
    layer3_outputs(7577) <= not((layer2_outputs(2780)) xor (layer2_outputs(4856)));
    layer3_outputs(7578) <= (layer2_outputs(4704)) and (layer2_outputs(5091));
    layer3_outputs(7579) <= not(layer2_outputs(3042)) or (layer2_outputs(4298));
    layer3_outputs(7580) <= (layer2_outputs(4512)) and not (layer2_outputs(270));
    layer3_outputs(7581) <= (layer2_outputs(1537)) and not (layer2_outputs(115));
    layer3_outputs(7582) <= not(layer2_outputs(2190));
    layer3_outputs(7583) <= '1';
    layer3_outputs(7584) <= '0';
    layer3_outputs(7585) <= layer2_outputs(3106);
    layer3_outputs(7586) <= not(layer2_outputs(2302));
    layer3_outputs(7587) <= layer2_outputs(2262);
    layer3_outputs(7588) <= (layer2_outputs(4329)) and not (layer2_outputs(759));
    layer3_outputs(7589) <= not((layer2_outputs(4643)) and (layer2_outputs(7173)));
    layer3_outputs(7590) <= not(layer2_outputs(6154)) or (layer2_outputs(465));
    layer3_outputs(7591) <= not((layer2_outputs(7568)) or (layer2_outputs(579)));
    layer3_outputs(7592) <= not(layer2_outputs(330)) or (layer2_outputs(7441));
    layer3_outputs(7593) <= not(layer2_outputs(4398));
    layer3_outputs(7594) <= not(layer2_outputs(1754));
    layer3_outputs(7595) <= layer2_outputs(3748);
    layer3_outputs(7596) <= not((layer2_outputs(2413)) and (layer2_outputs(4577)));
    layer3_outputs(7597) <= not(layer2_outputs(2454));
    layer3_outputs(7598) <= not(layer2_outputs(12));
    layer3_outputs(7599) <= (layer2_outputs(6221)) and not (layer2_outputs(4964));
    layer3_outputs(7600) <= not(layer2_outputs(5173)) or (layer2_outputs(3680));
    layer3_outputs(7601) <= layer2_outputs(404);
    layer3_outputs(7602) <= not(layer2_outputs(6604)) or (layer2_outputs(3034));
    layer3_outputs(7603) <= not((layer2_outputs(3220)) or (layer2_outputs(6619)));
    layer3_outputs(7604) <= (layer2_outputs(1445)) or (layer2_outputs(1632));
    layer3_outputs(7605) <= not(layer2_outputs(305)) or (layer2_outputs(497));
    layer3_outputs(7606) <= (layer2_outputs(3083)) and (layer2_outputs(1245));
    layer3_outputs(7607) <= (layer2_outputs(0)) and (layer2_outputs(976));
    layer3_outputs(7608) <= not((layer2_outputs(6580)) xor (layer2_outputs(168)));
    layer3_outputs(7609) <= not(layer2_outputs(6358));
    layer3_outputs(7610) <= '0';
    layer3_outputs(7611) <= '1';
    layer3_outputs(7612) <= '0';
    layer3_outputs(7613) <= (layer2_outputs(311)) xor (layer2_outputs(3425));
    layer3_outputs(7614) <= layer2_outputs(7176);
    layer3_outputs(7615) <= not((layer2_outputs(6443)) xor (layer2_outputs(4656)));
    layer3_outputs(7616) <= not((layer2_outputs(1136)) and (layer2_outputs(5264)));
    layer3_outputs(7617) <= layer2_outputs(3705);
    layer3_outputs(7618) <= (layer2_outputs(1014)) and not (layer2_outputs(4500));
    layer3_outputs(7619) <= (layer2_outputs(5309)) and (layer2_outputs(1562));
    layer3_outputs(7620) <= not(layer2_outputs(6896)) or (layer2_outputs(1091));
    layer3_outputs(7621) <= (layer2_outputs(3677)) and not (layer2_outputs(7477));
    layer3_outputs(7622) <= layer2_outputs(5814);
    layer3_outputs(7623) <= layer2_outputs(356);
    layer3_outputs(7624) <= layer2_outputs(4554);
    layer3_outputs(7625) <= (layer2_outputs(7094)) and not (layer2_outputs(5686));
    layer3_outputs(7626) <= '0';
    layer3_outputs(7627) <= (layer2_outputs(4812)) and (layer2_outputs(3685));
    layer3_outputs(7628) <= not((layer2_outputs(7674)) and (layer2_outputs(1097)));
    layer3_outputs(7629) <= not(layer2_outputs(4858)) or (layer2_outputs(2786));
    layer3_outputs(7630) <= '1';
    layer3_outputs(7631) <= layer2_outputs(7309);
    layer3_outputs(7632) <= (layer2_outputs(3951)) and not (layer2_outputs(4906));
    layer3_outputs(7633) <= not((layer2_outputs(7654)) or (layer2_outputs(841)));
    layer3_outputs(7634) <= not(layer2_outputs(1853));
    layer3_outputs(7635) <= not((layer2_outputs(810)) xor (layer2_outputs(3224)));
    layer3_outputs(7636) <= not(layer2_outputs(4839)) or (layer2_outputs(5251));
    layer3_outputs(7637) <= layer2_outputs(5234);
    layer3_outputs(7638) <= not(layer2_outputs(6098)) or (layer2_outputs(2968));
    layer3_outputs(7639) <= (layer2_outputs(4485)) and not (layer2_outputs(5503));
    layer3_outputs(7640) <= '0';
    layer3_outputs(7641) <= (layer2_outputs(5746)) and (layer2_outputs(5198));
    layer3_outputs(7642) <= layer2_outputs(225);
    layer3_outputs(7643) <= not(layer2_outputs(2842));
    layer3_outputs(7644) <= not(layer2_outputs(3237));
    layer3_outputs(7645) <= layer2_outputs(7031);
    layer3_outputs(7646) <= not(layer2_outputs(6328));
    layer3_outputs(7647) <= not(layer2_outputs(4328));
    layer3_outputs(7648) <= not((layer2_outputs(1743)) or (layer2_outputs(1919)));
    layer3_outputs(7649) <= not((layer2_outputs(7505)) xor (layer2_outputs(3148)));
    layer3_outputs(7650) <= layer2_outputs(1573);
    layer3_outputs(7651) <= not((layer2_outputs(1110)) xor (layer2_outputs(3142)));
    layer3_outputs(7652) <= not(layer2_outputs(6470)) or (layer2_outputs(3069));
    layer3_outputs(7653) <= not(layer2_outputs(6757));
    layer3_outputs(7654) <= (layer2_outputs(3715)) xor (layer2_outputs(104));
    layer3_outputs(7655) <= not(layer2_outputs(3997)) or (layer2_outputs(2211));
    layer3_outputs(7656) <= (layer2_outputs(5978)) and not (layer2_outputs(6286));
    layer3_outputs(7657) <= not(layer2_outputs(569));
    layer3_outputs(7658) <= not((layer2_outputs(134)) or (layer2_outputs(7079)));
    layer3_outputs(7659) <= layer2_outputs(1996);
    layer3_outputs(7660) <= (layer2_outputs(6931)) and not (layer2_outputs(4779));
    layer3_outputs(7661) <= layer2_outputs(3008);
    layer3_outputs(7662) <= not(layer2_outputs(2072));
    layer3_outputs(7663) <= layer2_outputs(1289);
    layer3_outputs(7664) <= (layer2_outputs(5006)) or (layer2_outputs(1407));
    layer3_outputs(7665) <= not(layer2_outputs(3404));
    layer3_outputs(7666) <= not(layer2_outputs(7334));
    layer3_outputs(7667) <= not(layer2_outputs(2916));
    layer3_outputs(7668) <= '0';
    layer3_outputs(7669) <= not(layer2_outputs(5861));
    layer3_outputs(7670) <= (layer2_outputs(399)) and (layer2_outputs(4922));
    layer3_outputs(7671) <= layer2_outputs(7069);
    layer3_outputs(7672) <= '1';
    layer3_outputs(7673) <= not((layer2_outputs(2910)) xor (layer2_outputs(266)));
    layer3_outputs(7674) <= (layer2_outputs(222)) xor (layer2_outputs(5169));
    layer3_outputs(7675) <= layer2_outputs(4222);
    layer3_outputs(7676) <= not(layer2_outputs(4208));
    layer3_outputs(7677) <= not(layer2_outputs(3158));
    layer3_outputs(7678) <= (layer2_outputs(2075)) and not (layer2_outputs(239));
    layer3_outputs(7679) <= (layer2_outputs(2858)) or (layer2_outputs(3658));
    layer4_outputs(0) <= layer3_outputs(2244);
    layer4_outputs(1) <= layer3_outputs(6995);
    layer4_outputs(2) <= not((layer3_outputs(1201)) and (layer3_outputs(1114)));
    layer4_outputs(3) <= layer3_outputs(1856);
    layer4_outputs(4) <= not(layer3_outputs(3473)) or (layer3_outputs(6109));
    layer4_outputs(5) <= layer3_outputs(5730);
    layer4_outputs(6) <= '1';
    layer4_outputs(7) <= layer3_outputs(7360);
    layer4_outputs(8) <= not(layer3_outputs(1504));
    layer4_outputs(9) <= layer3_outputs(1839);
    layer4_outputs(10) <= not((layer3_outputs(4967)) and (layer3_outputs(4376)));
    layer4_outputs(11) <= (layer3_outputs(7348)) xor (layer3_outputs(3109));
    layer4_outputs(12) <= (layer3_outputs(74)) and not (layer3_outputs(1130));
    layer4_outputs(13) <= layer3_outputs(4770);
    layer4_outputs(14) <= not((layer3_outputs(250)) xor (layer3_outputs(3221)));
    layer4_outputs(15) <= not((layer3_outputs(7419)) and (layer3_outputs(5082)));
    layer4_outputs(16) <= (layer3_outputs(5634)) xor (layer3_outputs(2901));
    layer4_outputs(17) <= (layer3_outputs(3936)) and (layer3_outputs(7116));
    layer4_outputs(18) <= layer3_outputs(3669);
    layer4_outputs(19) <= not((layer3_outputs(7488)) and (layer3_outputs(6270)));
    layer4_outputs(20) <= not(layer3_outputs(456));
    layer4_outputs(21) <= not(layer3_outputs(928));
    layer4_outputs(22) <= not(layer3_outputs(7053));
    layer4_outputs(23) <= layer3_outputs(871);
    layer4_outputs(24) <= not(layer3_outputs(568));
    layer4_outputs(25) <= not(layer3_outputs(6944));
    layer4_outputs(26) <= layer3_outputs(6812);
    layer4_outputs(27) <= (layer3_outputs(5868)) and not (layer3_outputs(7664));
    layer4_outputs(28) <= (layer3_outputs(247)) and (layer3_outputs(538));
    layer4_outputs(29) <= layer3_outputs(241);
    layer4_outputs(30) <= '1';
    layer4_outputs(31) <= layer3_outputs(3468);
    layer4_outputs(32) <= (layer3_outputs(5231)) and not (layer3_outputs(3644));
    layer4_outputs(33) <= not(layer3_outputs(2736));
    layer4_outputs(34) <= '0';
    layer4_outputs(35) <= '0';
    layer4_outputs(36) <= not((layer3_outputs(1741)) xor (layer3_outputs(2495)));
    layer4_outputs(37) <= not(layer3_outputs(5794));
    layer4_outputs(38) <= '0';
    layer4_outputs(39) <= not(layer3_outputs(4440));
    layer4_outputs(40) <= not(layer3_outputs(665));
    layer4_outputs(41) <= not(layer3_outputs(1355)) or (layer3_outputs(4352));
    layer4_outputs(42) <= not(layer3_outputs(1225));
    layer4_outputs(43) <= not((layer3_outputs(4427)) or (layer3_outputs(7546)));
    layer4_outputs(44) <= not((layer3_outputs(2193)) xor (layer3_outputs(4755)));
    layer4_outputs(45) <= not((layer3_outputs(403)) and (layer3_outputs(2045)));
    layer4_outputs(46) <= not((layer3_outputs(3192)) and (layer3_outputs(3185)));
    layer4_outputs(47) <= layer3_outputs(1958);
    layer4_outputs(48) <= '1';
    layer4_outputs(49) <= '1';
    layer4_outputs(50) <= not(layer3_outputs(5266));
    layer4_outputs(51) <= not(layer3_outputs(4393));
    layer4_outputs(52) <= not(layer3_outputs(2645));
    layer4_outputs(53) <= not(layer3_outputs(7573));
    layer4_outputs(54) <= not(layer3_outputs(2965));
    layer4_outputs(55) <= not((layer3_outputs(6523)) xor (layer3_outputs(2461)));
    layer4_outputs(56) <= not(layer3_outputs(785));
    layer4_outputs(57) <= '1';
    layer4_outputs(58) <= not(layer3_outputs(6737));
    layer4_outputs(59) <= (layer3_outputs(3110)) and (layer3_outputs(6067));
    layer4_outputs(60) <= layer3_outputs(5811);
    layer4_outputs(61) <= '1';
    layer4_outputs(62) <= (layer3_outputs(2900)) and not (layer3_outputs(3977));
    layer4_outputs(63) <= layer3_outputs(7355);
    layer4_outputs(64) <= (layer3_outputs(6243)) and (layer3_outputs(7067));
    layer4_outputs(65) <= not((layer3_outputs(784)) or (layer3_outputs(112)));
    layer4_outputs(66) <= not(layer3_outputs(700));
    layer4_outputs(67) <= not(layer3_outputs(6321));
    layer4_outputs(68) <= (layer3_outputs(4910)) or (layer3_outputs(1391));
    layer4_outputs(69) <= not(layer3_outputs(3674));
    layer4_outputs(70) <= not(layer3_outputs(669));
    layer4_outputs(71) <= '1';
    layer4_outputs(72) <= not(layer3_outputs(1561)) or (layer3_outputs(4794));
    layer4_outputs(73) <= not(layer3_outputs(2279)) or (layer3_outputs(7071));
    layer4_outputs(74) <= layer3_outputs(781);
    layer4_outputs(75) <= '0';
    layer4_outputs(76) <= (layer3_outputs(4424)) or (layer3_outputs(4334));
    layer4_outputs(77) <= not(layer3_outputs(4601)) or (layer3_outputs(174));
    layer4_outputs(78) <= not(layer3_outputs(7357)) or (layer3_outputs(3164));
    layer4_outputs(79) <= layer3_outputs(6411);
    layer4_outputs(80) <= not((layer3_outputs(49)) and (layer3_outputs(43)));
    layer4_outputs(81) <= not(layer3_outputs(1275)) or (layer3_outputs(6987));
    layer4_outputs(82) <= (layer3_outputs(3661)) and not (layer3_outputs(4990));
    layer4_outputs(83) <= not((layer3_outputs(6055)) or (layer3_outputs(6533)));
    layer4_outputs(84) <= not(layer3_outputs(1000));
    layer4_outputs(85) <= (layer3_outputs(4035)) and (layer3_outputs(4760));
    layer4_outputs(86) <= (layer3_outputs(3781)) and not (layer3_outputs(1667));
    layer4_outputs(87) <= not((layer3_outputs(92)) or (layer3_outputs(2622)));
    layer4_outputs(88) <= '0';
    layer4_outputs(89) <= layer3_outputs(1343);
    layer4_outputs(90) <= not((layer3_outputs(4058)) and (layer3_outputs(4031)));
    layer4_outputs(91) <= (layer3_outputs(2522)) and not (layer3_outputs(6049));
    layer4_outputs(92) <= not(layer3_outputs(300));
    layer4_outputs(93) <= not(layer3_outputs(2619));
    layer4_outputs(94) <= '1';
    layer4_outputs(95) <= layer3_outputs(5860);
    layer4_outputs(96) <= layer3_outputs(1218);
    layer4_outputs(97) <= (layer3_outputs(3264)) and not (layer3_outputs(6530));
    layer4_outputs(98) <= layer3_outputs(4649);
    layer4_outputs(99) <= layer3_outputs(4741);
    layer4_outputs(100) <= layer3_outputs(2920);
    layer4_outputs(101) <= not(layer3_outputs(6709));
    layer4_outputs(102) <= layer3_outputs(3828);
    layer4_outputs(103) <= not(layer3_outputs(6862));
    layer4_outputs(104) <= layer3_outputs(921);
    layer4_outputs(105) <= (layer3_outputs(2100)) or (layer3_outputs(4022));
    layer4_outputs(106) <= not(layer3_outputs(1684));
    layer4_outputs(107) <= not((layer3_outputs(4491)) xor (layer3_outputs(5818)));
    layer4_outputs(108) <= not(layer3_outputs(2546));
    layer4_outputs(109) <= '1';
    layer4_outputs(110) <= (layer3_outputs(6347)) xor (layer3_outputs(4387));
    layer4_outputs(111) <= (layer3_outputs(4609)) and not (layer3_outputs(5451));
    layer4_outputs(112) <= layer3_outputs(3436);
    layer4_outputs(113) <= layer3_outputs(3361);
    layer4_outputs(114) <= layer3_outputs(6490);
    layer4_outputs(115) <= not(layer3_outputs(1075));
    layer4_outputs(116) <= (layer3_outputs(7487)) and not (layer3_outputs(3468));
    layer4_outputs(117) <= (layer3_outputs(7229)) and (layer3_outputs(6710));
    layer4_outputs(118) <= layer3_outputs(5025);
    layer4_outputs(119) <= layer3_outputs(3496);
    layer4_outputs(120) <= not(layer3_outputs(4244));
    layer4_outputs(121) <= (layer3_outputs(4458)) and not (layer3_outputs(1523));
    layer4_outputs(122) <= layer3_outputs(2199);
    layer4_outputs(123) <= not((layer3_outputs(4196)) or (layer3_outputs(5114)));
    layer4_outputs(124) <= not(layer3_outputs(2794));
    layer4_outputs(125) <= layer3_outputs(6424);
    layer4_outputs(126) <= not((layer3_outputs(3139)) and (layer3_outputs(288)));
    layer4_outputs(127) <= not((layer3_outputs(1444)) and (layer3_outputs(4708)));
    layer4_outputs(128) <= not((layer3_outputs(5748)) and (layer3_outputs(680)));
    layer4_outputs(129) <= layer3_outputs(7089);
    layer4_outputs(130) <= layer3_outputs(382);
    layer4_outputs(131) <= (layer3_outputs(1550)) and not (layer3_outputs(4907));
    layer4_outputs(132) <= layer3_outputs(4790);
    layer4_outputs(133) <= not(layer3_outputs(2490)) or (layer3_outputs(2465));
    layer4_outputs(134) <= not(layer3_outputs(3907));
    layer4_outputs(135) <= not(layer3_outputs(502));
    layer4_outputs(136) <= (layer3_outputs(3381)) or (layer3_outputs(5554));
    layer4_outputs(137) <= (layer3_outputs(4317)) and not (layer3_outputs(7367));
    layer4_outputs(138) <= '1';
    layer4_outputs(139) <= (layer3_outputs(1514)) or (layer3_outputs(5910));
    layer4_outputs(140) <= (layer3_outputs(6518)) and not (layer3_outputs(4372));
    layer4_outputs(141) <= (layer3_outputs(2654)) and not (layer3_outputs(593));
    layer4_outputs(142) <= (layer3_outputs(6745)) and not (layer3_outputs(6458));
    layer4_outputs(143) <= not((layer3_outputs(320)) and (layer3_outputs(4632)));
    layer4_outputs(144) <= not(layer3_outputs(2925));
    layer4_outputs(145) <= not(layer3_outputs(1915)) or (layer3_outputs(7513));
    layer4_outputs(146) <= not(layer3_outputs(1305));
    layer4_outputs(147) <= layer3_outputs(4663);
    layer4_outputs(148) <= '1';
    layer4_outputs(149) <= not(layer3_outputs(309));
    layer4_outputs(150) <= not(layer3_outputs(2898));
    layer4_outputs(151) <= layer3_outputs(1260);
    layer4_outputs(152) <= layer3_outputs(1781);
    layer4_outputs(153) <= (layer3_outputs(6208)) and (layer3_outputs(2680));
    layer4_outputs(154) <= '1';
    layer4_outputs(155) <= not(layer3_outputs(4605)) or (layer3_outputs(7402));
    layer4_outputs(156) <= not((layer3_outputs(4690)) and (layer3_outputs(3721)));
    layer4_outputs(157) <= (layer3_outputs(4439)) and (layer3_outputs(6207));
    layer4_outputs(158) <= not(layer3_outputs(1990)) or (layer3_outputs(6387));
    layer4_outputs(159) <= not(layer3_outputs(4327));
    layer4_outputs(160) <= not(layer3_outputs(3290));
    layer4_outputs(161) <= not(layer3_outputs(2530));
    layer4_outputs(162) <= not(layer3_outputs(3996));
    layer4_outputs(163) <= not(layer3_outputs(459));
    layer4_outputs(164) <= (layer3_outputs(2512)) and (layer3_outputs(6818));
    layer4_outputs(165) <= not(layer3_outputs(4976));
    layer4_outputs(166) <= not((layer3_outputs(179)) or (layer3_outputs(5615)));
    layer4_outputs(167) <= not(layer3_outputs(3458));
    layer4_outputs(168) <= not(layer3_outputs(5909));
    layer4_outputs(169) <= layer3_outputs(6545);
    layer4_outputs(170) <= layer3_outputs(5550);
    layer4_outputs(171) <= (layer3_outputs(3575)) and not (layer3_outputs(4491));
    layer4_outputs(172) <= layer3_outputs(4533);
    layer4_outputs(173) <= not(layer3_outputs(1508));
    layer4_outputs(174) <= not(layer3_outputs(6066));
    layer4_outputs(175) <= layer3_outputs(5295);
    layer4_outputs(176) <= layer3_outputs(3066);
    layer4_outputs(177) <= '1';
    layer4_outputs(178) <= layer3_outputs(2122);
    layer4_outputs(179) <= layer3_outputs(5076);
    layer4_outputs(180) <= not(layer3_outputs(5647));
    layer4_outputs(181) <= not(layer3_outputs(6712)) or (layer3_outputs(3743));
    layer4_outputs(182) <= (layer3_outputs(5284)) xor (layer3_outputs(1382));
    layer4_outputs(183) <= not((layer3_outputs(2792)) or (layer3_outputs(4886)));
    layer4_outputs(184) <= not(layer3_outputs(2740));
    layer4_outputs(185) <= layer3_outputs(4131);
    layer4_outputs(186) <= '1';
    layer4_outputs(187) <= layer3_outputs(2377);
    layer4_outputs(188) <= not(layer3_outputs(1266));
    layer4_outputs(189) <= not(layer3_outputs(3503));
    layer4_outputs(190) <= layer3_outputs(6666);
    layer4_outputs(191) <= not((layer3_outputs(3441)) and (layer3_outputs(2170)));
    layer4_outputs(192) <= layer3_outputs(1102);
    layer4_outputs(193) <= layer3_outputs(4731);
    layer4_outputs(194) <= (layer3_outputs(602)) and not (layer3_outputs(3283));
    layer4_outputs(195) <= layer3_outputs(6154);
    layer4_outputs(196) <= layer3_outputs(3820);
    layer4_outputs(197) <= (layer3_outputs(4192)) and not (layer3_outputs(832));
    layer4_outputs(198) <= layer3_outputs(6749);
    layer4_outputs(199) <= (layer3_outputs(133)) and (layer3_outputs(5928));
    layer4_outputs(200) <= layer3_outputs(3226);
    layer4_outputs(201) <= (layer3_outputs(5622)) or (layer3_outputs(4396));
    layer4_outputs(202) <= not((layer3_outputs(3949)) and (layer3_outputs(3128)));
    layer4_outputs(203) <= (layer3_outputs(6316)) xor (layer3_outputs(4084));
    layer4_outputs(204) <= not(layer3_outputs(5210));
    layer4_outputs(205) <= (layer3_outputs(4015)) or (layer3_outputs(216));
    layer4_outputs(206) <= layer3_outputs(1045);
    layer4_outputs(207) <= layer3_outputs(5204);
    layer4_outputs(208) <= (layer3_outputs(4929)) and (layer3_outputs(5607));
    layer4_outputs(209) <= (layer3_outputs(1196)) and (layer3_outputs(6295));
    layer4_outputs(210) <= (layer3_outputs(1358)) and not (layer3_outputs(1381));
    layer4_outputs(211) <= layer3_outputs(7482);
    layer4_outputs(212) <= layer3_outputs(6760);
    layer4_outputs(213) <= layer3_outputs(2861);
    layer4_outputs(214) <= not((layer3_outputs(5038)) or (layer3_outputs(4721)));
    layer4_outputs(215) <= not(layer3_outputs(5027));
    layer4_outputs(216) <= layer3_outputs(900);
    layer4_outputs(217) <= layer3_outputs(2940);
    layer4_outputs(218) <= not(layer3_outputs(639));
    layer4_outputs(219) <= layer3_outputs(2405);
    layer4_outputs(220) <= not(layer3_outputs(7337));
    layer4_outputs(221) <= not(layer3_outputs(2292));
    layer4_outputs(222) <= not((layer3_outputs(1937)) xor (layer3_outputs(2455)));
    layer4_outputs(223) <= not((layer3_outputs(917)) or (layer3_outputs(4496)));
    layer4_outputs(224) <= not(layer3_outputs(6859)) or (layer3_outputs(1194));
    layer4_outputs(225) <= not(layer3_outputs(7459));
    layer4_outputs(226) <= (layer3_outputs(2284)) xor (layer3_outputs(2872));
    layer4_outputs(227) <= (layer3_outputs(3681)) and not (layer3_outputs(4855));
    layer4_outputs(228) <= layer3_outputs(5157);
    layer4_outputs(229) <= not((layer3_outputs(3490)) xor (layer3_outputs(7031)));
    layer4_outputs(230) <= not(layer3_outputs(2663));
    layer4_outputs(231) <= not(layer3_outputs(4019));
    layer4_outputs(232) <= '0';
    layer4_outputs(233) <= layer3_outputs(6833);
    layer4_outputs(234) <= layer3_outputs(1273);
    layer4_outputs(235) <= layer3_outputs(7475);
    layer4_outputs(236) <= not((layer3_outputs(2762)) xor (layer3_outputs(6703)));
    layer4_outputs(237) <= not(layer3_outputs(5929));
    layer4_outputs(238) <= not(layer3_outputs(4569)) or (layer3_outputs(4681));
    layer4_outputs(239) <= not(layer3_outputs(461));
    layer4_outputs(240) <= (layer3_outputs(4868)) and (layer3_outputs(6169));
    layer4_outputs(241) <= layer3_outputs(2428);
    layer4_outputs(242) <= (layer3_outputs(358)) or (layer3_outputs(7514));
    layer4_outputs(243) <= not(layer3_outputs(1361));
    layer4_outputs(244) <= not((layer3_outputs(7195)) xor (layer3_outputs(4038)));
    layer4_outputs(245) <= layer3_outputs(2842);
    layer4_outputs(246) <= not((layer3_outputs(2417)) or (layer3_outputs(4551)));
    layer4_outputs(247) <= layer3_outputs(2833);
    layer4_outputs(248) <= not((layer3_outputs(4341)) or (layer3_outputs(2888)));
    layer4_outputs(249) <= (layer3_outputs(477)) xor (layer3_outputs(5146));
    layer4_outputs(250) <= layer3_outputs(2958);
    layer4_outputs(251) <= layer3_outputs(1524);
    layer4_outputs(252) <= not(layer3_outputs(3176));
    layer4_outputs(253) <= not(layer3_outputs(5218)) or (layer3_outputs(1202));
    layer4_outputs(254) <= not(layer3_outputs(6618));
    layer4_outputs(255) <= not(layer3_outputs(5149)) or (layer3_outputs(1896));
    layer4_outputs(256) <= (layer3_outputs(6210)) and not (layer3_outputs(3086));
    layer4_outputs(257) <= (layer3_outputs(6763)) and (layer3_outputs(4407));
    layer4_outputs(258) <= not((layer3_outputs(2130)) xor (layer3_outputs(277)));
    layer4_outputs(259) <= layer3_outputs(3842);
    layer4_outputs(260) <= '1';
    layer4_outputs(261) <= (layer3_outputs(3443)) and not (layer3_outputs(1957));
    layer4_outputs(262) <= not(layer3_outputs(973));
    layer4_outputs(263) <= not((layer3_outputs(5368)) xor (layer3_outputs(1444)));
    layer4_outputs(264) <= layer3_outputs(5887);
    layer4_outputs(265) <= not(layer3_outputs(6761));
    layer4_outputs(266) <= not(layer3_outputs(6116));
    layer4_outputs(267) <= layer3_outputs(4581);
    layer4_outputs(268) <= layer3_outputs(7440);
    layer4_outputs(269) <= '1';
    layer4_outputs(270) <= not(layer3_outputs(3713));
    layer4_outputs(271) <= (layer3_outputs(6123)) or (layer3_outputs(4428));
    layer4_outputs(272) <= not((layer3_outputs(6476)) xor (layer3_outputs(7564)));
    layer4_outputs(273) <= not((layer3_outputs(3497)) or (layer3_outputs(5531)));
    layer4_outputs(274) <= (layer3_outputs(3505)) and not (layer3_outputs(6441));
    layer4_outputs(275) <= layer3_outputs(7603);
    layer4_outputs(276) <= (layer3_outputs(1457)) xor (layer3_outputs(1242));
    layer4_outputs(277) <= not(layer3_outputs(7306)) or (layer3_outputs(4926));
    layer4_outputs(278) <= not(layer3_outputs(3738)) or (layer3_outputs(252));
    layer4_outputs(279) <= not((layer3_outputs(810)) or (layer3_outputs(366)));
    layer4_outputs(280) <= layer3_outputs(3658);
    layer4_outputs(281) <= (layer3_outputs(4016)) xor (layer3_outputs(3843));
    layer4_outputs(282) <= not(layer3_outputs(4782));
    layer4_outputs(283) <= not(layer3_outputs(1148));
    layer4_outputs(284) <= not(layer3_outputs(7514));
    layer4_outputs(285) <= not(layer3_outputs(5788)) or (layer3_outputs(6885));
    layer4_outputs(286) <= not((layer3_outputs(400)) or (layer3_outputs(4821)));
    layer4_outputs(287) <= not(layer3_outputs(2846));
    layer4_outputs(288) <= not((layer3_outputs(3131)) and (layer3_outputs(1766)));
    layer4_outputs(289) <= not(layer3_outputs(4054)) or (layer3_outputs(4251));
    layer4_outputs(290) <= not(layer3_outputs(4767)) or (layer3_outputs(41));
    layer4_outputs(291) <= not(layer3_outputs(4258));
    layer4_outputs(292) <= not(layer3_outputs(6386)) or (layer3_outputs(3138));
    layer4_outputs(293) <= not(layer3_outputs(3674));
    layer4_outputs(294) <= layer3_outputs(3027);
    layer4_outputs(295) <= not((layer3_outputs(2040)) or (layer3_outputs(3770)));
    layer4_outputs(296) <= '0';
    layer4_outputs(297) <= (layer3_outputs(1524)) and not (layer3_outputs(1296));
    layer4_outputs(298) <= (layer3_outputs(2801)) and (layer3_outputs(6915));
    layer4_outputs(299) <= (layer3_outputs(4988)) xor (layer3_outputs(3285));
    layer4_outputs(300) <= not((layer3_outputs(120)) and (layer3_outputs(1386)));
    layer4_outputs(301) <= not(layer3_outputs(361));
    layer4_outputs(302) <= not(layer3_outputs(5350)) or (layer3_outputs(1357));
    layer4_outputs(303) <= layer3_outputs(536);
    layer4_outputs(304) <= not(layer3_outputs(4159));
    layer4_outputs(305) <= not(layer3_outputs(6303));
    layer4_outputs(306) <= not(layer3_outputs(3729));
    layer4_outputs(307) <= not(layer3_outputs(1994)) or (layer3_outputs(998));
    layer4_outputs(308) <= not((layer3_outputs(5845)) xor (layer3_outputs(5424)));
    layer4_outputs(309) <= not(layer3_outputs(1958));
    layer4_outputs(310) <= not(layer3_outputs(3781)) or (layer3_outputs(1892));
    layer4_outputs(311) <= not(layer3_outputs(4729));
    layer4_outputs(312) <= (layer3_outputs(3939)) or (layer3_outputs(7563));
    layer4_outputs(313) <= (layer3_outputs(5072)) and not (layer3_outputs(1816));
    layer4_outputs(314) <= not((layer3_outputs(6413)) xor (layer3_outputs(3082)));
    layer4_outputs(315) <= layer3_outputs(7098);
    layer4_outputs(316) <= not(layer3_outputs(6360)) or (layer3_outputs(3501));
    layer4_outputs(317) <= not(layer3_outputs(3515));
    layer4_outputs(318) <= not(layer3_outputs(741));
    layer4_outputs(319) <= layer3_outputs(346);
    layer4_outputs(320) <= '0';
    layer4_outputs(321) <= (layer3_outputs(6108)) and (layer3_outputs(482));
    layer4_outputs(322) <= not((layer3_outputs(4708)) or (layer3_outputs(291)));
    layer4_outputs(323) <= not(layer3_outputs(1962));
    layer4_outputs(324) <= (layer3_outputs(3327)) or (layer3_outputs(2669));
    layer4_outputs(325) <= '0';
    layer4_outputs(326) <= (layer3_outputs(4976)) and not (layer3_outputs(7659));
    layer4_outputs(327) <= not(layer3_outputs(5543)) or (layer3_outputs(1883));
    layer4_outputs(328) <= not(layer3_outputs(5449));
    layer4_outputs(329) <= (layer3_outputs(5175)) and not (layer3_outputs(1276));
    layer4_outputs(330) <= layer3_outputs(3784);
    layer4_outputs(331) <= (layer3_outputs(7087)) or (layer3_outputs(1675));
    layer4_outputs(332) <= layer3_outputs(428);
    layer4_outputs(333) <= not((layer3_outputs(74)) xor (layer3_outputs(1216)));
    layer4_outputs(334) <= not(layer3_outputs(5712));
    layer4_outputs(335) <= not(layer3_outputs(5161));
    layer4_outputs(336) <= (layer3_outputs(5627)) or (layer3_outputs(4616));
    layer4_outputs(337) <= (layer3_outputs(5648)) or (layer3_outputs(6882));
    layer4_outputs(338) <= '0';
    layer4_outputs(339) <= layer3_outputs(6287);
    layer4_outputs(340) <= not(layer3_outputs(7569));
    layer4_outputs(341) <= layer3_outputs(1604);
    layer4_outputs(342) <= (layer3_outputs(7408)) and (layer3_outputs(1259));
    layer4_outputs(343) <= not(layer3_outputs(3854));
    layer4_outputs(344) <= '1';
    layer4_outputs(345) <= layer3_outputs(3936);
    layer4_outputs(346) <= layer3_outputs(2554);
    layer4_outputs(347) <= layer3_outputs(7536);
    layer4_outputs(348) <= not((layer3_outputs(5148)) or (layer3_outputs(689)));
    layer4_outputs(349) <= not((layer3_outputs(7279)) and (layer3_outputs(5129)));
    layer4_outputs(350) <= '1';
    layer4_outputs(351) <= not(layer3_outputs(3476));
    layer4_outputs(352) <= layer3_outputs(4451);
    layer4_outputs(353) <= not(layer3_outputs(2341));
    layer4_outputs(354) <= '1';
    layer4_outputs(355) <= (layer3_outputs(5381)) or (layer3_outputs(4797));
    layer4_outputs(356) <= (layer3_outputs(7673)) and not (layer3_outputs(5935));
    layer4_outputs(357) <= (layer3_outputs(2431)) and (layer3_outputs(72));
    layer4_outputs(358) <= not(layer3_outputs(624));
    layer4_outputs(359) <= layer3_outputs(1002);
    layer4_outputs(360) <= not(layer3_outputs(6033));
    layer4_outputs(361) <= layer3_outputs(4261);
    layer4_outputs(362) <= (layer3_outputs(6888)) and not (layer3_outputs(2950));
    layer4_outputs(363) <= layer3_outputs(4746);
    layer4_outputs(364) <= not(layer3_outputs(5519));
    layer4_outputs(365) <= not(layer3_outputs(7202)) or (layer3_outputs(2927));
    layer4_outputs(366) <= not((layer3_outputs(4220)) xor (layer3_outputs(409)));
    layer4_outputs(367) <= '1';
    layer4_outputs(368) <= not(layer3_outputs(5216));
    layer4_outputs(369) <= (layer3_outputs(4433)) and (layer3_outputs(4824));
    layer4_outputs(370) <= '1';
    layer4_outputs(371) <= not(layer3_outputs(3300));
    layer4_outputs(372) <= layer3_outputs(1132);
    layer4_outputs(373) <= layer3_outputs(7004);
    layer4_outputs(374) <= not(layer3_outputs(1729)) or (layer3_outputs(3859));
    layer4_outputs(375) <= layer3_outputs(1826);
    layer4_outputs(376) <= not((layer3_outputs(333)) and (layer3_outputs(2687)));
    layer4_outputs(377) <= (layer3_outputs(6453)) and not (layer3_outputs(4431));
    layer4_outputs(378) <= (layer3_outputs(2087)) or (layer3_outputs(132));
    layer4_outputs(379) <= layer3_outputs(730);
    layer4_outputs(380) <= not(layer3_outputs(3879));
    layer4_outputs(381) <= (layer3_outputs(19)) and not (layer3_outputs(1144));
    layer4_outputs(382) <= not(layer3_outputs(2172));
    layer4_outputs(383) <= (layer3_outputs(2541)) or (layer3_outputs(4325));
    layer4_outputs(384) <= not(layer3_outputs(3394)) or (layer3_outputs(417));
    layer4_outputs(385) <= (layer3_outputs(1568)) and (layer3_outputs(2970));
    layer4_outputs(386) <= not(layer3_outputs(5730)) or (layer3_outputs(4052));
    layer4_outputs(387) <= not(layer3_outputs(56));
    layer4_outputs(388) <= layer3_outputs(513);
    layer4_outputs(389) <= '0';
    layer4_outputs(390) <= not(layer3_outputs(95)) or (layer3_outputs(3103));
    layer4_outputs(391) <= layer3_outputs(3133);
    layer4_outputs(392) <= (layer3_outputs(5882)) and (layer3_outputs(7170));
    layer4_outputs(393) <= layer3_outputs(4528);
    layer4_outputs(394) <= (layer3_outputs(5532)) and (layer3_outputs(3553));
    layer4_outputs(395) <= '0';
    layer4_outputs(396) <= layer3_outputs(7670);
    layer4_outputs(397) <= '1';
    layer4_outputs(398) <= not(layer3_outputs(6221));
    layer4_outputs(399) <= (layer3_outputs(2569)) and not (layer3_outputs(7623));
    layer4_outputs(400) <= layer3_outputs(2918);
    layer4_outputs(401) <= '0';
    layer4_outputs(402) <= not((layer3_outputs(830)) or (layer3_outputs(4322)));
    layer4_outputs(403) <= not(layer3_outputs(6375));
    layer4_outputs(404) <= not(layer3_outputs(2117));
    layer4_outputs(405) <= not(layer3_outputs(3620));
    layer4_outputs(406) <= (layer3_outputs(6057)) or (layer3_outputs(5397));
    layer4_outputs(407) <= not(layer3_outputs(1762));
    layer4_outputs(408) <= not((layer3_outputs(1662)) and (layer3_outputs(496)));
    layer4_outputs(409) <= not(layer3_outputs(7245));
    layer4_outputs(410) <= '0';
    layer4_outputs(411) <= (layer3_outputs(4120)) and not (layer3_outputs(2268));
    layer4_outputs(412) <= layer3_outputs(5195);
    layer4_outputs(413) <= not(layer3_outputs(7362));
    layer4_outputs(414) <= not(layer3_outputs(2438));
    layer4_outputs(415) <= not((layer3_outputs(1169)) and (layer3_outputs(4515)));
    layer4_outputs(416) <= layer3_outputs(1654);
    layer4_outputs(417) <= not(layer3_outputs(2428));
    layer4_outputs(418) <= not(layer3_outputs(1948));
    layer4_outputs(419) <= layer3_outputs(6581);
    layer4_outputs(420) <= not(layer3_outputs(6786));
    layer4_outputs(421) <= not(layer3_outputs(3398)) or (layer3_outputs(4822));
    layer4_outputs(422) <= not(layer3_outputs(180));
    layer4_outputs(423) <= layer3_outputs(6833);
    layer4_outputs(424) <= layer3_outputs(289);
    layer4_outputs(425) <= (layer3_outputs(1319)) and not (layer3_outputs(6508));
    layer4_outputs(426) <= layer3_outputs(4511);
    layer4_outputs(427) <= not(layer3_outputs(5006));
    layer4_outputs(428) <= not(layer3_outputs(3757)) or (layer3_outputs(1376));
    layer4_outputs(429) <= not(layer3_outputs(768));
    layer4_outputs(430) <= not(layer3_outputs(1749));
    layer4_outputs(431) <= '1';
    layer4_outputs(432) <= not(layer3_outputs(1543)) or (layer3_outputs(7487));
    layer4_outputs(433) <= (layer3_outputs(2920)) or (layer3_outputs(4765));
    layer4_outputs(434) <= not((layer3_outputs(5049)) or (layer3_outputs(136)));
    layer4_outputs(435) <= '0';
    layer4_outputs(436) <= not(layer3_outputs(5497));
    layer4_outputs(437) <= layer3_outputs(2489);
    layer4_outputs(438) <= not(layer3_outputs(4355));
    layer4_outputs(439) <= '1';
    layer4_outputs(440) <= not((layer3_outputs(481)) xor (layer3_outputs(2466)));
    layer4_outputs(441) <= not((layer3_outputs(4569)) or (layer3_outputs(6417)));
    layer4_outputs(442) <= not(layer3_outputs(3713)) or (layer3_outputs(5709));
    layer4_outputs(443) <= not(layer3_outputs(1963));
    layer4_outputs(444) <= layer3_outputs(1406);
    layer4_outputs(445) <= '0';
    layer4_outputs(446) <= layer3_outputs(5320);
    layer4_outputs(447) <= '1';
    layer4_outputs(448) <= layer3_outputs(1470);
    layer4_outputs(449) <= '0';
    layer4_outputs(450) <= (layer3_outputs(4197)) or (layer3_outputs(809));
    layer4_outputs(451) <= not(layer3_outputs(4847));
    layer4_outputs(452) <= (layer3_outputs(556)) and not (layer3_outputs(136));
    layer4_outputs(453) <= (layer3_outputs(4499)) and not (layer3_outputs(6451));
    layer4_outputs(454) <= not(layer3_outputs(2591)) or (layer3_outputs(70));
    layer4_outputs(455) <= layer3_outputs(314);
    layer4_outputs(456) <= not((layer3_outputs(4500)) and (layer3_outputs(1165)));
    layer4_outputs(457) <= (layer3_outputs(1891)) and (layer3_outputs(5023));
    layer4_outputs(458) <= layer3_outputs(5181);
    layer4_outputs(459) <= layer3_outputs(5244);
    layer4_outputs(460) <= layer3_outputs(2304);
    layer4_outputs(461) <= (layer3_outputs(903)) and not (layer3_outputs(566));
    layer4_outputs(462) <= layer3_outputs(2366);
    layer4_outputs(463) <= not(layer3_outputs(3522)) or (layer3_outputs(1113));
    layer4_outputs(464) <= (layer3_outputs(337)) and not (layer3_outputs(2736));
    layer4_outputs(465) <= layer3_outputs(585);
    layer4_outputs(466) <= '0';
    layer4_outputs(467) <= layer3_outputs(2530);
    layer4_outputs(468) <= (layer3_outputs(6565)) and not (layer3_outputs(6496));
    layer4_outputs(469) <= layer3_outputs(6672);
    layer4_outputs(470) <= not((layer3_outputs(4841)) or (layer3_outputs(778)));
    layer4_outputs(471) <= layer3_outputs(6543);
    layer4_outputs(472) <= layer3_outputs(2739);
    layer4_outputs(473) <= not(layer3_outputs(820));
    layer4_outputs(474) <= not(layer3_outputs(3756)) or (layer3_outputs(896));
    layer4_outputs(475) <= (layer3_outputs(6748)) and (layer3_outputs(5816));
    layer4_outputs(476) <= layer3_outputs(1176);
    layer4_outputs(477) <= (layer3_outputs(4764)) or (layer3_outputs(3177));
    layer4_outputs(478) <= layer3_outputs(927);
    layer4_outputs(479) <= (layer3_outputs(399)) or (layer3_outputs(5938));
    layer4_outputs(480) <= not(layer3_outputs(5980)) or (layer3_outputs(3346));
    layer4_outputs(481) <= not(layer3_outputs(41));
    layer4_outputs(482) <= not((layer3_outputs(344)) or (layer3_outputs(7162)));
    layer4_outputs(483) <= layer3_outputs(7508);
    layer4_outputs(484) <= not(layer3_outputs(5976));
    layer4_outputs(485) <= layer3_outputs(7170);
    layer4_outputs(486) <= not(layer3_outputs(3175)) or (layer3_outputs(4719));
    layer4_outputs(487) <= not(layer3_outputs(594));
    layer4_outputs(488) <= not((layer3_outputs(4548)) and (layer3_outputs(6424)));
    layer4_outputs(489) <= (layer3_outputs(4845)) or (layer3_outputs(3172));
    layer4_outputs(490) <= not(layer3_outputs(7077));
    layer4_outputs(491) <= (layer3_outputs(4993)) and not (layer3_outputs(2769));
    layer4_outputs(492) <= not((layer3_outputs(1557)) and (layer3_outputs(1617)));
    layer4_outputs(493) <= (layer3_outputs(1203)) and not (layer3_outputs(949));
    layer4_outputs(494) <= layer3_outputs(2060);
    layer4_outputs(495) <= layer3_outputs(5211);
    layer4_outputs(496) <= (layer3_outputs(1886)) and not (layer3_outputs(6924));
    layer4_outputs(497) <= '1';
    layer4_outputs(498) <= not(layer3_outputs(3978)) or (layer3_outputs(7644));
    layer4_outputs(499) <= not(layer3_outputs(4379));
    layer4_outputs(500) <= layer3_outputs(561);
    layer4_outputs(501) <= (layer3_outputs(2572)) and not (layer3_outputs(5391));
    layer4_outputs(502) <= (layer3_outputs(3155)) and (layer3_outputs(6865));
    layer4_outputs(503) <= (layer3_outputs(5405)) or (layer3_outputs(5635));
    layer4_outputs(504) <= not(layer3_outputs(550));
    layer4_outputs(505) <= not(layer3_outputs(2352));
    layer4_outputs(506) <= not(layer3_outputs(87)) or (layer3_outputs(3772));
    layer4_outputs(507) <= (layer3_outputs(1453)) or (layer3_outputs(4228));
    layer4_outputs(508) <= (layer3_outputs(3880)) and not (layer3_outputs(5674));
    layer4_outputs(509) <= layer3_outputs(6488);
    layer4_outputs(510) <= not((layer3_outputs(5440)) xor (layer3_outputs(6101)));
    layer4_outputs(511) <= not(layer3_outputs(2311));
    layer4_outputs(512) <= layer3_outputs(450);
    layer4_outputs(513) <= not((layer3_outputs(644)) xor (layer3_outputs(4649)));
    layer4_outputs(514) <= layer3_outputs(822);
    layer4_outputs(515) <= (layer3_outputs(572)) and (layer3_outputs(4670));
    layer4_outputs(516) <= layer3_outputs(5933);
    layer4_outputs(517) <= not(layer3_outputs(4234)) or (layer3_outputs(5694));
    layer4_outputs(518) <= (layer3_outputs(1843)) and not (layer3_outputs(4221));
    layer4_outputs(519) <= (layer3_outputs(2576)) xor (layer3_outputs(526));
    layer4_outputs(520) <= (layer3_outputs(2725)) and not (layer3_outputs(1048));
    layer4_outputs(521) <= (layer3_outputs(5142)) xor (layer3_outputs(6286));
    layer4_outputs(522) <= not((layer3_outputs(923)) and (layer3_outputs(2065)));
    layer4_outputs(523) <= not(layer3_outputs(1018)) or (layer3_outputs(2418));
    layer4_outputs(524) <= layer3_outputs(6366);
    layer4_outputs(525) <= layer3_outputs(1131);
    layer4_outputs(526) <= not(layer3_outputs(2165)) or (layer3_outputs(2577));
    layer4_outputs(527) <= not(layer3_outputs(3334)) or (layer3_outputs(5664));
    layer4_outputs(528) <= (layer3_outputs(5947)) and not (layer3_outputs(2192));
    layer4_outputs(529) <= (layer3_outputs(7241)) and (layer3_outputs(3903));
    layer4_outputs(530) <= (layer3_outputs(3582)) and (layer3_outputs(4939));
    layer4_outputs(531) <= not((layer3_outputs(4351)) xor (layer3_outputs(867)));
    layer4_outputs(532) <= not((layer3_outputs(5522)) or (layer3_outputs(299)));
    layer4_outputs(533) <= (layer3_outputs(7323)) or (layer3_outputs(5196));
    layer4_outputs(534) <= not(layer3_outputs(1845));
    layer4_outputs(535) <= layer3_outputs(4655);
    layer4_outputs(536) <= (layer3_outputs(1718)) and (layer3_outputs(7507));
    layer4_outputs(537) <= not((layer3_outputs(102)) or (layer3_outputs(5620)));
    layer4_outputs(538) <= not(layer3_outputs(1302));
    layer4_outputs(539) <= not((layer3_outputs(6170)) or (layer3_outputs(2703)));
    layer4_outputs(540) <= layer3_outputs(4360);
    layer4_outputs(541) <= not((layer3_outputs(5713)) and (layer3_outputs(7679)));
    layer4_outputs(542) <= (layer3_outputs(5538)) and (layer3_outputs(5924));
    layer4_outputs(543) <= (layer3_outputs(2509)) and not (layer3_outputs(7382));
    layer4_outputs(544) <= (layer3_outputs(2464)) and (layer3_outputs(5431));
    layer4_outputs(545) <= not(layer3_outputs(2204));
    layer4_outputs(546) <= not(layer3_outputs(2088)) or (layer3_outputs(7010));
    layer4_outputs(547) <= not(layer3_outputs(3837));
    layer4_outputs(548) <= not(layer3_outputs(2995));
    layer4_outputs(549) <= (layer3_outputs(7516)) or (layer3_outputs(4659));
    layer4_outputs(550) <= (layer3_outputs(3056)) xor (layer3_outputs(1081));
    layer4_outputs(551) <= (layer3_outputs(4540)) or (layer3_outputs(1679));
    layer4_outputs(552) <= (layer3_outputs(1770)) and (layer3_outputs(4482));
    layer4_outputs(553) <= not(layer3_outputs(4895)) or (layer3_outputs(1395));
    layer4_outputs(554) <= not((layer3_outputs(1023)) xor (layer3_outputs(6967)));
    layer4_outputs(555) <= not(layer3_outputs(5505)) or (layer3_outputs(6351));
    layer4_outputs(556) <= not(layer3_outputs(5236));
    layer4_outputs(557) <= layer3_outputs(1750);
    layer4_outputs(558) <= not(layer3_outputs(2386));
    layer4_outputs(559) <= (layer3_outputs(3075)) and (layer3_outputs(3543));
    layer4_outputs(560) <= layer3_outputs(4702);
    layer4_outputs(561) <= layer3_outputs(7368);
    layer4_outputs(562) <= not(layer3_outputs(3732));
    layer4_outputs(563) <= not(layer3_outputs(5360));
    layer4_outputs(564) <= layer3_outputs(2342);
    layer4_outputs(565) <= not(layer3_outputs(2479));
    layer4_outputs(566) <= not(layer3_outputs(3362)) or (layer3_outputs(5624));
    layer4_outputs(567) <= (layer3_outputs(5468)) xor (layer3_outputs(3295));
    layer4_outputs(568) <= not((layer3_outputs(823)) or (layer3_outputs(1233)));
    layer4_outputs(569) <= not(layer3_outputs(2484));
    layer4_outputs(570) <= '0';
    layer4_outputs(571) <= '1';
    layer4_outputs(572) <= not(layer3_outputs(573));
    layer4_outputs(573) <= layer3_outputs(5960);
    layer4_outputs(574) <= (layer3_outputs(4349)) and not (layer3_outputs(729));
    layer4_outputs(575) <= layer3_outputs(897);
    layer4_outputs(576) <= (layer3_outputs(2460)) and (layer3_outputs(5333));
    layer4_outputs(577) <= layer3_outputs(1527);
    layer4_outputs(578) <= not((layer3_outputs(5093)) or (layer3_outputs(4330)));
    layer4_outputs(579) <= (layer3_outputs(312)) xor (layer3_outputs(7617));
    layer4_outputs(580) <= layer3_outputs(7026);
    layer4_outputs(581) <= (layer3_outputs(307)) or (layer3_outputs(3231));
    layer4_outputs(582) <= layer3_outputs(1189);
    layer4_outputs(583) <= not(layer3_outputs(1025));
    layer4_outputs(584) <= (layer3_outputs(7349)) and (layer3_outputs(7520));
    layer4_outputs(585) <= '1';
    layer4_outputs(586) <= not((layer3_outputs(5881)) and (layer3_outputs(894)));
    layer4_outputs(587) <= not((layer3_outputs(1024)) xor (layer3_outputs(1614)));
    layer4_outputs(588) <= (layer3_outputs(5998)) or (layer3_outputs(6216));
    layer4_outputs(589) <= layer3_outputs(4246);
    layer4_outputs(590) <= (layer3_outputs(703)) or (layer3_outputs(1436));
    layer4_outputs(591) <= layer3_outputs(1754);
    layer4_outputs(592) <= (layer3_outputs(6953)) xor (layer3_outputs(6004));
    layer4_outputs(593) <= not(layer3_outputs(6168));
    layer4_outputs(594) <= (layer3_outputs(5028)) or (layer3_outputs(4301));
    layer4_outputs(595) <= (layer3_outputs(5348)) and not (layer3_outputs(3563));
    layer4_outputs(596) <= not(layer3_outputs(2635));
    layer4_outputs(597) <= not(layer3_outputs(6814));
    layer4_outputs(598) <= not(layer3_outputs(3774));
    layer4_outputs(599) <= '0';
    layer4_outputs(600) <= not((layer3_outputs(5355)) xor (layer3_outputs(5712)));
    layer4_outputs(601) <= layer3_outputs(6291);
    layer4_outputs(602) <= (layer3_outputs(3438)) or (layer3_outputs(1284));
    layer4_outputs(603) <= not(layer3_outputs(5065));
    layer4_outputs(604) <= layer3_outputs(883);
    layer4_outputs(605) <= (layer3_outputs(6133)) and (layer3_outputs(5201));
    layer4_outputs(606) <= not(layer3_outputs(6967)) or (layer3_outputs(7595));
    layer4_outputs(607) <= layer3_outputs(1659);
    layer4_outputs(608) <= (layer3_outputs(1739)) or (layer3_outputs(2520));
    layer4_outputs(609) <= (layer3_outputs(728)) and (layer3_outputs(1602));
    layer4_outputs(610) <= layer3_outputs(5513);
    layer4_outputs(611) <= layer3_outputs(1748);
    layer4_outputs(612) <= (layer3_outputs(2770)) and not (layer3_outputs(5562));
    layer4_outputs(613) <= layer3_outputs(3039);
    layer4_outputs(614) <= not(layer3_outputs(1910)) or (layer3_outputs(913));
    layer4_outputs(615) <= (layer3_outputs(3564)) and (layer3_outputs(7083));
    layer4_outputs(616) <= not(layer3_outputs(1890)) or (layer3_outputs(1723));
    layer4_outputs(617) <= layer3_outputs(6184);
    layer4_outputs(618) <= not(layer3_outputs(4916)) or (layer3_outputs(5259));
    layer4_outputs(619) <= not(layer3_outputs(1342));
    layer4_outputs(620) <= not(layer3_outputs(7613)) or (layer3_outputs(4422));
    layer4_outputs(621) <= not(layer3_outputs(5275));
    layer4_outputs(622) <= '0';
    layer4_outputs(623) <= '1';
    layer4_outputs(624) <= not(layer3_outputs(2745));
    layer4_outputs(625) <= (layer3_outputs(3255)) and (layer3_outputs(7499));
    layer4_outputs(626) <= not(layer3_outputs(3110));
    layer4_outputs(627) <= layer3_outputs(3390);
    layer4_outputs(628) <= '0';
    layer4_outputs(629) <= not((layer3_outputs(7201)) and (layer3_outputs(2078)));
    layer4_outputs(630) <= not(layer3_outputs(6467));
    layer4_outputs(631) <= '1';
    layer4_outputs(632) <= layer3_outputs(5976);
    layer4_outputs(633) <= (layer3_outputs(3950)) and not (layer3_outputs(6373));
    layer4_outputs(634) <= (layer3_outputs(4539)) and not (layer3_outputs(7544));
    layer4_outputs(635) <= '1';
    layer4_outputs(636) <= layer3_outputs(224);
    layer4_outputs(637) <= '1';
    layer4_outputs(638) <= not(layer3_outputs(5333));
    layer4_outputs(639) <= (layer3_outputs(2620)) and (layer3_outputs(3015));
    layer4_outputs(640) <= (layer3_outputs(5836)) and (layer3_outputs(5046));
    layer4_outputs(641) <= (layer3_outputs(2729)) and not (layer3_outputs(7416));
    layer4_outputs(642) <= (layer3_outputs(5452)) and (layer3_outputs(5975));
    layer4_outputs(643) <= (layer3_outputs(4417)) and not (layer3_outputs(5787));
    layer4_outputs(644) <= not(layer3_outputs(595));
    layer4_outputs(645) <= layer3_outputs(957);
    layer4_outputs(646) <= not(layer3_outputs(5760)) or (layer3_outputs(4524));
    layer4_outputs(647) <= not((layer3_outputs(2729)) xor (layer3_outputs(561)));
    layer4_outputs(648) <= layer3_outputs(3760);
    layer4_outputs(649) <= (layer3_outputs(5296)) and not (layer3_outputs(1084));
    layer4_outputs(650) <= (layer3_outputs(500)) and not (layer3_outputs(891));
    layer4_outputs(651) <= (layer3_outputs(1863)) and not (layer3_outputs(5078));
    layer4_outputs(652) <= layer3_outputs(5621);
    layer4_outputs(653) <= (layer3_outputs(7167)) or (layer3_outputs(969));
    layer4_outputs(654) <= not((layer3_outputs(6636)) and (layer3_outputs(3678)));
    layer4_outputs(655) <= not(layer3_outputs(2901));
    layer4_outputs(656) <= not(layer3_outputs(6006)) or (layer3_outputs(672));
    layer4_outputs(657) <= not(layer3_outputs(2803)) or (layer3_outputs(1840));
    layer4_outputs(658) <= not(layer3_outputs(5626));
    layer4_outputs(659) <= not((layer3_outputs(1330)) or (layer3_outputs(3383)));
    layer4_outputs(660) <= not(layer3_outputs(2830));
    layer4_outputs(661) <= '0';
    layer4_outputs(662) <= not((layer3_outputs(4638)) or (layer3_outputs(7596)));
    layer4_outputs(663) <= layer3_outputs(4413);
    layer4_outputs(664) <= layer3_outputs(6368);
    layer4_outputs(665) <= layer3_outputs(2792);
    layer4_outputs(666) <= (layer3_outputs(3130)) and not (layer3_outputs(6863));
    layer4_outputs(667) <= not(layer3_outputs(1040));
    layer4_outputs(668) <= not(layer3_outputs(7572));
    layer4_outputs(669) <= not(layer3_outputs(6232)) or (layer3_outputs(5586));
    layer4_outputs(670) <= (layer3_outputs(6580)) xor (layer3_outputs(3300));
    layer4_outputs(671) <= not(layer3_outputs(7465)) or (layer3_outputs(5894));
    layer4_outputs(672) <= not((layer3_outputs(3498)) and (layer3_outputs(6959)));
    layer4_outputs(673) <= layer3_outputs(3266);
    layer4_outputs(674) <= (layer3_outputs(7489)) and (layer3_outputs(2276));
    layer4_outputs(675) <= not((layer3_outputs(580)) and (layer3_outputs(1100)));
    layer4_outputs(676) <= not(layer3_outputs(3427)) or (layer3_outputs(4107));
    layer4_outputs(677) <= not(layer3_outputs(5463));
    layer4_outputs(678) <= not(layer3_outputs(4010));
    layer4_outputs(679) <= not(layer3_outputs(3155));
    layer4_outputs(680) <= layer3_outputs(2828);
    layer4_outputs(681) <= not(layer3_outputs(6080));
    layer4_outputs(682) <= not(layer3_outputs(4633));
    layer4_outputs(683) <= not(layer3_outputs(7607)) or (layer3_outputs(7441));
    layer4_outputs(684) <= not(layer3_outputs(2755));
    layer4_outputs(685) <= not((layer3_outputs(1882)) xor (layer3_outputs(4670)));
    layer4_outputs(686) <= layer3_outputs(3519);
    layer4_outputs(687) <= (layer3_outputs(5649)) xor (layer3_outputs(2278));
    layer4_outputs(688) <= not(layer3_outputs(3454));
    layer4_outputs(689) <= not(layer3_outputs(3211)) or (layer3_outputs(7334));
    layer4_outputs(690) <= not(layer3_outputs(432));
    layer4_outputs(691) <= not((layer3_outputs(2086)) and (layer3_outputs(1001)));
    layer4_outputs(692) <= '1';
    layer4_outputs(693) <= not((layer3_outputs(6809)) and (layer3_outputs(608)));
    layer4_outputs(694) <= layer3_outputs(3056);
    layer4_outputs(695) <= layer3_outputs(4426);
    layer4_outputs(696) <= not(layer3_outputs(5080));
    layer4_outputs(697) <= not(layer3_outputs(6220));
    layer4_outputs(698) <= not((layer3_outputs(7234)) and (layer3_outputs(7419)));
    layer4_outputs(699) <= not(layer3_outputs(1078));
    layer4_outputs(700) <= (layer3_outputs(6117)) xor (layer3_outputs(4216));
    layer4_outputs(701) <= (layer3_outputs(6619)) and (layer3_outputs(4488));
    layer4_outputs(702) <= not((layer3_outputs(2445)) or (layer3_outputs(127)));
    layer4_outputs(703) <= not((layer3_outputs(5608)) and (layer3_outputs(6189)));
    layer4_outputs(704) <= not(layer3_outputs(3507));
    layer4_outputs(705) <= not(layer3_outputs(7169));
    layer4_outputs(706) <= (layer3_outputs(3273)) and not (layer3_outputs(554));
    layer4_outputs(707) <= layer3_outputs(4972);
    layer4_outputs(708) <= not(layer3_outputs(1579));
    layer4_outputs(709) <= layer3_outputs(7422);
    layer4_outputs(710) <= not(layer3_outputs(3698)) or (layer3_outputs(717));
    layer4_outputs(711) <= layer3_outputs(1228);
    layer4_outputs(712) <= (layer3_outputs(6144)) and (layer3_outputs(6864));
    layer4_outputs(713) <= not(layer3_outputs(4389));
    layer4_outputs(714) <= not((layer3_outputs(4740)) or (layer3_outputs(4155)));
    layer4_outputs(715) <= (layer3_outputs(5139)) and not (layer3_outputs(2416));
    layer4_outputs(716) <= not((layer3_outputs(78)) or (layer3_outputs(663)));
    layer4_outputs(717) <= (layer3_outputs(5873)) and not (layer3_outputs(3704));
    layer4_outputs(718) <= not(layer3_outputs(32)) or (layer3_outputs(4409));
    layer4_outputs(719) <= not((layer3_outputs(3757)) and (layer3_outputs(7399)));
    layer4_outputs(720) <= '1';
    layer4_outputs(721) <= not((layer3_outputs(4000)) or (layer3_outputs(4739)));
    layer4_outputs(722) <= (layer3_outputs(3232)) and not (layer3_outputs(4269));
    layer4_outputs(723) <= not((layer3_outputs(7566)) and (layer3_outputs(6215)));
    layer4_outputs(724) <= layer3_outputs(3559);
    layer4_outputs(725) <= (layer3_outputs(7156)) or (layer3_outputs(3225));
    layer4_outputs(726) <= not(layer3_outputs(2032));
    layer4_outputs(727) <= layer3_outputs(2215);
    layer4_outputs(728) <= layer3_outputs(7591);
    layer4_outputs(729) <= (layer3_outputs(3844)) and not (layer3_outputs(2895));
    layer4_outputs(730) <= not(layer3_outputs(5412));
    layer4_outputs(731) <= not(layer3_outputs(4640));
    layer4_outputs(732) <= (layer3_outputs(811)) or (layer3_outputs(5776));
    layer4_outputs(733) <= not(layer3_outputs(1588));
    layer4_outputs(734) <= layer3_outputs(5595);
    layer4_outputs(735) <= (layer3_outputs(7499)) or (layer3_outputs(42));
    layer4_outputs(736) <= not(layer3_outputs(4747));
    layer4_outputs(737) <= not(layer3_outputs(7006));
    layer4_outputs(738) <= not(layer3_outputs(4368));
    layer4_outputs(739) <= (layer3_outputs(6705)) or (layer3_outputs(2020));
    layer4_outputs(740) <= not(layer3_outputs(3430));
    layer4_outputs(741) <= not((layer3_outputs(5213)) and (layer3_outputs(5545)));
    layer4_outputs(742) <= not(layer3_outputs(5163));
    layer4_outputs(743) <= not((layer3_outputs(1229)) or (layer3_outputs(3675)));
    layer4_outputs(744) <= (layer3_outputs(4166)) xor (layer3_outputs(3560));
    layer4_outputs(745) <= not(layer3_outputs(5188));
    layer4_outputs(746) <= not(layer3_outputs(2220));
    layer4_outputs(747) <= (layer3_outputs(4856)) and (layer3_outputs(7276));
    layer4_outputs(748) <= layer3_outputs(1278);
    layer4_outputs(749) <= (layer3_outputs(3872)) and not (layer3_outputs(7429));
    layer4_outputs(750) <= not(layer3_outputs(71));
    layer4_outputs(751) <= not(layer3_outputs(1624));
    layer4_outputs(752) <= '1';
    layer4_outputs(753) <= not(layer3_outputs(1827));
    layer4_outputs(754) <= not(layer3_outputs(1398));
    layer4_outputs(755) <= not(layer3_outputs(2362)) or (layer3_outputs(7599));
    layer4_outputs(756) <= not((layer3_outputs(6471)) and (layer3_outputs(3059)));
    layer4_outputs(757) <= (layer3_outputs(6799)) and not (layer3_outputs(2847));
    layer4_outputs(758) <= not((layer3_outputs(6444)) xor (layer3_outputs(4528)));
    layer4_outputs(759) <= not(layer3_outputs(226)) or (layer3_outputs(2426));
    layer4_outputs(760) <= (layer3_outputs(4140)) xor (layer3_outputs(1402));
    layer4_outputs(761) <= (layer3_outputs(2928)) xor (layer3_outputs(25));
    layer4_outputs(762) <= not(layer3_outputs(7227));
    layer4_outputs(763) <= not(layer3_outputs(1805));
    layer4_outputs(764) <= not(layer3_outputs(7282));
    layer4_outputs(765) <= (layer3_outputs(79)) and not (layer3_outputs(4181));
    layer4_outputs(766) <= not(layer3_outputs(1948));
    layer4_outputs(767) <= (layer3_outputs(945)) and not (layer3_outputs(2851));
    layer4_outputs(768) <= (layer3_outputs(196)) and not (layer3_outputs(221));
    layer4_outputs(769) <= not(layer3_outputs(306));
    layer4_outputs(770) <= '1';
    layer4_outputs(771) <= not(layer3_outputs(4677)) or (layer3_outputs(6637));
    layer4_outputs(772) <= layer3_outputs(5277);
    layer4_outputs(773) <= not(layer3_outputs(4419));
    layer4_outputs(774) <= (layer3_outputs(6103)) xor (layer3_outputs(7250));
    layer4_outputs(775) <= (layer3_outputs(7157)) xor (layer3_outputs(5484));
    layer4_outputs(776) <= layer3_outputs(1578);
    layer4_outputs(777) <= layer3_outputs(746);
    layer4_outputs(778) <= layer3_outputs(2184);
    layer4_outputs(779) <= (layer3_outputs(3012)) or (layer3_outputs(7109));
    layer4_outputs(780) <= not((layer3_outputs(7652)) or (layer3_outputs(1039)));
    layer4_outputs(781) <= not(layer3_outputs(207));
    layer4_outputs(782) <= not(layer3_outputs(5800));
    layer4_outputs(783) <= (layer3_outputs(1731)) and (layer3_outputs(4573));
    layer4_outputs(784) <= layer3_outputs(1054);
    layer4_outputs(785) <= (layer3_outputs(1060)) xor (layer3_outputs(4064));
    layer4_outputs(786) <= '1';
    layer4_outputs(787) <= (layer3_outputs(7107)) and not (layer3_outputs(2767));
    layer4_outputs(788) <= layer3_outputs(6017);
    layer4_outputs(789) <= not(layer3_outputs(3395));
    layer4_outputs(790) <= layer3_outputs(5744);
    layer4_outputs(791) <= not(layer3_outputs(3283));
    layer4_outputs(792) <= layer3_outputs(5267);
    layer4_outputs(793) <= not(layer3_outputs(2266)) or (layer3_outputs(590));
    layer4_outputs(794) <= (layer3_outputs(543)) and not (layer3_outputs(4794));
    layer4_outputs(795) <= '0';
    layer4_outputs(796) <= not(layer3_outputs(4808));
    layer4_outputs(797) <= (layer3_outputs(4604)) and not (layer3_outputs(3584));
    layer4_outputs(798) <= layer3_outputs(318);
    layer4_outputs(799) <= not(layer3_outputs(2104));
    layer4_outputs(800) <= layer3_outputs(3967);
    layer4_outputs(801) <= layer3_outputs(889);
    layer4_outputs(802) <= not(layer3_outputs(4870));
    layer4_outputs(803) <= (layer3_outputs(7055)) and (layer3_outputs(6335));
    layer4_outputs(804) <= not(layer3_outputs(4426));
    layer4_outputs(805) <= not(layer3_outputs(166));
    layer4_outputs(806) <= layer3_outputs(7449);
    layer4_outputs(807) <= layer3_outputs(1750);
    layer4_outputs(808) <= not(layer3_outputs(1088)) or (layer3_outputs(1179));
    layer4_outputs(809) <= layer3_outputs(4596);
    layer4_outputs(810) <= not((layer3_outputs(226)) xor (layer3_outputs(5430)));
    layer4_outputs(811) <= not(layer3_outputs(7044));
    layer4_outputs(812) <= (layer3_outputs(1368)) or (layer3_outputs(2321));
    layer4_outputs(813) <= not(layer3_outputs(205)) or (layer3_outputs(6604));
    layer4_outputs(814) <= layer3_outputs(57);
    layer4_outputs(815) <= not(layer3_outputs(2153));
    layer4_outputs(816) <= not(layer3_outputs(4978));
    layer4_outputs(817) <= not((layer3_outputs(3615)) or (layer3_outputs(7057)));
    layer4_outputs(818) <= not((layer3_outputs(5501)) or (layer3_outputs(4777)));
    layer4_outputs(819) <= not(layer3_outputs(5063)) or (layer3_outputs(3486));
    layer4_outputs(820) <= not(layer3_outputs(3616));
    layer4_outputs(821) <= not((layer3_outputs(5936)) and (layer3_outputs(57)));
    layer4_outputs(822) <= not((layer3_outputs(14)) and (layer3_outputs(6888)));
    layer4_outputs(823) <= (layer3_outputs(7645)) and not (layer3_outputs(7321));
    layer4_outputs(824) <= layer3_outputs(6517);
    layer4_outputs(825) <= '0';
    layer4_outputs(826) <= not(layer3_outputs(1298));
    layer4_outputs(827) <= not(layer3_outputs(4594)) or (layer3_outputs(469));
    layer4_outputs(828) <= not((layer3_outputs(5074)) xor (layer3_outputs(5754)));
    layer4_outputs(829) <= '1';
    layer4_outputs(830) <= layer3_outputs(3786);
    layer4_outputs(831) <= not(layer3_outputs(3658));
    layer4_outputs(832) <= '1';
    layer4_outputs(833) <= (layer3_outputs(1595)) and not (layer3_outputs(2044));
    layer4_outputs(834) <= not((layer3_outputs(6655)) and (layer3_outputs(6128)));
    layer4_outputs(835) <= '0';
    layer4_outputs(836) <= not((layer3_outputs(5009)) xor (layer3_outputs(1204)));
    layer4_outputs(837) <= (layer3_outputs(1098)) and not (layer3_outputs(506));
    layer4_outputs(838) <= (layer3_outputs(1535)) and not (layer3_outputs(4745));
    layer4_outputs(839) <= not((layer3_outputs(4651)) and (layer3_outputs(1365)));
    layer4_outputs(840) <= (layer3_outputs(3016)) and not (layer3_outputs(1464));
    layer4_outputs(841) <= not(layer3_outputs(6757)) or (layer3_outputs(1877));
    layer4_outputs(842) <= layer3_outputs(7301);
    layer4_outputs(843) <= not((layer3_outputs(8)) or (layer3_outputs(5685)));
    layer4_outputs(844) <= not(layer3_outputs(1307)) or (layer3_outputs(5310));
    layer4_outputs(845) <= '0';
    layer4_outputs(846) <= (layer3_outputs(4503)) xor (layer3_outputs(7158));
    layer4_outputs(847) <= layer3_outputs(5988);
    layer4_outputs(848) <= not(layer3_outputs(6350)) or (layer3_outputs(343));
    layer4_outputs(849) <= layer3_outputs(4565);
    layer4_outputs(850) <= (layer3_outputs(6521)) and not (layer3_outputs(7662));
    layer4_outputs(851) <= not(layer3_outputs(6297));
    layer4_outputs(852) <= (layer3_outputs(5452)) and not (layer3_outputs(3431));
    layer4_outputs(853) <= layer3_outputs(3599);
    layer4_outputs(854) <= not(layer3_outputs(6060));
    layer4_outputs(855) <= layer3_outputs(7252);
    layer4_outputs(856) <= layer3_outputs(1014);
    layer4_outputs(857) <= layer3_outputs(6928);
    layer4_outputs(858) <= not(layer3_outputs(6583));
    layer4_outputs(859) <= not(layer3_outputs(4865));
    layer4_outputs(860) <= not((layer3_outputs(1742)) xor (layer3_outputs(3294)));
    layer4_outputs(861) <= not(layer3_outputs(6925));
    layer4_outputs(862) <= not(layer3_outputs(3270)) or (layer3_outputs(1681));
    layer4_outputs(863) <= (layer3_outputs(7287)) xor (layer3_outputs(2562));
    layer4_outputs(864) <= layer3_outputs(4041);
    layer4_outputs(865) <= layer3_outputs(4043);
    layer4_outputs(866) <= layer3_outputs(7528);
    layer4_outputs(867) <= not((layer3_outputs(4280)) and (layer3_outputs(5681)));
    layer4_outputs(868) <= layer3_outputs(1779);
    layer4_outputs(869) <= not(layer3_outputs(6832)) or (layer3_outputs(7623));
    layer4_outputs(870) <= '1';
    layer4_outputs(871) <= layer3_outputs(2442);
    layer4_outputs(872) <= layer3_outputs(1912);
    layer4_outputs(873) <= not(layer3_outputs(6421));
    layer4_outputs(874) <= not((layer3_outputs(3974)) or (layer3_outputs(2338)));
    layer4_outputs(875) <= layer3_outputs(6930);
    layer4_outputs(876) <= not(layer3_outputs(1908));
    layer4_outputs(877) <= not((layer3_outputs(1870)) and (layer3_outputs(1936)));
    layer4_outputs(878) <= layer3_outputs(4012);
    layer4_outputs(879) <= not(layer3_outputs(6802)) or (layer3_outputs(6098));
    layer4_outputs(880) <= (layer3_outputs(4291)) and not (layer3_outputs(7272));
    layer4_outputs(881) <= not(layer3_outputs(839)) or (layer3_outputs(7264));
    layer4_outputs(882) <= not(layer3_outputs(3111));
    layer4_outputs(883) <= not(layer3_outputs(6227));
    layer4_outputs(884) <= not(layer3_outputs(7464));
    layer4_outputs(885) <= not(layer3_outputs(7478));
    layer4_outputs(886) <= (layer3_outputs(6990)) and not (layer3_outputs(2582));
    layer4_outputs(887) <= '0';
    layer4_outputs(888) <= not(layer3_outputs(6801));
    layer4_outputs(889) <= (layer3_outputs(3152)) or (layer3_outputs(1558));
    layer4_outputs(890) <= layer3_outputs(2819);
    layer4_outputs(891) <= not(layer3_outputs(140));
    layer4_outputs(892) <= not(layer3_outputs(6356)) or (layer3_outputs(2977));
    layer4_outputs(893) <= (layer3_outputs(7144)) and not (layer3_outputs(1880));
    layer4_outputs(894) <= not(layer3_outputs(3873));
    layer4_outputs(895) <= not(layer3_outputs(5962)) or (layer3_outputs(6165));
    layer4_outputs(896) <= not((layer3_outputs(6209)) and (layer3_outputs(4364)));
    layer4_outputs(897) <= (layer3_outputs(2337)) and not (layer3_outputs(2540));
    layer4_outputs(898) <= not(layer3_outputs(3318)) or (layer3_outputs(7525));
    layer4_outputs(899) <= (layer3_outputs(2397)) and (layer3_outputs(676));
    layer4_outputs(900) <= (layer3_outputs(837)) and not (layer3_outputs(880));
    layer4_outputs(901) <= (layer3_outputs(7492)) and not (layer3_outputs(2413));
    layer4_outputs(902) <= layer3_outputs(6609);
    layer4_outputs(903) <= not(layer3_outputs(4791)) or (layer3_outputs(6461));
    layer4_outputs(904) <= layer3_outputs(1666);
    layer4_outputs(905) <= not(layer3_outputs(4961));
    layer4_outputs(906) <= not(layer3_outputs(456));
    layer4_outputs(907) <= not(layer3_outputs(5325));
    layer4_outputs(908) <= '1';
    layer4_outputs(909) <= layer3_outputs(2054);
    layer4_outputs(910) <= not(layer3_outputs(5535));
    layer4_outputs(911) <= not(layer3_outputs(7424));
    layer4_outputs(912) <= (layer3_outputs(5883)) and (layer3_outputs(728));
    layer4_outputs(913) <= not((layer3_outputs(7021)) xor (layer3_outputs(1907)));
    layer4_outputs(914) <= not(layer3_outputs(4675)) or (layer3_outputs(3869));
    layer4_outputs(915) <= (layer3_outputs(7367)) and not (layer3_outputs(1466));
    layer4_outputs(916) <= layer3_outputs(3994);
    layer4_outputs(917) <= layer3_outputs(6841);
    layer4_outputs(918) <= (layer3_outputs(2094)) or (layer3_outputs(1947));
    layer4_outputs(919) <= not(layer3_outputs(5654));
    layer4_outputs(920) <= (layer3_outputs(2077)) and (layer3_outputs(2742));
    layer4_outputs(921) <= layer3_outputs(4482);
    layer4_outputs(922) <= layer3_outputs(913);
    layer4_outputs(923) <= '0';
    layer4_outputs(924) <= not((layer3_outputs(2598)) or (layer3_outputs(744)));
    layer4_outputs(925) <= not(layer3_outputs(6334));
    layer4_outputs(926) <= (layer3_outputs(3182)) and not (layer3_outputs(6226));
    layer4_outputs(927) <= not((layer3_outputs(4831)) or (layer3_outputs(4153)));
    layer4_outputs(928) <= (layer3_outputs(5754)) and not (layer3_outputs(6171));
    layer4_outputs(929) <= not(layer3_outputs(2992));
    layer4_outputs(930) <= not(layer3_outputs(4529)) or (layer3_outputs(2055));
    layer4_outputs(931) <= not(layer3_outputs(5996)) or (layer3_outputs(2835));
    layer4_outputs(932) <= layer3_outputs(820);
    layer4_outputs(933) <= not((layer3_outputs(7312)) and (layer3_outputs(3292)));
    layer4_outputs(934) <= layer3_outputs(4510);
    layer4_outputs(935) <= layer3_outputs(3129);
    layer4_outputs(936) <= not((layer3_outputs(342)) and (layer3_outputs(2474)));
    layer4_outputs(937) <= (layer3_outputs(2260)) xor (layer3_outputs(1503));
    layer4_outputs(938) <= not(layer3_outputs(65));
    layer4_outputs(939) <= layer3_outputs(188);
    layer4_outputs(940) <= not(layer3_outputs(3596));
    layer4_outputs(941) <= layer3_outputs(2867);
    layer4_outputs(942) <= (layer3_outputs(4264)) xor (layer3_outputs(7075));
    layer4_outputs(943) <= (layer3_outputs(4745)) xor (layer3_outputs(6765));
    layer4_outputs(944) <= layer3_outputs(201);
    layer4_outputs(945) <= not((layer3_outputs(5169)) or (layer3_outputs(3447)));
    layer4_outputs(946) <= not((layer3_outputs(4545)) and (layer3_outputs(5092)));
    layer4_outputs(947) <= '0';
    layer4_outputs(948) <= not((layer3_outputs(7022)) or (layer3_outputs(7179)));
    layer4_outputs(949) <= layer3_outputs(7523);
    layer4_outputs(950) <= '1';
    layer4_outputs(951) <= layer3_outputs(5652);
    layer4_outputs(952) <= (layer3_outputs(7350)) and (layer3_outputs(6840));
    layer4_outputs(953) <= not(layer3_outputs(4711));
    layer4_outputs(954) <= not(layer3_outputs(5773));
    layer4_outputs(955) <= layer3_outputs(5765);
    layer4_outputs(956) <= (layer3_outputs(2084)) and not (layer3_outputs(5153));
    layer4_outputs(957) <= (layer3_outputs(7539)) and not (layer3_outputs(1580));
    layer4_outputs(958) <= (layer3_outputs(3840)) and not (layer3_outputs(1207));
    layer4_outputs(959) <= not(layer3_outputs(473));
    layer4_outputs(960) <= not(layer3_outputs(7651));
    layer4_outputs(961) <= layer3_outputs(4710);
    layer4_outputs(962) <= (layer3_outputs(7430)) or (layer3_outputs(5293));
    layer4_outputs(963) <= (layer3_outputs(2135)) and (layer3_outputs(1379));
    layer4_outputs(964) <= layer3_outputs(1946);
    layer4_outputs(965) <= not(layer3_outputs(3055)) or (layer3_outputs(5439));
    layer4_outputs(966) <= (layer3_outputs(2016)) and not (layer3_outputs(103));
    layer4_outputs(967) <= not(layer3_outputs(4945)) or (layer3_outputs(1861));
    layer4_outputs(968) <= (layer3_outputs(3151)) or (layer3_outputs(6883));
    layer4_outputs(969) <= not((layer3_outputs(5951)) or (layer3_outputs(1665)));
    layer4_outputs(970) <= (layer3_outputs(7220)) and (layer3_outputs(439));
    layer4_outputs(971) <= '1';
    layer4_outputs(972) <= not((layer3_outputs(3767)) and (layer3_outputs(7466)));
    layer4_outputs(973) <= not(layer3_outputs(414));
    layer4_outputs(974) <= not(layer3_outputs(5274));
    layer4_outputs(975) <= not(layer3_outputs(4361));
    layer4_outputs(976) <= (layer3_outputs(5613)) xor (layer3_outputs(5987));
    layer4_outputs(977) <= (layer3_outputs(7081)) and not (layer3_outputs(3699));
    layer4_outputs(978) <= layer3_outputs(4534);
    layer4_outputs(979) <= not(layer3_outputs(6898));
    layer4_outputs(980) <= not(layer3_outputs(6087)) or (layer3_outputs(1826));
    layer4_outputs(981) <= (layer3_outputs(642)) and not (layer3_outputs(2956));
    layer4_outputs(982) <= not(layer3_outputs(1456));
    layer4_outputs(983) <= not(layer3_outputs(4128));
    layer4_outputs(984) <= not((layer3_outputs(5283)) or (layer3_outputs(668)));
    layer4_outputs(985) <= layer3_outputs(6025);
    layer4_outputs(986) <= (layer3_outputs(1210)) or (layer3_outputs(2564));
    layer4_outputs(987) <= (layer3_outputs(4034)) and not (layer3_outputs(1433));
    layer4_outputs(988) <= (layer3_outputs(629)) and not (layer3_outputs(2781));
    layer4_outputs(989) <= layer3_outputs(2883);
    layer4_outputs(990) <= not((layer3_outputs(7226)) and (layer3_outputs(5098)));
    layer4_outputs(991) <= not(layer3_outputs(3331));
    layer4_outputs(992) <= not(layer3_outputs(3094));
    layer4_outputs(993) <= layer3_outputs(618);
    layer4_outputs(994) <= layer3_outputs(5609);
    layer4_outputs(995) <= (layer3_outputs(1271)) and (layer3_outputs(3246));
    layer4_outputs(996) <= layer3_outputs(774);
    layer4_outputs(997) <= not(layer3_outputs(4688));
    layer4_outputs(998) <= (layer3_outputs(2297)) and (layer3_outputs(5553));
    layer4_outputs(999) <= (layer3_outputs(7356)) or (layer3_outputs(2790));
    layer4_outputs(1000) <= not((layer3_outputs(290)) or (layer3_outputs(5237)));
    layer4_outputs(1001) <= (layer3_outputs(2680)) xor (layer3_outputs(983));
    layer4_outputs(1002) <= not(layer3_outputs(3813));
    layer4_outputs(1003) <= (layer3_outputs(2937)) and not (layer3_outputs(5925));
    layer4_outputs(1004) <= (layer3_outputs(1907)) xor (layer3_outputs(5710));
    layer4_outputs(1005) <= not(layer3_outputs(3811)) or (layer3_outputs(582));
    layer4_outputs(1006) <= layer3_outputs(3913);
    layer4_outputs(1007) <= not(layer3_outputs(3105));
    layer4_outputs(1008) <= (layer3_outputs(1157)) and (layer3_outputs(1394));
    layer4_outputs(1009) <= layer3_outputs(1286);
    layer4_outputs(1010) <= not((layer3_outputs(4169)) or (layer3_outputs(4521)));
    layer4_outputs(1011) <= not(layer3_outputs(4750)) or (layer3_outputs(1537));
    layer4_outputs(1012) <= layer3_outputs(407);
    layer4_outputs(1013) <= not(layer3_outputs(5750));
    layer4_outputs(1014) <= (layer3_outputs(486)) and not (layer3_outputs(4517));
    layer4_outputs(1015) <= (layer3_outputs(1574)) and not (layer3_outputs(3455));
    layer4_outputs(1016) <= not((layer3_outputs(3419)) or (layer3_outputs(7677)));
    layer4_outputs(1017) <= layer3_outputs(6878);
    layer4_outputs(1018) <= not((layer3_outputs(3364)) xor (layer3_outputs(3755)));
    layer4_outputs(1019) <= layer3_outputs(6359);
    layer4_outputs(1020) <= not(layer3_outputs(6125)) or (layer3_outputs(2830));
    layer4_outputs(1021) <= (layer3_outputs(1674)) or (layer3_outputs(5759));
    layer4_outputs(1022) <= layer3_outputs(3350);
    layer4_outputs(1023) <= (layer3_outputs(3043)) and (layer3_outputs(524));
    layer4_outputs(1024) <= not((layer3_outputs(3806)) or (layer3_outputs(4623)));
    layer4_outputs(1025) <= not(layer3_outputs(4259));
    layer4_outputs(1026) <= layer3_outputs(4113);
    layer4_outputs(1027) <= layer3_outputs(7048);
    layer4_outputs(1028) <= not(layer3_outputs(5993)) or (layer3_outputs(1875));
    layer4_outputs(1029) <= not(layer3_outputs(1586)) or (layer3_outputs(1881));
    layer4_outputs(1030) <= (layer3_outputs(6704)) xor (layer3_outputs(154));
    layer4_outputs(1031) <= (layer3_outputs(1622)) and (layer3_outputs(6828));
    layer4_outputs(1032) <= not((layer3_outputs(1155)) or (layer3_outputs(3771)));
    layer4_outputs(1033) <= '1';
    layer4_outputs(1034) <= (layer3_outputs(702)) and (layer3_outputs(7008));
    layer4_outputs(1035) <= not(layer3_outputs(2821));
    layer4_outputs(1036) <= (layer3_outputs(5803)) or (layer3_outputs(4298));
    layer4_outputs(1037) <= '0';
    layer4_outputs(1038) <= (layer3_outputs(137)) and not (layer3_outputs(1501));
    layer4_outputs(1039) <= not((layer3_outputs(6848)) or (layer3_outputs(6361)));
    layer4_outputs(1040) <= (layer3_outputs(1719)) xor (layer3_outputs(2273));
    layer4_outputs(1041) <= layer3_outputs(6689);
    layer4_outputs(1042) <= not((layer3_outputs(503)) xor (layer3_outputs(549)));
    layer4_outputs(1043) <= layer3_outputs(3910);
    layer4_outputs(1044) <= '0';
    layer4_outputs(1045) <= not(layer3_outputs(6728)) or (layer3_outputs(2709));
    layer4_outputs(1046) <= not(layer3_outputs(7213)) or (layer3_outputs(2748));
    layer4_outputs(1047) <= '1';
    layer4_outputs(1048) <= not(layer3_outputs(537));
    layer4_outputs(1049) <= not(layer3_outputs(2550));
    layer4_outputs(1050) <= (layer3_outputs(1804)) and not (layer3_outputs(4606));
    layer4_outputs(1051) <= not((layer3_outputs(5799)) or (layer3_outputs(4354)));
    layer4_outputs(1052) <= layer3_outputs(6741);
    layer4_outputs(1053) <= not(layer3_outputs(1591));
    layer4_outputs(1054) <= not(layer3_outputs(2701)) or (layer3_outputs(4316));
    layer4_outputs(1055) <= not(layer3_outputs(1961));
    layer4_outputs(1056) <= layer3_outputs(954);
    layer4_outputs(1057) <= not(layer3_outputs(1923));
    layer4_outputs(1058) <= layer3_outputs(869);
    layer4_outputs(1059) <= not((layer3_outputs(4665)) and (layer3_outputs(6380)));
    layer4_outputs(1060) <= not(layer3_outputs(7466));
    layer4_outputs(1061) <= (layer3_outputs(2717)) and (layer3_outputs(1178));
    layer4_outputs(1062) <= layer3_outputs(7518);
    layer4_outputs(1063) <= (layer3_outputs(899)) and not (layer3_outputs(6285));
    layer4_outputs(1064) <= not(layer3_outputs(7374));
    layer4_outputs(1065) <= not((layer3_outputs(422)) and (layer3_outputs(525)));
    layer4_outputs(1066) <= '1';
    layer4_outputs(1067) <= layer3_outputs(2677);
    layer4_outputs(1068) <= (layer3_outputs(5328)) and not (layer3_outputs(5549));
    layer4_outputs(1069) <= layer3_outputs(5198);
    layer4_outputs(1070) <= layer3_outputs(3883);
    layer4_outputs(1071) <= layer3_outputs(451);
    layer4_outputs(1072) <= not(layer3_outputs(2287)) or (layer3_outputs(2896));
    layer4_outputs(1073) <= not(layer3_outputs(1163));
    layer4_outputs(1074) <= layer3_outputs(6150);
    layer4_outputs(1075) <= (layer3_outputs(7283)) or (layer3_outputs(5342));
    layer4_outputs(1076) <= layer3_outputs(1739);
    layer4_outputs(1077) <= (layer3_outputs(3928)) or (layer3_outputs(1516));
    layer4_outputs(1078) <= (layer3_outputs(1279)) and (layer3_outputs(4063));
    layer4_outputs(1079) <= not(layer3_outputs(1542)) or (layer3_outputs(4747));
    layer4_outputs(1080) <= not(layer3_outputs(2662));
    layer4_outputs(1081) <= not(layer3_outputs(6648)) or (layer3_outputs(393));
    layer4_outputs(1082) <= not((layer3_outputs(5010)) or (layer3_outputs(3860)));
    layer4_outputs(1083) <= layer3_outputs(6314);
    layer4_outputs(1084) <= layer3_outputs(4118);
    layer4_outputs(1085) <= '0';
    layer4_outputs(1086) <= (layer3_outputs(4608)) and (layer3_outputs(4376));
    layer4_outputs(1087) <= layer3_outputs(7059);
    layer4_outputs(1088) <= not(layer3_outputs(2825));
    layer4_outputs(1089) <= not((layer3_outputs(5832)) or (layer3_outputs(3317)));
    layer4_outputs(1090) <= (layer3_outputs(3649)) or (layer3_outputs(1110));
    layer4_outputs(1091) <= (layer3_outputs(2800)) and (layer3_outputs(483));
    layer4_outputs(1092) <= not(layer3_outputs(2404));
    layer4_outputs(1093) <= not(layer3_outputs(5812)) or (layer3_outputs(1836));
    layer4_outputs(1094) <= layer3_outputs(1262);
    layer4_outputs(1095) <= not(layer3_outputs(1147)) or (layer3_outputs(5129));
    layer4_outputs(1096) <= not((layer3_outputs(5996)) and (layer3_outputs(3391)));
    layer4_outputs(1097) <= not(layer3_outputs(6270));
    layer4_outputs(1098) <= (layer3_outputs(3599)) and not (layer3_outputs(3046));
    layer4_outputs(1099) <= '1';
    layer4_outputs(1100) <= not(layer3_outputs(6051));
    layer4_outputs(1101) <= (layer3_outputs(6009)) and not (layer3_outputs(4761));
    layer4_outputs(1102) <= not(layer3_outputs(2686)) or (layer3_outputs(1392));
    layer4_outputs(1103) <= not((layer3_outputs(1726)) and (layer3_outputs(4307)));
    layer4_outputs(1104) <= '0';
    layer4_outputs(1105) <= not(layer3_outputs(4854));
    layer4_outputs(1106) <= not(layer3_outputs(4925)) or (layer3_outputs(2097));
    layer4_outputs(1107) <= (layer3_outputs(104)) and not (layer3_outputs(699));
    layer4_outputs(1108) <= layer3_outputs(3906);
    layer4_outputs(1109) <= layer3_outputs(1521);
    layer4_outputs(1110) <= layer3_outputs(7575);
    layer4_outputs(1111) <= not(layer3_outputs(1455));
    layer4_outputs(1112) <= not((layer3_outputs(3186)) and (layer3_outputs(5362)));
    layer4_outputs(1113) <= not(layer3_outputs(106));
    layer4_outputs(1114) <= not((layer3_outputs(3285)) and (layer3_outputs(6500)));
    layer4_outputs(1115) <= not(layer3_outputs(3054));
    layer4_outputs(1116) <= not((layer3_outputs(2598)) and (layer3_outputs(5663)));
    layer4_outputs(1117) <= (layer3_outputs(747)) and not (layer3_outputs(2132));
    layer4_outputs(1118) <= not(layer3_outputs(1301)) or (layer3_outputs(7100));
    layer4_outputs(1119) <= not(layer3_outputs(2285)) or (layer3_outputs(2065));
    layer4_outputs(1120) <= layer3_outputs(3172);
    layer4_outputs(1121) <= (layer3_outputs(1618)) and not (layer3_outputs(5691));
    layer4_outputs(1122) <= '1';
    layer4_outputs(1123) <= not(layer3_outputs(7127)) or (layer3_outputs(1923));
    layer4_outputs(1124) <= layer3_outputs(3197);
    layer4_outputs(1125) <= not((layer3_outputs(6719)) and (layer3_outputs(1627)));
    layer4_outputs(1126) <= not(layer3_outputs(3876));
    layer4_outputs(1127) <= (layer3_outputs(1779)) or (layer3_outputs(6644));
    layer4_outputs(1128) <= (layer3_outputs(930)) xor (layer3_outputs(1789));
    layer4_outputs(1129) <= layer3_outputs(320);
    layer4_outputs(1130) <= not(layer3_outputs(5631));
    layer4_outputs(1131) <= (layer3_outputs(4253)) and not (layer3_outputs(2533));
    layer4_outputs(1132) <= not((layer3_outputs(3764)) and (layer3_outputs(6614)));
    layer4_outputs(1133) <= (layer3_outputs(3995)) or (layer3_outputs(6962));
    layer4_outputs(1134) <= (layer3_outputs(956)) and not (layer3_outputs(7047));
    layer4_outputs(1135) <= (layer3_outputs(6039)) or (layer3_outputs(656));
    layer4_outputs(1136) <= '1';
    layer4_outputs(1137) <= not(layer3_outputs(3105)) or (layer3_outputs(956));
    layer4_outputs(1138) <= (layer3_outputs(4785)) or (layer3_outputs(3334));
    layer4_outputs(1139) <= layer3_outputs(757);
    layer4_outputs(1140) <= not((layer3_outputs(2239)) and (layer3_outputs(7510)));
    layer4_outputs(1141) <= not((layer3_outputs(200)) and (layer3_outputs(5596)));
    layer4_outputs(1142) <= (layer3_outputs(1815)) xor (layer3_outputs(3628));
    layer4_outputs(1143) <= not(layer3_outputs(6425));
    layer4_outputs(1144) <= '1';
    layer4_outputs(1145) <= '0';
    layer4_outputs(1146) <= not(layer3_outputs(2187));
    layer4_outputs(1147) <= (layer3_outputs(3990)) and (layer3_outputs(6407));
    layer4_outputs(1148) <= '1';
    layer4_outputs(1149) <= (layer3_outputs(5372)) and not (layer3_outputs(3726));
    layer4_outputs(1150) <= (layer3_outputs(3916)) or (layer3_outputs(7457));
    layer4_outputs(1151) <= not(layer3_outputs(6536)) or (layer3_outputs(3004));
    layer4_outputs(1152) <= (layer3_outputs(5392)) and not (layer3_outputs(6869));
    layer4_outputs(1153) <= not((layer3_outputs(6333)) and (layer3_outputs(2636)));
    layer4_outputs(1154) <= layer3_outputs(280);
    layer4_outputs(1155) <= (layer3_outputs(1275)) and (layer3_outputs(5961));
    layer4_outputs(1156) <= (layer3_outputs(5255)) or (layer3_outputs(7144));
    layer4_outputs(1157) <= (layer3_outputs(7509)) and (layer3_outputs(4759));
    layer4_outputs(1158) <= '0';
    layer4_outputs(1159) <= not(layer3_outputs(7385)) or (layer3_outputs(5653));
    layer4_outputs(1160) <= (layer3_outputs(1482)) and (layer3_outputs(2212));
    layer4_outputs(1161) <= '1';
    layer4_outputs(1162) <= not(layer3_outputs(3725)) or (layer3_outputs(3329));
    layer4_outputs(1163) <= not(layer3_outputs(7569));
    layer4_outputs(1164) <= not(layer3_outputs(7100)) or (layer3_outputs(1127));
    layer4_outputs(1165) <= (layer3_outputs(1564)) and not (layer3_outputs(4174));
    layer4_outputs(1166) <= not(layer3_outputs(6548));
    layer4_outputs(1167) <= '1';
    layer4_outputs(1168) <= not(layer3_outputs(2279));
    layer4_outputs(1169) <= (layer3_outputs(5006)) and (layer3_outputs(4055));
    layer4_outputs(1170) <= not(layer3_outputs(7298));
    layer4_outputs(1171) <= (layer3_outputs(7368)) and (layer3_outputs(24));
    layer4_outputs(1172) <= not((layer3_outputs(64)) or (layer3_outputs(998)));
    layer4_outputs(1173) <= layer3_outputs(6087);
    layer4_outputs(1174) <= not(layer3_outputs(5479)) or (layer3_outputs(622));
    layer4_outputs(1175) <= layer3_outputs(978);
    layer4_outputs(1176) <= layer3_outputs(1637);
    layer4_outputs(1177) <= layer3_outputs(1909);
    layer4_outputs(1178) <= not((layer3_outputs(1323)) or (layer3_outputs(4751)));
    layer4_outputs(1179) <= layer3_outputs(2003);
    layer4_outputs(1180) <= not(layer3_outputs(3360)) or (layer3_outputs(5077));
    layer4_outputs(1181) <= not(layer3_outputs(1841));
    layer4_outputs(1182) <= (layer3_outputs(1399)) or (layer3_outputs(1990));
    layer4_outputs(1183) <= not((layer3_outputs(6056)) or (layer3_outputs(173)));
    layer4_outputs(1184) <= not(layer3_outputs(1624));
    layer4_outputs(1185) <= (layer3_outputs(6868)) and not (layer3_outputs(3821));
    layer4_outputs(1186) <= not(layer3_outputs(4859));
    layer4_outputs(1187) <= (layer3_outputs(4411)) xor (layer3_outputs(632));
    layer4_outputs(1188) <= (layer3_outputs(3394)) and not (layer3_outputs(2713));
    layer4_outputs(1189) <= not((layer3_outputs(3058)) and (layer3_outputs(5985)));
    layer4_outputs(1190) <= layer3_outputs(3782);
    layer4_outputs(1191) <= (layer3_outputs(6192)) and not (layer3_outputs(7160));
    layer4_outputs(1192) <= not(layer3_outputs(5672)) or (layer3_outputs(3959));
    layer4_outputs(1193) <= not(layer3_outputs(6468));
    layer4_outputs(1194) <= layer3_outputs(269);
    layer4_outputs(1195) <= not(layer3_outputs(7313));
    layer4_outputs(1196) <= (layer3_outputs(3315)) and (layer3_outputs(345));
    layer4_outputs(1197) <= (layer3_outputs(7423)) and not (layer3_outputs(438));
    layer4_outputs(1198) <= (layer3_outputs(1177)) and not (layer3_outputs(6418));
    layer4_outputs(1199) <= (layer3_outputs(470)) xor (layer3_outputs(878));
    layer4_outputs(1200) <= (layer3_outputs(939)) xor (layer3_outputs(546));
    layer4_outputs(1201) <= (layer3_outputs(2393)) xor (layer3_outputs(6336));
    layer4_outputs(1202) <= '0';
    layer4_outputs(1203) <= layer3_outputs(3057);
    layer4_outputs(1204) <= not((layer3_outputs(1807)) and (layer3_outputs(3166)));
    layer4_outputs(1205) <= (layer3_outputs(3946)) or (layer3_outputs(1873));
    layer4_outputs(1206) <= (layer3_outputs(1778)) and not (layer3_outputs(534));
    layer4_outputs(1207) <= not((layer3_outputs(1904)) and (layer3_outputs(7604)));
    layer4_outputs(1208) <= not(layer3_outputs(6610));
    layer4_outputs(1209) <= '1';
    layer4_outputs(1210) <= (layer3_outputs(7382)) or (layer3_outputs(717));
    layer4_outputs(1211) <= layer3_outputs(2802);
    layer4_outputs(1212) <= layer3_outputs(2347);
    layer4_outputs(1213) <= not(layer3_outputs(5924));
    layer4_outputs(1214) <= (layer3_outputs(4348)) and not (layer3_outputs(5125));
    layer4_outputs(1215) <= not(layer3_outputs(4744));
    layer4_outputs(1216) <= (layer3_outputs(5425)) or (layer3_outputs(6201));
    layer4_outputs(1217) <= not((layer3_outputs(7054)) and (layer3_outputs(278)));
    layer4_outputs(1218) <= layer3_outputs(1642);
    layer4_outputs(1219) <= not((layer3_outputs(5058)) and (layer3_outputs(7395)));
    layer4_outputs(1220) <= layer3_outputs(4248);
    layer4_outputs(1221) <= not(layer3_outputs(6617));
    layer4_outputs(1222) <= (layer3_outputs(2350)) and not (layer3_outputs(2834));
    layer4_outputs(1223) <= layer3_outputs(856);
    layer4_outputs(1224) <= (layer3_outputs(2347)) and not (layer3_outputs(3627));
    layer4_outputs(1225) <= not(layer3_outputs(6683));
    layer4_outputs(1226) <= (layer3_outputs(2566)) xor (layer3_outputs(6071));
    layer4_outputs(1227) <= (layer3_outputs(1386)) and (layer3_outputs(6856));
    layer4_outputs(1228) <= not(layer3_outputs(4188));
    layer4_outputs(1229) <= layer3_outputs(1885);
    layer4_outputs(1230) <= layer3_outputs(2987);
    layer4_outputs(1231) <= layer3_outputs(5241);
    layer4_outputs(1232) <= (layer3_outputs(546)) xor (layer3_outputs(6753));
    layer4_outputs(1233) <= layer3_outputs(4695);
    layer4_outputs(1234) <= not((layer3_outputs(6445)) and (layer3_outputs(995)));
    layer4_outputs(1235) <= (layer3_outputs(1420)) and not (layer3_outputs(7184));
    layer4_outputs(1236) <= not(layer3_outputs(760));
    layer4_outputs(1237) <= layer3_outputs(3859);
    layer4_outputs(1238) <= not((layer3_outputs(4048)) xor (layer3_outputs(3952)));
    layer4_outputs(1239) <= not(layer3_outputs(4549));
    layer4_outputs(1240) <= layer3_outputs(2092);
    layer4_outputs(1241) <= '0';
    layer4_outputs(1242) <= not(layer3_outputs(1324));
    layer4_outputs(1243) <= (layer3_outputs(2268)) or (layer3_outputs(3027));
    layer4_outputs(1244) <= (layer3_outputs(4672)) xor (layer3_outputs(7600));
    layer4_outputs(1245) <= (layer3_outputs(1162)) and (layer3_outputs(2180));
    layer4_outputs(1246) <= (layer3_outputs(5989)) and (layer3_outputs(2161));
    layer4_outputs(1247) <= '1';
    layer4_outputs(1248) <= layer3_outputs(6083);
    layer4_outputs(1249) <= (layer3_outputs(7583)) and not (layer3_outputs(708));
    layer4_outputs(1250) <= layer3_outputs(5157);
    layer4_outputs(1251) <= layer3_outputs(4496);
    layer4_outputs(1252) <= not(layer3_outputs(1931));
    layer4_outputs(1253) <= layer3_outputs(6318);
    layer4_outputs(1254) <= layer3_outputs(1296);
    layer4_outputs(1255) <= not(layer3_outputs(6893));
    layer4_outputs(1256) <= not(layer3_outputs(2197));
    layer4_outputs(1257) <= layer3_outputs(4425);
    layer4_outputs(1258) <= (layer3_outputs(1957)) xor (layer3_outputs(35));
    layer4_outputs(1259) <= not(layer3_outputs(3042));
    layer4_outputs(1260) <= (layer3_outputs(1390)) and (layer3_outputs(2099));
    layer4_outputs(1261) <= not((layer3_outputs(6754)) or (layer3_outputs(4145)));
    layer4_outputs(1262) <= layer3_outputs(698);
    layer4_outputs(1263) <= not(layer3_outputs(1969));
    layer4_outputs(1264) <= layer3_outputs(3735);
    layer4_outputs(1265) <= (layer3_outputs(3274)) and not (layer3_outputs(7562));
    layer4_outputs(1266) <= layer3_outputs(4508);
    layer4_outputs(1267) <= (layer3_outputs(1064)) xor (layer3_outputs(4281));
    layer4_outputs(1268) <= not((layer3_outputs(3026)) or (layer3_outputs(1299)));
    layer4_outputs(1269) <= not(layer3_outputs(6854)) or (layer3_outputs(5313));
    layer4_outputs(1270) <= not(layer3_outputs(109));
    layer4_outputs(1271) <= not(layer3_outputs(1384)) or (layer3_outputs(6688));
    layer4_outputs(1272) <= layer3_outputs(5490);
    layer4_outputs(1273) <= layer3_outputs(1986);
    layer4_outputs(1274) <= not(layer3_outputs(7192)) or (layer3_outputs(4354));
    layer4_outputs(1275) <= layer3_outputs(1532);
    layer4_outputs(1276) <= not((layer3_outputs(7147)) or (layer3_outputs(7553)));
    layer4_outputs(1277) <= not(layer3_outputs(7344));
    layer4_outputs(1278) <= not((layer3_outputs(2519)) and (layer3_outputs(5016)));
    layer4_outputs(1279) <= not(layer3_outputs(5584));
    layer4_outputs(1280) <= not(layer3_outputs(5966)) or (layer3_outputs(4187));
    layer4_outputs(1281) <= not((layer3_outputs(1677)) and (layer3_outputs(665)));
    layer4_outputs(1282) <= not((layer3_outputs(6149)) or (layer3_outputs(6746)));
    layer4_outputs(1283) <= layer3_outputs(5706);
    layer4_outputs(1284) <= not(layer3_outputs(7407)) or (layer3_outputs(1553));
    layer4_outputs(1285) <= not(layer3_outputs(3390));
    layer4_outputs(1286) <= layer3_outputs(3769);
    layer4_outputs(1287) <= not((layer3_outputs(3365)) or (layer3_outputs(952)));
    layer4_outputs(1288) <= (layer3_outputs(370)) or (layer3_outputs(3485));
    layer4_outputs(1289) <= layer3_outputs(7533);
    layer4_outputs(1290) <= (layer3_outputs(4935)) and not (layer3_outputs(7550));
    layer4_outputs(1291) <= not(layer3_outputs(1293)) or (layer3_outputs(3457));
    layer4_outputs(1292) <= not(layer3_outputs(2990));
    layer4_outputs(1293) <= layer3_outputs(3894);
    layer4_outputs(1294) <= not(layer3_outputs(164));
    layer4_outputs(1295) <= layer3_outputs(2463);
    layer4_outputs(1296) <= layer3_outputs(7265);
    layer4_outputs(1297) <= (layer3_outputs(5900)) xor (layer3_outputs(1404));
    layer4_outputs(1298) <= '1';
    layer4_outputs(1299) <= not(layer3_outputs(887));
    layer4_outputs(1300) <= not(layer3_outputs(4299));
    layer4_outputs(1301) <= (layer3_outputs(5382)) and not (layer3_outputs(3945));
    layer4_outputs(1302) <= (layer3_outputs(3744)) and not (layer3_outputs(2294));
    layer4_outputs(1303) <= (layer3_outputs(7460)) xor (layer3_outputs(6155));
    layer4_outputs(1304) <= (layer3_outputs(6950)) and (layer3_outputs(936));
    layer4_outputs(1305) <= (layer3_outputs(376)) and not (layer3_outputs(4668));
    layer4_outputs(1306) <= not(layer3_outputs(3243)) or (layer3_outputs(7025));
    layer4_outputs(1307) <= not(layer3_outputs(5782));
    layer4_outputs(1308) <= not(layer3_outputs(1554));
    layer4_outputs(1309) <= not(layer3_outputs(3029));
    layer4_outputs(1310) <= not((layer3_outputs(6080)) or (layer3_outputs(6397)));
    layer4_outputs(1311) <= not(layer3_outputs(1224));
    layer4_outputs(1312) <= layer3_outputs(6383);
    layer4_outputs(1313) <= (layer3_outputs(2626)) and (layer3_outputs(4709));
    layer4_outputs(1314) <= (layer3_outputs(6652)) and (layer3_outputs(6120));
    layer4_outputs(1315) <= layer3_outputs(1613);
    layer4_outputs(1316) <= not((layer3_outputs(3153)) or (layer3_outputs(430)));
    layer4_outputs(1317) <= (layer3_outputs(1249)) and (layer3_outputs(6896));
    layer4_outputs(1318) <= '0';
    layer4_outputs(1319) <= (layer3_outputs(4003)) and (layer3_outputs(383));
    layer4_outputs(1320) <= layer3_outputs(349);
    layer4_outputs(1321) <= not(layer3_outputs(2473));
    layer4_outputs(1322) <= (layer3_outputs(3443)) or (layer3_outputs(5245));
    layer4_outputs(1323) <= not((layer3_outputs(1416)) xor (layer3_outputs(5000)));
    layer4_outputs(1324) <= not((layer3_outputs(6333)) and (layer3_outputs(4304)));
    layer4_outputs(1325) <= not(layer3_outputs(347));
    layer4_outputs(1326) <= layer3_outputs(4765);
    layer4_outputs(1327) <= not(layer3_outputs(4435)) or (layer3_outputs(4740));
    layer4_outputs(1328) <= not((layer3_outputs(5637)) or (layer3_outputs(3817)));
    layer4_outputs(1329) <= not((layer3_outputs(1921)) or (layer3_outputs(375)));
    layer4_outputs(1330) <= not(layer3_outputs(6843)) or (layer3_outputs(1445));
    layer4_outputs(1331) <= layer3_outputs(5801);
    layer4_outputs(1332) <= layer3_outputs(2553);
    layer4_outputs(1333) <= not(layer3_outputs(2035));
    layer4_outputs(1334) <= not(layer3_outputs(5694)) or (layer3_outputs(2203));
    layer4_outputs(1335) <= not((layer3_outputs(64)) and (layer3_outputs(4460)));
    layer4_outputs(1336) <= not((layer3_outputs(2158)) and (layer3_outputs(5775)));
    layer4_outputs(1337) <= not(layer3_outputs(2205));
    layer4_outputs(1338) <= (layer3_outputs(4923)) or (layer3_outputs(4841));
    layer4_outputs(1339) <= not(layer3_outputs(6237));
    layer4_outputs(1340) <= not((layer3_outputs(7062)) xor (layer3_outputs(416)));
    layer4_outputs(1341) <= not(layer3_outputs(4642));
    layer4_outputs(1342) <= layer3_outputs(7252);
    layer4_outputs(1343) <= not((layer3_outputs(5132)) or (layer3_outputs(2474)));
    layer4_outputs(1344) <= not(layer3_outputs(1388));
    layer4_outputs(1345) <= (layer3_outputs(7164)) xor (layer3_outputs(1489));
    layer4_outputs(1346) <= (layer3_outputs(4694)) and not (layer3_outputs(1175));
    layer4_outputs(1347) <= (layer3_outputs(280)) and not (layer3_outputs(4968));
    layer4_outputs(1348) <= layer3_outputs(1584);
    layer4_outputs(1349) <= (layer3_outputs(5882)) or (layer3_outputs(2355));
    layer4_outputs(1350) <= not(layer3_outputs(6990));
    layer4_outputs(1351) <= not(layer3_outputs(6148));
    layer4_outputs(1352) <= '1';
    layer4_outputs(1353) <= layer3_outputs(453);
    layer4_outputs(1354) <= (layer3_outputs(4846)) and (layer3_outputs(4697));
    layer4_outputs(1355) <= not(layer3_outputs(357)) or (layer3_outputs(1421));
    layer4_outputs(1356) <= not(layer3_outputs(3013));
    layer4_outputs(1357) <= not((layer3_outputs(3656)) and (layer3_outputs(4494)));
    layer4_outputs(1358) <= not(layer3_outputs(169));
    layer4_outputs(1359) <= not((layer3_outputs(2516)) xor (layer3_outputs(2097)));
    layer4_outputs(1360) <= layer3_outputs(808);
    layer4_outputs(1361) <= layer3_outputs(563);
    layer4_outputs(1362) <= (layer3_outputs(3137)) and not (layer3_outputs(2899));
    layer4_outputs(1363) <= (layer3_outputs(2227)) and not (layer3_outputs(3039));
    layer4_outputs(1364) <= '0';
    layer4_outputs(1365) <= layer3_outputs(3578);
    layer4_outputs(1366) <= (layer3_outputs(5347)) and not (layer3_outputs(964));
    layer4_outputs(1367) <= (layer3_outputs(1439)) and not (layer3_outputs(5032));
    layer4_outputs(1368) <= '0';
    layer4_outputs(1369) <= '1';
    layer4_outputs(1370) <= not(layer3_outputs(1399));
    layer4_outputs(1371) <= not(layer3_outputs(1352));
    layer4_outputs(1372) <= not((layer3_outputs(3458)) or (layer3_outputs(1954)));
    layer4_outputs(1373) <= (layer3_outputs(3042)) and not (layer3_outputs(4035));
    layer4_outputs(1374) <= not(layer3_outputs(6266)) or (layer3_outputs(4827));
    layer4_outputs(1375) <= layer3_outputs(3549);
    layer4_outputs(1376) <= not(layer3_outputs(6765)) or (layer3_outputs(5097));
    layer4_outputs(1377) <= not(layer3_outputs(4252)) or (layer3_outputs(2253));
    layer4_outputs(1378) <= layer3_outputs(2240);
    layer4_outputs(1379) <= not((layer3_outputs(2185)) xor (layer3_outputs(4165)));
    layer4_outputs(1380) <= not(layer3_outputs(773));
    layer4_outputs(1381) <= (layer3_outputs(221)) and not (layer3_outputs(3030));
    layer4_outputs(1382) <= not(layer3_outputs(1585)) or (layer3_outputs(4825));
    layer4_outputs(1383) <= (layer3_outputs(7442)) and not (layer3_outputs(4271));
    layer4_outputs(1384) <= not((layer3_outputs(389)) xor (layer3_outputs(4876)));
    layer4_outputs(1385) <= not(layer3_outputs(5847));
    layer4_outputs(1386) <= layer3_outputs(5854);
    layer4_outputs(1387) <= layer3_outputs(7424);
    layer4_outputs(1388) <= (layer3_outputs(3332)) and (layer3_outputs(4346));
    layer4_outputs(1389) <= not(layer3_outputs(2466)) or (layer3_outputs(1182));
    layer4_outputs(1390) <= not((layer3_outputs(6515)) or (layer3_outputs(1269)));
    layer4_outputs(1391) <= not(layer3_outputs(2257));
    layer4_outputs(1392) <= not(layer3_outputs(6406)) or (layer3_outputs(4996));
    layer4_outputs(1393) <= layer3_outputs(3185);
    layer4_outputs(1394) <= not((layer3_outputs(3987)) and (layer3_outputs(7205)));
    layer4_outputs(1395) <= not((layer3_outputs(398)) and (layer3_outputs(6948)));
    layer4_outputs(1396) <= not(layer3_outputs(308)) or (layer3_outputs(496));
    layer4_outputs(1397) <= '1';
    layer4_outputs(1398) <= not(layer3_outputs(3309)) or (layer3_outputs(2771));
    layer4_outputs(1399) <= not(layer3_outputs(1808));
    layer4_outputs(1400) <= not(layer3_outputs(6630));
    layer4_outputs(1401) <= not(layer3_outputs(2177));
    layer4_outputs(1402) <= not((layer3_outputs(4277)) or (layer3_outputs(6454)));
    layer4_outputs(1403) <= not(layer3_outputs(2774));
    layer4_outputs(1404) <= '0';
    layer4_outputs(1405) <= not(layer3_outputs(402));
    layer4_outputs(1406) <= (layer3_outputs(975)) or (layer3_outputs(1283));
    layer4_outputs(1407) <= layer3_outputs(6179);
    layer4_outputs(1408) <= layer3_outputs(927);
    layer4_outputs(1409) <= not((layer3_outputs(4589)) and (layer3_outputs(5944)));
    layer4_outputs(1410) <= not(layer3_outputs(2056)) or (layer3_outputs(7103));
    layer4_outputs(1411) <= (layer3_outputs(6576)) and (layer3_outputs(4705));
    layer4_outputs(1412) <= not(layer3_outputs(3351));
    layer4_outputs(1413) <= layer3_outputs(2440);
    layer4_outputs(1414) <= '1';
    layer4_outputs(1415) <= layer3_outputs(725);
    layer4_outputs(1416) <= (layer3_outputs(5181)) or (layer3_outputs(6240));
    layer4_outputs(1417) <= not(layer3_outputs(3529));
    layer4_outputs(1418) <= not((layer3_outputs(3681)) xor (layer3_outputs(4701)));
    layer4_outputs(1419) <= not(layer3_outputs(5807));
    layer4_outputs(1420) <= not(layer3_outputs(4808));
    layer4_outputs(1421) <= layer3_outputs(1835);
    layer4_outputs(1422) <= (layer3_outputs(2542)) xor (layer3_outputs(3261));
    layer4_outputs(1423) <= (layer3_outputs(2101)) and not (layer3_outputs(7002));
    layer4_outputs(1424) <= (layer3_outputs(1480)) and not (layer3_outputs(4763));
    layer4_outputs(1425) <= not(layer3_outputs(4341)) or (layer3_outputs(26));
    layer4_outputs(1426) <= layer3_outputs(5629);
    layer4_outputs(1427) <= not((layer3_outputs(3637)) or (layer3_outputs(4126)));
    layer4_outputs(1428) <= not(layer3_outputs(4465)) or (layer3_outputs(5446));
    layer4_outputs(1429) <= (layer3_outputs(6792)) and not (layer3_outputs(5127));
    layer4_outputs(1430) <= not(layer3_outputs(6830));
    layer4_outputs(1431) <= not((layer3_outputs(4837)) and (layer3_outputs(3691)));
    layer4_outputs(1432) <= (layer3_outputs(4553)) and (layer3_outputs(6060));
    layer4_outputs(1433) <= not(layer3_outputs(1044)) or (layer3_outputs(3217));
    layer4_outputs(1434) <= not((layer3_outputs(5701)) or (layer3_outputs(2979)));
    layer4_outputs(1435) <= (layer3_outputs(6471)) and not (layer3_outputs(6435));
    layer4_outputs(1436) <= '1';
    layer4_outputs(1437) <= not(layer3_outputs(3653)) or (layer3_outputs(6544));
    layer4_outputs(1438) <= layer3_outputs(5240);
    layer4_outputs(1439) <= not((layer3_outputs(1148)) or (layer3_outputs(745)));
    layer4_outputs(1440) <= layer3_outputs(7507);
    layer4_outputs(1441) <= not((layer3_outputs(3259)) or (layer3_outputs(2723)));
    layer4_outputs(1442) <= not(layer3_outputs(1805));
    layer4_outputs(1443) <= (layer3_outputs(695)) or (layer3_outputs(4823));
    layer4_outputs(1444) <= not(layer3_outputs(5742)) or (layer3_outputs(6086));
    layer4_outputs(1445) <= not(layer3_outputs(5130));
    layer4_outputs(1446) <= '0';
    layer4_outputs(1447) <= not((layer3_outputs(4837)) xor (layer3_outputs(4061)));
    layer4_outputs(1448) <= '0';
    layer4_outputs(1449) <= layer3_outputs(7442);
    layer4_outputs(1450) <= not((layer3_outputs(955)) and (layer3_outputs(3263)));
    layer4_outputs(1451) <= not(layer3_outputs(2851));
    layer4_outputs(1452) <= not((layer3_outputs(6512)) or (layer3_outputs(5137)));
    layer4_outputs(1453) <= (layer3_outputs(422)) and not (layer3_outputs(50));
    layer4_outputs(1454) <= layer3_outputs(1464);
    layer4_outputs(1455) <= not(layer3_outputs(4834)) or (layer3_outputs(5537));
    layer4_outputs(1456) <= not((layer3_outputs(2143)) and (layer3_outputs(4907)));
    layer4_outputs(1457) <= not((layer3_outputs(3756)) and (layer3_outputs(1607)));
    layer4_outputs(1458) <= (layer3_outputs(3829)) and not (layer3_outputs(3656));
    layer4_outputs(1459) <= not(layer3_outputs(2969)) or (layer3_outputs(3286));
    layer4_outputs(1460) <= layer3_outputs(4474);
    layer4_outputs(1461) <= not((layer3_outputs(1058)) xor (layer3_outputs(7615)));
    layer4_outputs(1462) <= not((layer3_outputs(5563)) or (layer3_outputs(2639)));
    layer4_outputs(1463) <= not(layer3_outputs(6304));
    layer4_outputs(1464) <= not(layer3_outputs(2480));
    layer4_outputs(1465) <= not(layer3_outputs(6429));
    layer4_outputs(1466) <= not((layer3_outputs(5551)) xor (layer3_outputs(6583)));
    layer4_outputs(1467) <= (layer3_outputs(3165)) xor (layer3_outputs(864));
    layer4_outputs(1468) <= not(layer3_outputs(4593));
    layer4_outputs(1469) <= not((layer3_outputs(3884)) or (layer3_outputs(5529)));
    layer4_outputs(1470) <= not(layer3_outputs(445));
    layer4_outputs(1471) <= not(layer3_outputs(1467)) or (layer3_outputs(5781));
    layer4_outputs(1472) <= (layer3_outputs(898)) and not (layer3_outputs(948));
    layer4_outputs(1473) <= (layer3_outputs(2493)) and not (layer3_outputs(2361));
    layer4_outputs(1474) <= '1';
    layer4_outputs(1475) <= '0';
    layer4_outputs(1476) <= (layer3_outputs(6145)) or (layer3_outputs(2308));
    layer4_outputs(1477) <= layer3_outputs(5916);
    layer4_outputs(1478) <= not(layer3_outputs(846));
    layer4_outputs(1479) <= not(layer3_outputs(2424));
    layer4_outputs(1480) <= not(layer3_outputs(1789));
    layer4_outputs(1481) <= (layer3_outputs(3570)) or (layer3_outputs(3851));
    layer4_outputs(1482) <= (layer3_outputs(4183)) and (layer3_outputs(1297));
    layer4_outputs(1483) <= not(layer3_outputs(695));
    layer4_outputs(1484) <= layer3_outputs(374);
    layer4_outputs(1485) <= not(layer3_outputs(4129));
    layer4_outputs(1486) <= not(layer3_outputs(627)) or (layer3_outputs(6211));
    layer4_outputs(1487) <= layer3_outputs(7607);
    layer4_outputs(1488) <= layer3_outputs(111);
    layer4_outputs(1489) <= (layer3_outputs(1160)) and not (layer3_outputs(864));
    layer4_outputs(1490) <= layer3_outputs(2269);
    layer4_outputs(1491) <= (layer3_outputs(1753)) or (layer3_outputs(2983));
    layer4_outputs(1492) <= (layer3_outputs(5974)) and not (layer3_outputs(5174));
    layer4_outputs(1493) <= layer3_outputs(6524);
    layer4_outputs(1494) <= (layer3_outputs(706)) and not (layer3_outputs(245));
    layer4_outputs(1495) <= not((layer3_outputs(6135)) xor (layer3_outputs(1949)));
    layer4_outputs(1496) <= not(layer3_outputs(500));
    layer4_outputs(1497) <= (layer3_outputs(1736)) and (layer3_outputs(2171));
    layer4_outputs(1498) <= not(layer3_outputs(1893));
    layer4_outputs(1499) <= (layer3_outputs(4609)) and (layer3_outputs(1796));
    layer4_outputs(1500) <= not(layer3_outputs(353)) or (layer3_outputs(1502));
    layer4_outputs(1501) <= '0';
    layer4_outputs(1502) <= (layer3_outputs(362)) and not (layer3_outputs(6252));
    layer4_outputs(1503) <= layer3_outputs(6635);
    layer4_outputs(1504) <= not(layer3_outputs(3381));
    layer4_outputs(1505) <= (layer3_outputs(5389)) and (layer3_outputs(2173));
    layer4_outputs(1506) <= not((layer3_outputs(4262)) and (layer3_outputs(6054)));
    layer4_outputs(1507) <= (layer3_outputs(453)) and (layer3_outputs(5660));
    layer4_outputs(1508) <= (layer3_outputs(4582)) or (layer3_outputs(2511));
    layer4_outputs(1509) <= (layer3_outputs(6086)) and not (layer3_outputs(1433));
    layer4_outputs(1510) <= (layer3_outputs(1832)) and not (layer3_outputs(6836));
    layer4_outputs(1511) <= (layer3_outputs(1272)) and (layer3_outputs(1976));
    layer4_outputs(1512) <= layer3_outputs(6152);
    layer4_outputs(1513) <= layer3_outputs(981);
    layer4_outputs(1514) <= not(layer3_outputs(2235));
    layer4_outputs(1515) <= not(layer3_outputs(2756));
    layer4_outputs(1516) <= layer3_outputs(3456);
    layer4_outputs(1517) <= not((layer3_outputs(4315)) xor (layer3_outputs(2881)));
    layer4_outputs(1518) <= not((layer3_outputs(4944)) xor (layer3_outputs(882)));
    layer4_outputs(1519) <= not((layer3_outputs(3414)) or (layer3_outputs(850)));
    layer4_outputs(1520) <= not(layer3_outputs(783));
    layer4_outputs(1521) <= layer3_outputs(7473);
    layer4_outputs(1522) <= '0';
    layer4_outputs(1523) <= (layer3_outputs(1288)) and not (layer3_outputs(107));
    layer4_outputs(1524) <= layer3_outputs(905);
    layer4_outputs(1525) <= not(layer3_outputs(1134));
    layer4_outputs(1526) <= layer3_outputs(4546);
    layer4_outputs(1527) <= not((layer3_outputs(607)) or (layer3_outputs(7282)));
    layer4_outputs(1528) <= (layer3_outputs(1821)) and not (layer3_outputs(3180));
    layer4_outputs(1529) <= (layer3_outputs(7319)) xor (layer3_outputs(4862));
    layer4_outputs(1530) <= not(layer3_outputs(4939));
    layer4_outputs(1531) <= not(layer3_outputs(152)) or (layer3_outputs(39));
    layer4_outputs(1532) <= layer3_outputs(3495);
    layer4_outputs(1533) <= not(layer3_outputs(5307));
    layer4_outputs(1534) <= '1';
    layer4_outputs(1535) <= (layer3_outputs(4885)) and not (layer3_outputs(4539));
    layer4_outputs(1536) <= (layer3_outputs(7119)) and not (layer3_outputs(4896));
    layer4_outputs(1537) <= '0';
    layer4_outputs(1538) <= (layer3_outputs(576)) and (layer3_outputs(3685));
    layer4_outputs(1539) <= '1';
    layer4_outputs(1540) <= (layer3_outputs(3093)) and not (layer3_outputs(3447));
    layer4_outputs(1541) <= not(layer3_outputs(3815));
    layer4_outputs(1542) <= not((layer3_outputs(7411)) xor (layer3_outputs(1430)));
    layer4_outputs(1543) <= layer3_outputs(5488);
    layer4_outputs(1544) <= (layer3_outputs(999)) and (layer3_outputs(6371));
    layer4_outputs(1545) <= layer3_outputs(1183);
    layer4_outputs(1546) <= not(layer3_outputs(5296));
    layer4_outputs(1547) <= not(layer3_outputs(6955)) or (layer3_outputs(2681));
    layer4_outputs(1548) <= (layer3_outputs(4436)) or (layer3_outputs(7412));
    layer4_outputs(1549) <= '0';
    layer4_outputs(1550) <= not(layer3_outputs(2486)) or (layer3_outputs(4471));
    layer4_outputs(1551) <= layer3_outputs(1119);
    layer4_outputs(1552) <= layer3_outputs(583);
    layer4_outputs(1553) <= '1';
    layer4_outputs(1554) <= layer3_outputs(6115);
    layer4_outputs(1555) <= (layer3_outputs(1543)) and (layer3_outputs(4347));
    layer4_outputs(1556) <= not(layer3_outputs(108));
    layer4_outputs(1557) <= layer3_outputs(4305);
    layer4_outputs(1558) <= not(layer3_outputs(4467));
    layer4_outputs(1559) <= (layer3_outputs(5404)) and (layer3_outputs(1058));
    layer4_outputs(1560) <= (layer3_outputs(2731)) and not (layer3_outputs(7165));
    layer4_outputs(1561) <= not(layer3_outputs(1222)) or (layer3_outputs(6085));
    layer4_outputs(1562) <= not(layer3_outputs(4504));
    layer4_outputs(1563) <= not(layer3_outputs(3462)) or (layer3_outputs(3095));
    layer4_outputs(1564) <= (layer3_outputs(1174)) xor (layer3_outputs(2694));
    layer4_outputs(1565) <= not((layer3_outputs(5732)) xor (layer3_outputs(1814)));
    layer4_outputs(1566) <= not(layer3_outputs(2524)) or (layer3_outputs(6059));
    layer4_outputs(1567) <= not((layer3_outputs(815)) xor (layer3_outputs(2395)));
    layer4_outputs(1568) <= layer3_outputs(1042);
    layer4_outputs(1569) <= (layer3_outputs(2300)) xor (layer3_outputs(1143));
    layer4_outputs(1570) <= not((layer3_outputs(5424)) or (layer3_outputs(5207)));
    layer4_outputs(1571) <= not(layer3_outputs(4075)) or (layer3_outputs(3960));
    layer4_outputs(1572) <= layer3_outputs(1294);
    layer4_outputs(1573) <= '0';
    layer4_outputs(1574) <= '0';
    layer4_outputs(1575) <= layer3_outputs(4964);
    layer4_outputs(1576) <= (layer3_outputs(7653)) or (layer3_outputs(4718));
    layer4_outputs(1577) <= not(layer3_outputs(7622)) or (layer3_outputs(491));
    layer4_outputs(1578) <= (layer3_outputs(5782)) or (layer3_outputs(5977));
    layer4_outputs(1579) <= not((layer3_outputs(4584)) or (layer3_outputs(6007)));
    layer4_outputs(1580) <= not((layer3_outputs(1088)) or (layer3_outputs(1211)));
    layer4_outputs(1581) <= '1';
    layer4_outputs(1582) <= (layer3_outputs(5467)) and (layer3_outputs(6810));
    layer4_outputs(1583) <= not(layer3_outputs(3969)) or (layer3_outputs(2301));
    layer4_outputs(1584) <= not((layer3_outputs(383)) and (layer3_outputs(5252)));
    layer4_outputs(1585) <= not(layer3_outputs(3697)) or (layer3_outputs(7618));
    layer4_outputs(1586) <= not(layer3_outputs(6824)) or (layer3_outputs(6428));
    layer4_outputs(1587) <= not(layer3_outputs(2737));
    layer4_outputs(1588) <= layer3_outputs(2200);
    layer4_outputs(1589) <= not(layer3_outputs(1251));
    layer4_outputs(1590) <= not(layer3_outputs(857)) or (layer3_outputs(7600));
    layer4_outputs(1591) <= layer3_outputs(2943);
    layer4_outputs(1592) <= layer3_outputs(6935);
    layer4_outputs(1593) <= (layer3_outputs(1317)) and not (layer3_outputs(6363));
    layer4_outputs(1594) <= not(layer3_outputs(6375)) or (layer3_outputs(43));
    layer4_outputs(1595) <= (layer3_outputs(4487)) or (layer3_outputs(1811));
    layer4_outputs(1596) <= not(layer3_outputs(7339)) or (layer3_outputs(3433));
    layer4_outputs(1597) <= not((layer3_outputs(2291)) and (layer3_outputs(1074)));
    layer4_outputs(1598) <= '1';
    layer4_outputs(1599) <= layer3_outputs(21);
    layer4_outputs(1600) <= layer3_outputs(2544);
    layer4_outputs(1601) <= not((layer3_outputs(3608)) and (layer3_outputs(4838)));
    layer4_outputs(1602) <= not((layer3_outputs(364)) xor (layer3_outputs(5998)));
    layer4_outputs(1603) <= not(layer3_outputs(1749));
    layer4_outputs(1604) <= layer3_outputs(313);
    layer4_outputs(1605) <= not(layer3_outputs(178)) or (layer3_outputs(6976));
    layer4_outputs(1606) <= not(layer3_outputs(2949));
    layer4_outputs(1607) <= not(layer3_outputs(4452));
    layer4_outputs(1608) <= not((layer3_outputs(4029)) and (layer3_outputs(4591)));
    layer4_outputs(1609) <= not(layer3_outputs(4110));
    layer4_outputs(1610) <= layer3_outputs(4138);
    layer4_outputs(1611) <= layer3_outputs(1458);
    layer4_outputs(1612) <= (layer3_outputs(6970)) and not (layer3_outputs(3943));
    layer4_outputs(1613) <= layer3_outputs(7235);
    layer4_outputs(1614) <= not(layer3_outputs(7677));
    layer4_outputs(1615) <= (layer3_outputs(883)) and not (layer3_outputs(7076));
    layer4_outputs(1616) <= layer3_outputs(300);
    layer4_outputs(1617) <= layer3_outputs(3801);
    layer4_outputs(1618) <= not(layer3_outputs(1017)) or (layer3_outputs(2727));
    layer4_outputs(1619) <= not((layer3_outputs(1895)) xor (layer3_outputs(1754)));
    layer4_outputs(1620) <= not((layer3_outputs(6534)) and (layer3_outputs(4565)));
    layer4_outputs(1621) <= not(layer3_outputs(4894));
    layer4_outputs(1622) <= not((layer3_outputs(3311)) or (layer3_outputs(327)));
    layer4_outputs(1623) <= not(layer3_outputs(7657));
    layer4_outputs(1624) <= '1';
    layer4_outputs(1625) <= layer3_outputs(6777);
    layer4_outputs(1626) <= (layer3_outputs(5680)) and not (layer3_outputs(5565));
    layer4_outputs(1627) <= (layer3_outputs(3682)) and not (layer3_outputs(884));
    layer4_outputs(1628) <= not(layer3_outputs(3183));
    layer4_outputs(1629) <= (layer3_outputs(7105)) and (layer3_outputs(4108));
    layer4_outputs(1630) <= (layer3_outputs(2236)) and not (layer3_outputs(7150));
    layer4_outputs(1631) <= not(layer3_outputs(6673)) or (layer3_outputs(62));
    layer4_outputs(1632) <= layer3_outputs(2592);
    layer4_outputs(1633) <= (layer3_outputs(3943)) and (layer3_outputs(2909));
    layer4_outputs(1634) <= (layer3_outputs(5825)) and not (layer3_outputs(5067));
    layer4_outputs(1635) <= not((layer3_outputs(2534)) or (layer3_outputs(5566)));
    layer4_outputs(1636) <= not(layer3_outputs(3993)) or (layer3_outputs(1512));
    layer4_outputs(1637) <= (layer3_outputs(1355)) xor (layer3_outputs(5176));
    layer4_outputs(1638) <= not(layer3_outputs(5407)) or (layer3_outputs(2885));
    layer4_outputs(1639) <= (layer3_outputs(6869)) and not (layer3_outputs(2082));
    layer4_outputs(1640) <= not(layer3_outputs(4786)) or (layer3_outputs(6286));
    layer4_outputs(1641) <= layer3_outputs(1866);
    layer4_outputs(1642) <= not(layer3_outputs(7310)) or (layer3_outputs(1678));
    layer4_outputs(1643) <= layer3_outputs(6008);
    layer4_outputs(1644) <= not(layer3_outputs(3061));
    layer4_outputs(1645) <= not(layer3_outputs(1764)) or (layer3_outputs(6077));
    layer4_outputs(1646) <= (layer3_outputs(2415)) and not (layer3_outputs(3220));
    layer4_outputs(1647) <= not((layer3_outputs(5020)) and (layer3_outputs(6662)));
    layer4_outputs(1648) <= not(layer3_outputs(7286));
    layer4_outputs(1649) <= not((layer3_outputs(6390)) xor (layer3_outputs(7253)));
    layer4_outputs(1650) <= not(layer3_outputs(6692));
    layer4_outputs(1651) <= (layer3_outputs(3097)) or (layer3_outputs(2571));
    layer4_outputs(1652) <= layer3_outputs(2963);
    layer4_outputs(1653) <= (layer3_outputs(5960)) or (layer3_outputs(4554));
    layer4_outputs(1654) <= '1';
    layer4_outputs(1655) <= not(layer3_outputs(6341));
    layer4_outputs(1656) <= layer3_outputs(1389);
    layer4_outputs(1657) <= '0';
    layer4_outputs(1658) <= not((layer3_outputs(3323)) xor (layer3_outputs(6547)));
    layer4_outputs(1659) <= not(layer3_outputs(3663)) or (layer3_outputs(1304));
    layer4_outputs(1660) <= (layer3_outputs(4336)) or (layer3_outputs(4164));
    layer4_outputs(1661) <= not(layer3_outputs(7079)) or (layer3_outputs(2985));
    layer4_outputs(1662) <= not(layer3_outputs(2305)) or (layer3_outputs(578));
    layer4_outputs(1663) <= layer3_outputs(7201);
    layer4_outputs(1664) <= (layer3_outputs(5655)) and not (layer3_outputs(1034));
    layer4_outputs(1665) <= layer3_outputs(4079);
    layer4_outputs(1666) <= not(layer3_outputs(1494)) or (layer3_outputs(1365));
    layer4_outputs(1667) <= not(layer3_outputs(6819)) or (layer3_outputs(4607));
    layer4_outputs(1668) <= not(layer3_outputs(2935));
    layer4_outputs(1669) <= layer3_outputs(7591);
    layer4_outputs(1670) <= not(layer3_outputs(6589));
    layer4_outputs(1671) <= not(layer3_outputs(3144));
    layer4_outputs(1672) <= not(layer3_outputs(7587));
    layer4_outputs(1673) <= (layer3_outputs(6131)) or (layer3_outputs(5519));
    layer4_outputs(1674) <= not(layer3_outputs(1497));
    layer4_outputs(1675) <= not((layer3_outputs(2409)) and (layer3_outputs(6426)));
    layer4_outputs(1676) <= not(layer3_outputs(1200)) or (layer3_outputs(7679));
    layer4_outputs(1677) <= not(layer3_outputs(117)) or (layer3_outputs(6502));
    layer4_outputs(1678) <= layer3_outputs(5500);
    layer4_outputs(1679) <= not((layer3_outputs(7129)) and (layer3_outputs(3937)));
    layer4_outputs(1680) <= not((layer3_outputs(1107)) and (layer3_outputs(729)));
    layer4_outputs(1681) <= (layer3_outputs(7065)) and not (layer3_outputs(6984));
    layer4_outputs(1682) <= not(layer3_outputs(2774)) or (layer3_outputs(3953));
    layer4_outputs(1683) <= not(layer3_outputs(6362));
    layer4_outputs(1684) <= not(layer3_outputs(3171));
    layer4_outputs(1685) <= layer3_outputs(4776);
    layer4_outputs(1686) <= not(layer3_outputs(3856)) or (layer3_outputs(3660));
    layer4_outputs(1687) <= (layer3_outputs(4963)) and not (layer3_outputs(3540));
    layer4_outputs(1688) <= (layer3_outputs(1033)) and (layer3_outputs(2292));
    layer4_outputs(1689) <= (layer3_outputs(2526)) and not (layer3_outputs(4480));
    layer4_outputs(1690) <= (layer3_outputs(3875)) and not (layer3_outputs(3216));
    layer4_outputs(1691) <= layer3_outputs(2465);
    layer4_outputs(1692) <= not(layer3_outputs(4452));
    layer4_outputs(1693) <= (layer3_outputs(3372)) or (layer3_outputs(298));
    layer4_outputs(1694) <= '1';
    layer4_outputs(1695) <= not((layer3_outputs(7377)) or (layer3_outputs(87)));
    layer4_outputs(1696) <= not((layer3_outputs(7131)) and (layer3_outputs(5294)));
    layer4_outputs(1697) <= (layer3_outputs(5290)) or (layer3_outputs(866));
    layer4_outputs(1698) <= (layer3_outputs(2848)) xor (layer3_outputs(6867));
    layer4_outputs(1699) <= not(layer3_outputs(6982));
    layer4_outputs(1700) <= layer3_outputs(5205);
    layer4_outputs(1701) <= not(layer3_outputs(5444));
    layer4_outputs(1702) <= not(layer3_outputs(2382));
    layer4_outputs(1703) <= (layer3_outputs(2532)) xor (layer3_outputs(5980));
    layer4_outputs(1704) <= not(layer3_outputs(1025));
    layer4_outputs(1705) <= (layer3_outputs(2149)) and (layer3_outputs(1587));
    layer4_outputs(1706) <= not(layer3_outputs(596));
    layer4_outputs(1707) <= not(layer3_outputs(6747));
    layer4_outputs(1708) <= (layer3_outputs(6029)) xor (layer3_outputs(5574));
    layer4_outputs(1709) <= (layer3_outputs(2005)) and (layer3_outputs(4527));
    layer4_outputs(1710) <= not(layer3_outputs(7451)) or (layer3_outputs(35));
    layer4_outputs(1711) <= not((layer3_outputs(1138)) xor (layer3_outputs(2716)));
    layer4_outputs(1712) <= not((layer3_outputs(1769)) and (layer3_outputs(3970)));
    layer4_outputs(1713) <= not(layer3_outputs(5899));
    layer4_outputs(1714) <= (layer3_outputs(1173)) and not (layer3_outputs(1972));
    layer4_outputs(1715) <= not(layer3_outputs(6390));
    layer4_outputs(1716) <= not((layer3_outputs(2467)) and (layer3_outputs(3205)));
    layer4_outputs(1717) <= '1';
    layer4_outputs(1718) <= not((layer3_outputs(5615)) xor (layer3_outputs(2777)));
    layer4_outputs(1719) <= layer3_outputs(2959);
    layer4_outputs(1720) <= layer3_outputs(6523);
    layer4_outputs(1721) <= (layer3_outputs(4130)) and (layer3_outputs(2108));
    layer4_outputs(1722) <= (layer3_outputs(5777)) xor (layer3_outputs(4468));
    layer4_outputs(1723) <= (layer3_outputs(5473)) or (layer3_outputs(1842));
    layer4_outputs(1724) <= (layer3_outputs(4230)) or (layer3_outputs(306));
    layer4_outputs(1725) <= not((layer3_outputs(2705)) and (layer3_outputs(6762)));
    layer4_outputs(1726) <= (layer3_outputs(6727)) and (layer3_outputs(2767));
    layer4_outputs(1727) <= not(layer3_outputs(3572));
    layer4_outputs(1728) <= not(layer3_outputs(7311));
    layer4_outputs(1729) <= not(layer3_outputs(2449));
    layer4_outputs(1730) <= not((layer3_outputs(5897)) or (layer3_outputs(3395)));
    layer4_outputs(1731) <= layer3_outputs(2327);
    layer4_outputs(1732) <= (layer3_outputs(61)) and not (layer3_outputs(1621));
    layer4_outputs(1733) <= not((layer3_outputs(797)) and (layer3_outputs(6292)));
    layer4_outputs(1734) <= layer3_outputs(1336);
    layer4_outputs(1735) <= (layer3_outputs(5353)) and (layer3_outputs(7561));
    layer4_outputs(1736) <= (layer3_outputs(4053)) or (layer3_outputs(6011));
    layer4_outputs(1737) <= not((layer3_outputs(71)) and (layer3_outputs(4502)));
    layer4_outputs(1738) <= not(layer3_outputs(6239));
    layer4_outputs(1739) <= not(layer3_outputs(5528));
    layer4_outputs(1740) <= (layer3_outputs(3702)) xor (layer3_outputs(7531));
    layer4_outputs(1741) <= (layer3_outputs(3264)) and not (layer3_outputs(4932));
    layer4_outputs(1742) <= (layer3_outputs(3153)) or (layer3_outputs(611));
    layer4_outputs(1743) <= (layer3_outputs(1880)) or (layer3_outputs(3379));
    layer4_outputs(1744) <= (layer3_outputs(536)) xor (layer3_outputs(3465));
    layer4_outputs(1745) <= layer3_outputs(2169);
    layer4_outputs(1746) <= (layer3_outputs(7513)) or (layer3_outputs(259));
    layer4_outputs(1747) <= not((layer3_outputs(413)) and (layer3_outputs(1081)));
    layer4_outputs(1748) <= not(layer3_outputs(4292)) or (layer3_outputs(1578));
    layer4_outputs(1749) <= not(layer3_outputs(3136));
    layer4_outputs(1750) <= (layer3_outputs(4090)) and (layer3_outputs(6408));
    layer4_outputs(1751) <= not(layer3_outputs(68));
    layer4_outputs(1752) <= (layer3_outputs(6966)) and not (layer3_outputs(796));
    layer4_outputs(1753) <= not(layer3_outputs(3933)) or (layer3_outputs(934));
    layer4_outputs(1754) <= not(layer3_outputs(3617));
    layer4_outputs(1755) <= layer3_outputs(4302);
    layer4_outputs(1756) <= not((layer3_outputs(5316)) and (layer3_outputs(2317)));
    layer4_outputs(1757) <= layer3_outputs(3123);
    layer4_outputs(1758) <= layer3_outputs(731);
    layer4_outputs(1759) <= not(layer3_outputs(411)) or (layer3_outputs(4501));
    layer4_outputs(1760) <= layer3_outputs(2414);
    layer4_outputs(1761) <= (layer3_outputs(2995)) and (layer3_outputs(977));
    layer4_outputs(1762) <= layer3_outputs(5339);
    layer4_outputs(1763) <= (layer3_outputs(3282)) and (layer3_outputs(6997));
    layer4_outputs(1764) <= not(layer3_outputs(4045));
    layer4_outputs(1765) <= (layer3_outputs(3676)) and not (layer3_outputs(4394));
    layer4_outputs(1766) <= not(layer3_outputs(5904));
    layer4_outputs(1767) <= layer3_outputs(1657);
    layer4_outputs(1768) <= not((layer3_outputs(265)) xor (layer3_outputs(837)));
    layer4_outputs(1769) <= not((layer3_outputs(7612)) or (layer3_outputs(1851)));
    layer4_outputs(1770) <= layer3_outputs(1354);
    layer4_outputs(1771) <= not(layer3_outputs(5057));
    layer4_outputs(1772) <= layer3_outputs(2270);
    layer4_outputs(1773) <= not((layer3_outputs(2345)) xor (layer3_outputs(4683)));
    layer4_outputs(1774) <= layer3_outputs(384);
    layer4_outputs(1775) <= (layer3_outputs(4131)) and not (layer3_outputs(6092));
    layer4_outputs(1776) <= layer3_outputs(1253);
    layer4_outputs(1777) <= layer3_outputs(7427);
    layer4_outputs(1778) <= not(layer3_outputs(1825));
    layer4_outputs(1779) <= not(layer3_outputs(5313)) or (layer3_outputs(3343));
    layer4_outputs(1780) <= (layer3_outputs(6558)) and (layer3_outputs(6072));
    layer4_outputs(1781) <= not(layer3_outputs(2637)) or (layer3_outputs(3378));
    layer4_outputs(1782) <= layer3_outputs(5892);
    layer4_outputs(1783) <= (layer3_outputs(308)) and not (layer3_outputs(2373));
    layer4_outputs(1784) <= (layer3_outputs(5570)) and not (layer3_outputs(7260));
    layer4_outputs(1785) <= layer3_outputs(3411);
    layer4_outputs(1786) <= not(layer3_outputs(4318)) or (layer3_outputs(2951));
    layer4_outputs(1787) <= not(layer3_outputs(6892));
    layer4_outputs(1788) <= not(layer3_outputs(3497));
    layer4_outputs(1789) <= not(layer3_outputs(1532)) or (layer3_outputs(7658));
    layer4_outputs(1790) <= (layer3_outputs(1072)) and (layer3_outputs(1759));
    layer4_outputs(1791) <= layer3_outputs(1695);
    layer4_outputs(1792) <= (layer3_outputs(1837)) and not (layer3_outputs(5937));
    layer4_outputs(1793) <= layer3_outputs(4872);
    layer4_outputs(1794) <= not(layer3_outputs(6018));
    layer4_outputs(1795) <= not(layer3_outputs(2858));
    layer4_outputs(1796) <= (layer3_outputs(3047)) xor (layer3_outputs(840));
    layer4_outputs(1797) <= (layer3_outputs(3)) or (layer3_outputs(4417));
    layer4_outputs(1798) <= layer3_outputs(6557);
    layer4_outputs(1799) <= not((layer3_outputs(2220)) and (layer3_outputs(6665)));
    layer4_outputs(1800) <= not(layer3_outputs(6439));
    layer4_outputs(1801) <= not(layer3_outputs(5686));
    layer4_outputs(1802) <= not(layer3_outputs(3904));
    layer4_outputs(1803) <= not((layer3_outputs(6721)) xor (layer3_outputs(6727)));
    layer4_outputs(1804) <= not((layer3_outputs(123)) and (layer3_outputs(5531)));
    layer4_outputs(1805) <= not((layer3_outputs(5605)) and (layer3_outputs(1431)));
    layer4_outputs(1806) <= not(layer3_outputs(452)) or (layer3_outputs(3284));
    layer4_outputs(1807) <= (layer3_outputs(4288)) and not (layer3_outputs(3472));
    layer4_outputs(1808) <= layer3_outputs(5448);
    layer4_outputs(1809) <= layer3_outputs(3795);
    layer4_outputs(1810) <= not(layer3_outputs(791));
    layer4_outputs(1811) <= (layer3_outputs(3175)) xor (layer3_outputs(5719));
    layer4_outputs(1812) <= not(layer3_outputs(5643));
    layer4_outputs(1813) <= not(layer3_outputs(5365));
    layer4_outputs(1814) <= (layer3_outputs(2645)) and (layer3_outputs(5741));
    layer4_outputs(1815) <= (layer3_outputs(4684)) and not (layer3_outputs(1277));
    layer4_outputs(1816) <= (layer3_outputs(1582)) or (layer3_outputs(6982));
    layer4_outputs(1817) <= (layer3_outputs(5931)) and not (layer3_outputs(1855));
    layer4_outputs(1818) <= layer3_outputs(1928);
    layer4_outputs(1819) <= not(layer3_outputs(6038));
    layer4_outputs(1820) <= not(layer3_outputs(7203)) or (layer3_outputs(897));
    layer4_outputs(1821) <= not(layer3_outputs(6653)) or (layer3_outputs(5641));
    layer4_outputs(1822) <= not(layer3_outputs(4782)) or (layer3_outputs(7036));
    layer4_outputs(1823) <= (layer3_outputs(4004)) and not (layer3_outputs(6204));
    layer4_outputs(1824) <= not(layer3_outputs(3376));
    layer4_outputs(1825) <= not(layer3_outputs(1057));
    layer4_outputs(1826) <= not(layer3_outputs(6241));
    layer4_outputs(1827) <= not((layer3_outputs(7358)) and (layer3_outputs(3506)));
    layer4_outputs(1828) <= not(layer3_outputs(2889));
    layer4_outputs(1829) <= not(layer3_outputs(1177)) or (layer3_outputs(6611));
    layer4_outputs(1830) <= not(layer3_outputs(6044));
    layer4_outputs(1831) <= (layer3_outputs(7242)) and (layer3_outputs(1292));
    layer4_outputs(1832) <= '0';
    layer4_outputs(1833) <= not(layer3_outputs(7446));
    layer4_outputs(1834) <= (layer3_outputs(2913)) xor (layer3_outputs(4159));
    layer4_outputs(1835) <= not(layer3_outputs(5012)) or (layer3_outputs(4631));
    layer4_outputs(1836) <= not(layer3_outputs(7245)) or (layer3_outputs(3604));
    layer4_outputs(1837) <= (layer3_outputs(3210)) or (layer3_outputs(1374));
    layer4_outputs(1838) <= (layer3_outputs(2320)) and not (layer3_outputs(3377));
    layer4_outputs(1839) <= (layer3_outputs(4652)) and not (layer3_outputs(249));
    layer4_outputs(1840) <= '1';
    layer4_outputs(1841) <= not(layer3_outputs(7581)) or (layer3_outputs(6968));
    layer4_outputs(1842) <= layer3_outputs(6254);
    layer4_outputs(1843) <= not(layer3_outputs(4361)) or (layer3_outputs(3925));
    layer4_outputs(1844) <= layer3_outputs(2198);
    layer4_outputs(1845) <= not((layer3_outputs(6380)) xor (layer3_outputs(5283)));
    layer4_outputs(1846) <= not(layer3_outputs(1073));
    layer4_outputs(1847) <= (layer3_outputs(6986)) and (layer3_outputs(693));
    layer4_outputs(1848) <= not(layer3_outputs(3198));
    layer4_outputs(1849) <= layer3_outputs(1650);
    layer4_outputs(1850) <= '1';
    layer4_outputs(1851) <= (layer3_outputs(4168)) and (layer3_outputs(6034));
    layer4_outputs(1852) <= not((layer3_outputs(3511)) or (layer3_outputs(5270)));
    layer4_outputs(1853) <= not(layer3_outputs(5235));
    layer4_outputs(1854) <= not(layer3_outputs(1519));
    layer4_outputs(1855) <= not((layer3_outputs(2140)) and (layer3_outputs(2391)));
    layer4_outputs(1856) <= layer3_outputs(3600);
    layer4_outputs(1857) <= layer3_outputs(5995);
    layer4_outputs(1858) <= not((layer3_outputs(5055)) and (layer3_outputs(5455)));
    layer4_outputs(1859) <= (layer3_outputs(4229)) xor (layer3_outputs(795));
    layer4_outputs(1860) <= not(layer3_outputs(6598));
    layer4_outputs(1861) <= not((layer3_outputs(6117)) xor (layer3_outputs(3700)));
    layer4_outputs(1862) <= layer3_outputs(6428);
    layer4_outputs(1863) <= not(layer3_outputs(6403));
    layer4_outputs(1864) <= not(layer3_outputs(1900));
    layer4_outputs(1865) <= layer3_outputs(458);
    layer4_outputs(1866) <= not((layer3_outputs(3451)) and (layer3_outputs(3090)));
    layer4_outputs(1867) <= layer3_outputs(6105);
    layer4_outputs(1868) <= not(layer3_outputs(1384)) or (layer3_outputs(4490));
    layer4_outputs(1869) <= not(layer3_outputs(5184));
    layer4_outputs(1870) <= not(layer3_outputs(802));
    layer4_outputs(1871) <= (layer3_outputs(984)) and (layer3_outputs(5491));
    layer4_outputs(1872) <= not((layer3_outputs(3017)) or (layer3_outputs(6495)));
    layer4_outputs(1873) <= (layer3_outputs(3275)) and (layer3_outputs(294));
    layer4_outputs(1874) <= layer3_outputs(6470);
    layer4_outputs(1875) <= not(layer3_outputs(5834));
    layer4_outputs(1876) <= '0';
    layer4_outputs(1877) <= not((layer3_outputs(4244)) or (layer3_outputs(1115)));
    layer4_outputs(1878) <= (layer3_outputs(945)) and not (layer3_outputs(2686));
    layer4_outputs(1879) <= layer3_outputs(4339);
    layer4_outputs(1880) <= layer3_outputs(1594);
    layer4_outputs(1881) <= layer3_outputs(7085);
    layer4_outputs(1882) <= layer3_outputs(5118);
    layer4_outputs(1883) <= not(layer3_outputs(1071));
    layer4_outputs(1884) <= not(layer3_outputs(7199));
    layer4_outputs(1885) <= not((layer3_outputs(6127)) and (layer3_outputs(4044)));
    layer4_outputs(1886) <= '0';
    layer4_outputs(1887) <= layer3_outputs(4806);
    layer4_outputs(1888) <= (layer3_outputs(4158)) or (layer3_outputs(2505));
    layer4_outputs(1889) <= (layer3_outputs(4292)) xor (layer3_outputs(1259));
    layer4_outputs(1890) <= (layer3_outputs(4390)) and not (layer3_outputs(4519));
    layer4_outputs(1891) <= not(layer3_outputs(4460)) or (layer3_outputs(5651));
    layer4_outputs(1892) <= layer3_outputs(2752);
    layer4_outputs(1893) <= (layer3_outputs(5438)) or (layer3_outputs(5486));
    layer4_outputs(1894) <= layer3_outputs(5915);
    layer4_outputs(1895) <= (layer3_outputs(5578)) or (layer3_outputs(5292));
    layer4_outputs(1896) <= not(layer3_outputs(583));
    layer4_outputs(1897) <= not(layer3_outputs(817)) or (layer3_outputs(830));
    layer4_outputs(1898) <= (layer3_outputs(4052)) or (layer3_outputs(6122));
    layer4_outputs(1899) <= not(layer3_outputs(2958));
    layer4_outputs(1900) <= layer3_outputs(6350);
    layer4_outputs(1901) <= layer3_outputs(6975);
    layer4_outputs(1902) <= (layer3_outputs(5005)) and (layer3_outputs(2563));
    layer4_outputs(1903) <= not(layer3_outputs(1833));
    layer4_outputs(1904) <= '1';
    layer4_outputs(1905) <= (layer3_outputs(1550)) and not (layer3_outputs(491));
    layer4_outputs(1906) <= layer3_outputs(2528);
    layer4_outputs(1907) <= not((layer3_outputs(7236)) xor (layer3_outputs(3195)));
    layer4_outputs(1908) <= not((layer3_outputs(6804)) and (layer3_outputs(1751)));
    layer4_outputs(1909) <= not((layer3_outputs(543)) and (layer3_outputs(3906)));
    layer4_outputs(1910) <= '1';
    layer4_outputs(1911) <= not(layer3_outputs(7517));
    layer4_outputs(1912) <= layer3_outputs(4992);
    layer4_outputs(1913) <= (layer3_outputs(96)) or (layer3_outputs(2675));
    layer4_outputs(1914) <= not(layer3_outputs(4242));
    layer4_outputs(1915) <= (layer3_outputs(477)) and not (layer3_outputs(7068));
    layer4_outputs(1916) <= '1';
    layer4_outputs(1917) <= not(layer3_outputs(3179));
    layer4_outputs(1918) <= not(layer3_outputs(4780)) or (layer3_outputs(334));
    layer4_outputs(1919) <= layer3_outputs(939);
    layer4_outputs(1920) <= not(layer3_outputs(640)) or (layer3_outputs(4587));
    layer4_outputs(1921) <= not((layer3_outputs(1210)) or (layer3_outputs(4828)));
    layer4_outputs(1922) <= not((layer3_outputs(6607)) and (layer3_outputs(3193)));
    layer4_outputs(1923) <= '0';
    layer4_outputs(1924) <= not(layer3_outputs(5989)) or (layer3_outputs(5855));
    layer4_outputs(1925) <= not(layer3_outputs(3605));
    layer4_outputs(1926) <= '0';
    layer4_outputs(1927) <= (layer3_outputs(4618)) and not (layer3_outputs(4487));
    layer4_outputs(1928) <= layer3_outputs(5955);
    layer4_outputs(1929) <= (layer3_outputs(707)) and not (layer3_outputs(5698));
    layer4_outputs(1930) <= (layer3_outputs(426)) and not (layer3_outputs(1622));
    layer4_outputs(1931) <= not(layer3_outputs(4111)) or (layer3_outputs(6936));
    layer4_outputs(1932) <= not(layer3_outputs(2333)) or (layer3_outputs(2218));
    layer4_outputs(1933) <= (layer3_outputs(5571)) and (layer3_outputs(249));
    layer4_outputs(1934) <= not(layer3_outputs(2850)) or (layer3_outputs(6442));
    layer4_outputs(1935) <= not((layer3_outputs(7588)) and (layer3_outputs(2864)));
    layer4_outputs(1936) <= (layer3_outputs(6033)) and not (layer3_outputs(5927));
    layer4_outputs(1937) <= layer3_outputs(7602);
    layer4_outputs(1938) <= '1';
    layer4_outputs(1939) <= (layer3_outputs(666)) and (layer3_outputs(6933));
    layer4_outputs(1940) <= (layer3_outputs(1790)) and not (layer3_outputs(4895));
    layer4_outputs(1941) <= not(layer3_outputs(2501));
    layer4_outputs(1942) <= not((layer3_outputs(2434)) or (layer3_outputs(7121)));
    layer4_outputs(1943) <= layer3_outputs(5950);
    layer4_outputs(1944) <= (layer3_outputs(4950)) and (layer3_outputs(7471));
    layer4_outputs(1945) <= not(layer3_outputs(6866));
    layer4_outputs(1946) <= not(layer3_outputs(3239));
    layer4_outputs(1947) <= layer3_outputs(5018);
    layer4_outputs(1948) <= not(layer3_outputs(4129)) or (layer3_outputs(2679));
    layer4_outputs(1949) <= (layer3_outputs(6971)) xor (layer3_outputs(2525));
    layer4_outputs(1950) <= not((layer3_outputs(6176)) and (layer3_outputs(6416)));
    layer4_outputs(1951) <= (layer3_outputs(2176)) and not (layer3_outputs(1777));
    layer4_outputs(1952) <= not(layer3_outputs(3663));
    layer4_outputs(1953) <= (layer3_outputs(6021)) and (layer3_outputs(3630));
    layer4_outputs(1954) <= not(layer3_outputs(3112));
    layer4_outputs(1955) <= (layer3_outputs(3327)) and (layer3_outputs(6159));
    layer4_outputs(1956) <= layer3_outputs(4326);
    layer4_outputs(1957) <= not(layer3_outputs(6634));
    layer4_outputs(1958) <= (layer3_outputs(7652)) xor (layer3_outputs(6369));
    layer4_outputs(1959) <= layer3_outputs(2620);
    layer4_outputs(1960) <= not(layer3_outputs(1281));
    layer4_outputs(1961) <= '1';
    layer4_outputs(1962) <= not(layer3_outputs(6741));
    layer4_outputs(1963) <= layer3_outputs(5020);
    layer4_outputs(1964) <= not(layer3_outputs(5969)) or (layer3_outputs(363));
    layer4_outputs(1965) <= '0';
    layer4_outputs(1966) <= not((layer3_outputs(6773)) and (layer3_outputs(1719)));
    layer4_outputs(1967) <= layer3_outputs(6803);
    layer4_outputs(1968) <= (layer3_outputs(3296)) and not (layer3_outputs(1667));
    layer4_outputs(1969) <= not(layer3_outputs(412));
    layer4_outputs(1970) <= not((layer3_outputs(7533)) or (layer3_outputs(5911)));
    layer4_outputs(1971) <= layer3_outputs(653);
    layer4_outputs(1972) <= not((layer3_outputs(3796)) or (layer3_outputs(5314)));
    layer4_outputs(1973) <= not(layer3_outputs(2181));
    layer4_outputs(1974) <= not((layer3_outputs(2185)) or (layer3_outputs(2106)));
    layer4_outputs(1975) <= layer3_outputs(2339);
    layer4_outputs(1976) <= layer3_outputs(3083);
    layer4_outputs(1977) <= layer3_outputs(5299);
    layer4_outputs(1978) <= layer3_outputs(773);
    layer4_outputs(1979) <= not(layer3_outputs(5888));
    layer4_outputs(1980) <= not(layer3_outputs(1565));
    layer4_outputs(1981) <= not(layer3_outputs(5773)) or (layer3_outputs(862));
    layer4_outputs(1982) <= layer3_outputs(7396);
    layer4_outputs(1983) <= not((layer3_outputs(159)) and (layer3_outputs(2157)));
    layer4_outputs(1984) <= layer3_outputs(409);
    layer4_outputs(1985) <= not(layer3_outputs(3418));
    layer4_outputs(1986) <= layer3_outputs(1257);
    layer4_outputs(1987) <= not(layer3_outputs(955));
    layer4_outputs(1988) <= not(layer3_outputs(4435));
    layer4_outputs(1989) <= '1';
    layer4_outputs(1990) <= (layer3_outputs(4091)) xor (layer3_outputs(2809));
    layer4_outputs(1991) <= not(layer3_outputs(5695));
    layer4_outputs(1992) <= not((layer3_outputs(5339)) or (layer3_outputs(4636)));
    layer4_outputs(1993) <= (layer3_outputs(6931)) and not (layer3_outputs(4359));
    layer4_outputs(1994) <= (layer3_outputs(48)) and not (layer3_outputs(5369));
    layer4_outputs(1995) <= (layer3_outputs(7366)) or (layer3_outputs(4383));
    layer4_outputs(1996) <= layer3_outputs(7603);
    layer4_outputs(1997) <= not(layer3_outputs(4978));
    layer4_outputs(1998) <= (layer3_outputs(1336)) and not (layer3_outputs(3864));
    layer4_outputs(1999) <= layer3_outputs(459);
    layer4_outputs(2000) <= not(layer3_outputs(3516));
    layer4_outputs(2001) <= not(layer3_outputs(5096));
    layer4_outputs(2002) <= (layer3_outputs(4020)) xor (layer3_outputs(4157));
    layer4_outputs(2003) <= not(layer3_outputs(4206));
    layer4_outputs(2004) <= (layer3_outputs(6570)) and (layer3_outputs(2776));
    layer4_outputs(2005) <= not((layer3_outputs(2440)) and (layer3_outputs(262)));
    layer4_outputs(2006) <= not((layer3_outputs(6163)) or (layer3_outputs(6907)));
    layer4_outputs(2007) <= layer3_outputs(3117);
    layer4_outputs(2008) <= (layer3_outputs(5849)) xor (layer3_outputs(2119));
    layer4_outputs(2009) <= layer3_outputs(3230);
    layer4_outputs(2010) <= not(layer3_outputs(4672));
    layer4_outputs(2011) <= '0';
    layer4_outputs(2012) <= layer3_outputs(205);
    layer4_outputs(2013) <= (layer3_outputs(7366)) and not (layer3_outputs(2658));
    layer4_outputs(2014) <= not(layer3_outputs(4882));
    layer4_outputs(2015) <= layer3_outputs(2177);
    layer4_outputs(2016) <= '1';
    layer4_outputs(2017) <= (layer3_outputs(7040)) and not (layer3_outputs(7254));
    layer4_outputs(2018) <= '0';
    layer4_outputs(2019) <= not(layer3_outputs(1422)) or (layer3_outputs(6148));
    layer4_outputs(2020) <= not(layer3_outputs(3600));
    layer4_outputs(2021) <= (layer3_outputs(7678)) or (layer3_outputs(2161));
    layer4_outputs(2022) <= layer3_outputs(177);
    layer4_outputs(2023) <= not(layer3_outputs(985));
    layer4_outputs(2024) <= layer3_outputs(3602);
    layer4_outputs(2025) <= not((layer3_outputs(7056)) xor (layer3_outputs(4007)));
    layer4_outputs(2026) <= not((layer3_outputs(1302)) and (layer3_outputs(3006)));
    layer4_outputs(2027) <= (layer3_outputs(7568)) and not (layer3_outputs(7075));
    layer4_outputs(2028) <= not(layer3_outputs(2353));
    layer4_outputs(2029) <= not(layer3_outputs(192));
    layer4_outputs(2030) <= not(layer3_outputs(4852)) or (layer3_outputs(3030));
    layer4_outputs(2031) <= layer3_outputs(2306);
    layer4_outputs(2032) <= not(layer3_outputs(6023)) or (layer3_outputs(1429));
    layer4_outputs(2033) <= not((layer3_outputs(468)) or (layer3_outputs(7597)));
    layer4_outputs(2034) <= (layer3_outputs(1383)) and not (layer3_outputs(6303));
    layer4_outputs(2035) <= layer3_outputs(7494);
    layer4_outputs(2036) <= not((layer3_outputs(5959)) xor (layer3_outputs(122)));
    layer4_outputs(2037) <= (layer3_outputs(4224)) or (layer3_outputs(2138));
    layer4_outputs(2038) <= '1';
    layer4_outputs(2039) <= (layer3_outputs(929)) or (layer3_outputs(3052));
    layer4_outputs(2040) <= not((layer3_outputs(7448)) xor (layer3_outputs(6923)));
    layer4_outputs(2041) <= not(layer3_outputs(5298));
    layer4_outputs(2042) <= not((layer3_outputs(3262)) xor (layer3_outputs(4270)));
    layer4_outputs(2043) <= not(layer3_outputs(6791)) or (layer3_outputs(6941));
    layer4_outputs(2044) <= layer3_outputs(5645);
    layer4_outputs(2045) <= not((layer3_outputs(6001)) or (layer3_outputs(1273)));
    layer4_outputs(2046) <= (layer3_outputs(149)) and not (layer3_outputs(4399));
    layer4_outputs(2047) <= layer3_outputs(3568);
    layer4_outputs(2048) <= not(layer3_outputs(3775));
    layer4_outputs(2049) <= layer3_outputs(6516);
    layer4_outputs(2050) <= layer3_outputs(5838);
    layer4_outputs(2051) <= (layer3_outputs(5783)) and not (layer3_outputs(7317));
    layer4_outputs(2052) <= not(layer3_outputs(511)) or (layer3_outputs(4958));
    layer4_outputs(2053) <= not(layer3_outputs(804));
    layer4_outputs(2054) <= layer3_outputs(6940);
    layer4_outputs(2055) <= not((layer3_outputs(3986)) and (layer3_outputs(1413)));
    layer4_outputs(2056) <= (layer3_outputs(7271)) xor (layer3_outputs(5507));
    layer4_outputs(2057) <= not((layer3_outputs(2985)) xor (layer3_outputs(6260)));
    layer4_outputs(2058) <= (layer3_outputs(2750)) and not (layer3_outputs(462));
    layer4_outputs(2059) <= not(layer3_outputs(755));
    layer4_outputs(2060) <= (layer3_outputs(7171)) and (layer3_outputs(2383));
    layer4_outputs(2061) <= not(layer3_outputs(2285)) or (layer3_outputs(4581));
    layer4_outputs(2062) <= not((layer3_outputs(7562)) and (layer3_outputs(2334)));
    layer4_outputs(2063) <= layer3_outputs(7498);
    layer4_outputs(2064) <= not((layer3_outputs(3993)) and (layer3_outputs(5262)));
    layer4_outputs(2065) <= layer3_outputs(1672);
    layer4_outputs(2066) <= not((layer3_outputs(2186)) or (layer3_outputs(1919)));
    layer4_outputs(2067) <= not(layer3_outputs(2835)) or (layer3_outputs(1395));
    layer4_outputs(2068) <= layer3_outputs(2573);
    layer4_outputs(2069) <= not(layer3_outputs(6600)) or (layer3_outputs(1564));
    layer4_outputs(2070) <= '1';
    layer4_outputs(2071) <= (layer3_outputs(1504)) and not (layer3_outputs(6857));
    layer4_outputs(2072) <= not(layer3_outputs(285));
    layer4_outputs(2073) <= (layer3_outputs(7354)) and (layer3_outputs(4245));
    layer4_outputs(2074) <= (layer3_outputs(4980)) and not (layer3_outputs(2331));
    layer4_outputs(2075) <= not(layer3_outputs(7315));
    layer4_outputs(2076) <= (layer3_outputs(7019)) and not (layer3_outputs(5819));
    layer4_outputs(2077) <= not(layer3_outputs(2378));
    layer4_outputs(2078) <= layer3_outputs(5145);
    layer4_outputs(2079) <= (layer3_outputs(7556)) and (layer3_outputs(1388));
    layer4_outputs(2080) <= not(layer3_outputs(3696));
    layer4_outputs(2081) <= not((layer3_outputs(7467)) or (layer3_outputs(1095)));
    layer4_outputs(2082) <= not(layer3_outputs(6388));
    layer4_outputs(2083) <= layer3_outputs(3240);
    layer4_outputs(2084) <= (layer3_outputs(2954)) and not (layer3_outputs(329));
    layer4_outputs(2085) <= not(layer3_outputs(4152));
    layer4_outputs(2086) <= not(layer3_outputs(2162)) or (layer3_outputs(2351));
    layer4_outputs(2087) <= '0';
    layer4_outputs(2088) <= (layer3_outputs(3415)) and (layer3_outputs(7503));
    layer4_outputs(2089) <= layer3_outputs(5866);
    layer4_outputs(2090) <= '1';
    layer4_outputs(2091) <= not(layer3_outputs(2975));
    layer4_outputs(2092) <= (layer3_outputs(3001)) and not (layer3_outputs(508));
    layer4_outputs(2093) <= not(layer3_outputs(5483));
    layer4_outputs(2094) <= not(layer3_outputs(3319));
    layer4_outputs(2095) <= not(layer3_outputs(620));
    layer4_outputs(2096) <= layer3_outputs(6030);
    layer4_outputs(2097) <= (layer3_outputs(2053)) and not (layer3_outputs(4564));
    layer4_outputs(2098) <= not(layer3_outputs(1623)) or (layer3_outputs(1159));
    layer4_outputs(2099) <= (layer3_outputs(3707)) xor (layer3_outputs(5797));
    layer4_outputs(2100) <= not(layer3_outputs(1377));
    layer4_outputs(2101) <= not((layer3_outputs(5846)) xor (layer3_outputs(1699)));
    layer4_outputs(2102) <= not(layer3_outputs(3849));
    layer4_outputs(2103) <= not(layer3_outputs(4927));
    layer4_outputs(2104) <= not((layer3_outputs(2661)) and (layer3_outputs(527)));
    layer4_outputs(2105) <= not(layer3_outputs(1278));
    layer4_outputs(2106) <= layer3_outputs(5203);
    layer4_outputs(2107) <= not((layer3_outputs(950)) and (layer3_outputs(4182)));
    layer4_outputs(2108) <= not(layer3_outputs(4043));
    layer4_outputs(2109) <= layer3_outputs(3999);
    layer4_outputs(2110) <= (layer3_outputs(2846)) and (layer3_outputs(5802));
    layer4_outputs(2111) <= not((layer3_outputs(4505)) or (layer3_outputs(2878)));
    layer4_outputs(2112) <= (layer3_outputs(6508)) and not (layer3_outputs(7519));
    layer4_outputs(2113) <= layer3_outputs(11);
    layer4_outputs(2114) <= layer3_outputs(2778);
    layer4_outputs(2115) <= not((layer3_outputs(5274)) or (layer3_outputs(97)));
    layer4_outputs(2116) <= (layer3_outputs(1977)) xor (layer3_outputs(3278));
    layer4_outputs(2117) <= not(layer3_outputs(4235));
    layer4_outputs(2118) <= not(layer3_outputs(6173)) or (layer3_outputs(7029));
    layer4_outputs(2119) <= not(layer3_outputs(6175));
    layer4_outputs(2120) <= not(layer3_outputs(4915));
    layer4_outputs(2121) <= not(layer3_outputs(2314)) or (layer3_outputs(6040));
    layer4_outputs(2122) <= not(layer3_outputs(5068)) or (layer3_outputs(5458));
    layer4_outputs(2123) <= '0';
    layer4_outputs(2124) <= layer3_outputs(2290);
    layer4_outputs(2125) <= not((layer3_outputs(3739)) xor (layer3_outputs(1451)));
    layer4_outputs(2126) <= not((layer3_outputs(6720)) xor (layer3_outputs(371)));
    layer4_outputs(2127) <= layer3_outputs(3351);
    layer4_outputs(2128) <= '1';
    layer4_outputs(2129) <= (layer3_outputs(4722)) xor (layer3_outputs(3969));
    layer4_outputs(2130) <= not(layer3_outputs(6875));
    layer4_outputs(2131) <= layer3_outputs(3126);
    layer4_outputs(2132) <= layer3_outputs(4446);
    layer4_outputs(2133) <= not(layer3_outputs(3465));
    layer4_outputs(2134) <= not(layer3_outputs(7055));
    layer4_outputs(2135) <= not((layer3_outputs(259)) xor (layer3_outputs(5831)));
    layer4_outputs(2136) <= layer3_outputs(547);
    layer4_outputs(2137) <= not(layer3_outputs(248)) or (layer3_outputs(2557));
    layer4_outputs(2138) <= (layer3_outputs(6501)) xor (layer3_outputs(4321));
    layer4_outputs(2139) <= not((layer3_outputs(5372)) and (layer3_outputs(1197)));
    layer4_outputs(2140) <= not(layer3_outputs(7280));
    layer4_outputs(2141) <= not(layer3_outputs(5279));
    layer4_outputs(2142) <= (layer3_outputs(5486)) and (layer3_outputs(5104));
    layer4_outputs(2143) <= '0';
    layer4_outputs(2144) <= not((layer3_outputs(3765)) or (layer3_outputs(1108)));
    layer4_outputs(2145) <= layer3_outputs(6478);
    layer4_outputs(2146) <= layer3_outputs(5321);
    layer4_outputs(2147) <= (layer3_outputs(6918)) and not (layer3_outputs(4134));
    layer4_outputs(2148) <= (layer3_outputs(4795)) or (layer3_outputs(6446));
    layer4_outputs(2149) <= (layer3_outputs(2508)) or (layer3_outputs(2254));
    layer4_outputs(2150) <= not(layer3_outputs(959)) or (layer3_outputs(77));
    layer4_outputs(2151) <= (layer3_outputs(7078)) or (layer3_outputs(865));
    layer4_outputs(2152) <= not(layer3_outputs(7579));
    layer4_outputs(2153) <= '0';
    layer4_outputs(2154) <= (layer3_outputs(5121)) and (layer3_outputs(2914));
    layer4_outputs(2155) <= layer3_outputs(2277);
    layer4_outputs(2156) <= not(layer3_outputs(2547));
    layer4_outputs(2157) <= not(layer3_outputs(1997));
    layer4_outputs(2158) <= (layer3_outputs(1095)) or (layer3_outputs(664));
    layer4_outputs(2159) <= layer3_outputs(3596);
    layer4_outputs(2160) <= (layer3_outputs(3809)) and (layer3_outputs(1030));
    layer4_outputs(2161) <= '1';
    layer4_outputs(2162) <= layer3_outputs(3863);
    layer4_outputs(2163) <= not(layer3_outputs(6322));
    layer4_outputs(2164) <= not((layer3_outputs(4783)) xor (layer3_outputs(4)));
    layer4_outputs(2165) <= layer3_outputs(410);
    layer4_outputs(2166) <= (layer3_outputs(2989)) xor (layer3_outputs(4730));
    layer4_outputs(2167) <= not(layer3_outputs(1154));
    layer4_outputs(2168) <= not(layer3_outputs(1306));
    layer4_outputs(2169) <= layer3_outputs(1862);
    layer4_outputs(2170) <= not(layer3_outputs(1220)) or (layer3_outputs(1925));
    layer4_outputs(2171) <= (layer3_outputs(6445)) or (layer3_outputs(6335));
    layer4_outputs(2172) <= layer3_outputs(30);
    layer4_outputs(2173) <= '1';
    layer4_outputs(2174) <= (layer3_outputs(5264)) or (layer3_outputs(6486));
    layer4_outputs(2175) <= layer3_outputs(1601);
    layer4_outputs(2176) <= not(layer3_outputs(4612));
    layer4_outputs(2177) <= not((layer3_outputs(1158)) xor (layer3_outputs(1038)));
    layer4_outputs(2178) <= (layer3_outputs(5824)) xor (layer3_outputs(1875));
    layer4_outputs(2179) <= '0';
    layer4_outputs(2180) <= not(layer3_outputs(3927));
    layer4_outputs(2181) <= not(layer3_outputs(229)) or (layer3_outputs(5864));
    layer4_outputs(2182) <= layer3_outputs(3695);
    layer4_outputs(2183) <= '1';
    layer4_outputs(2184) <= not(layer3_outputs(822));
    layer4_outputs(2185) <= not((layer3_outputs(3529)) or (layer3_outputs(6829)));
    layer4_outputs(2186) <= (layer3_outputs(5809)) and (layer3_outputs(1811));
    layer4_outputs(2187) <= not((layer3_outputs(985)) and (layer3_outputs(3911)));
    layer4_outputs(2188) <= (layer3_outputs(3667)) and not (layer3_outputs(140));
    layer4_outputs(2189) <= not((layer3_outputs(6566)) xor (layer3_outputs(4748)));
    layer4_outputs(2190) <= (layer3_outputs(3809)) and (layer3_outputs(3437));
    layer4_outputs(2191) <= (layer3_outputs(2283)) xor (layer3_outputs(2735));
    layer4_outputs(2192) <= (layer3_outputs(1206)) and not (layer3_outputs(7413));
    layer4_outputs(2193) <= not((layer3_outputs(6307)) xor (layer3_outputs(6784)));
    layer4_outputs(2194) <= not((layer3_outputs(2531)) and (layer3_outputs(2875)));
    layer4_outputs(2195) <= (layer3_outputs(5258)) or (layer3_outputs(4650));
    layer4_outputs(2196) <= not(layer3_outputs(1330)) or (layer3_outputs(2506));
    layer4_outputs(2197) <= layer3_outputs(4800);
    layer4_outputs(2198) <= layer3_outputs(1419);
    layer4_outputs(2199) <= not(layer3_outputs(4260));
    layer4_outputs(2200) <= not(layer3_outputs(4843));
    layer4_outputs(2201) <= layer3_outputs(4083);
    layer4_outputs(2202) <= not(layer3_outputs(5767));
    layer4_outputs(2203) <= not((layer3_outputs(3396)) or (layer3_outputs(4223)));
    layer4_outputs(2204) <= (layer3_outputs(3430)) and not (layer3_outputs(7404));
    layer4_outputs(2205) <= (layer3_outputs(7117)) and not (layer3_outputs(5456));
    layer4_outputs(2206) <= not(layer3_outputs(5659));
    layer4_outputs(2207) <= layer3_outputs(3614);
    layer4_outputs(2208) <= not(layer3_outputs(5757)) or (layer3_outputs(2023));
    layer4_outputs(2209) <= layer3_outputs(1834);
    layer4_outputs(2210) <= not((layer3_outputs(2754)) or (layer3_outputs(5964)));
    layer4_outputs(2211) <= not(layer3_outputs(3694));
    layer4_outputs(2212) <= (layer3_outputs(5165)) and not (layer3_outputs(5337));
    layer4_outputs(2213) <= not((layer3_outputs(7218)) and (layer3_outputs(1240)));
    layer4_outputs(2214) <= (layer3_outputs(7166)) and not (layer3_outputs(83));
    layer4_outputs(2215) <= '1';
    layer4_outputs(2216) <= not((layer3_outputs(3109)) or (layer3_outputs(4851)));
    layer4_outputs(2217) <= not(layer3_outputs(2395)) or (layer3_outputs(6174));
    layer4_outputs(2218) <= not(layer3_outputs(1477)) or (layer3_outputs(1252));
    layer4_outputs(2219) <= not((layer3_outputs(7571)) and (layer3_outputs(3983)));
    layer4_outputs(2220) <= not(layer3_outputs(5325));
    layer4_outputs(2221) <= (layer3_outputs(3068)) and not (layer3_outputs(4175));
    layer4_outputs(2222) <= not(layer3_outputs(3819));
    layer4_outputs(2223) <= not(layer3_outputs(4879)) or (layer3_outputs(661));
    layer4_outputs(2224) <= not(layer3_outputs(2491));
    layer4_outputs(2225) <= (layer3_outputs(5636)) and not (layer3_outputs(7463));
    layer4_outputs(2226) <= not(layer3_outputs(6461));
    layer4_outputs(2227) <= not(layer3_outputs(4093));
    layer4_outputs(2228) <= (layer3_outputs(3423)) xor (layer3_outputs(4287));
    layer4_outputs(2229) <= not(layer3_outputs(2356));
    layer4_outputs(2230) <= not((layer3_outputs(2377)) or (layer3_outputs(5383)));
    layer4_outputs(2231) <= layer3_outputs(884);
    layer4_outputs(2232) <= not((layer3_outputs(3367)) and (layer3_outputs(7091)));
    layer4_outputs(2233) <= (layer3_outputs(2976)) and not (layer3_outputs(2827));
    layer4_outputs(2234) <= layer3_outputs(1482);
    layer4_outputs(2235) <= layer3_outputs(4832);
    layer4_outputs(2236) <= (layer3_outputs(6515)) and not (layer3_outputs(2182));
    layer4_outputs(2237) <= not((layer3_outputs(6402)) or (layer3_outputs(6082)));
    layer4_outputs(2238) <= layer3_outputs(2344);
    layer4_outputs(2239) <= not((layer3_outputs(4063)) and (layer3_outputs(3634)));
    layer4_outputs(2240) <= not(layer3_outputs(3364));
    layer4_outputs(2241) <= not(layer3_outputs(45));
    layer4_outputs(2242) <= (layer3_outputs(6552)) and not (layer3_outputs(3249));
    layer4_outputs(2243) <= not(layer3_outputs(1702));
    layer4_outputs(2244) <= (layer3_outputs(1332)) and not (layer3_outputs(2228));
    layer4_outputs(2245) <= (layer3_outputs(1406)) and (layer3_outputs(454));
    layer4_outputs(2246) <= layer3_outputs(4101);
    layer4_outputs(2247) <= not(layer3_outputs(3035)) or (layer3_outputs(3022));
    layer4_outputs(2248) <= not((layer3_outputs(7570)) or (layer3_outputs(5321)));
    layer4_outputs(2249) <= (layer3_outputs(5111)) and not (layer3_outputs(6389));
    layer4_outputs(2250) <= (layer3_outputs(1372)) or (layer3_outputs(1130));
    layer4_outputs(2251) <= not((layer3_outputs(1279)) or (layer3_outputs(5809)));
    layer4_outputs(2252) <= not(layer3_outputs(7508));
    layer4_outputs(2253) <= not(layer3_outputs(246));
    layer4_outputs(2254) <= (layer3_outputs(6631)) and (layer3_outputs(1312));
    layer4_outputs(2255) <= layer3_outputs(5903);
    layer4_outputs(2256) <= layer3_outputs(448);
    layer4_outputs(2257) <= not((layer3_outputs(3568)) and (layer3_outputs(3992)));
    layer4_outputs(2258) <= (layer3_outputs(802)) and not (layer3_outputs(6740));
    layer4_outputs(2259) <= not(layer3_outputs(6234));
    layer4_outputs(2260) <= (layer3_outputs(4686)) xor (layer3_outputs(2730));
    layer4_outputs(2261) <= not((layer3_outputs(4289)) and (layer3_outputs(2749)));
    layer4_outputs(2262) <= not(layer3_outputs(287));
    layer4_outputs(2263) <= not(layer3_outputs(4913)) or (layer3_outputs(859));
    layer4_outputs(2264) <= not(layer3_outputs(6567)) or (layer3_outputs(3088));
    layer4_outputs(2265) <= layer3_outputs(321);
    layer4_outputs(2266) <= (layer3_outputs(6532)) xor (layer3_outputs(13));
    layer4_outputs(2267) <= layer3_outputs(2159);
    layer4_outputs(2268) <= layer3_outputs(4513);
    layer4_outputs(2269) <= (layer3_outputs(4375)) and not (layer3_outputs(69));
    layer4_outputs(2270) <= not((layer3_outputs(1577)) and (layer3_outputs(128)));
    layer4_outputs(2271) <= not((layer3_outputs(2123)) and (layer3_outputs(5039)));
    layer4_outputs(2272) <= layer3_outputs(183);
    layer4_outputs(2273) <= not(layer3_outputs(4647));
    layer4_outputs(2274) <= not((layer3_outputs(6820)) and (layer3_outputs(4000)));
    layer4_outputs(2275) <= not((layer3_outputs(6352)) or (layer3_outputs(1652)));
    layer4_outputs(2276) <= (layer3_outputs(5347)) and not (layer3_outputs(1455));
    layer4_outputs(2277) <= layer3_outputs(3711);
    layer4_outputs(2278) <= not(layer3_outputs(1964)) or (layer3_outputs(295));
    layer4_outputs(2279) <= layer3_outputs(2005);
    layer4_outputs(2280) <= not(layer3_outputs(6301));
    layer4_outputs(2281) <= not(layer3_outputs(376));
    layer4_outputs(2282) <= layer3_outputs(594);
    layer4_outputs(2283) <= layer3_outputs(614);
    layer4_outputs(2284) <= not(layer3_outputs(3092)) or (layer3_outputs(3448));
    layer4_outputs(2285) <= not(layer3_outputs(7295));
    layer4_outputs(2286) <= not(layer3_outputs(4072));
    layer4_outputs(2287) <= not(layer3_outputs(3338)) or (layer3_outputs(1605));
    layer4_outputs(2288) <= (layer3_outputs(2246)) and not (layer3_outputs(6227));
    layer4_outputs(2289) <= layer3_outputs(5814);
    layer4_outputs(2290) <= not(layer3_outputs(1932));
    layer4_outputs(2291) <= not((layer3_outputs(312)) and (layer3_outputs(4040)));
    layer4_outputs(2292) <= layer3_outputs(261);
    layer4_outputs(2293) <= layer3_outputs(7286);
    layer4_outputs(2294) <= (layer3_outputs(1800)) and not (layer3_outputs(1755));
    layer4_outputs(2295) <= layer3_outputs(3492);
    layer4_outputs(2296) <= layer3_outputs(4853);
    layer4_outputs(2297) <= layer3_outputs(6034);
    layer4_outputs(2298) <= not(layer3_outputs(3992));
    layer4_outputs(2299) <= not(layer3_outputs(2163)) or (layer3_outputs(1822));
    layer4_outputs(2300) <= not((layer3_outputs(3882)) or (layer3_outputs(1542)));
    layer4_outputs(2301) <= not(layer3_outputs(541));
    layer4_outputs(2302) <= (layer3_outputs(1549)) and not (layer3_outputs(7051));
    layer4_outputs(2303) <= layer3_outputs(6559);
    layer4_outputs(2304) <= '1';
    layer4_outputs(2305) <= not(layer3_outputs(2528));
    layer4_outputs(2306) <= layer3_outputs(5862);
    layer4_outputs(2307) <= not((layer3_outputs(527)) and (layer3_outputs(3651)));
    layer4_outputs(2308) <= not((layer3_outputs(4124)) and (layer3_outputs(6663)));
    layer4_outputs(2309) <= '0';
    layer4_outputs(2310) <= layer3_outputs(7197);
    layer4_outputs(2311) <= not(layer3_outputs(6097));
    layer4_outputs(2312) <= not(layer3_outputs(1521)) or (layer3_outputs(6300));
    layer4_outputs(2313) <= not(layer3_outputs(4803)) or (layer3_outputs(7500));
    layer4_outputs(2314) <= layer3_outputs(7371);
    layer4_outputs(2315) <= not(layer3_outputs(5099));
    layer4_outputs(2316) <= layer3_outputs(2902);
    layer4_outputs(2317) <= not(layer3_outputs(6084)) or (layer3_outputs(3036));
    layer4_outputs(2318) <= not(layer3_outputs(3851)) or (layer3_outputs(2514));
    layer4_outputs(2319) <= not(layer3_outputs(4577)) or (layer3_outputs(5787));
    layer4_outputs(2320) <= not((layer3_outputs(3642)) and (layer3_outputs(6128)));
    layer4_outputs(2321) <= not((layer3_outputs(6905)) and (layer3_outputs(181)));
    layer4_outputs(2322) <= layer3_outputs(2422);
    layer4_outputs(2323) <= not((layer3_outputs(6522)) or (layer3_outputs(6815)));
    layer4_outputs(2324) <= (layer3_outputs(2696)) or (layer3_outputs(7291));
    layer4_outputs(2325) <= layer3_outputs(6222);
    layer4_outputs(2326) <= not(layer3_outputs(7378));
    layer4_outputs(2327) <= not(layer3_outputs(6218));
    layer4_outputs(2328) <= (layer3_outputs(1737)) and not (layer3_outputs(5932));
    layer4_outputs(2329) <= not(layer3_outputs(4028)) or (layer3_outputs(3412));
    layer4_outputs(2330) <= layer3_outputs(3168);
    layer4_outputs(2331) <= layer3_outputs(1099);
    layer4_outputs(2332) <= not(layer3_outputs(3543)) or (layer3_outputs(5940));
    layer4_outputs(2333) <= not(layer3_outputs(2336));
    layer4_outputs(2334) <= layer3_outputs(4226);
    layer4_outputs(2335) <= (layer3_outputs(5823)) or (layer3_outputs(2862));
    layer4_outputs(2336) <= not(layer3_outputs(471)) or (layer3_outputs(1438));
    layer4_outputs(2337) <= not(layer3_outputs(7258)) or (layer3_outputs(4024));
    layer4_outputs(2338) <= not(layer3_outputs(712));
    layer4_outputs(2339) <= not(layer3_outputs(5269));
    layer4_outputs(2340) <= not(layer3_outputs(3900));
    layer4_outputs(2341) <= not((layer3_outputs(3635)) and (layer3_outputs(2974)));
    layer4_outputs(2342) <= not(layer3_outputs(2762));
    layer4_outputs(2343) <= (layer3_outputs(7270)) xor (layer3_outputs(3979));
    layer4_outputs(2344) <= not(layer3_outputs(1540));
    layer4_outputs(2345) <= not(layer3_outputs(1070));
    layer4_outputs(2346) <= not(layer3_outputs(2032));
    layer4_outputs(2347) <= layer3_outputs(6098);
    layer4_outputs(2348) <= not((layer3_outputs(4432)) and (layer3_outputs(2457)));
    layer4_outputs(2349) <= not(layer3_outputs(6186));
    layer4_outputs(2350) <= not((layer3_outputs(5683)) xor (layer3_outputs(4092)));
    layer4_outputs(2351) <= not(layer3_outputs(982));
    layer4_outputs(2352) <= '0';
    layer4_outputs(2353) <= (layer3_outputs(1794)) and not (layer3_outputs(4335));
    layer4_outputs(2354) <= layer3_outputs(132);
    layer4_outputs(2355) <= (layer3_outputs(5913)) and not (layer3_outputs(3222));
    layer4_outputs(2356) <= not(layer3_outputs(7083)) or (layer3_outputs(2113));
    layer4_outputs(2357) <= not((layer3_outputs(7528)) or (layer3_outputs(6112)));
    layer4_outputs(2358) <= (layer3_outputs(7273)) or (layer3_outputs(4323));
    layer4_outputs(2359) <= (layer3_outputs(4796)) and (layer3_outputs(721));
    layer4_outputs(2360) <= not((layer3_outputs(6580)) or (layer3_outputs(4489)));
    layer4_outputs(2361) <= '1';
    layer4_outputs(2362) <= layer3_outputs(75);
    layer4_outputs(2363) <= layer3_outputs(922);
    layer4_outputs(2364) <= (layer3_outputs(1134)) and not (layer3_outputs(6752));
    layer4_outputs(2365) <= (layer3_outputs(5476)) and not (layer3_outputs(4804));
    layer4_outputs(2366) <= not(layer3_outputs(4902));
    layer4_outputs(2367) <= (layer3_outputs(4450)) or (layer3_outputs(5323));
    layer4_outputs(2368) <= layer3_outputs(5406);
    layer4_outputs(2369) <= (layer3_outputs(6301)) and (layer3_outputs(3561));
    layer4_outputs(2370) <= layer3_outputs(5774);
    layer4_outputs(2371) <= '0';
    layer4_outputs(2372) <= not(layer3_outputs(7339));
    layer4_outputs(2373) <= not((layer3_outputs(5601)) or (layer3_outputs(5567)));
    layer4_outputs(2374) <= not(layer3_outputs(6242));
    layer4_outputs(2375) <= '1';
    layer4_outputs(2376) <= layer3_outputs(5395);
    layer4_outputs(2377) <= (layer3_outputs(7463)) or (layer3_outputs(6629));
    layer4_outputs(2378) <= not(layer3_outputs(5829));
    layer4_outputs(2379) <= not((layer3_outputs(7149)) or (layer3_outputs(274)));
    layer4_outputs(2380) <= layer3_outputs(6484);
    layer4_outputs(2381) <= (layer3_outputs(1782)) and not (layer3_outputs(1325));
    layer4_outputs(2382) <= (layer3_outputs(4867)) or (layer3_outputs(3200));
    layer4_outputs(2383) <= layer3_outputs(6273);
    layer4_outputs(2384) <= not(layer3_outputs(3542));
    layer4_outputs(2385) <= layer3_outputs(2401);
    layer4_outputs(2386) <= (layer3_outputs(2209)) and (layer3_outputs(4102));
    layer4_outputs(2387) <= not(layer3_outputs(528));
    layer4_outputs(2388) <= not(layer3_outputs(1180));
    layer4_outputs(2389) <= not(layer3_outputs(4264)) or (layer3_outputs(3803));
    layer4_outputs(2390) <= not((layer3_outputs(6474)) or (layer3_outputs(33)));
    layer4_outputs(2391) <= (layer3_outputs(3121)) and not (layer3_outputs(381));
    layer4_outputs(2392) <= not(layer3_outputs(6757));
    layer4_outputs(2393) <= (layer3_outputs(337)) and (layer3_outputs(1364));
    layer4_outputs(2394) <= layer3_outputs(6759);
    layer4_outputs(2395) <= not(layer3_outputs(2579));
    layer4_outputs(2396) <= not(layer3_outputs(4889));
    layer4_outputs(2397) <= not((layer3_outputs(3773)) xor (layer3_outputs(767)));
    layer4_outputs(2398) <= '0';
    layer4_outputs(2399) <= layer3_outputs(7178);
    layer4_outputs(2400) <= (layer3_outputs(2503)) and (layer3_outputs(6802));
    layer4_outputs(2401) <= not(layer3_outputs(2630));
    layer4_outputs(2402) <= (layer3_outputs(3682)) or (layer3_outputs(4300));
    layer4_outputs(2403) <= not(layer3_outputs(1987));
    layer4_outputs(2404) <= (layer3_outputs(7457)) and (layer3_outputs(1360));
    layer4_outputs(2405) <= (layer3_outputs(4490)) and not (layer3_outputs(5244));
    layer4_outputs(2406) <= (layer3_outputs(142)) and (layer3_outputs(3401));
    layer4_outputs(2407) <= layer3_outputs(2021);
    layer4_outputs(2408) <= layer3_outputs(7318);
    layer4_outputs(2409) <= not(layer3_outputs(6184)) or (layer3_outputs(6417));
    layer4_outputs(2410) <= not((layer3_outputs(5848)) and (layer3_outputs(5090)));
    layer4_outputs(2411) <= not((layer3_outputs(156)) or (layer3_outputs(2107)));
    layer4_outputs(2412) <= (layer3_outputs(6295)) or (layer3_outputs(433));
    layer4_outputs(2413) <= not(layer3_outputs(4186));
    layer4_outputs(2414) <= not(layer3_outputs(5978)) or (layer3_outputs(6256));
    layer4_outputs(2415) <= layer3_outputs(5026);
    layer4_outputs(2416) <= not(layer3_outputs(7371));
    layer4_outputs(2417) <= layer3_outputs(1460);
    layer4_outputs(2418) <= not(layer3_outputs(1114));
    layer4_outputs(2419) <= (layer3_outputs(5844)) and (layer3_outputs(1280));
    layer4_outputs(2420) <= layer3_outputs(3591);
    layer4_outputs(2421) <= not(layer3_outputs(1518)) or (layer3_outputs(3732));
    layer4_outputs(2422) <= not(layer3_outputs(7593));
    layer4_outputs(2423) <= (layer3_outputs(544)) and not (layer3_outputs(1178));
    layer4_outputs(2424) <= (layer3_outputs(1942)) and (layer3_outputs(1469));
    layer4_outputs(2425) <= not(layer3_outputs(4810));
    layer4_outputs(2426) <= not((layer3_outputs(4206)) or (layer3_outputs(5044)));
    layer4_outputs(2427) <= (layer3_outputs(4171)) and not (layer3_outputs(2351));
    layer4_outputs(2428) <= (layer3_outputs(1925)) or (layer3_outputs(1994));
    layer4_outputs(2429) <= not((layer3_outputs(782)) and (layer3_outputs(5646)));
    layer4_outputs(2430) <= not(layer3_outputs(3298));
    layer4_outputs(2431) <= (layer3_outputs(2456)) and not (layer3_outputs(6481));
    layer4_outputs(2432) <= not(layer3_outputs(7656));
    layer4_outputs(2433) <= (layer3_outputs(80)) and not (layer3_outputs(4641));
    layer4_outputs(2434) <= layer3_outputs(1156);
    layer4_outputs(2435) <= (layer3_outputs(3228)) or (layer3_outputs(5535));
    layer4_outputs(2436) <= (layer3_outputs(1701)) and not (layer3_outputs(1322));
    layer4_outputs(2437) <= not((layer3_outputs(758)) xor (layer3_outputs(6761)));
    layer4_outputs(2438) <= (layer3_outputs(6346)) or (layer3_outputs(1676));
    layer4_outputs(2439) <= (layer3_outputs(6439)) xor (layer3_outputs(209));
    layer4_outputs(2440) <= not(layer3_outputs(4629));
    layer4_outputs(2441) <= layer3_outputs(415);
    layer4_outputs(2442) <= not((layer3_outputs(7561)) and (layer3_outputs(5779)));
    layer4_outputs(2443) <= not(layer3_outputs(2179));
    layer4_outputs(2444) <= (layer3_outputs(2136)) and not (layer3_outputs(2274));
    layer4_outputs(2445) <= layer3_outputs(4383);
    layer4_outputs(2446) <= not((layer3_outputs(6457)) xor (layer3_outputs(2929)));
    layer4_outputs(2447) <= (layer3_outputs(2414)) and not (layer3_outputs(1244));
    layer4_outputs(2448) <= not((layer3_outputs(2420)) xor (layer3_outputs(3504)));
    layer4_outputs(2449) <= not(layer3_outputs(5675));
    layer4_outputs(2450) <= not(layer3_outputs(2577)) or (layer3_outputs(5736));
    layer4_outputs(2451) <= '0';
    layer4_outputs(2452) <= not((layer3_outputs(2033)) and (layer3_outputs(2648)));
    layer4_outputs(2453) <= layer3_outputs(4908);
    layer4_outputs(2454) <= not(layer3_outputs(2497));
    layer4_outputs(2455) <= layer3_outputs(1810);
    layer4_outputs(2456) <= layer3_outputs(1531);
    layer4_outputs(2457) <= not(layer3_outputs(648)) or (layer3_outputs(4397));
    layer4_outputs(2458) <= (layer3_outputs(1510)) and (layer3_outputs(3869));
    layer4_outputs(2459) <= not(layer3_outputs(2728)) or (layer3_outputs(6895));
    layer4_outputs(2460) <= not(layer3_outputs(2973)) or (layer3_outputs(4314));
    layer4_outputs(2461) <= '0';
    layer4_outputs(2462) <= layer3_outputs(6456);
    layer4_outputs(2463) <= layer3_outputs(6685);
    layer4_outputs(2464) <= (layer3_outputs(46)) and not (layer3_outputs(240));
    layer4_outputs(2465) <= '0';
    layer4_outputs(2466) <= (layer3_outputs(6160)) xor (layer3_outputs(2764));
    layer4_outputs(2467) <= layer3_outputs(631);
    layer4_outputs(2468) <= not(layer3_outputs(4772));
    layer4_outputs(2469) <= not(layer3_outputs(7007));
    layer4_outputs(2470) <= not((layer3_outputs(516)) and (layer3_outputs(2388)));
    layer4_outputs(2471) <= not((layer3_outputs(999)) or (layer3_outputs(5308)));
    layer4_outputs(2472) <= '1';
    layer4_outputs(2473) <= not(layer3_outputs(2906)) or (layer3_outputs(3454));
    layer4_outputs(2474) <= (layer3_outputs(4028)) and (layer3_outputs(4030));
    layer4_outputs(2475) <= layer3_outputs(391);
    layer4_outputs(2476) <= '0';
    layer4_outputs(2477) <= layer3_outputs(2814);
    layer4_outputs(2478) <= (layer3_outputs(369)) xor (layer3_outputs(110));
    layer4_outputs(2479) <= '0';
    layer4_outputs(2480) <= (layer3_outputs(3667)) xor (layer3_outputs(713));
    layer4_outputs(2481) <= not(layer3_outputs(5758));
    layer4_outputs(2482) <= layer3_outputs(434);
    layer4_outputs(2483) <= not(layer3_outputs(6021)) or (layer3_outputs(6574));
    layer4_outputs(2484) <= layer3_outputs(2856);
    layer4_outputs(2485) <= (layer3_outputs(4830)) and (layer3_outputs(4691));
    layer4_outputs(2486) <= layer3_outputs(209);
    layer4_outputs(2487) <= (layer3_outputs(365)) or (layer3_outputs(6964));
    layer4_outputs(2488) <= not(layer3_outputs(673)) or (layer3_outputs(7009));
    layer4_outputs(2489) <= not(layer3_outputs(6266));
    layer4_outputs(2490) <= not(layer3_outputs(5857));
    layer4_outputs(2491) <= '1';
    layer4_outputs(2492) <= not((layer3_outputs(3635)) and (layer3_outputs(4778)));
    layer4_outputs(2493) <= not(layer3_outputs(4241)) or (layer3_outputs(3322));
    layer4_outputs(2494) <= layer3_outputs(966);
    layer4_outputs(2495) <= layer3_outputs(3133);
    layer4_outputs(2496) <= not(layer3_outputs(718));
    layer4_outputs(2497) <= layer3_outputs(5268);
    layer4_outputs(2498) <= layer3_outputs(6622);
    layer4_outputs(2499) <= not(layer3_outputs(6517));
    layer4_outputs(2500) <= not(layer3_outputs(3294)) or (layer3_outputs(1747));
    layer4_outputs(2501) <= not(layer3_outputs(4547));
    layer4_outputs(2502) <= (layer3_outputs(1588)) and not (layer3_outputs(7220));
    layer4_outputs(2503) <= '0';
    layer4_outputs(2504) <= (layer3_outputs(495)) xor (layer3_outputs(4984));
    layer4_outputs(2505) <= (layer3_outputs(2310)) and not (layer3_outputs(4833));
    layer4_outputs(2506) <= (layer3_outputs(32)) and not (layer3_outputs(3556));
    layer4_outputs(2507) <= (layer3_outputs(7180)) and not (layer3_outputs(3643));
    layer4_outputs(2508) <= layer3_outputs(5277);
    layer4_outputs(2509) <= (layer3_outputs(7431)) and (layer3_outputs(2358));
    layer4_outputs(2510) <= not(layer3_outputs(6376)) or (layer3_outputs(2865));
    layer4_outputs(2511) <= not(layer3_outputs(3074));
    layer4_outputs(2512) <= not((layer3_outputs(5472)) or (layer3_outputs(4735)));
    layer4_outputs(2513) <= (layer3_outputs(4036)) and not (layer3_outputs(4971));
    layer4_outputs(2514) <= (layer3_outputs(1903)) and not (layer3_outputs(5552));
    layer4_outputs(2515) <= (layer3_outputs(6809)) and not (layer3_outputs(1008));
    layer4_outputs(2516) <= (layer3_outputs(6200)) and (layer3_outputs(3182));
    layer4_outputs(2517) <= not(layer3_outputs(490)) or (layer3_outputs(446));
    layer4_outputs(2518) <= (layer3_outputs(4658)) or (layer3_outputs(1298));
    layer4_outputs(2519) <= layer3_outputs(2879);
    layer4_outputs(2520) <= not(layer3_outputs(4148));
    layer4_outputs(2521) <= not(layer3_outputs(7548)) or (layer3_outputs(3611));
    layer4_outputs(2522) <= (layer3_outputs(860)) and (layer3_outputs(343));
    layer4_outputs(2523) <= not((layer3_outputs(7000)) or (layer3_outputs(6975)));
    layer4_outputs(2524) <= layer3_outputs(5546);
    layer4_outputs(2525) <= not((layer3_outputs(4493)) and (layer3_outputs(3981)));
    layer4_outputs(2526) <= layer3_outputs(1998);
    layer4_outputs(2527) <= not(layer3_outputs(4768));
    layer4_outputs(2528) <= not((layer3_outputs(6810)) xor (layer3_outputs(4252)));
    layer4_outputs(2529) <= layer3_outputs(2139);
    layer4_outputs(2530) <= layer3_outputs(4588);
    layer4_outputs(2531) <= not((layer3_outputs(7297)) xor (layer3_outputs(6804)));
    layer4_outputs(2532) <= not(layer3_outputs(1890));
    layer4_outputs(2533) <= not(layer3_outputs(7311));
    layer4_outputs(2534) <= '1';
    layer4_outputs(2535) <= not((layer3_outputs(2915)) and (layer3_outputs(6657)));
    layer4_outputs(2536) <= layer3_outputs(1861);
    layer4_outputs(2537) <= layer3_outputs(1510);
    layer4_outputs(2538) <= (layer3_outputs(2522)) and (layer3_outputs(1289));
    layer4_outputs(2539) <= layer3_outputs(872);
    layer4_outputs(2540) <= '1';
    layer4_outputs(2541) <= not((layer3_outputs(6574)) or (layer3_outputs(3028)));
    layer4_outputs(2542) <= layer3_outputs(6240);
    layer4_outputs(2543) <= not(layer3_outputs(2931)) or (layer3_outputs(1716));
    layer4_outputs(2544) <= not(layer3_outputs(309));
    layer4_outputs(2545) <= not(layer3_outputs(6430));
    layer4_outputs(2546) <= (layer3_outputs(5931)) and not (layer3_outputs(2258));
    layer4_outputs(2547) <= not(layer3_outputs(3263)) or (layer3_outputs(3271));
    layer4_outputs(2548) <= (layer3_outputs(5633)) and (layer3_outputs(3044));
    layer4_outputs(2549) <= not((layer3_outputs(4807)) or (layer3_outputs(5589)));
    layer4_outputs(2550) <= layer3_outputs(2145);
    layer4_outputs(2551) <= (layer3_outputs(997)) and not (layer3_outputs(234));
    layer4_outputs(2552) <= layer3_outputs(3156);
    layer4_outputs(2553) <= not((layer3_outputs(6915)) or (layer3_outputs(3947)));
    layer4_outputs(2554) <= (layer3_outputs(4909)) and (layer3_outputs(1568));
    layer4_outputs(2555) <= layer3_outputs(6978);
    layer4_outputs(2556) <= not(layer3_outputs(1982));
    layer4_outputs(2557) <= (layer3_outputs(5879)) and not (layer3_outputs(3098));
    layer4_outputs(2558) <= not((layer3_outputs(4763)) xor (layer3_outputs(2486)));
    layer4_outputs(2559) <= not(layer3_outputs(6488));
    layer4_outputs(2560) <= (layer3_outputs(7400)) and (layer3_outputs(6849));
    layer4_outputs(2561) <= not(layer3_outputs(5109));
    layer4_outputs(2562) <= (layer3_outputs(6625)) and not (layer3_outputs(245));
    layer4_outputs(2563) <= layer3_outputs(2421);
    layer4_outputs(2564) <= not(layer3_outputs(4380));
    layer4_outputs(2565) <= not(layer3_outputs(7662)) or (layer3_outputs(2305));
    layer4_outputs(2566) <= not(layer3_outputs(4704)) or (layer3_outputs(5225));
    layer4_outputs(2567) <= '0';
    layer4_outputs(2568) <= (layer3_outputs(2558)) and not (layer3_outputs(5865));
    layer4_outputs(2569) <= '1';
    layer4_outputs(2570) <= (layer3_outputs(7129)) and (layer3_outputs(2768));
    layer4_outputs(2571) <= not(layer3_outputs(2951)) or (layer3_outputs(6427));
    layer4_outputs(2572) <= (layer3_outputs(1922)) and not (layer3_outputs(1207));
    layer4_outputs(2573) <= layer3_outputs(2664);
    layer4_outputs(2574) <= layer3_outputs(2787);
    layer4_outputs(2575) <= not(layer3_outputs(7388));
    layer4_outputs(2576) <= not(layer3_outputs(1186)) or (layer3_outputs(1465));
    layer4_outputs(2577) <= '1';
    layer4_outputs(2578) <= not(layer3_outputs(5183));
    layer4_outputs(2579) <= not((layer3_outputs(3363)) xor (layer3_outputs(2467)));
    layer4_outputs(2580) <= layer3_outputs(6863);
    layer4_outputs(2581) <= (layer3_outputs(3657)) and not (layer3_outputs(6140));
    layer4_outputs(2582) <= not(layer3_outputs(4894));
    layer4_outputs(2583) <= (layer3_outputs(2714)) or (layer3_outputs(1514));
    layer4_outputs(2584) <= (layer3_outputs(425)) and not (layer3_outputs(7043));
    layer4_outputs(2585) <= (layer3_outputs(2376)) or (layer3_outputs(6152));
    layer4_outputs(2586) <= (layer3_outputs(5060)) and (layer3_outputs(6288));
    layer4_outputs(2587) <= layer3_outputs(6314);
    layer4_outputs(2588) <= not((layer3_outputs(3076)) and (layer3_outputs(5423)));
    layer4_outputs(2589) <= layer3_outputs(4442);
    layer4_outputs(2590) <= layer3_outputs(5610);
    layer4_outputs(2591) <= (layer3_outputs(6032)) and not (layer3_outputs(4661));
    layer4_outputs(2592) <= layer3_outputs(3835);
    layer4_outputs(2593) <= not((layer3_outputs(5764)) or (layer3_outputs(6223)));
    layer4_outputs(2594) <= not((layer3_outputs(1663)) or (layer3_outputs(5539)));
    layer4_outputs(2595) <= layer3_outputs(7315);
    layer4_outputs(2596) <= (layer3_outputs(2286)) and not (layer3_outputs(752));
    layer4_outputs(2597) <= (layer3_outputs(1858)) and not (layer3_outputs(3217));
    layer4_outputs(2598) <= layer3_outputs(4757);
    layer4_outputs(2599) <= layer3_outputs(4610);
    layer4_outputs(2600) <= layer3_outputs(675);
    layer4_outputs(2601) <= (layer3_outputs(6902)) and not (layer3_outputs(6297));
    layer4_outputs(2602) <= not(layer3_outputs(3355)) or (layer3_outputs(3983));
    layer4_outputs(2603) <= (layer3_outputs(6590)) and not (layer3_outputs(970));
    layer4_outputs(2604) <= not(layer3_outputs(1468));
    layer4_outputs(2605) <= not(layer3_outputs(3466));
    layer4_outputs(2606) <= layer3_outputs(5238);
    layer4_outputs(2607) <= not((layer3_outputs(6472)) and (layer3_outputs(6545)));
    layer4_outputs(2608) <= not((layer3_outputs(2691)) and (layer3_outputs(663)));
    layer4_outputs(2609) <= layer3_outputs(2175);
    layer4_outputs(2610) <= not(layer3_outputs(5387));
    layer4_outputs(2611) <= not((layer3_outputs(5679)) or (layer3_outputs(3733)));
    layer4_outputs(2612) <= not((layer3_outputs(7072)) xor (layer3_outputs(5251)));
    layer4_outputs(2613) <= not(layer3_outputs(4381));
    layer4_outputs(2614) <= not(layer3_outputs(7320)) or (layer3_outputs(3423));
    layer4_outputs(2615) <= layer3_outputs(3571);
    layer4_outputs(2616) <= (layer3_outputs(6582)) and (layer3_outputs(924));
    layer4_outputs(2617) <= layer3_outputs(188);
    layer4_outputs(2618) <= not((layer3_outputs(3016)) or (layer3_outputs(7448)));
    layer4_outputs(2619) <= layer3_outputs(1153);
    layer4_outputs(2620) <= not(layer3_outputs(1970)) or (layer3_outputs(5606));
    layer4_outputs(2621) <= (layer3_outputs(7415)) and not (layer3_outputs(4624));
    layer4_outputs(2622) <= not(layer3_outputs(1616));
    layer4_outputs(2623) <= not((layer3_outputs(3450)) xor (layer3_outputs(5794)));
    layer4_outputs(2624) <= '1';
    layer4_outputs(2625) <= (layer3_outputs(5404)) and (layer3_outputs(4956));
    layer4_outputs(2626) <= not((layer3_outputs(7290)) and (layer3_outputs(919)));
    layer4_outputs(2627) <= not((layer3_outputs(5733)) and (layer3_outputs(6455)));
    layer4_outputs(2628) <= not(layer3_outputs(5668));
    layer4_outputs(2629) <= '0';
    layer4_outputs(2630) <= (layer3_outputs(5340)) and not (layer3_outputs(2054));
    layer4_outputs(2631) <= not(layer3_outputs(2670));
    layer4_outputs(2632) <= not((layer3_outputs(5171)) xor (layer3_outputs(407)));
    layer4_outputs(2633) <= layer3_outputs(3539);
    layer4_outputs(2634) <= layer3_outputs(4222);
    layer4_outputs(2635) <= (layer3_outputs(1024)) and not (layer3_outputs(1613));
    layer4_outputs(2636) <= not((layer3_outputs(7097)) xor (layer3_outputs(5607)));
    layer4_outputs(2637) <= not((layer3_outputs(4666)) and (layer3_outputs(6360)));
    layer4_outputs(2638) <= not(layer3_outputs(7558));
    layer4_outputs(2639) <= not((layer3_outputs(5148)) or (layer3_outputs(1746)));
    layer4_outputs(2640) <= not(layer3_outputs(2020));
    layer4_outputs(2641) <= not((layer3_outputs(6829)) and (layer3_outputs(5511)));
    layer4_outputs(2642) <= layer3_outputs(5422);
    layer4_outputs(2643) <= not(layer3_outputs(6520)) or (layer3_outputs(2891));
    layer4_outputs(2644) <= (layer3_outputs(3243)) and (layer3_outputs(3314));
    layer4_outputs(2645) <= (layer3_outputs(5414)) or (layer3_outputs(6968));
    layer4_outputs(2646) <= not((layer3_outputs(3520)) and (layer3_outputs(7670)));
    layer4_outputs(2647) <= '1';
    layer4_outputs(2648) <= (layer3_outputs(3045)) xor (layer3_outputs(6283));
    layer4_outputs(2649) <= not(layer3_outputs(3023));
    layer4_outputs(2650) <= (layer3_outputs(7481)) and not (layer3_outputs(1320));
    layer4_outputs(2651) <= (layer3_outputs(1995)) or (layer3_outputs(7543));
    layer4_outputs(2652) <= layer3_outputs(7028);
    layer4_outputs(2653) <= (layer3_outputs(4434)) xor (layer3_outputs(1002));
    layer4_outputs(2654) <= not(layer3_outputs(6116));
    layer4_outputs(2655) <= not((layer3_outputs(4526)) and (layer3_outputs(991)));
    layer4_outputs(2656) <= layer3_outputs(2319);
    layer4_outputs(2657) <= (layer3_outputs(6937)) and (layer3_outputs(621));
    layer4_outputs(2658) <= layer3_outputs(6200);
    layer4_outputs(2659) <= layer3_outputs(5440);
    layer4_outputs(2660) <= not(layer3_outputs(647)) or (layer3_outputs(7529));
    layer4_outputs(2661) <= not(layer3_outputs(643));
    layer4_outputs(2662) <= (layer3_outputs(7121)) or (layer3_outputs(3088));
    layer4_outputs(2663) <= layer3_outputs(4218);
    layer4_outputs(2664) <= not(layer3_outputs(636)) or (layer3_outputs(3065));
    layer4_outputs(2665) <= (layer3_outputs(2552)) or (layer3_outputs(5088));
    layer4_outputs(2666) <= not(layer3_outputs(356)) or (layer3_outputs(6527));
    layer4_outputs(2667) <= layer3_outputs(4207);
    layer4_outputs(2668) <= (layer3_outputs(2190)) xor (layer3_outputs(2250));
    layer4_outputs(2669) <= (layer3_outputs(3000)) and (layer3_outputs(4461));
    layer4_outputs(2670) <= (layer3_outputs(6856)) xor (layer3_outputs(2229));
    layer4_outputs(2671) <= (layer3_outputs(2938)) and (layer3_outputs(1509));
    layer4_outputs(2672) <= (layer3_outputs(7542)) and not (layer3_outputs(7493));
    layer4_outputs(2673) <= not(layer3_outputs(3479));
    layer4_outputs(2674) <= layer3_outputs(2096);
    layer4_outputs(2675) <= not(layer3_outputs(1290));
    layer4_outputs(2676) <= (layer3_outputs(5457)) and not (layer3_outputs(3625));
    layer4_outputs(2677) <= not(layer3_outputs(873)) or (layer3_outputs(216));
    layer4_outputs(2678) <= layer3_outputs(3670);
    layer4_outputs(2679) <= '0';
    layer4_outputs(2680) <= not(layer3_outputs(6280));
    layer4_outputs(2681) <= layer3_outputs(1505);
    layer4_outputs(2682) <= not(layer3_outputs(5126));
    layer4_outputs(2683) <= not(layer3_outputs(4532));
    layer4_outputs(2684) <= '0';
    layer4_outputs(2685) <= layer3_outputs(4296);
    layer4_outputs(2686) <= not(layer3_outputs(3790));
    layer4_outputs(2687) <= not(layer3_outputs(7249)) or (layer3_outputs(4932));
    layer4_outputs(2688) <= '0';
    layer4_outputs(2689) <= (layer3_outputs(4213)) and (layer3_outputs(3525));
    layer4_outputs(2690) <= not((layer3_outputs(101)) xor (layer3_outputs(3487)));
    layer4_outputs(2691) <= not(layer3_outputs(7133)) or (layer3_outputs(228));
    layer4_outputs(2692) <= not(layer3_outputs(3312));
    layer4_outputs(2693) <= '1';
    layer4_outputs(2694) <= layer3_outputs(1485);
    layer4_outputs(2695) <= '1';
    layer4_outputs(2696) <= '0';
    layer4_outputs(2697) <= (layer3_outputs(949)) and not (layer3_outputs(7096));
    layer4_outputs(2698) <= not((layer3_outputs(3083)) and (layer3_outputs(5041)));
    layer4_outputs(2699) <= not(layer3_outputs(5512));
    layer4_outputs(2700) <= (layer3_outputs(5791)) and (layer3_outputs(3791));
    layer4_outputs(2701) <= not((layer3_outputs(6815)) or (layer3_outputs(2359)));
    layer4_outputs(2702) <= not((layer3_outputs(267)) xor (layer3_outputs(5107)));
    layer4_outputs(2703) <= not(layer3_outputs(520)) or (layer3_outputs(6493));
    layer4_outputs(2704) <= not(layer3_outputs(1547));
    layer4_outputs(2705) <= not(layer3_outputs(1755)) or (layer3_outputs(6780));
    layer4_outputs(2706) <= (layer3_outputs(1441)) or (layer3_outputs(196));
    layer4_outputs(2707) <= not((layer3_outputs(6214)) or (layer3_outputs(1778)));
    layer4_outputs(2708) <= not(layer3_outputs(2695));
    layer4_outputs(2709) <= not((layer3_outputs(6755)) and (layer3_outputs(813)));
    layer4_outputs(2710) <= (layer3_outputs(3964)) and not (layer3_outputs(1371));
    layer4_outputs(2711) <= not((layer3_outputs(5229)) or (layer3_outputs(7475)));
    layer4_outputs(2712) <= not((layer3_outputs(5918)) or (layer3_outputs(2807)));
    layer4_outputs(2713) <= not(layer3_outputs(3130));
    layer4_outputs(2714) <= not((layer3_outputs(6120)) or (layer3_outputs(4934)));
    layer4_outputs(2715) <= (layer3_outputs(5683)) and not (layer3_outputs(2516));
    layer4_outputs(2716) <= layer3_outputs(3500);
    layer4_outputs(2717) <= not((layer3_outputs(1106)) and (layer3_outputs(6807)));
    layer4_outputs(2718) <= not((layer3_outputs(5265)) or (layer3_outputs(2717)));
    layer4_outputs(2719) <= layer3_outputs(3242);
    layer4_outputs(2720) <= (layer3_outputs(4285)) and (layer3_outputs(2659));
    layer4_outputs(2721) <= not(layer3_outputs(7632)) or (layer3_outputs(351));
    layer4_outputs(2722) <= not(layer3_outputs(4110));
    layer4_outputs(2723) <= '0';
    layer4_outputs(2724) <= '1';
    layer4_outputs(2725) <= (layer3_outputs(2381)) or (layer3_outputs(4830));
    layer4_outputs(2726) <= layer3_outputs(7035);
    layer4_outputs(2727) <= not(layer3_outputs(1956));
    layer4_outputs(2728) <= not(layer3_outputs(3038));
    layer4_outputs(2729) <= not((layer3_outputs(1625)) or (layer3_outputs(6703)));
    layer4_outputs(2730) <= layer3_outputs(1195);
    layer4_outputs(2731) <= not(layer3_outputs(574)) or (layer3_outputs(2141));
    layer4_outputs(2732) <= (layer3_outputs(5954)) and not (layer3_outputs(5227));
    layer4_outputs(2733) <= not(layer3_outputs(7421)) or (layer3_outputs(859));
    layer4_outputs(2734) <= '0';
    layer4_outputs(2735) <= not(layer3_outputs(3717));
    layer4_outputs(2736) <= not(layer3_outputs(3077));
    layer4_outputs(2737) <= layer3_outputs(1862);
    layer4_outputs(2738) <= (layer3_outputs(4963)) and not (layer3_outputs(4643));
    layer4_outputs(2739) <= (layer3_outputs(5252)) or (layer3_outputs(4310));
    layer4_outputs(2740) <= (layer3_outputs(7334)) and (layer3_outputs(3808));
    layer4_outputs(2741) <= not(layer3_outputs(4314));
    layer4_outputs(2742) <= not((layer3_outputs(3013)) or (layer3_outputs(3620)));
    layer4_outputs(2743) <= (layer3_outputs(1124)) and not (layer3_outputs(4212));
    layer4_outputs(2744) <= not(layer3_outputs(710)) or (layer3_outputs(3919));
    layer4_outputs(2745) <= not((layer3_outputs(2334)) or (layer3_outputs(2576)));
    layer4_outputs(2746) <= not((layer3_outputs(4585)) or (layer3_outputs(3448)));
    layer4_outputs(2747) <= layer3_outputs(5942);
    layer4_outputs(2748) <= layer3_outputs(3492);
    layer4_outputs(2749) <= not(layer3_outputs(5007));
    layer4_outputs(2750) <= not((layer3_outputs(7268)) and (layer3_outputs(1087)));
    layer4_outputs(2751) <= layer3_outputs(3777);
    layer4_outputs(2752) <= '1';
    layer4_outputs(2753) <= (layer3_outputs(7490)) or (layer3_outputs(5041));
    layer4_outputs(2754) <= not((layer3_outputs(5034)) and (layer3_outputs(173)));
    layer4_outputs(2755) <= not((layer3_outputs(5970)) or (layer3_outputs(5108)));
    layer4_outputs(2756) <= not(layer3_outputs(2673));
    layer4_outputs(2757) <= not(layer3_outputs(4541));
    layer4_outputs(2758) <= not(layer3_outputs(1007)) or (layer3_outputs(4047));
    layer4_outputs(2759) <= (layer3_outputs(5416)) and not (layer3_outputs(5619));
    layer4_outputs(2760) <= layer3_outputs(4570);
    layer4_outputs(2761) <= layer3_outputs(3885);
    layer4_outputs(2762) <= not(layer3_outputs(4638)) or (layer3_outputs(5400));
    layer4_outputs(2763) <= not(layer3_outputs(3460));
    layer4_outputs(2764) <= (layer3_outputs(2406)) xor (layer3_outputs(2001));
    layer4_outputs(2765) <= not((layer3_outputs(4645)) and (layer3_outputs(2190)));
    layer4_outputs(2766) <= not(layer3_outputs(2363)) or (layer3_outputs(4072));
    layer4_outputs(2767) <= not(layer3_outputs(2287));
    layer4_outputs(2768) <= not(layer3_outputs(2210));
    layer4_outputs(2769) <= not(layer3_outputs(6450));
    layer4_outputs(2770) <= not(layer3_outputs(7541));
    layer4_outputs(2771) <= not((layer3_outputs(2502)) or (layer3_outputs(6994)));
    layer4_outputs(2772) <= layer3_outputs(6447);
    layer4_outputs(2773) <= not((layer3_outputs(3377)) or (layer3_outputs(764)));
    layer4_outputs(2774) <= layer3_outputs(3690);
    layer4_outputs(2775) <= not(layer3_outputs(4856));
    layer4_outputs(2776) <= (layer3_outputs(5133)) and (layer3_outputs(3565));
    layer4_outputs(2777) <= (layer3_outputs(6963)) and not (layer3_outputs(7369));
    layer4_outputs(2778) <= (layer3_outputs(4256)) or (layer3_outputs(6904));
    layer4_outputs(2779) <= not(layer3_outputs(6693));
    layer4_outputs(2780) <= (layer3_outputs(2037)) and not (layer3_outputs(4238));
    layer4_outputs(2781) <= layer3_outputs(1692);
    layer4_outputs(2782) <= layer3_outputs(325);
    layer4_outputs(2783) <= not(layer3_outputs(7676));
    layer4_outputs(2784) <= (layer3_outputs(107)) and not (layer3_outputs(4840));
    layer4_outputs(2785) <= (layer3_outputs(6064)) or (layer3_outputs(2147));
    layer4_outputs(2786) <= not(layer3_outputs(229));
    layer4_outputs(2787) <= (layer3_outputs(5751)) and not (layer3_outputs(3564));
    layer4_outputs(2788) <= not(layer3_outputs(2656));
    layer4_outputs(2789) <= not((layer3_outputs(2986)) xor (layer3_outputs(4989)));
    layer4_outputs(2790) <= not(layer3_outputs(3418)) or (layer3_outputs(1715));
    layer4_outputs(2791) <= (layer3_outputs(3326)) and (layer3_outputs(5249));
    layer4_outputs(2792) <= not(layer3_outputs(1506));
    layer4_outputs(2793) <= (layer3_outputs(2355)) xor (layer3_outputs(2815));
    layer4_outputs(2794) <= not((layer3_outputs(4813)) and (layer3_outputs(2296)));
    layer4_outputs(2795) <= (layer3_outputs(3652)) and not (layer3_outputs(182));
    layer4_outputs(2796) <= (layer3_outputs(214)) and not (layer3_outputs(529));
    layer4_outputs(2797) <= (layer3_outputs(4618)) and not (layer3_outputs(4836));
    layer4_outputs(2798) <= not(layer3_outputs(4910));
    layer4_outputs(2799) <= not(layer3_outputs(4041));
    layer4_outputs(2800) <= not(layer3_outputs(424));
    layer4_outputs(2801) <= layer3_outputs(3288);
    layer4_outputs(2802) <= not(layer3_outputs(1676));
    layer4_outputs(2803) <= not(layer3_outputs(5847));
    layer4_outputs(2804) <= layer3_outputs(4966);
    layer4_outputs(2805) <= not((layer3_outputs(4229)) and (layer3_outputs(6143)));
    layer4_outputs(2806) <= '1';
    layer4_outputs(2807) <= layer3_outputs(633);
    layer4_outputs(2808) <= not(layer3_outputs(340));
    layer4_outputs(2809) <= (layer3_outputs(3139)) and not (layer3_outputs(2171));
    layer4_outputs(2810) <= not((layer3_outputs(7620)) or (layer3_outputs(800)));
    layer4_outputs(2811) <= (layer3_outputs(7296)) and not (layer3_outputs(5811));
    layer4_outputs(2812) <= not(layer3_outputs(5715));
    layer4_outputs(2813) <= (layer3_outputs(4079)) or (layer3_outputs(4415));
    layer4_outputs(2814) <= not(layer3_outputs(4318));
    layer4_outputs(2815) <= (layer3_outputs(372)) or (layer3_outputs(3703));
    layer4_outputs(2816) <= (layer3_outputs(1054)) and not (layer3_outputs(3389));
    layer4_outputs(2817) <= not(layer3_outputs(7638)) or (layer3_outputs(2636));
    layer4_outputs(2818) <= (layer3_outputs(5237)) or (layer3_outputs(5276));
    layer4_outputs(2819) <= not((layer3_outputs(1511)) or (layer3_outputs(6284)));
    layer4_outputs(2820) <= not(layer3_outputs(4996)) or (layer3_outputs(1117));
    layer4_outputs(2821) <= layer3_outputs(1072);
    layer4_outputs(2822) <= not(layer3_outputs(4651)) or (layer3_outputs(3695));
    layer4_outputs(2823) <= not(layer3_outputs(3730));
    layer4_outputs(2824) <= (layer3_outputs(4547)) and (layer3_outputs(6654));
    layer4_outputs(2825) <= not((layer3_outputs(2879)) and (layer3_outputs(1362)));
    layer4_outputs(2826) <= (layer3_outputs(367)) xor (layer3_outputs(4952));
    layer4_outputs(2827) <= not(layer3_outputs(58));
    layer4_outputs(2828) <= layer3_outputs(609);
    layer4_outputs(2829) <= '1';
    layer4_outputs(2830) <= (layer3_outputs(2365)) or (layer3_outputs(3919));
    layer4_outputs(2831) <= (layer3_outputs(5037)) xor (layer3_outputs(4942));
    layer4_outputs(2832) <= not((layer3_outputs(4497)) or (layer3_outputs(1359)));
    layer4_outputs(2833) <= (layer3_outputs(4934)) and not (layer3_outputs(739));
    layer4_outputs(2834) <= (layer3_outputs(3199)) and not (layer3_outputs(5682));
    layer4_outputs(2835) <= (layer3_outputs(7300)) and not (layer3_outputs(4962));
    layer4_outputs(2836) <= not(layer3_outputs(4850));
    layer4_outputs(2837) <= not((layer3_outputs(341)) and (layer3_outputs(3720)));
    layer4_outputs(2838) <= '1';
    layer4_outputs(2839) <= not((layer3_outputs(686)) and (layer3_outputs(4158)));
    layer4_outputs(2840) <= not(layer3_outputs(4954));
    layer4_outputs(2841) <= layer3_outputs(2010);
    layer4_outputs(2842) <= not((layer3_outputs(2360)) or (layer3_outputs(2006)));
    layer4_outputs(2843) <= layer3_outputs(6894);
    layer4_outputs(2844) <= layer3_outputs(6728);
    layer4_outputs(2845) <= layer3_outputs(3113);
    layer4_outputs(2846) <= layer3_outputs(3349);
    layer4_outputs(2847) <= not((layer3_outputs(904)) and (layer3_outputs(7624)));
    layer4_outputs(2848) <= (layer3_outputs(4324)) xor (layer3_outputs(2617));
    layer4_outputs(2849) <= '0';
    layer4_outputs(2850) <= not(layer3_outputs(5743)) or (layer3_outputs(1937));
    layer4_outputs(2851) <= not(layer3_outputs(2817)) or (layer3_outputs(3915));
    layer4_outputs(2852) <= not(layer3_outputs(148)) or (layer3_outputs(3689));
    layer4_outputs(2853) <= (layer3_outputs(6899)) xor (layer3_outputs(4637));
    layer4_outputs(2854) <= not(layer3_outputs(162));
    layer4_outputs(2855) <= not((layer3_outputs(2091)) or (layer3_outputs(430)));
    layer4_outputs(2856) <= (layer3_outputs(1187)) and (layer3_outputs(4251));
    layer4_outputs(2857) <= layer3_outputs(4236);
    layer4_outputs(2858) <= not(layer3_outputs(3748));
    layer4_outputs(2859) <= (layer3_outputs(7070)) and not (layer3_outputs(2536));
    layer4_outputs(2860) <= not(layer3_outputs(1358));
    layer4_outputs(2861) <= not(layer3_outputs(5828)) or (layer3_outputs(3227));
    layer4_outputs(2862) <= layer3_outputs(842);
    layer4_outputs(2863) <= layer3_outputs(3701);
    layer4_outputs(2864) <= not((layer3_outputs(3973)) xor (layer3_outputs(4509)));
    layer4_outputs(2865) <= layer3_outputs(2039);
    layer4_outputs(2866) <= not(layer3_outputs(4776)) or (layer3_outputs(7477));
    layer4_outputs(2867) <= (layer3_outputs(1163)) or (layer3_outputs(6394));
    layer4_outputs(2868) <= (layer3_outputs(904)) and (layer3_outputs(1874));
    layer4_outputs(2869) <= (layer3_outputs(1832)) and not (layer3_outputs(419));
    layer4_outputs(2870) <= not(layer3_outputs(6437));
    layer4_outputs(2871) <= '1';
    layer4_outputs(2872) <= layer3_outputs(3731);
    layer4_outputs(2873) <= layer3_outputs(1283);
    layer4_outputs(2874) <= (layer3_outputs(7527)) and not (layer3_outputs(1965));
    layer4_outputs(2875) <= not(layer3_outputs(3750));
    layer4_outputs(2876) <= not(layer3_outputs(6921)) or (layer3_outputs(2976));
    layer4_outputs(2877) <= not(layer3_outputs(1646));
    layer4_outputs(2878) <= layer3_outputs(1963);
    layer4_outputs(2879) <= '1';
    layer4_outputs(2880) <= layer3_outputs(4589);
    layer4_outputs(2881) <= not(layer3_outputs(5266));
    layer4_outputs(2882) <= not((layer3_outputs(3303)) xor (layer3_outputs(3256)));
    layer4_outputs(2883) <= not((layer3_outputs(2925)) xor (layer3_outputs(222)));
    layer4_outputs(2884) <= not(layer3_outputs(6960));
    layer4_outputs(2885) <= (layer3_outputs(2335)) and not (layer3_outputs(7563));
    layer4_outputs(2886) <= layer3_outputs(4086);
    layer4_outputs(2887) <= (layer3_outputs(3392)) and not (layer3_outputs(5007));
    layer4_outputs(2888) <= '1';
    layer4_outputs(2889) <= layer3_outputs(2063);
    layer4_outputs(2890) <= '1';
    layer4_outputs(2891) <= not((layer3_outputs(3102)) and (layer3_outputs(184)));
    layer4_outputs(2892) <= not((layer3_outputs(3693)) xor (layer3_outputs(5306)));
    layer4_outputs(2893) <= not(layer3_outputs(2683)) or (layer3_outputs(4279));
    layer4_outputs(2894) <= (layer3_outputs(7277)) xor (layer3_outputs(2308));
    layer4_outputs(2895) <= (layer3_outputs(3979)) and not (layer3_outputs(4289));
    layer4_outputs(2896) <= (layer3_outputs(6978)) and not (layer3_outputs(3474));
    layer4_outputs(2897) <= not(layer3_outputs(208)) or (layer3_outputs(2549));
    layer4_outputs(2898) <= not(layer3_outputs(6343)) or (layer3_outputs(4891));
    layer4_outputs(2899) <= not(layer3_outputs(5393)) or (layer3_outputs(5376));
    layer4_outputs(2900) <= '1';
    layer4_outputs(2901) <= layer3_outputs(3870);
    layer4_outputs(2902) <= layer3_outputs(1978);
    layer4_outputs(2903) <= layer3_outputs(4391);
    layer4_outputs(2904) <= not(layer3_outputs(4247));
    layer4_outputs(2905) <= layer3_outputs(5147);
    layer4_outputs(2906) <= not((layer3_outputs(4013)) or (layer3_outputs(5844)));
    layer4_outputs(2907) <= not(layer3_outputs(1871));
    layer4_outputs(2908) <= layer3_outputs(4197);
    layer4_outputs(2909) <= (layer3_outputs(5429)) xor (layer3_outputs(4444));
    layer4_outputs(2910) <= not(layer3_outputs(4498)) or (layer3_outputs(84));
    layer4_outputs(2911) <= not((layer3_outputs(6178)) and (layer3_outputs(2633)));
    layer4_outputs(2912) <= not(layer3_outputs(3662));
    layer4_outputs(2913) <= layer3_outputs(3212);
    layer4_outputs(2914) <= (layer3_outputs(5861)) and (layer3_outputs(2718));
    layer4_outputs(2915) <= not(layer3_outputs(247));
    layer4_outputs(2916) <= not(layer3_outputs(1057));
    layer4_outputs(2917) <= not((layer3_outputs(5166)) or (layer3_outputs(1031)));
    layer4_outputs(2918) <= layer3_outputs(5310);
    layer4_outputs(2919) <= not(layer3_outputs(5464)) or (layer3_outputs(7407));
    layer4_outputs(2920) <= not((layer3_outputs(433)) and (layer3_outputs(7581)));
    layer4_outputs(2921) <= (layer3_outputs(3545)) and not (layer3_outputs(7101));
    layer4_outputs(2922) <= (layer3_outputs(2040)) and (layer3_outputs(1136));
    layer4_outputs(2923) <= layer3_outputs(3814);
    layer4_outputs(2924) <= not(layer3_outputs(2678));
    layer4_outputs(2925) <= not((layer3_outputs(2221)) or (layer3_outputs(4409)));
    layer4_outputs(2926) <= (layer3_outputs(1127)) xor (layer3_outputs(6970));
    layer4_outputs(2927) <= '0';
    layer4_outputs(2928) <= layer3_outputs(1162);
    layer4_outputs(2929) <= layer3_outputs(7159);
    layer4_outputs(2930) <= not(layer3_outputs(2858)) or (layer3_outputs(5030));
    layer4_outputs(2931) <= layer3_outputs(7193);
    layer4_outputs(2932) <= (layer3_outputs(7049)) and (layer3_outputs(7230));
    layer4_outputs(2933) <= layer3_outputs(3010);
    layer4_outputs(2934) <= not((layer3_outputs(4362)) or (layer3_outputs(1052)));
    layer4_outputs(2935) <= not((layer3_outputs(1085)) or (layer3_outputs(5044)));
    layer4_outputs(2936) <= not(layer3_outputs(1213));
    layer4_outputs(2937) <= (layer3_outputs(4762)) xor (layer3_outputs(2591));
    layer4_outputs(2938) <= layer3_outputs(4355);
    layer4_outputs(2939) <= '0';
    layer4_outputs(2940) <= (layer3_outputs(3209)) or (layer3_outputs(217));
    layer4_outputs(2941) <= layer3_outputs(6024);
    layer4_outputs(2942) <= (layer3_outputs(1477)) and not (layer3_outputs(3289));
    layer4_outputs(2943) <= (layer3_outputs(2299)) xor (layer3_outputs(5545));
    layer4_outputs(2944) <= (layer3_outputs(2316)) or (layer3_outputs(1983));
    layer4_outputs(2945) <= '0';
    layer4_outputs(2946) <= not(layer3_outputs(530));
    layer4_outputs(2947) <= layer3_outputs(7329);
    layer4_outputs(2948) <= (layer3_outputs(5120)) and (layer3_outputs(1628));
    layer4_outputs(2949) <= layer3_outputs(6294);
    layer4_outputs(2950) <= not((layer3_outputs(2340)) and (layer3_outputs(2318)));
    layer4_outputs(2951) <= (layer3_outputs(387)) and not (layer3_outputs(2048));
    layer4_outputs(2952) <= layer3_outputs(1452);
    layer4_outputs(2953) <= not(layer3_outputs(610));
    layer4_outputs(2954) <= (layer3_outputs(2882)) xor (layer3_outputs(1902));
    layer4_outputs(2955) <= not((layer3_outputs(7609)) xor (layer3_outputs(6590)));
    layer4_outputs(2956) <= not(layer3_outputs(1683));
    layer4_outputs(2957) <= layer3_outputs(3576);
    layer4_outputs(2958) <= not(layer3_outputs(1060));
    layer4_outputs(2959) <= (layer3_outputs(1982)) xor (layer3_outputs(5521));
    layer4_outputs(2960) <= layer3_outputs(1800);
    layer4_outputs(2961) <= not(layer3_outputs(3727)) or (layer3_outputs(3301));
    layer4_outputs(2962) <= not(layer3_outputs(1525));
    layer4_outputs(2963) <= not(layer3_outputs(208));
    layer4_outputs(2964) <= '0';
    layer4_outputs(2965) <= not(layer3_outputs(2152)) or (layer3_outputs(3339));
    layer4_outputs(2966) <= layer3_outputs(2289);
    layer4_outputs(2967) <= not((layer3_outputs(2860)) or (layer3_outputs(3181)));
    layer4_outputs(2968) <= (layer3_outputs(878)) and (layer3_outputs(1610));
    layer4_outputs(2969) <= (layer3_outputs(6048)) xor (layer3_outputs(3971));
    layer4_outputs(2970) <= '0';
    layer4_outputs(2971) <= layer3_outputs(1849);
    layer4_outputs(2972) <= not(layer3_outputs(5419));
    layer4_outputs(2973) <= layer3_outputs(2109);
    layer4_outputs(2974) <= not(layer3_outputs(1304));
    layer4_outputs(2975) <= layer3_outputs(0);
    layer4_outputs(2976) <= not((layer3_outputs(6206)) and (layer3_outputs(1853)));
    layer4_outputs(2977) <= (layer3_outputs(5286)) and (layer3_outputs(7015));
    layer4_outputs(2978) <= (layer3_outputs(2597)) and not (layer3_outputs(4418));
    layer4_outputs(2979) <= (layer3_outputs(1345)) or (layer3_outputs(4057));
    layer4_outputs(2980) <= '0';
    layer4_outputs(2981) <= (layer3_outputs(1860)) and not (layer3_outputs(6315));
    layer4_outputs(2982) <= (layer3_outputs(6431)) and (layer3_outputs(1456));
    layer4_outputs(2983) <= (layer3_outputs(5346)) and not (layer3_outputs(3688));
    layer4_outputs(2984) <= layer3_outputs(3167);
    layer4_outputs(2985) <= not(layer3_outputs(4965));
    layer4_outputs(2986) <= (layer3_outputs(2965)) and not (layer3_outputs(2219));
    layer4_outputs(2987) <= (layer3_outputs(1187)) or (layer3_outputs(1236));
    layer4_outputs(2988) <= (layer3_outputs(7255)) and not (layer3_outputs(5073));
    layer4_outputs(2989) <= not((layer3_outputs(6758)) and (layer3_outputs(3647)));
    layer4_outputs(2990) <= not(layer3_outputs(1360));
    layer4_outputs(2991) <= (layer3_outputs(6789)) and not (layer3_outputs(1277));
    layer4_outputs(2992) <= layer3_outputs(818);
    layer4_outputs(2993) <= not(layer3_outputs(1487));
    layer4_outputs(2994) <= layer3_outputs(5124);
    layer4_outputs(2995) <= (layer3_outputs(3541)) and not (layer3_outputs(4352));
    layer4_outputs(2996) <= '1';
    layer4_outputs(2997) <= (layer3_outputs(2102)) xor (layer3_outputs(1496));
    layer4_outputs(2998) <= '0';
    layer4_outputs(2999) <= (layer3_outputs(5263)) or (layer3_outputs(1300));
    layer4_outputs(3000) <= not(layer3_outputs(1051));
    layer4_outputs(3001) <= (layer3_outputs(5092)) and (layer3_outputs(2537));
    layer4_outputs(3002) <= layer3_outputs(1254);
    layer4_outputs(3003) <= (layer3_outputs(4591)) and (layer3_outputs(4123));
    layer4_outputs(3004) <= '0';
    layer4_outputs(3005) <= (layer3_outputs(6153)) and (layer3_outputs(1886));
    layer4_outputs(3006) <= not(layer3_outputs(5322)) or (layer3_outputs(7238));
    layer4_outputs(3007) <= (layer3_outputs(5588)) and not (layer3_outputs(2829));
    layer4_outputs(3008) <= (layer3_outputs(2498)) or (layer3_outputs(2597));
    layer4_outputs(3009) <= not(layer3_outputs(2115));
    layer4_outputs(3010) <= '1';
    layer4_outputs(3011) <= (layer3_outputs(7257)) and not (layer3_outputs(547));
    layer4_outputs(3012) <= not((layer3_outputs(6593)) and (layer3_outputs(59)));
    layer4_outputs(3013) <= not(layer3_outputs(6871));
    layer4_outputs(3014) <= layer3_outputs(6790);
    layer4_outputs(3015) <= not(layer3_outputs(90));
    layer4_outputs(3016) <= not((layer3_outputs(6661)) or (layer3_outputs(873)));
    layer4_outputs(3017) <= layer3_outputs(751);
    layer4_outputs(3018) <= layer3_outputs(3638);
    layer4_outputs(3019) <= not(layer3_outputs(5514)) or (layer3_outputs(1501));
    layer4_outputs(3020) <= (layer3_outputs(5156)) and not (layer3_outputs(7109));
    layer4_outputs(3021) <= (layer3_outputs(3948)) and not (layer3_outputs(3570));
    layer4_outputs(3022) <= not((layer3_outputs(5288)) or (layer3_outputs(817)));
    layer4_outputs(3023) <= (layer3_outputs(2868)) or (layer3_outputs(840));
    layer4_outputs(3024) <= not((layer3_outputs(2862)) xor (layer3_outputs(103)));
    layer4_outputs(3025) <= (layer3_outputs(5465)) and not (layer3_outputs(853));
    layer4_outputs(3026) <= (layer3_outputs(3759)) and (layer3_outputs(3245));
    layer4_outputs(3027) <= layer3_outputs(6343);
    layer4_outputs(3028) <= (layer3_outputs(4196)) or (layer3_outputs(6484));
    layer4_outputs(3029) <= (layer3_outputs(801)) and not (layer3_outputs(6397));
    layer4_outputs(3030) <= not(layer3_outputs(562));
    layer4_outputs(3031) <= layer3_outputs(1571);
    layer4_outputs(3032) <= layer3_outputs(4831);
    layer4_outputs(3033) <= not(layer3_outputs(3204));
    layer4_outputs(3034) <= not(layer3_outputs(855)) or (layer3_outputs(6190));
    layer4_outputs(3035) <= not(layer3_outputs(3131));
    layer4_outputs(3036) <= layer3_outputs(4949);
    layer4_outputs(3037) <= layer3_outputs(2651);
    layer4_outputs(3038) <= layer3_outputs(2375);
    layer4_outputs(3039) <= not((layer3_outputs(2272)) or (layer3_outputs(588)));
    layer4_outputs(3040) <= layer3_outputs(2317);
    layer4_outputs(3041) <= not((layer3_outputs(5534)) or (layer3_outputs(4121)));
    layer4_outputs(3042) <= not(layer3_outputs(1195));
    layer4_outputs(3043) <= layer3_outputs(770);
    layer4_outputs(3044) <= not(layer3_outputs(2283)) or (layer3_outputs(920));
    layer4_outputs(3045) <= not(layer3_outputs(30));
    layer4_outputs(3046) <= layer3_outputs(4902);
    layer4_outputs(3047) <= '0';
    layer4_outputs(3048) <= not(layer3_outputs(3451)) or (layer3_outputs(3498));
    layer4_outputs(3049) <= not((layer3_outputs(5143)) and (layer3_outputs(23)));
    layer4_outputs(3050) <= not(layer3_outputs(3332));
    layer4_outputs(3051) <= not(layer3_outputs(3463));
    layer4_outputs(3052) <= not(layer3_outputs(2457)) or (layer3_outputs(3593));
    layer4_outputs(3053) <= not(layer3_outputs(624));
    layer4_outputs(3054) <= not((layer3_outputs(2302)) and (layer3_outputs(2850)));
    layer4_outputs(3055) <= not((layer3_outputs(686)) and (layer3_outputs(6038)));
    layer4_outputs(3056) <= not(layer3_outputs(5128));
    layer4_outputs(3057) <= not((layer3_outputs(3660)) and (layer3_outputs(2905)));
    layer4_outputs(3058) <= not(layer3_outputs(3654));
    layer4_outputs(3059) <= (layer3_outputs(81)) or (layer3_outputs(2128));
    layer4_outputs(3060) <= (layer3_outputs(4065)) or (layer3_outputs(3326));
    layer4_outputs(3061) <= not((layer3_outputs(7629)) or (layer3_outputs(2450)));
    layer4_outputs(3062) <= not(layer3_outputs(260));
    layer4_outputs(3063) <= not(layer3_outputs(3501));
    layer4_outputs(3064) <= not(layer3_outputs(3032));
    layer4_outputs(3065) <= layer3_outputs(3795);
    layer4_outputs(3066) <= (layer3_outputs(99)) xor (layer3_outputs(616));
    layer4_outputs(3067) <= not((layer3_outputs(5796)) and (layer3_outputs(4408)));
    layer4_outputs(3068) <= layer3_outputs(5353);
    layer4_outputs(3069) <= not(layer3_outputs(6349));
    layer4_outputs(3070) <= (layer3_outputs(2832)) and not (layer3_outputs(5655));
    layer4_outputs(3071) <= not(layer3_outputs(4016));
    layer4_outputs(3072) <= not((layer3_outputs(6903)) and (layer3_outputs(7058)));
    layer4_outputs(3073) <= layer3_outputs(552);
    layer4_outputs(3074) <= layer3_outputs(4518);
    layer4_outputs(3075) <= not(layer3_outputs(1190));
    layer4_outputs(3076) <= (layer3_outputs(3198)) and (layer3_outputs(3141));
    layer4_outputs(3077) <= layer3_outputs(1404);
    layer4_outputs(3078) <= layer3_outputs(2119);
    layer4_outputs(3079) <= '0';
    layer4_outputs(3080) <= not(layer3_outputs(5520));
    layer4_outputs(3081) <= not((layer3_outputs(7034)) and (layer3_outputs(3157)));
    layer4_outputs(3082) <= not(layer3_outputs(7066));
    layer4_outputs(3083) <= layer3_outputs(3846);
    layer4_outputs(3084) <= (layer3_outputs(2812)) or (layer3_outputs(4818));
    layer4_outputs(3085) <= (layer3_outputs(6407)) and not (layer3_outputs(3937));
    layer4_outputs(3086) <= layer3_outputs(1223);
    layer4_outputs(3087) <= (layer3_outputs(6153)) and not (layer3_outputs(1573));
    layer4_outputs(3088) <= not(layer3_outputs(1544));
    layer4_outputs(3089) <= (layer3_outputs(7625)) or (layer3_outputs(5527));
    layer4_outputs(3090) <= not((layer3_outputs(3358)) or (layer3_outputs(4152)));
    layer4_outputs(3091) <= (layer3_outputs(6138)) and not (layer3_outputs(3822));
    layer4_outputs(3092) <= '1';
    layer4_outputs(3093) <= '0';
    layer4_outputs(3094) <= layer3_outputs(1363);
    layer4_outputs(3095) <= not((layer3_outputs(6723)) xor (layer3_outputs(199)));
    layer4_outputs(3096) <= (layer3_outputs(694)) or (layer3_outputs(2567));
    layer4_outputs(3097) <= '0';
    layer4_outputs(3098) <= not(layer3_outputs(4660)) or (layer3_outputs(2345));
    layer4_outputs(3099) <= not(layer3_outputs(457));
    layer4_outputs(3100) <= (layer3_outputs(4969)) and not (layer3_outputs(7453));
    layer4_outputs(3101) <= not(layer3_outputs(7545));
    layer4_outputs(3102) <= not(layer3_outputs(792)) or (layer3_outputs(7290));
    layer4_outputs(3103) <= not(layer3_outputs(7338));
    layer4_outputs(3104) <= '0';
    layer4_outputs(3105) <= layer3_outputs(5207);
    layer4_outputs(3106) <= '0';
    layer4_outputs(3107) <= '1';
    layer4_outputs(3108) <= not((layer3_outputs(2344)) xor (layer3_outputs(6193)));
    layer4_outputs(3109) <= layer3_outputs(1338);
    layer4_outputs(3110) <= layer3_outputs(3807);
    layer4_outputs(3111) <= '0';
    layer4_outputs(3112) <= not((layer3_outputs(418)) or (layer3_outputs(3616)));
    layer4_outputs(3113) <= not(layer3_outputs(877));
    layer4_outputs(3114) <= (layer3_outputs(4272)) and not (layer3_outputs(7));
    layer4_outputs(3115) <= not(layer3_outputs(2126));
    layer4_outputs(3116) <= '0';
    layer4_outputs(3117) <= layer3_outputs(3415);
    layer4_outputs(3118) <= not(layer3_outputs(2521)) or (layer3_outputs(1916));
    layer4_outputs(3119) <= not(layer3_outputs(6135));
    layer4_outputs(3120) <= layer3_outputs(260);
    layer4_outputs(3121) <= not(layer3_outputs(3696));
    layer4_outputs(3122) <= (layer3_outputs(1121)) and (layer3_outputs(4390));
    layer4_outputs(3123) <= (layer3_outputs(1)) or (layer3_outputs(5411));
    layer4_outputs(3124) <= not((layer3_outputs(2696)) or (layer3_outputs(5437)));
    layer4_outputs(3125) <= (layer3_outputs(6016)) or (layer3_outputs(3344));
    layer4_outputs(3126) <= not(layer3_outputs(557));
    layer4_outputs(3127) <= layer3_outputs(4360);
    layer4_outputs(3128) <= (layer3_outputs(5450)) and not (layer3_outputs(281));
    layer4_outputs(3129) <= not((layer3_outputs(1078)) xor (layer3_outputs(687)));
    layer4_outputs(3130) <= '0';
    layer4_outputs(3131) <= layer3_outputs(4112);
    layer4_outputs(3132) <= layer3_outputs(6781);
    layer4_outputs(3133) <= (layer3_outputs(6860)) and not (layer3_outputs(4878));
    layer4_outputs(3134) <= (layer3_outputs(5036)) or (layer3_outputs(4600));
    layer4_outputs(3135) <= not(layer3_outputs(5037));
    layer4_outputs(3136) <= (layer3_outputs(5234)) and (layer3_outputs(6131));
    layer4_outputs(3137) <= not(layer3_outputs(351)) or (layer3_outputs(2947));
    layer4_outputs(3138) <= (layer3_outputs(3428)) or (layer3_outputs(1760));
    layer4_outputs(3139) <= not((layer3_outputs(5679)) or (layer3_outputs(1984)));
    layer4_outputs(3140) <= not(layer3_outputs(4464));
    layer4_outputs(3141) <= layer3_outputs(1552);
    layer4_outputs(3142) <= (layer3_outputs(3191)) and not (layer3_outputs(4432));
    layer4_outputs(3143) <= not(layer3_outputs(2206));
    layer4_outputs(3144) <= layer3_outputs(274);
    layer4_outputs(3145) <= layer3_outputs(4588);
    layer4_outputs(3146) <= (layer3_outputs(3989)) and not (layer3_outputs(7458));
    layer4_outputs(3147) <= not((layer3_outputs(296)) xor (layer3_outputs(4709)));
    layer4_outputs(3148) <= layer3_outputs(7175);
    layer4_outputs(3149) <= (layer3_outputs(5851)) and not (layer3_outputs(91));
    layer4_outputs(3150) <= layer3_outputs(270);
    layer4_outputs(3151) <= not(layer3_outputs(1344));
    layer4_outputs(3152) <= layer3_outputs(3408);
    layer4_outputs(3153) <= not((layer3_outputs(3122)) or (layer3_outputs(3029)));
    layer4_outputs(3154) <= (layer3_outputs(6298)) xor (layer3_outputs(4863));
    layer4_outputs(3155) <= not(layer3_outputs(5804));
    layer4_outputs(3156) <= not(layer3_outputs(2447)) or (layer3_outputs(1522));
    layer4_outputs(3157) <= layer3_outputs(329);
    layer4_outputs(3158) <= (layer3_outputs(6479)) and not (layer3_outputs(6497));
    layer4_outputs(3159) <= layer3_outputs(2655);
    layer4_outputs(3160) <= (layer3_outputs(1752)) or (layer3_outputs(2023));
    layer4_outputs(3161) <= (layer3_outputs(2458)) xor (layer3_outputs(4990));
    layer4_outputs(3162) <= not(layer3_outputs(736)) or (layer3_outputs(671));
    layer4_outputs(3163) <= (layer3_outputs(193)) and not (layer3_outputs(7080));
    layer4_outputs(3164) <= not((layer3_outputs(6091)) and (layer3_outputs(606)));
    layer4_outputs(3165) <= not(layer3_outputs(7080));
    layer4_outputs(3166) <= not(layer3_outputs(2052)) or (layer3_outputs(3966));
    layer4_outputs(3167) <= not(layer3_outputs(7544)) or (layer3_outputs(6339));
    layer4_outputs(3168) <= layer3_outputs(784);
    layer4_outputs(3169) <= (layer3_outputs(145)) or (layer3_outputs(3370));
    layer4_outputs(3170) <= layer3_outputs(125);
    layer4_outputs(3171) <= not(layer3_outputs(4143));
    layer4_outputs(3172) <= not(layer3_outputs(5113));
    layer4_outputs(3173) <= not((layer3_outputs(6485)) or (layer3_outputs(814)));
    layer4_outputs(3174) <= (layer3_outputs(3441)) and not (layer3_outputs(6751));
    layer4_outputs(3175) <= layer3_outputs(6277);
    layer4_outputs(3176) <= not((layer3_outputs(2369)) and (layer3_outputs(3249)));
    layer4_outputs(3177) <= layer3_outputs(6089);
    layer4_outputs(3178) <= not(layer3_outputs(2911)) or (layer3_outputs(4566));
    layer4_outputs(3179) <= layer3_outputs(5232);
    layer4_outputs(3180) <= not(layer3_outputs(6919)) or (layer3_outputs(5436));
    layer4_outputs(3181) <= not(layer3_outputs(25));
    layer4_outputs(3182) <= not((layer3_outputs(3422)) xor (layer3_outputs(5330)));
    layer4_outputs(3183) <= (layer3_outputs(5664)) or (layer3_outputs(328));
    layer4_outputs(3184) <= (layer3_outputs(1206)) and not (layer3_outputs(4414));
    layer4_outputs(3185) <= not(layer3_outputs(747));
    layer4_outputs(3186) <= not((layer3_outputs(775)) xor (layer3_outputs(6103)));
    layer4_outputs(3187) <= (layer3_outputs(658)) and not (layer3_outputs(5492));
    layer4_outputs(3188) <= not(layer3_outputs(6197));
    layer4_outputs(3189) <= layer3_outputs(3745);
    layer4_outputs(3190) <= (layer3_outputs(2926)) and not (layer3_outputs(2863));
    layer4_outputs(3191) <= (layer3_outputs(975)) or (layer3_outputs(1049));
    layer4_outputs(3192) <= not((layer3_outputs(4047)) or (layer3_outputs(3299)));
    layer4_outputs(3193) <= not((layer3_outputs(2247)) or (layer3_outputs(704)));
    layer4_outputs(3194) <= not(layer3_outputs(6313));
    layer4_outputs(3195) <= not(layer3_outputs(5478));
    layer4_outputs(3196) <= not(layer3_outputs(7489));
    layer4_outputs(3197) <= not(layer3_outputs(933)) or (layer3_outputs(4677));
    layer4_outputs(3198) <= (layer3_outputs(950)) and not (layer3_outputs(2699));
    layer4_outputs(3199) <= (layer3_outputs(3617)) or (layer3_outputs(5084));
    layer4_outputs(3200) <= '1';
    layer4_outputs(3201) <= not(layer3_outputs(6265));
    layer4_outputs(3202) <= layer3_outputs(2579);
    layer4_outputs(3203) <= (layer3_outputs(4680)) and (layer3_outputs(5676));
    layer4_outputs(3204) <= not((layer3_outputs(2384)) and (layer3_outputs(465)));
    layer4_outputs(3205) <= (layer3_outputs(2131)) and not (layer3_outputs(2860));
    layer4_outputs(3206) <= (layer3_outputs(2107)) and not (layer3_outputs(637));
    layer4_outputs(3207) <= not(layer3_outputs(5354));
    layer4_outputs(3208) <= (layer3_outputs(38)) and not (layer3_outputs(2935));
    layer4_outputs(3209) <= not(layer3_outputs(5511));
    layer4_outputs(3210) <= layer3_outputs(1780);
    layer4_outputs(3211) <= not(layer3_outputs(3385));
    layer4_outputs(3212) <= not(layer3_outputs(6729)) or (layer3_outputs(4194));
    layer4_outputs(3213) <= (layer3_outputs(2100)) or (layer3_outputs(5412));
    layer4_outputs(3214) <= (layer3_outputs(5190)) or (layer3_outputs(1704));
    layer4_outputs(3215) <= layer3_outputs(3734);
    layer4_outputs(3216) <= layer3_outputs(5061);
    layer4_outputs(3217) <= (layer3_outputs(7362)) and not (layer3_outputs(2916));
    layer4_outputs(3218) <= not(layer3_outputs(16));
    layer4_outputs(3219) <= not(layer3_outputs(2639));
    layer4_outputs(3220) <= not(layer3_outputs(2853));
    layer4_outputs(3221) <= not(layer3_outputs(2399));
    layer4_outputs(3222) <= not(layer3_outputs(7633)) or (layer3_outputs(2435));
    layer4_outputs(3223) <= not((layer3_outputs(5858)) and (layer3_outputs(1077)));
    layer4_outputs(3224) <= not(layer3_outputs(6355));
    layer4_outputs(3225) <= not((layer3_outputs(753)) xor (layer3_outputs(7453)));
    layer4_outputs(3226) <= not((layer3_outputs(4689)) or (layer3_outputs(5957)));
    layer4_outputs(3227) <= layer3_outputs(4964);
    layer4_outputs(3228) <= layer3_outputs(2893);
    layer4_outputs(3229) <= (layer3_outputs(1635)) and not (layer3_outputs(3619));
    layer4_outputs(3230) <= (layer3_outputs(410)) xor (layer3_outputs(1845));
    layer4_outputs(3231) <= not(layer3_outputs(3244)) or (layer3_outputs(3679));
    layer4_outputs(3232) <= (layer3_outputs(4312)) and not (layer3_outputs(184));
    layer4_outputs(3233) <= not(layer3_outputs(4486)) or (layer3_outputs(4410));
    layer4_outputs(3234) <= layer3_outputs(2327);
    layer4_outputs(3235) <= not(layer3_outputs(3866));
    layer4_outputs(3236) <= layer3_outputs(4271);
    layer4_outputs(3237) <= not(layer3_outputs(6736));
    layer4_outputs(3238) <= layer3_outputs(6910);
    layer4_outputs(3239) <= layer3_outputs(777);
    layer4_outputs(3240) <= layer3_outputs(1727);
    layer4_outputs(3241) <= not(layer3_outputs(5693)) or (layer3_outputs(1570));
    layer4_outputs(3242) <= layer3_outputs(4537);
    layer4_outputs(3243) <= layer3_outputs(1291);
    layer4_outputs(3244) <= not(layer3_outputs(542));
    layer4_outputs(3245) <= (layer3_outputs(761)) and (layer3_outputs(7439));
    layer4_outputs(3246) <= not((layer3_outputs(5084)) xor (layer3_outputs(5316)));
    layer4_outputs(3247) <= layer3_outputs(908);
    layer4_outputs(3248) <= (layer3_outputs(6121)) xor (layer3_outputs(2754));
    layer4_outputs(3249) <= not(layer3_outputs(28));
    layer4_outputs(3250) <= layer3_outputs(6963);
    layer4_outputs(3251) <= layer3_outputs(5163);
    layer4_outputs(3252) <= layer3_outputs(3353);
    layer4_outputs(3253) <= not(layer3_outputs(4369));
    layer4_outputs(3254) <= not(layer3_outputs(86)) or (layer3_outputs(6491));
    layer4_outputs(3255) <= not(layer3_outputs(1697));
    layer4_outputs(3256) <= (layer3_outputs(4815)) and not (layer3_outputs(6825));
    layer4_outputs(3257) <= not((layer3_outputs(6434)) xor (layer3_outputs(5021)));
    layer4_outputs(3258) <= '1';
    layer4_outputs(3259) <= (layer3_outputs(2751)) and (layer3_outputs(7182));
    layer4_outputs(3260) <= '0';
    layer4_outputs(3261) <= not(layer3_outputs(5416));
    layer4_outputs(3262) <= not(layer3_outputs(6880)) or (layer3_outputs(6248));
    layer4_outputs(3263) <= not((layer3_outputs(6198)) xor (layer3_outputs(3562)));
    layer4_outputs(3264) <= not(layer3_outputs(2262)) or (layer3_outputs(3918));
    layer4_outputs(3265) <= not(layer3_outputs(4639)) or (layer3_outputs(6879));
    layer4_outputs(3266) <= '0';
    layer4_outputs(3267) <= not((layer3_outputs(116)) xor (layer3_outputs(2634)));
    layer4_outputs(3268) <= (layer3_outputs(3154)) and not (layer3_outputs(6340));
    layer4_outputs(3269) <= layer3_outputs(4080);
    layer4_outputs(3270) <= (layer3_outputs(257)) and (layer3_outputs(6306));
    layer4_outputs(3271) <= layer3_outputs(5388);
    layer4_outputs(3272) <= (layer3_outputs(786)) and not (layer3_outputs(6526));
    layer4_outputs(3273) <= '0';
    layer4_outputs(3274) <= not(layer3_outputs(7316)) or (layer3_outputs(5355));
    layer4_outputs(3275) <= (layer3_outputs(3538)) and not (layer3_outputs(4386));
    layer4_outputs(3276) <= not(layer3_outputs(3607));
    layer4_outputs(3277) <= not(layer3_outputs(6707)) or (layer3_outputs(1579));
    layer4_outputs(3278) <= layer3_outputs(2430);
    layer4_outputs(3279) <= not(layer3_outputs(1878)) or (layer3_outputs(3653));
    layer4_outputs(3280) <= not((layer3_outputs(4955)) and (layer3_outputs(5397)));
    layer4_outputs(3281) <= not(layer3_outputs(6310)) or (layer3_outputs(4986));
    layer4_outputs(3282) <= not(layer3_outputs(7671)) or (layer3_outputs(7434));
    layer4_outputs(3283) <= '0';
    layer4_outputs(3284) <= (layer3_outputs(5701)) and not (layer3_outputs(1370));
    layer4_outputs(3285) <= not(layer3_outputs(1768));
    layer4_outputs(3286) <= layer3_outputs(3011);
    layer4_outputs(3287) <= not(layer3_outputs(7183));
    layer4_outputs(3288) <= (layer3_outputs(2979)) and (layer3_outputs(7324));
    layer4_outputs(3289) <= not(layer3_outputs(1913));
    layer4_outputs(3290) <= layer3_outputs(7013);
    layer4_outputs(3291) <= layer3_outputs(2491);
    layer4_outputs(3292) <= layer3_outputs(236);
    layer4_outputs(3293) <= layer3_outputs(6999);
    layer4_outputs(3294) <= layer3_outputs(6669);
    layer4_outputs(3295) <= not(layer3_outputs(2269));
    layer4_outputs(3296) <= (layer3_outputs(2543)) and not (layer3_outputs(1902));
    layer4_outputs(3297) <= layer3_outputs(5810);
    layer4_outputs(3298) <= not(layer3_outputs(3012)) or (layer3_outputs(2788));
    layer4_outputs(3299) <= (layer3_outputs(5219)) xor (layer3_outputs(3317));
    layer4_outputs(3300) <= (layer3_outputs(2422)) and not (layer3_outputs(317));
    layer4_outputs(3301) <= not((layer3_outputs(942)) and (layer3_outputs(6794)));
    layer4_outputs(3302) <= not(layer3_outputs(4899));
    layer4_outputs(3303) <= not((layer3_outputs(1212)) xor (layer3_outputs(6477)));
    layer4_outputs(3304) <= layer3_outputs(938);
    layer4_outputs(3305) <= not((layer3_outputs(16)) or (layer3_outputs(1891)));
    layer4_outputs(3306) <= layer3_outputs(6000);
    layer4_outputs(3307) <= not(layer3_outputs(7418));
    layer4_outputs(3308) <= not(layer3_outputs(1180));
    layer4_outputs(3309) <= not(layer3_outputs(856)) or (layer3_outputs(6980));
    layer4_outputs(3310) <= not((layer3_outputs(6104)) or (layer3_outputs(724)));
    layer4_outputs(3311) <= layer3_outputs(4842);
    layer4_outputs(3312) <= '0';
    layer4_outputs(3313) <= layer3_outputs(3594);
    layer4_outputs(3314) <= not(layer3_outputs(637)) or (layer3_outputs(6667));
    layer4_outputs(3315) <= layer3_outputs(4690);
    layer4_outputs(3316) <= not((layer3_outputs(5822)) or (layer3_outputs(7397)));
    layer4_outputs(3317) <= layer3_outputs(3955);
    layer4_outputs(3318) <= not(layer3_outputs(6973)) or (layer3_outputs(6081));
    layer4_outputs(3319) <= not(layer3_outputs(5291));
    layer4_outputs(3320) <= (layer3_outputs(3410)) and not (layer3_outputs(918));
    layer4_outputs(3321) <= layer3_outputs(5903);
    layer4_outputs(3322) <= (layer3_outputs(3413)) and not (layer3_outputs(4436));
    layer4_outputs(3323) <= not(layer3_outputs(7185));
    layer4_outputs(3324) <= not(layer3_outputs(3546));
    layer4_outputs(3325) <= not((layer3_outputs(6664)) or (layer3_outputs(2247)));
    layer4_outputs(3326) <= '0';
    layer4_outputs(3327) <= layer3_outputs(4854);
    layer4_outputs(3328) <= not((layer3_outputs(2367)) and (layer3_outputs(3424)));
    layer4_outputs(3329) <= not((layer3_outputs(1797)) and (layer3_outputs(7134)));
    layer4_outputs(3330) <= not(layer3_outputs(5457)) or (layer3_outputs(6282));
    layer4_outputs(3331) <= (layer3_outputs(1713)) and not (layer3_outputs(3527));
    layer4_outputs(3332) <= '0';
    layer4_outputs(3333) <= layer3_outputs(227);
    layer4_outputs(3334) <= not(layer3_outputs(5593));
    layer4_outputs(3335) <= not(layer3_outputs(5052));
    layer4_outputs(3336) <= not((layer3_outputs(5616)) or (layer3_outputs(6050)));
    layer4_outputs(3337) <= not((layer3_outputs(6642)) or (layer3_outputs(1255)));
    layer4_outputs(3338) <= layer3_outputs(4798);
    layer4_outputs(3339) <= (layer3_outputs(7398)) or (layer3_outputs(3587));
    layer4_outputs(3340) <= layer3_outputs(6307);
    layer4_outputs(3341) <= '0';
    layer4_outputs(3342) <= layer3_outputs(7420);
    layer4_outputs(3343) <= '0';
    layer4_outputs(3344) <= (layer3_outputs(2642)) or (layer3_outputs(2942));
    layer4_outputs(3345) <= not((layer3_outputs(4602)) xor (layer3_outputs(5863)));
    layer4_outputs(3346) <= (layer3_outputs(2759)) and not (layer3_outputs(1046));
    layer4_outputs(3347) <= not((layer3_outputs(5061)) xor (layer3_outputs(4215)));
    layer4_outputs(3348) <= layer3_outputs(6649);
    layer4_outputs(3349) <= (layer3_outputs(6281)) and not (layer3_outputs(5022));
    layer4_outputs(3350) <= not(layer3_outputs(5932)) or (layer3_outputs(3054));
    layer4_outputs(3351) <= layer3_outputs(4951);
    layer4_outputs(3352) <= layer3_outputs(4328);
    layer4_outputs(3353) <= (layer3_outputs(7602)) and not (layer3_outputs(1502));
    layer4_outputs(3354) <= '0';
    layer4_outputs(3355) <= not(layer3_outputs(1028)) or (layer3_outputs(1731));
    layer4_outputs(3356) <= not((layer3_outputs(5489)) and (layer3_outputs(2845)));
    layer4_outputs(3357) <= not((layer3_outputs(5285)) and (layer3_outputs(2027)));
    layer4_outputs(3358) <= not((layer3_outputs(6632)) or (layer3_outputs(5200)));
    layer4_outputs(3359) <= (layer3_outputs(390)) or (layer3_outputs(6796));
    layer4_outputs(3360) <= (layer3_outputs(2535)) and not (layer3_outputs(7549));
    layer4_outputs(3361) <= (layer3_outputs(6754)) and not (layer3_outputs(7256));
    layer4_outputs(3362) <= layer3_outputs(2727);
    layer4_outputs(3363) <= (layer3_outputs(7093)) and not (layer3_outputs(2402));
    layer4_outputs(3364) <= (layer3_outputs(6370)) and not (layer3_outputs(2003));
    layer4_outputs(3365) <= (layer3_outputs(3928)) or (layer3_outputs(5008));
    layer4_outputs(3366) <= not((layer3_outputs(1533)) and (layer3_outputs(137)));
    layer4_outputs(3367) <= '0';
    layer4_outputs(3368) <= not((layer3_outputs(6127)) xor (layer3_outputs(5187)));
    layer4_outputs(3369) <= (layer3_outputs(6239)) and not (layer3_outputs(6213));
    layer4_outputs(3370) <= not(layer3_outputs(3209));
    layer4_outputs(3371) <= layer3_outputs(3589);
    layer4_outputs(3372) <= '0';
    layer4_outputs(3373) <= not(layer3_outputs(7532)) or (layer3_outputs(2660));
    layer4_outputs(3374) <= layer3_outputs(6357);
    layer4_outputs(3375) <= layer3_outputs(5510);
    layer4_outputs(3376) <= (layer3_outputs(684)) and not (layer3_outputs(4987));
    layer4_outputs(3377) <= layer3_outputs(4809);
    layer4_outputs(3378) <= not(layer3_outputs(6902)) or (layer3_outputs(2937));
    layer4_outputs(3379) <= layer3_outputs(6690);
    layer4_outputs(3380) <= layer3_outputs(4995);
    layer4_outputs(3381) <= not((layer3_outputs(2241)) and (layer3_outputs(4345)));
    layer4_outputs(3382) <= not(layer3_outputs(5135)) or (layer3_outputs(5600));
    layer4_outputs(3383) <= (layer3_outputs(7151)) and not (layer3_outputs(5414));
    layer4_outputs(3384) <= layer3_outputs(1725);
    layer4_outputs(3385) <= layer3_outputs(6366);
    layer4_outputs(3386) <= '1';
    layer4_outputs(3387) <= layer3_outputs(6187);
    layer4_outputs(3388) <= layer3_outputs(2923);
    layer4_outputs(3389) <= not(layer3_outputs(4817));
    layer4_outputs(3390) <= layer3_outputs(2431);
    layer4_outputs(3391) <= not(layer3_outputs(1092));
    layer4_outputs(3392) <= layer3_outputs(4922);
    layer4_outputs(3393) <= not(layer3_outputs(31));
    layer4_outputs(3394) <= (layer3_outputs(3352)) and (layer3_outputs(2485));
    layer4_outputs(3395) <= not((layer3_outputs(6770)) xor (layer3_outputs(4999)));
    layer4_outputs(3396) <= layer3_outputs(3525);
    layer4_outputs(3397) <= not(layer3_outputs(3509));
    layer4_outputs(3398) <= '0';
    layer4_outputs(3399) <= layer3_outputs(4614);
    layer4_outputs(3400) <= (layer3_outputs(5241)) and not (layer3_outputs(5352));
    layer4_outputs(3401) <= (layer3_outputs(3922)) and not (layer3_outputs(1631));
    layer4_outputs(3402) <= (layer3_outputs(198)) and not (layer3_outputs(4074));
    layer4_outputs(3403) <= layer3_outputs(4400);
    layer4_outputs(3404) <= not(layer3_outputs(4476));
    layer4_outputs(3405) <= layer3_outputs(6681);
    layer4_outputs(3406) <= not((layer3_outputs(5360)) xor (layer3_outputs(1369)));
    layer4_outputs(3407) <= not((layer3_outputs(6596)) and (layer3_outputs(4559)));
    layer4_outputs(3408) <= not((layer3_outputs(3328)) xor (layer3_outputs(2222)));
    layer4_outputs(3409) <= not(layer3_outputs(6800));
    layer4_outputs(3410) <= layer3_outputs(5086);
    layer4_outputs(3411) <= '0';
    layer4_outputs(3412) <= not(layer3_outputs(4877)) or (layer3_outputs(2952));
    layer4_outputs(3413) <= not((layer3_outputs(3583)) or (layer3_outputs(1489)));
    layer4_outputs(3414) <= not((layer3_outputs(4313)) and (layer3_outputs(3951)));
    layer4_outputs(3415) <= (layer3_outputs(7598)) and (layer3_outputs(5644));
    layer4_outputs(3416) <= not(layer3_outputs(438));
    layer4_outputs(3417) <= (layer3_outputs(5363)) and not (layer3_outputs(751));
    layer4_outputs(3418) <= not(layer3_outputs(3558));
    layer4_outputs(3419) <= not(layer3_outputs(1311));
    layer4_outputs(3420) <= (layer3_outputs(3486)) and not (layer3_outputs(7062));
    layer4_outputs(3421) <= '0';
    layer4_outputs(3422) <= not(layer3_outputs(4991));
    layer4_outputs(3423) <= not((layer3_outputs(1814)) or (layer3_outputs(7369)));
    layer4_outputs(3424) <= (layer3_outputs(6542)) and not (layer3_outputs(3223));
    layer4_outputs(3425) <= not(layer3_outputs(4022));
    layer4_outputs(3426) <= (layer3_outputs(2578)) and (layer3_outputs(3595));
    layer4_outputs(3427) <= not((layer3_outputs(847)) xor (layer3_outputs(3650)));
    layer4_outputs(3428) <= not(layer3_outputs(4097));
    layer4_outputs(3429) <= layer3_outputs(5790);
    layer4_outputs(3430) <= not((layer3_outputs(6906)) and (layer3_outputs(6966)));
    layer4_outputs(3431) <= (layer3_outputs(7511)) and not (layer3_outputs(5415));
    layer4_outputs(3432) <= not(layer3_outputs(5572));
    layer4_outputs(3433) <= not(layer3_outputs(5739));
    layer4_outputs(3434) <= (layer3_outputs(4574)) and (layer3_outputs(1120));
    layer4_outputs(3435) <= not(layer3_outputs(804));
    layer4_outputs(3436) <= (layer3_outputs(633)) and not (layer3_outputs(6223));
    layer4_outputs(3437) <= not(layer3_outputs(7574));
    layer4_outputs(3438) <= not(layer3_outputs(1498));
    layer4_outputs(3439) <= not((layer3_outputs(600)) and (layer3_outputs(2062)));
    layer4_outputs(3440) <= (layer3_outputs(1015)) or (layer3_outputs(1416));
    layer4_outputs(3441) <= '0';
    layer4_outputs(3442) <= not((layer3_outputs(1703)) or (layer3_outputs(3709)));
    layer4_outputs(3443) <= not(layer3_outputs(1997));
    layer4_outputs(3444) <= '0';
    layer4_outputs(3445) <= not((layer3_outputs(5666)) xor (layer3_outputs(2492)));
    layer4_outputs(3446) <= not(layer3_outputs(7239));
    layer4_outputs(3447) <= layer3_outputs(11);
    layer4_outputs(3448) <= (layer3_outputs(2451)) and not (layer3_outputs(1868));
    layer4_outputs(3449) <= not(layer3_outputs(2064));
    layer4_outputs(3450) <= layer3_outputs(5714);
    layer4_outputs(3451) <= not((layer3_outputs(1743)) xor (layer3_outputs(2853)));
    layer4_outputs(3452) <= layer3_outputs(519);
    layer4_outputs(3453) <= layer3_outputs(2785);
    layer4_outputs(3454) <= not(layer3_outputs(4562)) or (layer3_outputs(4126));
    layer4_outputs(3455) <= (layer3_outputs(3385)) or (layer3_outputs(7120));
    layer4_outputs(3456) <= layer3_outputs(1036);
    layer4_outputs(3457) <= not(layer3_outputs(3147));
    layer4_outputs(3458) <= not(layer3_outputs(1312));
    layer4_outputs(3459) <= not(layer3_outputs(5642));
    layer4_outputs(3460) <= layer3_outputs(5192);
    layer4_outputs(3461) <= layer3_outputs(6404);
    layer4_outputs(3462) <= layer3_outputs(3212);
    layer4_outputs(3463) <= not(layer3_outputs(6950));
    layer4_outputs(3464) <= (layer3_outputs(5134)) and not (layer3_outputs(7483));
    layer4_outputs(3465) <= not(layer3_outputs(3156));
    layer4_outputs(3466) <= layer3_outputs(2921);
    layer4_outputs(3467) <= not((layer3_outputs(1961)) or (layer3_outputs(5941)));
    layer4_outputs(3468) <= not(layer3_outputs(6156));
    layer4_outputs(3469) <= (layer3_outputs(416)) xor (layer3_outputs(3006));
    layer4_outputs(3470) <= not((layer3_outputs(1718)) or (layer3_outputs(1481)));
    layer4_outputs(3471) <= (layer3_outputs(6704)) and (layer3_outputs(7402));
    layer4_outputs(3472) <= layer3_outputs(5999);
    layer4_outputs(3473) <= (layer3_outputs(1011)) and not (layer3_outputs(358));
    layer4_outputs(3474) <= (layer3_outputs(2446)) and (layer3_outputs(238));
    layer4_outputs(3475) <= not(layer3_outputs(495));
    layer4_outputs(3476) <= layer3_outputs(4632);
    layer4_outputs(3477) <= not(layer3_outputs(6085));
    layer4_outputs(3478) <= not(layer3_outputs(614));
    layer4_outputs(3479) <= layer3_outputs(6693);
    layer4_outputs(3480) <= layer3_outputs(5117);
    layer4_outputs(3481) <= layer3_outputs(3909);
    layer4_outputs(3482) <= layer3_outputs(5160);
    layer4_outputs(3483) <= not(layer3_outputs(225)) or (layer3_outputs(5158));
    layer4_outputs(3484) <= not(layer3_outputs(3544)) or (layer3_outputs(5640));
    layer4_outputs(3485) <= not(layer3_outputs(7389));
    layer4_outputs(3486) <= not((layer3_outputs(5361)) or (layer3_outputs(1332)));
    layer4_outputs(3487) <= not(layer3_outputs(5095));
    layer4_outputs(3488) <= not((layer3_outputs(2472)) and (layer3_outputs(4506)));
    layer4_outputs(3489) <= not(layer3_outputs(6260));
    layer4_outputs(3490) <= not(layer3_outputs(4293));
    layer4_outputs(3491) <= not(layer3_outputs(6852));
    layer4_outputs(3492) <= '0';
    layer4_outputs(3493) <= layer3_outputs(2845);
    layer4_outputs(3494) <= not((layer3_outputs(2824)) xor (layer3_outputs(1643)));
    layer4_outputs(3495) <= layer3_outputs(6647);
    layer4_outputs(3496) <= not(layer3_outputs(4571));
    layer4_outputs(3497) <= not(layer3_outputs(5228)) or (layer3_outputs(6167));
    layer4_outputs(3498) <= '0';
    layer4_outputs(3499) <= layer3_outputs(890);
    layer4_outputs(3500) <= (layer3_outputs(7020)) and (layer3_outputs(2833));
    layer4_outputs(3501) <= layer3_outputs(5841);
    layer4_outputs(3502) <= not((layer3_outputs(4210)) or (layer3_outputs(5464)));
    layer4_outputs(3503) <= '1';
    layer4_outputs(3504) <= layer3_outputs(1500);
    layer4_outputs(3505) <= (layer3_outputs(5239)) xor (layer3_outputs(5678));
    layer4_outputs(3506) <= (layer3_outputs(7173)) and not (layer3_outputs(6076));
    layer4_outputs(3507) <= (layer3_outputs(3751)) and not (layer3_outputs(158));
    layer4_outputs(3508) <= not(layer3_outputs(7364)) or (layer3_outputs(5874));
    layer4_outputs(3509) <= layer3_outputs(1996);
    layer4_outputs(3510) <= not(layer3_outputs(908)) or (layer3_outputs(5401));
    layer4_outputs(3511) <= layer3_outputs(4149);
    layer4_outputs(3512) <= not(layer3_outputs(303)) or (layer3_outputs(7169));
    layer4_outputs(3513) <= not(layer3_outputs(5091));
    layer4_outputs(3514) <= not(layer3_outputs(3416));
    layer4_outputs(3515) <= '0';
    layer4_outputs(3516) <= layer3_outputs(2343);
    layer4_outputs(3517) <= layer3_outputs(3797);
    layer4_outputs(3518) <= '1';
    layer4_outputs(3519) <= layer3_outputs(6589);
    layer4_outputs(3520) <= (layer3_outputs(5663)) and not (layer3_outputs(1320));
    layer4_outputs(3521) <= '0';
    layer4_outputs(3522) <= layer3_outputs(5671);
    layer4_outputs(3523) <= not(layer3_outputs(6730)) or (layer3_outputs(3084));
    layer4_outputs(3524) <= layer3_outputs(559);
    layer4_outputs(3525) <= not((layer3_outputs(779)) and (layer3_outputs(4333)));
    layer4_outputs(3526) <= not(layer3_outputs(4276));
    layer4_outputs(3527) <= (layer3_outputs(6729)) or (layer3_outputs(4051));
    layer4_outputs(3528) <= not(layer3_outputs(347));
    layer4_outputs(3529) <= not(layer3_outputs(4448)) or (layer3_outputs(4630));
    layer4_outputs(3530) <= not(layer3_outputs(6151)) or (layer3_outputs(5341));
    layer4_outputs(3531) <= not((layer3_outputs(2195)) and (layer3_outputs(115)));
    layer4_outputs(3532) <= not(layer3_outputs(3318)) or (layer3_outputs(7531));
    layer4_outputs(3533) <= layer3_outputs(4555);
    layer4_outputs(3534) <= not(layer3_outputs(6202));
    layer4_outputs(3535) <= layer3_outputs(3489);
    layer4_outputs(3536) <= (layer3_outputs(5597)) or (layer3_outputs(553));
    layer4_outputs(3537) <= layer3_outputs(6344);
    layer4_outputs(3538) <= layer3_outputs(7512);
    layer4_outputs(3539) <= not(layer3_outputs(775));
    layer4_outputs(3540) <= not(layer3_outputs(994));
    layer4_outputs(3541) <= not(layer3_outputs(4903));
    layer4_outputs(3542) <= not((layer3_outputs(1556)) xor (layer3_outputs(3549)));
    layer4_outputs(3543) <= (layer3_outputs(3565)) or (layer3_outputs(2663));
    layer4_outputs(3544) <= '1';
    layer4_outputs(3545) <= (layer3_outputs(6565)) and (layer3_outputs(279));
    layer4_outputs(3546) <= not(layer3_outputs(4700)) or (layer3_outputs(854));
    layer4_outputs(3547) <= not(layer3_outputs(2752));
    layer4_outputs(3548) <= '1';
    layer4_outputs(3549) <= (layer3_outputs(5644)) or (layer3_outputs(3143));
    layer4_outputs(3550) <= not(layer3_outputs(4931));
    layer4_outputs(3551) <= not((layer3_outputs(3857)) or (layer3_outputs(3100)));
    layer4_outputs(3552) <= layer3_outputs(3589);
    layer4_outputs(3553) <= not((layer3_outputs(6956)) or (layer3_outputs(6554)));
    layer4_outputs(3554) <= (layer3_outputs(4059)) and (layer3_outputs(3246));
    layer4_outputs(3555) <= (layer3_outputs(1644)) and not (layer3_outputs(2529));
    layer4_outputs(3556) <= not((layer3_outputs(5329)) or (layer3_outputs(190)));
    layer4_outputs(3557) <= not((layer3_outputs(7041)) or (layer3_outputs(1357)));
    layer4_outputs(3558) <= not(layer3_outputs(2585)) or (layer3_outputs(2216));
    layer4_outputs(3559) <= (layer3_outputs(3178)) and not (layer3_outputs(1129));
    layer4_outputs(3560) <= not(layer3_outputs(6205));
    layer4_outputs(3561) <= not(layer3_outputs(1968));
    layer4_outputs(3562) <= not(layer3_outputs(5298));
    layer4_outputs(3563) <= (layer3_outputs(3857)) and not (layer3_outputs(6235));
    layer4_outputs(3564) <= (layer3_outputs(1919)) or (layer3_outputs(1507));
    layer4_outputs(3565) <= not(layer3_outputs(5523));
    layer4_outputs(3566) <= layer3_outputs(6507);
    layer4_outputs(3567) <= layer3_outputs(6324);
    layer4_outputs(3568) <= layer3_outputs(3987);
    layer4_outputs(3569) <= not(layer3_outputs(6681)) or (layer3_outputs(7299));
    layer4_outputs(3570) <= not((layer3_outputs(4095)) or (layer3_outputs(3382)));
    layer4_outputs(3571) <= layer3_outputs(5367);
    layer4_outputs(3572) <= not((layer3_outputs(2339)) or (layer3_outputs(3118)));
    layer4_outputs(3573) <= not(layer3_outputs(286)) or (layer3_outputs(5089));
    layer4_outputs(3574) <= not((layer3_outputs(5871)) xor (layer3_outputs(5395)));
    layer4_outputs(3575) <= layer3_outputs(6870);
    layer4_outputs(3576) <= not((layer3_outputs(7285)) and (layer3_outputs(2019)));
    layer4_outputs(3577) <= layer3_outputs(2199);
    layer4_outputs(3578) <= not(layer3_outputs(7225));
    layer4_outputs(3579) <= not((layer3_outputs(2449)) or (layer3_outputs(6115)));
    layer4_outputs(3580) <= not((layer3_outputs(6393)) or (layer3_outputs(1636)));
    layer4_outputs(3581) <= (layer3_outputs(6944)) xor (layer3_outputs(4739));
    layer4_outputs(3582) <= layer3_outputs(5621);
    layer4_outputs(3583) <= (layer3_outputs(4572)) or (layer3_outputs(7103));
    layer4_outputs(3584) <= (layer3_outputs(1599)) and not (layer3_outputs(4560));
    layer4_outputs(3585) <= not(layer3_outputs(5315));
    layer4_outputs(3586) <= '0';
    layer4_outputs(3587) <= not((layer3_outputs(2765)) and (layer3_outputs(7115)));
    layer4_outputs(3588) <= layer3_outputs(6064);
    layer4_outputs(3589) <= not(layer3_outputs(1986));
    layer4_outputs(3590) <= (layer3_outputs(2791)) and not (layer3_outputs(406));
    layer4_outputs(3591) <= not(layer3_outputs(2346));
    layer4_outputs(3592) <= layer3_outputs(2483);
    layer4_outputs(3593) <= not((layer3_outputs(6795)) and (layer3_outputs(7278)));
    layer4_outputs(3594) <= not((layer3_outputs(5579)) or (layer3_outputs(5053)));
    layer4_outputs(3595) <= layer3_outputs(4105);
    layer4_outputs(3596) <= not(layer3_outputs(7172));
    layer4_outputs(3597) <= (layer3_outputs(4316)) or (layer3_outputs(6952));
    layer4_outputs(3598) <= not((layer3_outputs(4759)) xor (layer3_outputs(5329)));
    layer4_outputs(3599) <= not(layer3_outputs(4388));
    layer4_outputs(3600) <= (layer3_outputs(4538)) or (layer3_outputs(7410));
    layer4_outputs(3601) <= (layer3_outputs(4664)) and (layer3_outputs(4081));
    layer4_outputs(3602) <= not((layer3_outputs(2967)) or (layer3_outputs(3736)));
    layer4_outputs(3603) <= not((layer3_outputs(2224)) and (layer3_outputs(4984)));
    layer4_outputs(3604) <= not((layer3_outputs(4637)) xor (layer3_outputs(4660)));
    layer4_outputs(3605) <= (layer3_outputs(6494)) and not (layer3_outputs(3793));
    layer4_outputs(3606) <= (layer3_outputs(4302)) or (layer3_outputs(604));
    layer4_outputs(3607) <= layer3_outputs(6842);
    layer4_outputs(3608) <= layer3_outputs(4738);
    layer4_outputs(3609) <= layer3_outputs(370);
    layer4_outputs(3610) <= not(layer3_outputs(6717)) or (layer3_outputs(4406));
    layer4_outputs(3611) <= not((layer3_outputs(2459)) and (layer3_outputs(6659)));
    layer4_outputs(3612) <= layer3_outputs(2456);
    layer4_outputs(3613) <= not(layer3_outputs(3073)) or (layer3_outputs(2827));
    layer4_outputs(3614) <= layer3_outputs(4720);
    layer4_outputs(3615) <= layer3_outputs(4203);
    layer4_outputs(3616) <= (layer3_outputs(3289)) and not (layer3_outputs(2048));
    layer4_outputs(3617) <= layer3_outputs(7665);
    layer4_outputs(3618) <= layer3_outputs(47);
    layer4_outputs(3619) <= (layer3_outputs(5197)) and not (layer3_outputs(2444));
    layer4_outputs(3620) <= (layer3_outputs(2241)) and (layer3_outputs(113));
    layer4_outputs(3621) <= not((layer3_outputs(3701)) or (layer3_outputs(7354)));
    layer4_outputs(3622) <= (layer3_outputs(5481)) and not (layer3_outputs(3787));
    layer4_outputs(3623) <= not((layer3_outputs(7433)) and (layer3_outputs(6379)));
    layer4_outputs(3624) <= layer3_outputs(1495);
    layer4_outputs(3625) <= not(layer3_outputs(3208));
    layer4_outputs(3626) <= (layer3_outputs(6322)) xor (layer3_outputs(3397));
    layer4_outputs(3627) <= not((layer3_outputs(6926)) or (layer3_outputs(4335)));
    layer4_outputs(3628) <= layer3_outputs(2802);
    layer4_outputs(3629) <= '1';
    layer4_outputs(3630) <= (layer3_outputs(6999)) and not (layer3_outputs(55));
    layer4_outputs(3631) <= (layer3_outputs(3462)) xor (layer3_outputs(5389));
    layer4_outputs(3632) <= not((layer3_outputs(4039)) or (layer3_outputs(7079)));
    layer4_outputs(3633) <= '0';
    layer4_outputs(3634) <= not((layer3_outputs(838)) and (layer3_outputs(6945)));
    layer4_outputs(3635) <= not((layer3_outputs(605)) xor (layer3_outputs(5214)));
    layer4_outputs(3636) <= not(layer3_outputs(6976));
    layer4_outputs(3637) <= (layer3_outputs(391)) and not (layer3_outputs(6658));
    layer4_outputs(3638) <= not(layer3_outputs(2672)) or (layer3_outputs(7123));
    layer4_outputs(3639) <= layer3_outputs(3316);
    layer4_outputs(3640) <= (layer3_outputs(1313)) and not (layer3_outputs(1239));
    layer4_outputs(3641) <= not(layer3_outputs(264));
    layer4_outputs(3642) <= (layer3_outputs(276)) and not (layer3_outputs(3839));
    layer4_outputs(3643) <= not((layer3_outputs(3551)) and (layer3_outputs(2784)));
    layer4_outputs(3644) <= (layer3_outputs(6107)) and not (layer3_outputs(2013));
    layer4_outputs(3645) <= (layer3_outputs(880)) or (layer3_outputs(2004));
    layer4_outputs(3646) <= not(layer3_outputs(5762)) or (layer3_outputs(1132));
    layer4_outputs(3647) <= not((layer3_outputs(6205)) and (layer3_outputs(6664)));
    layer4_outputs(3648) <= not(layer3_outputs(6927));
    layer4_outputs(3649) <= not(layer3_outputs(6992)) or (layer3_outputs(1804));
    layer4_outputs(3650) <= (layer3_outputs(4813)) and not (layer3_outputs(2988));
    layer4_outputs(3651) <= not(layer3_outputs(803));
    layer4_outputs(3652) <= '0';
    layer4_outputs(3653) <= not((layer3_outputs(4029)) xor (layer3_outputs(5986)));
    layer4_outputs(3654) <= '0';
    layer4_outputs(3655) <= not(layer3_outputs(7675)) or (layer3_outputs(5421));
    layer4_outputs(3656) <= not(layer3_outputs(4108));
    layer4_outputs(3657) <= layer3_outputs(2392);
    layer4_outputs(3658) <= not((layer3_outputs(3174)) and (layer3_outputs(3080)));
    layer4_outputs(3659) <= layer3_outputs(220);
    layer4_outputs(3660) <= '0';
    layer4_outputs(3661) <= not(layer3_outputs(1526)) or (layer3_outputs(4524));
    layer4_outputs(3662) <= layer3_outputs(3004);
    layer4_outputs(3663) <= not(layer3_outputs(4687));
    layer4_outputs(3664) <= not(layer3_outputs(877));
    layer4_outputs(3665) <= not(layer3_outputs(2214)) or (layer3_outputs(5828));
    layer4_outputs(3666) <= layer3_outputs(4141);
    layer4_outputs(3667) <= (layer3_outputs(1540)) and not (layer3_outputs(271));
    layer4_outputs(3668) <= layer3_outputs(5737);
    layer4_outputs(3669) <= layer3_outputs(5684);
    layer4_outputs(3670) <= not(layer3_outputs(6044));
    layer4_outputs(3671) <= not((layer3_outputs(355)) or (layer3_outputs(4378)));
    layer4_outputs(3672) <= (layer3_outputs(5569)) or (layer3_outputs(4408));
    layer4_outputs(3673) <= (layer3_outputs(2674)) and (layer3_outputs(1328));
    layer4_outputs(3674) <= '1';
    layer4_outputs(3675) <= '1';
    layer4_outputs(3676) <= not((layer3_outputs(742)) or (layer3_outputs(1047)));
    layer4_outputs(3677) <= (layer3_outputs(6903)) or (layer3_outputs(2504));
    layer4_outputs(3678) <= not(layer3_outputs(6077)) or (layer3_outputs(1679));
    layer4_outputs(3679) <= (layer3_outputs(5026)) or (layer3_outputs(4200));
    layer4_outputs(3680) <= not(layer3_outputs(1854));
    layer4_outputs(3681) <= not(layer3_outputs(5866)) or (layer3_outputs(7301));
    layer4_outputs(3682) <= layer3_outputs(1887);
    layer4_outputs(3683) <= layer3_outputs(212);
    layer4_outputs(3684) <= (layer3_outputs(6396)) and not (layer3_outputs(6378));
    layer4_outputs(3685) <= (layer3_outputs(4835)) or (layer3_outputs(4574));
    layer4_outputs(3686) <= (layer3_outputs(1479)) and (layer3_outputs(6939));
    layer4_outputs(3687) <= (layer3_outputs(6088)) or (layer3_outputs(3927));
    layer4_outputs(3688) <= not(layer3_outputs(4617)) or (layer3_outputs(4529));
    layer4_outputs(3689) <= not((layer3_outputs(6070)) xor (layer3_outputs(5559)));
    layer4_outputs(3690) <= (layer3_outputs(6381)) xor (layer3_outputs(4357));
    layer4_outputs(3691) <= (layer3_outputs(6577)) xor (layer3_outputs(613));
    layer4_outputs(3692) <= (layer3_outputs(4643)) and (layer3_outputs(592));
    layer4_outputs(3693) <= not((layer3_outputs(6706)) or (layer3_outputs(3585)));
    layer4_outputs(3694) <= not(layer3_outputs(3216));
    layer4_outputs(3695) <= '1';
    layer4_outputs(3696) <= layer3_outputs(5045);
    layer4_outputs(3697) <= (layer3_outputs(1136)) and not (layer3_outputs(7349));
    layer4_outputs(3698) <= (layer3_outputs(3237)) xor (layer3_outputs(6132));
    layer4_outputs(3699) <= (layer3_outputs(6102)) xor (layer3_outputs(2155));
    layer4_outputs(3700) <= not((layer3_outputs(5611)) and (layer3_outputs(6855)));
    layer4_outputs(3701) <= not(layer3_outputs(1788));
    layer4_outputs(3702) <= layer3_outputs(968);
    layer4_outputs(3703) <= not((layer3_outputs(3310)) or (layer3_outputs(5176)));
    layer4_outputs(3704) <= (layer3_outputs(3914)) or (layer3_outputs(4793));
    layer4_outputs(3705) <= not(layer3_outputs(319)) or (layer3_outputs(2233));
    layer4_outputs(3706) <= not((layer3_outputs(3944)) or (layer3_outputs(203)));
    layer4_outputs(3707) <= (layer3_outputs(3799)) or (layer3_outputs(5217));
    layer4_outputs(3708) <= (layer3_outputs(870)) and not (layer3_outputs(6777));
    layer4_outputs(3709) <= '1';
    layer4_outputs(3710) <= (layer3_outputs(3437)) and not (layer3_outputs(3361));
    layer4_outputs(3711) <= not((layer3_outputs(2250)) or (layer3_outputs(318)));
    layer4_outputs(3712) <= not(layer3_outputs(1863));
    layer4_outputs(3713) <= (layer3_outputs(6299)) or (layer3_outputs(6793));
    layer4_outputs(3714) <= layer3_outputs(678);
    layer4_outputs(3715) <= (layer3_outputs(5149)) and (layer3_outputs(2575));
    layer4_outputs(3716) <= not(layer3_outputs(6510));
    layer4_outputs(3717) <= layer3_outputs(3598);
    layer4_outputs(3718) <= (layer3_outputs(1545)) or (layer3_outputs(2246));
    layer4_outputs(3719) <= (layer3_outputs(2747)) or (layer3_outputs(609));
    layer4_outputs(3720) <= (layer3_outputs(5426)) and not (layer3_outputs(6465));
    layer4_outputs(3721) <= layer3_outputs(7516);
    layer4_outputs(3722) <= not(layer3_outputs(3378));
    layer4_outputs(3723) <= not(layer3_outputs(4168));
    layer4_outputs(3724) <= '1';
    layer4_outputs(3725) <= (layer3_outputs(1746)) xor (layer3_outputs(2234));
    layer4_outputs(3726) <= layer3_outputs(5217);
    layer4_outputs(3727) <= not(layer3_outputs(5727));
    layer4_outputs(3728) <= not((layer3_outputs(7042)) xor (layer3_outputs(1446)));
    layer4_outputs(3729) <= not((layer3_outputs(976)) and (layer3_outputs(3668)));
    layer4_outputs(3730) <= not(layer3_outputs(5865)) or (layer3_outputs(6673));
    layer4_outputs(3731) <= not((layer3_outputs(748)) or (layer3_outputs(4536)));
    layer4_outputs(3732) <= (layer3_outputs(917)) and not (layer3_outputs(3452));
    layer4_outputs(3733) <= not(layer3_outputs(6551));
    layer4_outputs(3734) <= (layer3_outputs(7365)) or (layer3_outputs(5698));
    layer4_outputs(3735) <= not((layer3_outputs(3531)) or (layer3_outputs(1217)));
    layer4_outputs(3736) <= not(layer3_outputs(554));
    layer4_outputs(3737) <= layer3_outputs(1629);
    layer4_outputs(3738) <= not(layer3_outputs(1812));
    layer4_outputs(3739) <= (layer3_outputs(990)) or (layer3_outputs(1834));
    layer4_outputs(3740) <= (layer3_outputs(2240)) and (layer3_outputs(2993));
    layer4_outputs(3741) <= '1';
    layer4_outputs(3742) <= layer3_outputs(1551);
    layer4_outputs(3743) <= not((layer3_outputs(2573)) or (layer3_outputs(2897)));
    layer4_outputs(3744) <= not(layer3_outputs(5330)) or (layer3_outputs(2629));
    layer4_outputs(3745) <= layer3_outputs(808);
    layer4_outputs(3746) <= layer3_outputs(4805);
    layer4_outputs(3747) <= not((layer3_outputs(449)) xor (layer3_outputs(6062)));
    layer4_outputs(3748) <= not(layer3_outputs(58));
    layer4_outputs(3749) <= not(layer3_outputs(3479));
    layer4_outputs(3750) <= not(layer3_outputs(5877));
    layer4_outputs(3751) <= not(layer3_outputs(1066));
    layer4_outputs(3752) <= not(layer3_outputs(3555));
    layer4_outputs(3753) <= not(layer3_outputs(5556)) or (layer3_outputs(870));
    layer4_outputs(3754) <= not((layer3_outputs(6954)) or (layer3_outputs(6563)));
    layer4_outputs(3755) <= layer3_outputs(235);
    layer4_outputs(3756) <= (layer3_outputs(7036)) and not (layer3_outputs(2058));
    layer4_outputs(3757) <= not(layer3_outputs(2711));
    layer4_outputs(3758) <= layer3_outputs(2433);
    layer4_outputs(3759) <= not((layer3_outputs(6252)) or (layer3_outputs(1380)));
    layer4_outputs(3760) <= not((layer3_outputs(7008)) xor (layer3_outputs(7520)));
    layer4_outputs(3761) <= layer3_outputs(966);
    layer4_outputs(3762) <= (layer3_outputs(4291)) and not (layer3_outputs(3953));
    layer4_outputs(3763) <= not(layer3_outputs(4344));
    layer4_outputs(3764) <= not(layer3_outputs(4155));
    layer4_outputs(3765) <= not(layer3_outputs(1854));
    layer4_outputs(3766) <= not(layer3_outputs(7320));
    layer4_outputs(3767) <= not(layer3_outputs(4898));
    layer4_outputs(3768) <= (layer3_outputs(7011)) and not (layer3_outputs(574));
    layer4_outputs(3769) <= layer3_outputs(3330);
    layer4_outputs(3770) <= '0';
    layer4_outputs(3771) <= not(layer3_outputs(1270)) or (layer3_outputs(3626));
    layer4_outputs(3772) <= not(layer3_outputs(7283));
    layer4_outputs(3773) <= not(layer3_outputs(3818)) or (layer3_outputs(958));
    layer4_outputs(3774) <= layer3_outputs(4109);
    layer4_outputs(3775) <= (layer3_outputs(2267)) xor (layer3_outputs(2621));
    layer4_outputs(3776) <= (layer3_outputs(1068)) and (layer3_outputs(6675));
    layer4_outputs(3777) <= not(layer3_outputs(113));
    layer4_outputs(3778) <= (layer3_outputs(7333)) and not (layer3_outputs(5391));
    layer4_outputs(3779) <= not(layer3_outputs(467)) or (layer3_outputs(4443));
    layer4_outputs(3780) <= (layer3_outputs(465)) and not (layer3_outputs(4888));
    layer4_outputs(3781) <= layer3_outputs(5956);
    layer4_outputs(3782) <= '1';
    layer4_outputs(3783) <= (layer3_outputs(3613)) and (layer3_outputs(2070));
    layer4_outputs(3784) <= layer3_outputs(6594);
    layer4_outputs(3785) <= not((layer3_outputs(953)) xor (layer3_outputs(6811)));
    layer4_outputs(3786) <= layer3_outputs(222);
    layer4_outputs(3787) <= not((layer3_outputs(4132)) and (layer3_outputs(7414)));
    layer4_outputs(3788) <= '1';
    layer4_outputs(3789) <= (layer3_outputs(6775)) or (layer3_outputs(5842));
    layer4_outputs(3790) <= layer3_outputs(7438);
    layer4_outputs(3791) <= (layer3_outputs(160)) and (layer3_outputs(408));
    layer4_outputs(3792) <= (layer3_outputs(807)) and (layer3_outputs(6726));
    layer4_outputs(3793) <= not(layer3_outputs(2498));
    layer4_outputs(3794) <= (layer3_outputs(3162)) and (layer3_outputs(4994));
    layer4_outputs(3795) <= not((layer3_outputs(2926)) or (layer3_outputs(4749)));
    layer4_outputs(3796) <= (layer3_outputs(5375)) and not (layer3_outputs(3931));
    layer4_outputs(3797) <= not((layer3_outputs(1724)) and (layer3_outputs(6936)));
    layer4_outputs(3798) <= not(layer3_outputs(1634)) or (layer3_outputs(7636));
    layer4_outputs(3799) <= '1';
    layer4_outputs(3800) <= layer3_outputs(2031);
    layer4_outputs(3801) <= (layer3_outputs(3481)) or (layer3_outputs(12));
    layer4_outputs(3802) <= '1';
    layer4_outputs(3803) <= (layer3_outputs(6998)) xor (layer3_outputs(4918));
    layer4_outputs(3804) <= (layer3_outputs(5707)) or (layer3_outputs(4676));
    layer4_outputs(3805) <= (layer3_outputs(3091)) or (layer3_outputs(1658));
    layer4_outputs(3806) <= not(layer3_outputs(6607)) or (layer3_outputs(4870));
    layer4_outputs(3807) <= not(layer3_outputs(1933));
    layer4_outputs(3808) <= (layer3_outputs(5630)) and not (layer3_outputs(1449));
    layer4_outputs(3809) <= not(layer3_outputs(5682));
    layer4_outputs(3810) <= layer3_outputs(2867);
    layer4_outputs(3811) <= layer3_outputs(5648);
    layer4_outputs(3812) <= (layer3_outputs(1103)) xor (layer3_outputs(753));
    layer4_outputs(3813) <= not(layer3_outputs(6391));
    layer4_outputs(3814) <= (layer3_outputs(3526)) xor (layer3_outputs(3845));
    layer4_outputs(3815) <= not((layer3_outputs(7111)) or (layer3_outputs(4515)));
    layer4_outputs(3816) <= not(layer3_outputs(1022));
    layer4_outputs(3817) <= (layer3_outputs(3975)) and not (layer3_outputs(86));
    layer4_outputs(3818) <= not((layer3_outputs(3106)) or (layer3_outputs(3405)));
    layer4_outputs(3819) <= layer3_outputs(1518);
    layer4_outputs(3820) <= layer3_outputs(6242);
    layer4_outputs(3821) <= '1';
    layer4_outputs(3822) <= (layer3_outputs(767)) and not (layer3_outputs(1696));
    layer4_outputs(3823) <= not((layer3_outputs(6528)) and (layer3_outputs(1490)));
    layer4_outputs(3824) <= (layer3_outputs(3466)) and not (layer3_outputs(2213));
    layer4_outputs(3825) <= (layer3_outputs(1154)) and not (layer3_outputs(4069));
    layer4_outputs(3826) <= (layer3_outputs(5369)) and not (layer3_outputs(4180));
    layer4_outputs(3827) <= layer3_outputs(906);
    layer4_outputs(3828) <= not(layer3_outputs(1463)) or (layer3_outputs(6267));
    layer4_outputs(3829) <= (layer3_outputs(364)) and not (layer3_outputs(6462));
    layer4_outputs(3830) <= not(layer3_outputs(6419));
    layer4_outputs(3831) <= layer3_outputs(2201);
    layer4_outputs(3832) <= not(layer3_outputs(419)) or (layer3_outputs(5566));
    layer4_outputs(3833) <= (layer3_outputs(4193)) or (layer3_outputs(7484));
    layer4_outputs(3834) <= not((layer3_outputs(440)) xor (layer3_outputs(6506)));
    layer4_outputs(3835) <= not((layer3_outputs(3107)) and (layer3_outputs(1062)));
    layer4_outputs(3836) <= '1';
    layer4_outputs(3837) <= (layer3_outputs(1688)) and (layer3_outputs(4828));
    layer4_outputs(3838) <= layer3_outputs(5840);
    layer4_outputs(3839) <= (layer3_outputs(4986)) and not (layer3_outputs(1762));
    layer4_outputs(3840) <= not(layer3_outputs(4319));
    layer4_outputs(3841) <= '1';
    layer4_outputs(3842) <= '0';
    layer4_outputs(3843) <= not((layer3_outputs(649)) or (layer3_outputs(2278)));
    layer4_outputs(3844) <= (layer3_outputs(4144)) and not (layer3_outputs(4946));
    layer4_outputs(3845) <= not(layer3_outputs(3459));
    layer4_outputs(3846) <= not(layer3_outputs(235)) or (layer3_outputs(3305));
    layer4_outputs(3847) <= not(layer3_outputs(5755));
    layer4_outputs(3848) <= (layer3_outputs(5905)) and not (layer3_outputs(1975));
    layer4_outputs(3849) <= layer3_outputs(1765);
    layer4_outputs(3850) <= not(layer3_outputs(2329)) or (layer3_outputs(5451));
    layer4_outputs(3851) <= layer3_outputs(1077);
    layer4_outputs(3852) <= not(layer3_outputs(1630));
    layer4_outputs(3853) <= (layer3_outputs(7537)) and not (layer3_outputs(2611));
    layer4_outputs(3854) <= layer3_outputs(3104);
    layer4_outputs(3855) <= '1';
    layer4_outputs(3856) <= (layer3_outputs(2565)) and (layer3_outputs(1222));
    layer4_outputs(3857) <= (layer3_outputs(1876)) and (layer3_outputs(4303));
    layer4_outputs(3858) <= not(layer3_outputs(3895));
    layer4_outputs(3859) <= not((layer3_outputs(7551)) or (layer3_outputs(3484)));
    layer4_outputs(3860) <= layer3_outputs(5795);
    layer4_outputs(3861) <= not(layer3_outputs(5031));
    layer4_outputs(3862) <= not(layer3_outputs(3287));
    layer4_outputs(3863) <= not(layer3_outputs(4710)) or (layer3_outputs(2));
    layer4_outputs(3864) <= not(layer3_outputs(3335));
    layer4_outputs(3865) <= not(layer3_outputs(2059)) or (layer3_outputs(442));
    layer4_outputs(3866) <= not(layer3_outputs(4227)) or (layer3_outputs(3510));
    layer4_outputs(3867) <= not(layer3_outputs(601));
    layer4_outputs(3868) <= not((layer3_outputs(3839)) xor (layer3_outputs(4775)));
    layer4_outputs(3869) <= not(layer3_outputs(6816));
    layer4_outputs(3870) <= (layer3_outputs(2389)) and not (layer3_outputs(3646));
    layer4_outputs(3871) <= (layer3_outputs(1824)) and not (layer3_outputs(4511));
    layer4_outputs(3872) <= layer3_outputs(6645);
    layer4_outputs(3873) <= layer3_outputs(4725);
    layer4_outputs(3874) <= (layer3_outputs(5065)) and (layer3_outputs(1665));
    layer4_outputs(3875) <= not(layer3_outputs(3668)) or (layer3_outputs(3071));
    layer4_outputs(3876) <= not((layer3_outputs(145)) or (layer3_outputs(5441)));
    layer4_outputs(3877) <= layer3_outputs(1572);
    layer4_outputs(3878) <= not((layer3_outputs(483)) and (layer3_outputs(3643)));
    layer4_outputs(3879) <= not((layer3_outputs(5497)) and (layer3_outputs(5919)));
    layer4_outputs(3880) <= not(layer3_outputs(7565));
    layer4_outputs(3881) <= (layer3_outputs(1326)) and not (layer3_outputs(1061));
    layer4_outputs(3882) <= not((layer3_outputs(5018)) or (layer3_outputs(6552)));
    layer4_outputs(3883) <= not((layer3_outputs(4032)) or (layer3_outputs(37)));
    layer4_outputs(3884) <= not((layer3_outputs(2235)) and (layer3_outputs(289)));
    layer4_outputs(3885) <= not(layer3_outputs(4456)) or (layer3_outputs(4042));
    layer4_outputs(3886) <= not(layer3_outputs(6276));
    layer4_outputs(3887) <= not(layer3_outputs(6603));
    layer4_outputs(3888) <= '1';
    layer4_outputs(3889) <= not((layer3_outputs(4147)) xor (layer3_outputs(5696)));
    layer4_outputs(3890) <= not((layer3_outputs(3188)) and (layer3_outputs(7308)));
    layer4_outputs(3891) <= not(layer3_outputs(75)) or (layer3_outputs(1541));
    layer4_outputs(3892) <= (layer3_outputs(1261)) and not (layer3_outputs(3976));
    layer4_outputs(3893) <= (layer3_outputs(5332)) and (layer3_outputs(7422));
    layer4_outputs(3894) <= (layer3_outputs(3865)) or (layer3_outputs(298));
    layer4_outputs(3895) <= (layer3_outputs(2601)) and not (layer3_outputs(960));
    layer4_outputs(3896) <= layer3_outputs(3850);
    layer4_outputs(3897) <= layer3_outputs(6226);
    layer4_outputs(3898) <= not(layer3_outputs(1857));
    layer4_outputs(3899) <= not(layer3_outputs(5119));
    layer4_outputs(3900) <= '1';
    layer4_outputs(3901) <= layer3_outputs(6656);
    layer4_outputs(3902) <= layer3_outputs(7658);
    layer4_outputs(3903) <= layer3_outputs(7325);
    layer4_outputs(3904) <= not(layer3_outputs(4065));
    layer4_outputs(3905) <= layer3_outputs(7443);
    layer4_outputs(3906) <= (layer3_outputs(1738)) or (layer3_outputs(7222));
    layer4_outputs(3907) <= not(layer3_outputs(2695));
    layer4_outputs(3908) <= layer3_outputs(2423);
    layer4_outputs(3909) <= layer3_outputs(5408);
    layer4_outputs(3910) <= '1';
    layer4_outputs(3911) <= layer3_outputs(662);
    layer4_outputs(3912) <= layer3_outputs(769);
    layer4_outputs(3913) <= not(layer3_outputs(3409));
    layer4_outputs(3914) <= '1';
    layer4_outputs(3915) <= not(layer3_outputs(1678));
    layer4_outputs(3916) <= not(layer3_outputs(3850));
    layer4_outputs(3917) <= layer3_outputs(2811);
    layer4_outputs(3918) <= not(layer3_outputs(1321));
    layer4_outputs(3919) <= not((layer3_outputs(6486)) xor (layer3_outputs(664)));
    layer4_outputs(3920) <= not((layer3_outputs(3420)) and (layer3_outputs(2761)));
    layer4_outputs(3921) <= '1';
    layer4_outputs(3922) <= (layer3_outputs(2000)) xor (layer3_outputs(1446));
    layer4_outputs(3923) <= not(layer3_outputs(3297)) or (layer3_outputs(2594));
    layer4_outputs(3924) <= '0';
    layer4_outputs(3925) <= not((layer3_outputs(5715)) xor (layer3_outputs(3699)));
    layer4_outputs(3926) <= not(layer3_outputs(6969));
    layer4_outputs(3927) <= not(layer3_outputs(6690)) or (layer3_outputs(2607));
    layer4_outputs(3928) <= not((layer3_outputs(5820)) and (layer3_outputs(5656)));
    layer4_outputs(3929) <= (layer3_outputs(4992)) or (layer3_outputs(3747));
    layer4_outputs(3930) <= '1';
    layer4_outputs(3931) <= (layer3_outputs(5618)) or (layer3_outputs(2545));
    layer4_outputs(3932) <= not(layer3_outputs(1571));
    layer4_outputs(3933) <= not(layer3_outputs(254)) or (layer3_outputs(5575));
    layer4_outputs(3934) <= not(layer3_outputs(2684)) or (layer3_outputs(211));
    layer4_outputs(3935) <= not(layer3_outputs(3816));
    layer4_outputs(3936) <= layer3_outputs(3009);
    layer4_outputs(3937) <= not(layer3_outputs(3804));
    layer4_outputs(3938) <= not(layer3_outputs(3988));
    layer4_outputs(3939) <= not(layer3_outputs(1070));
    layer4_outputs(3940) <= layer3_outputs(2523);
    layer4_outputs(3941) <= (layer3_outputs(2318)) xor (layer3_outputs(7643));
    layer4_outputs(3942) <= not((layer3_outputs(5869)) or (layer3_outputs(1198)));
    layer4_outputs(3943) <= layer3_outputs(545);
    layer4_outputs(3944) <= '0';
    layer4_outputs(3945) <= not((layer3_outputs(7586)) xor (layer3_outputs(4626)));
    layer4_outputs(3946) <= (layer3_outputs(3003)) and (layer3_outputs(2539));
    layer4_outputs(3947) <= '0';
    layer4_outputs(3948) <= not(layer3_outputs(1274));
    layer4_outputs(3949) <= not((layer3_outputs(3886)) xor (layer3_outputs(5034)));
    layer4_outputs(3950) <= (layer3_outputs(7547)) and not (layer3_outputs(3324));
    layer4_outputs(3951) <= not((layer3_outputs(2874)) or (layer3_outputs(3609)));
    layer4_outputs(3952) <= not(layer3_outputs(6556)) or (layer3_outputs(3057));
    layer4_outputs(3953) <= layer3_outputs(6615);
    layer4_outputs(3954) <= not((layer3_outputs(6278)) and (layer3_outputs(5977)));
    layer4_outputs(3955) <= (layer3_outputs(2116)) and (layer3_outputs(6498));
    layer4_outputs(3956) <= not((layer3_outputs(3000)) xor (layer3_outputs(1128)));
    layer4_outputs(3957) <= not((layer3_outputs(1315)) or (layer3_outputs(3033)));
    layer4_outputs(3958) <= (layer3_outputs(1704)) or (layer3_outputs(3214));
    layer4_outputs(3959) <= layer3_outputs(1841);
    layer4_outputs(3960) <= not(layer3_outputs(5528));
    layer4_outputs(3961) <= (layer3_outputs(1041)) and not (layer3_outputs(3279));
    layer4_outputs(3962) <= not((layer3_outputs(5945)) and (layer3_outputs(4422)));
    layer4_outputs(3963) <= not((layer3_outputs(6858)) and (layer3_outputs(5902)));
    layer4_outputs(3964) <= '0';
    layer4_outputs(3965) <= layer3_outputs(5067);
    layer4_outputs(3966) <= (layer3_outputs(2115)) and not (layer3_outputs(6423));
    layer4_outputs(3967) <= (layer3_outputs(4025)) and not (layer3_outputs(162));
    layer4_outputs(3968) <= '1';
    layer4_outputs(3969) <= not(layer3_outputs(2561));
    layer4_outputs(3970) <= not(layer3_outputs(5837));
    layer4_outputs(3971) <= not(layer3_outputs(5216));
    layer4_outputs(3972) <= not(layer3_outputs(7073)) or (layer3_outputs(650));
    layer4_outputs(3973) <= not(layer3_outputs(4903));
    layer4_outputs(3974) <= not(layer3_outputs(3870));
    layer4_outputs(3975) <= (layer3_outputs(3935)) and (layer3_outputs(2141));
    layer4_outputs(3976) <= layer3_outputs(1866);
    layer4_outputs(3977) <= not((layer3_outputs(2478)) or (layer3_outputs(2281)));
    layer4_outputs(3978) <= (layer3_outputs(6698)) and not (layer3_outputs(6513));
    layer4_outputs(3979) <= not((layer3_outputs(67)) and (layer3_outputs(3265)));
    layer4_outputs(3980) <= (layer3_outputs(6696)) and (layer3_outputs(4071));
    layer4_outputs(3981) <= layer3_outputs(7356);
    layer4_outputs(3982) <= not(layer3_outputs(3495));
    layer4_outputs(3983) <= layer3_outputs(2889);
    layer4_outputs(3984) <= not(layer3_outputs(2960));
    layer4_outputs(3985) <= layer3_outputs(5949);
    layer4_outputs(3986) <= '1';
    layer4_outputs(3987) <= (layer3_outputs(6374)) or (layer3_outputs(5623));
    layer4_outputs(3988) <= not(layer3_outputs(2229)) or (layer3_outputs(4198));
    layer4_outputs(3989) <= not(layer3_outputs(1664));
    layer4_outputs(3990) <= not(layer3_outputs(4243));
    layer4_outputs(3991) <= (layer3_outputs(5967)) xor (layer3_outputs(2784));
    layer4_outputs(3992) <= not((layer3_outputs(7332)) and (layer3_outputs(368)));
    layer4_outputs(3993) <= (layer3_outputs(947)) and not (layer3_outputs(3349));
    layer4_outputs(3994) <= not((layer3_outputs(3050)) or (layer3_outputs(1812)));
    layer4_outputs(3995) <= not(layer3_outputs(6628));
    layer4_outputs(3996) <= not(layer3_outputs(1030)) or (layer3_outputs(4046));
    layer4_outputs(3997) <= not(layer3_outputs(5445));
    layer4_outputs(3998) <= not((layer3_outputs(4873)) and (layer3_outputs(3604)));
    layer4_outputs(3999) <= not(layer3_outputs(1520));
    layer4_outputs(4000) <= (layer3_outputs(3232)) and not (layer3_outputs(5393));
    layer4_outputs(4001) <= not((layer3_outputs(378)) or (layer3_outputs(5772)));
    layer4_outputs(4002) <= not(layer3_outputs(1884)) or (layer3_outputs(6478));
    layer4_outputs(4003) <= not(layer3_outputs(1864));
    layer4_outputs(4004) <= not((layer3_outputs(1603)) and (layer3_outputs(6048)));
    layer4_outputs(4005) <= not((layer3_outputs(7034)) and (layer3_outputs(7274)));
    layer4_outputs(4006) <= (layer3_outputs(6945)) and (layer3_outputs(4716));
    layer4_outputs(4007) <= not((layer3_outputs(3456)) and (layer3_outputs(2664)));
    layer4_outputs(4008) <= layer3_outputs(2025);
    layer4_outputs(4009) <= layer3_outputs(6631);
    layer4_outputs(4010) <= not(layer3_outputs(2089));
    layer4_outputs(4011) <= not(layer3_outputs(4822));
    layer4_outputs(4012) <= (layer3_outputs(151)) and not (layer3_outputs(5875));
    layer4_outputs(4013) <= layer3_outputs(5442);
    layer4_outputs(4014) <= layer3_outputs(1145);
    layer4_outputs(4015) <= not(layer3_outputs(4684)) or (layer3_outputs(6911));
    layer4_outputs(4016) <= not(layer3_outputs(7347)) or (layer3_outputs(570));
    layer4_outputs(4017) <= (layer3_outputs(5786)) and (layer3_outputs(3502));
    layer4_outputs(4018) <= layer3_outputs(6182);
    layer4_outputs(4019) <= '1';
    layer4_outputs(4020) <= not(layer3_outputs(5493)) or (layer3_outputs(6124));
    layer4_outputs(4021) <= not(layer3_outputs(4132));
    layer4_outputs(4022) <= layer3_outputs(2446);
    layer4_outputs(4023) <= layer3_outputs(34);
    layer4_outputs(4024) <= (layer3_outputs(4018)) or (layer3_outputs(1807));
    layer4_outputs(4025) <= (layer3_outputs(2332)) and (layer3_outputs(1503));
    layer4_outputs(4026) <= '0';
    layer4_outputs(4027) <= (layer3_outputs(6470)) and (layer3_outputs(1394));
    layer4_outputs(4028) <= not(layer3_outputs(1236));
    layer4_outputs(4029) <= layer3_outputs(2743);
    layer4_outputs(4030) <= not(layer3_outputs(2387));
    layer4_outputs(4031) <= not(layer3_outputs(2070)) or (layer3_outputs(4520));
    layer4_outputs(4032) <= not(layer3_outputs(3459)) or (layer3_outputs(4472));
    layer4_outputs(4033) <= '1';
    layer4_outputs(4034) <= not((layer3_outputs(3961)) and (layer3_outputs(851)));
    layer4_outputs(4035) <= layer3_outputs(6733);
    layer4_outputs(4036) <= (layer3_outputs(6608)) and not (layer3_outputs(6188));
    layer4_outputs(4037) <= not(layer3_outputs(855)) or (layer3_outputs(3567));
    layer4_outputs(4038) <= layer3_outputs(3649);
    layer4_outputs(4039) <= not(layer3_outputs(6663)) or (layer3_outputs(1706));
    layer4_outputs(4040) <= layer3_outputs(2497);
    layer4_outputs(4041) <= layer3_outputs(1460);
    layer4_outputs(4042) <= not((layer3_outputs(1179)) and (layer3_outputs(6519)));
    layer4_outputs(4043) <= layer3_outputs(1515);
    layer4_outputs(4044) <= (layer3_outputs(874)) xor (layer3_outputs(4788));
    layer4_outputs(4045) <= layer3_outputs(6411);
    layer4_outputs(4046) <= not(layer3_outputs(4180));
    layer4_outputs(4047) <= (layer3_outputs(4141)) and not (layer3_outputs(5900));
    layer4_outputs(4048) <= '1';
    layer4_outputs(4049) <= (layer3_outputs(6509)) and not (layer3_outputs(798));
    layer4_outputs(4050) <= not((layer3_outputs(3146)) and (layer3_outputs(1286)));
    layer4_outputs(4051) <= not(layer3_outputs(3277));
    layer4_outputs(4052) <= not((layer3_outputs(5326)) xor (layer3_outputs(112)));
    layer4_outputs(4053) <= not(layer3_outputs(4761)) or (layer3_outputs(2120));
    layer4_outputs(4054) <= not(layer3_outputs(6006));
    layer4_outputs(4055) <= not(layer3_outputs(457));
    layer4_outputs(4056) <= layer3_outputs(7592);
    layer4_outputs(4057) <= (layer3_outputs(854)) xor (layer3_outputs(1164));
    layer4_outputs(4058) <= layer3_outputs(7542);
    layer4_outputs(4059) <= layer3_outputs(2164);
    layer4_outputs(4060) <= not((layer3_outputs(3142)) and (layer3_outputs(5477)));
    layer4_outputs(4061) <= not(layer3_outputs(1223)) or (layer3_outputs(7648));
    layer4_outputs(4062) <= layer3_outputs(4507);
    layer4_outputs(4063) <= not(layer3_outputs(3306)) or (layer3_outputs(7146));
    layer4_outputs(4064) <= (layer3_outputs(4785)) and not (layer3_outputs(2609));
    layer4_outputs(4065) <= not(layer3_outputs(986));
    layer4_outputs(4066) <= not((layer3_outputs(2067)) or (layer3_outputs(2978)));
    layer4_outputs(4067) <= layer3_outputs(1089);
    layer4_outputs(4068) <= not(layer3_outputs(2000));
    layer4_outputs(4069) <= (layer3_outputs(3761)) or (layer3_outputs(4117));
    layer4_outputs(4070) <= not(layer3_outputs(3778)) or (layer3_outputs(331));
    layer4_outputs(4071) <= '0';
    layer4_outputs(4072) <= (layer3_outputs(4083)) and (layer3_outputs(2902));
    layer4_outputs(4073) <= layer3_outputs(3858);
    layer4_outputs(4074) <= not(layer3_outputs(1417));
    layer4_outputs(4075) <= (layer3_outputs(5015)) xor (layer3_outputs(4425));
    layer4_outputs(4076) <= layer3_outputs(3040);
    layer4_outputs(4077) <= (layer3_outputs(5377)) xor (layer3_outputs(1539));
    layer4_outputs(4078) <= layer3_outputs(1728);
    layer4_outputs(4079) <= not((layer3_outputs(3546)) or (layer3_outputs(1418)));
    layer4_outputs(4080) <= (layer3_outputs(7535)) and not (layer3_outputs(6985));
    layer4_outputs(4081) <= not(layer3_outputs(2917));
    layer4_outputs(4082) <= not((layer3_outputs(6568)) and (layer3_outputs(4237)));
    layer4_outputs(4083) <= layer3_outputs(3723);
    layer4_outputs(4084) <= (layer3_outputs(275)) and not (layer3_outputs(4836));
    layer4_outputs(4085) <= '1';
    layer4_outputs(4086) <= (layer3_outputs(7003)) or (layer3_outputs(7211));
    layer4_outputs(4087) <= not(layer3_outputs(4127));
    layer4_outputs(4088) <= not(layer3_outputs(2026));
    layer4_outputs(4089) <= not(layer3_outputs(4377)) or (layer3_outputs(6409));
    layer4_outputs(4090) <= not((layer3_outputs(7518)) and (layer3_outputs(4295)));
    layer4_outputs(4091) <= '1';
    layer4_outputs(4092) <= layer3_outputs(3639);
    layer4_outputs(4093) <= not(layer3_outputs(144));
    layer4_outputs(4094) <= layer3_outputs(935);
    layer4_outputs(4095) <= layer3_outputs(886);
    layer4_outputs(4096) <= (layer3_outputs(3520)) xor (layer3_outputs(4098));
    layer4_outputs(4097) <= not(layer3_outputs(7176));
    layer4_outputs(4098) <= (layer3_outputs(6147)) and not (layer3_outputs(265));
    layer4_outputs(4099) <= not(layer3_outputs(794));
    layer4_outputs(4100) <= layer3_outputs(3450);
    layer4_outputs(4101) <= not((layer3_outputs(2844)) or (layer3_outputs(4019)));
    layer4_outputs(4102) <= not(layer3_outputs(3402));
    layer4_outputs(4103) <= not(layer3_outputs(7238));
    layer4_outputs(4104) <= layer3_outputs(6666);
    layer4_outputs(4105) <= not(layer3_outputs(3755)) or (layer3_outputs(3312));
    layer4_outputs(4106) <= '0';
    layer4_outputs(4107) <= not(layer3_outputs(4850));
    layer4_outputs(4108) <= not(layer3_outputs(6247)) or (layer3_outputs(6930));
    layer4_outputs(4109) <= (layer3_outputs(5443)) and (layer3_outputs(3248));
    layer4_outputs(4110) <= (layer3_outputs(4900)) xor (layer3_outputs(3097));
    layer4_outputs(4111) <= not(layer3_outputs(2891)) or (layer3_outputs(4675));
    layer4_outputs(4112) <= not(layer3_outputs(943));
    layer4_outputs(4113) <= (layer3_outputs(6466)) and (layer3_outputs(2549));
    layer4_outputs(4114) <= '1';
    layer4_outputs(4115) <= '0';
    layer4_outputs(4116) <= not(layer3_outputs(2548));
    layer4_outputs(4117) <= layer3_outputs(3005);
    layer4_outputs(4118) <= (layer3_outputs(2225)) and not (layer3_outputs(1673));
    layer4_outputs(4119) <= '1';
    layer4_outputs(4120) <= not(layer3_outputs(3971));
    layer4_outputs(4121) <= not(layer3_outputs(1425));
    layer4_outputs(4122) <= layer3_outputs(3676);
    layer4_outputs(4123) <= not((layer3_outputs(6722)) xor (layer3_outputs(5151)));
    layer4_outputs(4124) <= '0';
    layer4_outputs(4125) <= not(layer3_outputs(2277));
    layer4_outputs(4126) <= not(layer3_outputs(6883)) or (layer3_outputs(4066));
    layer4_outputs(4127) <= (layer3_outputs(766)) xor (layer3_outputs(6483));
    layer4_outputs(4128) <= not(layer3_outputs(4717));
    layer4_outputs(4129) <= '0';
    layer4_outputs(4130) <= not((layer3_outputs(2257)) or (layer3_outputs(1511)));
    layer4_outputs(4131) <= not(layer3_outputs(1487));
    layer4_outputs(4132) <= (layer3_outputs(6145)) or (layer3_outputs(4007));
    layer4_outputs(4133) <= not(layer3_outputs(4476));
    layer4_outputs(4134) <= not(layer3_outputs(2615));
    layer4_outputs(4135) <= (layer3_outputs(353)) and not (layer3_outputs(5356));
    layer4_outputs(4136) <= layer3_outputs(1371);
    layer4_outputs(4137) <= not(layer3_outputs(5136));
    layer4_outputs(4138) <= not(layer3_outputs(6139));
    layer4_outputs(4139) <= not(layer3_outputs(4567)) or (layer3_outputs(2633));
    layer4_outputs(4140) <= not(layer3_outputs(1347)) or (layer3_outputs(1729));
    layer4_outputs(4141) <= '0';
    layer4_outputs(4142) <= layer3_outputs(3442);
    layer4_outputs(4143) <= (layer3_outputs(2555)) xor (layer3_outputs(114));
    layer4_outputs(4144) <= (layer3_outputs(4223)) and not (layer3_outputs(3411));
    layer4_outputs(4145) <= layer3_outputs(7156);
    layer4_outputs(4146) <= not(layer3_outputs(5072)) or (layer3_outputs(4384));
    layer4_outputs(4147) <= not(layer3_outputs(4693));
    layer4_outputs(4148) <= not(layer3_outputs(3511)) or (layer3_outputs(80));
    layer4_outputs(4149) <= (layer3_outputs(5608)) and (layer3_outputs(3343));
    layer4_outputs(4150) <= layer3_outputs(1979);
    layer4_outputs(4151) <= (layer3_outputs(1338)) and not (layer3_outputs(4236));
    layer4_outputs(4152) <= not(layer3_outputs(6577));
    layer4_outputs(4153) <= not(layer3_outputs(566)) or (layer3_outputs(5042));
    layer4_outputs(4154) <= layer3_outputs(4263);
    layer4_outputs(4155) <= layer3_outputs(2504);
    layer4_outputs(4156) <= layer3_outputs(3215);
    layer4_outputs(4157) <= not(layer3_outputs(7411)) or (layer3_outputs(7576));
    layer4_outputs(4158) <= '1';
    layer4_outputs(4159) <= not(layer3_outputs(1605));
    layer4_outputs(4160) <= not((layer3_outputs(4971)) or (layer3_outputs(4401)));
    layer4_outputs(4161) <= '1';
    layer4_outputs(4162) <= '0';
    layer4_outputs(4163) <= not(layer3_outputs(1138));
    layer4_outputs(4164) <= (layer3_outputs(790)) or (layer3_outputs(762));
    layer4_outputs(4165) <= (layer3_outputs(6308)) and not (layer3_outputs(723));
    layer4_outputs(4166) <= (layer3_outputs(2315)) and (layer3_outputs(1535));
    layer4_outputs(4167) <= layer3_outputs(6256);
    layer4_outputs(4168) <= not(layer3_outputs(2372));
    layer4_outputs(4169) <= layer3_outputs(6687);
    layer4_outputs(4170) <= (layer3_outputs(1428)) and not (layer3_outputs(1097));
    layer4_outputs(4171) <= (layer3_outputs(1668)) and (layer3_outputs(3480));
    layer4_outputs(4172) <= (layer3_outputs(236)) and not (layer3_outputs(2002));
    layer4_outputs(4173) <= not(layer3_outputs(6004)) or (layer3_outputs(7577));
    layer4_outputs(4174) <= '0';
    layer4_outputs(4175) <= layer3_outputs(6695);
    layer4_outputs(4176) <= (layer3_outputs(6718)) and (layer3_outputs(4011));
    layer4_outputs(4177) <= not(layer3_outputs(381)) or (layer3_outputs(6940));
    layer4_outputs(4178) <= (layer3_outputs(2720)) and not (layer3_outputs(5830));
    layer4_outputs(4179) <= not((layer3_outputs(2953)) and (layer3_outputs(3991)));
    layer4_outputs(4180) <= not((layer3_outputs(681)) or (layer3_outputs(4246)));
    layer4_outputs(4181) <= (layer3_outputs(6384)) and not (layer3_outputs(4607));
    layer4_outputs(4182) <= (layer3_outputs(1083)) and (layer3_outputs(2772));
    layer4_outputs(4183) <= not((layer3_outputs(4150)) and (layer3_outputs(3683)));
    layer4_outputs(4184) <= layer3_outputs(5543);
    layer4_outputs(4185) <= layer3_outputs(7391);
    layer4_outputs(4186) <= (layer3_outputs(593)) or (layer3_outputs(6953));
    layer4_outputs(4187) <= not(layer3_outputs(992)) or (layer3_outputs(6168));
    layer4_outputs(4188) <= layer3_outputs(6742);
    layer4_outputs(4189) <= (layer3_outputs(5800)) xor (layer3_outputs(3435));
    layer4_outputs(4190) <= (layer3_outputs(3386)) and not (layer3_outputs(7555));
    layer4_outputs(4191) <= not((layer3_outputs(6985)) and (layer3_outputs(6961)));
    layer4_outputs(4192) <= (layer3_outputs(6646)) or (layer3_outputs(3276));
    layer4_outputs(4193) <= (layer3_outputs(1785)) and not (layer3_outputs(2596));
    layer4_outputs(4194) <= not(layer3_outputs(5762)) or (layer3_outputs(3022));
    layer4_outputs(4195) <= layer3_outputs(656);
    layer4_outputs(4196) <= not((layer3_outputs(3738)) and (layer3_outputs(1294)));
    layer4_outputs(4197) <= not(layer3_outputs(231));
    layer4_outputs(4198) <= not((layer3_outputs(5)) and (layer3_outputs(5555)));
    layer4_outputs(4199) <= not((layer3_outputs(3673)) xor (layer3_outputs(4003)));
    layer4_outputs(4200) <= not((layer3_outputs(2603)) and (layer3_outputs(1437)));
    layer4_outputs(4201) <= (layer3_outputs(2652)) and not (layer3_outputs(4195));
    layer4_outputs(4202) <= layer3_outputs(2134);
    layer4_outputs(4203) <= not(layer3_outputs(1139));
    layer4_outputs(4204) <= not((layer3_outputs(2595)) and (layer3_outputs(1100)));
    layer4_outputs(4205) <= '1';
    layer4_outputs(4206) <= layer3_outputs(7529);
    layer4_outputs(4207) <= not((layer3_outputs(3762)) and (layer3_outputs(7618)));
    layer4_outputs(4208) <= (layer3_outputs(1906)) and (layer3_outputs(1971));
    layer4_outputs(4209) <= not((layer3_outputs(3280)) and (layer3_outputs(3800)));
    layer4_outputs(4210) <= '0';
    layer4_outputs(4211) <= layer3_outputs(3487);
    layer4_outputs(4212) <= not(layer3_outputs(1441));
    layer4_outputs(4213) <= (layer3_outputs(7110)) and (layer3_outputs(3785));
    layer4_outputs(4214) <= (layer3_outputs(1137)) or (layer3_outputs(5260));
    layer4_outputs(4215) <= not(layer3_outputs(4176));
    layer4_outputs(4216) <= (layer3_outputs(1235)) and not (layer3_outputs(4160));
    layer4_outputs(4217) <= not(layer3_outputs(1693));
    layer4_outputs(4218) <= layer3_outputs(1992);
    layer4_outputs(4219) <= (layer3_outputs(2221)) xor (layer3_outputs(7377));
    layer4_outputs(4220) <= (layer3_outputs(7610)) and not (layer3_outputs(4793));
    layer4_outputs(4221) <= not(layer3_outputs(7360));
    layer4_outputs(4222) <= not(layer3_outputs(989)) or (layer3_outputs(7661));
    layer4_outputs(4223) <= layer3_outputs(6620);
    layer4_outputs(4224) <= not(layer3_outputs(5118));
    layer4_outputs(4225) <= not(layer3_outputs(940));
    layer4_outputs(4226) <= layer3_outputs(926);
    layer4_outputs(4227) <= layer3_outputs(6499);
    layer4_outputs(4228) <= not(layer3_outputs(6691));
    layer4_outputs(4229) <= layer3_outputs(7445);
    layer4_outputs(4230) <= layer3_outputs(4378);
    layer4_outputs(4231) <= not(layer3_outputs(4001));
    layer4_outputs(4232) <= layer3_outputs(6537);
    layer4_outputs(4233) <= not(layer3_outputs(281)) or (layer3_outputs(4774));
    layer4_outputs(4234) <= (layer3_outputs(5269)) and not (layer3_outputs(726));
    layer4_outputs(4235) <= (layer3_outputs(6955)) and (layer3_outputs(1539));
    layer4_outputs(4236) <= not(layer3_outputs(780));
    layer4_outputs(4237) <= (layer3_outputs(4370)) or (layer3_outputs(1703));
    layer4_outputs(4238) <= not(layer3_outputs(2398)) or (layer3_outputs(657));
    layer4_outputs(4239) <= layer3_outputs(2197);
    layer4_outputs(4240) <= not(layer3_outputs(3972));
    layer4_outputs(4241) <= layer3_outputs(1802);
    layer4_outputs(4242) <= not((layer3_outputs(509)) xor (layer3_outputs(5040)));
    layer4_outputs(4243) <= (layer3_outputs(4558)) xor (layer3_outputs(1457));
    layer4_outputs(4244) <= (layer3_outputs(5004)) and not (layer3_outputs(4100));
    layer4_outputs(4245) <= (layer3_outputs(2081)) and (layer3_outputs(4898));
    layer4_outputs(4246) <= not((layer3_outputs(6628)) and (layer3_outputs(5319)));
    layer4_outputs(4247) <= not(layer3_outputs(3724));
    layer4_outputs(4248) <= (layer3_outputs(1111)) and (layer3_outputs(1850));
    layer4_outputs(4249) <= not(layer3_outputs(6639));
    layer4_outputs(4250) <= not(layer3_outputs(2342));
    layer4_outputs(4251) <= (layer3_outputs(2520)) and not (layer3_outputs(310));
    layer4_outputs(4252) <= layer3_outputs(5215);
    layer4_outputs(4253) <= layer3_outputs(5877);
    layer4_outputs(4254) <= (layer3_outputs(2072)) and not (layer3_outputs(7495));
    layer4_outputs(4255) <= layer3_outputs(4320);
    layer4_outputs(4256) <= not(layer3_outputs(3215)) or (layer3_outputs(2066));
    layer4_outputs(4257) <= not(layer3_outputs(4328)) or (layer3_outputs(5939));
    layer4_outputs(4258) <= not(layer3_outputs(5934)) or (layer3_outputs(5843));
    layer4_outputs(4259) <= not(layer3_outputs(6105)) or (layer3_outputs(449));
    layer4_outputs(4260) <= not(layer3_outputs(7495));
    layer4_outputs(4261) <= (layer3_outputs(3379)) and (layer3_outputs(1644));
    layer4_outputs(4262) <= layer3_outputs(1819);
    layer4_outputs(4263) <= (layer3_outputs(7203)) and (layer3_outputs(3792));
    layer4_outputs(4264) <= not(layer3_outputs(2962));
    layer4_outputs(4265) <= layer3_outputs(3531);
    layer4_outputs(4266) <= layer3_outputs(4156);
    layer4_outputs(4267) <= layer3_outputs(3717);
    layer4_outputs(4268) <= not(layer3_outputs(965)) or (layer3_outputs(3990));
    layer4_outputs(4269) <= not(layer3_outputs(7136)) or (layer3_outputs(1916));
    layer4_outputs(4270) <= not(layer3_outputs(1375));
    layer4_outputs(4271) <= not(layer3_outputs(3836)) or (layer3_outputs(6676));
    layer4_outputs(4272) <= not(layer3_outputs(5725));
    layer4_outputs(4273) <= (layer3_outputs(5100)) or (layer3_outputs(2490));
    layer4_outputs(4274) <= not(layer3_outputs(5923));
    layer4_outputs(4275) <= not((layer3_outputs(1561)) xor (layer3_outputs(4826)));
    layer4_outputs(4276) <= (layer3_outputs(3878)) and not (layer3_outputs(1318));
    layer4_outputs(4277) <= (layer3_outputs(1853)) and (layer3_outputs(6416));
    layer4_outputs(4278) <= not(layer3_outputs(641)) or (layer3_outputs(1391));
    layer4_outputs(4279) <= '1';
    layer4_outputs(4280) <= '0';
    layer4_outputs(4281) <= not(layer3_outputs(3868)) or (layer3_outputs(2362));
    layer4_outputs(4282) <= not(layer3_outputs(623));
    layer4_outputs(4283) <= not(layer3_outputs(2245));
    layer4_outputs(4284) <= not(layer3_outputs(6626));
    layer4_outputs(4285) <= layer3_outputs(1199);
    layer4_outputs(4286) <= layer3_outputs(1040);
    layer4_outputs(4287) <= (layer3_outputs(1964)) xor (layer3_outputs(5657));
    layer4_outputs(4288) <= not(layer3_outputs(4232));
    layer4_outputs(4289) <= not(layer3_outputs(738)) or (layer3_outputs(4995));
    layer4_outputs(4290) <= not(layer3_outputs(6685)) or (layer3_outputs(6114));
    layer4_outputs(4291) <= not(layer3_outputs(1055));
    layer4_outputs(4292) <= layer3_outputs(1190);
    layer4_outputs(4293) <= not(layer3_outputs(3631)) or (layer3_outputs(2291));
    layer4_outputs(4294) <= layer3_outputs(4522);
    layer4_outputs(4295) <= not((layer3_outputs(692)) and (layer3_outputs(1763)));
    layer4_outputs(4296) <= layer3_outputs(3463);
    layer4_outputs(4297) <= layer3_outputs(951);
    layer4_outputs(4298) <= not(layer3_outputs(4122)) or (layer3_outputs(7295));
    layer4_outputs(4299) <= (layer3_outputs(1786)) and not (layer3_outputs(4284));
    layer4_outputs(4300) <= layer3_outputs(7390);
    layer4_outputs(4301) <= (layer3_outputs(2789)) and (layer3_outputs(4307));
    layer4_outputs(4302) <= not((layer3_outputs(1135)) xor (layer3_outputs(4026)));
    layer4_outputs(4303) <= not(layer3_outputs(3812));
    layer4_outputs(4304) <= not((layer3_outputs(480)) xor (layer3_outputs(4410)));
    layer4_outputs(4305) <= not(layer3_outputs(812)) or (layer3_outputs(3863));
    layer4_outputs(4306) <= not(layer3_outputs(5934));
    layer4_outputs(4307) <= not(layer3_outputs(1771));
    layer4_outputs(4308) <= layer3_outputs(3037);
    layer4_outputs(4309) <= layer3_outputs(5178);
    layer4_outputs(4310) <= layer3_outputs(951);
    layer4_outputs(4311) <= (layer3_outputs(5890)) and not (layer3_outputs(3475));
    layer4_outputs(4312) <= (layer3_outputs(5599)) and not (layer3_outputs(3079));
    layer4_outputs(4313) <= (layer3_outputs(3055)) or (layer3_outputs(7304));
    layer4_outputs(4314) <= layer3_outputs(5758);
    layer4_outputs(4315) <= layer3_outputs(3007);
    layer4_outputs(4316) <= not(layer3_outputs(1047));
    layer4_outputs(4317) <= layer3_outputs(7425);
    layer4_outputs(4318) <= layer3_outputs(3982);
    layer4_outputs(4319) <= not(layer3_outputs(1681));
    layer4_outputs(4320) <= (layer3_outputs(2652)) xor (layer3_outputs(2412));
    layer4_outputs(4321) <= not(layer3_outputs(421));
    layer4_outputs(4322) <= layer3_outputs(5229);
    layer4_outputs(4323) <= (layer3_outputs(7332)) or (layer3_outputs(2980));
    layer4_outputs(4324) <= not((layer3_outputs(4189)) xor (layer3_outputs(6688)));
    layer4_outputs(4325) <= not((layer3_outputs(512)) and (layer3_outputs(5123)));
    layer4_outputs(4326) <= not((layer3_outputs(1560)) and (layer3_outputs(3661)));
    layer4_outputs(4327) <= not(layer3_outputs(1198)) or (layer3_outputs(7505));
    layer4_outputs(4328) <= (layer3_outputs(6172)) and (layer3_outputs(6762));
    layer4_outputs(4329) <= layer3_outputs(2132);
    layer4_outputs(4330) <= '0';
    layer4_outputs(4331) <= layer3_outputs(2682);
    layer4_outputs(4332) <= not((layer3_outputs(6538)) or (layer3_outputs(7522)));
    layer4_outputs(4333) <= '1';
    layer4_outputs(4334) <= '0';
    layer4_outputs(4335) <= not(layer3_outputs(2376));
    layer4_outputs(4336) <= not((layer3_outputs(4015)) and (layer3_outputs(3329)));
    layer4_outputs(4337) <= (layer3_outputs(5390)) and (layer3_outputs(7625));
    layer4_outputs(4338) <= (layer3_outputs(7251)) and not (layer3_outputs(1769));
    layer4_outputs(4339) <= (layer3_outputs(5220)) and not (layer3_outputs(379));
    layer4_outputs(4340) <= layer3_outputs(3393);
    layer4_outputs(4341) <= '1';
    layer4_outputs(4342) <= not(layer3_outputs(2057));
    layer4_outputs(4343) <= '0';
    layer4_outputs(4344) <= not(layer3_outputs(6063)) or (layer3_outputs(4350));
    layer4_outputs(4345) <= layer3_outputs(3705);
    layer4_outputs(4346) <= (layer3_outputs(1001)) and not (layer3_outputs(1640));
    layer4_outputs(4347) <= layer3_outputs(7353);
    layer4_outputs(4348) <= (layer3_outputs(5373)) and not (layer3_outputs(6778));
    layer4_outputs(4349) <= not(layer3_outputs(2022));
    layer4_outputs(4350) <= '1';
    layer4_outputs(4351) <= not(layer3_outputs(2610));
    layer4_outputs(4352) <= (layer3_outputs(5343)) and not (layer3_outputs(6231));
    layer4_outputs(4353) <= (layer3_outputs(1227)) and not (layer3_outputs(2008));
    layer4_outputs(4354) <= layer3_outputs(6222);
    layer4_outputs(4355) <= '0';
    layer4_outputs(4356) <= layer3_outputs(705);
    layer4_outputs(4357) <= not(layer3_outputs(590));
    layer4_outputs(4358) <= (layer3_outputs(3692)) and not (layer3_outputs(4149));
    layer4_outputs(4359) <= not(layer3_outputs(6318));
    layer4_outputs(4360) <= (layer3_outputs(4283)) xor (layer3_outputs(7409));
    layer4_outputs(4361) <= not(layer3_outputs(7643));
    layer4_outputs(4362) <= not(layer3_outputs(170)) or (layer3_outputs(7511));
    layer4_outputs(4363) <= (layer3_outputs(4579)) and not (layer3_outputs(5152));
    layer4_outputs(4364) <= not(layer3_outputs(4319));
    layer4_outputs(4365) <= not(layer3_outputs(874));
    layer4_outputs(4366) <= '1';
    layer4_outputs(4367) <= not(layer3_outputs(5154));
    layer4_outputs(4368) <= not(layer3_outputs(2251)) or (layer3_outputs(3356));
    layer4_outputs(4369) <= (layer3_outputs(3592)) and (layer3_outputs(4173));
    layer4_outputs(4370) <= not(layer3_outputs(6838)) or (layer3_outputs(4241));
    layer4_outputs(4371) <= not(layer3_outputs(4530));
    layer4_outputs(4372) <= layer3_outputs(1567);
    layer4_outputs(4373) <= (layer3_outputs(759)) and not (layer3_outputs(829));
    layer4_outputs(4374) <= (layer3_outputs(6384)) and (layer3_outputs(5917));
    layer4_outputs(4375) <= not((layer3_outputs(6731)) or (layer3_outputs(3528)));
    layer4_outputs(4376) <= not(layer3_outputs(3607));
    layer4_outputs(4377) <= not(layer3_outputs(898));
    layer4_outputs(4378) <= not((layer3_outputs(2202)) xor (layer3_outputs(5521)));
    layer4_outputs(4379) <= layer3_outputs(4531);
    layer4_outputs(4380) <= (layer3_outputs(2676)) and not (layer3_outputs(3321));
    layer4_outputs(4381) <= layer3_outputs(2338);
    layer4_outputs(4382) <= '1';
    layer4_outputs(4383) <= not(layer3_outputs(666)) or (layer3_outputs(4568));
    layer4_outputs(4384) <= (layer3_outputs(7496)) or (layer3_outputs(1027));
    layer4_outputs(4385) <= layer3_outputs(5307);
    layer4_outputs(4386) <= (layer3_outputs(4685)) and (layer3_outputs(6177));
    layer4_outputs(4387) <= (layer3_outputs(5746)) and not (layer3_outputs(6361));
    layer4_outputs(4388) <= (layer3_outputs(7327)) or (layer3_outputs(523));
    layer4_outputs(4389) <= layer3_outputs(4770);
    layer4_outputs(4390) <= '1';
    layer4_outputs(4391) <= layer3_outputs(2479);
    layer4_outputs(4392) <= not((layer3_outputs(6096)) or (layer3_outputs(2408)));
    layer4_outputs(4393) <= (layer3_outputs(535)) and not (layer3_outputs(4111));
    layer4_outputs(4394) <= (layer3_outputs(6344)) and not (layer3_outputs(6656));
    layer4_outputs(4395) <= (layer3_outputs(5248)) and not (layer3_outputs(2200));
    layer4_outputs(4396) <= (layer3_outputs(2873)) or (layer3_outputs(28));
    layer4_outputs(4397) <= not((layer3_outputs(7174)) or (layer3_outputs(7130)));
    layer4_outputs(4398) <= not(layer3_outputs(626));
    layer4_outputs(4399) <= not((layer3_outputs(4941)) xor (layer3_outputs(180)));
    layer4_outputs(4400) <= not(layer3_outputs(174));
    layer4_outputs(4401) <= (layer3_outputs(5239)) xor (layer3_outputs(5670));
    layer4_outputs(4402) <= layer3_outputs(2153);
    layer4_outputs(4403) <= (layer3_outputs(6878)) and not (layer3_outputs(1988));
    layer4_outputs(4404) <= not(layer3_outputs(4395));
    layer4_outputs(4405) <= not((layer3_outputs(1869)) xor (layer3_outputs(4070)));
    layer4_outputs(4406) <= '0';
    layer4_outputs(4407) <= (layer3_outputs(1334)) or (layer3_outputs(1851));
    layer4_outputs(4408) <= layer3_outputs(7324);
    layer4_outputs(4409) <= not(layer3_outputs(1116));
    layer4_outputs(4410) <= not(layer3_outputs(3192)) or (layer3_outputs(5901));
    layer4_outputs(4411) <= not(layer3_outputs(7037));
    layer4_outputs(4412) <= layer3_outputs(3277);
    layer4_outputs(4413) <= not(layer3_outputs(5206));
    layer4_outputs(4414) <= (layer3_outputs(935)) or (layer3_outputs(4294));
    layer4_outputs(4415) <= not(layer3_outputs(671));
    layer4_outputs(4416) <= layer3_outputs(5338);
    layer4_outputs(4417) <= (layer3_outputs(3445)) and (layer3_outputs(1204));
    layer4_outputs(4418) <= not(layer3_outputs(4006));
    layer4_outputs(4419) <= not(layer3_outputs(1817));
    layer4_outputs(4420) <= not(layer3_outputs(1215));
    layer4_outputs(4421) <= not((layer3_outputs(2396)) xor (layer3_outputs(5136)));
    layer4_outputs(4422) <= not(layer3_outputs(6129));
    layer4_outputs(4423) <= layer3_outputs(3715);
    layer4_outputs(4424) <= (layer3_outputs(5433)) or (layer3_outputs(4365));
    layer4_outputs(4425) <= not((layer3_outputs(2808)) or (layer3_outputs(986)));
    layer4_outputs(4426) <= (layer3_outputs(6995)) and not (layer3_outputs(359));
    layer4_outputs(4427) <= layer3_outputs(2034);
    layer4_outputs(4428) <= not(layer3_outputs(6811)) or (layer3_outputs(6913));
    layer4_outputs(4429) <= (layer3_outputs(2811)) and not (layer3_outputs(2643));
    layer4_outputs(4430) <= (layer3_outputs(2489)) and not (layer3_outputs(4227));
    layer4_outputs(4431) <= (layer3_outputs(5116)) or (layer3_outputs(1654));
    layer4_outputs(4432) <= (layer3_outputs(681)) and not (layer3_outputs(7064));
    layer4_outputs(4433) <= not(layer3_outputs(3482));
    layer4_outputs(4434) <= layer3_outputs(2616);
    layer4_outputs(4435) <= (layer3_outputs(378)) and not (layer3_outputs(94));
    layer4_outputs(4436) <= layer3_outputs(4913);
    layer4_outputs(4437) <= layer3_outputs(3062);
    layer4_outputs(4438) <= '0';
    layer4_outputs(4439) <= not((layer3_outputs(5791)) and (layer3_outputs(6726)));
    layer4_outputs(4440) <= (layer3_outputs(3801)) xor (layer3_outputs(3204));
    layer4_outputs(4441) <= (layer3_outputs(2439)) and not (layer3_outputs(4179));
    layer4_outputs(4442) <= (layer3_outputs(1707)) or (layer3_outputs(1557));
    layer4_outputs(4443) <= layer3_outputs(3357);
    layer4_outputs(4444) <= not(layer3_outputs(5320));
    layer4_outputs(4445) <= not(layer3_outputs(6041));
    layer4_outputs(4446) <= not(layer3_outputs(769));
    layer4_outputs(4447) <= not(layer3_outputs(5303));
    layer4_outputs(4448) <= not((layer3_outputs(5105)) or (layer3_outputs(464)));
    layer4_outputs(4449) <= not(layer3_outputs(2809));
    layer4_outputs(4450) <= layer3_outputs(1383);
    layer4_outputs(4451) <= (layer3_outputs(138)) xor (layer3_outputs(78));
    layer4_outputs(4452) <= (layer3_outputs(2711)) and not (layer3_outputs(7019));
    layer4_outputs(4453) <= not(layer3_outputs(3772)) or (layer3_outputs(5530));
    layer4_outputs(4454) <= (layer3_outputs(5783)) and not (layer3_outputs(2238));
    layer4_outputs(4455) <= layer3_outputs(2580);
    layer4_outputs(4456) <= (layer3_outputs(3623)) or (layer3_outputs(6834));
    layer4_outputs(4457) <= not(layer3_outputs(5335));
    layer4_outputs(4458) <= layer3_outputs(4013);
    layer4_outputs(4459) <= not((layer3_outputs(4098)) and (layer3_outputs(6599)));
    layer4_outputs(4460) <= layer3_outputs(3250);
    layer4_outputs(4461) <= layer3_outputs(323);
    layer4_outputs(4462) <= '0';
    layer4_outputs(4463) <= (layer3_outputs(6255)) and not (layer3_outputs(6692));
    layer4_outputs(4464) <= not(layer3_outputs(4217));
    layer4_outputs(4465) <= '0';
    layer4_outputs(4466) <= not(layer3_outputs(6535));
    layer4_outputs(4467) <= '0';
    layer4_outputs(4468) <= (layer3_outputs(6905)) and (layer3_outputs(902));
    layer4_outputs(4469) <= layer3_outputs(100);
    layer4_outputs(4470) <= not(layer3_outputs(772)) or (layer3_outputs(4882));
    layer4_outputs(4471) <= not(layer3_outputs(2205));
    layer4_outputs(4472) <= not(layer3_outputs(4085));
    layer4_outputs(4473) <= not(layer3_outputs(6884));
    layer4_outputs(4474) <= not(layer3_outputs(5894));
    layer4_outputs(4475) <= not((layer3_outputs(171)) and (layer3_outputs(5916)));
    layer4_outputs(4476) <= not((layer3_outputs(5766)) or (layer3_outputs(2038)));
    layer4_outputs(4477) <= not(layer3_outputs(1043));
    layer4_outputs(4478) <= not(layer3_outputs(2397));
    layer4_outputs(4479) <= '1';
    layer4_outputs(4480) <= not(layer3_outputs(2587));
    layer4_outputs(4481) <= (layer3_outputs(4119)) or (layer3_outputs(5793));
    layer4_outputs(4482) <= not((layer3_outputs(5541)) xor (layer3_outputs(879)));
    layer4_outputs(4483) <= layer3_outputs(3633);
    layer4_outputs(4484) <= not(layer3_outputs(3474)) or (layer3_outputs(2433));
    layer4_outputs(4485) <= not((layer3_outputs(5870)) xor (layer3_outputs(1743)));
    layer4_outputs(4486) <= not(layer3_outputs(1993)) or (layer3_outputs(3123));
    layer4_outputs(4487) <= (layer3_outputs(4267)) and not (layer3_outputs(6192));
    layer4_outputs(4488) <= not(layer3_outputs(2210));
    layer4_outputs(4489) <= '1';
    layer4_outputs(4490) <= not((layer3_outputs(5697)) and (layer3_outputs(7393)));
    layer4_outputs(4491) <= (layer3_outputs(7497)) and not (layer3_outputs(5294));
    layer4_outputs(4492) <= (layer3_outputs(6164)) and not (layer3_outputs(6877));
    layer4_outputs(4493) <= layer3_outputs(5579);
    layer4_outputs(4494) <= not(layer3_outputs(5299)) or (layer3_outputs(6095));
    layer4_outputs(4495) <= '0';
    layer4_outputs(4496) <= not((layer3_outputs(3852)) or (layer3_outputs(7390)));
    layer4_outputs(4497) <= layer3_outputs(2443);
    layer4_outputs(4498) <= layer3_outputs(6480);
    layer4_outputs(4499) <= '0';
    layer4_outputs(4500) <= not((layer3_outputs(4686)) and (layer3_outputs(5797)));
    layer4_outputs(4501) <= not(layer3_outputs(3672));
    layer4_outputs(4502) <= not(layer3_outputs(2282)) or (layer3_outputs(4911));
    layer4_outputs(4503) <= not(layer3_outputs(711));
    layer4_outputs(4504) <= layer3_outputs(722);
    layer4_outputs(4505) <= layer3_outputs(6745);
    layer4_outputs(4506) <= not(layer3_outputs(3581)) or (layer3_outputs(2195));
    layer4_outputs(4507) <= layer3_outputs(6735);
    layer4_outputs(4508) <= layer3_outputs(5731);
    layer4_outputs(4509) <= (layer3_outputs(5476)) xor (layer3_outputs(3387));
    layer4_outputs(4510) <= not(layer3_outputs(5000));
    layer4_outputs(4511) <= (layer3_outputs(5659)) or (layer3_outputs(7660));
    layer4_outputs(4512) <= not(layer3_outputs(2233));
    layer4_outputs(4513) <= not((layer3_outputs(6020)) or (layer3_outputs(111)));
    layer4_outputs(4514) <= not((layer3_outputs(5547)) or (layer3_outputs(2166)));
    layer4_outputs(4515) <= not(layer3_outputs(6911));
    layer4_outputs(4516) <= not(layer3_outputs(1584));
    layer4_outputs(4517) <= '1';
    layer4_outputs(4518) <= not((layer3_outputs(4577)) or (layer3_outputs(3908)));
    layer4_outputs(4519) <= (layer3_outputs(6234)) and (layer3_outputs(1219));
    layer4_outputs(4520) <= not((layer3_outputs(952)) or (layer3_outputs(7142)));
    layer4_outputs(4521) <= layer3_outputs(5985);
    layer4_outputs(4522) <= layer3_outputs(7663);
    layer4_outputs(4523) <= layer3_outputs(155);
    layer4_outputs(4524) <= (layer3_outputs(5846)) and not (layer3_outputs(5901));
    layer4_outputs(4525) <= not((layer3_outputs(3165)) or (layer3_outputs(1793)));
    layer4_outputs(4526) <= (layer3_outputs(4847)) or (layer3_outputs(961));
    layer4_outputs(4527) <= not(layer3_outputs(99));
    layer4_outputs(4528) <= layer3_outputs(2884);
    layer4_outputs(4529) <= not(layer3_outputs(1686));
    layer4_outputs(4530) <= not(layer3_outputs(4217));
    layer4_outputs(4531) <= not(layer3_outputs(6363));
    layer4_outputs(4532) <= '0';
    layer4_outputs(4533) <= (layer3_outputs(4805)) and (layer3_outputs(5835));
    layer4_outputs(4534) <= not(layer3_outputs(5054));
    layer4_outputs(4535) <= (layer3_outputs(7543)) and (layer3_outputs(4748));
    layer4_outputs(4536) <= not(layer3_outputs(2942));
    layer4_outputs(4537) <= not(layer3_outputs(5302));
    layer4_outputs(4538) <= not((layer3_outputs(2910)) and (layer3_outputs(6659)));
    layer4_outputs(4539) <= not(layer3_outputs(833));
    layer4_outputs(4540) <= not(layer3_outputs(5279));
    layer4_outputs(4541) <= layer3_outputs(3774);
    layer4_outputs(4542) <= layer3_outputs(3550);
    layer4_outputs(4543) <= not(layer3_outputs(6539));
    layer4_outputs(4544) <= layer3_outputs(1513);
    layer4_outputs(4545) <= (layer3_outputs(2232)) and (layer3_outputs(4562));
    layer4_outputs(4546) <= (layer3_outputs(3142)) xor (layer3_outputs(6564));
    layer4_outputs(4547) <= not((layer3_outputs(7476)) and (layer3_outputs(6849)));
    layer4_outputs(4548) <= not(layer3_outputs(3127)) or (layer3_outputs(2677));
    layer4_outputs(4549) <= not(layer3_outputs(2118));
    layer4_outputs(4550) <= (layer3_outputs(3566)) and not (layer3_outputs(569));
    layer4_outputs(4551) <= not((layer3_outputs(0)) and (layer3_outputs(6463)));
    layer4_outputs(4552) <= layer3_outputs(1797);
    layer4_outputs(4553) <= not(layer3_outputs(269));
    layer4_outputs(4554) <= not(layer3_outputs(4968)) or (layer3_outputs(1295));
    layer4_outputs(4555) <= (layer3_outputs(2813)) or (layer3_outputs(2477));
    layer4_outputs(4556) <= '0';
    layer4_outputs(4557) <= layer3_outputs(4901);
    layer4_outputs(4558) <= (layer3_outputs(2348)) or (layer3_outputs(5243));
    layer4_outputs(4559) <= not(layer3_outputs(6913));
    layer4_outputs(4560) <= (layer3_outputs(7482)) or (layer3_outputs(3679));
    layer4_outputs(4561) <= (layer3_outputs(7340)) and not (layer3_outputs(4505));
    layer4_outputs(4562) <= not(layer3_outputs(2770));
    layer4_outputs(4563) <= (layer3_outputs(1939)) and not (layer3_outputs(5780));
    layer4_outputs(4564) <= not(layer3_outputs(4447));
    layer4_outputs(4565) <= (layer3_outputs(1185)) xor (layer3_outputs(7248));
    layer4_outputs(4566) <= '0';
    layer4_outputs(4567) <= layer3_outputs(691);
    layer4_outputs(4568) <= not(layer3_outputs(1972)) or (layer3_outputs(5125));
    layer4_outputs(4569) <= (layer3_outputs(943)) and not (layer3_outputs(2364));
    layer4_outputs(4570) <= layer3_outputs(6326);
    layer4_outputs(4571) <= (layer3_outputs(4087)) and (layer3_outputs(4758));
    layer4_outputs(4572) <= not((layer3_outputs(220)) xor (layer3_outputs(5087)));
    layer4_outputs(4573) <= (layer3_outputs(7579)) and not (layer3_outputs(3874));
    layer4_outputs(4574) <= not(layer3_outputs(4137));
    layer4_outputs(4575) <= '1';
    layer4_outputs(4576) <= (layer3_outputs(6755)) xor (layer3_outputs(938));
    layer4_outputs(4577) <= layer3_outputs(3127);
    layer4_outputs(4578) <= (layer3_outputs(6848)) and not (layer3_outputs(2159));
    layer4_outputs(4579) <= not((layer3_outputs(2095)) xor (layer3_outputs(6753)));
    layer4_outputs(4580) <= not(layer3_outputs(849));
    layer4_outputs(4581) <= (layer3_outputs(5474)) xor (layer3_outputs(7624));
    layer4_outputs(4582) <= not(layer3_outputs(2080));
    layer4_outputs(4583) <= not((layer3_outputs(4268)) or (layer3_outputs(6090)));
    layer4_outputs(4584) <= not((layer3_outputs(7468)) or (layer3_outputs(2939)));
    layer4_outputs(4585) <= layer3_outputs(426);
    layer4_outputs(4586) <= (layer3_outputs(3965)) xor (layer3_outputs(3138));
    layer4_outputs(4587) <= layer3_outputs(4842);
    layer4_outputs(4588) <= layer3_outputs(1264);
    layer4_outputs(4589) <= (layer3_outputs(2647)) and not (layer3_outputs(4595));
    layer4_outputs(4590) <= (layer3_outputs(2795)) or (layer3_outputs(2468));
    layer4_outputs(4591) <= (layer3_outputs(1065)) and (layer3_outputs(1402));
    layer4_outputs(4592) <= layer3_outputs(5526);
    layer4_outputs(4593) <= not(layer3_outputs(3912));
    layer4_outputs(4594) <= layer3_outputs(3512);
    layer4_outputs(4595) <= not(layer3_outputs(1381));
    layer4_outputs(4596) <= not(layer3_outputs(415));
    layer4_outputs(4597) <= not((layer3_outputs(1499)) and (layer3_outputs(3991)));
    layer4_outputs(4598) <= layer3_outputs(6838);
    layer4_outputs(4599) <= (layer3_outputs(4278)) and (layer3_outputs(596));
    layer4_outputs(4600) <= not(layer3_outputs(3933));
    layer4_outputs(4601) <= '1';
    layer4_outputs(4602) <= (layer3_outputs(6772)) and not (layer3_outputs(6180));
    layer4_outputs(4603) <= layer3_outputs(2547);
    layer4_outputs(4604) <= layer3_outputs(4773);
    layer4_outputs(4605) <= '1';
    layer4_outputs(4606) <= not(layer3_outputs(2732));
    layer4_outputs(4607) <= layer3_outputs(3697);
    layer4_outputs(4608) <= not(layer3_outputs(6351)) or (layer3_outputs(732));
    layer4_outputs(4609) <= not(layer3_outputs(4290)) or (layer3_outputs(3889));
    layer4_outputs(4610) <= '1';
    layer4_outputs(4611) <= not(layer3_outputs(6800));
    layer4_outputs(4612) <= layer3_outputs(3989);
    layer4_outputs(4613) <= not(layer3_outputs(5019)) or (layer3_outputs(7126));
    layer4_outputs(4614) <= layer3_outputs(1272);
    layer4_outputs(4615) <= not(layer3_outputs(475)) or (layer3_outputs(1440));
    layer4_outputs(4616) <= (layer3_outputs(5533)) xor (layer3_outputs(6211));
    layer4_outputs(4617) <= (layer3_outputs(3121)) or (layer3_outputs(7237));
    layer4_outputs(4618) <= not((layer3_outputs(4861)) or (layer3_outputs(2359)));
    layer4_outputs(4619) <= layer3_outputs(375);
    layer4_outputs(4620) <= layer3_outputs(3997);
    layer4_outputs(4621) <= not(layer3_outputs(5576));
    layer4_outputs(4622) <= (layer3_outputs(7125)) and not (layer3_outputs(2368));
    layer4_outputs(4623) <= not(layer3_outputs(1829));
    layer4_outputs(4624) <= (layer3_outputs(2168)) or (layer3_outputs(6233));
    layer4_outputs(4625) <= layer3_outputs(7446);
    layer4_outputs(4626) <= (layer3_outputs(2529)) or (layer3_outputs(4483));
    layer4_outputs(4627) <= layer3_outputs(6921);
    layer4_outputs(4628) <= not(layer3_outputs(5807));
    layer4_outputs(4629) <= layer3_outputs(4598);
    layer4_outputs(4630) <= not((layer3_outputs(2521)) xor (layer3_outputs(2281)));
    layer4_outputs(4631) <= not((layer3_outputs(1146)) and (layer3_outputs(6711)));
    layer4_outputs(4632) <= layer3_outputs(2148);
    layer4_outputs(4633) <= not((layer3_outputs(2971)) and (layer3_outputs(155)));
    layer4_outputs(4634) <= not(layer3_outputs(2502));
    layer4_outputs(4635) <= layer3_outputs(1037);
    layer4_outputs(4636) <= (layer3_outputs(4182)) and not (layer3_outputs(474));
    layer4_outputs(4637) <= not(layer3_outputs(826));
    layer4_outputs(4638) <= not(layer3_outputs(1208)) or (layer3_outputs(1730));
    layer4_outputs(4639) <= layer3_outputs(5164);
    layer4_outputs(4640) <= (layer3_outputs(5891)) and not (layer3_outputs(1314));
    layer4_outputs(4641) <= not(layer3_outputs(214)) or (layer3_outputs(2588));
    layer4_outputs(4642) <= layer3_outputs(3854);
    layer4_outputs(4643) <= '0';
    layer4_outputs(4644) <= (layer3_outputs(252)) xor (layer3_outputs(2841));
    layer4_outputs(4645) <= (layer3_outputs(7188)) and not (layer3_outputs(141));
    layer4_outputs(4646) <= (layer3_outputs(7032)) and not (layer3_outputs(2904));
    layer4_outputs(4647) <= not(layer3_outputs(7413)) or (layer3_outputs(2139));
    layer4_outputs(4648) <= layer3_outputs(578);
    layer4_outputs(4649) <= not(layer3_outputs(2255));
    layer4_outputs(4650) <= '0';
    layer4_outputs(4651) <= not(layer3_outputs(5609));
    layer4_outputs(4652) <= layer3_outputs(2259);
    layer4_outputs(4653) <= not(layer3_outputs(6550));
    layer4_outputs(4654) <= not(layer3_outputs(460)) or (layer3_outputs(1245));
    layer4_outputs(4655) <= (layer3_outputs(5577)) and not (layer3_outputs(4428));
    layer4_outputs(4656) <= layer3_outputs(7294);
    layer4_outputs(4657) <= (layer3_outputs(3439)) or (layer3_outputs(1968));
    layer4_outputs(4658) <= not(layer3_outputs(4039)) or (layer3_outputs(7094));
    layer4_outputs(4659) <= '1';
    layer4_outputs(4660) <= not((layer3_outputs(3444)) and (layer3_outputs(264)));
    layer4_outputs(4661) <= (layer3_outputs(4655)) or (layer3_outputs(2772));
    layer4_outputs(4662) <= not((layer3_outputs(6193)) or (layer3_outputs(23)));
    layer4_outputs(4663) <= layer3_outputs(888);
    layer4_outputs(4664) <= not(layer3_outputs(885)) or (layer3_outputs(1344));
    layer4_outputs(4665) <= layer3_outputs(1237);
    layer4_outputs(4666) <= not(layer3_outputs(5929));
    layer4_outputs(4667) <= layer3_outputs(6436);
    layer4_outputs(4668) <= not(layer3_outputs(616));
    layer4_outputs(4669) <= not(layer3_outputs(4262));
    layer4_outputs(4670) <= not(layer3_outputs(2930));
    layer4_outputs(4671) <= layer3_outputs(3515);
    layer4_outputs(4672) <= not((layer3_outputs(7641)) or (layer3_outputs(4448)));
    layer4_outputs(4673) <= not(layer3_outputs(1366));
    layer4_outputs(4674) <= '0';
    layer4_outputs(4675) <= not((layer3_outputs(3286)) or (layer3_outputs(4190)));
    layer4_outputs(4676) <= '0';
    layer4_outputs(4677) <= not(layer3_outputs(7504));
    layer4_outputs(4678) <= (layer3_outputs(893)) and not (layer3_outputs(4466));
    layer4_outputs(4679) <= not(layer3_outputs(4372));
    layer4_outputs(4680) <= '0';
    layer4_outputs(4681) <= not((layer3_outputs(3968)) and (layer3_outputs(1419)));
    layer4_outputs(4682) <= not(layer3_outputs(1732)) or (layer3_outputs(3768));
    layer4_outputs(4683) <= (layer3_outputs(7274)) and (layer3_outputs(2778));
    layer4_outputs(4684) <= not(layer3_outputs(545));
    layer4_outputs(4685) <= not(layer3_outputs(5908));
    layer4_outputs(4686) <= layer3_outputs(7515);
    layer4_outputs(4687) <= not(layer3_outputs(27));
    layer4_outputs(4688) <= not(layer3_outputs(4922));
    layer4_outputs(4689) <= layer3_outputs(149);
    layer4_outputs(4690) <= layer3_outputs(2280);
    layer4_outputs(4691) <= not(layer3_outputs(7640));
    layer4_outputs(4692) <= '0';
    layer4_outputs(4693) <= layer3_outputs(2276);
    layer4_outputs(4694) <= layer3_outputs(1056);
    layer4_outputs(4695) <= layer3_outputs(2616);
    layer4_outputs(4696) <= '0';
    layer4_outputs(4697) <= not(layer3_outputs(3099)) or (layer3_outputs(282));
    layer4_outputs(4698) <= layer3_outputs(3470);
    layer4_outputs(4699) <= layer3_outputs(2570);
    layer4_outputs(4700) <= '1';
    layer4_outputs(4701) <= not((layer3_outputs(7065)) or (layer3_outputs(4092)));
    layer4_outputs(4702) <= layer3_outputs(6831);
    layer4_outputs(4703) <= layer3_outputs(7574);
    layer4_outputs(4704) <= not((layer3_outputs(1113)) or (layer3_outputs(4169)));
    layer4_outputs(4705) <= (layer3_outputs(5921)) and (layer3_outputs(7345));
    layer4_outputs(4706) <= layer3_outputs(6510);
    layer4_outputs(4707) <= not((layer3_outputs(389)) or (layer3_outputs(4604)));
    layer4_outputs(4708) <= (layer3_outputs(1351)) and (layer3_outputs(2527));
    layer4_outputs(4709) <= not((layer3_outputs(2441)) or (layer3_outputs(5247)));
    layer4_outputs(4710) <= (layer3_outputs(7155)) xor (layer3_outputs(5368));
    layer4_outputs(4711) <= not(layer3_outputs(501)) or (layer3_outputs(7649));
    layer4_outputs(4712) <= (layer3_outputs(3574)) xor (layer3_outputs(5262));
    layer4_outputs(4713) <= not(layer3_outputs(135));
    layer4_outputs(4714) <= (layer3_outputs(4553)) and not (layer3_outputs(1770));
    layer4_outputs(4715) <= (layer3_outputs(3750)) and not (layer3_outputs(369));
    layer4_outputs(4716) <= (layer3_outputs(4629)) and (layer3_outputs(3048));
    layer4_outputs(4717) <= not(layer3_outputs(6282));
    layer4_outputs(4718) <= not(layer3_outputs(2014));
    layer4_outputs(4719) <= '0';
    layer4_outputs(4720) <= '0';
    layer4_outputs(4721) <= not(layer3_outputs(3659)) or (layer3_outputs(3023));
    layer4_outputs(4722) <= layer3_outputs(5892);
    layer4_outputs(4723) <= not((layer3_outputs(6909)) and (layer3_outputs(2337)));
    layer4_outputs(4724) <= (layer3_outputs(4205)) or (layer3_outputs(4552));
    layer4_outputs(4725) <= layer3_outputs(5097);
    layer4_outputs(4726) <= not(layer3_outputs(5733));
    layer4_outputs(4727) <= (layer3_outputs(3864)) and not (layer3_outputs(2813));
    layer4_outputs(4728) <= not(layer3_outputs(7363));
    layer4_outputs(4729) <= not(layer3_outputs(6943));
    layer4_outputs(4730) <= layer3_outputs(1346);
    layer4_outputs(4731) <= not((layer3_outputs(6806)) xor (layer3_outputs(326)));
    layer4_outputs(4732) <= layer3_outputs(1620);
    layer4_outputs(4733) <= (layer3_outputs(5069)) or (layer3_outputs(4617));
    layer4_outputs(4734) <= not(layer3_outputs(172));
    layer4_outputs(4735) <= not(layer3_outputs(3254));
    layer4_outputs(4736) <= not(layer3_outputs(7325));
    layer4_outputs(4737) <= layer3_outputs(3163);
    layer4_outputs(4738) <= layer3_outputs(1248);
    layer4_outputs(4739) <= layer3_outputs(3469);
    layer4_outputs(4740) <= layer3_outputs(6166);
    layer4_outputs(4741) <= layer3_outputs(1985);
    layer4_outputs(4742) <= not(layer3_outputs(5257)) or (layer3_outputs(508));
    layer4_outputs(4743) <= not(layer3_outputs(4427));
    layer4_outputs(4744) <= (layer3_outputs(4478)) or (layer3_outputs(2154));
    layer4_outputs(4745) <= not(layer3_outputs(4125)) or (layer3_outputs(7153));
    layer4_outputs(4746) <= layer3_outputs(5691);
    layer4_outputs(4747) <= (layer3_outputs(40)) and not (layer3_outputs(5047));
    layer4_outputs(4748) <= not(layer3_outputs(6553)) or (layer3_outputs(441));
    layer4_outputs(4749) <= not(layer3_outputs(6195));
    layer4_outputs(4750) <= not((layer3_outputs(6576)) xor (layer3_outputs(1378)));
    layer4_outputs(4751) <= not((layer3_outputs(2275)) and (layer3_outputs(3768)));
    layer4_outputs(4752) <= (layer3_outputs(3940)) and (layer3_outputs(2127));
    layer4_outputs(4753) <= not((layer3_outputs(354)) and (layer3_outputs(2931)));
    layer4_outputs(4754) <= (layer3_outputs(1050)) or (layer3_outputs(607));
    layer4_outputs(4755) <= not((layer3_outputs(2961)) xor (layer3_outputs(4816)));
    layer4_outputs(4756) <= (layer3_outputs(2782)) and not (layer3_outputs(5523));
    layer4_outputs(4757) <= layer3_outputs(5305);
    layer4_outputs(4758) <= layer3_outputs(2823);
    layer4_outputs(4759) <= layer3_outputs(6560);
    layer4_outputs(4760) <= layer3_outputs(2206);
    layer4_outputs(4761) <= (layer3_outputs(251)) and not (layer3_outputs(2755));
    layer4_outputs(4762) <= layer3_outputs(7488);
    layer4_outputs(4763) <= (layer3_outputs(4556)) xor (layer3_outputs(2296));
    layer4_outputs(4764) <= '0';
    layer4_outputs(4765) <= not(layer3_outputs(4798)) or (layer3_outputs(7191));
    layer4_outputs(4766) <= layer3_outputs(7041);
    layer4_outputs(4767) <= layer3_outputs(5029);
    layer4_outputs(4768) <= not(layer3_outputs(5911));
    layer4_outputs(4769) <= not(layer3_outputs(1828)) or (layer3_outputs(4600));
    layer4_outputs(4770) <= layer3_outputs(33);
    layer4_outputs(4771) <= layer3_outputs(73);
    layer4_outputs(4772) <= (layer3_outputs(7233)) xor (layer3_outputs(1492));
    layer4_outputs(4773) <= layer3_outputs(6868);
    layer4_outputs(4774) <= (layer3_outputs(5402)) and (layer3_outputs(4087));
    layer4_outputs(4775) <= '1';
    layer4_outputs(4776) <= not(layer3_outputs(6674)) or (layer3_outputs(1282));
    layer4_outputs(4777) <= '0';
    layer4_outputs(4778) <= not(layer3_outputs(6203)) or (layer3_outputs(3485));
    layer4_outputs(4779) <= not(layer3_outputs(6012));
    layer4_outputs(4780) <= layer3_outputs(1612);
    layer4_outputs(4781) <= layer3_outputs(1421);
    layer4_outputs(4782) <= layer3_outputs(6669);
    layer4_outputs(4783) <= '1';
    layer4_outputs(4784) <= layer3_outputs(6130);
    layer4_outputs(4785) <= not(layer3_outputs(620)) or (layer3_outputs(799));
    layer4_outputs(4786) <= not(layer3_outputs(3513));
    layer4_outputs(4787) <= not((layer3_outputs(980)) xor (layer3_outputs(4332)));
    layer4_outputs(4788) <= (layer3_outputs(7549)) and (layer3_outputs(7215));
    layer4_outputs(4789) <= not(layer3_outputs(4023)) or (layer3_outputs(967));
    layer4_outputs(4790) <= (layer3_outputs(1926)) and not (layer3_outputs(2824));
    layer4_outputs(4791) <= (layer3_outputs(5839)) and not (layer3_outputs(937));
    layer4_outputs(4792) <= not((layer3_outputs(2861)) or (layer3_outputs(7517)));
    layer4_outputs(4793) <= (layer3_outputs(708)) and (layer3_outputs(7415));
    layer4_outputs(4794) <= not(layer3_outputs(6732));
    layer4_outputs(4795) <= not(layer3_outputs(3461));
    layer4_outputs(4796) <= (layer3_outputs(5308)) and not (layer3_outputs(5304));
    layer4_outputs(4797) <= not(layer3_outputs(1785));
    layer4_outputs(4798) <= (layer3_outputs(1567)) and not (layer3_outputs(984));
    layer4_outputs(4799) <= not(layer3_outputs(3745));
    layer4_outputs(4800) <= layer3_outputs(4389);
    layer4_outputs(4801) <= (layer3_outputs(4587)) and not (layer3_outputs(466));
    layer4_outputs(4802) <= not(layer3_outputs(7557)) or (layer3_outputs(531));
    layer4_outputs(4803) <= '0';
    layer4_outputs(4804) <= (layer3_outputs(6890)) and not (layer3_outputs(2074));
    layer4_outputs(4805) <= (layer3_outputs(6697)) xor (layer3_outputs(277));
    layer4_outputs(4806) <= (layer3_outputs(7093)) or (layer3_outputs(1326));
    layer4_outputs(4807) <= layer3_outputs(1945);
    layer4_outputs(4808) <= not((layer3_outputs(1103)) and (layer3_outputs(597)));
    layer4_outputs(4809) <= (layer3_outputs(4998)) and (layer3_outputs(7394));
    layer4_outputs(4810) <= (layer3_outputs(5487)) and not (layer3_outputs(4441));
    layer4_outputs(4811) <= not(layer3_outputs(1212));
    layer4_outputs(4812) <= (layer3_outputs(3586)) and not (layer3_outputs(5696));
    layer4_outputs(4813) <= (layer3_outputs(4875)) or (layer3_outputs(2401));
    layer4_outputs(4814) <= (layer3_outputs(4884)) and not (layer3_outputs(27));
    layer4_outputs(4815) <= layer3_outputs(5098);
    layer4_outputs(4816) <= layer3_outputs(5919);
    layer4_outputs(4817) <= (layer3_outputs(7230)) and not (layer3_outputs(7105));
    layer4_outputs(4818) <= (layer3_outputs(2816)) or (layer3_outputs(4088));
    layer4_outputs(4819) <= layer3_outputs(2869);
    layer4_outputs(4820) <= not((layer3_outputs(2008)) and (layer3_outputs(5193)));
    layer4_outputs(4821) <= not(layer3_outputs(1261));
    layer4_outputs(4822) <= layer3_outputs(1835);
    layer4_outputs(4823) <= layer3_outputs(241);
    layer4_outputs(4824) <= not(layer3_outputs(5856)) or (layer3_outputs(6835));
    layer4_outputs(4825) <= (layer3_outputs(6094)) and (layer3_outputs(2069));
    layer4_outputs(4826) <= (layer3_outputs(2592)) xor (layer3_outputs(3997));
    layer4_outputs(4827) <= layer3_outputs(734);
    layer4_outputs(4828) <= (layer3_outputs(1626)) and not (layer3_outputs(231));
    layer4_outputs(4829) <= (layer3_outputs(5907)) and not (layer3_outputs(1635));
    layer4_outputs(4830) <= (layer3_outputs(2806)) xor (layer3_outputs(6238));
    layer4_outputs(4831) <= layer3_outputs(1339);
    layer4_outputs(4832) <= layer3_outputs(7656);
    layer4_outputs(4833) <= not(layer3_outputs(7644)) or (layer3_outputs(3601));
    layer4_outputs(4834) <= not(layer3_outputs(3120));
    layer4_outputs(4835) <= layer3_outputs(6277);
    layer4_outputs(4836) <= layer3_outputs(452);
    layer4_outputs(4837) <= '1';
    layer4_outputs(4838) <= layer3_outputs(6321);
    layer4_outputs(4839) <= not((layer3_outputs(2500)) and (layer3_outputs(5952)));
    layer4_outputs(4840) <= not((layer3_outputs(7501)) xor (layer3_outputs(3762)));
    layer4_outputs(4841) <= (layer3_outputs(924)) and (layer3_outputs(4572));
    layer4_outputs(4842) <= (layer3_outputs(7024)) xor (layer3_outputs(1795));
    layer4_outputs(4843) <= not((layer3_outputs(4276)) or (layer3_outputs(4193)));
    layer4_outputs(4844) <= not(layer3_outputs(2187));
    layer4_outputs(4845) <= layer3_outputs(5737);
    layer4_outputs(4846) <= not((layer3_outputs(1711)) and (layer3_outputs(7318)));
    layer4_outputs(4847) <= (layer3_outputs(3838)) and (layer3_outputs(675));
    layer4_outputs(4848) <= layer3_outputs(4973);
    layer4_outputs(4849) <= (layer3_outputs(2118)) and not (layer3_outputs(4322));
    layer4_outputs(4850) <= layer3_outputs(3354);
    layer4_outputs(4851) <= (layer3_outputs(7009)) xor (layer3_outputs(7233));
    layer4_outputs(4852) <= (layer3_outputs(7038)) or (layer3_outputs(5834));
    layer4_outputs(4853) <= not(layer3_outputs(2612));
    layer4_outputs(4854) <= (layer3_outputs(3628)) xor (layer3_outputs(6296));
    layer4_outputs(4855) <= not(layer3_outputs(2024));
    layer4_outputs(4856) <= not(layer3_outputs(6376));
    layer4_outputs(4857) <= not(layer3_outputs(3999)) or (layer3_outputs(5687));
    layer4_outputs(4858) <= (layer3_outputs(3959)) and not (layer3_outputs(6782));
    layer4_outputs(4859) <= '1';
    layer4_outputs(4860) <= not(layer3_outputs(1973));
    layer4_outputs(4861) <= (layer3_outputs(6713)) xor (layer3_outputs(6805));
    layer4_outputs(4862) <= not(layer3_outputs(4580));
    layer4_outputs(4863) <= layer3_outputs(3578);
    layer4_outputs(4864) <= not(layer3_outputs(2906)) or (layer3_outputs(3926));
    layer4_outputs(4865) <= '0';
    layer4_outputs(4866) <= not((layer3_outputs(7148)) xor (layer3_outputs(6807)));
    layer4_outputs(4867) <= (layer3_outputs(6896)) and not (layer3_outputs(1478));
    layer4_outputs(4868) <= layer3_outputs(4396);
    layer4_outputs(4869) <= (layer3_outputs(3761)) and not (layer3_outputs(3018));
    layer4_outputs(4870) <= (layer3_outputs(940)) and not (layer3_outputs(4563));
    layer4_outputs(4871) <= not((layer3_outputs(1967)) or (layer3_outputs(6325)));
    layer4_outputs(4872) <= not(layer3_outputs(4826));
    layer4_outputs(4873) <= '1';
    layer4_outputs(4874) <= (layer3_outputs(4561)) and not (layer3_outputs(509));
    layer4_outputs(4875) <= layer3_outputs(5558);
    layer4_outputs(4876) <= (layer3_outputs(5127)) and not (layer3_outputs(2882));
    layer4_outputs(4877) <= not(layer3_outputs(3827));
    layer4_outputs(4878) <= (layer3_outputs(718)) and (layer3_outputs(7061));
    layer4_outputs(4879) <= not(layer3_outputs(5540));
    layer4_outputs(4880) <= not(layer3_outputs(5617)) or (layer3_outputs(1337));
    layer4_outputs(4881) <= not(layer3_outputs(2957));
    layer4_outputs(4882) <= '0';
    layer4_outputs(4883) <= layer3_outputs(5261);
    layer4_outputs(4884) <= (layer3_outputs(42)) and (layer3_outputs(5923));
    layer4_outputs(4885) <= not((layer3_outputs(4420)) xor (layer3_outputs(7118)));
    layer4_outputs(4886) <= layer3_outputs(4237);
    layer4_outputs(4887) <= not(layer3_outputs(6010)) or (layer3_outputs(7030));
    layer4_outputs(4888) <= layer3_outputs(1617);
    layer4_outputs(4889) <= not(layer3_outputs(6837));
    layer4_outputs(4890) <= not(layer3_outputs(1337));
    layer4_outputs(4891) <= (layer3_outputs(7331)) and not (layer3_outputs(3078));
    layer4_outputs(4892) <= (layer3_outputs(6787)) and (layer3_outputs(239));
    layer4_outputs(4893) <= layer3_outputs(7605);
    layer4_outputs(4894) <= not(layer3_outputs(1626));
    layer4_outputs(4895) <= (layer3_outputs(4929)) and not (layer3_outputs(4628));
    layer4_outputs(4896) <= not((layer3_outputs(4815)) or (layer3_outputs(4100)));
    layer4_outputs(4897) <= (layer3_outputs(988)) or (layer3_outputs(3680));
    layer4_outputs(4898) <= not((layer3_outputs(4642)) xor (layer3_outputs(439)));
    layer4_outputs(4899) <= layer3_outputs(4204);
    layer4_outputs(4900) <= (layer3_outputs(2615)) and (layer3_outputs(5432));
    layer4_outputs(4901) <= layer3_outputs(60);
    layer4_outputs(4902) <= layer3_outputs(5876);
    layer4_outputs(4903) <= (layer3_outputs(3794)) and not (layer3_outputs(2650));
    layer4_outputs(4904) <= layer3_outputs(5057);
    layer4_outputs(4905) <= layer3_outputs(5390);
    layer4_outputs(4906) <= (layer3_outputs(2602)) and (layer3_outputs(7218));
    layer4_outputs(4907) <= not(layer3_outputs(4293));
    layer4_outputs(4908) <= not(layer3_outputs(3431));
    layer4_outputs(4909) <= (layer3_outputs(6872)) xor (layer3_outputs(2231));
    layer4_outputs(4910) <= not(layer3_outputs(3176));
    layer4_outputs(4911) <= not(layer3_outputs(911));
    layer4_outputs(4912) <= not(layer3_outputs(1310));
    layer4_outputs(4913) <= not(layer3_outputs(2174));
    layer4_outputs(4914) <= not(layer3_outputs(7224)) or (layer3_outputs(4861));
    layer4_outputs(4915) <= (layer3_outputs(6678)) and not (layer3_outputs(552));
    layer4_outputs(4916) <= '1';
    layer4_outputs(4917) <= not(layer3_outputs(6228));
    layer4_outputs(4918) <= layer3_outputs(4208);
    layer4_outputs(4919) <= layer3_outputs(7042);
    layer4_outputs(4920) <= not(layer3_outputs(5936));
    layer4_outputs(4921) <= not(layer3_outputs(7435)) or (layer3_outputs(6881));
    layer4_outputs(4922) <= (layer3_outputs(2638)) or (layer3_outputs(1596));
    layer4_outputs(4923) <= not(layer3_outputs(5918));
    layer4_outputs(4924) <= not(layer3_outputs(5070));
    layer4_outputs(4925) <= (layer3_outputs(470)) xor (layer3_outputs(5047));
    layer4_outputs(4926) <= (layer3_outputs(2852)) and not (layer3_outputs(1137));
    layer4_outputs(4927) <= (layer3_outputs(4283)) and (layer3_outputs(3115));
    layer4_outputs(4928) <= not(layer3_outputs(819));
    layer4_outputs(4929) <= (layer3_outputs(915)) and not (layer3_outputs(5326));
    layer4_outputs(4930) <= not((layer3_outputs(7078)) or (layer3_outputs(5004)));
    layer4_outputs(4931) <= not((layer3_outputs(5997)) xor (layer3_outputs(5327)));
    layer4_outputs(4932) <= not(layer3_outputs(2814));
    layer4_outputs(4933) <= not(layer3_outputs(4919)) or (layer3_outputs(3322));
    layer4_outputs(4934) <= layer3_outputs(1559);
    layer4_outputs(4935) <= not(layer3_outputs(3340));
    layer4_outputs(4936) <= not(layer3_outputs(721));
    layer4_outputs(4937) <= (layer3_outputs(3986)) and (layer3_outputs(1155));
    layer4_outputs(4938) <= not((layer3_outputs(4033)) xor (layer3_outputs(7540)));
    layer4_outputs(4939) <= not(layer3_outputs(1799)) or (layer3_outputs(2932));
    layer4_outputs(4940) <= (layer3_outputs(141)) and not (layer3_outputs(4165));
    layer4_outputs(4941) <= layer3_outputs(5660);
    layer4_outputs(4942) <= (layer3_outputs(3373)) and (layer3_outputs(2917));
    layer4_outputs(4943) <= not((layer3_outputs(4731)) xor (layer3_outputs(5386)));
    layer4_outputs(4944) <= not(layer3_outputs(3368));
    layer4_outputs(4945) <= not(layer3_outputs(2368)) or (layer3_outputs(4866));
    layer4_outputs(4946) <= not(layer3_outputs(7328)) or (layer3_outputs(5541));
    layer4_outputs(4947) <= not(layer3_outputs(961));
    layer4_outputs(4948) <= layer3_outputs(5344);
    layer4_outputs(4949) <= not(layer3_outputs(5675));
    layer4_outputs(4950) <= '0';
    layer4_outputs(4951) <= not((layer3_outputs(7309)) and (layer3_outputs(4255)));
    layer4_outputs(4952) <= layer3_outputs(4009);
    layer4_outputs(4953) <= (layer3_outputs(2984)) and not (layer3_outputs(1827));
    layer4_outputs(4954) <= not((layer3_outputs(4611)) xor (layer3_outputs(5250)));
    layer4_outputs(4955) <= layer3_outputs(2627);
    layer4_outputs(4956) <= (layer3_outputs(7584)) and not (layer3_outputs(2264));
    layer4_outputs(4957) <= layer3_outputs(2369);
    layer4_outputs(4958) <= not(layer3_outputs(1908));
    layer4_outputs(4959) <= not(layer3_outputs(3655));
    layer4_outputs(4960) <= layer3_outputs(3238);
    layer4_outputs(4961) <= not(layer3_outputs(564)) or (layer3_outputs(3323));
    layer4_outputs(4962) <= not(layer3_outputs(7335)) or (layer3_outputs(4857));
    layer4_outputs(4963) <= not((layer3_outputs(6884)) xor (layer3_outputs(3645)));
    layer4_outputs(4964) <= (layer3_outputs(3831)) or (layer3_outputs(1325));
    layer4_outputs(4965) <= (layer3_outputs(5306)) or (layer3_outputs(1959));
    layer4_outputs(4966) <= not((layer3_outputs(7261)) or (layer3_outputs(6643)));
    layer4_outputs(4967) <= not(layer3_outputs(6889)) or (layer3_outputs(3389));
    layer4_outputs(4968) <= (layer3_outputs(7106)) or (layer3_outputs(2857));
    layer4_outputs(4969) <= not(layer3_outputs(5114));
    layer4_outputs(4970) <= layer3_outputs(2857);
    layer4_outputs(4971) <= layer3_outputs(6070);
    layer4_outputs(4972) <= not(layer3_outputs(3360));
    layer4_outputs(4973) <= not((layer3_outputs(1317)) and (layer3_outputs(7122)));
    layer4_outputs(4974) <= not(layer3_outputs(2204));
    layer4_outputs(4975) <= layer3_outputs(1096);
    layer4_outputs(4976) <= not(layer3_outputs(3128));
    layer4_outputs(4977) <= layer3_outputs(4418);
    layer4_outputs(4978) <= layer3_outputs(3975);
    layer4_outputs(4979) <= layer3_outputs(6677);
    layer4_outputs(4980) <= (layer3_outputs(6623)) and (layer3_outputs(1776));
    layer4_outputs(4981) <= layer3_outputs(7486);
    layer4_outputs(4982) <= (layer3_outputs(5130)) and not (layer3_outputs(6900));
    layer4_outputs(4983) <= layer3_outputs(5417);
    layer4_outputs(4984) <= not(layer3_outputs(5966));
    layer4_outputs(4985) <= not((layer3_outputs(515)) and (layer3_outputs(5591)));
    layer4_outputs(4986) <= not(layer3_outputs(677));
    layer4_outputs(4987) <= not(layer3_outputs(6161)) or (layer3_outputs(3606));
    layer4_outputs(4988) <= not(layer3_outputs(4769));
    layer4_outputs(4989) <= (layer3_outputs(3779)) and not (layer3_outputs(7604));
    layer4_outputs(4990) <= not((layer3_outputs(3852)) xor (layer3_outputs(7491)));
    layer4_outputs(4991) <= layer3_outputs(1015);
    layer4_outputs(4992) <= layer3_outputs(6686);
    layer4_outputs(4993) <= (layer3_outputs(7108)) and (layer3_outputs(4374));
    layer4_outputs(4994) <= (layer3_outputs(1563)) and (layer3_outputs(563));
    layer4_outputs(4995) <= not(layer3_outputs(1476));
    layer4_outputs(4996) <= not((layer3_outputs(5673)) xor (layer3_outputs(5060)));
    layer4_outputs(4997) <= not(layer3_outputs(6330));
    layer4_outputs(4998) <= not((layer3_outputs(258)) xor (layer3_outputs(6319)));
    layer4_outputs(4999) <= layer3_outputs(5151);
    layer4_outputs(5000) <= layer3_outputs(2189);
    layer4_outputs(5001) <= (layer3_outputs(1116)) and not (layer3_outputs(4199));
    layer4_outputs(5002) <= '1';
    layer4_outputs(5003) <= (layer3_outputs(4546)) or (layer3_outputs(3651));
    layer4_outputs(5004) <= not(layer3_outputs(2908));
    layer4_outputs(5005) <= not(layer3_outputs(6248));
    layer4_outputs(5006) <= (layer3_outputs(6642)) and not (layer3_outputs(3173));
    layer4_outputs(5007) <= layer3_outputs(6839);
    layer4_outputs(5008) <= not(layer3_outputs(2228)) or (layer3_outputs(5979));
    layer4_outputs(5009) <= not(layer3_outputs(7165)) or (layer3_outputs(4889));
    layer4_outputs(5010) <= (layer3_outputs(4988)) xor (layer3_outputs(1228));
    layer4_outputs(5011) <= (layer3_outputs(6682)) and not (layer3_outputs(2299));
    layer4_outputs(5012) <= (layer3_outputs(3321)) and (layer3_outputs(4799));
    layer4_outputs(5013) <= '1';
    layer4_outputs(5014) <= (layer3_outputs(3890)) and not (layer3_outputs(4412));
    layer4_outputs(5015) <= layer3_outputs(5751);
    layer4_outputs(5016) <= not(layer3_outputs(1713)) or (layer3_outputs(1980));
    layer4_outputs(5017) <= (layer3_outputs(1492)) xor (layer3_outputs(3070));
    layer4_outputs(5018) <= (layer3_outputs(2140)) or (layer3_outputs(5001));
    layer4_outputs(5019) <= layer3_outputs(1133);
    layer4_outputs(5020) <= layer3_outputs(463);
    layer4_outputs(5021) <= (layer3_outputs(4926)) or (layer3_outputs(770));
    layer4_outputs(5022) <= layer3_outputs(4723);
    layer4_outputs(5023) <= (layer3_outputs(3872)) and not (layer3_outputs(6789));
    layer4_outputs(5024) <= (layer3_outputs(3638)) and not (layer3_outputs(1230));
    layer4_outputs(5025) <= not(layer3_outputs(3336)) or (layer3_outputs(5388));
    layer4_outputs(5026) <= '1';
    layer4_outputs(5027) <= (layer3_outputs(1631)) xor (layer3_outputs(4068));
    layer4_outputs(5028) <= (layer3_outputs(3714)) and not (layer3_outputs(1423));
    layer4_outputs(5029) <= '1';
    layer4_outputs(5030) <= (layer3_outputs(5011)) and (layer3_outputs(7074));
    layer4_outputs(5031) <= (layer3_outputs(2745)) or (layer3_outputs(6039));
    layer4_outputs(5032) <= (layer3_outputs(5580)) xor (layer3_outputs(4960));
    layer4_outputs(5033) <= (layer3_outputs(2022)) xor (layer3_outputs(1004));
    layer4_outputs(5034) <= '1';
    layer4_outputs(5035) <= not(layer3_outputs(6402));
    layer4_outputs(5036) <= not((layer3_outputs(7666)) and (layer3_outputs(7234)));
    layer4_outputs(5037) <= not((layer3_outputs(4985)) or (layer3_outputs(114)));
    layer4_outputs(5038) <= not(layer3_outputs(1932)) or (layer3_outputs(2585));
    layer4_outputs(5039) <= not(layer3_outputs(3170));
    layer4_outputs(5040) <= (layer3_outputs(5396)) and (layer3_outputs(1086));
    layer4_outputs(5041) <= not(layer3_outputs(4954));
    layer4_outputs(5042) <= (layer3_outputs(827)) and not (layer3_outputs(4500));
    layer4_outputs(5043) <= layer3_outputs(6225);
    layer4_outputs(5044) <= layer3_outputs(6353);
    layer4_outputs(5045) <= (layer3_outputs(2036)) and (layer3_outputs(1461));
    layer4_outputs(5046) <= layer3_outputs(1705);
    layer4_outputs(5047) <= not(layer3_outputs(1153));
    layer4_outputs(5048) <= not((layer3_outputs(3258)) and (layer3_outputs(7429)));
    layer4_outputs(5049) <= (layer3_outputs(6143)) and not (layer3_outputs(3150));
    layer4_outputs(5050) <= not((layer3_outputs(562)) and (layer3_outputs(5384)));
    layer4_outputs(5051) <= layer3_outputs(2082);
    layer4_outputs(5052) <= not((layer3_outputs(1566)) and (layer3_outputs(1411)));
    layer4_outputs(5053) <= layer3_outputs(7392);
    layer4_outputs(5054) <= layer3_outputs(1005);
    layer4_outputs(5055) <= not(layer3_outputs(3914)) or (layer3_outputs(1589));
    layer4_outputs(5056) <= not(layer3_outputs(2708));
    layer4_outputs(5057) <= (layer3_outputs(3866)) and not (layer3_outputs(472));
    layer4_outputs(5058) <= not(layer3_outputs(5417));
    layer4_outputs(5059) <= not((layer3_outputs(2307)) xor (layer3_outputs(1431)));
    layer4_outputs(5060) <= not(layer3_outputs(980)) or (layer3_outputs(3867));
    layer4_outputs(5061) <= not(layer3_outputs(4375));
    layer4_outputs(5062) <= '0';
    layer4_outputs(5063) <= not((layer3_outputs(6711)) or (layer3_outputs(5749)));
    layer4_outputs(5064) <= not(layer3_outputs(7478));
    layer4_outputs(5065) <= not(layer3_outputs(3670));
    layer4_outputs(5066) <= layer3_outputs(3460);
    layer4_outputs(5067) <= layer3_outputs(1519);
    layer4_outputs(5068) <= layer3_outputs(223);
    layer4_outputs(5069) <= not(layer3_outputs(6665));
    layer4_outputs(5070) <= (layer3_outputs(3254)) and not (layer3_outputs(1924));
    layer4_outputs(5071) <= not(layer3_outputs(1361));
    layer4_outputs(5072) <= layer3_outputs(7343);
    layer4_outputs(5073) <= not(layer3_outputs(1823));
    layer4_outputs(5074) <= not((layer3_outputs(4190)) and (layer3_outputs(5897)));
    layer4_outputs(5075) <= '0';
    layer4_outputs(5076) <= not(layer3_outputs(1596));
    layer4_outputs(5077) <= not(layer3_outputs(3201)) or (layer3_outputs(5138));
    layer4_outputs(5078) <= not(layer3_outputs(6134));
    layer4_outputs(5079) <= not(layer3_outputs(5525)) or (layer3_outputs(4201));
    layer4_outputs(5080) <= layer3_outputs(7251);
    layer4_outputs(5081) <= '1';
    layer4_outputs(5082) <= (layer3_outputs(1288)) and (layer3_outputs(3284));
    layer4_outputs(5083) <= layer3_outputs(6364);
    layer4_outputs(5084) <= not((layer3_outputs(6480)) xor (layer3_outputs(6106)));
    layer4_outputs(5085) <= (layer3_outputs(3069)) or (layer3_outputs(7014));
    layer4_outputs(5086) <= '1';
    layer4_outputs(5087) <= layer3_outputs(6974);
    layer4_outputs(5088) <= not((layer3_outputs(6342)) or (layer3_outputs(2822)));
    layer4_outputs(5089) <= not(layer3_outputs(1723));
    layer4_outputs(5090) <= not((layer3_outputs(5999)) xor (layer3_outputs(2131)));
    layer4_outputs(5091) <= (layer3_outputs(5010)) and not (layer3_outputs(2019));
    layer4_outputs(5092) <= layer3_outputs(2574);
    layer4_outputs(5093) <= (layer3_outputs(3512)) or (layer3_outputs(1995));
    layer4_outputs(5094) <= (layer3_outputs(2154)) and not (layer3_outputs(5598));
    layer4_outputs(5095) <= not((layer3_outputs(2657)) or (layer3_outputs(1110)));
    layer4_outputs(5096) <= (layer3_outputs(1555)) or (layer3_outputs(7177));
    layer4_outputs(5097) <= (layer3_outputs(971)) and not (layer3_outputs(4513));
    layer4_outputs(5098) <= '1';
    layer4_outputs(5099) <= (layer3_outputs(5594)) and not (layer3_outputs(5161));
    layer4_outputs(5100) <= (layer3_outputs(1993)) or (layer3_outputs(1652));
    layer4_outputs(5101) <= not(layer3_outputs(4943)) or (layer3_outputs(2794));
    layer4_outputs(5102) <= layer3_outputs(2163);
    layer4_outputs(5103) <= (layer3_outputs(3255)) and not (layer3_outputs(1630));
    layer4_outputs(5104) <= (layer3_outputs(5209)) and not (layer3_outputs(1790));
    layer4_outputs(5105) <= not(layer3_outputs(238));
    layer4_outputs(5106) <= not(layer3_outputs(6036));
    layer4_outputs(5107) <= not(layer3_outputs(6420));
    layer4_outputs(5108) <= '0';
    layer4_outputs(5109) <= not((layer3_outputs(7341)) and (layer3_outputs(2849)));
    layer4_outputs(5110) <= not(layer3_outputs(5815));
    layer4_outputs(5111) <= (layer3_outputs(2728)) and (layer3_outputs(7521));
    layer4_outputs(5112) <= layer3_outputs(1189);
    layer4_outputs(5113) <= (layer3_outputs(4203)) and not (layer3_outputs(4133));
    layer4_outputs(5114) <= layer3_outputs(4288);
    layer4_outputs(5115) <= layer3_outputs(2716);
    layer4_outputs(5116) <= not(layer3_outputs(6218));
    layer4_outputs(5117) <= not(layer3_outputs(6790));
    layer4_outputs(5118) <= not((layer3_outputs(7229)) xor (layer3_outputs(5875)));
    layer4_outputs(5119) <= not((layer3_outputs(3236)) or (layer3_outputs(469)));
    layer4_outputs(5120) <= not((layer3_outputs(5734)) xor (layer3_outputs(3405)));
    layer4_outputs(5121) <= layer3_outputs(6887);
    layer4_outputs(5122) <= not(layer3_outputs(332));
    layer4_outputs(5123) <= layer3_outputs(6156);
    layer4_outputs(5124) <= '1';
    layer4_outputs(5125) <= not(layer3_outputs(6547));
    layer4_outputs(5126) <= (layer3_outputs(6001)) or (layer3_outputs(6460));
    layer4_outputs(5127) <= (layer3_outputs(586)) and (layer3_outputs(3562));
    layer4_outputs(5128) <= layer3_outputs(7253);
    layer4_outputs(5129) <= (layer3_outputs(2033)) or (layer3_outputs(4345));
    layer4_outputs(5130) <= not((layer3_outputs(1316)) and (layer3_outputs(3432)));
    layer4_outputs(5131) <= layer3_outputs(2352);
    layer4_outputs(5132) <= not(layer3_outputs(1120));
    layer4_outputs(5133) <= (layer3_outputs(2387)) or (layer3_outputs(733));
    layer4_outputs(5134) <= (layer3_outputs(4824)) and not (layer3_outputs(2646));
    layer4_outputs(5135) <= not(layer3_outputs(5340));
    layer4_outputs(5136) <= '1';
    layer4_outputs(5137) <= not((layer3_outputs(6637)) and (layer3_outputs(339)));
    layer4_outputs(5138) <= not(layer3_outputs(4779)) or (layer3_outputs(3532));
    layer4_outputs(5139) <= not((layer3_outputs(7522)) xor (layer3_outputs(5550)));
    layer4_outputs(5140) <= '0';
    layer4_outputs(5141) <= (layer3_outputs(6412)) and not (layer3_outputs(3219));
    layer4_outputs(5142) <= layer3_outputs(1282);
    layer4_outputs(5143) <= not((layer3_outputs(5300)) or (layer3_outputs(7431)));
    layer4_outputs(5144) <= not(layer3_outputs(6074));
    layer4_outputs(5145) <= layer3_outputs(499);
    layer4_outputs(5146) <= '1';
    layer4_outputs(5147) <= not((layer3_outputs(779)) and (layer3_outputs(697)));
    layer4_outputs(5148) <= not(layer3_outputs(1243)) or (layer3_outputs(2886));
    layer4_outputs(5149) <= layer3_outputs(4025);
    layer4_outputs(5150) <= not((layer3_outputs(7439)) or (layer3_outputs(7610)));
    layer4_outputs(5151) <= layer3_outputs(3534);
    layer4_outputs(5152) <= not(layer3_outputs(1417));
    layer4_outputs(5153) <= not(layer3_outputs(5813));
    layer4_outputs(5154) <= not(layer3_outputs(4347));
    layer4_outputs(5155) <= '1';
    layer4_outputs(5156) <= not(layer3_outputs(7548));
    layer4_outputs(5157) <= not(layer3_outputs(1412));
    layer4_outputs(5158) <= (layer3_outputs(2919)) and not (layer3_outputs(5494));
    layer4_outputs(5159) <= layer3_outputs(4644);
    layer4_outputs(5160) <= not(layer3_outputs(6377));
    layer4_outputs(5161) <= not(layer3_outputs(3505));
    layer4_outputs(5162) <= not(layer3_outputs(175)) or (layer3_outputs(2865));
    layer4_outputs(5163) <= not(layer3_outputs(6185));
    layer4_outputs(5164) <= not(layer3_outputs(3333)) or (layer3_outputs(5830));
    layer4_outputs(5165) <= not((layer3_outputs(2104)) and (layer3_outputs(2758)));
    layer4_outputs(5166) <= not(layer3_outputs(6263));
    layer4_outputs(5167) <= not(layer3_outputs(4320));
    layer4_outputs(5168) <= not(layer3_outputs(6477));
    layer4_outputs(5169) <= (layer3_outputs(4823)) and (layer3_outputs(3626));
    layer4_outputs(5170) <= (layer3_outputs(5827)) and not (layer3_outputs(1852));
    layer4_outputs(5171) <= '0';
    layer4_outputs(5172) <= layer3_outputs(793);
    layer4_outputs(5173) <= (layer3_outputs(6522)) or (layer3_outputs(512));
    layer4_outputs(5174) <= not(layer3_outputs(4605)) or (layer3_outputs(4364));
    layer4_outputs(5175) <= (layer3_outputs(3902)) and not (layer3_outputs(492));
    layer4_outputs(5176) <= not(layer3_outputs(5723));
    layer4_outputs(5177) <= not(layer3_outputs(6202));
    layer4_outputs(5178) <= layer3_outputs(3409);
    layer4_outputs(5179) <= not((layer3_outputs(5938)) and (layer3_outputs(6232)));
    layer4_outputs(5180) <= layer3_outputs(6613);
    layer4_outputs(5181) <= (layer3_outputs(2707)) and not (layer3_outputs(5272));
    layer4_outputs(5182) <= layer3_outputs(3523);
    layer4_outputs(5183) <= not(layer3_outputs(7653));
    layer4_outputs(5184) <= layer3_outputs(7428);
    layer4_outputs(5185) <= layer3_outputs(5853);
    layer4_outputs(5186) <= layer3_outputs(2949);
    layer4_outputs(5187) <= not(layer3_outputs(6005));
    layer4_outputs(5188) <= (layer3_outputs(7299)) xor (layer3_outputs(3241));
    layer4_outputs(5189) <= layer3_outputs(1245);
    layer4_outputs(5190) <= not(layer3_outputs(134));
    layer4_outputs(5191) <= not(layer3_outputs(3162));
    layer4_outputs(5192) <= (layer3_outputs(3974)) and (layer3_outputs(730));
    layer4_outputs(5193) <= layer3_outputs(584);
    layer4_outputs(5194) <= not((layer3_outputs(1133)) xor (layer3_outputs(2993)));
    layer4_outputs(5195) <= layer3_outputs(4542);
    layer4_outputs(5196) <= (layer3_outputs(1474)) and not (layer3_outputs(7111));
    layer4_outputs(5197) <= '0';
    layer4_outputs(5198) <= (layer3_outputs(3871)) or (layer3_outputs(657));
    layer4_outputs(5199) <= (layer3_outputs(7646)) and not (layer3_outputs(341));
    layer4_outputs(5200) <= not(layer3_outputs(2927)) or (layer3_outputs(2289));
    layer4_outputs(5201) <= not(layer3_outputs(2267));
    layer4_outputs(5202) <= layer3_outputs(5642);
    layer4_outputs(5203) <= not(layer3_outputs(6864)) or (layer3_outputs(6463));
    layer4_outputs(5204) <= layer3_outputs(5588);
    layer4_outputs(5205) <= (layer3_outputs(365)) or (layer3_outputs(6529));
    layer4_outputs(5206) <= not((layer3_outputs(4760)) xor (layer3_outputs(3700)));
    layer4_outputs(5207) <= not((layer3_outputs(2363)) or (layer3_outputs(287)));
    layer4_outputs(5208) <= not(layer3_outputs(4865));
    layer4_outputs(5209) <= not(layer3_outputs(5695));
    layer4_outputs(5210) <= not(layer3_outputs(548));
    layer4_outputs(5211) <= layer3_outputs(7269);
    layer4_outputs(5212) <= (layer3_outputs(6170)) xor (layer3_outputs(6359));
    layer4_outputs(5213) <= not(layer3_outputs(2708));
    layer4_outputs(5214) <= (layer3_outputs(7576)) and not (layer3_outputs(3654));
    layer4_outputs(5215) <= not((layer3_outputs(1171)) and (layer3_outputs(1461)));
    layer4_outputs(5216) <= layer3_outputs(324);
    layer4_outputs(5217) <= (layer3_outputs(5504)) and not (layer3_outputs(7583));
    layer4_outputs(5218) <= (layer3_outputs(7357)) and not (layer3_outputs(403));
    layer4_outputs(5219) <= (layer3_outputs(4652)) and not (layer3_outputs(1744));
    layer4_outputs(5220) <= not(layer3_outputs(6827)) or (layer3_outputs(6650));
    layer4_outputs(5221) <= layer3_outputs(5896);
    layer4_outputs(5222) <= (layer3_outputs(7087)) xor (layer3_outputs(5260));
    layer4_outputs(5223) <= not(layer3_outputs(1266));
    layer4_outputs(5224) <= (layer3_outputs(3925)) and (layer3_outputs(4764));
    layer4_outputs(5225) <= (layer3_outputs(2545)) or (layer3_outputs(4222));
    layer4_outputs(5226) <= not(layer3_outputs(6447));
    layer4_outputs(5227) <= not((layer3_outputs(4097)) or (layer3_outputs(2572)));
    layer4_outputs(5228) <= not(layer3_outputs(5512));
    layer4_outputs(5229) <= (layer3_outputs(5820)) and (layer3_outputs(6413));
    layer4_outputs(5230) <= layer3_outputs(1352);
    layer4_outputs(5231) <= '1';
    layer4_outputs(5232) <= layer3_outputs(928);
    layer4_outputs(5233) <= not(layer3_outputs(4713)) or (layer3_outputs(3064));
    layer4_outputs(5234) <= not((layer3_outputs(895)) xor (layer3_outputs(5771)));
    layer4_outputs(5235) <= (layer3_outputs(4357)) or (layer3_outputs(2419));
    layer4_outputs(5236) <= (layer3_outputs(3826)) or (layer3_outputs(7176));
    layer4_outputs(5237) <= (layer3_outputs(3218)) and (layer3_outputs(2385));
    layer4_outputs(5238) <= layer3_outputs(3352);
    layer4_outputs(5239) <= not(layer3_outputs(1258));
    layer4_outputs(5240) <= (layer3_outputs(3369)) or (layer3_outputs(7498));
    layer4_outputs(5241) <= layer3_outputs(1347);
    layer4_outputs(5242) <= layer3_outputs(6708);
    layer4_outputs(5243) <= not(layer3_outputs(5427));
    layer4_outputs(5244) <= (layer3_outputs(498)) and (layer3_outputs(1865));
    layer4_outputs(5245) <= not(layer3_outputs(1295));
    layer4_outputs(5246) <= not(layer3_outputs(144));
    layer4_outputs(5247) <= (layer3_outputs(6339)) and (layer3_outputs(7477));
    layer4_outputs(5248) <= not(layer3_outputs(1591));
    layer4_outputs(5249) <= layer3_outputs(4729);
    layer4_outputs(5250) <= not(layer3_outputs(5173));
    layer4_outputs(5251) <= not((layer3_outputs(6959)) and (layer3_outputs(6065)));
    layer4_outputs(5252) <= '1';
    layer4_outputs(5253) <= (layer3_outputs(5780)) and not (layer3_outputs(386));
    layer4_outputs(5254) <= layer3_outputs(5710);
    layer4_outputs(5255) <= layer3_outputs(1716);
    layer4_outputs(5256) <= not((layer3_outputs(5515)) and (layer3_outputs(6003)));
    layer4_outputs(5257) <= '0';
    layer4_outputs(5258) <= not(layer3_outputs(694));
    layer4_outputs(5259) <= (layer3_outputs(7580)) and (layer3_outputs(2234));
    layer4_outputs(5260) <= (layer3_outputs(1599)) and (layer3_outputs(7152));
    layer4_outputs(5261) <= not((layer3_outputs(833)) and (layer3_outputs(2870)));
    layer4_outputs(5262) <= layer3_outputs(89);
    layer4_outputs(5263) <= not(layer3_outputs(5453));
    layer4_outputs(5264) <= not(layer3_outputs(3161)) or (layer3_outputs(6937));
    layer4_outputs(5265) <= (layer3_outputs(3229)) and (layer3_outputs(693));
    layer4_outputs(5266) <= not(layer3_outputs(5869));
    layer4_outputs(5267) <= not((layer3_outputs(6744)) xor (layer3_outputs(6313)));
    layer4_outputs(5268) <= not(layer3_outputs(5848)) or (layer3_outputs(7208));
    layer4_outputs(5269) <= not(layer3_outputs(3140)) or (layer3_outputs(6609));
    layer4_outputs(5270) <= layer3_outputs(6750);
    layer4_outputs(5271) <= (layer3_outputs(2800)) xor (layer3_outputs(424));
    layer4_outputs(5272) <= (layer3_outputs(5062)) and not (layer3_outputs(2239));
    layer4_outputs(5273) <= not(layer3_outputs(124)) or (layer3_outputs(4327));
    layer4_outputs(5274) <= layer3_outputs(4930);
    layer4_outputs(5275) <= '1';
    layer4_outputs(5276) <= not(layer3_outputs(5027));
    layer4_outputs(5277) <= (layer3_outputs(6349)) and (layer3_outputs(4615));
    layer4_outputs(5278) <= (layer3_outputs(3239)) xor (layer3_outputs(3478));
    layer4_outputs(5279) <= (layer3_outputs(3024)) or (layer3_outputs(3167));
    layer4_outputs(5280) <= (layer3_outputs(3893)) or (layer3_outputs(4648));
    layer4_outputs(5281) <= not(layer3_outputs(6257));
    layer4_outputs(5282) <= (layer3_outputs(7312)) or (layer3_outputs(7321));
    layer4_outputs(5283) <= (layer3_outputs(3417)) and not (layer3_outputs(7003));
    layer4_outputs(5284) <= layer3_outputs(5045);
    layer4_outputs(5285) <= not((layer3_outputs(868)) and (layer3_outputs(4471)));
    layer4_outputs(5286) <= not(layer3_outputs(5688)) or (layer3_outputs(6453));
    layer4_outputs(5287) <= layer3_outputs(2047);
    layer4_outputs(5288) <= '1';
    layer4_outputs(5289) <= layer3_outputs(1472);
    layer4_outputs(5290) <= not(layer3_outputs(1660)) or (layer3_outputs(7673));
    layer4_outputs(5291) <= layer3_outputs(240);
    layer4_outputs(5292) <= (layer3_outputs(700)) and (layer3_outputs(2606));
    layer4_outputs(5293) <= '1';
    layer4_outputs(5294) <= not((layer3_outputs(4646)) or (layer3_outputs(3811)));
    layer4_outputs(5295) <= layer3_outputs(3665);
    layer4_outputs(5296) <= not(layer3_outputs(4405));
    layer4_outputs(5297) <= (layer3_outputs(5590)) and (layer3_outputs(2319));
    layer4_outputs(5298) <= layer3_outputs(3957);
    layer4_outputs(5299) <= (layer3_outputs(6280)) and not (layer3_outputs(1112));
    layer4_outputs(5300) <= not(layer3_outputs(1313)) or (layer3_outputs(6541));
    layer4_outputs(5301) <= layer3_outputs(2254);
    layer4_outputs(5302) <= (layer3_outputs(5658)) and not (layer3_outputs(6734));
    layer4_outputs(5303) <= (layer3_outputs(5872)) xor (layer3_outputs(1721));
    layer4_outputs(5304) <= not(layer3_outputs(3090));
    layer4_outputs(5305) <= not(layer3_outputs(6136));
    layer4_outputs(5306) <= (layer3_outputs(6540)) and (layer3_outputs(227));
    layer4_outputs(5307) <= layer3_outputs(6140);
    layer4_outputs(5308) <= not((layer3_outputs(530)) and (layer3_outputs(6183)));
    layer4_outputs(5309) <= not((layer3_outputs(2432)) and (layer3_outputs(1931)));
    layer4_outputs(5310) <= not((layer3_outputs(2625)) or (layer3_outputs(7594)));
    layer4_outputs(5311) <= '0';
    layer4_outputs(5312) <= (layer3_outputs(1397)) and not (layer3_outputs(6213));
    layer4_outputs(5313) <= (layer3_outputs(122)) and not (layer3_outputs(5150));
    layer4_outputs(5314) <= (layer3_outputs(5577)) and not (layer3_outputs(4756));
    layer4_outputs(5315) <= not(layer3_outputs(6365)) or (layer3_outputs(1226));
    layer4_outputs(5316) <= layer3_outputs(6247);
    layer4_outputs(5317) <= layer3_outputs(3187);
    layer4_outputs(5318) <= not(layer3_outputs(3365)) or (layer3_outputs(36));
    layer4_outputs(5319) <= not(layer3_outputs(3917)) or (layer3_outputs(5141));
    layer4_outputs(5320) <= layer3_outputs(7336);
    layer4_outputs(5321) <= (layer3_outputs(3421)) and not (layer3_outputs(6624));
    layer4_outputs(5322) <= (layer3_outputs(1809)) and not (layer3_outputs(5714));
    layer4_outputs(5323) <= not(layer3_outputs(6839)) or (layer3_outputs(4985));
    layer4_outputs(5324) <= layer3_outputs(821);
    layer4_outputs(5325) <= layer3_outputs(7076);
    layer4_outputs(5326) <= not((layer3_outputs(1903)) xor (layer3_outputs(683)));
    layer4_outputs(5327) <= (layer3_outputs(2580)) and (layer3_outputs(6530));
    layer4_outputs(5328) <= not(layer3_outputs(4200));
    layer4_outputs(5329) <= not(layer3_outputs(6274));
    layer4_outputs(5330) <= not(layer3_outputs(2447)) or (layer3_outputs(4725));
    layer4_outputs(5331) <= not(layer3_outputs(4350));
    layer4_outputs(5332) <= not((layer3_outputs(7589)) or (layer3_outputs(3513)));
    layer4_outputs(5333) <= (layer3_outputs(5993)) xor (layer3_outputs(4650));
    layer4_outputs(5334) <= not(layer3_outputs(2482));
    layer4_outputs(5335) <= layer3_outputs(4062);
    layer4_outputs(5336) <= layer3_outputs(1186);
    layer4_outputs(5337) <= layer3_outputs(3776);
    layer4_outputs(5338) <= layer3_outputs(3310);
    layer4_outputs(5339) <= (layer3_outputs(1799)) and (layer3_outputs(5081));
    layer4_outputs(5340) <= not((layer3_outputs(1823)) and (layer3_outputs(2404)));
    layer4_outputs(5341) <= '0';
    layer4_outputs(5342) <= layer3_outputs(3951);
    layer4_outputs(5343) <= layer3_outputs(3873);
    layer4_outputs(5344) <= not(layer3_outputs(2106));
    layer4_outputs(5345) <= (layer3_outputs(6764)) xor (layer3_outputs(6394));
    layer4_outputs(5346) <= layer3_outputs(7432);
    layer4_outputs(5347) <= not(layer3_outputs(1668)) or (layer3_outputs(3502));
    layer4_outputs(5348) <= not(layer3_outputs(6721));
    layer4_outputs(5349) <= layer3_outputs(742);
    layer4_outputs(5350) <= (layer3_outputs(5581)) and not (layer3_outputs(116));
    layer4_outputs(5351) <= layer3_outputs(2869);
    layer4_outputs(5352) <= (layer3_outputs(5837)) and not (layer3_outputs(5864));
    layer4_outputs(5353) <= (layer3_outputs(6398)) xor (layer3_outputs(6385));
    layer4_outputs(5354) <= (layer3_outputs(4379)) or (layer3_outputs(6310));
    layer4_outputs(5355) <= not(layer3_outputs(2137));
    layer4_outputs(5356) <= (layer3_outputs(7281)) and (layer3_outputs(7609));
    layer4_outputs(5357) <= not(layer3_outputs(4900));
    layer4_outputs(5358) <= layer3_outputs(333);
    layer4_outputs(5359) <= (layer3_outputs(402)) xor (layer3_outputs(858));
    layer4_outputs(5360) <= (layer3_outputs(7214)) xor (layer3_outputs(7526));
    layer4_outputs(5361) <= (layer3_outputs(1094)) and not (layer3_outputs(1813));
    layer4_outputs(5362) <= layer3_outputs(82);
    layer4_outputs(5363) <= not(layer3_outputs(1742));
    layer4_outputs(5364) <= not(layer3_outputs(3477));
    layer4_outputs(5365) <= not(layer3_outputs(6616));
    layer4_outputs(5366) <= layer3_outputs(2372);
    layer4_outputs(5367) <= not(layer3_outputs(4697));
    layer4_outputs(5368) <= not(layer3_outputs(2946));
    layer4_outputs(5369) <= layer3_outputs(5893);
    layer4_outputs(5370) <= not(layer3_outputs(688));
    layer4_outputs(5371) <= (layer3_outputs(6191)) and (layer3_outputs(3050));
    layer4_outputs(5372) <= (layer3_outputs(6037)) xor (layer3_outputs(6516));
    layer4_outputs(5373) <= not(layer3_outputs(6816));
    layer4_outputs(5374) <= layer3_outputs(533);
    layer4_outputs(5375) <= not(layer3_outputs(3401));
    layer4_outputs(5376) <= (layer3_outputs(3119)) and not (layer3_outputs(5461));
    layer4_outputs(5377) <= not(layer3_outputs(4873));
    layer4_outputs(5378) <= layer3_outputs(5635);
    layer4_outputs(5379) <= not(layer3_outputs(911));
    layer4_outputs(5380) <= not(layer3_outputs(5884));
    layer4_outputs(5381) <= '0';
    layer4_outputs(5382) <= not(layer3_outputs(3708));
    layer4_outputs(5383) <= not(layer3_outputs(654)) or (layer3_outputs(4936));
    layer4_outputs(5384) <= '0';
    layer4_outputs(5385) <= (layer3_outputs(7405)) and not (layer3_outputs(1691));
    layer4_outputs(5386) <= not(layer3_outputs(2399));
    layer4_outputs(5387) <= (layer3_outputs(5431)) and not (layer3_outputs(4571));
    layer4_outputs(5388) <= not(layer3_outputs(2188));
    layer4_outputs(5389) <= not(layer3_outputs(3640));
    layer4_outputs(5390) <= '1';
    layer4_outputs(5391) <= layer3_outputs(5191);
    layer4_outputs(5392) <= (layer3_outputs(7417)) and not (layer3_outputs(5582));
    layer4_outputs(5393) <= not(layer3_outputs(7153));
    layer4_outputs(5394) <= not(layer3_outputs(4224)) or (layer3_outputs(6462));
    layer4_outputs(5395) <= not(layer3_outputs(5872));
    layer4_outputs(5396) <= layer3_outputs(1142);
    layer4_outputs(5397) <= '1';
    layer4_outputs(5398) <= not(layer3_outputs(5221));
    layer4_outputs(5399) <= not(layer3_outputs(5587)) or (layer3_outputs(737));
    layer4_outputs(5400) <= layer3_outputs(2284);
    layer4_outputs(5401) <= (layer3_outputs(361)) or (layer3_outputs(5949));
    layer4_outputs(5402) <= (layer3_outputs(5439)) and (layer3_outputs(2888));
    layer4_outputs(5403) <= (layer3_outputs(5126)) and not (layer3_outputs(3958));
    layer4_outputs(5404) <= not(layer3_outputs(7280));
    layer4_outputs(5405) <= not((layer3_outputs(6311)) and (layer3_outputs(4430)));
    layer4_outputs(5406) <= layer3_outputs(187);
    layer4_outputs(5407) <= not(layer3_outputs(6320));
    layer4_outputs(5408) <= '0';
    layer4_outputs(5409) <= (layer3_outputs(2328)) and not (layer3_outputs(7130));
    layer4_outputs(5410) <= not((layer3_outputs(5374)) xor (layer3_outputs(4405)));
    layer4_outputs(5411) <= '1';
    layer4_outputs(5412) <= layer3_outputs(6806);
    layer4_outputs(5413) <= not(layer3_outputs(3077));
    layer4_outputs(5414) <= not(layer3_outputs(6686));
    layer4_outputs(5415) <= (layer3_outputs(6284)) and not (layer3_outputs(2997));
    layer4_outputs(5416) <= '1';
    layer4_outputs(5417) <= '1';
    layer4_outputs(5418) <= layer3_outputs(4771);
    layer4_outputs(5419) <= (layer3_outputs(5852)) and (layer3_outputs(5400));
    layer4_outputs(5420) <= layer3_outputs(6821);
    layer4_outputs(5421) <= layer3_outputs(4412);
    layer4_outputs(5422) <= not(layer3_outputs(6739));
    layer4_outputs(5423) <= not(layer3_outputs(5166)) or (layer3_outputs(2144));
    layer4_outputs(5424) <= not((layer3_outputs(890)) and (layer3_outputs(4481)));
    layer4_outputs(5425) <= not(layer3_outputs(1331));
    layer4_outputs(5426) <= (layer3_outputs(4441)) and (layer3_outputs(1217));
    layer4_outputs(5427) <= layer3_outputs(2189);
    layer4_outputs(5428) <= not(layer3_outputs(1508));
    layer4_outputs(5429) <= (layer3_outputs(6278)) or (layer3_outputs(812));
    layer4_outputs(5430) <= not((layer3_outputs(1161)) and (layer3_outputs(6768)));
    layer4_outputs(5431) <= (layer3_outputs(1708)) and not (layer3_outputs(6774));
    layer4_outputs(5432) <= layer3_outputs(732);
    layer4_outputs(5433) <= not((layer3_outputs(6719)) or (layer3_outputs(6573)));
    layer4_outputs(5434) <= not(layer3_outputs(571)) or (layer3_outputs(5085));
    layer4_outputs(5435) <= not((layer3_outputs(5083)) or (layer3_outputs(4139)));
    layer4_outputs(5436) <= layer3_outputs(1372);
    layer4_outputs(5437) <= not((layer3_outputs(1522)) or (layer3_outputs(1590)));
    layer4_outputs(5438) <= layer3_outputs(4443);
    layer4_outputs(5439) <= layer3_outputs(740);
    layer4_outputs(5440) <= layer3_outputs(6279);
    layer4_outputs(5441) <= not(layer3_outputs(5456));
    layer4_outputs(5442) <= not((layer3_outputs(996)) or (layer3_outputs(6182)));
    layer4_outputs(5443) <= (layer3_outputs(994)) and not (layer3_outputs(4768));
    layer4_outputs(5444) <= (layer3_outputs(1651)) or (layer3_outputs(4140));
    layer4_outputs(5445) <= layer3_outputs(6415);
    layer4_outputs(5446) <= '1';
    layer4_outputs(5447) <= not(layer3_outputs(576));
    layer4_outputs(5448) <= (layer3_outputs(6578)) and (layer3_outputs(2427));
    layer4_outputs(5449) <= layer3_outputs(4634);
    layer4_outputs(5450) <= not(layer3_outputs(1311)) or (layer3_outputs(304));
    layer4_outputs(5451) <= not((layer3_outputs(6770)) and (layer3_outputs(6873)));
    layer4_outputs(5452) <= '1';
    layer4_outputs(5453) <= (layer3_outputs(3528)) and not (layer3_outputs(6167));
    layer4_outputs(5454) <= not(layer3_outputs(3347)) or (layer3_outputs(4921));
    layer4_outputs(5455) <= not((layer3_outputs(6469)) or (layer3_outputs(6938)));
    layer4_outputs(5456) <= not(layer3_outputs(1193));
    layer4_outputs(5457) <= not(layer3_outputs(3785)) or (layer3_outputs(1303));
    layer4_outputs(5458) <= layer3_outputs(4091);
    layer4_outputs(5459) <= not(layer3_outputs(186));
    layer4_outputs(5460) <= '0';
    layer4_outputs(5461) <= layer3_outputs(2001);
    layer4_outputs(5462) <= (layer3_outputs(577)) and not (layer3_outputs(3560));
    layer4_outputs(5463) <= (layer3_outputs(204)) xor (layer3_outputs(53));
    layer4_outputs(5464) <= (layer3_outputs(219)) and (layer3_outputs(643));
    layer4_outputs(5465) <= not((layer3_outputs(5673)) or (layer3_outputs(1122)));
    layer4_outputs(5466) <= (layer3_outputs(4734)) or (layer3_outputs(6633));
    layer4_outputs(5467) <= not(layer3_outputs(659));
    layer4_outputs(5468) <= not(layer3_outputs(2720)) or (layer3_outputs(1348));
    layer4_outputs(5469) <= layer3_outputs(669);
    layer4_outputs(5470) <= layer3_outputs(3810);
    layer4_outputs(5471) <= not(layer3_outputs(45));
    layer4_outputs(5472) <= layer3_outputs(2329);
    layer4_outputs(5473) <= (layer3_outputs(5378)) or (layer3_outputs(5073));
    layer4_outputs(5474) <= '1';
    layer4_outputs(5475) <= not(layer3_outputs(5653));
    layer4_outputs(5476) <= (layer3_outputs(1638)) and (layer3_outputs(7020));
    layer4_outputs(5477) <= layer3_outputs(5574);
    layer4_outputs(5478) <= (layer3_outputs(255)) and (layer3_outputs(6831));
    layer4_outputs(5479) <= not(layer3_outputs(7291)) or (layer3_outputs(5228));
    layer4_outputs(5480) <= not(layer3_outputs(7418));
    layer4_outputs(5481) <= not((layer3_outputs(2105)) and (layer3_outputs(5012)));
    layer4_outputs(5482) <= not(layer3_outputs(7206)) or (layer3_outputs(6108));
    layer4_outputs(5483) <= (layer3_outputs(6473)) or (layer3_outputs(7337));
    layer4_outputs(5484) <= not(layer3_outputs(7227)) or (layer3_outputs(4983));
    layer4_outputs(5485) <= (layer3_outputs(6926)) or (layer3_outputs(1068));
    layer4_outputs(5486) <= (layer3_outputs(5833)) xor (layer3_outputs(3271));
    layer4_outputs(5487) <= not((layer3_outputs(2212)) and (layer3_outputs(5495)));
    layer4_outputs(5488) <= (layer3_outputs(302)) and not (layer3_outputs(5542));
    layer4_outputs(5489) <= (layer3_outputs(1913)) and not (layer3_outputs(6533));
    layer4_outputs(5490) <= not(layer3_outputs(3913));
    layer4_outputs(5491) <= not(layer3_outputs(7399));
    layer4_outputs(5492) <= '1';
    layer4_outputs(5493) <= (layer3_outputs(3798)) and not (layer3_outputs(6448));
    layer4_outputs(5494) <= (layer3_outputs(2148)) or (layer3_outputs(1559));
    layer4_outputs(5495) <= (layer3_outputs(2365)) and (layer3_outputs(6126));
    layer4_outputs(5496) <= not(layer3_outputs(4082));
    layer4_outputs(5497) <= not(layer3_outputs(5915));
    layer4_outputs(5498) <= layer3_outputs(922);
    layer4_outputs(5499) <= not(layer3_outputs(3819));
    layer4_outputs(5500) <= (layer3_outputs(6065)) or (layer3_outputs(712));
    layer4_outputs(5501) <= (layer3_outputs(2624)) and (layer3_outputs(1434));
    layer4_outputs(5502) <= layer3_outputs(3834);
    layer4_outputs(5503) <= not(layer3_outputs(2974));
    layer4_outputs(5504) <= layer3_outputs(6840);
    layer4_outputs(5505) <= '1';
    layer4_outputs(5506) <= not(layer3_outputs(6358)) or (layer3_outputs(3065));
    layer4_outputs(5507) <= '1';
    layer4_outputs(5508) <= '1';
    layer4_outputs(5509) <= layer3_outputs(738);
    layer4_outputs(5510) <= not(layer3_outputs(2231));
    layer4_outputs(5511) <= layer3_outputs(4419);
    layer4_outputs(5512) <= not(layer3_outputs(763)) or (layer3_outputs(5371));
    layer4_outputs(5513) <= not(layer3_outputs(1576));
    layer4_outputs(5514) <= not((layer3_outputs(6600)) xor (layer3_outputs(5764)));
    layer4_outputs(5515) <= not((layer3_outputs(7500)) xor (layer3_outputs(5317)));
    layer4_outputs(5516) <= layer3_outputs(5614);
    layer4_outputs(5517) <= not(layer3_outputs(2886));
    layer4_outputs(5518) <= layer3_outputs(1574);
    layer4_outputs(5519) <= not(layer3_outputs(2817));
    layer4_outputs(5520) <= (layer3_outputs(2550)) and not (layer3_outputs(3737));
    layer4_outputs(5521) <= not(layer3_outputs(273));
    layer4_outputs(5522) <= (layer3_outputs(4325)) or (layer3_outputs(2012));
    layer4_outputs(5523) <= (layer3_outputs(3522)) and (layer3_outputs(399));
    layer4_outputs(5524) <= (layer3_outputs(2757)) or (layer3_outputs(6449));
    layer4_outputs(5525) <= not(layer3_outputs(192));
    layer4_outputs(5526) <= '0';
    layer4_outputs(5527) <= (layer3_outputs(6612)) and (layer3_outputs(3144));
    layer4_outputs(5528) <= '1';
    layer4_outputs(5529) <= not(layer3_outputs(5509));
    layer4_outputs(5530) <= not(layer3_outputs(7273)) or (layer3_outputs(3551));
    layer4_outputs(5531) <= layer3_outputs(1551);
    layer4_outputs(5532) <= (layer3_outputs(2335)) and not (layer3_outputs(56));
    layer4_outputs(5533) <= not(layer3_outputs(2230));
    layer4_outputs(5534) <= (layer3_outputs(1067)) or (layer3_outputs(1788));
    layer4_outputs(5535) <= (layer3_outputs(1079)) and (layer3_outputs(3901));
    layer4_outputs(5536) <= (layer3_outputs(3101)) and not (layer3_outputs(4148));
    layer4_outputs(5537) <= not(layer3_outputs(1318));
    layer4_outputs(5538) <= not(layer3_outputs(5442));
    layer4_outputs(5539) <= (layer3_outputs(1669)) and not (layer3_outputs(7678));
    layer4_outputs(5540) <= (layer3_outputs(3844)) and (layer3_outputs(1499));
    layer4_outputs(5541) <= '1';
    layer4_outputs(5542) <= not(layer3_outputs(326)) or (layer3_outputs(7135));
    layer4_outputs(5543) <= layer3_outputs(1918);
    layer4_outputs(5544) <= (layer3_outputs(4975)) and not (layer3_outputs(4544));
    layer4_outputs(5545) <= not(layer3_outputs(5145)) or (layer3_outputs(2966));
    layer4_outputs(5546) <= layer3_outputs(6962);
    layer4_outputs(5547) <= not(layer3_outputs(4191));
    layer4_outputs(5548) <= layer3_outputs(232);
    layer4_outputs(5549) <= layer3_outputs(2142);
    layer4_outputs(5550) <= layer3_outputs(1205);
    layer4_outputs(5551) <= layer3_outputs(6432);
    layer4_outputs(5552) <= not((layer3_outputs(3519)) and (layer3_outputs(6668)));
    layer4_outputs(5553) <= not((layer3_outputs(1471)) and (layer3_outputs(6294)));
    layer4_outputs(5554) <= not(layer3_outputs(6700));
    layer4_outputs(5555) <= (layer3_outputs(2876)) and (layer3_outputs(3051));
    layer4_outputs(5556) <= not(layer3_outputs(335)) or (layer3_outputs(6676));
    layer4_outputs(5557) <= not(layer3_outputs(3258)) or (layer3_outputs(4715));
    layer4_outputs(5558) <= layer3_outputs(5539);
    layer4_outputs(5559) <= not((layer3_outputs(3931)) and (layer3_outputs(821)));
    layer4_outputs(5560) <= (layer3_outputs(4446)) and (layer3_outputs(1820));
    layer4_outputs(5561) <= (layer3_outputs(2609)) and not (layer3_outputs(905));
    layer4_outputs(5562) <= layer3_outputs(4344);
    layer4_outputs(5563) <= not((layer3_outputs(5463)) and (layer3_outputs(892)));
    layer4_outputs(5564) <= not((layer3_outputs(5822)) xor (layer3_outputs(1585)));
    layer4_outputs(5565) <= not(layer3_outputs(4308)) or (layer3_outputs(4498));
    layer4_outputs(5566) <= layer3_outputs(1872);
    layer4_outputs(5567) <= not(layer3_outputs(3018));
    layer4_outputs(5568) <= not(layer3_outputs(1944));
    layer4_outputs(5569) <= '1';
    layer4_outputs(5570) <= (layer3_outputs(2394)) and not (layer3_outputs(3749));
    layer4_outputs(5571) <= layer3_outputs(1566);
    layer4_outputs(5572) <= '1';
    layer4_outputs(5573) <= not(layer3_outputs(4204));
    layer4_outputs(5574) <= (layer3_outputs(3078)) and not (layer3_outputs(3742));
    layer4_outputs(5575) <= not(layer3_outputs(4367));
    layer4_outputs(5576) <= layer3_outputs(4273);
    layer4_outputs(5577) <= (layer3_outputs(5793)) or (layer3_outputs(4789));
    layer4_outputs(5578) <= (layer3_outputs(1614)) and not (layer3_outputs(2742));
    layer4_outputs(5579) <= not((layer3_outputs(2897)) or (layer3_outputs(1546)));
    layer4_outputs(5580) <= not((layer3_outputs(5591)) and (layer3_outputs(861)));
    layer4_outputs(5581) <= not(layer3_outputs(6655)) or (layer3_outputs(3802));
    layer4_outputs(5582) <= (layer3_outputs(4403)) and not (layer3_outputs(619));
    layer4_outputs(5583) <= layer3_outputs(2555);
    layer4_outputs(5584) <= (layer3_outputs(4890)) and (layer3_outputs(1200));
    layer4_outputs(5585) <= not((layer3_outputs(1246)) or (layer3_outputs(5681)));
    layer4_outputs(5586) <= not(layer3_outputs(6144)) or (layer3_outputs(7150));
    layer4_outputs(5587) <= layer3_outputs(2756);
    layer4_outputs(5588) <= not(layer3_outputs(5570));
    layer4_outputs(5589) <= layer3_outputs(1414);
    layer4_outputs(5590) <= not((layer3_outputs(5336)) xor (layer3_outputs(1234)));
    layer4_outputs(5591) <= (layer3_outputs(6964)) and (layer3_outputs(685));
    layer4_outputs(5592) <= (layer3_outputs(336)) and not (layer3_outputs(1753));
    layer4_outputs(5593) <= layer3_outputs(3253);
    layer4_outputs(5594) <= '1';
    layer4_outputs(5595) <= (layer3_outputs(1038)) xor (layer3_outputs(534));
    layer4_outputs(5596) <= not(layer3_outputs(7550));
    layer4_outputs(5597) <= (layer3_outputs(254)) and not (layer3_outputs(6354));
    layer4_outputs(5598) <= not(layer3_outputs(1546));
    layer4_outputs(5599) <= layer3_outputs(2356);
    layer4_outputs(5600) <= not(layer3_outputs(4791));
    layer4_outputs(5601) <= '1';
    layer4_outputs(5602) <= not(layer3_outputs(6485)) or (layer3_outputs(556));
    layer4_outputs(5603) <= not((layer3_outputs(3548)) xor (layer3_outputs(7421)));
    layer4_outputs(5604) <= not((layer3_outputs(3374)) or (layer3_outputs(1229)));
    layer4_outputs(5605) <= (layer3_outputs(6846)) and not (layer3_outputs(1756));
    layer4_outputs(5606) <= not((layer3_outputs(979)) and (layer3_outputs(6123)));
    layer4_outputs(5607) <= (layer3_outputs(1231)) and not (layer3_outputs(6922));
    layer4_outputs(5608) <= (layer3_outputs(3234)) or (layer3_outputs(5652));
    layer4_outputs(5609) <= not(layer3_outputs(6042));
    layer4_outputs(5610) <= not(layer3_outputs(2916));
    layer4_outputs(5611) <= (layer3_outputs(6891)) and not (layer3_outputs(3753));
    layer4_outputs(5612) <= not(layer3_outputs(5992));
    layer4_outputs(5613) <= not(layer3_outputs(920)) or (layer3_outputs(7256));
    layer4_outputs(5614) <= not(layer3_outputs(2184)) or (layer3_outputs(6356));
    layer4_outputs(5615) <= (layer3_outputs(3015)) or (layer3_outputs(5350));
    layer4_outputs(5616) <= not(layer3_outputs(510)) or (layer3_outputs(6980));
    layer4_outputs(5617) <= '0';
    layer4_outputs(5618) <= layer3_outputs(3527);
    layer4_outputs(5619) <= layer3_outputs(6176);
    layer4_outputs(5620) <= not(layer3_outputs(4967));
    layer4_outputs(5621) <= not(layer3_outputs(6465));
    layer4_outputs(5622) <= (layer3_outputs(6548)) and not (layer3_outputs(6157));
    layer4_outputs(5623) <= not(layer3_outputs(6300));
    layer4_outputs(5624) <= (layer3_outputs(476)) and not (layer3_outputs(6520));
    layer4_outputs(5625) <= not(layer3_outputs(335)) or (layer3_outputs(7400));
    layer4_outputs(5626) <= not((layer3_outputs(431)) and (layer3_outputs(1632)));
    layer4_outputs(5627) <= (layer3_outputs(1947)) and (layer3_outputs(1415));
    layer4_outputs(5628) <= not(layer3_outputs(4342)) or (layer3_outputs(6346));
    layer4_outputs(5629) <= layer3_outputs(481);
    layer4_outputs(5630) <= (layer3_outputs(2613)) and not (layer3_outputs(3962));
    layer4_outputs(5631) <= (layer3_outputs(863)) and (layer3_outputs(1900));
    layer4_outputs(5632) <= layer3_outputs(6981);
    layer4_outputs(5633) <= not((layer3_outputs(5946)) or (layer3_outputs(2322)));
    layer4_outputs(5634) <= '0';
    layer4_outputs(5635) <= (layer3_outputs(1476)) and not (layer3_outputs(7061));
    layer4_outputs(5636) <= not(layer3_outputs(639));
    layer4_outputs(5637) <= not((layer3_outputs(4566)) or (layer3_outputs(3752)));
    layer4_outputs(5638) <= not(layer3_outputs(7566)) or (layer3_outputs(1801));
    layer4_outputs(5639) <= not(layer3_outputs(5595));
    layer4_outputs(5640) <= not(layer3_outputs(4663)) or (layer3_outputs(7447));
    layer4_outputs(5641) <= not(layer3_outputs(7650)) or (layer3_outputs(279));
    layer4_outputs(5642) <= (layer3_outputs(6920)) and (layer3_outputs(2684));
    layer4_outputs(5643) <= not(layer3_outputs(2026));
    layer4_outputs(5644) <= (layer3_outputs(1647)) xor (layer3_outputs(5331));
    layer4_outputs(5645) <= (layer3_outputs(947)) xor (layer3_outputs(3714));
    layer4_outputs(5646) <= not(layer3_outputs(1809));
    layer4_outputs(5647) <= layer3_outputs(2274);
    layer4_outputs(5648) <= not(layer3_outputs(4326)) or (layer3_outputs(1575));
    layer4_outputs(5649) <= (layer3_outputs(251)) and not (layer3_outputs(5173));
    layer4_outputs(5650) <= layer3_outputs(4231);
    layer4_outputs(5651) <= not(layer3_outputs(442));
    layer4_outputs(5652) <= not((layer3_outputs(6219)) xor (layer3_outputs(5759)));
    layer4_outputs(5653) <= not(layer3_outputs(7194)) or (layer3_outputs(5460));
    layer4_outputs(5654) <= layer3_outputs(1418);
    layer4_outputs(5655) <= '1';
    layer4_outputs(5656) <= layer3_outputs(3930);
    layer4_outputs(5657) <= layer3_outputs(800);
    layer4_outputs(5658) <= layer3_outputs(524);
    layer4_outputs(5659) <= (layer3_outputs(6237)) and (layer3_outputs(641));
    layer4_outputs(5660) <= not(layer3_outputs(2057)) or (layer3_outputs(7018));
    layer4_outputs(5661) <= not(layer3_outputs(6328));
    layer4_outputs(5662) <= not(layer3_outputs(2805));
    layer4_outputs(5663) <= layer3_outputs(6224);
    layer4_outputs(5664) <= not((layer3_outputs(159)) or (layer3_outputs(592)));
    layer4_outputs(5665) <= (layer3_outputs(7122)) or (layer3_outputs(6253));
    layer4_outputs(5666) <= (layer3_outputs(7217)) and not (layer3_outputs(5560));
    layer4_outputs(5667) <= layer3_outputs(6529);
    layer4_outputs(5668) <= '1';
    layer4_outputs(5669) <= layer3_outputs(151);
    layer4_outputs(5670) <= not((layer3_outputs(2271)) or (layer3_outputs(1935)));
    layer4_outputs(5671) <= not(layer3_outputs(1079));
    layer4_outputs(5672) <= (layer3_outputs(4521)) or (layer3_outputs(4147));
    layer4_outputs(5673) <= not((layer3_outputs(2093)) and (layer3_outputs(4367)));
    layer4_outputs(5674) <= not((layer3_outputs(1887)) or (layer3_outputs(5546)));
    layer4_outputs(5675) <= not(layer3_outputs(26));
    layer4_outputs(5676) <= (layer3_outputs(4442)) and (layer3_outputs(6886));
    layer4_outputs(5677) <= layer3_outputs(4736);
    layer4_outputs(5678) <= not((layer3_outputs(793)) and (layer3_outputs(2641)));
    layer4_outputs(5679) <= (layer3_outputs(522)) or (layer3_outputs(3789));
    layer4_outputs(5680) <= layer3_outputs(5445);
    layer4_outputs(5681) <= layer3_outputs(4338);
    layer4_outputs(5682) <= not(layer3_outputs(3346));
    layer4_outputs(5683) <= layer3_outputs(2261);
    layer4_outputs(5684) <= not(layer3_outputs(3279)) or (layer3_outputs(3115));
    layer4_outputs(5685) <= not(layer3_outputs(4818)) or (layer3_outputs(5795));
    layer4_outputs(5686) <= not(layer3_outputs(4744));
    layer4_outputs(5687) <= (layer3_outputs(246)) xor (layer3_outputs(588));
    layer4_outputs(5688) <= not(layer3_outputs(3707));
    layer4_outputs(5689) <= not(layer3_outputs(621));
    layer4_outputs(5690) <= (layer3_outputs(4594)) or (layer3_outputs(7289));
    layer4_outputs(5691) <= not(layer3_outputs(2568)) or (layer3_outputs(5678));
    layer4_outputs(5692) <= not(layer3_outputs(3251)) or (layer3_outputs(2627));
    layer4_outputs(5693) <= not((layer3_outputs(4703)) or (layer3_outputs(2126)));
    layer4_outputs(5694) <= not(layer3_outputs(4279));
    layer4_outputs(5695) <= not((layer3_outputs(7239)) or (layer3_outputs(3631)));
    layer4_outputs(5696) <= (layer3_outputs(4458)) and (layer3_outputs(2666));
    layer4_outputs(5697) <= not(layer3_outputs(5427)) or (layer3_outputs(531));
    layer4_outputs(5698) <= '0';
    layer4_outputs(5699) <= not(layer3_outputs(1687));
    layer4_outputs(5700) <= layer3_outputs(3281);
    layer4_outputs(5701) <= (layer3_outputs(2010)) and not (layer3_outputs(484));
    layer4_outputs(5702) <= layer3_outputs(5544);
    layer4_outputs(5703) <= (layer3_outputs(1894)) and not (layer3_outputs(1139));
    layer4_outputs(5704) <= not(layer3_outputs(2991)) or (layer3_outputs(4619));
    layer4_outputs(5705) <= (layer3_outputs(6026)) and (layer3_outputs(1099));
    layer4_outputs(5706) <= (layer3_outputs(13)) and not (layer3_outputs(4778));
    layer4_outputs(5707) <= not(layer3_outputs(5586)) or (layer3_outputs(3746));
    layer4_outputs(5708) <= layer3_outputs(4334);
    layer4_outputs(5709) <= (layer3_outputs(4308)) xor (layer3_outputs(3169));
    layer4_outputs(5710) <= (layer3_outputs(6744)) and (layer3_outputs(1974));
    layer4_outputs(5711) <= not(layer3_outputs(3028));
    layer4_outputs(5712) <= not(layer3_outputs(185));
    layer4_outputs(5713) <= layer3_outputs(6233);
    layer4_outputs(5714) <= (layer3_outputs(2688)) and not (layer3_outputs(1105));
    layer4_outputs(5715) <= (layer3_outputs(352)) and (layer3_outputs(5914));
    layer4_outputs(5716) <= not(layer3_outputs(1696));
    layer4_outputs(5717) <= not((layer3_outputs(572)) or (layer3_outputs(608)));
    layer4_outputs(5718) <= layer3_outputs(7297);
    layer4_outputs(5719) <= (layer3_outputs(3421)) xor (layer3_outputs(2568));
    layer4_outputs(5720) <= not(layer3_outputs(6534)) or (layer3_outputs(6989));
    layer4_outputs(5721) <= not((layer3_outputs(2791)) and (layer3_outputs(3888)));
    layer4_outputs(5722) <= layer3_outputs(1946);
    layer4_outputs(5723) <= layer3_outputs(7095);
    layer4_outputs(5724) <= (layer3_outputs(2062)) and not (layer3_outputs(7128));
    layer4_outputs(5725) <= layer3_outputs(5520);
    layer4_outputs(5726) <= (layer3_outputs(539)) and not (layer3_outputs(1237));
    layer4_outputs(5727) <= not((layer3_outputs(2361)) and (layer3_outputs(4917)));
    layer4_outputs(5728) <= (layer3_outputs(7559)) and not (layer3_outputs(7479));
    layer4_outputs(5729) <= not(layer3_outputs(1408));
    layer4_outputs(5730) <= not((layer3_outputs(4342)) xor (layer3_outputs(311)));
    layer4_outputs(5731) <= (layer3_outputs(1020)) and not (layer3_outputs(1989));
    layer4_outputs(5732) <= layer3_outputs(2050);
    layer4_outputs(5733) <= not(layer3_outputs(6861));
    layer4_outputs(5734) <= not(layer3_outputs(7002));
    layer4_outputs(5735) <= not(layer3_outputs(3244));
    layer4_outputs(5736) <= not(layer3_outputs(1706));
    layer4_outputs(5737) <= not(layer3_outputs(4398)) or (layer3_outputs(5910));
    layer4_outputs(5738) <= (layer3_outputs(5447)) and (layer3_outputs(4749));
    layer4_outputs(5739) <= (layer3_outputs(3690)) or (layer3_outputs(268));
    layer4_outputs(5740) <= (layer3_outputs(4977)) and not (layer3_outputs(1252));
    layer4_outputs(5741) <= not(layer3_outputs(1978)) or (layer3_outputs(642));
    layer4_outputs(5742) <= layer3_outputs(7190);
    layer4_outputs(5743) <= not((layer3_outputs(915)) and (layer3_outputs(4104)));
    layer4_outputs(5744) <= not((layer3_outputs(3158)) or (layer3_outputs(5070)));
    layer4_outputs(5745) <= layer3_outputs(5723);
    layer4_outputs(5746) <= not(layer3_outputs(5769));
    layer4_outputs(5747) <= not(layer3_outputs(1231));
    layer4_outputs(5748) <= (layer3_outputs(4714)) and not (layer3_outputs(7027));
    layer4_outputs(5749) <= not(layer3_outputs(3374));
    layer4_outputs(5750) <= (layer3_outputs(2946)) or (layer3_outputs(5912));
    layer4_outputs(5751) <= not(layer3_outputs(1734)) or (layer3_outputs(2215));
    layer4_outputs(5752) <= (layer3_outputs(6506)) xor (layer3_outputs(1694));
    layer4_outputs(5753) <= not((layer3_outputs(1619)) and (layer3_outputs(582)));
    layer4_outputs(5754) <= (layer3_outputs(1638)) and not (layer3_outputs(5853));
    layer4_outputs(5755) <= not((layer3_outputs(7011)) or (layer3_outputs(4151)));
    layer4_outputs(5756) <= not(layer3_outputs(3828));
    layer4_outputs(5757) <= (layer3_outputs(3373)) and (layer3_outputs(5626));
    layer4_outputs(5758) <= not((layer3_outputs(1424)) and (layer3_outputs(301)));
    layer4_outputs(5759) <= not((layer3_outputs(6929)) or (layer3_outputs(6399)));
    layer4_outputs(5760) <= not(layer3_outputs(2182));
    layer4_outputs(5761) <= layer3_outputs(7015);
    layer4_outputs(5762) <= not(layer3_outputs(3010)) or (layer3_outputs(3609));
    layer4_outputs(5763) <= layer3_outputs(627);
    layer4_outputs(5764) <= not(layer3_outputs(5083));
    layer4_outputs(5765) <= (layer3_outputs(5995)) xor (layer3_outputs(754));
    layer4_outputs(5766) <= (layer3_outputs(7032)) and (layer3_outputs(2977));
    layer4_outputs(5767) <= not((layer3_outputs(1967)) and (layer3_outputs(3309)));
    layer4_outputs(5768) <= layer3_outputs(2819);
    layer4_outputs(5769) <= layer3_outputs(3554);
    layer4_outputs(5770) <= '0';
    layer4_outputs(5771) <= not((layer3_outputs(2236)) and (layer3_outputs(6093)));
    layer4_outputs(5772) <= layer3_outputs(2225);
    layer4_outputs(5773) <= not((layer3_outputs(1520)) and (layer3_outputs(6934)));
    layer4_outputs(5774) <= (layer3_outputs(2469)) and not (layer3_outputs(5366));
    layer4_outputs(5775) <= (layer3_outputs(5604)) and not (layer3_outputs(501));
    layer4_outputs(5776) <= layer3_outputs(786);
    layer4_outputs(5777) <= '1';
    layer4_outputs(5778) <= (layer3_outputs(5380)) and not (layer3_outputs(3763));
    layer4_outputs(5779) <= not(layer3_outputs(1094)) or (layer3_outputs(3758));
    layer4_outputs(5780) <= (layer3_outputs(540)) or (layer3_outputs(2697));
    layer4_outputs(5781) <= (layer3_outputs(6497)) xor (layer3_outputs(1483));
    layer4_outputs(5782) <= (layer3_outputs(3159)) xor (layer3_outputs(4470));
    layer4_outputs(5783) <= not(layer3_outputs(5297)) or (layer3_outputs(1724));
    layer4_outputs(5784) <= '1';
    layer4_outputs(5785) <= not((layer3_outputs(474)) xor (layer3_outputs(3629)));
    layer4_outputs(5786) <= not(layer3_outputs(5371)) or (layer3_outputs(5742));
    layer4_outputs(5787) <= (layer3_outputs(4756)) or (layer3_outputs(832));
    layer4_outputs(5788) <= not((layer3_outputs(514)) or (layer3_outputs(7650)));
    layer4_outputs(5789) <= not(layer3_outputs(4621));
    layer4_outputs(5790) <= not(layer3_outputs(1773));
    layer4_outputs(5791) <= layer3_outputs(5735);
    layer4_outputs(5792) <= (layer3_outputs(1118)) and not (layer3_outputs(4295));
    layer4_outputs(5793) <= not(layer3_outputs(6165)) or (layer3_outputs(2948));
    layer4_outputs(5794) <= (layer3_outputs(3440)) and not (layer3_outputs(118));
    layer4_outputs(5795) <= not(layer3_outputs(1610));
    layer4_outputs(5796) <= (layer3_outputs(1517)) or (layer3_outputs(6090));
    layer4_outputs(5797) <= (layer3_outputs(6792)) xor (layer3_outputs(4712));
    layer4_outputs(5798) <= not(layer3_outputs(3190)) or (layer3_outputs(5618));
    layer4_outputs(5799) <= '1';
    layer4_outputs(5800) <= not(layer3_outputs(1846));
    layer4_outputs(5801) <= layer3_outputs(4612);
    layer4_outputs(5802) <= layer3_outputs(67);
    layer4_outputs(5803) <= not(layer3_outputs(5421)) or (layer3_outputs(6591));
    layer4_outputs(5804) <= (layer3_outputs(2460)) and not (layer3_outputs(2178));
    layer4_outputs(5805) <= not((layer3_outputs(3406)) or (layer3_outputs(313)));
    layer4_outputs(5806) <= not((layer3_outputs(6769)) and (layer3_outputs(2599)));
    layer4_outputs(5807) <= not(layer3_outputs(7375));
    layer4_outputs(5808) <= not(layer3_outputs(2895));
    layer4_outputs(5809) <= '0';
    layer4_outputs(5810) <= not((layer3_outputs(5102)) xor (layer3_outputs(5599)));
    layer4_outputs(5811) <= layer3_outputs(108);
    layer4_outputs(5812) <= layer3_outputs(6571);
    layer4_outputs(5813) <= not(layer3_outputs(5435));
    layer4_outputs(5814) <= not(layer3_outputs(1496));
    layer4_outputs(5815) <= (layer3_outputs(6257)) and not (layer3_outputs(6767));
    layer4_outputs(5816) <= layer3_outputs(5351);
    layer4_outputs(5817) <= not(layer3_outputs(7212)) or (layer3_outputs(3948));
    layer4_outputs(5818) <= (layer3_outputs(7031)) or (layer3_outputs(242));
    layer4_outputs(5819) <= layer3_outputs(4066);
    layer4_outputs(5820) <= layer3_outputs(3320);
    layer4_outputs(5821) <= layer3_outputs(3434);
    layer4_outputs(5822) <= not(layer3_outputs(4386)) or (layer3_outputs(1717));
    layer4_outputs(5823) <= (layer3_outputs(6740)) and (layer3_outputs(5419));
    layer4_outputs(5824) <= not(layer3_outputs(2783));
    layer4_outputs(5825) <= '1';
    layer4_outputs(5826) <= not(layer3_outputs(4541));
    layer4_outputs(5827) <= layer3_outputs(7384);
    layer4_outputs(5828) <= layer3_outputs(2242);
    layer4_outputs(5829) <= (layer3_outputs(7257)) and (layer3_outputs(6608));
    layer4_outputs(5830) <= not(layer3_outputs(6012));
    layer4_outputs(5831) <= layer3_outputs(239);
    layer4_outputs(5832) <= not(layer3_outputs(3603)) or (layer3_outputs(4150));
    layer4_outputs(5833) <= not(layer3_outputs(7118));
    layer4_outputs(5834) <= not(layer3_outputs(5516));
    layer4_outputs(5835) <= (layer3_outputs(4758)) or (layer3_outputs(2565));
    layer4_outputs(5836) <= not(layer3_outputs(1105));
    layer4_outputs(5837) <= not((layer3_outputs(2907)) and (layer3_outputs(4300)));
    layer4_outputs(5838) <= (layer3_outputs(3452)) and (layer3_outputs(5101));
    layer4_outputs(5839) <= layer3_outputs(3816);
    layer4_outputs(5840) <= layer3_outputs(1955);
    layer4_outputs(5841) <= layer3_outputs(7515);
    layer4_outputs(5842) <= (layer3_outputs(4444)) and not (layer3_outputs(7535));
    layer4_outputs(5843) <= not((layer3_outputs(2776)) and (layer3_outputs(6570)));
    layer4_outputs(5844) <= not(layer3_outputs(3569)) or (layer3_outputs(5394));
    layer4_outputs(5845) <= layer3_outputs(5494);
    layer4_outputs(5846) <= not(layer3_outputs(3234));
    layer4_outputs(5847) <= not((layer3_outputs(1244)) xor (layer3_outputs(7596)));
    layer4_outputs(5848) <= layer3_outputs(2706);
    layer4_outputs(5849) <= layer3_outputs(374);
    layer4_outputs(5850) <= (layer3_outputs(5219)) or (layer3_outputs(4362));
    layer4_outputs(5851) <= not(layer3_outputs(5101)) or (layer3_outputs(701));
    layer4_outputs(5852) <= layer3_outputs(5968);
    layer4_outputs(5853) <= '0';
    layer4_outputs(5854) <= layer3_outputs(752);
    layer4_outputs(5855) <= '1';
    layer4_outputs(5856) <= (layer3_outputs(5185)) xor (layer3_outputs(1500));
    layer4_outputs(5857) <= not(layer3_outputs(7384));
    layer4_outputs(5858) <= '1';
    layer4_outputs(5859) <= '0';
    layer4_outputs(5860) <= layer3_outputs(5596);
    layer4_outputs(5861) <= not(layer3_outputs(7191));
    layer4_outputs(5862) <= not(layer3_outputs(589));
    layer4_outputs(5863) <= not(layer3_outputs(2348));
    layer4_outputs(5864) <= not((layer3_outputs(6502)) and (layer3_outputs(3073)));
    layer4_outputs(5865) <= layer3_outputs(5538);
    layer4_outputs(5866) <= '1';
    layer4_outputs(5867) <= not((layer3_outputs(4916)) xor (layer3_outputs(7317)));
    layer4_outputs(5868) <= not(layer3_outputs(1562));
    layer4_outputs(5869) <= (layer3_outputs(6785)) and not (layer3_outputs(6441));
    layer4_outputs(5870) <= not(layer3_outputs(6013));
    layer4_outputs(5871) <= not(layer3_outputs(2837));
    layer4_outputs(5872) <= (layer3_outputs(3934)) or (layer3_outputs(843));
    layer4_outputs(5873) <= not(layer3_outputs(5031));
    layer4_outputs(5874) <= not(layer3_outputs(1035)) or (layer3_outputs(2051));
    layer4_outputs(5875) <= (layer3_outputs(172)) and not (layer3_outputs(5418));
    layer4_outputs(5876) <= not(layer3_outputs(6446)) or (layer3_outputs(7263));
    layer4_outputs(5877) <= layer3_outputs(1430);
    layer4_outputs(5878) <= not(layer3_outputs(1709)) or (layer3_outputs(3558));
    layer4_outputs(5879) <= layer3_outputs(3141);
    layer4_outputs(5880) <= layer3_outputs(6797);
    layer4_outputs(5881) <= '1';
    layer4_outputs(5882) <= not((layer3_outputs(7386)) and (layer3_outputs(3477)));
    layer4_outputs(5883) <= layer3_outputs(3069);
    layer4_outputs(5884) <= not(layer3_outputs(185));
    layer4_outputs(5885) <= '1';
    layer4_outputs(5886) <= layer3_outputs(3514);
    layer4_outputs(5887) <= (layer3_outputs(2333)) or (layer3_outputs(5718));
    layer4_outputs(5888) <= (layer3_outputs(5050)) and (layer3_outputs(1044));
    layer4_outputs(5889) <= not(layer3_outputs(6194)) or (layer3_outputs(3262));
    layer4_outputs(5890) <= not(layer3_outputs(7560)) or (layer3_outputs(1768));
    layer4_outputs(5891) <= not(layer3_outputs(4106));
    layer4_outputs(5892) <= not(layer3_outputs(2394)) or (layer3_outputs(7619));
    layer4_outputs(5893) <= not(layer3_outputs(4048)) or (layer3_outputs(2134));
    layer4_outputs(5894) <= '1';
    layer4_outputs(5895) <= not((layer3_outputs(6426)) xor (layer3_outputs(3473)));
    layer4_outputs(5896) <= not((layer3_outputs(1784)) xor (layer3_outputs(7460)));
    layer4_outputs(5897) <= layer3_outputs(7634);
    layer4_outputs(5898) <= not((layer3_outputs(1998)) or (layer3_outputs(4440)));
    layer4_outputs(5899) <= not(layer3_outputs(7651));
    layer4_outputs(5900) <= not((layer3_outputs(2855)) and (layer3_outputs(3920)));
    layer4_outputs(5901) <= layer3_outputs(987);
    layer4_outputs(5902) <= not(layer3_outputs(2432));
    layer4_outputs(5903) <= not(layer3_outputs(5948));
    layer4_outputs(5904) <= (layer3_outputs(1859)) xor (layer3_outputs(5878));
    layer4_outputs(5905) <= layer3_outputs(4470);
    layer4_outputs(5906) <= layer3_outputs(611);
    layer4_outputs(5907) <= (layer3_outputs(1268)) and (layer3_outputs(54));
    layer4_outputs(5908) <= not(layer3_outputs(3613));
    layer4_outputs(5909) <= '1';
    layer4_outputs(5910) <= layer3_outputs(4330);
    layer4_outputs(5911) <= not((layer3_outputs(4720)) xor (layer3_outputs(5573)));
    layer4_outputs(5912) <= layer3_outputs(4956);
    layer4_outputs(5913) <= '1';
    layer4_outputs(5914) <= not((layer3_outputs(953)) and (layer3_outputs(2611)));
    layer4_outputs(5915) <= not(layer3_outputs(4876));
    layer4_outputs(5916) <= not(layer3_outputs(2838)) or (layer3_outputs(6194));
    layer4_outputs(5917) <= not((layer3_outputs(565)) and (layer3_outputs(754)));
    layer4_outputs(5918) <= layer3_outputs(7088);
    layer4_outputs(5919) <= not((layer3_outputs(5344)) and (layer3_outputs(3048)));
    layer4_outputs(5920) <= '0';
    layer4_outputs(5921) <= (layer3_outputs(6586)) xor (layer3_outputs(6325));
    layer4_outputs(5922) <= layer3_outputs(6195);
    layer4_outputs(5923) <= '1';
    layer4_outputs(5924) <= not(layer3_outputs(1205)) or (layer3_outputs(3877));
    layer4_outputs(5925) <= '0';
    layer4_outputs(5926) <= layer3_outputs(6897);
    layer4_outputs(5927) <= not(layer3_outputs(4195));
    layer4_outputs(5928) <= not(layer3_outputs(3905)) or (layer3_outputs(186));
    layer4_outputs(5929) <= not(layer3_outputs(5632)) or (layer3_outputs(4069));
    layer4_outputs(5930) <= not(layer3_outputs(2989));
    layer4_outputs(5931) <= not((layer3_outputs(2108)) or (layer3_outputs(7119)));
    layer4_outputs(5932) <= (layer3_outputs(3718)) and not (layer3_outputs(4478));
    layer4_outputs(5933) <= not(layer3_outputs(4495));
    layer4_outputs(5934) <= '0';
    layer4_outputs(5935) <= layer3_outputs(3161);
    layer4_outputs(5936) <= (layer3_outputs(4467)) and not (layer3_outputs(1366));
    layer4_outputs(5937) <= not(layer3_outputs(587));
    layer4_outputs(5938) <= not(layer3_outputs(1513));
    layer4_outputs(5939) <= not(layer3_outputs(5890));
    layer4_outputs(5940) <= not(layer3_outputs(713));
    layer4_outputs(5941) <= (layer3_outputs(1260)) and not (layer3_outputs(434));
    layer4_outputs(5942) <= '0';
    layer4_outputs(5943) <= (layer3_outputs(6263)) and not (layer3_outputs(6722));
    layer4_outputs(5944) <= not(layer3_outputs(4406));
    layer4_outputs(5945) <= not(layer3_outputs(825)) or (layer3_outputs(6893));
    layer4_outputs(5946) <= not(layer3_outputs(3045));
    layer4_outputs(5947) <= not((layer3_outputs(2741)) or (layer3_outputs(3794)));
    layer4_outputs(5948) <= (layer3_outputs(5317)) and not (layer3_outputs(314));
    layer4_outputs(5949) <= not((layer3_outputs(1653)) or (layer3_outputs(94)));
    layer4_outputs(5950) <= layer3_outputs(7586);
    layer4_outputs(5951) <= not((layer3_outputs(1848)) and (layer3_outputs(7636)));
    layer4_outputs(5952) <= (layer3_outputs(5051)) or (layer3_outputs(2595));
    layer4_outputs(5953) <= not(layer3_outputs(6157));
    layer4_outputs(5954) <= not((layer3_outputs(4373)) xor (layer3_outputs(4211)));
    layer4_outputs(5955) <= (layer3_outputs(2838)) and (layer3_outputs(2477));
    layer4_outputs(5956) <= not(layer3_outputs(1473)) or (layer3_outputs(7039));
    layer4_outputs(5957) <= (layer3_outputs(4991)) and not (layer3_outputs(3814));
    layer4_outputs(5958) <= not(layer3_outputs(7095));
    layer4_outputs(5959) <= not((layer3_outputs(7616)) or (layer3_outputs(1380)));
    layer4_outputs(5960) <= not(layer3_outputs(4004)) or (layer3_outputs(4820));
    layer4_outputs(5961) <= layer3_outputs(19);
    layer4_outputs(5962) <= not(layer3_outputs(4475)) or (layer3_outputs(6943));
    layer4_outputs(5963) <= layer3_outputs(3384);
    layer4_outputs(5964) <= (layer3_outputs(6910)) and not (layer3_outputs(7582));
    layer4_outputs(5965) <= not(layer3_outputs(5544));
    layer4_outputs(5966) <= not((layer3_outputs(6259)) xor (layer3_outputs(4625)));
    layer4_outputs(5967) <= layer3_outputs(2203);
    layer4_outputs(5968) <= (layer3_outputs(1356)) or (layer3_outputs(5422));
    layer4_outputs(5969) <= not((layer3_outputs(2475)) and (layer3_outputs(1341)));
    layer4_outputs(5970) <= not(layer3_outputs(4679)) or (layer3_outputs(7388));
    layer4_outputs(5971) <= (layer3_outputs(5150)) and not (layer3_outputs(5883));
    layer4_outputs(5972) <= not(layer3_outputs(3273)) or (layer3_outputs(485));
    layer4_outputs(5973) <= not((layer3_outputs(5771)) or (layer3_outputs(560)));
    layer4_outputs(5974) <= not(layer3_outputs(1714)) or (layer3_outputs(1803));
    layer4_outputs(5975) <= layer3_outputs(3338);
    layer4_outputs(5976) <= not((layer3_outputs(70)) or (layer3_outputs(2712)));
    layer4_outputs(5977) <= not((layer3_outputs(3998)) or (layer3_outputs(7141)));
    layer4_outputs(5978) <= not(layer3_outputs(7254)) or (layer3_outputs(7436));
    layer4_outputs(5979) <= not(layer3_outputs(4056));
    layer4_outputs(5980) <= not(layer3_outputs(6850));
    layer4_outputs(5981) <= layer3_outputs(5968);
    layer4_outputs(5982) <= (layer3_outputs(6199)) and not (layer3_outputs(7486));
    layer4_outputs(5983) <= not(layer3_outputs(5779));
    layer4_outputs(5984) <= not(layer3_outputs(7054));
    layer4_outputs(5985) <= not(layer3_outputs(4407));
    layer4_outputs(5986) <= not(layer3_outputs(156));
    layer4_outputs(5987) <= layer3_outputs(2673);
    layer4_outputs(5988) <= not((layer3_outputs(5580)) and (layer3_outputs(494)));
    layer4_outputs(5989) <= '0';
    layer4_outputs(5990) <= '0';
    layer4_outputs(5991) <= not(layer3_outputs(6081));
    layer4_outputs(5992) <= not(layer3_outputs(4008));
    layer4_outputs(5993) <= not((layer3_outputs(3722)) xor (layer3_outputs(4733)));
    layer4_outputs(5994) <= layer3_outputs(3407);
    layer4_outputs(5995) <= layer3_outputs(5030);
    layer4_outputs(5996) <= not(layer3_outputs(1090));
    layer4_outputs(5997) <= layer3_outputs(6798);
    layer4_outputs(5998) <= not((layer3_outputs(7126)) or (layer3_outputs(6912)));
    layer4_outputs(5999) <= not(layer3_outputs(794));
    layer4_outputs(6000) <= not(layer3_outputs(5909)) or (layer3_outputs(6647));
    layer4_outputs(6001) <= layer3_outputs(6050);
    layer4_outputs(6002) <= layer3_outputs(3207);
    layer4_outputs(6003) <= (layer3_outputs(3625)) or (layer3_outputs(273));
    layer4_outputs(6004) <= (layer3_outputs(6160)) and not (layer3_outputs(2127));
    layer4_outputs(6005) <= not((layer3_outputs(6680)) and (layer3_outputs(5309)));
    layer4_outputs(6006) <= not(layer3_outputs(5799));
    layer4_outputs(6007) <= (layer3_outputs(6468)) and (layer3_outputs(4848));
    layer4_outputs(6008) <= (layer3_outputs(5226)) and not (layer3_outputs(5142));
    layer4_outputs(6009) <= not((layer3_outputs(5164)) xor (layer3_outputs(2178)));
    layer4_outputs(6010) <= not(layer3_outputs(7192)) or (layer3_outputs(6853));
    layer4_outputs(6011) <= (layer3_outputs(6068)) and not (layer3_outputs(4027));
    layer4_outputs(6012) <= not((layer3_outputs(2149)) and (layer3_outputs(7622)));
    layer4_outputs(6013) <= (layer3_outputs(6207)) xor (layer3_outputs(4481));
    layer4_outputs(6014) <= (layer3_outputs(5071)) and (layer3_outputs(3575));
    layer4_outputs(6015) <= (layer3_outputs(202)) xor (layer3_outputs(3910));
    layer4_outputs(6016) <= not(layer3_outputs(1608)) or (layer3_outputs(7584));
    layer4_outputs(6017) <= '0';
    layer4_outputs(6018) <= not(layer3_outputs(5508));
    layer4_outputs(6019) <= layer3_outputs(1062);
    layer4_outputs(6020) <= not(layer3_outputs(2170)) or (layer3_outputs(2741));
    layer4_outputs(6021) <= '0';
    layer4_outputs(6022) <= not(layer3_outputs(1151));
    layer4_outputs(6023) <= (layer3_outputs(4329)) and (layer3_outputs(2932));
    layer4_outputs(6024) <= not((layer3_outputs(6249)) and (layer3_outputs(3957)));
    layer4_outputs(6025) <= '0';
    layer4_outputs(6026) <= not((layer3_outputs(2110)) or (layer3_outputs(6306)));
    layer4_outputs(6027) <= not(layer3_outputs(6701)) or (layer3_outputs(602));
    layer4_outputs(6028) <= '0';
    layer4_outputs(6029) <= not(layer3_outputs(540)) or (layer3_outputs(2452));
    layer4_outputs(6030) <= not(layer3_outputs(783)) or (layer3_outputs(6712));
    layer4_outputs(6031) <= not((layer3_outputs(2144)) and (layer3_outputs(244)));
    layer4_outputs(6032) <= layer3_outputs(2043);
    layer4_outputs(6033) <= (layer3_outputs(4792)) and (layer3_outputs(4272));
    layer4_outputs(6034) <= (layer3_outputs(4757)) and not (layer3_outputs(2894));
    layer4_outputs(6035) <= layer3_outputs(4702);
    layer4_outputs(6036) <= not(layer3_outputs(2263)) or (layer3_outputs(5280));
    layer4_outputs(6037) <= not(layer3_outputs(2391)) or (layer3_outputs(1658));
    layer4_outputs(6038) <= (layer3_outputs(4754)) and (layer3_outputs(6204));
    layer4_outputs(6039) <= (layer3_outputs(3404)) or (layer3_outputs(3845));
    layer4_outputs(6040) <= not((layer3_outputs(6774)) or (layer3_outputs(1226)));
    layer4_outputs(6041) <= layer3_outputs(218);
    layer4_outputs(6042) <= (layer3_outputs(6764)) and not (layer3_outputs(1051));
    layer4_outputs(6043) <= not(layer3_outputs(1602));
    layer4_outputs(6044) <= (layer3_outputs(2941)) and not (layer3_outputs(6991));
    layer4_outputs(6045) <= not((layer3_outputs(6779)) or (layer3_outputs(2968)));
    layer4_outputs(6046) <= (layer3_outputs(4621)) and (layer3_outputs(3995));
    layer4_outputs(6047) <= not(layer3_outputs(3618));
    layer4_outputs(6048) <= layer3_outputs(194);
    layer4_outputs(6049) <= not(layer3_outputs(1379)) or (layer3_outputs(2112));
    layer4_outputs(6050) <= not(layer3_outputs(4871));
    layer4_outputs(6051) <= not((layer3_outputs(7268)) and (layer3_outputs(2385)));
    layer4_outputs(6052) <= not((layer3_outputs(839)) and (layer3_outputs(7240)));
    layer4_outputs(6053) <= not(layer3_outputs(4306));
    layer4_outputs(6054) <= layer3_outputs(2662);
    layer4_outputs(6055) <= not(layer3_outputs(7524));
    layer4_outputs(6056) <= layer3_outputs(5629);
    layer4_outputs(6057) <= (layer3_outputs(4959)) or (layer3_outputs(7665));
    layer4_outputs(6058) <= (layer3_outputs(2146)) and not (layer3_outputs(962));
    layer4_outputs(6059) <= not(layer3_outputs(3632));
    layer4_outputs(6060) <= not(layer3_outputs(5572));
    layer4_outputs(6061) <= layer3_outputs(1628);
    layer4_outputs(6062) <= '1';
    layer4_outputs(6063) <= (layer3_outputs(2910)) and not (layer3_outputs(4415));
    layer4_outputs(6064) <= layer3_outputs(3669);
    layer4_outputs(6065) <= not(layer3_outputs(4469));
    layer4_outputs(6066) <= not(layer3_outputs(1938)) or (layer3_outputs(5123));
    layer4_outputs(6067) <= '0';
    layer4_outputs(6068) <= not((layer3_outputs(5081)) and (layer3_outputs(5345)));
    layer4_outputs(6069) <= '0';
    layer4_outputs(6070) <= (layer3_outputs(5880)) and not (layer3_outputs(4904));
    layer4_outputs(6071) <= not((layer3_outputs(232)) xor (layer3_outputs(2554)));
    layer4_outputs(6072) <= not(layer3_outputs(1722));
    layer4_outputs(6073) <= not(layer3_outputs(292));
    layer4_outputs(6074) <= not(layer3_outputs(5132)) or (layer3_outputs(6290));
    layer4_outputs(6075) <= (layer3_outputs(7379)) or (layer3_outputs(2196));
    layer4_outputs(6076) <= not(layer3_outputs(1101));
    layer4_outputs(6077) <= not(layer3_outputs(511)) or (layer3_outputs(865));
    layer4_outputs(6078) <= (layer3_outputs(4401)) and (layer3_outputs(706));
    layer4_outputs(6079) <= not(layer3_outputs(1700)) or (layer3_outputs(4209));
    layer4_outputs(6080) <= not(layer3_outputs(7459));
    layer4_outputs(6081) <= not((layer3_outputs(907)) or (layer3_outputs(230)));
    layer4_outputs(6082) <= layer3_outputs(7178);
    layer4_outputs(6083) <= layer3_outputs(5551);
    layer4_outputs(6084) <= not(layer3_outputs(1906));
    layer4_outputs(6085) <= layer3_outputs(768);
    layer4_outputs(6086) <= not(layer3_outputs(2424));
    layer4_outputs(6087) <= (layer3_outputs(2980)) and not (layer3_outputs(1450));
    layer4_outputs(6088) <= not(layer3_outputs(119)) or (layer3_outputs(4590));
    layer4_outputs(6089) <= layer3_outputs(5802);
    layer4_outputs(6090) <= (layer3_outputs(6986)) and (layer3_outputs(2429));
    layer4_outputs(6091) <= not(layer3_outputs(1767));
    layer4_outputs(6092) <= layer3_outputs(3402);
    layer4_outputs(6093) <= (layer3_outputs(843)) xor (layer3_outputs(1738));
    layer4_outputs(6094) <= (layer3_outputs(1528)) and not (layer3_outputs(5808));
    layer4_outputs(6095) <= not(layer3_outputs(632));
    layer4_outputs(6096) <= layer3_outputs(539);
    layer4_outputs(6097) <= layer3_outputs(5788);
    layer4_outputs(6098) <= not((layer3_outputs(5208)) xor (layer3_outputs(5449)));
    layer4_outputs(6099) <= layer3_outputs(7401);
    layer4_outputs(6100) <= layer3_outputs(3516);
    layer4_outputs(6101) <= not(layer3_outputs(4797));
    layer4_outputs(6102) <= not((layer3_outputs(4917)) or (layer3_outputs(850)));
    layer4_outputs(6103) <= '0';
    layer4_outputs(6104) <= layer3_outputs(2443);
    layer4_outputs(6105) <= (layer3_outputs(5143)) and not (layer3_outputs(5189));
    layer4_outputs(6106) <= (layer3_outputs(3894)) and (layer3_outputs(4509));
    layer4_outputs(6107) <= '1';
    layer4_outputs(6108) <= not((layer3_outputs(5705)) xor (layer3_outputs(3689)));
    layer4_outputs(6109) <= (layer3_outputs(1960)) and (layer3_outputs(5304));
    layer4_outputs(6110) <= not((layer3_outputs(5134)) or (layer3_outputs(3748)));
    layer4_outputs(6111) <= (layer3_outputs(4343)) and (layer3_outputs(6635));
    layer4_outputs(6112) <= (layer3_outputs(635)) and not (layer3_outputs(727));
    layer4_outputs(6113) <= (layer3_outputs(3371)) and not (layer3_outputs(5223));
    layer4_outputs(6114) <= not((layer3_outputs(5282)) and (layer3_outputs(5858)));
    layer4_outputs(6115) <= not(layer3_outputs(2471));
    layer4_outputs(6116) <= not((layer3_outputs(3892)) and (layer3_outputs(2681)));
    layer4_outputs(6117) <= layer3_outputs(3840);
    layer4_outputs(6118) <= (layer3_outputs(662)) or (layer3_outputs(871));
    layer4_outputs(6119) <= (layer3_outputs(1606)) and not (layer3_outputs(4429));
    layer4_outputs(6120) <= not(layer3_outputs(3082));
    layer4_outputs(6121) <= not(layer3_outputs(3929));
    layer4_outputs(6122) <= not((layer3_outputs(1775)) xor (layer3_outputs(6272)));
    layer4_outputs(6123) <= not((layer3_outputs(1603)) xor (layer3_outputs(7527)));
    layer4_outputs(6124) <= not((layer3_outputs(460)) and (layer3_outputs(824)));
    layer4_outputs(6125) <= (layer3_outputs(4488)) and not (layer3_outputs(526));
    layer4_outputs(6126) <= not(layer3_outputs(2079));
    layer4_outputs(6127) <= not((layer3_outputs(3896)) and (layer3_outputs(538)));
    layer4_outputs(6128) <= layer3_outputs(1844);
    layer4_outputs(6129) <= (layer3_outputs(6766)) and (layer3_outputs(3319));
    layer4_outputs(6130) <= layer3_outputs(6391);
    layer4_outputs(6131) <= layer3_outputs(4802);
    layer4_outputs(6132) <= layer3_outputs(6735);
    layer4_outputs(6133) <= layer3_outputs(4801);
    layer4_outputs(6134) <= layer3_outputs(3934);
    layer4_outputs(6135) <= not(layer3_outputs(2145));
    layer4_outputs(6136) <= not((layer3_outputs(3553)) and (layer3_outputs(7437)));
    layer4_outputs(6137) <= not(layer3_outputs(1901));
    layer4_outputs(6138) <= '1';
    layer4_outputs(6139) <= not(layer3_outputs(2510));
    layer4_outputs(6140) <= (layer3_outputs(1327)) xor (layer3_outputs(4388));
    layer4_outputs(6141) <= not(layer3_outputs(1921));
    layer4_outputs(6142) <= (layer3_outputs(1403)) and not (layer3_outputs(4134));
    layer4_outputs(6143) <= (layer3_outputs(4260)) and (layer3_outputs(3043));
    layer4_outputs(6144) <= (layer3_outputs(6525)) or (layer3_outputs(1844));
    layer4_outputs(6145) <= not(layer3_outputs(7263));
    layer4_outputs(6146) <= not(layer3_outputs(5769));
    layer4_outputs(6147) <= (layer3_outputs(6606)) and not (layer3_outputs(1398));
    layer4_outputs(6148) <= '1';
    layer4_outputs(6149) <= (layer3_outputs(6579)) and not (layer3_outputs(6507));
    layer4_outputs(6150) <= (layer3_outputs(2111)) and not (layer3_outputs(2668));
    layer4_outputs(6151) <= (layer3_outputs(2856)) or (layer3_outputs(7536));
    layer4_outputs(6152) <= (layer3_outputs(4377)) and not (layer3_outputs(6329));
    layer4_outputs(6153) <= not(layer3_outputs(6977));
    layer4_outputs(6154) <= not(layer3_outputs(2191));
    layer4_outputs(6155) <= '0';
    layer4_outputs(6156) <= not((layer3_outputs(7)) and (layer3_outputs(4160)));
    layer4_outputs(6157) <= layer3_outputs(6229);
    layer4_outputs(6158) <= '0';
    layer4_outputs(6159) <= not(layer3_outputs(4599));
    layer4_outputs(6160) <= not(layer3_outputs(3764));
    layer4_outputs(6161) <= not(layer3_outputs(4430)) or (layer3_outputs(4213));
    layer4_outputs(6162) <= not(layer3_outputs(2999));
    layer4_outputs(6163) <= (layer3_outputs(1041)) and not (layer3_outputs(200));
    layer4_outputs(6164) <= not((layer3_outputs(3582)) or (layer3_outputs(6269)));
    layer4_outputs(6165) <= '0';
    layer4_outputs(6166) <= not(layer3_outputs(5468));
    layer4_outputs(6167) <= not(layer3_outputs(5808)) or (layer3_outputs(5354));
    layer4_outputs(6168) <= (layer3_outputs(5194)) and not (layer3_outputs(396));
    layer4_outputs(6169) <= layer3_outputs(5505);
    layer4_outputs(6170) <= not(layer3_outputs(4309)) or (layer3_outputs(5552));
    layer4_outputs(6171) <= not(layer3_outputs(1661)) or (layer3_outputs(3190));
    layer4_outputs(6172) <= not(layer3_outputs(7631));
    layer4_outputs(6173) <= not(layer3_outputs(6487));
    layer4_outputs(6174) <= (layer3_outputs(5862)) xor (layer3_outputs(3311));
    layer4_outputs(6175) <= (layer3_outputs(3573)) and (layer3_outputs(1097));
    layer4_outputs(6176) <= '1';
    layer4_outputs(6177) <= layer3_outputs(6743);
    layer4_outputs(6178) <= (layer3_outputs(2737)) and not (layer3_outputs(6076));
    layer4_outputs(6179) <= not(layer3_outputs(4208));
    layer4_outputs(6180) <= not(layer3_outputs(5117));
    layer4_outputs(6181) <= not(layer3_outputs(6799));
    layer4_outputs(6182) <= not((layer3_outputs(570)) and (layer3_outputs(6514)));
    layer4_outputs(6183) <= '1';
    layer4_outputs(6184) <= layer3_outputs(2726);
    layer4_outputs(6185) <= layer3_outputs(655);
    layer4_outputs(6186) <= (layer3_outputs(4001)) and not (layer3_outputs(6146));
    layer4_outputs(6187) <= not(layer3_outputs(5052));
    layer4_outputs(6188) <= layer3_outputs(2194);
    layer4_outputs(6189) <= (layer3_outputs(1747)) xor (layer3_outputs(4231));
    layer4_outputs(6190) <= not(layer3_outputs(1485));
    layer4_outputs(6191) <= not(layer3_outputs(6898)) or (layer3_outputs(1639));
    layer4_outputs(6192) <= not(layer3_outputs(7260));
    layer4_outputs(6193) <= (layer3_outputs(4947)) and not (layer3_outputs(4485));
    layer4_outputs(6194) <= (layer3_outputs(7608)) and not (layer3_outputs(1734));
    layer4_outputs(6195) <= (layer3_outputs(667)) or (layer3_outputs(560));
    layer4_outputs(6196) <= layer3_outputs(7322);
    layer4_outputs(6197) <= layer3_outputs(7599);
    layer4_outputs(6198) <= not(layer3_outputs(7435));
    layer4_outputs(6199) <= '1';
    layer4_outputs(6200) <= '0';
    layer4_outputs(6201) <= not(layer3_outputs(925));
    layer4_outputs(6202) <= '0';
    layer4_outputs(6203) <= not(layer3_outputs(6776));
    layer4_outputs(6204) <= '1';
    layer4_outputs(6205) <= layer3_outputs(860);
    layer4_outputs(6206) <= not(layer3_outputs(6073));
    layer4_outputs(6207) <= (layer3_outputs(791)) and (layer3_outputs(3158));
    layer4_outputs(6208) <= not(layer3_outputs(5271)) or (layer3_outputs(388));
    layer4_outputs(6209) <= (layer3_outputs(275)) and not (layer3_outputs(6289));
    layer4_outputs(6210) <= not((layer3_outputs(6597)) and (layer3_outputs(4473)));
    layer4_outputs(6211) <= not(layer3_outputs(6249));
    layer4_outputs(6212) <= (layer3_outputs(2007)) xor (layer3_outputs(6106));
    layer4_outputs(6213) <= (layer3_outputs(3455)) and not (layer3_outputs(2655));
    layer4_outputs(6214) <= not(layer3_outputs(1309));
    layer4_outputs(6215) <= layer3_outputs(3393);
    layer4_outputs(6216) <= (layer3_outputs(4800)) and not (layer3_outputs(1940));
    layer4_outputs(6217) <= layer3_outputs(3362);
    layer4_outputs(6218) <= not(layer3_outputs(7626)) or (layer3_outputs(2705));
    layer4_outputs(6219) <= (layer3_outputs(7351)) xor (layer3_outputs(7614));
    layer4_outputs(6220) <= not((layer3_outputs(1061)) xor (layer3_outputs(4538)));
    layer4_outputs(6221) <= layer3_outputs(5201);
    layer4_outputs(6222) <= '1';
    layer4_outputs(6223) <= not(layer3_outputs(2098)) or (layer3_outputs(2924));
    layer4_outputs(6224) <= layer3_outputs(6987);
    layer4_outputs(6225) <= (layer3_outputs(4477)) or (layer3_outputs(1554));
    layer4_outputs(6226) <= '1';
    layer4_outputs(6227) <= not(layer3_outputs(828));
    layer4_outputs(6228) <= not((layer3_outputs(7023)) and (layer3_outputs(2871)));
    layer4_outputs(6229) <= not(layer3_outputs(7397));
    layer4_outputs(6230) <= layer3_outputs(210);
    layer4_outputs(6231) <= not(layer3_outputs(253));
    layer4_outputs(6232) <= (layer3_outputs(5867)) xor (layer3_outputs(6354));
    layer4_outputs(6233) <= (layer3_outputs(4453)) and not (layer3_outputs(3871));
    layer4_outputs(6234) <= (layer3_outputs(7132)) or (layer3_outputs(4535));
    layer4_outputs(6235) <= '0';
    layer4_outputs(6236) <= not(layer3_outputs(2948));
    layer4_outputs(6237) <= (layer3_outputs(3550)) and (layer3_outputs(2380));
    layer4_outputs(6238) <= layer3_outputs(7530);
    layer4_outputs(6239) <= (layer3_outputs(3964)) and not (layer3_outputs(2715));
    layer4_outputs(6240) <= (layer3_outputs(3196)) and (layer3_outputs(1410));
    layer4_outputs(6241) <= not(layer3_outputs(2924)) or (layer3_outputs(503));
    layer4_outputs(6242) <= layer3_outputs(2037);
    layer4_outputs(6243) <= not((layer3_outputs(1498)) or (layer3_outputs(5855)));
    layer4_outputs(6244) <= '1';
    layer4_outputs(6245) <= (layer3_outputs(4285)) or (layer3_outputs(5533));
    layer4_outputs(6246) <= (layer3_outputs(6392)) and (layer3_outputs(1831));
    layer4_outputs(6247) <= not(layer3_outputs(673)) or (layer3_outputs(2613));
    layer4_outputs(6248) <= not(layer3_outputs(4721));
    layer4_outputs(6249) <= not(layer3_outputs(3662)) or (layer3_outputs(6906));
    layer4_outputs(6250) <= not(layer3_outputs(1783)) or (layer3_outputs(6002));
    layer4_outputs(6251) <= '1';
    layer4_outputs(6252) <= layer3_outputs(4501);
    layer4_outputs(6253) <= layer3_outputs(5781);
    layer4_outputs(6254) <= not(layer3_outputs(2244));
    layer4_outputs(6255) <= layer3_outputs(3442);
    layer4_outputs(6256) <= layer3_outputs(900);
    layer4_outputs(6257) <= (layer3_outputs(1774)) xor (layer3_outputs(2330));
    layer4_outputs(6258) <= '0';
    layer4_outputs(6259) <= not(layer3_outputs(6028)) or (layer3_outputs(5665));
    layer4_outputs(6260) <= (layer3_outputs(720)) xor (layer3_outputs(6113));
    layer4_outputs(6261) <= layer3_outputs(5232);
    layer4_outputs(6262) <= (layer3_outputs(2896)) xor (layer3_outputs(3384));
    layer4_outputs(6263) <= (layer3_outputs(1396)) and not (layer3_outputs(5871));
    layer4_outputs(6264) <= not((layer3_outputs(597)) and (layer3_outputs(436)));
    layer4_outputs(6265) <= layer3_outputs(4857);
    layer4_outputs(6266) <= not(layer3_outputs(1975));
    layer4_outputs(6267) <= not((layer3_outputs(4358)) or (layer3_outputs(5210)));
    layer4_outputs(6268) <= not(layer3_outputs(2890)) or (layer3_outputs(6166));
    layer4_outputs(6269) <= (layer3_outputs(4348)) and (layer3_outputs(1773));
    layer4_outputs(6270) <= not(layer3_outputs(1090));
    layer4_outputs(6271) <= (layer3_outputs(6889)) and not (layer3_outputs(6079));
    layer4_outputs(6272) <= (layer3_outputs(3383)) and not (layer3_outputs(4192));
    layer4_outputs(6273) <= layer3_outputs(6933);
    layer4_outputs(6274) <= not(layer3_outputs(5124));
    layer4_outputs(6275) <= (layer3_outputs(5761)) and (layer3_outputs(2496));
    layer4_outputs(6276) <= (layer3_outputs(3744)) and not (layer3_outputs(5066));
    layer4_outputs(6277) <= not(layer3_outputs(5319));
    layer4_outputs(6278) <= '0';
    layer4_outputs(6279) <= not((layer3_outputs(1671)) and (layer3_outputs(6965)));
    layer4_outputs(6280) <= not(layer3_outputs(4972));
    layer4_outputs(6281) <= layer3_outputs(5370);
    layer4_outputs(6282) <= layer3_outputs(7168);
    layer4_outputs(6283) <= not(layer3_outputs(3307));
    layer4_outputs(6284) <= not((layer3_outputs(2061)) and (layer3_outputs(2098)));
    layer4_outputs(6285) <= not(layer3_outputs(2217));
    layer4_outputs(6286) <= '0';
    layer4_outputs(6287) <= (layer3_outputs(7552)) and not (layer3_outputs(7654));
    layer4_outputs(6288) <= not((layer3_outputs(6560)) or (layer3_outputs(2719)));
    layer4_outputs(6289) <= (layer3_outputs(6827)) and not (layer3_outputs(6362));
    layer4_outputs(6290) <= (layer3_outputs(189)) and not (layer3_outputs(6830));
    layer4_outputs(6291) <= not(layer3_outputs(5801));
    layer4_outputs(6292) <= '0';
    layer4_outputs(6293) <= layer3_outputs(6312);
    layer4_outputs(6294) <= (layer3_outputs(1349)) and (layer3_outputs(4305));
    layer4_outputs(6295) <= not((layer3_outputs(5466)) or (layer3_outputs(1942)));
    layer4_outputs(6296) <= layer3_outputs(6305);
    layer4_outputs(6297) <= not(layer3_outputs(2103));
    layer4_outputs(6298) <= layer3_outputs(2563);
    layer4_outputs(6299) <= (layer3_outputs(4037)) and (layer3_outputs(1849));
    layer4_outputs(6300) <= (layer3_outputs(6043)) and not (layer3_outputs(2303));
    layer4_outputs(6301) <= (layer3_outputs(4786)) and not (layer3_outputs(5813));
    layer4_outputs(6302) <= (layer3_outputs(3367)) and not (layer3_outputs(4321));
    layer4_outputs(6303) <= not(layer3_outputs(3947)) or (layer3_outputs(2952));
    layer4_outputs(6304) <= layer3_outputs(5937);
    layer4_outputs(6305) <= not((layer3_outputs(787)) and (layer3_outputs(4136)));
    layer4_outputs(6306) <= not(layer3_outputs(1065));
    layer4_outputs(6307) <= not(layer3_outputs(3861)) or (layer3_outputs(5752));
    layer4_outputs(6308) <= not((layer3_outputs(158)) and (layer3_outputs(7198)));
    layer4_outputs(6309) <= '1';
    layer4_outputs(6310) <= layer3_outputs(5517);
    layer4_outputs(6311) <= layer3_outputs(7241);
    layer4_outputs(6312) <= (layer3_outputs(7322)) and (layer3_outputs(2470));
    layer4_outputs(6313) <= not((layer3_outputs(1102)) or (layer3_outputs(2086)));
    layer4_outputs(6314) <= layer3_outputs(4693);
    layer4_outputs(6315) <= not(layer3_outputs(6543));
    layer4_outputs(6316) <= (layer3_outputs(7361)) and not (layer3_outputs(5816));
    layer4_outputs(6317) <= layer3_outputs(2997);
    layer4_outputs(6318) <= not((layer3_outputs(5495)) xor (layer3_outputs(5434)));
    layer4_outputs(6319) <= not(layer3_outputs(6134));
    layer4_outputs(6320) <= (layer3_outputs(2843)) or (layer3_outputs(5920));
    layer4_outputs(6321) <= layer3_outputs(3858);
    layer4_outputs(6322) <= not(layer3_outputs(44));
    layer4_outputs(6323) <= (layer3_outputs(5983)) and not (layer3_outputs(521));
    layer4_outputs(6324) <= layer3_outputs(3098);
    layer4_outputs(6325) <= not(layer3_outputs(5821));
    layer4_outputs(6326) <= (layer3_outputs(5485)) and not (layer3_outputs(5342));
    layer4_outputs(6327) <= '1';
    layer4_outputs(6328) <= (layer3_outputs(4453)) or (layer3_outputs(6496));
    layer4_outputs(6329) <= '0';
    layer4_outputs(6330) <= not((layer3_outputs(4256)) or (layer3_outputs(2868)));
    layer4_outputs(6331) <= (layer3_outputs(6851)) xor (layer3_outputs(7223));
    layer4_outputs(6332) <= not(layer3_outputs(1409));
    layer4_outputs(6333) <= not(layer3_outputs(5222));
    layer4_outputs(6334) <= layer3_outputs(451);
    layer4_outputs(6335) <= layer3_outputs(3075);
    layer4_outputs(6336) <= layer3_outputs(3905);
    layer4_outputs(6337) <= (layer3_outputs(2425)) and not (layer3_outputs(1453));
    layer4_outputs(6338) <= layer3_outputs(4062);
    layer4_outputs(6339) <= (layer3_outputs(1848)) and not (layer3_outputs(7085));
    layer4_outputs(6340) <= not((layer3_outputs(6382)) and (layer3_outputs(2323)));
    layer4_outputs(6341) <= not((layer3_outputs(5590)) or (layer3_outputs(1615)));
    layer4_outputs(6342) <= not((layer3_outputs(4950)) and (layer3_outputs(1929)));
    layer4_outputs(6343) <= layer3_outputs(2484);
    layer4_outputs(6344) <= not(layer3_outputs(7123));
    layer4_outputs(6345) <= layer3_outputs(7406);
    layer4_outputs(6346) <= not((layer3_outputs(489)) xor (layer3_outputs(4011)));
    layer4_outputs(6347) <= layer3_outputs(4620);
    layer4_outputs(6348) <= (layer3_outputs(5517)) xor (layer3_outputs(6684));
    layer4_outputs(6349) <= not(layer3_outputs(3475)) or (layer3_outputs(1440));
    layer4_outputs(6350) <= not(layer3_outputs(601));
    layer4_outputs(6351) <= (layer3_outputs(6616)) xor (layer3_outputs(3790));
    layer4_outputs(6352) <= not(layer3_outputs(3062));
    layer4_outputs(6353) <= not(layer3_outputs(6328));
    layer4_outputs(6354) <= (layer3_outputs(7293)) or (layer3_outputs(7350));
    layer4_outputs(6355) <= not(layer3_outputs(3646));
    layer4_outputs(6356) <= (layer3_outputs(1411)) and not (layer3_outputs(1833));
    layer4_outputs(6357) <= layer3_outputs(680);
    layer4_outputs(6358) <= (layer3_outputs(4274)) and not (layer3_outputs(4833));
    layer4_outputs(6359) <= layer3_outputs(3530);
    layer4_outputs(6360) <= (layer3_outputs(233)) or (layer3_outputs(5917));
    layer4_outputs(6361) <= not((layer3_outputs(2669)) xor (layer3_outputs(2222)));
    layer4_outputs(6362) <= layer3_outputs(6187);
    layer4_outputs(6363) <= layer3_outputs(3824);
    layer4_outputs(6364) <= not((layer3_outputs(7243)) and (layer3_outputs(537)));
    layer4_outputs(6365) <= layer3_outputs(6475);
    layer4_outputs(6366) <= not(layer3_outputs(6159)) or (layer3_outputs(7472));
    layer4_outputs(6367) <= layer3_outputs(7342);
    layer4_outputs(6368) <= not(layer3_outputs(3269));
    layer4_outputs(6369) <= not(layer3_outputs(447)) or (layer3_outputs(6444));
    layer4_outputs(6370) <= not(layer3_outputs(667));
    layer4_outputs(6371) <= (layer3_outputs(5805)) and (layer3_outputs(2312));
    layer4_outputs(6372) <= (layer3_outputs(2839)) and (layer3_outputs(6110));
    layer4_outputs(6373) <= not(layer3_outputs(7112));
    layer4_outputs(6374) <= not(layer3_outputs(7455));
    layer4_outputs(6375) <= not(layer3_outputs(5169));
    layer4_outputs(6376) <= (layer3_outputs(2564)) and (layer3_outputs(4829));
    layer4_outputs(6377) <= not((layer3_outputs(5945)) and (layer3_outputs(5884)));
    layer4_outputs(6378) <= not(layer3_outputs(1101)) or (layer3_outputs(6938));
    layer4_outputs(6379) <= not(layer3_outputs(5458));
    layer4_outputs(6380) <= '0';
    layer4_outputs(6381) <= layer3_outputs(1871);
    layer4_outputs(6382) <= not(layer3_outputs(5534)) or (layer3_outputs(2494));
    layer4_outputs(6383) <= (layer3_outputs(2831)) xor (layer3_outputs(1160));
    layer4_outputs(6384) <= not((layer3_outputs(661)) and (layer3_outputs(5592)));
    layer4_outputs(6385) <= not((layer3_outputs(636)) and (layer3_outputs(5186)));
    layer4_outputs(6386) <= not(layer3_outputs(4852));
    layer4_outputs(6387) <= '1';
    layer4_outputs(6388) <= layer3_outputs(4551);
    layer4_outputs(6389) <= not(layer3_outputs(580));
    layer4_outputs(6390) <= (layer3_outputs(4602)) or (layer3_outputs(2515));
    layer4_outputs(6391) <= not(layer3_outputs(3168));
    layer4_outputs(6392) <= layer3_outputs(4620);
    layer4_outputs(6393) <= not(layer3_outputs(5203));
    layer4_outputs(6394) <= not(layer3_outputs(2069)) or (layer3_outputs(1486));
    layer4_outputs(6395) <= not(layer3_outputs(1339));
    layer4_outputs(6396) <= not((layer3_outputs(3499)) and (layer3_outputs(1004)));
    layer4_outputs(6397) <= '1';
    layer4_outputs(6398) <= not((layer3_outputs(5904)) and (layer3_outputs(4864)));
    layer4_outputs(6399) <= '1';
    layer4_outputs(6400) <= (layer3_outputs(5606)) or (layer3_outputs(2961));
    layer4_outputs(6401) <= (layer3_outputs(4275)) and not (layer3_outputs(1191));
    layer4_outputs(6402) <= not((layer3_outputs(5700)) and (layer3_outputs(5337)));
    layer4_outputs(6403) <= not(layer3_outputs(1468)) or (layer3_outputs(3912));
    layer4_outputs(6404) <= not(layer3_outputs(2649)) or (layer3_outputs(2556));
    layer4_outputs(6405) <= (layer3_outputs(5587)) and not (layer3_outputs(5261));
    layer4_outputs(6406) <= not(layer3_outputs(4404)) or (layer3_outputs(7503));
    layer4_outputs(6407) <= not((layer3_outputs(4671)) and (layer3_outputs(4653)));
    layer4_outputs(6408) <= layer3_outputs(2439);
    layer4_outputs(6409) <= (layer3_outputs(2892)) and not (layer3_outputs(3211));
    layer4_outputs(6410) <= not((layer3_outputs(2049)) or (layer3_outputs(7396)));
    layer4_outputs(6411) <= not((layer3_outputs(6049)) or (layer3_outputs(1821)));
    layer4_outputs(6412) <= not(layer3_outputs(6275));
    layer4_outputs(6413) <= layer3_outputs(2768);
    layer4_outputs(6414) <= layer3_outputs(6409);
    layer4_outputs(6415) <= not((layer3_outputs(6014)) or (layer3_outputs(5064)));
    layer4_outputs(6416) <= (layer3_outputs(1370)) and not (layer3_outputs(6649));
    layer4_outputs(6417) <= (layer3_outputs(6566)) and not (layer3_outputs(2892));
    layer4_outputs(6418) <= (layer3_outputs(6042)) or (layer3_outputs(3763));
    layer4_outputs(6419) <= not((layer3_outputs(2730)) xor (layer3_outputs(2061)));
    layer4_outputs(6420) <= not(layer3_outputs(1238)) or (layer3_outputs(5413));
    layer4_outputs(6421) <= not(layer3_outputs(2731));
    layer4_outputs(6422) <= layer3_outputs(194);
    layer4_outputs(6423) <= (layer3_outputs(4202)) and not (layer3_outputs(7417));
    layer4_outputs(6424) <= layer3_outputs(3893);
    layer4_outputs(6425) <= not(layer3_outputs(2542));
    layer4_outputs(6426) <= not(layer3_outputs(3020));
    layer4_outputs(6427) <= layer3_outputs(5979);
    layer4_outputs(6428) <= (layer3_outputs(4914)) and (layer3_outputs(1962));
    layer4_outputs(6429) <= not(layer3_outputs(1583)) or (layer3_outputs(5641));
    layer4_outputs(6430) <= layer3_outputs(2450);
    layer4_outputs(6431) <= '1';
    layer4_outputs(6432) <= layer3_outputs(5576);
    layer4_outputs(6433) <= not(layer3_outputs(5177));
    layer4_outputs(6434) <= (layer3_outputs(2298)) or (layer3_outputs(290));
    layer4_outputs(6435) <= (layer3_outputs(6078)) and not (layer3_outputs(5986));
    layer4_outputs(6436) <= not((layer3_outputs(7189)) and (layer3_outputs(6743)));
    layer4_outputs(6437) <= not(layer3_outputs(646));
    layer4_outputs(6438) <= (layer3_outputs(2049)) and not (layer3_outputs(4145));
    layer4_outputs(6439) <= layer3_outputs(889);
    layer4_outputs(6440) <= not(layer3_outputs(5898));
    layer4_outputs(6441) <= not((layer3_outputs(5638)) or (layer3_outputs(4243)));
    layer4_outputs(6442) <= not((layer3_outputs(7660)) and (layer3_outputs(6141)));
    layer4_outputs(6443) <= (layer3_outputs(2691)) and not (layer3_outputs(6847));
    layer4_outputs(6444) <= (layer3_outputs(2253)) or (layer3_outputs(2947));
    layer4_outputs(6445) <= layer3_outputs(6482);
    layer4_outputs(6446) <= (layer3_outputs(7504)) and not (layer3_outputs(4366));
    layer4_outputs(6447) <= layer3_outputs(3593);
    layer4_outputs(6448) <= layer3_outputs(7667);
    layer4_outputs(6449) <= layer3_outputs(6304);
    layer4_outputs(6450) <= layer3_outputs(6632);
    layer4_outputs(6451) <= layer3_outputs(5122);
    layer4_outputs(6452) <= layer3_outputs(5206);
    layer4_outputs(6453) <= layer3_outputs(1018);
    layer4_outputs(6454) <= '0';
    layer4_outputs(6455) <= not(layer3_outputs(330)) or (layer3_outputs(1593));
    layer4_outputs(6456) <= (layer3_outputs(4240)) and not (layer3_outputs(4728));
    layer4_outputs(6457) <= '0';
    layer4_outputs(6458) <= not((layer3_outputs(1698)) or (layer3_outputs(7141)));
    layer4_outputs(6459) <= (layer3_outputs(5194)) or (layer3_outputs(7148));
    layer4_outputs(6460) <= (layer3_outputs(3302)) and not (layer3_outputs(6291));
    layer4_outputs(6461) <= layer3_outputs(2196);
    layer4_outputs(6462) <= not((layer3_outputs(3380)) and (layer3_outputs(5963)));
    layer4_outputs(6463) <= not((layer3_outputs(5856)) and (layer3_outputs(4812)));
    layer4_outputs(6464) <= not(layer3_outputs(6061));
    layer4_outputs(6465) <= (layer3_outputs(3998)) and not (layer3_outputs(5433));
    layer4_outputs(6466) <= not((layer3_outputs(7655)) or (layer3_outputs(146)));
    layer4_outputs(6467) <= (layer3_outputs(331)) and (layer3_outputs(1822));
    layer4_outputs(6468) <= layer3_outputs(5193);
    layer4_outputs(6469) <= layer3_outputs(5189);
    layer4_outputs(6470) <= not(layer3_outputs(1270));
    layer4_outputs(6471) <= not(layer3_outputs(6786));
    layer4_outputs(6472) <= (layer3_outputs(3146)) and not (layer3_outputs(3060));
    layer4_outputs(6473) <= (layer3_outputs(4597)) and (layer3_outputs(3119));
    layer4_outputs(6474) <= layer3_outputs(5536);
    layer4_outputs(6475) <= layer3_outputs(3561);
    layer4_outputs(6476) <= (layer3_outputs(4634)) and not (layer3_outputs(7558));
    layer4_outputs(6477) <= layer3_outputs(6217);
    layer4_outputs(6478) <= (layer3_outputs(6459)) or (layer3_outputs(4615));
    layer4_outputs(6479) <= not(layer3_outputs(7590));
    layer4_outputs(6480) <= not(layer3_outputs(3846));
    layer4_outputs(6481) <= not(layer3_outputs(1122));
    layer4_outputs(6482) <= (layer3_outputs(4834)) and (layer3_outputs(4021));
    layer4_outputs(6483) <= layer3_outputs(3426);
    layer4_outputs(6484) <= (layer3_outputs(4579)) xor (layer3_outputs(735));
    layer4_outputs(6485) <= layer3_outputs(3618);
    layer4_outputs(6486) <= (layer3_outputs(5611)) xor (layer3_outputs(3770));
    layer4_outputs(6487) <= layer3_outputs(5613);
    layer4_outputs(6488) <= (layer3_outputs(7264)) and not (layer3_outputs(6531));
    layer4_outputs(6489) <= (layer3_outputs(4199)) and not (layer3_outputs(1965));
    layer4_outputs(6490) <= not(layer3_outputs(2907));
    layer4_outputs(6491) <= not(layer3_outputs(3201));
    layer4_outputs(6492) <= layer3_outputs(568);
    layer4_outputs(6493) <= not((layer3_outputs(1636)) xor (layer3_outputs(638)));
    layer4_outputs(6494) <= not(layer3_outputs(5957));
    layer4_outputs(6495) <= '1';
    layer4_outputs(6496) <= layer3_outputs(167);
    layer4_outputs(6497) <= '1';
    layer4_outputs(6498) <= not(layer3_outputs(7236));
    layer4_outputs(6499) <= not((layer3_outputs(1708)) and (layer3_outputs(5475)));
    layer4_outputs(6500) <= (layer3_outputs(4463)) and (layer3_outputs(284));
    layer4_outputs(6501) <= layer3_outputs(2354);
    layer4_outputs(6502) <= (layer3_outputs(7509)) and (layer3_outputs(5195));
    layer4_outputs(6503) <= not(layer3_outputs(4076)) or (layer3_outputs(478));
    layer4_outputs(6504) <= '0';
    layer4_outputs(6505) <= not((layer3_outputs(2293)) or (layer3_outputs(1952)));
    layer4_outputs(6506) <= not(layer3_outputs(2709)) or (layer3_outputs(7310));
    layer4_outputs(6507) <= not((layer3_outputs(1442)) xor (layer3_outputs(1182)));
    layer4_outputs(6508) <= not((layer3_outputs(7005)) and (layer3_outputs(4338)));
    layer4_outputs(6509) <= layer3_outputs(1170);
    layer4_outputs(6510) <= not(layer3_outputs(6961)) or (layer3_outputs(6954));
    layer4_outputs(6511) <= not(layer3_outputs(2169));
    layer4_outputs(6512) <= layer3_outputs(3252);
    layer4_outputs(6513) <= layer3_outputs(1117);
    layer4_outputs(6514) <= (layer3_outputs(5058)) and not (layer3_outputs(3537));
    layer4_outputs(6515) <= not((layer3_outputs(5314)) xor (layer3_outputs(6834)));
    layer4_outputs(6516) <= not(layer3_outputs(4248)) or (layer3_outputs(53));
    layer4_outputs(6517) <= (layer3_outputs(2859)) or (layer3_outputs(1648));
    layer4_outputs(6518) <= not(layer3_outputs(4365));
    layer4_outputs(6519) <= layer3_outputs(2544);
    layer4_outputs(6520) <= (layer3_outputs(2866)) and not (layer3_outputs(513));
    layer4_outputs(6521) <= layer3_outputs(2637);
    layer4_outputs(6522) <= not((layer3_outputs(4919)) or (layer3_outputs(3132)));
    layer4_outputs(6523) <= '1';
    layer4_outputs(6524) <= (layer3_outputs(6008)) or (layer3_outputs(5273));
    layer4_outputs(6525) <= layer3_outputs(6179);
    layer4_outputs(6526) <= '1';
    layer4_outputs(6527) <= not(layer3_outputs(7133)) or (layer3_outputs(3594));
    layer4_outputs(6528) <= not((layer3_outputs(4402)) xor (layer3_outputs(5075)));
    layer4_outputs(6529) <= not(layer3_outputs(2232)) or (layer3_outputs(932));
    layer4_outputs(6530) <= not(layer3_outputs(6874));
    layer4_outputs(6531) <= '0';
    layer4_outputs(6532) <= (layer3_outputs(901)) and (layer3_outputs(7316));
    layer4_outputs(6533) <= (layer3_outputs(3803)) and not (layer3_outputs(6002));
    layer4_outputs(6534) <= not(layer3_outputs(2764)) or (layer3_outputs(6949));
    layer4_outputs(6535) <= not(layer3_outputs(978)) or (layer3_outputs(499));
    layer4_outputs(6536) <= layer3_outputs(654);
    layer4_outputs(6537) <= layer3_outputs(746);
    layer4_outputs(6538) <= not((layer3_outputs(3096)) xor (layer3_outputs(4286)));
    layer4_outputs(6539) <= not(layer3_outputs(163)) or (layer3_outputs(4232));
    layer4_outputs(6540) <= '1';
    layer4_outputs(6541) <= not(layer3_outputs(3820));
    layer4_outputs(6542) <= (layer3_outputs(3422)) and not (layer3_outputs(5984));
    layer4_outputs(6543) <= not((layer3_outputs(7617)) or (layer3_outputs(203)));
    layer4_outputs(6544) <= not(layer3_outputs(2593));
    layer4_outputs(6545) <= '1';
    layer4_outputs(6546) <= layer3_outputs(3269);
    layer4_outputs(6547) <= not((layer3_outputs(2653)) xor (layer3_outputs(6147)));
    layer4_outputs(6548) <= layer3_outputs(7181);
    layer4_outputs(6549) <= (layer3_outputs(5958)) and not (layer3_outputs(1645));
    layer4_outputs(6550) <= layer3_outputs(4616);
    layer4_outputs(6551) <= (layer3_outputs(3849)) and (layer3_outputs(5265));
    layer4_outputs(6552) <= not((layer3_outputs(4904)) xor (layer3_outputs(7630)));
    layer4_outputs(6553) <= (layer3_outputs(6705)) and not (layer3_outputs(3883));
    layer4_outputs(6554) <= (layer3_outputs(3114)) xor (layer3_outputs(4874));
    layer4_outputs(6555) <= layer3_outputs(4239);
    layer4_outputs(6556) <= not((layer3_outputs(1662)) xor (layer3_outputs(1432)));
    layer4_outputs(6557) <= (layer3_outputs(1424)) and not (layer3_outputs(3242));
    layer4_outputs(6558) <= not(layer3_outputs(5849)) or (layer3_outputs(919));
    layer4_outputs(6559) <= not(layer3_outputs(5886)) or (layer3_outputs(4336));
    layer4_outputs(6560) <= (layer3_outputs(7410)) and (layer3_outputs(6430));
    layer4_outputs(6561) <= (layer3_outputs(2488)) xor (layer3_outputs(4211));
    layer4_outputs(6562) <= not(layer3_outputs(4504)) or (layer3_outputs(6567));
    layer4_outputs(6563) <= (layer3_outputs(6648)) and not (layer3_outputs(404));
    layer4_outputs(6564) <= (layer3_outputs(1249)) and not (layer3_outputs(2766));
    layer4_outputs(6565) <= not(layer3_outputs(1970));
    layer4_outputs(6566) <= not((layer3_outputs(7279)) or (layer3_outputs(2379)));
    layer4_outputs(6567) <= not(layer3_outputs(1782));
    layer4_outputs(6568) <= layer3_outputs(863);
    layer4_outputs(6569) <= not((layer3_outputs(3896)) and (layer3_outputs(5033)));
    layer4_outputs(6570) <= (layer3_outputs(1879)) or (layer3_outputs(348));
    layer4_outputs(6571) <= layer3_outputs(3230);
    layer4_outputs(6572) <= (layer3_outputs(4457)) and not (layer3_outputs(4946));
    layer4_outputs(6573) <= layer3_outputs(3939);
    layer4_outputs(6574) <= layer3_outputs(493);
    layer4_outputs(6575) <= layer3_outputs(5556);
    layer4_outputs(6576) <= not(layer3_outputs(2312));
    layer4_outputs(6577) <= not((layer3_outputs(5666)) or (layer3_outputs(5336)));
    layer4_outputs(6578) <= not(layer3_outputs(3671));
    layer4_outputs(6579) <= '1';
    layer4_outputs(6580) <= (layer3_outputs(3407)) or (layer3_outputs(2050));
    layer4_outputs(6581) <= layer3_outputs(696);
    layer4_outputs(6582) <= (layer3_outputs(1926)) or (layer3_outputs(5651));
    layer4_outputs(6583) <= (layer3_outputs(3875)) xor (layer3_outputs(5756));
    layer4_outputs(6584) <= layer3_outputs(5233);
    layer4_outputs(6585) <= not((layer3_outputs(4692)) and (layer3_outputs(1185)));
    layer4_outputs(6586) <= (layer3_outputs(4439)) and not (layer3_outputs(7425));
    layer4_outputs(6587) <= layer3_outputs(3009);
    layer4_outputs(6588) <= not((layer3_outputs(6443)) and (layer3_outputs(5878)));
    layer4_outputs(6589) <= not((layer3_outputs(6410)) and (layer3_outputs(6415)));
    layer4_outputs(6590) <= not((layer3_outputs(861)) xor (layer3_outputs(2349)));
    layer4_outputs(6591) <= not(layer3_outputs(2214));
    layer4_outputs(6592) <= not(layer3_outputs(2111));
    layer4_outputs(6593) <= not(layer3_outputs(5387));
    layer4_outputs(6594) <= layer3_outputs(5231);
    layer4_outputs(6595) <= not(layer3_outputs(5432)) or (layer3_outputs(6922));
    layer4_outputs(6596) <= (layer3_outputs(7204)) or (layer3_outputs(1741));
    layer4_outputs(6597) <= not(layer3_outputs(2534)) or (layer3_outputs(2408));
    layer4_outputs(6598) <= not((layer3_outputs(2798)) or (layer3_outputs(6555)));
    layer4_outputs(6599) <= layer3_outputs(1413);
    layer4_outputs(6600) <= (layer3_outputs(3081)) and not (layer3_outputs(6161));
    layer4_outputs(6601) <= (layer3_outputs(6595)) or (layer3_outputs(3305));
    layer4_outputs(6602) <= not(layer3_outputs(2421));
    layer4_outputs(6603) <= not(layer3_outputs(2406)) or (layer3_outputs(3723));
    layer4_outputs(6604) <= (layer3_outputs(5677)) and not (layer3_outputs(4905));
    layer4_outputs(6605) <= '1';
    layer4_outputs(6606) <= not(layer3_outputs(2540)) or (layer3_outputs(5592));
    layer4_outputs(6607) <= layer3_outputs(4820);
    layer4_outputs(6608) <= not(layer3_outputs(818)) or (layer3_outputs(4210));
    layer4_outputs(6609) <= not(layer3_outputs(3760));
    layer4_outputs(6610) <= '0';
    layer4_outputs(6611) <= not(layer3_outputs(3728));
    layer4_outputs(6612) <= not((layer3_outputs(4403)) and (layer3_outputs(5496)));
    layer4_outputs(6613) <= layer3_outputs(5356);
    layer4_outputs(6614) <= not(layer3_outputs(6981));
    layer4_outputs(6615) <= (layer3_outputs(2748)) xor (layer3_outputs(4880));
    layer4_outputs(6616) <= layer3_outputs(1659);
    layer4_outputs(6617) <= not(layer3_outputs(3206));
    layer4_outputs(6618) <= not((layer3_outputs(5662)) and (layer3_outputs(93)));
    layer4_outputs(6619) <= layer3_outputs(285);
    layer4_outputs(6620) <= (layer3_outputs(7484)) xor (layer3_outputs(3170));
    layer4_outputs(6621) <= (layer3_outputs(3518)) or (layer3_outputs(3293));
    layer4_outputs(6622) <= (layer3_outputs(7606)) xor (layer3_outputs(4172));
    layer4_outputs(6623) <= not(layer3_outputs(4860));
    layer4_outputs(6624) <= (layer3_outputs(63)) xor (layer3_outputs(157));
    layer4_outputs(6625) <= not(layer3_outputs(5208));
    layer4_outputs(6626) <= layer3_outputs(6357);
    layer4_outputs(6627) <= not(layer3_outputs(1894)) or (layer3_outputs(6019));
    layer4_outputs(6628) <= layer3_outputs(7647);
    layer4_outputs(6629) <= (layer3_outputs(3403)) and (layer3_outputs(5493));
    layer4_outputs(6630) <= not(layer3_outputs(1780));
    layer4_outputs(6631) <= not((layer3_outputs(3089)) and (layer3_outputs(6024)));
    layer4_outputs(6632) <= not(layer3_outputs(7288)) or (layer3_outputs(2420));
    layer4_outputs(6633) <= layer3_outputs(6708);
    layer4_outputs(6634) <= (layer3_outputs(1920)) or (layer3_outputs(5379));
    layer4_outputs(6635) <= '1';
    layer4_outputs(6636) <= layer3_outputs(3563);
    layer4_outputs(6637) <= not(layer3_outputs(6373));
    layer4_outputs(6638) <= (layer3_outputs(3907)) and not (layer3_outputs(5964));
    layer4_outputs(6639) <= (layer3_outputs(7250)) or (layer3_outputs(2690));
    layer4_outputs(6640) <= (layer3_outputs(4733)) xor (layer3_outputs(2751));
    layer4_outputs(6641) <= layer3_outputs(1598);
    layer4_outputs(6642) <= layer3_outputs(4164);
    layer4_outputs(6643) <= not(layer3_outputs(4474)) or (layer3_outputs(3219));
    layer4_outputs(6644) <= '1';
    layer4_outputs(6645) <= not(layer3_outputs(6505)) or (layer3_outputs(2175));
    layer4_outputs(6646) <= (layer3_outputs(7372)) and not (layer3_outputs(1135));
    layer4_outputs(6647) <= (layer3_outputs(100)) or (layer3_outputs(1824));
    layer4_outputs(6648) <= not(layer3_outputs(3340)) or (layer3_outputs(1316));
    layer4_outputs(6649) <= layer3_outputs(2623);
    layer4_outputs(6650) <= (layer3_outputs(516)) and not (layer3_outputs(3490));
    layer4_outputs(6651) <= layer3_outputs(4127);
    layer4_outputs(6652) <= not(layer3_outputs(128));
    layer4_outputs(6653) <= (layer3_outputs(6216)) xor (layer3_outputs(4701));
    layer4_outputs(6654) <= not((layer3_outputs(1666)) or (layer3_outputs(906)));
    layer4_outputs(6655) <= not(layer3_outputs(1350));
    layer4_outputs(6656) <= not((layer3_outputs(4219)) and (layer3_outputs(7270)));
    layer4_outputs(6657) <= not(layer3_outputs(1281));
    layer4_outputs(6658) <= not(layer3_outputs(3074));
    layer4_outputs(6659) <= '1';
    layer4_outputs(6660) <= not((layer3_outputs(1677)) or (layer3_outputs(6912)));
    layer4_outputs(6661) <= (layer3_outputs(7608)) xor (layer3_outputs(5987));
    layer4_outputs(6662) <= (layer3_outputs(1917)) and (layer3_outputs(1888));
    layer4_outputs(6663) <= layer3_outputs(6716);
    layer4_outputs(6664) <= not(layer3_outputs(4611));
    layer4_outputs(6665) <= layer3_outputs(1794);
    layer4_outputs(6666) <= not((layer3_outputs(1763)) or (layer3_outputs(2437)));
    layer4_outputs(6667) <= '0';
    layer4_outputs(6668) <= layer3_outputs(6592);
    layer4_outputs(6669) <= (layer3_outputs(5272)) and (layer3_outputs(294));
    layer4_outputs(6670) <= (layer3_outputs(5805)) or (layer3_outputs(7376));
    layer4_outputs(6671) <= (layer3_outputs(2248)) or (layer3_outputs(5056));
    layer4_outputs(6672) <= layer3_outputs(6698);
    layer4_outputs(6673) <= not(layer3_outputs(388));
    layer4_outputs(6674) <= not(layer3_outputs(7140));
    layer4_outputs(6675) <= not(layer3_outputs(3557));
    layer4_outputs(6676) <= '0';
    layer4_outputs(6677) <= (layer3_outputs(931)) and not (layer3_outputs(5236));
    layer4_outputs(6678) <= '1';
    layer4_outputs(6679) <= layer3_outputs(2628);
    layer4_outputs(6680) <= not((layer3_outputs(5514)) and (layer3_outputs(3725)));
    layer4_outputs(6681) <= not(layer3_outputs(6265)) or (layer3_outputs(2007));
    layer4_outputs(6682) <= not((layer3_outputs(166)) and (layer3_outputs(3339)));
    layer4_outputs(6683) <= (layer3_outputs(5736)) and (layer3_outputs(377));
    layer4_outputs(6684) <= not(layer3_outputs(2324)) or (layer3_outputs(4112));
    layer4_outputs(6685) <= not((layer3_outputs(1633)) and (layer3_outputs(6525)));
    layer4_outputs(6686) <= (layer3_outputs(6093)) and not (layer3_outputs(1553));
    layer4_outputs(6687) <= layer3_outputs(5752);
    layer4_outputs(6688) <= (layer3_outputs(5569)) and not (layer3_outputs(6783));
    layer4_outputs(6689) <= layer3_outputs(2548);
    layer4_outputs(6690) <= (layer3_outputs(1959)) or (layer3_outputs(2226));
    layer4_outputs(6691) <= '0';
    layer4_outputs(6692) <= layer3_outputs(4351);
    layer4_outputs(6693) <= not(layer3_outputs(2933));
    layer4_outputs(6694) <= layer3_outputs(2513);
    layer4_outputs(6695) <= (layer3_outputs(6235)) and not (layer3_outputs(7335));
    layer4_outputs(6696) <= layer3_outputs(6499);
    layer4_outputs(6697) <= (layer3_outputs(3125)) and (layer3_outputs(7187));
    layer4_outputs(6698) <= '0';
    layer4_outputs(6699) <= not((layer3_outputs(6037)) and (layer3_outputs(2763)));
    layer4_outputs(6700) <= not(layer3_outputs(2994)) or (layer3_outputs(3888));
    layer4_outputs(6701) <= not((layer3_outputs(2832)) or (layer3_outputs(5209)));
    layer4_outputs(6702) <= not(layer3_outputs(3178)) or (layer3_outputs(5482));
    layer4_outputs(6703) <= layer3_outputs(3233);
    layer4_outputs(6704) <= (layer3_outputs(6699)) and not (layer3_outputs(2193));
    layer4_outputs(6705) <= layer3_outputs(3189);
    layer4_outputs(6706) <= not(layer3_outputs(3988));
    layer4_outputs(6707) <= layer3_outputs(2518);
    layer4_outputs(6708) <= '0';
    layer4_outputs(6709) <= not((layer3_outputs(5492)) xor (layer3_outputs(3684)));
    layer4_outputs(6710) <= '1';
    layer4_outputs(6711) <= layer3_outputs(1922);
    layer4_outputs(6712) <= not((layer3_outputs(5312)) xor (layer3_outputs(1530)));
    layer4_outputs(6713) <= not(layer3_outputs(2064));
    layer4_outputs(6714) <= (layer3_outputs(4331)) and not (layer3_outputs(7577));
    layer4_outputs(6715) <= not(layer3_outputs(6874)) or (layer3_outputs(2293));
    layer4_outputs(6716) <= not((layer3_outputs(960)) and (layer3_outputs(3113)));
    layer4_outputs(6717) <= layer3_outputs(1757);
    layer4_outputs(6718) <= not(layer3_outputs(518)) or (layer3_outputs(5267));
    layer4_outputs(6719) <= layer3_outputs(1953);
    layer4_outputs(6720) <= layer3_outputs(6275);
    layer4_outputs(6721) <= not(layer3_outputs(555));
    layer4_outputs(6722) <= layer3_outputs(7196);
    layer4_outputs(6723) <= not(layer3_outputs(6594)) or (layer3_outputs(3853));
    layer4_outputs(6724) <= layer3_outputs(5370);
    layer4_outputs(6725) <= not((layer3_outputs(3403)) or (layer3_outputs(1846)));
    layer4_outputs(6726) <= not(layer3_outputs(2634)) or (layer3_outputs(5948));
    layer4_outputs(6727) <= (layer3_outputs(2619)) or (layer3_outputs(5289));
    layer4_outputs(6728) <= not(layer3_outputs(3147)) or (layer3_outputs(6916));
    layer4_outputs(6729) <= not(layer3_outputs(4040)) or (layer3_outputs(3923));
    layer4_outputs(6730) <= (layer3_outputs(2493)) and (layer3_outputs(4974));
    layer4_outputs(6731) <= '1';
    layer4_outputs(6732) <= not(layer3_outputs(1939));
    layer4_outputs(6733) <= '0';
    layer4_outputs(6734) <= not((layer3_outputs(6640)) or (layer3_outputs(4678)));
    layer4_outputs(6735) <= (layer3_outputs(3337)) and not (layer3_outputs(992));
    layer4_outputs(6736) <= not((layer3_outputs(5674)) xor (layer3_outputs(6670)));
    layer4_outputs(6737) <= not(layer3_outputs(3363));
    layer4_outputs(6738) <= '0';
    layer4_outputs(6739) <= layer3_outputs(5436);
    layer4_outputs(6740) <= (layer3_outputs(5050)) and (layer3_outputs(2912));
    layer4_outputs(6741) <= (layer3_outputs(6798)) and not (layer3_outputs(7330));
    layer4_outputs(6742) <= not(layer3_outputs(4402)) or (layer3_outputs(6925));
    layer4_outputs(6743) <= not(layer3_outputs(4750)) or (layer3_outputs(4557));
    layer4_outputs(6744) <= not(layer3_outputs(1150));
    layer4_outputs(6745) <= not(layer3_outputs(2721)) or (layer3_outputs(1027));
    layer4_outputs(6746) <= layer3_outputs(2237);
    layer4_outputs(6747) <= not(layer3_outputs(1020)) or (layer3_outputs(6951));
    layer4_outputs(6748) <= (layer3_outputs(6031)) and (layer3_outputs(3634));
    layer4_outputs(6749) <= not(layer3_outputs(3484));
    layer4_outputs(6750) <= layer3_outputs(5374);
    layer4_outputs(6751) <= (layer3_outputs(5453)) xor (layer3_outputs(3524));
    layer4_outputs(6752) <= not(layer3_outputs(5197));
    layer4_outputs(6753) <= not(layer3_outputs(7657));
    layer4_outputs(6754) <= not(layer3_outputs(448)) or (layer3_outputs(4226));
    layer4_outputs(6755) <= not(layer3_outputs(2058));
    layer4_outputs(6756) <= layer3_outputs(1979);
    layer4_outputs(6757) <= (layer3_outputs(5688)) and not (layer3_outputs(4582));
    layer4_outputs(6758) <= (layer3_outputs(7556)) and not (layer3_outputs(4287));
    layer4_outputs(6759) <= not(layer3_outputs(95));
    layer4_outputs(6760) <= not(layer3_outputs(3259));
    layer4_outputs(6761) <= not(layer3_outputs(2605)) or (layer3_outputs(4732));
    layer4_outputs(6762) <= not(layer3_outputs(3712));
    layer4_outputs(6763) <= '1';
    layer4_outputs(6764) <= not((layer3_outputs(396)) and (layer3_outputs(1815)));
    layer4_outputs(6765) <= not(layer3_outputs(4380)) or (layer3_outputs(4799));
    layer4_outputs(6766) <= layer3_outputs(5687);
    layer4_outputs(6767) <= layer3_outputs(4045);
    layer4_outputs(6768) <= not(layer3_outputs(4358)) or (layer3_outputs(3388));
    layer4_outputs(6769) <= not((layer3_outputs(510)) and (layer3_outputs(3457)));
    layer4_outputs(6770) <= not(layer3_outputs(7007));
    layer4_outputs(6771) <= (layer3_outputs(6958)) xor (layer3_outputs(3632));
    layer4_outputs(6772) <= not(layer3_outputs(6584));
    layer4_outputs(6773) <= layer3_outputs(3453);
    layer4_outputs(6774) <= not((layer3_outputs(7361)) or (layer3_outputs(5859)));
    layer4_outputs(6775) <= layer3_outputs(5357);
    layer4_outputs(6776) <= layer3_outputs(4340);
    layer4_outputs(6777) <= not(layer3_outputs(7106)) or (layer3_outputs(4494));
    layer4_outputs(6778) <= not(layer3_outputs(1594));
    layer4_outputs(6779) <= not(layer3_outputs(4489));
    layer4_outputs(6780) <= not(layer3_outputs(5792)) or (layer3_outputs(6549));
    layer4_outputs(6781) <= not(layer3_outputs(129)) or (layer3_outputs(2842));
    layer4_outputs(6782) <= layer3_outputs(2510);
    layer4_outputs(6783) <= layer3_outputs(901);
    layer4_outputs(6784) <= layer3_outputs(2124);
    layer4_outputs(6785) <= layer3_outputs(397);
    layer4_outputs(6786) <= not((layer3_outputs(5418)) or (layer3_outputs(7160)));
    layer4_outputs(6787) <= '1';
    layer4_outputs(6788) <= not(layer3_outputs(5133));
    layer4_outputs(6789) <= (layer3_outputs(6382)) and not (layer3_outputs(2820));
    layer4_outputs(6790) <= not(layer3_outputs(3503));
    layer4_outputs(6791) <= not(layer3_outputs(749));
    layer4_outputs(6792) <= not(layer3_outputs(3727)) or (layer3_outputs(5638));
    layer4_outputs(6793) <= (layer3_outputs(6822)) or (layer3_outputs(7552));
    layer4_outputs(6794) <= layer3_outputs(1220);
    layer4_outputs(6795) <= not((layer3_outputs(3148)) or (layer3_outputs(2514)));
    layer4_outputs(6796) <= (layer3_outputs(4928)) and not (layer3_outputs(4373));
    layer4_outputs(6797) <= not(layer3_outputs(6615));
    layer4_outputs(6798) <= '1';
    layer4_outputs(6799) <= (layer3_outputs(6290)) and not (layer3_outputs(1589));
    layer4_outputs(6800) <= layer3_outputs(7162);
    layer4_outputs(6801) <= (layer3_outputs(1305)) xor (layer3_outputs(6952));
    layer4_outputs(6802) <= not(layer3_outputs(893));
    layer4_outputs(6803) <= layer3_outputs(4705);
    layer4_outputs(6804) <= not((layer3_outputs(1893)) and (layer3_outputs(88)));
    layer4_outputs(6805) <= not((layer3_outputs(6620)) or (layer3_outputs(4259)));
    layer4_outputs(6806) <= (layer3_outputs(744)) and (layer3_outputs(5069));
    layer4_outputs(6807) <= not(layer3_outputs(2366)) or (layer3_outputs(848));
    layer4_outputs(6808) <= not(layer3_outputs(2878)) or (layer3_outputs(7043));
    layer4_outputs(6809) <= (layer3_outputs(5509)) xor (layer3_outputs(1745));
    layer4_outputs(6810) <= not((layer3_outputs(7380)) and (layer3_outputs(6096)));
    layer4_outputs(6811) <= not((layer3_outputs(579)) and (layer3_outputs(1450)));
    layer4_outputs(6812) <= not(layer3_outputs(7288)) or (layer3_outputs(2044));
    layer4_outputs(6813) <= not(layer3_outputs(6618));
    layer4_outputs(6814) <= not(layer3_outputs(2703));
    layer4_outputs(6815) <= '0';
    layer4_outputs(6816) <= not((layer3_outputs(3739)) xor (layer3_outputs(6643)));
    layer4_outputs(6817) <= layer3_outputs(7292);
    layer4_outputs(6818) <= layer3_outputs(2841);
    layer4_outputs(6819) <= not(layer3_outputs(6768));
    layer4_outputs(6820) <= not((layer3_outputs(405)) or (layer3_outputs(3899)));
    layer4_outputs(6821) <= (layer3_outputs(2757)) and not (layer3_outputs(6561));
    layer4_outputs(6822) <= '1';
    layer4_outputs(6823) <= not(layer3_outputs(6969)) or (layer3_outputs(7161));
    layer4_outputs(6824) <= not(layer3_outputs(1806)) or (layer3_outputs(805));
    layer4_outputs(6825) <= not(layer3_outputs(5767));
    layer4_outputs(6826) <= '1';
    layer4_outputs(6827) <= not(layer3_outputs(5021));
    layer4_outputs(6828) <= (layer3_outputs(6670)) and not (layer3_outputs(936));
    layer4_outputs(6829) <= '1';
    layer4_outputs(6830) <= '0';
    layer4_outputs(6831) <= not(layer3_outputs(6289)) or (layer3_outputs(2021));
    layer4_outputs(6832) <= not(layer3_outputs(7050));
    layer4_outputs(6833) <= not((layer3_outputs(5953)) or (layer3_outputs(2110)));
    layer4_outputs(6834) <= '0';
    layer4_outputs(6835) <= not(layer3_outputs(3001));
    layer4_outputs(6836) <= not((layer3_outputs(2589)) and (layer3_outputs(2766)));
    layer4_outputs(6837) <= not(layer3_outputs(5426)) or (layer3_outputs(4627));
    layer4_outputs(6838) <= not((layer3_outputs(944)) and (layer3_outputs(5860)));
    layer4_outputs(6839) <= not((layer3_outputs(1104)) and (layer3_outputs(6627)));
    layer4_outputs(6840) <= not((layer3_outputs(4736)) and (layer3_outputs(2209)));
    layer4_outputs(6841) <= layer3_outputs(4603);
    layer4_outputs(6842) <= not((layer3_outputs(4153)) or (layer3_outputs(1303)));
    layer4_outputs(6843) <= not(layer3_outputs(771));
    layer4_outputs(6844) <= layer3_outputs(1787);
    layer4_outputs(6845) <= not(layer3_outputs(2701)) or (layer3_outputs(814));
    layer4_outputs(6846) <= not(layer3_outputs(2999));
    layer4_outputs(6847) <= layer3_outputs(4940);
    layer4_outputs(6848) <= (layer3_outputs(2390)) and (layer3_outputs(828));
    layer4_outputs(6849) <= '1';
    layer4_outputs(6850) <= not((layer3_outputs(2571)) and (layer3_outputs(6383)));
    layer4_outputs(6851) <= (layer3_outputs(349)) and (layer3_outputs(581));
    layer4_outputs(6852) <= not(layer3_outputs(2053)) or (layer3_outputs(5941));
    layer4_outputs(6853) <= (layer3_outputs(81)) or (layer3_outputs(1992));
    layer4_outputs(6854) <= (layer3_outputs(1466)) or (layer3_outputs(1733));
    layer4_outputs(6855) <= (layer3_outputs(5684)) or (layer3_outputs(5982));
    layer4_outputs(6856) <= not(layer3_outputs(969));
    layer4_outputs(6857) <= not((layer3_outputs(4810)) and (layer3_outputs(2524)));
    layer4_outputs(6858) <= not((layer3_outputs(6535)) and (layer3_outputs(1246)));
    layer4_outputs(6859) <= not(layer3_outputs(223));
    layer4_outputs(6860) <= layer3_outputs(7049);
    layer4_outputs(6861) <= not(layer3_outputs(4437));
    layer4_outputs(6862) <= '1';
    layer4_outputs(6863) <= layer3_outputs(7313);
    layer4_outputs(6864) <= layer3_outputs(6287);
    layer4_outputs(6865) <= not(layer3_outputs(6332));
    layer4_outputs(6866) <= not((layer3_outputs(1819)) and (layer3_outputs(5043)));
    layer4_outputs(6867) <= not(layer3_outputs(1003)) or (layer3_outputs(3087));
    layer4_outputs(6868) <= not(layer3_outputs(6100));
    layer4_outputs(6869) <= not(layer3_outputs(5734));
    layer4_outputs(6870) <= layer3_outputs(4434);
    layer4_outputs(6871) <= not(layer3_outputs(4198));
    layer4_outputs(6872) <= layer3_outputs(3275);
    layer4_outputs(6873) <= layer3_outputs(7262);
    layer4_outputs(6874) <= (layer3_outputs(1643)) and not (layer3_outputs(4176));
    layer4_outputs(6875) <= not(layer3_outputs(2694));
    layer4_outputs(6876) <= (layer3_outputs(323)) or (layer3_outputs(4146));
    layer4_outputs(6877) <= (layer3_outputs(2518)) xor (layer3_outputs(3375));
    layer4_outputs(6878) <= not(layer3_outputs(6273)) or (layer3_outputs(5043));
    layer4_outputs(6879) <= layer3_outputs(4057);
    layer4_outputs(6880) <= not(layer3_outputs(5757));
    layer4_outputs(6881) <= not(layer3_outputs(741));
    layer4_outputs(6882) <= not(layer3_outputs(3102));
    layer4_outputs(6883) <= '0';
    layer4_outputs(6884) <= not((layer3_outputs(6795)) and (layer3_outputs(5507)));
    layer4_outputs(6885) <= '0';
    layer4_outputs(6886) <= (layer3_outputs(7021)) and (layer3_outputs(2818));
    layer4_outputs(6887) <= (layer3_outputs(5271)) xor (layer3_outputs(284));
    layer4_outputs(6888) <= not(layer3_outputs(7447));
    layer4_outputs(6889) <= layer3_outputs(2750);
    layer4_outputs(6890) <= not(layer3_outputs(3320));
    layer4_outputs(6891) <= layer3_outputs(5196);
    layer4_outputs(6892) <= not(layer3_outputs(2331)) or (layer3_outputs(7248));
    layer4_outputs(6893) <= not((layer3_outputs(1008)) or (layer3_outputs(2411)));
    layer4_outputs(6894) <= (layer3_outputs(2599)) and not (layer3_outputs(4752));
    layer4_outputs(6895) <= (layer3_outputs(3282)) and (layer3_outputs(6842));
    layer4_outputs(6896) <= not((layer3_outputs(4667)) xor (layer3_outputs(617)));
    layer4_outputs(6897) <= not((layer3_outputs(3499)) or (layer3_outputs(1954)));
    layer4_outputs(6898) <= (layer3_outputs(3874)) and (layer3_outputs(1581));
    layer4_outputs(6899) <= layer3_outputs(6308);
    layer4_outputs(6900) <= not(layer3_outputs(6149)) or (layer3_outputs(6316));
    layer4_outputs(6901) <= '1';
    layer4_outputs(6902) <= not(layer3_outputs(2685)) or (layer3_outputs(360));
    layer4_outputs(6903) <= not((layer3_outputs(3640)) and (layer3_outputs(653)));
    layer4_outputs(6904) <= (layer3_outputs(3096)) and not (layer3_outputs(1118));
    layer4_outputs(6905) <= not(layer3_outputs(3597));
    layer4_outputs(6906) <= layer3_outputs(4849);
    layer4_outputs(6907) <= (layer3_outputs(5328)) and not (layer3_outputs(5003));
    layer4_outputs(6908) <= not(layer3_outputs(6)) or (layer3_outputs(5636));
    layer4_outputs(6909) <= (layer3_outputs(5946)) and not (layer3_outputs(7438));
    layer4_outputs(6910) <= not((layer3_outputs(6053)) xor (layer3_outputs(3980)));
    layer4_outputs(6911) <= (layer3_outputs(1013)) and not (layer3_outputs(6329));
    layer4_outputs(6912) <= not((layer3_outputs(4059)) or (layer3_outputs(1692)));
    layer4_outputs(6913) <= '0';
    layer4_outputs(6914) <= layer3_outputs(7450);
    layer4_outputs(6915) <= not((layer3_outputs(2265)) xor (layer3_outputs(3280)));
    layer4_outputs(6916) <= (layer3_outputs(1046)) and not (layer3_outputs(5077));
    layer4_outputs(6917) <= not(layer3_outputs(6892));
    layer4_outputs(6918) <= layer3_outputs(3743);
    layer4_outputs(6919) <= not(layer3_outputs(2790));
    layer4_outputs(6920) <= layer3_outputs(1829);
    layer4_outputs(6921) <= not(layer3_outputs(1690));
    layer4_outputs(6922) <= '1';
    layer4_outputs(6923) <= layer3_outputs(743);
    layer4_outputs(6924) <= (layer3_outputs(5646)) and (layer3_outputs(4240));
    layer4_outputs(6925) <= not(layer3_outputs(3480)) or (layer3_outputs(2963));
    layer4_outputs(6926) <= (layer3_outputs(1066)) or (layer3_outputs(3449));
    layer4_outputs(6927) <= not(layer3_outputs(3304)) or (layer3_outputs(2194));
    layer4_outputs(6928) <= '1';
    layer4_outputs(6929) <= layer3_outputs(2024);
    layer4_outputs(6930) <= (layer3_outputs(7330)) and (layer3_outputs(2954));
    layer4_outputs(6931) <= layer3_outputs(7307);
    layer4_outputs(6932) <= not(layer3_outputs(6317));
    layer4_outputs(6933) <= (layer3_outputs(4931)) or (layer3_outputs(6758));
    layer4_outputs(6934) <= not(layer3_outputs(319)) or (layer3_outputs(4673));
    layer4_outputs(6935) <= (layer3_outputs(6541)) and not (layer3_outputs(1285));
    layer4_outputs(6936) <= (layer3_outputs(3677)) xor (layer3_outputs(4061));
    layer4_outputs(6937) <= (layer3_outputs(1353)) and not (layer3_outputs(7372));
    layer4_outputs(6938) <= layer3_outputs(6956);
    layer4_outputs(6939) <= layer3_outputs(968);
    layer4_outputs(6940) <= layer3_outputs(1974);
    layer4_outputs(6941) <= not(layer3_outputs(4183));
    layer4_outputs(6942) <= not((layer3_outputs(5804)) and (layer3_outputs(3521)));
    layer4_outputs(6943) <= (layer3_outputs(3493)) or (layer3_outputs(1775));
    layer4_outputs(6944) <= (layer3_outputs(4038)) xor (layer3_outputs(385));
    layer4_outputs(6945) <= (layer3_outputs(2840)) or (layer3_outputs(1872));
    layer4_outputs(6946) <= not(layer3_outputs(3024));
    layer4_outputs(6947) <= (layer3_outputs(2381)) and (layer3_outputs(2649));
    layer4_outputs(6948) <= (layer3_outputs(1647)) and (layer3_outputs(7306));
    layer4_outputs(6949) <= not(layer3_outputs(1104));
    layer4_outputs(6950) <= not(layer3_outputs(187));
    layer4_outputs(6951) <= not(layer3_outputs(7277)) or (layer3_outputs(1243));
    layer4_outputs(6952) <= (layer3_outputs(1758)) and (layer3_outputs(2911));
    layer4_outputs(6953) <= layer3_outputs(4909);
    layer4_outputs(6954) <= (layer3_outputs(2434)) xor (layer3_outputs(4948));
    layer4_outputs(6955) <= layer3_outputs(3126);
    layer4_outputs(6956) <= not(layer3_outputs(5095)) or (layer3_outputs(4951));
    layer4_outputs(6957) <= layer3_outputs(1238);
    layer4_outputs(6958) <= not((layer3_outputs(3783)) and (layer3_outputs(2666)));
    layer4_outputs(6959) <= (layer3_outputs(1538)) or (layer3_outputs(4005));
    layer4_outputs(6960) <= (layer3_outputs(2733)) and not (layer3_outputs(1265));
    layer4_outputs(6961) <= not(layer3_outputs(429));
    layer4_outputs(6962) <= not(layer3_outputs(4006)) or (layer3_outputs(7117));
    layer4_outputs(6963) <= not(layer3_outputs(371)) or (layer3_outputs(3805));
    layer4_outputs(6964) <= layer3_outputs(3598);
    layer4_outputs(6965) <= not(layer3_outputs(7639));
    layer4_outputs(6966) <= (layer3_outputs(6271)) and not (layer3_outputs(5202));
    layer4_outputs(6967) <= not((layer3_outputs(1247)) or (layer3_outputs(7146)));
    layer4_outputs(6968) <= not(layer3_outputs(168));
    layer4_outputs(6969) <= (layer3_outputs(1914)) and not (layer3_outputs(1353));
    layer4_outputs(6970) <= layer3_outputs(765);
    layer4_outputs(6971) <= layer3_outputs(2125);
    layer4_outputs(6972) <= layer3_outputs(6581);
    layer4_outputs(6973) <= '1';
    layer4_outputs(6974) <= layer3_outputs(6068);
    layer4_outputs(6975) <= not(layer3_outputs(3135));
    layer4_outputs(6976) <= layer3_outputs(3143);
    layer4_outputs(6977) <= (layer3_outputs(3337)) xor (layer3_outputs(4892));
    layer4_outputs(6978) <= layer3_outputs(2887);
    layer4_outputs(6979) <= not(layer3_outputs(130)) or (layer3_outputs(7209));
    layer4_outputs(6980) <= not((layer3_outputs(3798)) and (layer3_outputs(6016)));
    layer4_outputs(6981) <= (layer3_outputs(3830)) and not (layer3_outputs(2973));
    layer4_outputs(6982) <= layer3_outputs(6352);
    layer4_outputs(6983) <= not((layer3_outputs(6163)) or (layer3_outputs(2606)));
    layer4_outputs(6984) <= not(layer3_outputs(5824));
    layer4_outputs(6985) <= not(layer3_outputs(1010));
    layer4_outputs(6986) <= not(layer3_outputs(2047));
    layer4_outputs(6987) <= not((layer3_outputs(5639)) or (layer3_outputs(7179)));
    layer4_outputs(6988) <= not(layer3_outputs(4216));
    layer4_outputs(6989) <= not(layer3_outputs(3108));
    layer4_outputs(6990) <= layer3_outputs(1183);
    layer4_outputs(6991) <= not((layer3_outputs(2718)) or (layer3_outputs(5051)));
    layer4_outputs(6992) <= not((layer3_outputs(4734)) or (layer3_outputs(6544)));
    layer4_outputs(6993) <= (layer3_outputs(6236)) and not (layer3_outputs(2765));
    layer4_outputs(6994) <= not(layer3_outputs(2698));
    layer4_outputs(6995) <= not(layer3_outputs(3965)) or (layer3_outputs(7186));
    layer4_outputs(6996) <= layer3_outputs(3507);
    layer4_outputs(6997) <= (layer3_outputs(6571)) and not (layer3_outputs(5255));
    layer4_outputs(6998) <= (layer3_outputs(7294)) and not (layer3_outputs(283));
    layer4_outputs(6999) <= not(layer3_outputs(3672));
    layer4_outputs(7000) <= not(layer3_outputs(2546)) or (layer3_outputs(48));
    layer4_outputs(7001) <= not(layer3_outputs(3140));
    layer4_outputs(7002) <= layer3_outputs(6575);
    layer4_outputs(7003) <= (layer3_outputs(4525)) and not (layer3_outputs(6993));
    layer4_outputs(7004) <= not(layer3_outputs(46)) or (layer3_outputs(5407));
    layer4_outputs(7005) <= (layer3_outputs(6440)) and not (layer3_outputs(6857));
    layer4_outputs(7006) <= not(layer3_outputs(6493));
    layer4_outputs(7007) <= layer3_outputs(59);
    layer4_outputs(7008) <= layer3_outputs(1910);
    layer4_outputs(7009) <= (layer3_outputs(124)) and not (layer3_outputs(37));
    layer4_outputs(7010) <= not(layer3_outputs(2618));
    layer4_outputs(7011) <= layer3_outputs(3041);
    layer4_outputs(7012) <= not(layer3_outputs(4726)) or (layer3_outputs(4814));
    layer4_outputs(7013) <= not((layer3_outputs(959)) and (layer3_outputs(2350)));
    layer4_outputs(7014) <= layer3_outputs(3611);
    layer4_outputs(7015) <= layer3_outputs(4883);
    layer4_outputs(7016) <= layer3_outputs(1838);
    layer4_outputs(7017) <= layer3_outputs(5704);
    layer4_outputs(7018) <= not(layer3_outputs(213));
    layer4_outputs(7019) <= layer3_outputs(2712);
    layer4_outputs(7020) <= layer3_outputs(6881);
    layer4_outputs(7021) <= layer3_outputs(3921);
    layer4_outputs(7022) <= layer3_outputs(4235);
    layer4_outputs(7023) <= '1';
    layer4_outputs(7024) <= layer3_outputs(2560);
    layer4_outputs(7025) <= (layer3_outputs(338)) or (layer3_outputs(1125));
    layer4_outputs(7026) <= '0';
    layer4_outputs(7027) <= (layer3_outputs(3588)) or (layer3_outputs(2578));
    layer4_outputs(7028) <= not(layer3_outputs(599)) or (layer3_outputs(2371));
    layer4_outputs(7029) <= not((layer3_outputs(4886)) and (layer3_outputs(6714)));
    layer4_outputs(7030) <= '1';
    layer4_outputs(7031) <= not(layer3_outputs(2581)) or (layer3_outputs(2208));
    layer4_outputs(7032) <= not(layer3_outputs(2429)) or (layer3_outputs(5110));
    layer4_outputs(7033) <= (layer3_outputs(4254)) and (layer3_outputs(2797));
    layer4_outputs(7034) <= not((layer3_outputs(1971)) and (layer3_outputs(1733)));
    layer4_outputs(7035) <= not(layer3_outputs(4008));
    layer4_outputs(7036) <= (layer3_outputs(4094)) and not (layer3_outputs(6782));
    layer4_outputs(7037) <= not(layer3_outputs(6342)) or (layer3_outputs(2759));
    layer4_outputs(7038) <= not(layer3_outputs(6890)) or (layer3_outputs(4945));
    layer4_outputs(7039) <= not((layer3_outputs(3426)) or (layer3_outputs(2046)));
    layer4_outputs(7040) <= '1';
    layer4_outputs(7041) <= (layer3_outputs(1410)) and (layer3_outputs(2656));
    layer4_outputs(7042) <= not(layer3_outputs(967)) or (layer3_outputs(3576));
    layer4_outputs(7043) <= not(layer3_outputs(5639)) or (layer3_outputs(400));
    layer4_outputs(7044) <= not((layer3_outputs(66)) and (layer3_outputs(5093)));
    layer4_outputs(7045) <= not((layer3_outputs(2971)) or (layer3_outputs(5212)));
    layer4_outputs(7046) <= not(layer3_outputs(6904));
    layer4_outputs(7047) <= not((layer3_outputs(1560)) xor (layer3_outputs(7403)));
    layer4_outputs(7048) <= layer3_outputs(6403);
    layer4_outputs(7049) <= (layer3_outputs(3429)) and (layer3_outputs(1241));
    layer4_outputs(7050) <= layer3_outputs(979);
    layer4_outputs(7051) <= (layer3_outputs(4135)) xor (layer3_outputs(2480));
    layer4_outputs(7052) <= (layer3_outputs(4843)) or (layer3_outputs(7347));
    layer4_outputs(7053) <= layer3_outputs(5191);
    layer4_outputs(7054) <= layer3_outputs(5631);
    layer4_outputs(7055) <= not((layer3_outputs(3425)) and (layer3_outputs(535)));
    layer4_outputs(7056) <= (layer3_outputs(7669)) or (layer3_outputs(441));
    layer4_outputs(7057) <= (layer3_outputs(3977)) and not (layer3_outputs(5461));
    layer4_outputs(7058) <= not(layer3_outputs(5650)) or (layer3_outputs(3026));
    layer4_outputs(7059) <= not((layer3_outputs(6100)) and (layer3_outputs(2326)));
    layer4_outputs(7060) <= layer3_outputs(62);
    layer4_outputs(7061) <= not(layer3_outputs(5704));
    layer4_outputs(7062) <= not((layer3_outputs(6546)) and (layer3_outputs(1791)));
    layer4_outputs(7063) <= layer3_outputs(2966);
    layer4_outputs(7064) <= layer3_outputs(7443);
    layer4_outputs(7065) <= layer3_outputs(1436);
    layer4_outputs(7066) <= layer3_outputs(6947);
    layer4_outputs(7067) <= layer3_outputs(7143);
    layer4_outputs(7068) <= (layer3_outputs(4337)) and not (layer3_outputs(881));
    layer4_outputs(7069) <= (layer3_outputs(7458)) or (layer3_outputs(195));
    layer4_outputs(7070) <= not(layer3_outputs(6738));
    layer4_outputs(7071) <= not((layer3_outputs(4930)) and (layer3_outputs(1771)));
    layer4_outputs(7072) <= (layer3_outputs(1914)) and (layer3_outputs(1538));
    layer4_outputs(7073) <= not(layer3_outputs(5253));
    layer4_outputs(7074) <= not(layer3_outputs(4218));
    layer4_outputs(7075) <= not((layer3_outputs(5459)) or (layer3_outputs(6550)));
    layer4_outputs(7076) <= layer3_outputs(5211);
    layer4_outputs(7077) <= layer3_outputs(4698);
    layer4_outputs(7078) <= not((layer3_outputs(1143)) or (layer3_outputs(3180)));
    layer4_outputs(7079) <= layer3_outputs(4973);
    layer4_outputs(7080) <= not((layer3_outputs(4309)) xor (layer3_outputs(1435)));
    layer4_outputs(7081) <= layer3_outputs(4094);
    layer4_outputs(7082) <= (layer3_outputs(6957)) xor (layer3_outputs(1949));
    layer4_outputs(7083) <= not((layer3_outputs(5107)) or (layer3_outputs(7029)));
    layer4_outputs(7084) <= not(layer3_outputs(5571));
    layer4_outputs(7085) <= not(layer3_outputs(519));
    layer4_outputs(7086) <= not(layer3_outputs(4506));
    layer4_outputs(7087) <= layer3_outputs(5981);
    layer4_outputs(7088) <= not(layer3_outputs(1850)) or (layer3_outputs(1218));
    layer4_outputs(7089) <= layer3_outputs(1544);
    layer4_outputs(7090) <= not(layer3_outputs(5481));
    layer4_outputs(7091) <= not(layer3_outputs(6658)) or (layer3_outputs(3052));
    layer4_outputs(7092) <= layer3_outputs(6337);
    layer4_outputs(7093) <= layer3_outputs(350);
    layer4_outputs(7094) <= layer3_outputs(7351);
    layer4_outputs(7095) <= (layer3_outputs(2080)) or (layer3_outputs(3818));
    layer4_outputs(7096) <= not((layer3_outputs(7340)) or (layer3_outputs(1984)));
    layer4_outputs(7097) <= not((layer3_outputs(1345)) or (layer3_outputs(6996)));
    layer4_outputs(7098) <= not(layer3_outputs(3797));
    layer4_outputs(7099) <= '1';
    layer4_outputs(7100) <= not(layer3_outputs(6495)) or (layer3_outputs(7070));
    layer4_outputs(7101) <= (layer3_outputs(3890)) or (layer3_outputs(4687));
    layer4_outputs(7102) <= not(layer3_outputs(4416)) or (layer3_outputs(3747));
    layer4_outputs(7103) <= '0';
    layer4_outputs(7104) <= layer3_outputs(6452);
    layer4_outputs(7105) <= not(layer3_outputs(1080));
    layer4_outputs(7106) <= (layer3_outputs(4892)) and not (layer3_outputs(7063));
    layer4_outputs(7107) <= (layer3_outputs(3228)) and not (layer3_outputs(6562));
    layer4_outputs(7108) <= layer3_outputs(5251);
    layer4_outputs(7109) <= layer3_outputs(2915);
    layer4_outputs(7110) <= (layer3_outputs(6887)) and not (layer3_outputs(3040));
    layer4_outputs(7111) <= not((layer3_outputs(6454)) and (layer3_outputs(6825)));
    layer4_outputs(7112) <= not(layer3_outputs(1400)) or (layer3_outputs(2828));
    layer4_outputs(7113) <= '1';
    layer4_outputs(7114) <= layer3_outputs(6697);
    layer4_outputs(7115) <= layer3_outputs(5398);
    layer4_outputs(7116) <= (layer3_outputs(5583)) and not (layer3_outputs(5732));
    layer4_outputs(7117) <= not((layer3_outputs(3208)) or (layer3_outputs(2702)));
    layer4_outputs(7118) <= (layer3_outputs(6010)) or (layer3_outputs(6025));
    layer4_outputs(7119) <= not(layer3_outputs(1232));
    layer4_outputs(7120) <= '0';
    layer4_outputs(7121) <= not((layer3_outputs(6126)) and (layer3_outputs(2039)));
    layer4_outputs(7122) <= not(layer3_outputs(5023));
    layer4_outputs(7123) <= layer3_outputs(330);
    layer4_outputs(7124) <= (layer3_outputs(6714)) and not (layer3_outputs(7594));
    layer4_outputs(7125) <= layer3_outputs(5137);
    layer4_outputs(7126) <= not(layer3_outputs(2795));
    layer4_outputs(7127) <= layer3_outputs(6422);
    layer4_outputs(7128) <= not(layer3_outputs(143));
    layer4_outputs(7129) <= not((layer3_outputs(1756)) or (layer3_outputs(7240)));
    layer4_outputs(7130) <= not(layer3_outputs(931));
    layer4_outputs(7131) <= layer3_outputs(4510);
    layer4_outputs(7132) <= not(layer3_outputs(1287));
    layer4_outputs(7133) <= not(layer3_outputs(916)) or (layer3_outputs(5703));
    layer4_outputs(7134) <= layer3_outputs(2464);
    layer4_outputs(7135) <= not((layer3_outputs(6043)) or (layer3_outputs(4167)));
    layer4_outputs(7136) <= (layer3_outputs(2207)) or (layer3_outputs(3684));
    layer4_outputs(7137) <= layer3_outputs(7454);
    layer4_outputs(7138) <= layer3_outputs(2783);
    layer4_outputs(7139) <= not(layer3_outputs(2661));
    layer4_outputs(7140) <= not((layer3_outputs(1053)) or (layer3_outputs(18)));
    layer4_outputs(7141) <= not(layer3_outputs(6948)) or (layer3_outputs(3967));
    layer4_outputs(7142) <= (layer3_outputs(4664)) xor (layer3_outputs(5334));
    layer4_outputs(7143) <= (layer3_outputs(7069)) xor (layer3_outputs(5766));
    layer4_outputs(7144) <= not(layer3_outputs(4239));
    layer4_outputs(7145) <= not(layer3_outputs(579)) or (layer3_outputs(121));
    layer4_outputs(7146) <= not(layer3_outputs(5908));
    layer4_outputs(7147) <= layer3_outputs(5102);
    layer4_outputs(7148) <= not(layer3_outputs(447)) or (layer3_outputs(7538));
    layer4_outputs(7149) <= (layer3_outputs(831)) or (layer3_outputs(386));
    layer4_outputs(7150) <= not(layer3_outputs(2031));
    layer4_outputs(7151) <= (layer3_outputs(4753)) and not (layer3_outputs(2260));
    layer4_outputs(7152) <= layer3_outputs(1709);
    layer4_outputs(7153) <= not(layer3_outputs(2596)) or (layer3_outputs(1454));
    layer4_outputs(7154) <= '0';
    layer4_outputs(7155) <= not(layer3_outputs(569));
    layer4_outputs(7156) <= (layer3_outputs(1314)) and (layer3_outputs(723));
    layer4_outputs(7157) <= not(layer3_outputs(5146));
    layer4_outputs(7158) <= layer3_outputs(3556);
    layer4_outputs(7159) <= (layer3_outputs(1720)) and not (layer3_outputs(6026));
    layer4_outputs(7160) <= (layer3_outputs(6058)) and not (layer3_outputs(7135));
    layer4_outputs(7161) <= not((layer3_outputs(925)) and (layer3_outputs(532)));
    layer4_outputs(7162) <= not(layer3_outputs(1573));
    layer4_outputs(7163) <= (layer3_outputs(6231)) and not (layer3_outputs(4463));
    layer4_outputs(7164) <= (layer3_outputs(3787)) and not (layer3_outputs(5944));
    layer4_outputs(7165) <= (layer3_outputs(5925)) and not (layer3_outputs(3659));
    layer4_outputs(7166) <= layer3_outputs(1247);
    layer4_outputs(7167) <= layer3_outputs(5246);
    layer4_outputs(7168) <= '1';
    layer4_outputs(7169) <= not(layer3_outputs(6750));
    layer4_outputs(7170) <= '0';
    layer4_outputs(7171) <= layer3_outputs(4622);
    layer4_outputs(7172) <= not(layer3_outputs(395)) or (layer3_outputs(6865));
    layer4_outputs(7173) <= '0';
    layer4_outputs(7174) <= not((layer3_outputs(1193)) xor (layer3_outputs(7086)));
    layer4_outputs(7175) <= not((layer3_outputs(6677)) or (layer3_outputs(6479)));
    layer4_outputs(7176) <= layer3_outputs(69);
    layer4_outputs(7177) <= not(layer3_outputs(3932)) or (layer3_outputs(6661));
    layer4_outputs(7178) <= layer3_outputs(1870);
    layer4_outputs(7179) <= layer3_outputs(7491);
    layer4_outputs(7180) <= not(layer3_outputs(7184)) or (layer3_outputs(4537));
    layer4_outputs(7181) <= layer3_outputs(1287);
    layer4_outputs(7182) <= (layer3_outputs(4479)) and not (layer3_outputs(4578));
    layer4_outputs(7183) <= (layer3_outputs(2398)) and not (layer3_outputs(3915));
    layer4_outputs(7184) <= not(layer3_outputs(5005));
    layer4_outputs(7185) <= (layer3_outputs(1005)) and not (layer3_outputs(3666));
    layer4_outputs(7186) <= layer3_outputs(2632);
    layer4_outputs(7187) <= layer3_outputs(6652);
    layer4_outputs(7188) <= layer3_outputs(4273);
    layer4_outputs(7189) <= not(layer3_outputs(3235)) or (layer3_outputs(1687));
    layer4_outputs(7190) <= (layer3_outputs(2822)) and not (layer3_outputs(4623));
    layer4_outputs(7191) <= not(layer3_outputs(3889));
    layer4_outputs(7192) <= not(layer3_outputs(7004)) or (layer3_outputs(4267));
    layer4_outputs(7193) <= not(layer3_outputs(2029)) or (layer3_outputs(85));
    layer4_outputs(7194) <= not(layer3_outputs(2091)) or (layer3_outputs(679));
    layer4_outputs(7195) <= (layer3_outputs(1682)) and (layer3_outputs(6587));
    layer4_outputs(7196) <= not(layer3_outputs(6118)) or (layer3_outputs(6734));
    layer4_outputs(7197) <= '1';
    layer4_outputs(7198) <= (layer3_outputs(3205)) xor (layer3_outputs(3780));
    layer4_outputs(7199) <= not((layer3_outputs(658)) and (layer3_outputs(887)));
    layer4_outputs(7200) <= (layer3_outputs(3061)) and not (layer3_outputs(6283));
    layer4_outputs(7201) <= not(layer3_outputs(7416)) or (layer3_outputs(256));
    layer4_outputs(7202) <= (layer3_outputs(2601)) or (layer3_outputs(1575));
    layer4_outputs(7203) <= '0';
    layer4_outputs(7204) <= layer3_outputs(1009);
    layer4_outputs(7205) <= (layer3_outputs(1911)) xor (layer3_outputs(3540));
    layer4_outputs(7206) <= (layer3_outputs(443)) and not (layer3_outputs(76));
    layer4_outputs(7207) <= not(layer3_outputs(1945));
    layer4_outputs(7208) <= layer3_outputs(2605);
    layer4_outputs(7209) <= not((layer3_outputs(3924)) xor (layer3_outputs(3471)));
    layer4_outputs(7210) <= not((layer3_outputs(1761)) or (layer3_outputs(6285)));
    layer4_outputs(7211) <= (layer3_outputs(390)) and not (layer3_outputs(4975));
    layer4_outputs(7212) <= not((layer3_outputs(1331)) or (layer3_outputs(2512)));
    layer4_outputs(7213) <= not(layer3_outputs(6965));
    layer4_outputs(7214) <= not((layer3_outputs(2410)) and (layer3_outputs(6793)));
    layer4_outputs(7215) <= not(layer3_outputs(2700));
    layer4_outputs(7216) <= (layer3_outputs(4459)) and not (layer3_outputs(3509));
    layer4_outputs(7217) <= (layer3_outputs(4103)) and not (layer3_outputs(2265));
    layer4_outputs(7218) <= (layer3_outputs(4076)) and not (layer3_outputs(2747));
    layer4_outputs(7219) <= layer3_outputs(3841);
    layer4_outputs(7220) <= not((layer3_outputs(5359)) or (layer3_outputs(4177)));
    layer4_outputs(7221) <= layer3_outputs(2496);
    layer4_outputs(7222) <= not(layer3_outputs(7131));
    layer4_outputs(7223) <= (layer3_outputs(2659)) and (layer3_outputs(7672));
    layer4_outputs(7224) <= (layer3_outputs(6653)) and not (layer3_outputs(1976));
    layer4_outputs(7225) <= not((layer3_outputs(7289)) xor (layer3_outputs(3260)));
    layer4_outputs(7226) <= (layer3_outputs(983)) or (layer3_outputs(3046));
    layer4_outputs(7227) <= not(layer3_outputs(4312));
    layer4_outputs(7228) <= not((layer3_outputs(2320)) or (layer3_outputs(2511)));
    layer4_outputs(7229) <= '1';
    layer4_outputs(7230) <= not(layer3_outputs(2986));
    layer4_outputs(7231) <= (layer3_outputs(3508)) and (layer3_outputs(6040));
    layer4_outputs(7232) <= layer3_outputs(2035);
    layer4_outputs(7233) <= not(layer3_outputs(2844));
    layer4_outputs(7234) <= (layer3_outputs(2325)) and not (layer3_outputs(660));
    layer4_outputs(7235) <= layer3_outputs(414);
    layer4_outputs(7236) <= not(layer3_outputs(5806));
    layer4_outputs(7237) <= (layer3_outputs(1199)) and not (layer3_outputs(6448));
    layer4_outputs(7238) <= not(layer3_outputs(2674));
    layer4_outputs(7239) <= layer3_outputs(2120);
    layer4_outputs(7240) <= not(layer3_outputs(4036)) or (layer3_outputs(7022));
    layer4_outputs(7241) <= not(layer3_outputs(5859)) or (layer3_outputs(3601));
    layer4_outputs(7242) <= layer3_outputs(745);
    layer4_outputs(7243) <= not((layer3_outputs(6347)) or (layer3_outputs(5821)));
    layer4_outputs(7244) <= layer3_outputs(4088);
    layer4_outputs(7245) <= (layer3_outputs(1166)) and not (layer3_outputs(507));
    layer4_outputs(7246) <= not(layer3_outputs(7216)) or (layer3_outputs(4941));
    layer4_outputs(7247) <= not((layer3_outputs(7138)) or (layer3_outputs(4382)));
    layer4_outputs(7248) <= (layer3_outputs(4636)) and not (layer3_outputs(5270));
    layer4_outputs(7249) <= layer3_outputs(4438);
    layer4_outputs(7250) <= (layer3_outputs(133)) and not (layer3_outputs(3996));
    layer4_outputs(7251) <= not(layer3_outputs(824)) or (layer3_outputs(1401));
    layer4_outputs(7252) <= not((layer3_outputs(7091)) or (layer3_outputs(934)));
    layer4_outputs(7253) <= not((layer3_outputs(7242)) or (layer3_outputs(3664)));
    layer4_outputs(7254) <= (layer3_outputs(3341)) or (layer3_outputs(7355));
    layer4_outputs(7255) <= layer3_outputs(6780);
    layer4_outputs(7256) <= layer3_outputs(3483);
    layer4_outputs(7257) <= (layer3_outputs(6749)) and not (layer3_outputs(5902));
    layer4_outputs(7258) <= not((layer3_outputs(2224)) or (layer3_outputs(4018)));
    layer4_outputs(7259) <= '1';
    layer4_outputs(7260) <= not(layer3_outputs(2492)) or (layer3_outputs(3253));
    layer4_outputs(7261) <= not((layer3_outputs(7445)) xor (layer3_outputs(401)));
    layer4_outputs(7262) <= not(layer3_outputs(2996)) or (layer3_outputs(766));
    layer4_outputs(7263) <= not(layer3_outputs(4699));
    layer4_outputs(7264) <= (layer3_outputs(7139)) and not (layer3_outputs(2167));
    layer4_outputs(7265) <= (layer3_outputs(6368)) or (layer3_outputs(3420));
    layer4_outputs(7266) <= not(layer3_outputs(5268));
    layer4_outputs(7267) <= not(layer3_outputs(2541));
    layer4_outputs(7268) <= (layer3_outputs(7094)) and not (layer3_outputs(5285));
    layer4_outputs(7269) <= not(layer3_outputs(2600));
    layer4_outputs(7270) <= (layer3_outputs(3537)) xor (layer3_outputs(4142));
    layer4_outputs(7271) <= layer3_outputs(3414);
    layer4_outputs(7272) <= layer3_outputs(3581);
    layer4_outputs(7273) <= layer3_outputs(7619);
    layer4_outputs(7274) <= (layer3_outputs(1526)) or (layer3_outputs(4653));
    layer4_outputs(7275) <= not(layer3_outputs(4762)) or (layer3_outputs(7182));
    layer4_outputs(7276) <= (layer3_outputs(4989)) xor (layer3_outputs(2030));
    layer4_outputs(7277) <= not((layer3_outputs(1860)) and (layer3_outputs(7026)));
    layer4_outputs(7278) <= layer3_outputs(342);
    layer4_outputs(7279) <= layer3_outputs(4576);
    layer4_outputs(7280) <= (layer3_outputs(7395)) and not (layer3_outputs(4887));
    layer4_outputs(7281) <= (layer3_outputs(4712)) or (layer3_outputs(3533));
    layer4_outputs(7282) <= not(layer3_outputs(558)) or (layer3_outputs(6781));
    layer4_outputs(7283) <= not(layer3_outputs(1936));
    layer4_outputs(7284) <= not((layer3_outputs(1149)) or (layer3_outputs(2608)));
    layer4_outputs(7285) <= (layer3_outputs(5810)) and not (layer3_outputs(1898));
    layer4_outputs(7286) <= layer3_outputs(5401);
    layer4_outputs(7287) <= not((layer3_outputs(7198)) and (layer3_outputs(4527)));
    layer4_outputs(7288) <= (layer3_outputs(6345)) and not (layer3_outputs(292));
    layer4_outputs(7289) <= (layer3_outputs(3946)) and not (layer3_outputs(7336));
    layer4_outputs(7290) <= not(layer3_outputs(4559));
    layer4_outputs(7291) <= (layer3_outputs(5748)) and not (layer3_outputs(1147));
    layer4_outputs(7292) <= (layer3_outputs(7575)) and (layer3_outputs(5103));
    layer4_outputs(7293) <= layer3_outputs(2180);
    layer4_outputs(7294) <= (layer3_outputs(716)) and not (layer3_outputs(4371));
    layer4_outputs(7295) <= (layer3_outputs(7420)) or (layer3_outputs(5224));
    layer4_outputs(7296) <= layer3_outputs(2263);
    layer4_outputs(7297) <= layer3_outputs(5498);
    layer4_outputs(7298) <= '1';
    layer4_outputs(7299) <= (layer3_outputs(5188)) and not (layer3_outputs(4492));
    layer4_outputs(7300) <= (layer3_outputs(4531)) and (layer3_outputs(3994));
    layer4_outputs(7301) <= (layer3_outputs(4139)) and not (layer3_outputs(5111));
    layer4_outputs(7302) <= layer3_outputs(3853);
    layer4_outputs(7303) <= (layer3_outputs(4627)) and (layer3_outputs(4106));
    layer4_outputs(7304) <= layer3_outputs(1407);
    layer4_outputs(7305) <= (layer3_outputs(1409)) and not (layer3_outputs(5435));
    layer4_outputs(7306) <= layer3_outputs(1350);
    layer4_outputs(7307) <= not(layer3_outputs(7099));
    layer4_outputs(7308) <= layer3_outputs(4534);
    layer4_outputs(7309) <= layer3_outputs(2252);
    layer4_outputs(7310) <= (layer3_outputs(5965)) and not (layer3_outputs(6215));
    layer4_outputs(7311) <= not(layer3_outputs(4949));
    layer4_outputs(7312) <= not((layer3_outputs(4479)) and (layer3_outputs(5106)));
    layer4_outputs(7313) <= not(layer3_outputs(5760));
    layer4_outputs(7314) <= not(layer3_outputs(4067));
    layer4_outputs(7315) <= not(layer3_outputs(4070));
    layer4_outputs(7316) <= not(layer3_outputs(60)) or (layer3_outputs(4997));
    layer4_outputs(7317) <= not(layer3_outputs(4738));
    layer4_outputs(7318) <= layer3_outputs(3924);
    layer4_outputs(7319) <= not(layer3_outputs(2459));
    layer4_outputs(7320) <= not((layer3_outputs(5053)) and (layer3_outputs(4906)));
    layer4_outputs(7321) <= not(layer3_outputs(4966));
    layer4_outputs(7322) <= not((layer3_outputs(6932)) xor (layer3_outputs(1940)));
    layer4_outputs(7323) <= (layer3_outputs(6511)) and (layer3_outputs(5536));
    layer4_outputs(7324) <= layer3_outputs(5789);
    layer4_outputs(7325) <= layer3_outputs(6208);
    layer4_outputs(7326) <= layer3_outputs(4249);
    layer4_outputs(7327) <= (layer3_outputs(2852)) xor (layer3_outputs(3081));
    layer4_outputs(7328) <= not(layer3_outputs(6593)) or (layer3_outputs(4010));
    layer4_outputs(7329) <= (layer3_outputs(3406)) and not (layer3_outputs(4516));
    layer4_outputs(7330) <= '1';
    layer4_outputs(7331) <= layer3_outputs(5933);
    layer4_outputs(7332) <= not(layer3_outputs(1632));
    layer4_outputs(7333) <= not(layer3_outputs(1996));
    layer4_outputs(7334) <= not(layer3_outputs(1757));
    layer4_outputs(7335) <= (layer3_outputs(6374)) and (layer3_outputs(4844));
    layer4_outputs(7336) <= not(layer3_outputs(3929));
    layer4_outputs(7337) <= not(layer3_outputs(1885));
    layer4_outputs(7338) <= (layer3_outputs(1493)) and (layer3_outputs(4167));
    layer4_outputs(7339) <= not(layer3_outputs(1736));
    layer4_outputs(7340) <= '1';
    layer4_outputs(7341) <= not(layer3_outputs(478));
    layer4_outputs(7342) <= not((layer3_outputs(716)) and (layer3_outputs(1952)));
    layer4_outputs(7343) <= not((layer3_outputs(7145)) or (layer3_outputs(5470)));
    layer4_outputs(7344) <= layer3_outputs(3064);
    layer4_outputs(7345) <= (layer3_outputs(1408)) and (layer3_outputs(4674));
    layer4_outputs(7346) <= (layer3_outputs(4550)) and not (layer3_outputs(2617));
    layer4_outputs(7347) <= layer3_outputs(6082);
    layer4_outputs(7348) <= (layer3_outputs(2009)) xor (layer3_outputs(3387));
    layer4_outputs(7349) <= not(layer3_outputs(586));
    layer4_outputs(7350) <= '0';
    layer4_outputs(7351) <= layer3_outputs(4862);
    layer4_outputs(7352) <= layer3_outputs(394);
    layer4_outputs(7353) <= not((layer3_outputs(2323)) and (layer3_outputs(336)));
    layer4_outputs(7354) <= (layer3_outputs(4969)) and (layer3_outputs(4901));
    layer4_outputs(7355) <= not(layer3_outputs(2678));
    layer4_outputs(7356) <= (layer3_outputs(2604)) and not (layer3_outputs(1653));
    layer4_outputs(7357) <= (layer3_outputs(1726)) xor (layer3_outputs(5088));
    layer4_outputs(7358) <= '1';
    layer4_outputs(7359) <= not(layer3_outputs(6526)) or (layer3_outputs(6604));
    layer4_outputs(7360) <= not(layer3_outputs(3500)) or (layer3_outputs(5059));
    layer4_outputs(7361) <= (layer3_outputs(5243)) and not (layer3_outputs(3843));
    layer4_outputs(7362) <= (layer3_outputs(6598)) and not (layer3_outputs(5454));
    layer4_outputs(7363) <= '0';
    layer4_outputs(7364) <= layer3_outputs(4306);
    layer4_outputs(7365) <= not(layer3_outputs(7572));
    layer4_outputs(7366) <= not(layer3_outputs(366)) or (layer3_outputs(5324));
    layer4_outputs(7367) <= (layer3_outputs(7261)) and not (layer3_outputs(6393));
    layer4_outputs(7368) <= (layer3_outputs(3035)) xor (layer3_outputs(3926));
    layer4_outputs(7369) <= '0';
    layer4_outputs(7370) <= (layer3_outputs(5454)) and not (layer3_outputs(1448));
    layer4_outputs(7371) <= layer3_outputs(6336);
    layer4_outputs(7372) <= (layer3_outputs(3777)) and not (layer3_outputs(1912));
    layer4_outputs(7373) <= not(layer3_outputs(237));
    layer4_outputs(7374) <= (layer3_outputs(3807)) and not (layer3_outputs(4277));
    layer4_outputs(7375) <= layer3_outputs(5489);
    layer4_outputs(7376) <= not(layer3_outputs(4105));
    layer4_outputs(7377) <= '1';
    layer4_outputs(7378) <= layer3_outputs(6960);
    layer4_outputs(7379) <= (layer3_outputs(1082)) and (layer3_outputs(5585));
    layer4_outputs(7380) <= not(layer3_outputs(505));
    layer4_outputs(7381) <= not(layer3_outputs(7554));
    layer4_outputs(7382) <= (layer3_outputs(7132)) or (layer3_outputs(809));
    layer4_outputs(7383) <= not((layer3_outputs(4257)) xor (layer3_outputs(7255)));
    layer4_outputs(7384) <= not(layer3_outputs(487));
    layer4_outputs(7385) <= not(layer3_outputs(2780)) or (layer3_outputs(7110));
    layer4_outputs(7386) <= '0';
    layer4_outputs(7387) <= layer3_outputs(5699);
    layer4_outputs(7388) <= (layer3_outputs(1483)) and not (layer3_outputs(2936));
    layer4_outputs(7389) <= not(layer3_outputs(5971));
    layer4_outputs(7390) <= layer3_outputs(868);
    layer4_outputs(7391) <= (layer3_outputs(4073)) and not (layer3_outputs(435));
    layer4_outputs(7392) <= layer3_outputs(2527);
    layer4_outputs(7393) <= layer3_outputs(5863);
    layer4_outputs(7394) <= layer3_outputs(3120);
    layer4_outputs(7395) <= (layer3_outputs(3226)) and (layer3_outputs(7173));
    layer4_outputs(7396) <= not(layer3_outputs(5056));
    layer4_outputs(7397) <= not(layer3_outputs(77));
    layer4_outputs(7398) <= (layer3_outputs(7089)) or (layer3_outputs(7060));
    layer4_outputs(7399) <= not(layer3_outputs(324));
    layer4_outputs(7400) <= layer3_outputs(715);
    layer4_outputs(7401) <= not(layer3_outputs(4385));
    layer4_outputs(7402) <= not(layer3_outputs(5480));
    layer4_outputs(7403) <= not(layer3_outputs(5402));
    layer4_outputs(7404) <= not(layer3_outputs(4645));
    layer4_outputs(7405) <= not((layer3_outputs(5526)) or (layer3_outputs(2472)));
    layer4_outputs(7406) <= (layer3_outputs(7638)) xor (layer3_outputs(6519));
    layer4_outputs(7407) <= layer3_outputs(3011);
    layer4_outputs(7408) <= (layer3_outputs(3615)) and not (layer3_outputs(4728));
    layer4_outputs(7409) <= not(layer3_outputs(1838)) or (layer3_outputs(5829));
    layer4_outputs(7410) <= layer3_outputs(5172);
    layer4_outputs(7411) <= not(layer3_outputs(1577)) or (layer3_outputs(2444));
    layer4_outputs(7412) <= not((layer3_outputs(6372)) and (layer3_outputs(1548)));
    layer4_outputs(7413) <= (layer3_outputs(1126)) and not (layer3_outputs(6052));
    layer4_outputs(7414) <= not(layer3_outputs(92)) or (layer3_outputs(2066));
    layer4_outputs(7415) <= not(layer3_outputs(5365)) or (layer3_outputs(5215));
    layer4_outputs(7416) <= not(layer3_outputs(1531));
    layer4_outputs(7417) <= layer3_outputs(4866);
    layer4_outputs(7418) <= not(layer3_outputs(7597));
    layer4_outputs(7419) <= layer3_outputs(3769);
    layer4_outputs(7420) <= not((layer3_outputs(3702)) or (layer3_outputs(3904)));
    layer4_outputs(7421) <= (layer3_outputs(5138)) and not (layer3_outputs(5506));
    layer4_outputs(7422) <= not((layer3_outputs(2693)) xor (layer3_outputs(748)));
    layer4_outputs(7423) <= layer3_outputs(2216);
    layer4_outputs(7424) <= not(layer3_outputs(5537));
    layer4_outputs(7425) <= not(layer3_outputs(3372));
    layer4_outputs(7426) <= not(layer3_outputs(7547)) or (layer3_outputs(1459));
    layer4_outputs(7427) <= not(layer3_outputs(1740)) or (layer3_outputs(3855));
    layer4_outputs(7428) <= (layer3_outputs(7598)) and not (layer3_outputs(4598));
    layer4_outputs(7429) <= layer3_outputs(1014);
    layer4_outputs(7430) <= (layer3_outputs(1141)) and not (layer3_outputs(6528));
    layer4_outputs(7431) <= '1';
    layer4_outputs(7432) <= not((layer3_outputs(4023)) and (layer3_outputs(344)));
    layer4_outputs(7433) <= not(layer3_outputs(6672));
    layer4_outputs(7434) <= not(layer3_outputs(6651));
    layer4_outputs(7435) <= (layer3_outputs(1541)) and not (layer3_outputs(5322));
    layer4_outputs(7436) <= not(layer3_outputs(6958));
    layer4_outputs(7437) <= (layer3_outputs(4933)) or (layer3_outputs(628));
    layer4_outputs(7438) <= not((layer3_outputs(3918)) or (layer3_outputs(6886)));
    layer4_outputs(7439) <= not(layer3_outputs(3555));
    layer4_outputs(7440) <= not(layer3_outputs(5140)) or (layer3_outputs(5225));
    layer4_outputs(7441) <= not(layer3_outputs(941));
    layer4_outputs(7442) <= (layer3_outputs(4332)) and not (layer3_outputs(2959));
    layer4_outputs(7443) <= '0';
    layer4_outputs(7444) <= (layer3_outputs(3579)) and not (layer3_outputs(6870));
    layer4_outputs(7445) <= (layer3_outputs(6475)) xor (layer3_outputs(3229));
    layer4_outputs(7446) <= not(layer3_outputs(932)) or (layer3_outputs(5525));
    layer4_outputs(7447) <= layer3_outputs(631);
    layer4_outputs(7448) <= not(layer3_outputs(3941)) or (layer3_outputs(4647));
    layer4_outputs(7449) <= not(layer3_outputs(7305));
    layer4_outputs(7450) <= (layer3_outputs(6467)) and not (layer3_outputs(692));
    layer4_outputs(7451) <= not((layer3_outputs(3044)) and (layer3_outputs(6456)));
    layer4_outputs(7452) <= not(layer3_outputs(755));
    layer4_outputs(7453) <= layer3_outputs(2042);
    layer4_outputs(7454) <= layer3_outputs(5082);
    layer4_outputs(7455) <= (layer3_outputs(6769)) or (layer3_outputs(1587));
    layer4_outputs(7456) <= not(layer3_outputs(5982)) or (layer3_outputs(5434));
    layer4_outputs(7457) <= layer3_outputs(51);
    layer4_outputs(7458) <= not((layer3_outputs(7293)) or (layer3_outputs(2587)));
    layer4_outputs(7459) <= '0';
    layer4_outputs(7460) <= not((layer3_outputs(1172)) xor (layer3_outputs(5700)));
    layer4_outputs(7461) <= '0';
    layer4_outputs(7462) <= not((layer3_outputs(3085)) and (layer3_outputs(7570)));
    layer4_outputs(7463) <= not((layer3_outputs(4981)) xor (layer3_outputs(4249)));
    layer4_outputs(7464) <= not(layer3_outputs(2734));
    layer4_outputs(7465) <= (layer3_outputs(7134)) and not (layer3_outputs(4017));
    layer4_outputs(7466) <= not((layer3_outputs(3966)) xor (layer3_outputs(6591)));
    layer4_outputs(7467) <= '0';
    layer4_outputs(7468) <= not((layer3_outputs(1784)) xor (layer3_outputs(517)));
    layer4_outputs(7469) <= '1';
    layer4_outputs(7470) <= not(layer3_outputs(7428));
    layer4_outputs(7471) <= not(layer3_outputs(2721)) or (layer3_outputs(7145));
    layer4_outputs(7472) <= (layer3_outputs(5450)) and (layer3_outputs(1322));
    layer4_outputs(7473) <= not(layer3_outputs(3548)) or (layer3_outputs(6737));
    layer4_outputs(7474) <= not(layer3_outputs(4032));
    layer4_outputs(7475) <= (layer3_outputs(6422)) and (layer3_outputs(354));
    layer4_outputs(7476) <= (layer3_outputs(3788)) and not (layer3_outputs(1558));
    layer4_outputs(7477) <= layer3_outputs(2753);
    layer4_outputs(7478) <= not(layer3_outputs(6142));
    layer4_outputs(7479) <= (layer3_outputs(1625)) and not (layer3_outputs(3399));
    layer4_outputs(7480) <= layer3_outputs(3313);
    layer4_outputs(7481) <= not((layer3_outputs(5068)) and (layer3_outputs(6599)));
    layer4_outputs(7482) <= (layer3_outputs(5741)) and not (layer3_outputs(1240));
    layer4_outputs(7483) <= not(layer3_outputs(6942));
    layer4_outputs(7484) <= not(layer3_outputs(6399)) or (layer3_outputs(2854));
    layer4_outputs(7485) <= not((layer3_outputs(4431)) xor (layer3_outputs(4723)));
    layer4_outputs(7486) <= not(layer3_outputs(2463));
    layer4_outputs(7487) <= not((layer3_outputs(5647)) or (layer3_outputs(6337)));
    layer4_outputs(7488) <= not(layer3_outputs(4811)) or (layer3_outputs(355));
    layer4_outputs(7489) <= not(layer3_outputs(3084));
    layer4_outputs(7490) <= layer3_outputs(4580);
    layer4_outputs(7491) <= (layer3_outputs(163)) and not (layer3_outputs(815));
    layer4_outputs(7492) <= layer3_outputs(6083);
    layer4_outputs(7493) <= layer3_outputs(1387);
    layer4_outputs(7494) <= not((layer3_outputs(6099)) or (layer3_outputs(4713)));
    layer4_outputs(7495) <= not(layer3_outputs(3199));
    layer4_outputs(7496) <= '0';
    layer4_outputs(7497) <= layer3_outputs(1368);
    layer4_outputs(7498) <= not(layer3_outputs(1545));
    layer4_outputs(7499) <= not((layer3_outputs(4121)) and (layer3_outputs(7628)));
    layer4_outputs(7500) <= '1';
    layer4_outputs(7501) <= layer3_outputs(7329);
    layer4_outputs(7502) <= (layer3_outputs(6088)) xor (layer3_outputs(6973));
    layer4_outputs(7503) <= layer3_outputs(3899);
    layer4_outputs(7504) <= not((layer3_outputs(1701)) or (layer3_outputs(2407)));
    layer4_outputs(7505) <= not(layer3_outputs(4370));
    layer4_outputs(7506) <= (layer3_outputs(1480)) and not (layer3_outputs(5728));
    layer4_outputs(7507) <= layer3_outputs(5833);
    layer4_outputs(7508) <= layer3_outputs(7587);
    layer4_outputs(7509) <= not(layer3_outputs(3652));
    layer4_outputs(7510) <= not(layer3_outputs(7444));
    layer4_outputs(7511) <= (layer3_outputs(4024)) and (layer3_outputs(3359));
    layer4_outputs(7512) <= layer3_outputs(2885);
    layer4_outputs(7513) <= (layer3_outputs(1787)) and not (layer3_outputs(2282));
    layer4_outputs(7514) <= (layer3_outputs(4166)) and not (layer3_outputs(6395));
    layer4_outputs(7515) <= not(layer3_outputs(1698));
    layer4_outputs(7516) <= '0';
    layer4_outputs(7517) <= layer3_outputs(101);
    layer4_outputs(7518) <= (layer3_outputs(5722)) and not (layer3_outputs(4669));
    layer4_outputs(7519) <= '1';
    layer4_outputs(7520) <= layer3_outputs(7232);
    layer4_outputs(7521) <= not(layer3_outputs(4424));
    layer4_outputs(7522) <= not((layer3_outputs(6709)) or (layer3_outputs(5475)));
    layer4_outputs(7523) <= layer3_outputs(5218);
    layer4_outputs(7524) <= (layer3_outputs(1348)) and not (layer3_outputs(5501));
    layer4_outputs(7525) <= layer3_outputs(7663);
    layer4_outputs(7526) <= (layer3_outputs(849)) and not (layer3_outputs(3706));
    layer4_outputs(7527) <= not(layer3_outputs(4970)) or (layer3_outputs(4340));
    layer4_outputs(7528) <= layer3_outputs(5561);
    layer4_outputs(7529) <= (layer3_outputs(4214)) or (layer3_outputs(3116));
    layer4_outputs(7530) <= layer3_outputs(7060);
    layer4_outputs(7531) <= not(layer3_outputs(5616));
    layer4_outputs(7532) <= not(layer3_outputs(5343)) or (layer3_outputs(7469));
    layer4_outputs(7533) <= '0';
    layer4_outputs(7534) <= layer3_outputs(6229);
    layer4_outputs(7535) <= layer3_outputs(3692);
    layer4_outputs(7536) <= not((layer3_outputs(1529)) and (layer3_outputs(3942)));
    layer4_outputs(7537) <= not(layer3_outputs(7044)) or (layer3_outputs(170));
    layer4_outputs(7538) <= (layer3_outputs(4654)) and (layer3_outputs(5706));
    layer4_outputs(7539) <= not(layer3_outputs(3094));
    layer4_outputs(7540) <= layer3_outputs(5410);
    layer4_outputs(7541) <= not(layer3_outputs(6679)) or (layer3_outputs(4648));
    layer4_outputs(7542) <= not(layer3_outputs(4545)) or (layer3_outputs(2483));
    layer4_outputs(7543) <= (layer3_outputs(1144)) and (layer3_outputs(461));
    layer4_outputs(7544) <= not(layer3_outputs(6578));
    layer4_outputs(7545) <= not((layer3_outputs(4413)) or (layer3_outputs(5854)));
    layer4_outputs(7546) <= (layer3_outputs(5738)) and not (layer3_outputs(7519));
    layer4_outputs(7547) <= not(layer3_outputs(3086));
    layer4_outputs(7548) <= (layer3_outputs(6438)) and not (layer3_outputs(7502));
    layer4_outputs(7549) <= not((layer3_outputs(1766)) and (layer3_outputs(2017)));
    layer4_outputs(7550) <= not(layer3_outputs(5708)) or (layer3_outputs(847));
    layer4_outputs(7551) <= not(layer3_outputs(2340));
    layer4_outputs(7552) <= layer3_outputs(909);
    layer4_outputs(7553) <= (layer3_outputs(3861)) and (layer3_outputs(197));
    layer4_outputs(7554) <= layer3_outputs(3898);
    layer4_outputs(7555) <= layer3_outputs(5598);
    layer4_outputs(7556) <= layer3_outputs(297);
    layer4_outputs(7557) <= (layer3_outputs(5558)) xor (layer3_outputs(3590));
    layer4_outputs(7558) <= layer3_outputs(2909);
    layer4_outputs(7559) <= (layer3_outputs(866)) and (layer3_outputs(4297));
    layer4_outputs(7560) <= (layer3_outputs(3897)) and not (layer3_outputs(234));
    layer4_outputs(7561) <= layer3_outputs(7208);
    layer4_outputs(7562) <= not((layer3_outputs(3118)) xor (layer3_outputs(3071)));
    layer4_outputs(7563) <= not(layer3_outputs(5961));
    layer4_outputs(7564) <= '0';
    layer4_outputs(7565) <= layer3_outputs(6919);
    layer4_outputs(7566) <= (layer3_outputs(6136)) xor (layer3_outputs(6406));
    layer4_outputs(7567) <= (layer3_outputs(3789)) xor (layer3_outputs(2295));
    layer4_outputs(7568) <= not(layer3_outputs(3709));
    layer4_outputs(7569) <= not((layer3_outputs(1865)) and (layer3_outputs(6582)));
    layer4_outputs(7570) <= not(layer3_outputs(1493)) or (layer3_outputs(5784));
    layer4_outputs(7571) <= not(layer3_outputs(3238));
    layer4_outputs(7572) <= not(layer3_outputs(2043));
    layer4_outputs(7573) <= not(layer3_outputs(7479));
    layer4_outputs(7574) <= not((layer3_outputs(1392)) or (layer3_outputs(1595)));
    layer4_outputs(7575) <= not(layer3_outputs(5338)) or (layer3_outputs(3730));
    layer4_outputs(7576) <= layer3_outputs(2453);
    layer4_outputs(7577) <= not(layer3_outputs(2914));
    layer4_outputs(7578) <= '0';
    layer4_outputs(7579) <= (layer3_outputs(2071)) and not (layer3_outputs(1905));
    layer4_outputs(7580) <= (layer3_outputs(6820)) or (layer3_outputs(1141));
    layer4_outputs(7581) <= '0';
    layer4_outputs(7582) <= layer3_outputs(2781);
    layer4_outputs(7583) <= not(layer3_outputs(6636));
    layer4_outputs(7584) <= (layer3_outputs(1297)) and not (layer3_outputs(1486));
    layer4_outputs(7585) <= not(layer3_outputs(1700)) or (layer3_outputs(3650));
    layer4_outputs(7586) <= layer3_outputs(1655);
    layer4_outputs(7587) <= not(layer3_outputs(2584));
    layer4_outputs(7588) <= not((layer3_outputs(2559)) and (layer3_outputs(7084)));
    layer4_outputs(7589) <= not(layer3_outputs(5301)) or (layer3_outputs(5392));
    layer4_outputs(7590) <= layer3_outputs(3398);
    layer4_outputs(7591) <= not(layer3_outputs(6588));
    layer4_outputs(7592) <= (layer3_outputs(2074)) or (layer3_outputs(2202));
    layer4_outputs(7593) <= not(layer3_outputs(7097)) or (layer3_outputs(5403));
    layer4_outputs(7594) <= layer3_outputs(7471);
    layer4_outputs(7595) <= not(layer3_outputs(1401));
    layer4_outputs(7596) <= layer3_outputs(88);
    layer4_outputs(7597) <= layer3_outputs(674);
    layer4_outputs(7598) <= layer3_outputs(2075);
    layer4_outputs(7599) <= layer3_outputs(3584);
    layer4_outputs(7600) <= not((layer3_outputs(6432)) or (layer3_outputs(54)));
    layer4_outputs(7601) <= not((layer3_outputs(202)) or (layer3_outputs(6113)));
    layer4_outputs(7602) <= layer3_outputs(5836);
    layer4_outputs(7603) <= layer3_outputs(6296);
    layer4_outputs(7604) <= layer3_outputs(5160);
    layer4_outputs(7605) <= not(layer3_outputs(3641)) or (layer3_outputs(3419));
    layer4_outputs(7606) <= not(layer3_outputs(7190)) or (layer3_outputs(1888));
    layer4_outputs(7607) <= not((layer3_outputs(909)) or (layer3_outputs(310)));
    layer4_outputs(7608) <= not(layer3_outputs(2724));
    layer4_outputs(7609) <= layer3_outputs(455);
    layer4_outputs(7610) <= '0';
    layer4_outputs(7611) <= layer3_outputs(2025);
    layer4_outputs(7612) <= not(layer3_outputs(1740));
    layer4_outputs(7613) <= layer3_outputs(2945);
    layer4_outputs(7614) <= not(layer3_outputs(6992));
    layer4_outputs(7615) <= (layer3_outputs(7580)) and (layer3_outputs(488));
    layer4_outputs(7616) <= layer3_outputs(5654);
    layer4_outputs(7617) <= layer3_outputs(5035);
    layer4_outputs(7618) <= (layer3_outputs(629)) and (layer3_outputs(5745));
    layer4_outputs(7619) <= not((layer3_outputs(792)) or (layer3_outputs(3014)));
    layer4_outputs(7620) <= not(layer3_outputs(4359));
    layer4_outputs(7621) <= not((layer3_outputs(3758)) and (layer3_outputs(7593)));
    layer4_outputs(7622) <= not(layer3_outputs(5895)) or (layer3_outputs(581));
    layer4_outputs(7623) <= (layer3_outputs(5981)) and not (layer3_outputs(3892));
    layer4_outputs(7624) <= not(layer3_outputs(5055)) or (layer3_outputs(6731));
    layer4_outputs(7625) <= (layer3_outputs(1351)) and not (layer3_outputs(286));
    layer4_outputs(7626) <= not(layer3_outputs(5351));
    layer4_outputs(7627) <= (layer3_outputs(2960)) and (layer3_outputs(2955));
    layer4_outputs(7628) <= not((layer3_outputs(160)) and (layer3_outputs(6934)));
    layer4_outputs(7629) <= not(layer3_outputs(3759)) or (layer3_outputs(5078));
    layer4_outputs(7630) <= not((layer3_outputs(2905)) xor (layer3_outputs(191)));
    layer4_outputs(7631) <= not((layer3_outputs(2096)) xor (layer3_outputs(3784)));
    layer4_outputs(7632) <= (layer3_outputs(6613)) xor (layer3_outputs(6684));
    layer4_outputs(7633) <= not((layer3_outputs(6988)) or (layer3_outputs(2936)));
    layer4_outputs(7634) <= (layer3_outputs(5428)) and not (layer3_outputs(6539));
    layer4_outputs(7635) <= not(layer3_outputs(2430));
    layer4_outputs(7636) <= not(layer3_outputs(3922));
    layer4_outputs(7637) <= not(layer3_outputs(6000));
    layer4_outputs(7638) <= (layer3_outputs(3624)) or (layer3_outputs(4311));
    layer4_outputs(7639) <= not((layer3_outputs(3324)) xor (layer3_outputs(7237)));
    layer4_outputs(7640) <= not((layer3_outputs(5667)) or (layer3_outputs(161)));
    layer4_outputs(7641) <= not((layer3_outputs(7092)) xor (layer3_outputs(6941)));
    layer4_outputs(7642) <= (layer3_outputs(6623)) and (layer3_outputs(5870));
    layer4_outputs(7643) <= layer3_outputs(3720);
    layer4_outputs(7644) <= not((layer3_outputs(5385)) and (layer3_outputs(380)));
    layer4_outputs(7645) <= layer3_outputs(4613);
    layer4_outputs(7646) <= layer3_outputs(393);
    layer4_outputs(7647) <= layer3_outputs(6671);
    layer4_outputs(7648) <= layer3_outputs(7637);
    layer4_outputs(7649) <= not(layer3_outputs(2558));
    layer4_outputs(7650) <= (layer3_outputs(176)) and (layer3_outputs(6027));
    layer4_outputs(7651) <= (layer3_outputs(150)) and not (layer3_outputs(2870));
    layer4_outputs(7652) <= (layer3_outputs(829)) and (layer3_outputs(1050));
    layer4_outputs(7653) <= not(layer3_outputs(4034));
    layer4_outputs(7654) <= (layer3_outputs(4993)) and not (layer3_outputs(4503));
    layer4_outputs(7655) <= (layer3_outputs(3521)) and not (layer3_outputs(5765));
    layer4_outputs(7656) <= not(layer3_outputs(6489));
    layer4_outputs(7657) <= not((layer3_outputs(3014)) and (layer3_outputs(5956)));
    layer4_outputs(7658) <= '1';
    layer4_outputs(7659) <= not((layer3_outputs(726)) xor (layer3_outputs(1093)));
    layer4_outputs(7660) <= not(layer3_outputs(7606)) or (layer3_outputs(2941));
    layer4_outputs(7661) <= (layer3_outputs(703)) and not (layer3_outputs(2697));
    layer4_outputs(7662) <= not((layer3_outputs(485)) xor (layer3_outputs(3019)));
    layer4_outputs(7663) <= layer3_outputs(1428);
    layer4_outputs(7664) <= (layer3_outputs(4445)) and not (layer3_outputs(3518));
    layer4_outputs(7665) <= not(layer3_outputs(4517)) or (layer3_outputs(5622));
    layer4_outputs(7666) <= not(layer3_outputs(3657));
    layer4_outputs(7667) <= not((layer3_outputs(7114)) and (layer3_outputs(2016)));
    layer4_outputs(7668) <= layer3_outputs(2983);
    layer4_outputs(7669) <= layer3_outputs(841);
    layer4_outputs(7670) <= not(layer3_outputs(3775));
    layer4_outputs(7671) <= not((layer3_outputs(1181)) or (layer3_outputs(807)));
    layer4_outputs(7672) <= (layer3_outputs(7267)) or (layer3_outputs(4263));
    layer4_outputs(7673) <= layer3_outputs(3472);
    layer4_outputs(7674) <= layer3_outputs(676);
    layer4_outputs(7675) <= not(layer3_outputs(5318));
    layer4_outputs(7676) <= layer3_outputs(3791);
    layer4_outputs(7677) <= (layer3_outputs(6320)) and not (layer3_outputs(6775));
    layer4_outputs(7678) <= not(layer3_outputs(2672)) or (layer3_outputs(412));
    layer4_outputs(7679) <= not(layer3_outputs(130));
    layer5_outputs(0) <= (layer4_outputs(6837)) and not (layer4_outputs(4098));
    layer5_outputs(1) <= not((layer4_outputs(2558)) xor (layer4_outputs(1537)));
    layer5_outputs(2) <= layer4_outputs(5535);
    layer5_outputs(3) <= not((layer4_outputs(4512)) xor (layer4_outputs(1705)));
    layer5_outputs(4) <= (layer4_outputs(5978)) xor (layer4_outputs(1342));
    layer5_outputs(5) <= not(layer4_outputs(7035));
    layer5_outputs(6) <= not(layer4_outputs(6152));
    layer5_outputs(7) <= not(layer4_outputs(712));
    layer5_outputs(8) <= (layer4_outputs(970)) and (layer4_outputs(4714));
    layer5_outputs(9) <= (layer4_outputs(5087)) and not (layer4_outputs(89));
    layer5_outputs(10) <= not(layer4_outputs(6771));
    layer5_outputs(11) <= not((layer4_outputs(5508)) xor (layer4_outputs(6428)));
    layer5_outputs(12) <= layer4_outputs(6727);
    layer5_outputs(13) <= not(layer4_outputs(6134));
    layer5_outputs(14) <= '0';
    layer5_outputs(15) <= layer4_outputs(6803);
    layer5_outputs(16) <= not((layer4_outputs(2405)) and (layer4_outputs(7496)));
    layer5_outputs(17) <= layer4_outputs(4482);
    layer5_outputs(18) <= layer4_outputs(509);
    layer5_outputs(19) <= not((layer4_outputs(4253)) xor (layer4_outputs(4009)));
    layer5_outputs(20) <= layer4_outputs(6825);
    layer5_outputs(21) <= layer4_outputs(7548);
    layer5_outputs(22) <= not((layer4_outputs(6545)) xor (layer4_outputs(3732)));
    layer5_outputs(23) <= not((layer4_outputs(3546)) or (layer4_outputs(5616)));
    layer5_outputs(24) <= not(layer4_outputs(6520));
    layer5_outputs(25) <= not(layer4_outputs(3483)) or (layer4_outputs(1768));
    layer5_outputs(26) <= not((layer4_outputs(7633)) and (layer4_outputs(7124)));
    layer5_outputs(27) <= layer4_outputs(5054);
    layer5_outputs(28) <= (layer4_outputs(4548)) and not (layer4_outputs(3743));
    layer5_outputs(29) <= not(layer4_outputs(511));
    layer5_outputs(30) <= not(layer4_outputs(4674)) or (layer4_outputs(6184));
    layer5_outputs(31) <= layer4_outputs(1796);
    layer5_outputs(32) <= (layer4_outputs(5379)) and (layer4_outputs(3951));
    layer5_outputs(33) <= layer4_outputs(1893);
    layer5_outputs(34) <= layer4_outputs(1607);
    layer5_outputs(35) <= not(layer4_outputs(3787));
    layer5_outputs(36) <= (layer4_outputs(331)) or (layer4_outputs(7200));
    layer5_outputs(37) <= not(layer4_outputs(685)) or (layer4_outputs(762));
    layer5_outputs(38) <= '0';
    layer5_outputs(39) <= '0';
    layer5_outputs(40) <= layer4_outputs(3636);
    layer5_outputs(41) <= not((layer4_outputs(2242)) xor (layer4_outputs(3438)));
    layer5_outputs(42) <= not(layer4_outputs(2188));
    layer5_outputs(43) <= (layer4_outputs(456)) xor (layer4_outputs(5194));
    layer5_outputs(44) <= not(layer4_outputs(198));
    layer5_outputs(45) <= (layer4_outputs(5701)) or (layer4_outputs(6869));
    layer5_outputs(46) <= not(layer4_outputs(6692));
    layer5_outputs(47) <= layer4_outputs(7394);
    layer5_outputs(48) <= (layer4_outputs(2397)) and not (layer4_outputs(2799));
    layer5_outputs(49) <= not(layer4_outputs(92));
    layer5_outputs(50) <= (layer4_outputs(3922)) and not (layer4_outputs(5421));
    layer5_outputs(51) <= not(layer4_outputs(4924));
    layer5_outputs(52) <= not(layer4_outputs(5192)) or (layer4_outputs(5083));
    layer5_outputs(53) <= not((layer4_outputs(2325)) xor (layer4_outputs(3589)));
    layer5_outputs(54) <= not(layer4_outputs(4222));
    layer5_outputs(55) <= not(layer4_outputs(2273));
    layer5_outputs(56) <= (layer4_outputs(6071)) or (layer4_outputs(6006));
    layer5_outputs(57) <= not((layer4_outputs(2141)) or (layer4_outputs(6036)));
    layer5_outputs(58) <= (layer4_outputs(6402)) and not (layer4_outputs(58));
    layer5_outputs(59) <= not(layer4_outputs(6600));
    layer5_outputs(60) <= (layer4_outputs(835)) or (layer4_outputs(6218));
    layer5_outputs(61) <= (layer4_outputs(820)) and (layer4_outputs(466));
    layer5_outputs(62) <= (layer4_outputs(2534)) or (layer4_outputs(710));
    layer5_outputs(63) <= (layer4_outputs(1254)) and not (layer4_outputs(4850));
    layer5_outputs(64) <= not(layer4_outputs(4491)) or (layer4_outputs(6727));
    layer5_outputs(65) <= layer4_outputs(6804);
    layer5_outputs(66) <= layer4_outputs(215);
    layer5_outputs(67) <= (layer4_outputs(1987)) xor (layer4_outputs(5110));
    layer5_outputs(68) <= (layer4_outputs(218)) and (layer4_outputs(3056));
    layer5_outputs(69) <= not(layer4_outputs(5750)) or (layer4_outputs(6248));
    layer5_outputs(70) <= not(layer4_outputs(6850));
    layer5_outputs(71) <= not(layer4_outputs(2110));
    layer5_outputs(72) <= (layer4_outputs(7079)) or (layer4_outputs(3589));
    layer5_outputs(73) <= (layer4_outputs(1640)) or (layer4_outputs(3212));
    layer5_outputs(74) <= not(layer4_outputs(1387)) or (layer4_outputs(6764));
    layer5_outputs(75) <= layer4_outputs(3955);
    layer5_outputs(76) <= layer4_outputs(6001);
    layer5_outputs(77) <= layer4_outputs(3943);
    layer5_outputs(78) <= not(layer4_outputs(4983));
    layer5_outputs(79) <= (layer4_outputs(7609)) and not (layer4_outputs(1556));
    layer5_outputs(80) <= layer4_outputs(4552);
    layer5_outputs(81) <= not(layer4_outputs(4327));
    layer5_outputs(82) <= layer4_outputs(786);
    layer5_outputs(83) <= layer4_outputs(3315);
    layer5_outputs(84) <= (layer4_outputs(2471)) and (layer4_outputs(983));
    layer5_outputs(85) <= not(layer4_outputs(2009)) or (layer4_outputs(6912));
    layer5_outputs(86) <= layer4_outputs(2480);
    layer5_outputs(87) <= layer4_outputs(1952);
    layer5_outputs(88) <= not(layer4_outputs(935)) or (layer4_outputs(5914));
    layer5_outputs(89) <= layer4_outputs(4266);
    layer5_outputs(90) <= (layer4_outputs(7227)) or (layer4_outputs(2715));
    layer5_outputs(91) <= not((layer4_outputs(2321)) or (layer4_outputs(4032)));
    layer5_outputs(92) <= not(layer4_outputs(4561));
    layer5_outputs(93) <= (layer4_outputs(5218)) and not (layer4_outputs(3692));
    layer5_outputs(94) <= (layer4_outputs(2431)) or (layer4_outputs(6564));
    layer5_outputs(95) <= (layer4_outputs(977)) and not (layer4_outputs(2569));
    layer5_outputs(96) <= not(layer4_outputs(3430));
    layer5_outputs(97) <= (layer4_outputs(2746)) and (layer4_outputs(911));
    layer5_outputs(98) <= not(layer4_outputs(2136)) or (layer4_outputs(2719));
    layer5_outputs(99) <= layer4_outputs(4521);
    layer5_outputs(100) <= (layer4_outputs(5257)) xor (layer4_outputs(601));
    layer5_outputs(101) <= layer4_outputs(2888);
    layer5_outputs(102) <= layer4_outputs(7014);
    layer5_outputs(103) <= not(layer4_outputs(5600));
    layer5_outputs(104) <= layer4_outputs(2567);
    layer5_outputs(105) <= not(layer4_outputs(1866));
    layer5_outputs(106) <= (layer4_outputs(2925)) and not (layer4_outputs(1444));
    layer5_outputs(107) <= layer4_outputs(6589);
    layer5_outputs(108) <= not(layer4_outputs(5328)) or (layer4_outputs(5574));
    layer5_outputs(109) <= not((layer4_outputs(1088)) xor (layer4_outputs(5581)));
    layer5_outputs(110) <= layer4_outputs(2260);
    layer5_outputs(111) <= layer4_outputs(1106);
    layer5_outputs(112) <= not((layer4_outputs(4560)) and (layer4_outputs(7568)));
    layer5_outputs(113) <= layer4_outputs(142);
    layer5_outputs(114) <= not(layer4_outputs(7191));
    layer5_outputs(115) <= not((layer4_outputs(4844)) and (layer4_outputs(3794)));
    layer5_outputs(116) <= (layer4_outputs(4292)) and not (layer4_outputs(6110));
    layer5_outputs(117) <= (layer4_outputs(7189)) xor (layer4_outputs(6853));
    layer5_outputs(118) <= (layer4_outputs(3275)) or (layer4_outputs(2357));
    layer5_outputs(119) <= not((layer4_outputs(5665)) xor (layer4_outputs(6)));
    layer5_outputs(120) <= not(layer4_outputs(5689));
    layer5_outputs(121) <= '1';
    layer5_outputs(122) <= (layer4_outputs(1331)) xor (layer4_outputs(7312));
    layer5_outputs(123) <= not(layer4_outputs(1531));
    layer5_outputs(124) <= layer4_outputs(4833);
    layer5_outputs(125) <= (layer4_outputs(4117)) xor (layer4_outputs(4428));
    layer5_outputs(126) <= not(layer4_outputs(3116));
    layer5_outputs(127) <= layer4_outputs(352);
    layer5_outputs(128) <= not(layer4_outputs(3285));
    layer5_outputs(129) <= not(layer4_outputs(973));
    layer5_outputs(130) <= layer4_outputs(378);
    layer5_outputs(131) <= not(layer4_outputs(6583));
    layer5_outputs(132) <= not(layer4_outputs(3070));
    layer5_outputs(133) <= (layer4_outputs(1323)) and not (layer4_outputs(984));
    layer5_outputs(134) <= layer4_outputs(2320);
    layer5_outputs(135) <= layer4_outputs(4934);
    layer5_outputs(136) <= not(layer4_outputs(5615));
    layer5_outputs(137) <= (layer4_outputs(4075)) and not (layer4_outputs(5482));
    layer5_outputs(138) <= layer4_outputs(1014);
    layer5_outputs(139) <= (layer4_outputs(7588)) and not (layer4_outputs(1274));
    layer5_outputs(140) <= not((layer4_outputs(641)) and (layer4_outputs(5778)));
    layer5_outputs(141) <= not(layer4_outputs(7241));
    layer5_outputs(142) <= not(layer4_outputs(5481));
    layer5_outputs(143) <= not(layer4_outputs(1329));
    layer5_outputs(144) <= (layer4_outputs(1350)) and not (layer4_outputs(1477));
    layer5_outputs(145) <= layer4_outputs(4847);
    layer5_outputs(146) <= not((layer4_outputs(6869)) or (layer4_outputs(2728)));
    layer5_outputs(147) <= not(layer4_outputs(5489));
    layer5_outputs(148) <= (layer4_outputs(4628)) and not (layer4_outputs(196));
    layer5_outputs(149) <= (layer4_outputs(2027)) and (layer4_outputs(3875));
    layer5_outputs(150) <= not(layer4_outputs(7236));
    layer5_outputs(151) <= (layer4_outputs(7024)) and not (layer4_outputs(416));
    layer5_outputs(152) <= not(layer4_outputs(3566)) or (layer4_outputs(3363));
    layer5_outputs(153) <= not(layer4_outputs(3069));
    layer5_outputs(154) <= not(layer4_outputs(6171));
    layer5_outputs(155) <= not((layer4_outputs(1175)) and (layer4_outputs(7575)));
    layer5_outputs(156) <= not((layer4_outputs(6011)) xor (layer4_outputs(83)));
    layer5_outputs(157) <= not((layer4_outputs(319)) xor (layer4_outputs(4118)));
    layer5_outputs(158) <= not(layer4_outputs(4233)) or (layer4_outputs(3818));
    layer5_outputs(159) <= layer4_outputs(1118);
    layer5_outputs(160) <= layer4_outputs(2043);
    layer5_outputs(161) <= not(layer4_outputs(4186));
    layer5_outputs(162) <= not(layer4_outputs(6230));
    layer5_outputs(163) <= (layer4_outputs(5619)) and (layer4_outputs(6263));
    layer5_outputs(164) <= not(layer4_outputs(6876));
    layer5_outputs(165) <= layer4_outputs(6417);
    layer5_outputs(166) <= not(layer4_outputs(4144));
    layer5_outputs(167) <= layer4_outputs(3758);
    layer5_outputs(168) <= not(layer4_outputs(3711));
    layer5_outputs(169) <= (layer4_outputs(903)) xor (layer4_outputs(2020));
    layer5_outputs(170) <= layer4_outputs(2683);
    layer5_outputs(171) <= layer4_outputs(3071);
    layer5_outputs(172) <= not((layer4_outputs(2637)) xor (layer4_outputs(1415)));
    layer5_outputs(173) <= not((layer4_outputs(5112)) and (layer4_outputs(5947)));
    layer5_outputs(174) <= (layer4_outputs(7617)) xor (layer4_outputs(2311));
    layer5_outputs(175) <= not(layer4_outputs(2515));
    layer5_outputs(176) <= not((layer4_outputs(1375)) xor (layer4_outputs(3553)));
    layer5_outputs(177) <= (layer4_outputs(1671)) and not (layer4_outputs(2240));
    layer5_outputs(178) <= not((layer4_outputs(1679)) and (layer4_outputs(4867)));
    layer5_outputs(179) <= layer4_outputs(5975);
    layer5_outputs(180) <= (layer4_outputs(7424)) or (layer4_outputs(5115));
    layer5_outputs(181) <= (layer4_outputs(7494)) and (layer4_outputs(4186));
    layer5_outputs(182) <= layer4_outputs(6581);
    layer5_outputs(183) <= not(layer4_outputs(5312));
    layer5_outputs(184) <= not(layer4_outputs(2002)) or (layer4_outputs(193));
    layer5_outputs(185) <= not(layer4_outputs(631));
    layer5_outputs(186) <= not((layer4_outputs(7067)) xor (layer4_outputs(4729)));
    layer5_outputs(187) <= layer4_outputs(3271);
    layer5_outputs(188) <= not(layer4_outputs(4243)) or (layer4_outputs(2419));
    layer5_outputs(189) <= (layer4_outputs(5273)) and (layer4_outputs(1179));
    layer5_outputs(190) <= not(layer4_outputs(2963));
    layer5_outputs(191) <= layer4_outputs(1133);
    layer5_outputs(192) <= (layer4_outputs(3814)) and not (layer4_outputs(6679));
    layer5_outputs(193) <= not((layer4_outputs(5186)) or (layer4_outputs(2270)));
    layer5_outputs(194) <= not(layer4_outputs(5018)) or (layer4_outputs(7121));
    layer5_outputs(195) <= layer4_outputs(4734);
    layer5_outputs(196) <= (layer4_outputs(6436)) xor (layer4_outputs(4083));
    layer5_outputs(197) <= not(layer4_outputs(6793)) or (layer4_outputs(427));
    layer5_outputs(198) <= not(layer4_outputs(1653)) or (layer4_outputs(332));
    layer5_outputs(199) <= layer4_outputs(3042);
    layer5_outputs(200) <= not(layer4_outputs(5068));
    layer5_outputs(201) <= not((layer4_outputs(5038)) xor (layer4_outputs(1463)));
    layer5_outputs(202) <= not((layer4_outputs(4456)) xor (layer4_outputs(5522)));
    layer5_outputs(203) <= (layer4_outputs(3475)) or (layer4_outputs(5673));
    layer5_outputs(204) <= not(layer4_outputs(3517));
    layer5_outputs(205) <= not(layer4_outputs(4615));
    layer5_outputs(206) <= layer4_outputs(6836);
    layer5_outputs(207) <= not(layer4_outputs(5375));
    layer5_outputs(208) <= not(layer4_outputs(318));
    layer5_outputs(209) <= layer4_outputs(7202);
    layer5_outputs(210) <= not(layer4_outputs(4743));
    layer5_outputs(211) <= not(layer4_outputs(3935)) or (layer4_outputs(5361));
    layer5_outputs(212) <= not(layer4_outputs(1108)) or (layer4_outputs(7044));
    layer5_outputs(213) <= (layer4_outputs(966)) and not (layer4_outputs(1234));
    layer5_outputs(214) <= (layer4_outputs(4447)) and (layer4_outputs(6954));
    layer5_outputs(215) <= (layer4_outputs(3486)) and (layer4_outputs(4817));
    layer5_outputs(216) <= not(layer4_outputs(6775));
    layer5_outputs(217) <= not(layer4_outputs(1559)) or (layer4_outputs(6382));
    layer5_outputs(218) <= not((layer4_outputs(4242)) and (layer4_outputs(6168)));
    layer5_outputs(219) <= '1';
    layer5_outputs(220) <= not((layer4_outputs(3013)) and (layer4_outputs(926)));
    layer5_outputs(221) <= layer4_outputs(5190);
    layer5_outputs(222) <= not(layer4_outputs(6347));
    layer5_outputs(223) <= not(layer4_outputs(7642));
    layer5_outputs(224) <= not((layer4_outputs(339)) or (layer4_outputs(5709)));
    layer5_outputs(225) <= layer4_outputs(4997);
    layer5_outputs(226) <= not(layer4_outputs(2418));
    layer5_outputs(227) <= not(layer4_outputs(5628));
    layer5_outputs(228) <= layer4_outputs(7119);
    layer5_outputs(229) <= layer4_outputs(809);
    layer5_outputs(230) <= layer4_outputs(4775);
    layer5_outputs(231) <= not((layer4_outputs(5633)) and (layer4_outputs(7176)));
    layer5_outputs(232) <= not(layer4_outputs(3386)) or (layer4_outputs(6896));
    layer5_outputs(233) <= not(layer4_outputs(2960)) or (layer4_outputs(586));
    layer5_outputs(234) <= not((layer4_outputs(947)) and (layer4_outputs(2129)));
    layer5_outputs(235) <= not(layer4_outputs(7111));
    layer5_outputs(236) <= not(layer4_outputs(66));
    layer5_outputs(237) <= not((layer4_outputs(3872)) xor (layer4_outputs(4444)));
    layer5_outputs(238) <= not((layer4_outputs(7245)) or (layer4_outputs(3656)));
    layer5_outputs(239) <= (layer4_outputs(5892)) and not (layer4_outputs(3837));
    layer5_outputs(240) <= layer4_outputs(6296);
    layer5_outputs(241) <= not(layer4_outputs(241)) or (layer4_outputs(2516));
    layer5_outputs(242) <= not((layer4_outputs(5162)) xor (layer4_outputs(1248)));
    layer5_outputs(243) <= not((layer4_outputs(5155)) xor (layer4_outputs(1401)));
    layer5_outputs(244) <= not(layer4_outputs(3978));
    layer5_outputs(245) <= not((layer4_outputs(4953)) and (layer4_outputs(90)));
    layer5_outputs(246) <= (layer4_outputs(1088)) and not (layer4_outputs(1745));
    layer5_outputs(247) <= not((layer4_outputs(941)) and (layer4_outputs(602)));
    layer5_outputs(248) <= layer4_outputs(3046);
    layer5_outputs(249) <= layer4_outputs(2078);
    layer5_outputs(250) <= not((layer4_outputs(6923)) and (layer4_outputs(620)));
    layer5_outputs(251) <= not(layer4_outputs(5449)) or (layer4_outputs(2177));
    layer5_outputs(252) <= (layer4_outputs(812)) and (layer4_outputs(6003));
    layer5_outputs(253) <= '1';
    layer5_outputs(254) <= not((layer4_outputs(6734)) xor (layer4_outputs(6097)));
    layer5_outputs(255) <= not(layer4_outputs(363));
    layer5_outputs(256) <= layer4_outputs(4576);
    layer5_outputs(257) <= not(layer4_outputs(4319)) or (layer4_outputs(1190));
    layer5_outputs(258) <= not(layer4_outputs(6906));
    layer5_outputs(259) <= layer4_outputs(7352);
    layer5_outputs(260) <= not((layer4_outputs(1587)) xor (layer4_outputs(1084)));
    layer5_outputs(261) <= (layer4_outputs(3204)) and not (layer4_outputs(2114));
    layer5_outputs(262) <= not(layer4_outputs(5414));
    layer5_outputs(263) <= layer4_outputs(251);
    layer5_outputs(264) <= layer4_outputs(5310);
    layer5_outputs(265) <= (layer4_outputs(6301)) xor (layer4_outputs(4712));
    layer5_outputs(266) <= not((layer4_outputs(1599)) xor (layer4_outputs(1462)));
    layer5_outputs(267) <= '0';
    layer5_outputs(268) <= not(layer4_outputs(6403));
    layer5_outputs(269) <= not(layer4_outputs(6158)) or (layer4_outputs(7040));
    layer5_outputs(270) <= not((layer4_outputs(7280)) xor (layer4_outputs(3448)));
    layer5_outputs(271) <= not(layer4_outputs(2633)) or (layer4_outputs(4309));
    layer5_outputs(272) <= layer4_outputs(281);
    layer5_outputs(273) <= layer4_outputs(1996);
    layer5_outputs(274) <= not((layer4_outputs(5064)) xor (layer4_outputs(2991)));
    layer5_outputs(275) <= not(layer4_outputs(4183));
    layer5_outputs(276) <= not(layer4_outputs(5057));
    layer5_outputs(277) <= not(layer4_outputs(7041));
    layer5_outputs(278) <= not(layer4_outputs(829));
    layer5_outputs(279) <= not(layer4_outputs(579));
    layer5_outputs(280) <= (layer4_outputs(2839)) or (layer4_outputs(2699));
    layer5_outputs(281) <= not(layer4_outputs(3105));
    layer5_outputs(282) <= layer4_outputs(5371);
    layer5_outputs(283) <= layer4_outputs(5425);
    layer5_outputs(284) <= not(layer4_outputs(7627)) or (layer4_outputs(7205));
    layer5_outputs(285) <= layer4_outputs(197);
    layer5_outputs(286) <= not(layer4_outputs(6066));
    layer5_outputs(287) <= layer4_outputs(2056);
    layer5_outputs(288) <= not((layer4_outputs(6026)) xor (layer4_outputs(5094)));
    layer5_outputs(289) <= layer4_outputs(3940);
    layer5_outputs(290) <= not(layer4_outputs(3130));
    layer5_outputs(291) <= not(layer4_outputs(2475));
    layer5_outputs(292) <= (layer4_outputs(5632)) xor (layer4_outputs(5831));
    layer5_outputs(293) <= layer4_outputs(5409);
    layer5_outputs(294) <= not((layer4_outputs(3756)) or (layer4_outputs(4141)));
    layer5_outputs(295) <= (layer4_outputs(5814)) and not (layer4_outputs(7478));
    layer5_outputs(296) <= not(layer4_outputs(3346)) or (layer4_outputs(1244));
    layer5_outputs(297) <= not(layer4_outputs(3967));
    layer5_outputs(298) <= layer4_outputs(3671);
    layer5_outputs(299) <= not((layer4_outputs(5711)) or (layer4_outputs(3574)));
    layer5_outputs(300) <= not(layer4_outputs(3821));
    layer5_outputs(301) <= layer4_outputs(2478);
    layer5_outputs(302) <= layer4_outputs(1337);
    layer5_outputs(303) <= layer4_outputs(327);
    layer5_outputs(304) <= not(layer4_outputs(3362));
    layer5_outputs(305) <= layer4_outputs(5524);
    layer5_outputs(306) <= (layer4_outputs(1145)) and not (layer4_outputs(3330));
    layer5_outputs(307) <= not(layer4_outputs(5705)) or (layer4_outputs(7023));
    layer5_outputs(308) <= (layer4_outputs(7173)) xor (layer4_outputs(4081));
    layer5_outputs(309) <= not(layer4_outputs(308));
    layer5_outputs(310) <= layer4_outputs(7291);
    layer5_outputs(311) <= layer4_outputs(5469);
    layer5_outputs(312) <= layer4_outputs(5402);
    layer5_outputs(313) <= not((layer4_outputs(3079)) or (layer4_outputs(6777)));
    layer5_outputs(314) <= layer4_outputs(6356);
    layer5_outputs(315) <= layer4_outputs(6345);
    layer5_outputs(316) <= layer4_outputs(4113);
    layer5_outputs(317) <= (layer4_outputs(1374)) and not (layer4_outputs(1072));
    layer5_outputs(318) <= not(layer4_outputs(2073));
    layer5_outputs(319) <= not((layer4_outputs(6735)) xor (layer4_outputs(1036)));
    layer5_outputs(320) <= layer4_outputs(1174);
    layer5_outputs(321) <= (layer4_outputs(3280)) or (layer4_outputs(5172));
    layer5_outputs(322) <= layer4_outputs(4880);
    layer5_outputs(323) <= not((layer4_outputs(2649)) or (layer4_outputs(7107)));
    layer5_outputs(324) <= layer4_outputs(190);
    layer5_outputs(325) <= not(layer4_outputs(7396));
    layer5_outputs(326) <= not((layer4_outputs(1591)) or (layer4_outputs(3252)));
    layer5_outputs(327) <= not(layer4_outputs(1107));
    layer5_outputs(328) <= not(layer4_outputs(227));
    layer5_outputs(329) <= not((layer4_outputs(1450)) xor (layer4_outputs(1971)));
    layer5_outputs(330) <= not(layer4_outputs(5819));
    layer5_outputs(331) <= not(layer4_outputs(6115)) or (layer4_outputs(2758));
    layer5_outputs(332) <= not((layer4_outputs(7539)) xor (layer4_outputs(2154)));
    layer5_outputs(333) <= not(layer4_outputs(1896));
    layer5_outputs(334) <= not((layer4_outputs(1028)) xor (layer4_outputs(4806)));
    layer5_outputs(335) <= not((layer4_outputs(3300)) xor (layer4_outputs(6611)));
    layer5_outputs(336) <= (layer4_outputs(6861)) or (layer4_outputs(5092));
    layer5_outputs(337) <= (layer4_outputs(4250)) or (layer4_outputs(3947));
    layer5_outputs(338) <= not((layer4_outputs(273)) or (layer4_outputs(5410)));
    layer5_outputs(339) <= not(layer4_outputs(393));
    layer5_outputs(340) <= layer4_outputs(6107);
    layer5_outputs(341) <= not(layer4_outputs(1516)) or (layer4_outputs(1474));
    layer5_outputs(342) <= layer4_outputs(5209);
    layer5_outputs(343) <= not(layer4_outputs(3547));
    layer5_outputs(344) <= (layer4_outputs(4142)) and not (layer4_outputs(1828));
    layer5_outputs(345) <= (layer4_outputs(157)) and not (layer4_outputs(2493));
    layer5_outputs(346) <= not(layer4_outputs(6725));
    layer5_outputs(347) <= not(layer4_outputs(3372));
    layer5_outputs(348) <= (layer4_outputs(6478)) or (layer4_outputs(2062));
    layer5_outputs(349) <= layer4_outputs(663);
    layer5_outputs(350) <= not(layer4_outputs(4848));
    layer5_outputs(351) <= '0';
    layer5_outputs(352) <= (layer4_outputs(5550)) and not (layer4_outputs(865));
    layer5_outputs(353) <= (layer4_outputs(2769)) or (layer4_outputs(290));
    layer5_outputs(354) <= not((layer4_outputs(1682)) and (layer4_outputs(18)));
    layer5_outputs(355) <= not(layer4_outputs(5833));
    layer5_outputs(356) <= not(layer4_outputs(2691));
    layer5_outputs(357) <= layer4_outputs(4918);
    layer5_outputs(358) <= (layer4_outputs(339)) and (layer4_outputs(3288));
    layer5_outputs(359) <= layer4_outputs(6720);
    layer5_outputs(360) <= not(layer4_outputs(3996)) or (layer4_outputs(3234));
    layer5_outputs(361) <= not(layer4_outputs(4058));
    layer5_outputs(362) <= not(layer4_outputs(1776));
    layer5_outputs(363) <= not((layer4_outputs(3715)) and (layer4_outputs(1268)));
    layer5_outputs(364) <= not((layer4_outputs(4542)) and (layer4_outputs(640)));
    layer5_outputs(365) <= layer4_outputs(7479);
    layer5_outputs(366) <= layer4_outputs(650);
    layer5_outputs(367) <= not(layer4_outputs(5014)) or (layer4_outputs(2203));
    layer5_outputs(368) <= not((layer4_outputs(4348)) or (layer4_outputs(1919)));
    layer5_outputs(369) <= not((layer4_outputs(6141)) and (layer4_outputs(7016)));
    layer5_outputs(370) <= layer4_outputs(6105);
    layer5_outputs(371) <= not((layer4_outputs(1353)) xor (layer4_outputs(3250)));
    layer5_outputs(372) <= (layer4_outputs(4646)) and not (layer4_outputs(4068));
    layer5_outputs(373) <= not((layer4_outputs(2115)) or (layer4_outputs(7308)));
    layer5_outputs(374) <= (layer4_outputs(6349)) and not (layer4_outputs(4915));
    layer5_outputs(375) <= layer4_outputs(2282);
    layer5_outputs(376) <= not((layer4_outputs(3935)) xor (layer4_outputs(1950)));
    layer5_outputs(377) <= layer4_outputs(1211);
    layer5_outputs(378) <= layer4_outputs(2223);
    layer5_outputs(379) <= layer4_outputs(4655);
    layer5_outputs(380) <= not((layer4_outputs(1246)) xor (layer4_outputs(5028)));
    layer5_outputs(381) <= not(layer4_outputs(4619)) or (layer4_outputs(2968));
    layer5_outputs(382) <= layer4_outputs(3340);
    layer5_outputs(383) <= not((layer4_outputs(4486)) and (layer4_outputs(889)));
    layer5_outputs(384) <= not((layer4_outputs(113)) xor (layer4_outputs(5354)));
    layer5_outputs(385) <= (layer4_outputs(5039)) or (layer4_outputs(3583));
    layer5_outputs(386) <= not((layer4_outputs(7679)) and (layer4_outputs(7156)));
    layer5_outputs(387) <= layer4_outputs(1045);
    layer5_outputs(388) <= layer4_outputs(6721);
    layer5_outputs(389) <= not(layer4_outputs(1763));
    layer5_outputs(390) <= (layer4_outputs(4539)) and (layer4_outputs(2816));
    layer5_outputs(391) <= not(layer4_outputs(7199));
    layer5_outputs(392) <= layer4_outputs(1243);
    layer5_outputs(393) <= (layer4_outputs(5291)) and not (layer4_outputs(1968));
    layer5_outputs(394) <= layer4_outputs(1882);
    layer5_outputs(395) <= not(layer4_outputs(155));
    layer5_outputs(396) <= layer4_outputs(3649);
    layer5_outputs(397) <= not((layer4_outputs(6685)) and (layer4_outputs(1975)));
    layer5_outputs(398) <= layer4_outputs(5813);
    layer5_outputs(399) <= (layer4_outputs(2956)) and not (layer4_outputs(6145));
    layer5_outputs(400) <= layer4_outputs(2124);
    layer5_outputs(401) <= not(layer4_outputs(1161));
    layer5_outputs(402) <= not(layer4_outputs(329));
    layer5_outputs(403) <= not((layer4_outputs(5927)) and (layer4_outputs(1230)));
    layer5_outputs(404) <= not(layer4_outputs(4621));
    layer5_outputs(405) <= layer4_outputs(3681);
    layer5_outputs(406) <= not((layer4_outputs(2517)) or (layer4_outputs(2947)));
    layer5_outputs(407) <= layer4_outputs(2407);
    layer5_outputs(408) <= (layer4_outputs(5887)) and (layer4_outputs(7531));
    layer5_outputs(409) <= not(layer4_outputs(4110));
    layer5_outputs(410) <= '1';
    layer5_outputs(411) <= not(layer4_outputs(7286));
    layer5_outputs(412) <= not(layer4_outputs(4501));
    layer5_outputs(413) <= not((layer4_outputs(3677)) and (layer4_outputs(873)));
    layer5_outputs(414) <= layer4_outputs(3566);
    layer5_outputs(415) <= not(layer4_outputs(1991)) or (layer4_outputs(6293));
    layer5_outputs(416) <= not((layer4_outputs(3121)) or (layer4_outputs(200)));
    layer5_outputs(417) <= not((layer4_outputs(5698)) and (layer4_outputs(5292)));
    layer5_outputs(418) <= (layer4_outputs(2635)) and not (layer4_outputs(6509));
    layer5_outputs(419) <= not((layer4_outputs(2057)) or (layer4_outputs(825)));
    layer5_outputs(420) <= not(layer4_outputs(373));
    layer5_outputs(421) <= layer4_outputs(1437);
    layer5_outputs(422) <= (layer4_outputs(6515)) and not (layer4_outputs(7106));
    layer5_outputs(423) <= not(layer4_outputs(2846));
    layer5_outputs(424) <= not(layer4_outputs(3454)) or (layer4_outputs(6533));
    layer5_outputs(425) <= layer4_outputs(2106);
    layer5_outputs(426) <= not(layer4_outputs(872));
    layer5_outputs(427) <= not(layer4_outputs(6336)) or (layer4_outputs(450));
    layer5_outputs(428) <= not((layer4_outputs(5821)) xor (layer4_outputs(1810)));
    layer5_outputs(429) <= not(layer4_outputs(5360));
    layer5_outputs(430) <= layer4_outputs(3700);
    layer5_outputs(431) <= layer4_outputs(5519);
    layer5_outputs(432) <= not(layer4_outputs(4904));
    layer5_outputs(433) <= layer4_outputs(2134);
    layer5_outputs(434) <= layer4_outputs(576);
    layer5_outputs(435) <= layer4_outputs(1892);
    layer5_outputs(436) <= not((layer4_outputs(2744)) xor (layer4_outputs(7611)));
    layer5_outputs(437) <= not((layer4_outputs(4151)) or (layer4_outputs(3485)));
    layer5_outputs(438) <= (layer4_outputs(3302)) xor (layer4_outputs(412));
    layer5_outputs(439) <= not(layer4_outputs(423));
    layer5_outputs(440) <= layer4_outputs(3939);
    layer5_outputs(441) <= not(layer4_outputs(188));
    layer5_outputs(442) <= layer4_outputs(563);
    layer5_outputs(443) <= (layer4_outputs(5080)) and not (layer4_outputs(4102));
    layer5_outputs(444) <= (layer4_outputs(4742)) and not (layer4_outputs(554));
    layer5_outputs(445) <= not((layer4_outputs(2999)) xor (layer4_outputs(4280)));
    layer5_outputs(446) <= (layer4_outputs(7266)) and not (layer4_outputs(5016));
    layer5_outputs(447) <= layer4_outputs(6075);
    layer5_outputs(448) <= not((layer4_outputs(5698)) xor (layer4_outputs(6699)));
    layer5_outputs(449) <= not(layer4_outputs(3202));
    layer5_outputs(450) <= not(layer4_outputs(1464));
    layer5_outputs(451) <= layer4_outputs(4585);
    layer5_outputs(452) <= (layer4_outputs(3626)) and not (layer4_outputs(1026));
    layer5_outputs(453) <= not(layer4_outputs(4849)) or (layer4_outputs(3209));
    layer5_outputs(454) <= not(layer4_outputs(1210));
    layer5_outputs(455) <= not((layer4_outputs(3567)) or (layer4_outputs(1624)));
    layer5_outputs(456) <= not(layer4_outputs(7384));
    layer5_outputs(457) <= not(layer4_outputs(686)) or (layer4_outputs(7264));
    layer5_outputs(458) <= layer4_outputs(1060);
    layer5_outputs(459) <= layer4_outputs(516);
    layer5_outputs(460) <= '1';
    layer5_outputs(461) <= not(layer4_outputs(672));
    layer5_outputs(462) <= layer4_outputs(2353);
    layer5_outputs(463) <= not(layer4_outputs(3815)) or (layer4_outputs(6349));
    layer5_outputs(464) <= (layer4_outputs(5065)) and not (layer4_outputs(6446));
    layer5_outputs(465) <= (layer4_outputs(2257)) xor (layer4_outputs(1988));
    layer5_outputs(466) <= layer4_outputs(2698);
    layer5_outputs(467) <= (layer4_outputs(6096)) or (layer4_outputs(5949));
    layer5_outputs(468) <= (layer4_outputs(6543)) and not (layer4_outputs(2499));
    layer5_outputs(469) <= '0';
    layer5_outputs(470) <= (layer4_outputs(6602)) or (layer4_outputs(3826));
    layer5_outputs(471) <= (layer4_outputs(3149)) and not (layer4_outputs(6957));
    layer5_outputs(472) <= not(layer4_outputs(6127)) or (layer4_outputs(7653));
    layer5_outputs(473) <= layer4_outputs(4877);
    layer5_outputs(474) <= (layer4_outputs(7478)) or (layer4_outputs(7282));
    layer5_outputs(475) <= not(layer4_outputs(7345));
    layer5_outputs(476) <= layer4_outputs(3477);
    layer5_outputs(477) <= not((layer4_outputs(2809)) and (layer4_outputs(5188)));
    layer5_outputs(478) <= not((layer4_outputs(946)) xor (layer4_outputs(5732)));
    layer5_outputs(479) <= not(layer4_outputs(2913)) or (layer4_outputs(6187));
    layer5_outputs(480) <= layer4_outputs(4688);
    layer5_outputs(481) <= layer4_outputs(5975);
    layer5_outputs(482) <= (layer4_outputs(5060)) and (layer4_outputs(3155));
    layer5_outputs(483) <= not(layer4_outputs(3614)) or (layer4_outputs(7068));
    layer5_outputs(484) <= layer4_outputs(1009);
    layer5_outputs(485) <= not(layer4_outputs(4289));
    layer5_outputs(486) <= not(layer4_outputs(2660));
    layer5_outputs(487) <= (layer4_outputs(4679)) and not (layer4_outputs(3268));
    layer5_outputs(488) <= layer4_outputs(2931);
    layer5_outputs(489) <= not((layer4_outputs(6468)) xor (layer4_outputs(4090)));
    layer5_outputs(490) <= not(layer4_outputs(1898)) or (layer4_outputs(6786));
    layer5_outputs(491) <= (layer4_outputs(2265)) xor (layer4_outputs(2040));
    layer5_outputs(492) <= layer4_outputs(3304);
    layer5_outputs(493) <= not(layer4_outputs(3222)) or (layer4_outputs(1728));
    layer5_outputs(494) <= not(layer4_outputs(7339)) or (layer4_outputs(5192));
    layer5_outputs(495) <= layer4_outputs(6616);
    layer5_outputs(496) <= not((layer4_outputs(2871)) and (layer4_outputs(4261)));
    layer5_outputs(497) <= not(layer4_outputs(7165)) or (layer4_outputs(5612));
    layer5_outputs(498) <= (layer4_outputs(1453)) and (layer4_outputs(6544));
    layer5_outputs(499) <= (layer4_outputs(5011)) and not (layer4_outputs(6292));
    layer5_outputs(500) <= layer4_outputs(1767);
    layer5_outputs(501) <= not(layer4_outputs(3046));
    layer5_outputs(502) <= not(layer4_outputs(5202)) or (layer4_outputs(3637));
    layer5_outputs(503) <= '0';
    layer5_outputs(504) <= not((layer4_outputs(1414)) or (layer4_outputs(5474)));
    layer5_outputs(505) <= not(layer4_outputs(3468));
    layer5_outputs(506) <= layer4_outputs(6080);
    layer5_outputs(507) <= (layer4_outputs(6458)) xor (layer4_outputs(5931));
    layer5_outputs(508) <= (layer4_outputs(4097)) and not (layer4_outputs(1475));
    layer5_outputs(509) <= not((layer4_outputs(14)) and (layer4_outputs(3171)));
    layer5_outputs(510) <= not(layer4_outputs(4768));
    layer5_outputs(511) <= (layer4_outputs(7386)) xor (layer4_outputs(1061));
    layer5_outputs(512) <= (layer4_outputs(2296)) xor (layer4_outputs(6228));
    layer5_outputs(513) <= not(layer4_outputs(575));
    layer5_outputs(514) <= (layer4_outputs(6390)) and (layer4_outputs(1447));
    layer5_outputs(515) <= not((layer4_outputs(874)) and (layer4_outputs(741)));
    layer5_outputs(516) <= not((layer4_outputs(7371)) or (layer4_outputs(1099)));
    layer5_outputs(517) <= not(layer4_outputs(748));
    layer5_outputs(518) <= '0';
    layer5_outputs(519) <= not(layer4_outputs(4229));
    layer5_outputs(520) <= not(layer4_outputs(6882));
    layer5_outputs(521) <= (layer4_outputs(1323)) and (layer4_outputs(7245));
    layer5_outputs(522) <= not(layer4_outputs(5581)) or (layer4_outputs(139));
    layer5_outputs(523) <= (layer4_outputs(1653)) and not (layer4_outputs(188));
    layer5_outputs(524) <= (layer4_outputs(3670)) and not (layer4_outputs(2221));
    layer5_outputs(525) <= layer4_outputs(6431);
    layer5_outputs(526) <= not(layer4_outputs(2958));
    layer5_outputs(527) <= not((layer4_outputs(2076)) and (layer4_outputs(2438)));
    layer5_outputs(528) <= not((layer4_outputs(6447)) or (layer4_outputs(167)));
    layer5_outputs(529) <= layer4_outputs(403);
    layer5_outputs(530) <= (layer4_outputs(1793)) and not (layer4_outputs(2266));
    layer5_outputs(531) <= not(layer4_outputs(3318));
    layer5_outputs(532) <= layer4_outputs(7596);
    layer5_outputs(533) <= not(layer4_outputs(3476)) or (layer4_outputs(7391));
    layer5_outputs(534) <= not(layer4_outputs(2560));
    layer5_outputs(535) <= (layer4_outputs(831)) and not (layer4_outputs(918));
    layer5_outputs(536) <= (layer4_outputs(7120)) and (layer4_outputs(6738));
    layer5_outputs(537) <= layer4_outputs(4450);
    layer5_outputs(538) <= layer4_outputs(7390);
    layer5_outputs(539) <= not(layer4_outputs(1538));
    layer5_outputs(540) <= layer4_outputs(2550);
    layer5_outputs(541) <= layer4_outputs(5893);
    layer5_outputs(542) <= not(layer4_outputs(4987)) or (layer4_outputs(702));
    layer5_outputs(543) <= not((layer4_outputs(2285)) xor (layer4_outputs(2206)));
    layer5_outputs(544) <= layer4_outputs(7172);
    layer5_outputs(545) <= layer4_outputs(5393);
    layer5_outputs(546) <= (layer4_outputs(2202)) xor (layer4_outputs(5987));
    layer5_outputs(547) <= not(layer4_outputs(3242));
    layer5_outputs(548) <= (layer4_outputs(5528)) and not (layer4_outputs(2276));
    layer5_outputs(549) <= (layer4_outputs(3606)) and not (layer4_outputs(1079));
    layer5_outputs(550) <= layer4_outputs(6202);
    layer5_outputs(551) <= (layer4_outputs(3611)) and not (layer4_outputs(2441));
    layer5_outputs(552) <= not((layer4_outputs(1288)) or (layer4_outputs(354)));
    layer5_outputs(553) <= (layer4_outputs(671)) and not (layer4_outputs(2438));
    layer5_outputs(554) <= not((layer4_outputs(3880)) xor (layer4_outputs(5927)));
    layer5_outputs(555) <= (layer4_outputs(4369)) and not (layer4_outputs(642));
    layer5_outputs(556) <= (layer4_outputs(2209)) and not (layer4_outputs(6616));
    layer5_outputs(557) <= not((layer4_outputs(1272)) xor (layer4_outputs(3570)));
    layer5_outputs(558) <= layer4_outputs(5899);
    layer5_outputs(559) <= not(layer4_outputs(5956));
    layer5_outputs(560) <= (layer4_outputs(216)) and not (layer4_outputs(6111));
    layer5_outputs(561) <= not(layer4_outputs(3256));
    layer5_outputs(562) <= layer4_outputs(769);
    layer5_outputs(563) <= (layer4_outputs(1168)) and (layer4_outputs(1596));
    layer5_outputs(564) <= layer4_outputs(5480);
    layer5_outputs(565) <= layer4_outputs(3008);
    layer5_outputs(566) <= not(layer4_outputs(2724));
    layer5_outputs(567) <= not(layer4_outputs(3441));
    layer5_outputs(568) <= (layer4_outputs(3863)) and not (layer4_outputs(2134));
    layer5_outputs(569) <= layer4_outputs(768);
    layer5_outputs(570) <= layer4_outputs(4562);
    layer5_outputs(571) <= layer4_outputs(343);
    layer5_outputs(572) <= not(layer4_outputs(6365)) or (layer4_outputs(1821));
    layer5_outputs(573) <= not(layer4_outputs(3271)) or (layer4_outputs(5836));
    layer5_outputs(574) <= (layer4_outputs(279)) and (layer4_outputs(3325));
    layer5_outputs(575) <= layer4_outputs(2751);
    layer5_outputs(576) <= not(layer4_outputs(6999));
    layer5_outputs(577) <= (layer4_outputs(2574)) xor (layer4_outputs(3382));
    layer5_outputs(578) <= not(layer4_outputs(2549));
    layer5_outputs(579) <= not((layer4_outputs(813)) and (layer4_outputs(2083)));
    layer5_outputs(580) <= (layer4_outputs(515)) xor (layer4_outputs(5606));
    layer5_outputs(581) <= (layer4_outputs(5134)) and not (layer4_outputs(5759));
    layer5_outputs(582) <= not(layer4_outputs(3973));
    layer5_outputs(583) <= not(layer4_outputs(3039));
    layer5_outputs(584) <= not(layer4_outputs(4553));
    layer5_outputs(585) <= not(layer4_outputs(2354));
    layer5_outputs(586) <= not((layer4_outputs(5601)) xor (layer4_outputs(6485)));
    layer5_outputs(587) <= layer4_outputs(2341);
    layer5_outputs(588) <= (layer4_outputs(1069)) xor (layer4_outputs(5299));
    layer5_outputs(589) <= not(layer4_outputs(2091));
    layer5_outputs(590) <= (layer4_outputs(4130)) and (layer4_outputs(6270));
    layer5_outputs(591) <= not((layer4_outputs(6810)) and (layer4_outputs(5857)));
    layer5_outputs(592) <= not((layer4_outputs(6021)) xor (layer4_outputs(1678)));
    layer5_outputs(593) <= layer4_outputs(3528);
    layer5_outputs(594) <= layer4_outputs(4449);
    layer5_outputs(595) <= not(layer4_outputs(5420));
    layer5_outputs(596) <= (layer4_outputs(2785)) and not (layer4_outputs(6233));
    layer5_outputs(597) <= layer4_outputs(3463);
    layer5_outputs(598) <= (layer4_outputs(3991)) xor (layer4_outputs(1251));
    layer5_outputs(599) <= (layer4_outputs(2975)) and not (layer4_outputs(6573));
    layer5_outputs(600) <= not(layer4_outputs(4535));
    layer5_outputs(601) <= '1';
    layer5_outputs(602) <= layer4_outputs(1523);
    layer5_outputs(603) <= (layer4_outputs(5244)) and not (layer4_outputs(3685));
    layer5_outputs(604) <= (layer4_outputs(285)) and (layer4_outputs(484));
    layer5_outputs(605) <= not(layer4_outputs(7100));
    layer5_outputs(606) <= not(layer4_outputs(7437));
    layer5_outputs(607) <= not((layer4_outputs(157)) xor (layer4_outputs(6269)));
    layer5_outputs(608) <= not(layer4_outputs(5210));
    layer5_outputs(609) <= (layer4_outputs(6762)) or (layer4_outputs(7574));
    layer5_outputs(610) <= not(layer4_outputs(1563));
    layer5_outputs(611) <= not((layer4_outputs(3811)) or (layer4_outputs(6967)));
    layer5_outputs(612) <= (layer4_outputs(6434)) and not (layer4_outputs(1419));
    layer5_outputs(613) <= not((layer4_outputs(6276)) xor (layer4_outputs(7034)));
    layer5_outputs(614) <= layer4_outputs(5260);
    layer5_outputs(615) <= (layer4_outputs(6750)) xor (layer4_outputs(6170));
    layer5_outputs(616) <= (layer4_outputs(5151)) and not (layer4_outputs(3538));
    layer5_outputs(617) <= layer4_outputs(2330);
    layer5_outputs(618) <= (layer4_outputs(6801)) and not (layer4_outputs(2068));
    layer5_outputs(619) <= layer4_outputs(5313);
    layer5_outputs(620) <= layer4_outputs(459);
    layer5_outputs(621) <= not(layer4_outputs(4230));
    layer5_outputs(622) <= (layer4_outputs(3424)) and (layer4_outputs(1362));
    layer5_outputs(623) <= layer4_outputs(5461);
    layer5_outputs(624) <= (layer4_outputs(3684)) or (layer4_outputs(346));
    layer5_outputs(625) <= not(layer4_outputs(6549)) or (layer4_outputs(367));
    layer5_outputs(626) <= layer4_outputs(1659);
    layer5_outputs(627) <= not(layer4_outputs(327));
    layer5_outputs(628) <= (layer4_outputs(4063)) or (layer4_outputs(6188));
    layer5_outputs(629) <= layer4_outputs(2463);
    layer5_outputs(630) <= layer4_outputs(1703);
    layer5_outputs(631) <= layer4_outputs(3035);
    layer5_outputs(632) <= not(layer4_outputs(5079)) or (layer4_outputs(839));
    layer5_outputs(633) <= layer4_outputs(7171);
    layer5_outputs(634) <= not(layer4_outputs(2767));
    layer5_outputs(635) <= not(layer4_outputs(2708));
    layer5_outputs(636) <= not(layer4_outputs(4123));
    layer5_outputs(637) <= not(layer4_outputs(4758)) or (layer4_outputs(3143));
    layer5_outputs(638) <= (layer4_outputs(4320)) and not (layer4_outputs(572));
    layer5_outputs(639) <= layer4_outputs(946);
    layer5_outputs(640) <= not((layer4_outputs(1136)) xor (layer4_outputs(4501)));
    layer5_outputs(641) <= (layer4_outputs(3957)) or (layer4_outputs(3506));
    layer5_outputs(642) <= layer4_outputs(2680);
    layer5_outputs(643) <= not(layer4_outputs(7037));
    layer5_outputs(644) <= (layer4_outputs(5605)) and not (layer4_outputs(1904));
    layer5_outputs(645) <= (layer4_outputs(3050)) and not (layer4_outputs(4571));
    layer5_outputs(646) <= not(layer4_outputs(6612));
    layer5_outputs(647) <= not((layer4_outputs(3718)) or (layer4_outputs(4625)));
    layer5_outputs(648) <= (layer4_outputs(2562)) or (layer4_outputs(6355));
    layer5_outputs(649) <= layer4_outputs(6767);
    layer5_outputs(650) <= not((layer4_outputs(4412)) and (layer4_outputs(5531)));
    layer5_outputs(651) <= (layer4_outputs(7321)) or (layer4_outputs(1496));
    layer5_outputs(652) <= not(layer4_outputs(1455));
    layer5_outputs(653) <= not(layer4_outputs(5069));
    layer5_outputs(654) <= (layer4_outputs(2576)) and not (layer4_outputs(1016));
    layer5_outputs(655) <= not(layer4_outputs(1722)) or (layer4_outputs(6951));
    layer5_outputs(656) <= (layer4_outputs(6214)) and not (layer4_outputs(3556));
    layer5_outputs(657) <= layer4_outputs(29);
    layer5_outputs(658) <= not((layer4_outputs(4240)) xor (layer4_outputs(2187)));
    layer5_outputs(659) <= layer4_outputs(4005);
    layer5_outputs(660) <= layer4_outputs(6232);
    layer5_outputs(661) <= layer4_outputs(6785);
    layer5_outputs(662) <= (layer4_outputs(5045)) and not (layer4_outputs(4360));
    layer5_outputs(663) <= not(layer4_outputs(179)) or (layer4_outputs(7061));
    layer5_outputs(664) <= layer4_outputs(1604);
    layer5_outputs(665) <= layer4_outputs(2263);
    layer5_outputs(666) <= not(layer4_outputs(699));
    layer5_outputs(667) <= layer4_outputs(7249);
    layer5_outputs(668) <= not((layer4_outputs(130)) xor (layer4_outputs(3629)));
    layer5_outputs(669) <= not(layer4_outputs(823)) or (layer4_outputs(1206));
    layer5_outputs(670) <= not(layer4_outputs(2056));
    layer5_outputs(671) <= (layer4_outputs(3034)) and not (layer4_outputs(3800));
    layer5_outputs(672) <= not(layer4_outputs(5699));
    layer5_outputs(673) <= layer4_outputs(236);
    layer5_outputs(674) <= (layer4_outputs(568)) and not (layer4_outputs(3269));
    layer5_outputs(675) <= layer4_outputs(2476);
    layer5_outputs(676) <= (layer4_outputs(7559)) xor (layer4_outputs(4311));
    layer5_outputs(677) <= '0';
    layer5_outputs(678) <= (layer4_outputs(648)) and not (layer4_outputs(4704));
    layer5_outputs(679) <= (layer4_outputs(1967)) and not (layer4_outputs(7471));
    layer5_outputs(680) <= '0';
    layer5_outputs(681) <= not(layer4_outputs(2124)) or (layer4_outputs(6868));
    layer5_outputs(682) <= (layer4_outputs(1061)) and not (layer4_outputs(4606));
    layer5_outputs(683) <= not(layer4_outputs(4061));
    layer5_outputs(684) <= layer4_outputs(2826);
    layer5_outputs(685) <= (layer4_outputs(7670)) and not (layer4_outputs(3516));
    layer5_outputs(686) <= layer4_outputs(4515);
    layer5_outputs(687) <= not(layer4_outputs(1884));
    layer5_outputs(688) <= (layer4_outputs(2001)) and not (layer4_outputs(7141));
    layer5_outputs(689) <= not(layer4_outputs(4943));
    layer5_outputs(690) <= '1';
    layer5_outputs(691) <= not(layer4_outputs(3585));
    layer5_outputs(692) <= not(layer4_outputs(1159));
    layer5_outputs(693) <= layer4_outputs(6991);
    layer5_outputs(694) <= not(layer4_outputs(3821));
    layer5_outputs(695) <= not((layer4_outputs(3055)) or (layer4_outputs(1700)));
    layer5_outputs(696) <= (layer4_outputs(4045)) and not (layer4_outputs(1163));
    layer5_outputs(697) <= layer4_outputs(7212);
    layer5_outputs(698) <= layer4_outputs(2453);
    layer5_outputs(699) <= layer4_outputs(1863);
    layer5_outputs(700) <= layer4_outputs(824);
    layer5_outputs(701) <= not((layer4_outputs(3183)) and (layer4_outputs(5529)));
    layer5_outputs(702) <= not((layer4_outputs(4228)) xor (layer4_outputs(5066)));
    layer5_outputs(703) <= layer4_outputs(4698);
    layer5_outputs(704) <= not((layer4_outputs(2909)) xor (layer4_outputs(464)));
    layer5_outputs(705) <= layer4_outputs(6111);
    layer5_outputs(706) <= (layer4_outputs(1680)) and not (layer4_outputs(4086));
    layer5_outputs(707) <= not(layer4_outputs(5333)) or (layer4_outputs(926));
    layer5_outputs(708) <= not(layer4_outputs(4509));
    layer5_outputs(709) <= not(layer4_outputs(6458)) or (layer4_outputs(7463));
    layer5_outputs(710) <= layer4_outputs(1960);
    layer5_outputs(711) <= layer4_outputs(4393);
    layer5_outputs(712) <= layer4_outputs(2538);
    layer5_outputs(713) <= layer4_outputs(5349);
    layer5_outputs(714) <= '0';
    layer5_outputs(715) <= not(layer4_outputs(4189));
    layer5_outputs(716) <= not(layer4_outputs(4922));
    layer5_outputs(717) <= layer4_outputs(460);
    layer5_outputs(718) <= layer4_outputs(2976);
    layer5_outputs(719) <= not(layer4_outputs(2102));
    layer5_outputs(720) <= not(layer4_outputs(275));
    layer5_outputs(721) <= (layer4_outputs(6557)) and (layer4_outputs(2316));
    layer5_outputs(722) <= (layer4_outputs(6307)) and (layer4_outputs(2566));
    layer5_outputs(723) <= not((layer4_outputs(1007)) and (layer4_outputs(3091)));
    layer5_outputs(724) <= layer4_outputs(4923);
    layer5_outputs(725) <= (layer4_outputs(2233)) and not (layer4_outputs(3435));
    layer5_outputs(726) <= not(layer4_outputs(446));
    layer5_outputs(727) <= (layer4_outputs(2073)) or (layer4_outputs(6325));
    layer5_outputs(728) <= layer4_outputs(6681);
    layer5_outputs(729) <= not(layer4_outputs(3390));
    layer5_outputs(730) <= not(layer4_outputs(2387));
    layer5_outputs(731) <= (layer4_outputs(2402)) and (layer4_outputs(3074));
    layer5_outputs(732) <= (layer4_outputs(5631)) or (layer4_outputs(5305));
    layer5_outputs(733) <= layer4_outputs(5697);
    layer5_outputs(734) <= not((layer4_outputs(6574)) xor (layer4_outputs(469)));
    layer5_outputs(735) <= not((layer4_outputs(1606)) or (layer4_outputs(3858)));
    layer5_outputs(736) <= not(layer4_outputs(5443)) or (layer4_outputs(276));
    layer5_outputs(737) <= layer4_outputs(5510);
    layer5_outputs(738) <= not(layer4_outputs(3329));
    layer5_outputs(739) <= '1';
    layer5_outputs(740) <= not(layer4_outputs(229)) or (layer4_outputs(1923));
    layer5_outputs(741) <= layer4_outputs(1184);
    layer5_outputs(742) <= not((layer4_outputs(3886)) or (layer4_outputs(6156)));
    layer5_outputs(743) <= not(layer4_outputs(178));
    layer5_outputs(744) <= not(layer4_outputs(7437)) or (layer4_outputs(5248));
    layer5_outputs(745) <= not(layer4_outputs(417));
    layer5_outputs(746) <= (layer4_outputs(5692)) or (layer4_outputs(955));
    layer5_outputs(747) <= not((layer4_outputs(3296)) xor (layer4_outputs(66)));
    layer5_outputs(748) <= (layer4_outputs(7045)) or (layer4_outputs(2501));
    layer5_outputs(749) <= layer4_outputs(5123);
    layer5_outputs(750) <= not(layer4_outputs(3449));
    layer5_outputs(751) <= layer4_outputs(1777);
    layer5_outputs(752) <= (layer4_outputs(802)) xor (layer4_outputs(4479));
    layer5_outputs(753) <= (layer4_outputs(4936)) or (layer4_outputs(2986));
    layer5_outputs(754) <= not(layer4_outputs(4693));
    layer5_outputs(755) <= not(layer4_outputs(5411)) or (layer4_outputs(3620));
    layer5_outputs(756) <= not(layer4_outputs(7604));
    layer5_outputs(757) <= not(layer4_outputs(3000));
    layer5_outputs(758) <= not(layer4_outputs(6282));
    layer5_outputs(759) <= layer4_outputs(316);
    layer5_outputs(760) <= layer4_outputs(2269);
    layer5_outputs(761) <= not(layer4_outputs(5111)) or (layer4_outputs(177));
    layer5_outputs(762) <= not(layer4_outputs(2766));
    layer5_outputs(763) <= (layer4_outputs(5729)) or (layer4_outputs(6973));
    layer5_outputs(764) <= layer4_outputs(2657);
    layer5_outputs(765) <= layer4_outputs(843);
    layer5_outputs(766) <= layer4_outputs(2380);
    layer5_outputs(767) <= not(layer4_outputs(697));
    layer5_outputs(768) <= layer4_outputs(2671);
    layer5_outputs(769) <= (layer4_outputs(1128)) and not (layer4_outputs(2774));
    layer5_outputs(770) <= layer4_outputs(4283);
    layer5_outputs(771) <= '1';
    layer5_outputs(772) <= (layer4_outputs(1421)) xor (layer4_outputs(903));
    layer5_outputs(773) <= not((layer4_outputs(3218)) and (layer4_outputs(5856)));
    layer5_outputs(774) <= layer4_outputs(828);
    layer5_outputs(775) <= not(layer4_outputs(219));
    layer5_outputs(776) <= (layer4_outputs(1558)) and not (layer4_outputs(6675));
    layer5_outputs(777) <= layer4_outputs(2031);
    layer5_outputs(778) <= layer4_outputs(5087);
    layer5_outputs(779) <= not(layer4_outputs(2769));
    layer5_outputs(780) <= layer4_outputs(6732);
    layer5_outputs(781) <= '1';
    layer5_outputs(782) <= not(layer4_outputs(7582)) or (layer4_outputs(4235));
    layer5_outputs(783) <= (layer4_outputs(4185)) xor (layer4_outputs(7077));
    layer5_outputs(784) <= not((layer4_outputs(1150)) xor (layer4_outputs(1073)));
    layer5_outputs(785) <= not(layer4_outputs(1775));
    layer5_outputs(786) <= layer4_outputs(4911);
    layer5_outputs(787) <= layer4_outputs(1383);
    layer5_outputs(788) <= '0';
    layer5_outputs(789) <= not((layer4_outputs(3532)) and (layer4_outputs(646)));
    layer5_outputs(790) <= not((layer4_outputs(5713)) or (layer4_outputs(5763)));
    layer5_outputs(791) <= '1';
    layer5_outputs(792) <= not(layer4_outputs(5106));
    layer5_outputs(793) <= layer4_outputs(4981);
    layer5_outputs(794) <= not((layer4_outputs(2789)) and (layer4_outputs(2158)));
    layer5_outputs(795) <= not(layer4_outputs(6482)) or (layer4_outputs(7443));
    layer5_outputs(796) <= not(layer4_outputs(2825)) or (layer4_outputs(6575));
    layer5_outputs(797) <= (layer4_outputs(6149)) and not (layer4_outputs(2024));
    layer5_outputs(798) <= not(layer4_outputs(6670)) or (layer4_outputs(2782));
    layer5_outputs(799) <= (layer4_outputs(1480)) xor (layer4_outputs(13));
    layer5_outputs(800) <= not(layer4_outputs(433));
    layer5_outputs(801) <= layer4_outputs(2071);
    layer5_outputs(802) <= not((layer4_outputs(4349)) and (layer4_outputs(7049)));
    layer5_outputs(803) <= (layer4_outputs(2585)) and not (layer4_outputs(1928));
    layer5_outputs(804) <= (layer4_outputs(1182)) and not (layer4_outputs(67));
    layer5_outputs(805) <= not(layer4_outputs(487));
    layer5_outputs(806) <= layer4_outputs(5910);
    layer5_outputs(807) <= layer4_outputs(2294);
    layer5_outputs(808) <= (layer4_outputs(5308)) xor (layer4_outputs(5708));
    layer5_outputs(809) <= layer4_outputs(5011);
    layer5_outputs(810) <= layer4_outputs(6663);
    layer5_outputs(811) <= not(layer4_outputs(2001));
    layer5_outputs(812) <= not(layer4_outputs(7172));
    layer5_outputs(813) <= not(layer4_outputs(5882));
    layer5_outputs(814) <= (layer4_outputs(2807)) and not (layer4_outputs(3894));
    layer5_outputs(815) <= (layer4_outputs(7370)) and (layer4_outputs(376));
    layer5_outputs(816) <= not((layer4_outputs(741)) or (layer4_outputs(3466)));
    layer5_outputs(817) <= not((layer4_outputs(2707)) or (layer4_outputs(1892)));
    layer5_outputs(818) <= (layer4_outputs(2600)) xor (layer4_outputs(1970));
    layer5_outputs(819) <= not(layer4_outputs(2009));
    layer5_outputs(820) <= not(layer4_outputs(1479)) or (layer4_outputs(5969));
    layer5_outputs(821) <= not((layer4_outputs(4352)) xor (layer4_outputs(1711)));
    layer5_outputs(822) <= layer4_outputs(1344);
    layer5_outputs(823) <= (layer4_outputs(4465)) and not (layer4_outputs(5048));
    layer5_outputs(824) <= (layer4_outputs(7601)) xor (layer4_outputs(6599));
    layer5_outputs(825) <= layer4_outputs(3899);
    layer5_outputs(826) <= (layer4_outputs(2882)) and not (layer4_outputs(2531));
    layer5_outputs(827) <= not((layer4_outputs(4964)) or (layer4_outputs(900)));
    layer5_outputs(828) <= not(layer4_outputs(2694));
    layer5_outputs(829) <= not(layer4_outputs(503)) or (layer4_outputs(5178));
    layer5_outputs(830) <= not(layer4_outputs(4497));
    layer5_outputs(831) <= not(layer4_outputs(7058));
    layer5_outputs(832) <= not(layer4_outputs(405));
    layer5_outputs(833) <= layer4_outputs(6995);
    layer5_outputs(834) <= layer4_outputs(5022);
    layer5_outputs(835) <= (layer4_outputs(5598)) and not (layer4_outputs(3682));
    layer5_outputs(836) <= (layer4_outputs(5718)) and not (layer4_outputs(5178));
    layer5_outputs(837) <= not(layer4_outputs(1957)) or (layer4_outputs(6559));
    layer5_outputs(838) <= not((layer4_outputs(6929)) xor (layer4_outputs(4144)));
    layer5_outputs(839) <= not(layer4_outputs(2870)) or (layer4_outputs(6568));
    layer5_outputs(840) <= layer4_outputs(6581);
    layer5_outputs(841) <= not(layer4_outputs(6081)) or (layer4_outputs(5762));
    layer5_outputs(842) <= (layer4_outputs(599)) and not (layer4_outputs(6945));
    layer5_outputs(843) <= (layer4_outputs(1552)) xor (layer4_outputs(1182));
    layer5_outputs(844) <= (layer4_outputs(3813)) and not (layer4_outputs(1245));
    layer5_outputs(845) <= not(layer4_outputs(5084));
    layer5_outputs(846) <= not((layer4_outputs(4854)) and (layer4_outputs(6612)));
    layer5_outputs(847) <= (layer4_outputs(2700)) xor (layer4_outputs(1869));
    layer5_outputs(848) <= layer4_outputs(4542);
    layer5_outputs(849) <= not(layer4_outputs(2297)) or (layer4_outputs(1742));
    layer5_outputs(850) <= layer4_outputs(4305);
    layer5_outputs(851) <= not(layer4_outputs(781));
    layer5_outputs(852) <= not(layer4_outputs(1937));
    layer5_outputs(853) <= not(layer4_outputs(1875)) or (layer4_outputs(1812));
    layer5_outputs(854) <= (layer4_outputs(765)) xor (layer4_outputs(6782));
    layer5_outputs(855) <= layer4_outputs(7108);
    layer5_outputs(856) <= not(layer4_outputs(2065));
    layer5_outputs(857) <= (layer4_outputs(4211)) xor (layer4_outputs(5124));
    layer5_outputs(858) <= not(layer4_outputs(1405));
    layer5_outputs(859) <= layer4_outputs(7581);
    layer5_outputs(860) <= layer4_outputs(4221);
    layer5_outputs(861) <= not((layer4_outputs(5402)) xor (layer4_outputs(5110)));
    layer5_outputs(862) <= not(layer4_outputs(6748));
    layer5_outputs(863) <= layer4_outputs(1361);
    layer5_outputs(864) <= not(layer4_outputs(1504));
    layer5_outputs(865) <= not(layer4_outputs(2833)) or (layer4_outputs(2520));
    layer5_outputs(866) <= (layer4_outputs(2883)) and not (layer4_outputs(3662));
    layer5_outputs(867) <= not((layer4_outputs(1897)) xor (layer4_outputs(7527)));
    layer5_outputs(868) <= not(layer4_outputs(6767));
    layer5_outputs(869) <= not(layer4_outputs(6215));
    layer5_outputs(870) <= layer4_outputs(111);
    layer5_outputs(871) <= not((layer4_outputs(2086)) xor (layer4_outputs(1018)));
    layer5_outputs(872) <= layer4_outputs(4208);
    layer5_outputs(873) <= (layer4_outputs(2541)) and not (layer4_outputs(6268));
    layer5_outputs(874) <= not(layer4_outputs(4399)) or (layer4_outputs(3153));
    layer5_outputs(875) <= (layer4_outputs(4220)) xor (layer4_outputs(6824));
    layer5_outputs(876) <= not(layer4_outputs(416)) or (layer4_outputs(6596));
    layer5_outputs(877) <= not(layer4_outputs(5103));
    layer5_outputs(878) <= not((layer4_outputs(2213)) and (layer4_outputs(4269)));
    layer5_outputs(879) <= not(layer4_outputs(3762));
    layer5_outputs(880) <= (layer4_outputs(6990)) or (layer4_outputs(581));
    layer5_outputs(881) <= '0';
    layer5_outputs(882) <= not(layer4_outputs(7116)) or (layer4_outputs(2492));
    layer5_outputs(883) <= not(layer4_outputs(4588)) or (layer4_outputs(93));
    layer5_outputs(884) <= not((layer4_outputs(5919)) xor (layer4_outputs(485)));
    layer5_outputs(885) <= (layer4_outputs(3686)) xor (layer4_outputs(1819));
    layer5_outputs(886) <= (layer4_outputs(5121)) and not (layer4_outputs(2787));
    layer5_outputs(887) <= not((layer4_outputs(3032)) xor (layer4_outputs(5437)));
    layer5_outputs(888) <= layer4_outputs(5772);
    layer5_outputs(889) <= (layer4_outputs(7021)) and (layer4_outputs(4424));
    layer5_outputs(890) <= not((layer4_outputs(7427)) xor (layer4_outputs(1714)));
    layer5_outputs(891) <= not(layer4_outputs(1976));
    layer5_outputs(892) <= not((layer4_outputs(1322)) or (layer4_outputs(2288)));
    layer5_outputs(893) <= layer4_outputs(1373);
    layer5_outputs(894) <= (layer4_outputs(4136)) and (layer4_outputs(5967));
    layer5_outputs(895) <= not((layer4_outputs(785)) or (layer4_outputs(3012)));
    layer5_outputs(896) <= not(layer4_outputs(4613)) or (layer4_outputs(5664));
    layer5_outputs(897) <= (layer4_outputs(3491)) and (layer4_outputs(2801));
    layer5_outputs(898) <= layer4_outputs(3938);
    layer5_outputs(899) <= (layer4_outputs(3168)) and not (layer4_outputs(5774));
    layer5_outputs(900) <= not((layer4_outputs(3952)) xor (layer4_outputs(247)));
    layer5_outputs(901) <= layer4_outputs(4067);
    layer5_outputs(902) <= not(layer4_outputs(2905));
    layer5_outputs(903) <= not(layer4_outputs(4488));
    layer5_outputs(904) <= layer4_outputs(1349);
    layer5_outputs(905) <= not(layer4_outputs(6177));
    layer5_outputs(906) <= (layer4_outputs(1931)) and not (layer4_outputs(4324));
    layer5_outputs(907) <= (layer4_outputs(5921)) and not (layer4_outputs(3076));
    layer5_outputs(908) <= (layer4_outputs(5610)) xor (layer4_outputs(2322));
    layer5_outputs(909) <= not(layer4_outputs(6909)) or (layer4_outputs(302));
    layer5_outputs(910) <= not(layer4_outputs(3043));
    layer5_outputs(911) <= not(layer4_outputs(4023));
    layer5_outputs(912) <= (layer4_outputs(6423)) xor (layer4_outputs(6154));
    layer5_outputs(913) <= (layer4_outputs(3366)) or (layer4_outputs(1807));
    layer5_outputs(914) <= (layer4_outputs(1238)) xor (layer4_outputs(944));
    layer5_outputs(915) <= not(layer4_outputs(5010)) or (layer4_outputs(6313));
    layer5_outputs(916) <= not(layer4_outputs(4725)) or (layer4_outputs(4926));
    layer5_outputs(917) <= (layer4_outputs(3528)) and not (layer4_outputs(3425));
    layer5_outputs(918) <= layer4_outputs(6169);
    layer5_outputs(919) <= layer4_outputs(6998);
    layer5_outputs(920) <= (layer4_outputs(1255)) or (layer4_outputs(4511));
    layer5_outputs(921) <= not((layer4_outputs(2478)) xor (layer4_outputs(105)));
    layer5_outputs(922) <= not(layer4_outputs(5491));
    layer5_outputs(923) <= (layer4_outputs(5464)) or (layer4_outputs(71));
    layer5_outputs(924) <= layer4_outputs(4413);
    layer5_outputs(925) <= layer4_outputs(4878);
    layer5_outputs(926) <= not(layer4_outputs(3011));
    layer5_outputs(927) <= (layer4_outputs(2058)) xor (layer4_outputs(5906));
    layer5_outputs(928) <= not((layer4_outputs(5250)) xor (layer4_outputs(5033)));
    layer5_outputs(929) <= not(layer4_outputs(6661));
    layer5_outputs(930) <= layer4_outputs(4832);
    layer5_outputs(931) <= (layer4_outputs(531)) and not (layer4_outputs(2586));
    layer5_outputs(932) <= not(layer4_outputs(6532)) or (layer4_outputs(2322));
    layer5_outputs(933) <= layer4_outputs(7302);
    layer5_outputs(934) <= (layer4_outputs(3117)) and not (layer4_outputs(6060));
    layer5_outputs(935) <= layer4_outputs(4889);
    layer5_outputs(936) <= layer4_outputs(6909);
    layer5_outputs(937) <= layer4_outputs(1642);
    layer5_outputs(938) <= not((layer4_outputs(3089)) xor (layer4_outputs(22)));
    layer5_outputs(939) <= (layer4_outputs(3535)) and not (layer4_outputs(7544));
    layer5_outputs(940) <= not(layer4_outputs(3167)) or (layer4_outputs(3610));
    layer5_outputs(941) <= (layer4_outputs(3298)) and not (layer4_outputs(4675));
    layer5_outputs(942) <= not((layer4_outputs(4767)) xor (layer4_outputs(1800)));
    layer5_outputs(943) <= not(layer4_outputs(4239));
    layer5_outputs(944) <= not(layer4_outputs(6511)) or (layer4_outputs(5871));
    layer5_outputs(945) <= (layer4_outputs(6559)) and not (layer4_outputs(4097));
    layer5_outputs(946) <= layer4_outputs(4224);
    layer5_outputs(947) <= not((layer4_outputs(4027)) and (layer4_outputs(1631)));
    layer5_outputs(948) <= layer4_outputs(1648);
    layer5_outputs(949) <= layer4_outputs(6562);
    layer5_outputs(950) <= not(layer4_outputs(738));
    layer5_outputs(951) <= not(layer4_outputs(5348)) or (layer4_outputs(2505));
    layer5_outputs(952) <= (layer4_outputs(6461)) xor (layer4_outputs(1074));
    layer5_outputs(953) <= not(layer4_outputs(3142));
    layer5_outputs(954) <= layer4_outputs(6538);
    layer5_outputs(955) <= not(layer4_outputs(4087));
    layer5_outputs(956) <= layer4_outputs(4364);
    layer5_outputs(957) <= not(layer4_outputs(6064)) or (layer4_outputs(3867));
    layer5_outputs(958) <= layer4_outputs(5252);
    layer5_outputs(959) <= (layer4_outputs(3462)) and (layer4_outputs(7073));
    layer5_outputs(960) <= not(layer4_outputs(6244));
    layer5_outputs(961) <= not((layer4_outputs(6499)) xor (layer4_outputs(5872)));
    layer5_outputs(962) <= layer4_outputs(1658);
    layer5_outputs(963) <= (layer4_outputs(2312)) xor (layer4_outputs(2755));
    layer5_outputs(964) <= (layer4_outputs(3124)) xor (layer4_outputs(1429));
    layer5_outputs(965) <= not((layer4_outputs(5236)) or (layer4_outputs(3879)));
    layer5_outputs(966) <= (layer4_outputs(6043)) xor (layer4_outputs(5931));
    layer5_outputs(967) <= layer4_outputs(860);
    layer5_outputs(968) <= (layer4_outputs(3751)) or (layer4_outputs(110));
    layer5_outputs(969) <= layer4_outputs(4312);
    layer5_outputs(970) <= not((layer4_outputs(6913)) xor (layer4_outputs(3847)));
    layer5_outputs(971) <= layer4_outputs(6950);
    layer5_outputs(972) <= layer4_outputs(1797);
    layer5_outputs(973) <= not(layer4_outputs(758));
    layer5_outputs(974) <= not((layer4_outputs(6389)) or (layer4_outputs(6078)));
    layer5_outputs(975) <= layer4_outputs(4938);
    layer5_outputs(976) <= layer4_outputs(4302);
    layer5_outputs(977) <= layer4_outputs(5099);
    layer5_outputs(978) <= not(layer4_outputs(4390)) or (layer4_outputs(5392));
    layer5_outputs(979) <= layer4_outputs(31);
    layer5_outputs(980) <= not((layer4_outputs(6915)) or (layer4_outputs(3873)));
    layer5_outputs(981) <= not(layer4_outputs(335));
    layer5_outputs(982) <= layer4_outputs(3096);
    layer5_outputs(983) <= (layer4_outputs(5211)) xor (layer4_outputs(6891));
    layer5_outputs(984) <= (layer4_outputs(225)) and not (layer4_outputs(3371));
    layer5_outputs(985) <= not(layer4_outputs(3120));
    layer5_outputs(986) <= layer4_outputs(3031);
    layer5_outputs(987) <= '1';
    layer5_outputs(988) <= not(layer4_outputs(950));
    layer5_outputs(989) <= layer4_outputs(1542);
    layer5_outputs(990) <= not(layer4_outputs(7428)) or (layer4_outputs(1939));
    layer5_outputs(991) <= (layer4_outputs(7624)) or (layer4_outputs(4295));
    layer5_outputs(992) <= not(layer4_outputs(699));
    layer5_outputs(993) <= not(layer4_outputs(5223));
    layer5_outputs(994) <= not(layer4_outputs(647)) or (layer4_outputs(6132));
    layer5_outputs(995) <= (layer4_outputs(6765)) and not (layer4_outputs(4546));
    layer5_outputs(996) <= (layer4_outputs(4540)) xor (layer4_outputs(3354));
    layer5_outputs(997) <= layer4_outputs(6433);
    layer5_outputs(998) <= not(layer4_outputs(4551));
    layer5_outputs(999) <= not((layer4_outputs(5446)) xor (layer4_outputs(1705)));
    layer5_outputs(1000) <= not((layer4_outputs(1675)) or (layer4_outputs(7544)));
    layer5_outputs(1001) <= not((layer4_outputs(7558)) xor (layer4_outputs(3099)));
    layer5_outputs(1002) <= layer4_outputs(7411);
    layer5_outputs(1003) <= not(layer4_outputs(2378));
    layer5_outputs(1004) <= layer4_outputs(41);
    layer5_outputs(1005) <= '0';
    layer5_outputs(1006) <= not((layer4_outputs(1107)) or (layer4_outputs(2764)));
    layer5_outputs(1007) <= layer4_outputs(1355);
    layer5_outputs(1008) <= not(layer4_outputs(6334));
    layer5_outputs(1009) <= not(layer4_outputs(2172));
    layer5_outputs(1010) <= not(layer4_outputs(2138));
    layer5_outputs(1011) <= not(layer4_outputs(1813));
    layer5_outputs(1012) <= layer4_outputs(1755);
    layer5_outputs(1013) <= '1';
    layer5_outputs(1014) <= (layer4_outputs(6185)) and not (layer4_outputs(1992));
    layer5_outputs(1015) <= not(layer4_outputs(3819));
    layer5_outputs(1016) <= (layer4_outputs(4289)) xor (layer4_outputs(3714));
    layer5_outputs(1017) <= not(layer4_outputs(6262));
    layer5_outputs(1018) <= (layer4_outputs(2796)) or (layer4_outputs(3091));
    layer5_outputs(1019) <= not(layer4_outputs(3916)) or (layer4_outputs(1769));
    layer5_outputs(1020) <= not(layer4_outputs(4219));
    layer5_outputs(1021) <= not(layer4_outputs(4917));
    layer5_outputs(1022) <= not(layer4_outputs(1829));
    layer5_outputs(1023) <= not(layer4_outputs(5746));
    layer5_outputs(1024) <= not(layer4_outputs(4381));
    layer5_outputs(1025) <= layer4_outputs(6174);
    layer5_outputs(1026) <= (layer4_outputs(2146)) and not (layer4_outputs(1086));
    layer5_outputs(1027) <= layer4_outputs(6121);
    layer5_outputs(1028) <= (layer4_outputs(3683)) and (layer4_outputs(2840));
    layer5_outputs(1029) <= not(layer4_outputs(5968));
    layer5_outputs(1030) <= not(layer4_outputs(3228));
    layer5_outputs(1031) <= not(layer4_outputs(4802));
    layer5_outputs(1032) <= not((layer4_outputs(1715)) or (layer4_outputs(2061)));
    layer5_outputs(1033) <= not(layer4_outputs(1189));
    layer5_outputs(1034) <= layer4_outputs(5649);
    layer5_outputs(1035) <= not(layer4_outputs(6201)) or (layer4_outputs(3496));
    layer5_outputs(1036) <= not(layer4_outputs(5357));
    layer5_outputs(1037) <= not((layer4_outputs(1027)) xor (layer4_outputs(7529)));
    layer5_outputs(1038) <= not((layer4_outputs(7195)) and (layer4_outputs(472)));
    layer5_outputs(1039) <= not(layer4_outputs(96));
    layer5_outputs(1040) <= layer4_outputs(4212);
    layer5_outputs(1041) <= (layer4_outputs(77)) or (layer4_outputs(7265));
    layer5_outputs(1042) <= layer4_outputs(5344);
    layer5_outputs(1043) <= (layer4_outputs(1237)) and not (layer4_outputs(2792));
    layer5_outputs(1044) <= layer4_outputs(3810);
    layer5_outputs(1045) <= '0';
    layer5_outputs(1046) <= not(layer4_outputs(2045));
    layer5_outputs(1047) <= not(layer4_outputs(5453));
    layer5_outputs(1048) <= (layer4_outputs(2776)) or (layer4_outputs(4430));
    layer5_outputs(1049) <= (layer4_outputs(258)) or (layer4_outputs(7612));
    layer5_outputs(1050) <= not(layer4_outputs(5096));
    layer5_outputs(1051) <= (layer4_outputs(120)) and not (layer4_outputs(747));
    layer5_outputs(1052) <= (layer4_outputs(6056)) and (layer4_outputs(6733));
    layer5_outputs(1053) <= not(layer4_outputs(1328));
    layer5_outputs(1054) <= not(layer4_outputs(2764));
    layer5_outputs(1055) <= not((layer4_outputs(5)) and (layer4_outputs(1564)));
    layer5_outputs(1056) <= not(layer4_outputs(1536));
    layer5_outputs(1057) <= not((layer4_outputs(5070)) and (layer4_outputs(1450)));
    layer5_outputs(1058) <= not(layer4_outputs(1908));
    layer5_outputs(1059) <= not((layer4_outputs(4410)) and (layer4_outputs(7087)));
    layer5_outputs(1060) <= not(layer4_outputs(4945));
    layer5_outputs(1061) <= (layer4_outputs(1147)) and not (layer4_outputs(2281));
    layer5_outputs(1062) <= (layer4_outputs(3526)) and (layer4_outputs(3097));
    layer5_outputs(1063) <= layer4_outputs(4256);
    layer5_outputs(1064) <= not(layer4_outputs(3483));
    layer5_outputs(1065) <= not(layer4_outputs(5677));
    layer5_outputs(1066) <= layer4_outputs(7295);
    layer5_outputs(1067) <= (layer4_outputs(6655)) and (layer4_outputs(3547));
    layer5_outputs(1068) <= not(layer4_outputs(1246));
    layer5_outputs(1069) <= (layer4_outputs(5859)) xor (layer4_outputs(6839));
    layer5_outputs(1070) <= not((layer4_outputs(5961)) xor (layer4_outputs(911)));
    layer5_outputs(1071) <= not(layer4_outputs(2052));
    layer5_outputs(1072) <= not((layer4_outputs(58)) xor (layer4_outputs(2765)));
    layer5_outputs(1073) <= (layer4_outputs(1769)) or (layer4_outputs(1222));
    layer5_outputs(1074) <= not(layer4_outputs(4272));
    layer5_outputs(1075) <= (layer4_outputs(3024)) xor (layer4_outputs(2194));
    layer5_outputs(1076) <= (layer4_outputs(7510)) and (layer4_outputs(6056));
    layer5_outputs(1077) <= not(layer4_outputs(2411));
    layer5_outputs(1078) <= not(layer4_outputs(3230));
    layer5_outputs(1079) <= layer4_outputs(927);
    layer5_outputs(1080) <= (layer4_outputs(6555)) and not (layer4_outputs(754));
    layer5_outputs(1081) <= not((layer4_outputs(3208)) xor (layer4_outputs(274)));
    layer5_outputs(1082) <= layer4_outputs(3401);
    layer5_outputs(1083) <= not((layer4_outputs(2025)) or (layer4_outputs(20)));
    layer5_outputs(1084) <= not(layer4_outputs(5629));
    layer5_outputs(1085) <= (layer4_outputs(7257)) xor (layer4_outputs(7401));
    layer5_outputs(1086) <= '0';
    layer5_outputs(1087) <= not(layer4_outputs(4010));
    layer5_outputs(1088) <= not((layer4_outputs(7442)) or (layer4_outputs(1053)));
    layer5_outputs(1089) <= layer4_outputs(1732);
    layer5_outputs(1090) <= layer4_outputs(2059);
    layer5_outputs(1091) <= not((layer4_outputs(7018)) or (layer4_outputs(800)));
    layer5_outputs(1092) <= not((layer4_outputs(505)) xor (layer4_outputs(5945)));
    layer5_outputs(1093) <= not(layer4_outputs(1978));
    layer5_outputs(1094) <= not(layer4_outputs(773)) or (layer4_outputs(488));
    layer5_outputs(1095) <= not(layer4_outputs(3203));
    layer5_outputs(1096) <= layer4_outputs(6968);
    layer5_outputs(1097) <= layer4_outputs(2482);
    layer5_outputs(1098) <= (layer4_outputs(3560)) xor (layer4_outputs(6997));
    layer5_outputs(1099) <= not(layer4_outputs(734));
    layer5_outputs(1100) <= layer4_outputs(1413);
    layer5_outputs(1101) <= not(layer4_outputs(6344));
    layer5_outputs(1102) <= layer4_outputs(213);
    layer5_outputs(1103) <= not(layer4_outputs(3814));
    layer5_outputs(1104) <= (layer4_outputs(6905)) and (layer4_outputs(7615));
    layer5_outputs(1105) <= layer4_outputs(7393);
    layer5_outputs(1106) <= (layer4_outputs(6384)) and (layer4_outputs(5720));
    layer5_outputs(1107) <= (layer4_outputs(5485)) xor (layer4_outputs(304));
    layer5_outputs(1108) <= layer4_outputs(2502);
    layer5_outputs(1109) <= not(layer4_outputs(3471));
    layer5_outputs(1110) <= (layer4_outputs(3579)) or (layer4_outputs(6347));
    layer5_outputs(1111) <= layer4_outputs(1452);
    layer5_outputs(1112) <= not((layer4_outputs(2778)) xor (layer4_outputs(1598)));
    layer5_outputs(1113) <= layer4_outputs(417);
    layer5_outputs(1114) <= layer4_outputs(1627);
    layer5_outputs(1115) <= layer4_outputs(2168);
    layer5_outputs(1116) <= (layer4_outputs(6688)) and not (layer4_outputs(6081));
    layer5_outputs(1117) <= (layer4_outputs(2012)) and not (layer4_outputs(1443));
    layer5_outputs(1118) <= not(layer4_outputs(4345)) or (layer4_outputs(1179));
    layer5_outputs(1119) <= layer4_outputs(802);
    layer5_outputs(1120) <= (layer4_outputs(1022)) or (layer4_outputs(514));
    layer5_outputs(1121) <= (layer4_outputs(5637)) xor (layer4_outputs(4697));
    layer5_outputs(1122) <= not(layer4_outputs(6698));
    layer5_outputs(1123) <= layer4_outputs(4315);
    layer5_outputs(1124) <= not(layer4_outputs(3722));
    layer5_outputs(1125) <= '1';
    layer5_outputs(1126) <= not(layer4_outputs(2150));
    layer5_outputs(1127) <= not((layer4_outputs(7205)) xor (layer4_outputs(3764)));
    layer5_outputs(1128) <= (layer4_outputs(6286)) and (layer4_outputs(3174));
    layer5_outputs(1129) <= layer4_outputs(5806);
    layer5_outputs(1130) <= layer4_outputs(4228);
    layer5_outputs(1131) <= layer4_outputs(695);
    layer5_outputs(1132) <= layer4_outputs(6217);
    layer5_outputs(1133) <= (layer4_outputs(2604)) and (layer4_outputs(2337));
    layer5_outputs(1134) <= not(layer4_outputs(6898));
    layer5_outputs(1135) <= layer4_outputs(4435);
    layer5_outputs(1136) <= not((layer4_outputs(79)) xor (layer4_outputs(5298)));
    layer5_outputs(1137) <= layer4_outputs(2283);
    layer5_outputs(1138) <= not(layer4_outputs(6703));
    layer5_outputs(1139) <= not(layer4_outputs(1000));
    layer5_outputs(1140) <= not(layer4_outputs(2940));
    layer5_outputs(1141) <= (layer4_outputs(1858)) and (layer4_outputs(1969));
    layer5_outputs(1142) <= (layer4_outputs(6916)) and (layer4_outputs(1326));
    layer5_outputs(1143) <= not(layer4_outputs(3534));
    layer5_outputs(1144) <= not(layer4_outputs(6643));
    layer5_outputs(1145) <= (layer4_outputs(1259)) and not (layer4_outputs(6259));
    layer5_outputs(1146) <= not(layer4_outputs(2262)) or (layer4_outputs(4154));
    layer5_outputs(1147) <= (layer4_outputs(6859)) or (layer4_outputs(4583));
    layer5_outputs(1148) <= (layer4_outputs(7488)) or (layer4_outputs(3243));
    layer5_outputs(1149) <= not((layer4_outputs(5030)) xor (layer4_outputs(235)));
    layer5_outputs(1150) <= not(layer4_outputs(4361));
    layer5_outputs(1151) <= not((layer4_outputs(5746)) and (layer4_outputs(4844)));
    layer5_outputs(1152) <= not(layer4_outputs(1470));
    layer5_outputs(1153) <= layer4_outputs(4939);
    layer5_outputs(1154) <= (layer4_outputs(4802)) and (layer4_outputs(63));
    layer5_outputs(1155) <= (layer4_outputs(737)) and (layer4_outputs(2592));
    layer5_outputs(1156) <= not((layer4_outputs(3873)) xor (layer4_outputs(3440)));
    layer5_outputs(1157) <= (layer4_outputs(5429)) and (layer4_outputs(781));
    layer5_outputs(1158) <= (layer4_outputs(2500)) or (layer4_outputs(4827));
    layer5_outputs(1159) <= not(layer4_outputs(6391)) or (layer4_outputs(3689));
    layer5_outputs(1160) <= (layer4_outputs(7435)) or (layer4_outputs(4571));
    layer5_outputs(1161) <= not((layer4_outputs(2983)) xor (layer4_outputs(286)));
    layer5_outputs(1162) <= not(layer4_outputs(3185));
    layer5_outputs(1163) <= not(layer4_outputs(316)) or (layer4_outputs(4607));
    layer5_outputs(1164) <= (layer4_outputs(6937)) or (layer4_outputs(311));
    layer5_outputs(1165) <= (layer4_outputs(2654)) and not (layer4_outputs(4649));
    layer5_outputs(1166) <= (layer4_outputs(5512)) or (layer4_outputs(129));
    layer5_outputs(1167) <= layer4_outputs(6652);
    layer5_outputs(1168) <= not((layer4_outputs(4939)) xor (layer4_outputs(2519)));
    layer5_outputs(1169) <= not(layer4_outputs(6885)) or (layer4_outputs(1021));
    layer5_outputs(1170) <= (layer4_outputs(3369)) xor (layer4_outputs(3920));
    layer5_outputs(1171) <= not((layer4_outputs(986)) xor (layer4_outputs(2586)));
    layer5_outputs(1172) <= not(layer4_outputs(4378));
    layer5_outputs(1173) <= not(layer4_outputs(7198)) or (layer4_outputs(5861));
    layer5_outputs(1174) <= not((layer4_outputs(333)) xor (layer4_outputs(5105)));
    layer5_outputs(1175) <= not(layer4_outputs(5648)) or (layer4_outputs(1199));
    layer5_outputs(1176) <= layer4_outputs(4865);
    layer5_outputs(1177) <= not(layer4_outputs(4167));
    layer5_outputs(1178) <= not((layer4_outputs(6057)) and (layer4_outputs(2907)));
    layer5_outputs(1179) <= (layer4_outputs(4706)) and not (layer4_outputs(3353));
    layer5_outputs(1180) <= '0';
    layer5_outputs(1181) <= layer4_outputs(1434);
    layer5_outputs(1182) <= not(layer4_outputs(4467));
    layer5_outputs(1183) <= not(layer4_outputs(3272));
    layer5_outputs(1184) <= (layer4_outputs(3702)) and not (layer4_outputs(4354));
    layer5_outputs(1185) <= not(layer4_outputs(7121));
    layer5_outputs(1186) <= not(layer4_outputs(2697)) or (layer4_outputs(5551));
    layer5_outputs(1187) <= layer4_outputs(2617);
    layer5_outputs(1188) <= not(layer4_outputs(5470)) or (layer4_outputs(4398));
    layer5_outputs(1189) <= not((layer4_outputs(1818)) or (layer4_outputs(1508)));
    layer5_outputs(1190) <= not((layer4_outputs(3790)) and (layer4_outputs(261)));
    layer5_outputs(1191) <= (layer4_outputs(543)) and not (layer4_outputs(1369));
    layer5_outputs(1192) <= layer4_outputs(995);
    layer5_outputs(1193) <= (layer4_outputs(2417)) or (layer4_outputs(3843));
    layer5_outputs(1194) <= not(layer4_outputs(7492));
    layer5_outputs(1195) <= (layer4_outputs(5867)) xor (layer4_outputs(4291));
    layer5_outputs(1196) <= '1';
    layer5_outputs(1197) <= not(layer4_outputs(4635));
    layer5_outputs(1198) <= not(layer4_outputs(1074)) or (layer4_outputs(4320));
    layer5_outputs(1199) <= (layer4_outputs(7023)) or (layer4_outputs(3845));
    layer5_outputs(1200) <= (layer4_outputs(1891)) and (layer4_outputs(5686));
    layer5_outputs(1201) <= not((layer4_outputs(1540)) and (layer4_outputs(5994)));
    layer5_outputs(1202) <= layer4_outputs(878);
    layer5_outputs(1203) <= not(layer4_outputs(4384));
    layer5_outputs(1204) <= not(layer4_outputs(3803));
    layer5_outputs(1205) <= layer4_outputs(7277);
    layer5_outputs(1206) <= layer4_outputs(1850);
    layer5_outputs(1207) <= layer4_outputs(3857);
    layer5_outputs(1208) <= not((layer4_outputs(5567)) and (layer4_outputs(1355)));
    layer5_outputs(1209) <= not(layer4_outputs(3676));
    layer5_outputs(1210) <= (layer4_outputs(415)) xor (layer4_outputs(217));
    layer5_outputs(1211) <= layer4_outputs(209);
    layer5_outputs(1212) <= (layer4_outputs(5914)) xor (layer4_outputs(4455));
    layer5_outputs(1213) <= layer4_outputs(2621);
    layer5_outputs(1214) <= (layer4_outputs(2104)) or (layer4_outputs(5552));
    layer5_outputs(1215) <= not(layer4_outputs(4903));
    layer5_outputs(1216) <= layer4_outputs(1225);
    layer5_outputs(1217) <= not(layer4_outputs(808)) or (layer4_outputs(6579));
    layer5_outputs(1218) <= (layer4_outputs(3646)) or (layer4_outputs(7004));
    layer5_outputs(1219) <= layer4_outputs(7385);
    layer5_outputs(1220) <= (layer4_outputs(6203)) and (layer4_outputs(6278));
    layer5_outputs(1221) <= not(layer4_outputs(6827)) or (layer4_outputs(750));
    layer5_outputs(1222) <= not(layer4_outputs(5595));
    layer5_outputs(1223) <= not(layer4_outputs(6186));
    layer5_outputs(1224) <= layer4_outputs(1215);
    layer5_outputs(1225) <= not(layer4_outputs(4800));
    layer5_outputs(1226) <= not(layer4_outputs(687));
    layer5_outputs(1227) <= layer4_outputs(3067);
    layer5_outputs(1228) <= not((layer4_outputs(4598)) xor (layer4_outputs(4208)));
    layer5_outputs(1229) <= layer4_outputs(2346);
    layer5_outputs(1230) <= (layer4_outputs(3525)) and (layer4_outputs(1651));
    layer5_outputs(1231) <= (layer4_outputs(6818)) and (layer4_outputs(1842));
    layer5_outputs(1232) <= not(layer4_outputs(5075));
    layer5_outputs(1233) <= not((layer4_outputs(4037)) xor (layer4_outputs(1512)));
    layer5_outputs(1234) <= (layer4_outputs(1090)) xor (layer4_outputs(6112));
    layer5_outputs(1235) <= layer4_outputs(3620);
    layer5_outputs(1236) <= not(layer4_outputs(1721));
    layer5_outputs(1237) <= '1';
    layer5_outputs(1238) <= not(layer4_outputs(4468)) or (layer4_outputs(2076));
    layer5_outputs(1239) <= layer4_outputs(5716);
    layer5_outputs(1240) <= not((layer4_outputs(2250)) xor (layer4_outputs(959)));
    layer5_outputs(1241) <= not((layer4_outputs(7220)) and (layer4_outputs(7307)));
    layer5_outputs(1242) <= not((layer4_outputs(3594)) and (layer4_outputs(4985)));
    layer5_outputs(1243) <= not(layer4_outputs(264)) or (layer4_outputs(19));
    layer5_outputs(1244) <= not((layer4_outputs(3549)) and (layer4_outputs(2046)));
    layer5_outputs(1245) <= not(layer4_outputs(794)) or (layer4_outputs(1180));
    layer5_outputs(1246) <= (layer4_outputs(6239)) xor (layer4_outputs(6435));
    layer5_outputs(1247) <= not((layer4_outputs(1435)) xor (layer4_outputs(470)));
    layer5_outputs(1248) <= not(layer4_outputs(462)) or (layer4_outputs(6302));
    layer5_outputs(1249) <= not((layer4_outputs(6363)) xor (layer4_outputs(1162)));
    layer5_outputs(1250) <= (layer4_outputs(102)) or (layer4_outputs(1402));
    layer5_outputs(1251) <= not(layer4_outputs(5778)) or (layer4_outputs(4484));
    layer5_outputs(1252) <= not(layer4_outputs(4765));
    layer5_outputs(1253) <= layer4_outputs(3983);
    layer5_outputs(1254) <= not(layer4_outputs(4057)) or (layer4_outputs(1728));
    layer5_outputs(1255) <= not(layer4_outputs(5826));
    layer5_outputs(1256) <= (layer4_outputs(3092)) or (layer4_outputs(5204));
    layer5_outputs(1257) <= layer4_outputs(4352);
    layer5_outputs(1258) <= not((layer4_outputs(1003)) or (layer4_outputs(3621)));
    layer5_outputs(1259) <= layer4_outputs(4258);
    layer5_outputs(1260) <= not(layer4_outputs(6747));
    layer5_outputs(1261) <= (layer4_outputs(5844)) xor (layer4_outputs(634));
    layer5_outputs(1262) <= layer4_outputs(7352);
    layer5_outputs(1263) <= not(layer4_outputs(4263));
    layer5_outputs(1264) <= not(layer4_outputs(6963));
    layer5_outputs(1265) <= not((layer4_outputs(5754)) and (layer4_outputs(3565)));
    layer5_outputs(1266) <= layer4_outputs(7586);
    layer5_outputs(1267) <= not(layer4_outputs(4708));
    layer5_outputs(1268) <= not((layer4_outputs(2509)) or (layer4_outputs(1194)));
    layer5_outputs(1269) <= (layer4_outputs(3986)) xor (layer4_outputs(770));
    layer5_outputs(1270) <= not(layer4_outputs(280));
    layer5_outputs(1271) <= not(layer4_outputs(4686));
    layer5_outputs(1272) <= (layer4_outputs(7610)) and not (layer4_outputs(2215));
    layer5_outputs(1273) <= not(layer4_outputs(1955)) or (layer4_outputs(6977));
    layer5_outputs(1274) <= not(layer4_outputs(7631)) or (layer4_outputs(1125));
    layer5_outputs(1275) <= (layer4_outputs(4788)) and (layer4_outputs(5847));
    layer5_outputs(1276) <= layer4_outputs(1255);
    layer5_outputs(1277) <= '1';
    layer5_outputs(1278) <= (layer4_outputs(4287)) or (layer4_outputs(4068));
    layer5_outputs(1279) <= not(layer4_outputs(7029));
    layer5_outputs(1280) <= (layer4_outputs(4963)) or (layer4_outputs(1183));
    layer5_outputs(1281) <= not((layer4_outputs(5977)) or (layer4_outputs(4689)));
    layer5_outputs(1282) <= not((layer4_outputs(251)) xor (layer4_outputs(2115)));
    layer5_outputs(1283) <= layer4_outputs(2706);
    layer5_outputs(1284) <= not((layer4_outputs(5776)) xor (layer4_outputs(4733)));
    layer5_outputs(1285) <= layer4_outputs(4760);
    layer5_outputs(1286) <= not(layer4_outputs(7539));
    layer5_outputs(1287) <= not(layer4_outputs(300));
    layer5_outputs(1288) <= not(layer4_outputs(4314));
    layer5_outputs(1289) <= not(layer4_outputs(213));
    layer5_outputs(1290) <= layer4_outputs(2234);
    layer5_outputs(1291) <= not(layer4_outputs(2425));
    layer5_outputs(1292) <= (layer4_outputs(7374)) and not (layer4_outputs(6884));
    layer5_outputs(1293) <= (layer4_outputs(3618)) xor (layer4_outputs(4706));
    layer5_outputs(1294) <= (layer4_outputs(6032)) or (layer4_outputs(3506));
    layer5_outputs(1295) <= not((layer4_outputs(4526)) xor (layer4_outputs(5911)));
    layer5_outputs(1296) <= '1';
    layer5_outputs(1297) <= layer4_outputs(3692);
    layer5_outputs(1298) <= (layer4_outputs(4969)) and (layer4_outputs(2123));
    layer5_outputs(1299) <= layer4_outputs(481);
    layer5_outputs(1300) <= (layer4_outputs(5878)) and (layer4_outputs(4355));
    layer5_outputs(1301) <= not((layer4_outputs(3472)) and (layer4_outputs(1146)));
    layer5_outputs(1302) <= not((layer4_outputs(2159)) or (layer4_outputs(2096)));
    layer5_outputs(1303) <= (layer4_outputs(3668)) and (layer4_outputs(1890));
    layer5_outputs(1304) <= (layer4_outputs(2483)) and not (layer4_outputs(3598));
    layer5_outputs(1305) <= not(layer4_outputs(4831));
    layer5_outputs(1306) <= not(layer4_outputs(3323));
    layer5_outputs(1307) <= layer4_outputs(6247);
    layer5_outputs(1308) <= not(layer4_outputs(3276));
    layer5_outputs(1309) <= not(layer4_outputs(7194)) or (layer4_outputs(3693));
    layer5_outputs(1310) <= not(layer4_outputs(3148)) or (layer4_outputs(5411));
    layer5_outputs(1311) <= not(layer4_outputs(500));
    layer5_outputs(1312) <= not(layer4_outputs(387)) or (layer4_outputs(3635));
    layer5_outputs(1313) <= (layer4_outputs(4274)) and (layer4_outputs(4113));
    layer5_outputs(1314) <= layer4_outputs(958);
    layer5_outputs(1315) <= not(layer4_outputs(2942)) or (layer4_outputs(5230));
    layer5_outputs(1316) <= not(layer4_outputs(7423));
    layer5_outputs(1317) <= (layer4_outputs(6833)) xor (layer4_outputs(789));
    layer5_outputs(1318) <= not(layer4_outputs(147));
    layer5_outputs(1319) <= layer4_outputs(219);
    layer5_outputs(1320) <= not(layer4_outputs(1267));
    layer5_outputs(1321) <= layer4_outputs(5586);
    layer5_outputs(1322) <= not(layer4_outputs(4660));
    layer5_outputs(1323) <= layer4_outputs(7088);
    layer5_outputs(1324) <= (layer4_outputs(6463)) or (layer4_outputs(4038));
    layer5_outputs(1325) <= (layer4_outputs(4135)) and not (layer4_outputs(6648));
    layer5_outputs(1326) <= (layer4_outputs(7635)) or (layer4_outputs(159));
    layer5_outputs(1327) <= '1';
    layer5_outputs(1328) <= not((layer4_outputs(5283)) and (layer4_outputs(5634)));
    layer5_outputs(1329) <= layer4_outputs(4423);
    layer5_outputs(1330) <= (layer4_outputs(4331)) and not (layer4_outputs(2559));
    layer5_outputs(1331) <= not(layer4_outputs(3154)) or (layer4_outputs(1035));
    layer5_outputs(1332) <= not(layer4_outputs(3691));
    layer5_outputs(1333) <= not(layer4_outputs(2448));
    layer5_outputs(1334) <= not(layer4_outputs(4905));
    layer5_outputs(1335) <= (layer4_outputs(7408)) and not (layer4_outputs(3204));
    layer5_outputs(1336) <= not(layer4_outputs(1572));
    layer5_outputs(1337) <= not(layer4_outputs(4074)) or (layer4_outputs(4473));
    layer5_outputs(1338) <= not(layer4_outputs(4002));
    layer5_outputs(1339) <= (layer4_outputs(5688)) or (layer4_outputs(5669));
    layer5_outputs(1340) <= not(layer4_outputs(2517)) or (layer4_outputs(5575));
    layer5_outputs(1341) <= not(layer4_outputs(5691));
    layer5_outputs(1342) <= (layer4_outputs(2733)) and not (layer4_outputs(6421));
    layer5_outputs(1343) <= not((layer4_outputs(369)) or (layer4_outputs(2740)));
    layer5_outputs(1344) <= not(layer4_outputs(2329));
    layer5_outputs(1345) <= not(layer4_outputs(3098));
    layer5_outputs(1346) <= '1';
    layer5_outputs(1347) <= layer4_outputs(3108);
    layer5_outputs(1348) <= (layer4_outputs(1164)) xor (layer4_outputs(1338));
    layer5_outputs(1349) <= not(layer4_outputs(3988));
    layer5_outputs(1350) <= not((layer4_outputs(5917)) xor (layer4_outputs(2160)));
    layer5_outputs(1351) <= layer4_outputs(2342);
    layer5_outputs(1352) <= not(layer4_outputs(872));
    layer5_outputs(1353) <= layer4_outputs(6066);
    layer5_outputs(1354) <= (layer4_outputs(4153)) and not (layer4_outputs(5969));
    layer5_outputs(1355) <= '0';
    layer5_outputs(1356) <= not(layer4_outputs(552)) or (layer4_outputs(5086));
    layer5_outputs(1357) <= not(layer4_outputs(44));
    layer5_outputs(1358) <= not(layer4_outputs(3249));
    layer5_outputs(1359) <= layer4_outputs(545);
    layer5_outputs(1360) <= not(layer4_outputs(402));
    layer5_outputs(1361) <= (layer4_outputs(1101)) or (layer4_outputs(4404));
    layer5_outputs(1362) <= not(layer4_outputs(2209));
    layer5_outputs(1363) <= layer4_outputs(2337);
    layer5_outputs(1364) <= not(layer4_outputs(7132));
    layer5_outputs(1365) <= layer4_outputs(4506);
    layer5_outputs(1366) <= (layer4_outputs(5488)) and (layer4_outputs(1673));
    layer5_outputs(1367) <= layer4_outputs(27);
    layer5_outputs(1368) <= not(layer4_outputs(3788));
    layer5_outputs(1369) <= not(layer4_outputs(6351));
    layer5_outputs(1370) <= not((layer4_outputs(4009)) and (layer4_outputs(6908)));
    layer5_outputs(1371) <= layer4_outputs(4816);
    layer5_outputs(1372) <= not((layer4_outputs(1603)) xor (layer4_outputs(6178)));
    layer5_outputs(1373) <= layer4_outputs(2746);
    layer5_outputs(1374) <= (layer4_outputs(2370)) xor (layer4_outputs(3736));
    layer5_outputs(1375) <= not(layer4_outputs(1862));
    layer5_outputs(1376) <= not((layer4_outputs(1903)) xor (layer4_outputs(1531)));
    layer5_outputs(1377) <= not((layer4_outputs(3407)) and (layer4_outputs(6763)));
    layer5_outputs(1378) <= layer4_outputs(6233);
    layer5_outputs(1379) <= (layer4_outputs(1030)) or (layer4_outputs(6108));
    layer5_outputs(1380) <= not((layer4_outputs(5025)) or (layer4_outputs(6570)));
    layer5_outputs(1381) <= layer4_outputs(1667);
    layer5_outputs(1382) <= not(layer4_outputs(2356)) or (layer4_outputs(5292));
    layer5_outputs(1383) <= not(layer4_outputs(709));
    layer5_outputs(1384) <= not(layer4_outputs(553));
    layer5_outputs(1385) <= layer4_outputs(3822);
    layer5_outputs(1386) <= (layer4_outputs(5460)) and (layer4_outputs(69));
    layer5_outputs(1387) <= not(layer4_outputs(5725));
    layer5_outputs(1388) <= (layer4_outputs(6143)) and not (layer4_outputs(409));
    layer5_outputs(1389) <= layer4_outputs(5225);
    layer5_outputs(1390) <= not(layer4_outputs(7561)) or (layer4_outputs(3795));
    layer5_outputs(1391) <= not((layer4_outputs(4813)) or (layer4_outputs(7348)));
    layer5_outputs(1392) <= not(layer4_outputs(7020));
    layer5_outputs(1393) <= not(layer4_outputs(7483));
    layer5_outputs(1394) <= not(layer4_outputs(3449));
    layer5_outputs(1395) <= (layer4_outputs(2618)) and (layer4_outputs(7025));
    layer5_outputs(1396) <= layer4_outputs(906);
    layer5_outputs(1397) <= layer4_outputs(7572);
    layer5_outputs(1398) <= not(layer4_outputs(3292)) or (layer4_outputs(200));
    layer5_outputs(1399) <= not(layer4_outputs(7093));
    layer5_outputs(1400) <= layer4_outputs(1778);
    layer5_outputs(1401) <= not(layer4_outputs(3322)) or (layer4_outputs(6304));
    layer5_outputs(1402) <= (layer4_outputs(5175)) xor (layer4_outputs(7502));
    layer5_outputs(1403) <= (layer4_outputs(3349)) and not (layer4_outputs(1029));
    layer5_outputs(1404) <= (layer4_outputs(3802)) xor (layer4_outputs(5423));
    layer5_outputs(1405) <= (layer4_outputs(6739)) and (layer4_outputs(7460));
    layer5_outputs(1406) <= not(layer4_outputs(5166));
    layer5_outputs(1407) <= layer4_outputs(5242);
    layer5_outputs(1408) <= not(layer4_outputs(2332));
    layer5_outputs(1409) <= not(layer4_outputs(1541));
    layer5_outputs(1410) <= not(layer4_outputs(6298));
    layer5_outputs(1411) <= '1';
    layer5_outputs(1412) <= not(layer4_outputs(6297));
    layer5_outputs(1413) <= '1';
    layer5_outputs(1414) <= layer4_outputs(3340);
    layer5_outputs(1415) <= not(layer4_outputs(677));
    layer5_outputs(1416) <= layer4_outputs(496);
    layer5_outputs(1417) <= layer4_outputs(1230);
    layer5_outputs(1418) <= (layer4_outputs(2472)) xor (layer4_outputs(1738));
    layer5_outputs(1419) <= layer4_outputs(7489);
    layer5_outputs(1420) <= not(layer4_outputs(2222)) or (layer4_outputs(6720));
    layer5_outputs(1421) <= not((layer4_outputs(1693)) xor (layer4_outputs(2053)));
    layer5_outputs(1422) <= (layer4_outputs(3930)) and not (layer4_outputs(1076));
    layer5_outputs(1423) <= (layer4_outputs(2696)) and not (layer4_outputs(6303));
    layer5_outputs(1424) <= layer4_outputs(862);
    layer5_outputs(1425) <= layer4_outputs(6062);
    layer5_outputs(1426) <= not((layer4_outputs(4947)) and (layer4_outputs(3013)));
    layer5_outputs(1427) <= not(layer4_outputs(5750));
    layer5_outputs(1428) <= not(layer4_outputs(5391));
    layer5_outputs(1429) <= not(layer4_outputs(150));
    layer5_outputs(1430) <= not(layer4_outputs(3954));
    layer5_outputs(1431) <= (layer4_outputs(4797)) or (layer4_outputs(3106));
    layer5_outputs(1432) <= '0';
    layer5_outputs(1433) <= (layer4_outputs(6424)) and not (layer4_outputs(4240));
    layer5_outputs(1434) <= not(layer4_outputs(1302)) or (layer4_outputs(6093));
    layer5_outputs(1435) <= (layer4_outputs(3233)) xor (layer4_outputs(5304));
    layer5_outputs(1436) <= layer4_outputs(1468);
    layer5_outputs(1437) <= (layer4_outputs(6133)) and not (layer4_outputs(7587));
    layer5_outputs(1438) <= layer4_outputs(2521);
    layer5_outputs(1439) <= not(layer4_outputs(5484));
    layer5_outputs(1440) <= (layer4_outputs(115)) and not (layer4_outputs(5304));
    layer5_outputs(1441) <= not(layer4_outputs(1226)) or (layer4_outputs(2324));
    layer5_outputs(1442) <= not(layer4_outputs(4441)) or (layer4_outputs(6707));
    layer5_outputs(1443) <= layer4_outputs(6410);
    layer5_outputs(1444) <= layer4_outputs(2095);
    layer5_outputs(1445) <= not((layer4_outputs(2081)) or (layer4_outputs(1919)));
    layer5_outputs(1446) <= layer4_outputs(5014);
    layer5_outputs(1447) <= '1';
    layer5_outputs(1448) <= not((layer4_outputs(3993)) xor (layer4_outputs(2712)));
    layer5_outputs(1449) <= (layer4_outputs(5878)) and not (layer4_outputs(6135));
    layer5_outputs(1450) <= not(layer4_outputs(52));
    layer5_outputs(1451) <= not(layer4_outputs(934));
    layer5_outputs(1452) <= not(layer4_outputs(2776));
    layer5_outputs(1453) <= (layer4_outputs(7063)) and not (layer4_outputs(3934));
    layer5_outputs(1454) <= not(layer4_outputs(1129)) or (layer4_outputs(7664));
    layer5_outputs(1455) <= (layer4_outputs(1466)) and not (layer4_outputs(2568));
    layer5_outputs(1456) <= layer4_outputs(1493);
    layer5_outputs(1457) <= (layer4_outputs(877)) and (layer4_outputs(2110));
    layer5_outputs(1458) <= not(layer4_outputs(4715)) or (layer4_outputs(5936));
    layer5_outputs(1459) <= (layer4_outputs(1339)) or (layer4_outputs(5710));
    layer5_outputs(1460) <= (layer4_outputs(2910)) xor (layer4_outputs(3448));
    layer5_outputs(1461) <= not((layer4_outputs(6868)) and (layer4_outputs(5653)));
    layer5_outputs(1462) <= not(layer4_outputs(1924));
    layer5_outputs(1463) <= '0';
    layer5_outputs(1464) <= '1';
    layer5_outputs(1465) <= (layer4_outputs(4297)) and not (layer4_outputs(5591));
    layer5_outputs(1466) <= not(layer4_outputs(3187)) or (layer4_outputs(243));
    layer5_outputs(1467) <= not((layer4_outputs(5349)) and (layer4_outputs(4679)));
    layer5_outputs(1468) <= '1';
    layer5_outputs(1469) <= layer4_outputs(6682);
    layer5_outputs(1470) <= not(layer4_outputs(6599)) or (layer4_outputs(1621));
    layer5_outputs(1471) <= not(layer4_outputs(1751));
    layer5_outputs(1472) <= layer4_outputs(5066);
    layer5_outputs(1473) <= not((layer4_outputs(2622)) xor (layer4_outputs(443)));
    layer5_outputs(1474) <= layer4_outputs(5498);
    layer5_outputs(1475) <= (layer4_outputs(4330)) xor (layer4_outputs(3594));
    layer5_outputs(1476) <= (layer4_outputs(7600)) and (layer4_outputs(2669));
    layer5_outputs(1477) <= (layer4_outputs(7645)) and not (layer4_outputs(5532));
    layer5_outputs(1478) <= layer4_outputs(2198);
    layer5_outputs(1479) <= (layer4_outputs(5643)) xor (layer4_outputs(7677));
    layer5_outputs(1480) <= not((layer4_outputs(2739)) and (layer4_outputs(4295)));
    layer5_outputs(1481) <= not(layer4_outputs(7376));
    layer5_outputs(1482) <= not(layer4_outputs(5671));
    layer5_outputs(1483) <= layer4_outputs(4901);
    layer5_outputs(1484) <= not((layer4_outputs(2748)) xor (layer4_outputs(4448)));
    layer5_outputs(1485) <= not(layer4_outputs(3032));
    layer5_outputs(1486) <= not(layer4_outputs(6771));
    layer5_outputs(1487) <= not(layer4_outputs(4434));
    layer5_outputs(1488) <= layer4_outputs(1264);
    layer5_outputs(1489) <= not(layer4_outputs(2508)) or (layer4_outputs(1721));
    layer5_outputs(1490) <= layer4_outputs(3868);
    layer5_outputs(1491) <= not(layer4_outputs(4149));
    layer5_outputs(1492) <= not((layer4_outputs(5508)) xor (layer4_outputs(6724)));
    layer5_outputs(1493) <= layer4_outputs(5724);
    layer5_outputs(1494) <= layer4_outputs(590);
    layer5_outputs(1495) <= (layer4_outputs(265)) and (layer4_outputs(182));
    layer5_outputs(1496) <= not(layer4_outputs(3054));
    layer5_outputs(1497) <= not(layer4_outputs(3810));
    layer5_outputs(1498) <= layer4_outputs(4984);
    layer5_outputs(1499) <= not(layer4_outputs(2703));
    layer5_outputs(1500) <= layer4_outputs(7373);
    layer5_outputs(1501) <= not(layer4_outputs(1111)) or (layer4_outputs(4375));
    layer5_outputs(1502) <= layer4_outputs(5212);
    layer5_outputs(1503) <= (layer4_outputs(4529)) and not (layer4_outputs(2568));
    layer5_outputs(1504) <= not(layer4_outputs(7062));
    layer5_outputs(1505) <= not(layer4_outputs(4936));
    layer5_outputs(1506) <= (layer4_outputs(4447)) xor (layer4_outputs(310));
    layer5_outputs(1507) <= layer4_outputs(2540);
    layer5_outputs(1508) <= layer4_outputs(2937);
    layer5_outputs(1509) <= not(layer4_outputs(1930));
    layer5_outputs(1510) <= layer4_outputs(973);
    layer5_outputs(1511) <= layer4_outputs(1690);
    layer5_outputs(1512) <= not(layer4_outputs(3363));
    layer5_outputs(1513) <= not((layer4_outputs(6430)) xor (layer4_outputs(369)));
    layer5_outputs(1514) <= layer4_outputs(3469);
    layer5_outputs(1515) <= (layer4_outputs(3572)) and not (layer4_outputs(6813));
    layer5_outputs(1516) <= (layer4_outputs(7328)) xor (layer4_outputs(6094));
    layer5_outputs(1517) <= not(layer4_outputs(2386)) or (layer4_outputs(2985));
    layer5_outputs(1518) <= (layer4_outputs(5079)) and not (layer4_outputs(116));
    layer5_outputs(1519) <= not(layer4_outputs(3075));
    layer5_outputs(1520) <= (layer4_outputs(5436)) and (layer4_outputs(5821));
    layer5_outputs(1521) <= not(layer4_outputs(398));
    layer5_outputs(1522) <= (layer4_outputs(7041)) and not (layer4_outputs(6882));
    layer5_outputs(1523) <= not(layer4_outputs(1618));
    layer5_outputs(1524) <= (layer4_outputs(7552)) and not (layer4_outputs(5835));
    layer5_outputs(1525) <= (layer4_outputs(991)) and not (layer4_outputs(559));
    layer5_outputs(1526) <= not((layer4_outputs(5363)) and (layer4_outputs(572)));
    layer5_outputs(1527) <= layer4_outputs(5769);
    layer5_outputs(1528) <= layer4_outputs(4822);
    layer5_outputs(1529) <= not(layer4_outputs(5107)) or (layer4_outputs(7017));
    layer5_outputs(1530) <= not(layer4_outputs(2790));
    layer5_outputs(1531) <= layer4_outputs(6652);
    layer5_outputs(1532) <= (layer4_outputs(6719)) and (layer4_outputs(7666));
    layer5_outputs(1533) <= layer4_outputs(6776);
    layer5_outputs(1534) <= not(layer4_outputs(827)) or (layer4_outputs(5165));
    layer5_outputs(1535) <= not(layer4_outputs(436));
    layer5_outputs(1536) <= (layer4_outputs(4765)) and not (layer4_outputs(913));
    layer5_outputs(1537) <= not(layer4_outputs(215));
    layer5_outputs(1538) <= not((layer4_outputs(1937)) or (layer4_outputs(4757)));
    layer5_outputs(1539) <= (layer4_outputs(3342)) and not (layer4_outputs(5123));
    layer5_outputs(1540) <= not(layer4_outputs(3331));
    layer5_outputs(1541) <= (layer4_outputs(6099)) and not (layer4_outputs(4383));
    layer5_outputs(1542) <= '1';
    layer5_outputs(1543) <= not((layer4_outputs(6680)) and (layer4_outputs(3078)));
    layer5_outputs(1544) <= not(layer4_outputs(3862));
    layer5_outputs(1545) <= not((layer4_outputs(7520)) xor (layer4_outputs(6429)));
    layer5_outputs(1546) <= not(layer4_outputs(1619)) or (layer4_outputs(2010));
    layer5_outputs(1547) <= (layer4_outputs(6413)) and (layer4_outputs(4237));
    layer5_outputs(1548) <= not(layer4_outputs(3966)) or (layer4_outputs(5938));
    layer5_outputs(1549) <= not((layer4_outputs(638)) xor (layer4_outputs(3505)));
    layer5_outputs(1550) <= '0';
    layer5_outputs(1551) <= not(layer4_outputs(1070));
    layer5_outputs(1552) <= (layer4_outputs(1903)) and not (layer4_outputs(1646));
    layer5_outputs(1553) <= (layer4_outputs(3302)) xor (layer4_outputs(6832));
    layer5_outputs(1554) <= not(layer4_outputs(5703));
    layer5_outputs(1555) <= not(layer4_outputs(4110)) or (layer4_outputs(5050));
    layer5_outputs(1556) <= not(layer4_outputs(4392)) or (layer4_outputs(4115));
    layer5_outputs(1557) <= not((layer4_outputs(4463)) and (layer4_outputs(6549)));
    layer5_outputs(1558) <= (layer4_outputs(1949)) or (layer4_outputs(4104));
    layer5_outputs(1559) <= not(layer4_outputs(536));
    layer5_outputs(1560) <= layer4_outputs(1664);
    layer5_outputs(1561) <= (layer4_outputs(725)) and not (layer4_outputs(7407));
    layer5_outputs(1562) <= not(layer4_outputs(2791));
    layer5_outputs(1563) <= (layer4_outputs(2606)) and (layer4_outputs(1729));
    layer5_outputs(1564) <= (layer4_outputs(6267)) xor (layer4_outputs(672));
    layer5_outputs(1565) <= not(layer4_outputs(3778));
    layer5_outputs(1566) <= layer4_outputs(2498);
    layer5_outputs(1567) <= not((layer4_outputs(4868)) xor (layer4_outputs(5433)));
    layer5_outputs(1568) <= (layer4_outputs(5447)) xor (layer4_outputs(119));
    layer5_outputs(1569) <= '0';
    layer5_outputs(1570) <= not(layer4_outputs(895));
    layer5_outputs(1571) <= not(layer4_outputs(3259));
    layer5_outputs(1572) <= (layer4_outputs(5849)) and not (layer4_outputs(65));
    layer5_outputs(1573) <= layer4_outputs(6762);
    layer5_outputs(1574) <= (layer4_outputs(123)) and not (layer4_outputs(3442));
    layer5_outputs(1575) <= not((layer4_outputs(3907)) and (layer4_outputs(2651)));
    layer5_outputs(1576) <= layer4_outputs(4179);
    layer5_outputs(1577) <= layer4_outputs(6485);
    layer5_outputs(1578) <= (layer4_outputs(2017)) and not (layer4_outputs(1569));
    layer5_outputs(1579) <= not(layer4_outputs(2834));
    layer5_outputs(1580) <= not(layer4_outputs(2469));
    layer5_outputs(1581) <= not(layer4_outputs(2770));
    layer5_outputs(1582) <= not((layer4_outputs(5630)) xor (layer4_outputs(3533)));
    layer5_outputs(1583) <= layer4_outputs(745);
    layer5_outputs(1584) <= '0';
    layer5_outputs(1585) <= not(layer4_outputs(7560));
    layer5_outputs(1586) <= not(layer4_outputs(6257));
    layer5_outputs(1587) <= not(layer4_outputs(7444));
    layer5_outputs(1588) <= (layer4_outputs(6552)) and not (layer4_outputs(2723));
    layer5_outputs(1589) <= layer4_outputs(3726);
    layer5_outputs(1590) <= not(layer4_outputs(4012));
    layer5_outputs(1591) <= layer4_outputs(3336);
    layer5_outputs(1592) <= not(layer4_outputs(3519));
    layer5_outputs(1593) <= not(layer4_outputs(6460));
    layer5_outputs(1594) <= not(layer4_outputs(3509));
    layer5_outputs(1595) <= layer4_outputs(2550);
    layer5_outputs(1596) <= not(layer4_outputs(6956));
    layer5_outputs(1597) <= not(layer4_outputs(7537)) or (layer4_outputs(619));
    layer5_outputs(1598) <= (layer4_outputs(7361)) and not (layer4_outputs(5483));
    layer5_outputs(1599) <= not(layer4_outputs(3214));
    layer5_outputs(1600) <= not(layer4_outputs(1169));
    layer5_outputs(1601) <= not(layer4_outputs(4653)) or (layer4_outputs(2367));
    layer5_outputs(1602) <= layer4_outputs(6993);
    layer5_outputs(1603) <= not(layer4_outputs(4875));
    layer5_outputs(1604) <= not(layer4_outputs(6968));
    layer5_outputs(1605) <= layer4_outputs(2365);
    layer5_outputs(1606) <= layer4_outputs(2687);
    layer5_outputs(1607) <= layer4_outputs(1838);
    layer5_outputs(1608) <= not(layer4_outputs(1194));
    layer5_outputs(1609) <= layer4_outputs(5309);
    layer5_outputs(1610) <= not((layer4_outputs(2592)) or (layer4_outputs(7529)));
    layer5_outputs(1611) <= layer4_outputs(1989);
    layer5_outputs(1612) <= layer4_outputs(1439);
    layer5_outputs(1613) <= layer4_outputs(2526);
    layer5_outputs(1614) <= not(layer4_outputs(5815)) or (layer4_outputs(6901));
    layer5_outputs(1615) <= layer4_outputs(4656);
    layer5_outputs(1616) <= (layer4_outputs(2016)) and not (layer4_outputs(5189));
    layer5_outputs(1617) <= not(layer4_outputs(252));
    layer5_outputs(1618) <= layer4_outputs(6800);
    layer5_outputs(1619) <= not(layer4_outputs(6798)) or (layer4_outputs(1685));
    layer5_outputs(1620) <= '1';
    layer5_outputs(1621) <= not(layer4_outputs(3930)) or (layer4_outputs(2090));
    layer5_outputs(1622) <= layer4_outputs(3206);
    layer5_outputs(1623) <= layer4_outputs(682);
    layer5_outputs(1624) <= layer4_outputs(748);
    layer5_outputs(1625) <= (layer4_outputs(3239)) and not (layer4_outputs(4798));
    layer5_outputs(1626) <= '1';
    layer5_outputs(1627) <= layer4_outputs(2556);
    layer5_outputs(1628) <= layer4_outputs(769);
    layer5_outputs(1629) <= not(layer4_outputs(4310));
    layer5_outputs(1630) <= not(layer4_outputs(2859)) or (layer4_outputs(3531));
    layer5_outputs(1631) <= (layer4_outputs(2096)) and not (layer4_outputs(5007));
    layer5_outputs(1632) <= not(layer4_outputs(5781));
    layer5_outputs(1633) <= layer4_outputs(987);
    layer5_outputs(1634) <= not(layer4_outputs(2120)) or (layer4_outputs(2485));
    layer5_outputs(1635) <= layer4_outputs(4262);
    layer5_outputs(1636) <= layer4_outputs(1);
    layer5_outputs(1637) <= layer4_outputs(320);
    layer5_outputs(1638) <= '0';
    layer5_outputs(1639) <= not((layer4_outputs(647)) and (layer4_outputs(355)));
    layer5_outputs(1640) <= layer4_outputs(1692);
    layer5_outputs(1641) <= (layer4_outputs(486)) xor (layer4_outputs(6322));
    layer5_outputs(1642) <= not((layer4_outputs(449)) xor (layer4_outputs(2760)));
    layer5_outputs(1643) <= layer4_outputs(6773);
    layer5_outputs(1644) <= layer4_outputs(1581);
    layer5_outputs(1645) <= layer4_outputs(6887);
    layer5_outputs(1646) <= layer4_outputs(7649);
    layer5_outputs(1647) <= (layer4_outputs(6519)) and not (layer4_outputs(767));
    layer5_outputs(1648) <= layer4_outputs(4690);
    layer5_outputs(1649) <= layer4_outputs(5968);
    layer5_outputs(1650) <= layer4_outputs(1707);
    layer5_outputs(1651) <= layer4_outputs(4746);
    layer5_outputs(1652) <= not(layer4_outputs(939));
    layer5_outputs(1653) <= not(layer4_outputs(524)) or (layer4_outputs(6243));
    layer5_outputs(1654) <= '0';
    layer5_outputs(1655) <= (layer4_outputs(528)) and not (layer4_outputs(522));
    layer5_outputs(1656) <= layer4_outputs(3519);
    layer5_outputs(1657) <= layer4_outputs(6146);
    layer5_outputs(1658) <= (layer4_outputs(7174)) and not (layer4_outputs(5572));
    layer5_outputs(1659) <= not((layer4_outputs(3687)) xor (layer4_outputs(5539)));
    layer5_outputs(1660) <= not(layer4_outputs(5173)) or (layer4_outputs(5830));
    layer5_outputs(1661) <= not((layer4_outputs(5278)) or (layer4_outputs(5791)));
    layer5_outputs(1662) <= not(layer4_outputs(6005));
    layer5_outputs(1663) <= not((layer4_outputs(4339)) and (layer4_outputs(7059)));
    layer5_outputs(1664) <= (layer4_outputs(1916)) or (layer4_outputs(2919));
    layer5_outputs(1665) <= not(layer4_outputs(5445));
    layer5_outputs(1666) <= not(layer4_outputs(1276)) or (layer4_outputs(109));
    layer5_outputs(1667) <= not((layer4_outputs(912)) or (layer4_outputs(7675)));
    layer5_outputs(1668) <= (layer4_outputs(3270)) and not (layer4_outputs(1611));
    layer5_outputs(1669) <= (layer4_outputs(6584)) and not (layer4_outputs(194));
    layer5_outputs(1670) <= not(layer4_outputs(7142));
    layer5_outputs(1671) <= not(layer4_outputs(6737));
    layer5_outputs(1672) <= not((layer4_outputs(6509)) or (layer4_outputs(2409)));
    layer5_outputs(1673) <= (layer4_outputs(5648)) and not (layer4_outputs(3877));
    layer5_outputs(1674) <= (layer4_outputs(7406)) and not (layer4_outputs(3602));
    layer5_outputs(1675) <= layer4_outputs(1682);
    layer5_outputs(1676) <= (layer4_outputs(5695)) and not (layer4_outputs(6872));
    layer5_outputs(1677) <= layer4_outputs(3558);
    layer5_outputs(1678) <= not(layer4_outputs(441)) or (layer4_outputs(3294));
    layer5_outputs(1679) <= not(layer4_outputs(667)) or (layer4_outputs(6505));
    layer5_outputs(1680) <= '1';
    layer5_outputs(1681) <= not(layer4_outputs(3372));
    layer5_outputs(1682) <= '1';
    layer5_outputs(1683) <= not(layer4_outputs(1534)) or (layer4_outputs(4683));
    layer5_outputs(1684) <= not(layer4_outputs(480));
    layer5_outputs(1685) <= not((layer4_outputs(301)) and (layer4_outputs(5599)));
    layer5_outputs(1686) <= not((layer4_outputs(930)) and (layer4_outputs(1168)));
    layer5_outputs(1687) <= (layer4_outputs(2341)) and not (layer4_outputs(3725));
    layer5_outputs(1688) <= layer4_outputs(7005);
    layer5_outputs(1689) <= layer4_outputs(4121);
    layer5_outputs(1690) <= not(layer4_outputs(2274));
    layer5_outputs(1691) <= not(layer4_outputs(4713));
    layer5_outputs(1692) <= not(layer4_outputs(7208));
    layer5_outputs(1693) <= layer4_outputs(1190);
    layer5_outputs(1694) <= not(layer4_outputs(5323));
    layer5_outputs(1695) <= '1';
    layer5_outputs(1696) <= (layer4_outputs(494)) and (layer4_outputs(711));
    layer5_outputs(1697) <= (layer4_outputs(2271)) xor (layer4_outputs(2686));
    layer5_outputs(1698) <= not((layer4_outputs(3262)) or (layer4_outputs(4114)));
    layer5_outputs(1699) <= layer4_outputs(6926);
    layer5_outputs(1700) <= not((layer4_outputs(5930)) xor (layer4_outputs(3121)));
    layer5_outputs(1701) <= (layer4_outputs(6315)) and not (layer4_outputs(7014));
    layer5_outputs(1702) <= layer4_outputs(6275);
    layer5_outputs(1703) <= (layer4_outputs(6795)) xor (layer4_outputs(2717));
    layer5_outputs(1704) <= not((layer4_outputs(7451)) xor (layer4_outputs(7558)));
    layer5_outputs(1705) <= (layer4_outputs(3917)) xor (layer4_outputs(2041));
    layer5_outputs(1706) <= (layer4_outputs(3741)) and not (layer4_outputs(848));
    layer5_outputs(1707) <= not((layer4_outputs(4570)) xor (layer4_outputs(4859)));
    layer5_outputs(1708) <= (layer4_outputs(1814)) xor (layer4_outputs(930));
    layer5_outputs(1709) <= not(layer4_outputs(5200)) or (layer4_outputs(1071));
    layer5_outputs(1710) <= layer4_outputs(1333);
    layer5_outputs(1711) <= layer4_outputs(3065);
    layer5_outputs(1712) <= not((layer4_outputs(1273)) or (layer4_outputs(2845)));
    layer5_outputs(1713) <= layer4_outputs(3701);
    layer5_outputs(1714) <= not(layer4_outputs(2116));
    layer5_outputs(1715) <= (layer4_outputs(1628)) and not (layer4_outputs(7655));
    layer5_outputs(1716) <= (layer4_outputs(3999)) and not (layer4_outputs(5444));
    layer5_outputs(1717) <= not((layer4_outputs(7220)) and (layer4_outputs(6154)));
    layer5_outputs(1718) <= (layer4_outputs(4916)) or (layer4_outputs(656));
    layer5_outputs(1719) <= layer4_outputs(1382);
    layer5_outputs(1720) <= (layer4_outputs(23)) or (layer4_outputs(3698));
    layer5_outputs(1721) <= (layer4_outputs(5585)) and (layer4_outputs(6922));
    layer5_outputs(1722) <= layer4_outputs(4751);
    layer5_outputs(1723) <= layer4_outputs(3875);
    layer5_outputs(1724) <= not(layer4_outputs(653));
    layer5_outputs(1725) <= layer4_outputs(3974);
    layer5_outputs(1726) <= layer4_outputs(3278);
    layer5_outputs(1727) <= not((layer4_outputs(1157)) or (layer4_outputs(4439)));
    layer5_outputs(1728) <= (layer4_outputs(1535)) and not (layer4_outputs(755));
    layer5_outputs(1729) <= layer4_outputs(3648);
    layer5_outputs(1730) <= not(layer4_outputs(3277));
    layer5_outputs(1731) <= not(layer4_outputs(5473));
    layer5_outputs(1732) <= not(layer4_outputs(3313));
    layer5_outputs(1733) <= not(layer4_outputs(422));
    layer5_outputs(1734) <= (layer4_outputs(375)) or (layer4_outputs(4875));
    layer5_outputs(1735) <= (layer4_outputs(4700)) and not (layer4_outputs(7131));
    layer5_outputs(1736) <= layer4_outputs(1752);
    layer5_outputs(1737) <= (layer4_outputs(6363)) and not (layer4_outputs(1890));
    layer5_outputs(1738) <= not(layer4_outputs(1862));
    layer5_outputs(1739) <= layer4_outputs(6391);
    layer5_outputs(1740) <= layer4_outputs(3508);
    layer5_outputs(1741) <= not(layer4_outputs(7436));
    layer5_outputs(1742) <= (layer4_outputs(2133)) and not (layer4_outputs(4897));
    layer5_outputs(1743) <= (layer4_outputs(7581)) or (layer4_outputs(195));
    layer5_outputs(1744) <= '0';
    layer5_outputs(1745) <= not(layer4_outputs(2880));
    layer5_outputs(1746) <= not(layer4_outputs(4855));
    layer5_outputs(1747) <= not((layer4_outputs(7538)) or (layer4_outputs(2697)));
    layer5_outputs(1748) <= not(layer4_outputs(3526)) or (layer4_outputs(6196));
    layer5_outputs(1749) <= not(layer4_outputs(3242)) or (layer4_outputs(7049));
    layer5_outputs(1750) <= layer4_outputs(6448);
    layer5_outputs(1751) <= (layer4_outputs(5036)) and not (layer4_outputs(3274));
    layer5_outputs(1752) <= (layer4_outputs(3960)) and not (layer4_outputs(1362));
    layer5_outputs(1753) <= not(layer4_outputs(7647));
    layer5_outputs(1754) <= '0';
    layer5_outputs(1755) <= layer4_outputs(4131);
    layer5_outputs(1756) <= (layer4_outputs(3172)) and not (layer4_outputs(1760));
    layer5_outputs(1757) <= layer4_outputs(70);
    layer5_outputs(1758) <= layer4_outputs(5935);
    layer5_outputs(1759) <= not(layer4_outputs(3321));
    layer5_outputs(1760) <= (layer4_outputs(7452)) xor (layer4_outputs(2005));
    layer5_outputs(1761) <= (layer4_outputs(2618)) xor (layer4_outputs(4264));
    layer5_outputs(1762) <= not(layer4_outputs(3757));
    layer5_outputs(1763) <= layer4_outputs(1801);
    layer5_outputs(1764) <= layer4_outputs(4391);
    layer5_outputs(1765) <= not(layer4_outputs(3280));
    layer5_outputs(1766) <= layer4_outputs(7336);
    layer5_outputs(1767) <= not(layer4_outputs(4891)) or (layer4_outputs(1665));
    layer5_outputs(1768) <= layer4_outputs(7104);
    layer5_outputs(1769) <= not(layer4_outputs(3066));
    layer5_outputs(1770) <= '1';
    layer5_outputs(1771) <= (layer4_outputs(4595)) or (layer4_outputs(7674));
    layer5_outputs(1772) <= not(layer4_outputs(2326)) or (layer4_outputs(909));
    layer5_outputs(1773) <= (layer4_outputs(986)) and not (layer4_outputs(4303));
    layer5_outputs(1774) <= not(layer4_outputs(2384)) or (layer4_outputs(1421));
    layer5_outputs(1775) <= (layer4_outputs(1377)) and not (layer4_outputs(5832));
    layer5_outputs(1776) <= (layer4_outputs(3592)) or (layer4_outputs(5999));
    layer5_outputs(1777) <= not((layer4_outputs(5296)) and (layer4_outputs(76)));
    layer5_outputs(1778) <= not(layer4_outputs(7312)) or (layer4_outputs(6859));
    layer5_outputs(1779) <= layer4_outputs(6603);
    layer5_outputs(1780) <= not(layer4_outputs(6790));
    layer5_outputs(1781) <= not(layer4_outputs(5426));
    layer5_outputs(1782) <= layer4_outputs(4685);
    layer5_outputs(1783) <= not(layer4_outputs(7067));
    layer5_outputs(1784) <= layer4_outputs(402);
    layer5_outputs(1785) <= (layer4_outputs(6717)) and not (layer4_outputs(294));
    layer5_outputs(1786) <= not((layer4_outputs(6057)) and (layer4_outputs(2345)));
    layer5_outputs(1787) <= not((layer4_outputs(2193)) xor (layer4_outputs(6332)));
    layer5_outputs(1788) <= not(layer4_outputs(4414));
    layer5_outputs(1789) <= layer4_outputs(1348);
    layer5_outputs(1790) <= layer4_outputs(6875);
    layer5_outputs(1791) <= not(layer4_outputs(3324));
    layer5_outputs(1792) <= not((layer4_outputs(4478)) xor (layer4_outputs(607)));
    layer5_outputs(1793) <= (layer4_outputs(6238)) xor (layer4_outputs(4177));
    layer5_outputs(1794) <= not((layer4_outputs(3484)) and (layer4_outputs(2055)));
    layer5_outputs(1795) <= not((layer4_outputs(7032)) xor (layer4_outputs(1677)));
    layer5_outputs(1796) <= not(layer4_outputs(5457)) or (layer4_outputs(7554));
    layer5_outputs(1797) <= not(layer4_outputs(1947));
    layer5_outputs(1798) <= layer4_outputs(3089);
    layer5_outputs(1799) <= layer4_outputs(2822);
    layer5_outputs(1800) <= (layer4_outputs(4)) and (layer4_outputs(7479));
    layer5_outputs(1801) <= not((layer4_outputs(2079)) and (layer4_outputs(6504)));
    layer5_outputs(1802) <= not(layer4_outputs(6054));
    layer5_outputs(1803) <= not(layer4_outputs(7653)) or (layer4_outputs(1105));
    layer5_outputs(1804) <= not(layer4_outputs(4605)) or (layer4_outputs(4803));
    layer5_outputs(1805) <= not(layer4_outputs(426));
    layer5_outputs(1806) <= not((layer4_outputs(1313)) xor (layer4_outputs(1161)));
    layer5_outputs(1807) <= not(layer4_outputs(4470));
    layer5_outputs(1808) <= '0';
    layer5_outputs(1809) <= not(layer4_outputs(5183));
    layer5_outputs(1810) <= layer4_outputs(6160);
    layer5_outputs(1811) <= not(layer4_outputs(2742));
    layer5_outputs(1812) <= not(layer4_outputs(4275)) or (layer4_outputs(3151));
    layer5_outputs(1813) <= '1';
    layer5_outputs(1814) <= (layer4_outputs(4215)) or (layer4_outputs(6261));
    layer5_outputs(1815) <= layer4_outputs(7641);
    layer5_outputs(1816) <= (layer4_outputs(140)) and (layer4_outputs(6368));
    layer5_outputs(1817) <= layer4_outputs(301);
    layer5_outputs(1818) <= not((layer4_outputs(5373)) xor (layer4_outputs(4300)));
    layer5_outputs(1819) <= (layer4_outputs(1626)) and not (layer4_outputs(1520));
    layer5_outputs(1820) <= layer4_outputs(4543);
    layer5_outputs(1821) <= not(layer4_outputs(1718)) or (layer4_outputs(2837));
    layer5_outputs(1822) <= (layer4_outputs(3081)) and not (layer4_outputs(7609));
    layer5_outputs(1823) <= layer4_outputs(1521);
    layer5_outputs(1824) <= (layer4_outputs(6814)) xor (layer4_outputs(4545));
    layer5_outputs(1825) <= '0';
    layer5_outputs(1826) <= not(layer4_outputs(6975));
    layer5_outputs(1827) <= not((layer4_outputs(465)) or (layer4_outputs(3514)));
    layer5_outputs(1828) <= layer4_outputs(1794);
    layer5_outputs(1829) <= layer4_outputs(1816);
    layer5_outputs(1830) <= not(layer4_outputs(5085));
    layer5_outputs(1831) <= (layer4_outputs(749)) or (layer4_outputs(3229));
    layer5_outputs(1832) <= layer4_outputs(2528);
    layer5_outputs(1833) <= (layer4_outputs(3992)) or (layer4_outputs(2415));
    layer5_outputs(1834) <= (layer4_outputs(7135)) xor (layer4_outputs(3825));
    layer5_outputs(1835) <= not(layer4_outputs(2440));
    layer5_outputs(1836) <= (layer4_outputs(7606)) or (layer4_outputs(799));
    layer5_outputs(1837) <= (layer4_outputs(6539)) or (layer4_outputs(1717));
    layer5_outputs(1838) <= '0';
    layer5_outputs(1839) <= layer4_outputs(5523);
    layer5_outputs(1840) <= not((layer4_outputs(6378)) and (layer4_outputs(4563)));
    layer5_outputs(1841) <= not(layer4_outputs(965)) or (layer4_outputs(1638));
    layer5_outputs(1842) <= not(layer4_outputs(3127));
    layer5_outputs(1843) <= (layer4_outputs(6819)) or (layer4_outputs(875));
    layer5_outputs(1844) <= not((layer4_outputs(2139)) xor (layer4_outputs(2930)));
    layer5_outputs(1845) <= '0';
    layer5_outputs(1846) <= not(layer4_outputs(6919)) or (layer4_outputs(3913));
    layer5_outputs(1847) <= (layer4_outputs(5491)) or (layer4_outputs(2661));
    layer5_outputs(1848) <= layer4_outputs(4112);
    layer5_outputs(1849) <= not(layer4_outputs(6122));
    layer5_outputs(1850) <= not(layer4_outputs(6726)) or (layer4_outputs(2653));
    layer5_outputs(1851) <= layer4_outputs(4514);
    layer5_outputs(1852) <= (layer4_outputs(4777)) xor (layer4_outputs(2581));
    layer5_outputs(1853) <= (layer4_outputs(576)) and not (layer4_outputs(5042));
    layer5_outputs(1854) <= layer4_outputs(6627);
    layer5_outputs(1855) <= layer4_outputs(1963);
    layer5_outputs(1856) <= not(layer4_outputs(2510)) or (layer4_outputs(6306));
    layer5_outputs(1857) <= not((layer4_outputs(170)) xor (layer4_outputs(1868)));
    layer5_outputs(1858) <= not(layer4_outputs(7181)) or (layer4_outputs(4732));
    layer5_outputs(1859) <= not(layer4_outputs(7663));
    layer5_outputs(1860) <= '0';
    layer5_outputs(1861) <= (layer4_outputs(3320)) xor (layer4_outputs(6860));
    layer5_outputs(1862) <= not(layer4_outputs(1927));
    layer5_outputs(1863) <= not(layer4_outputs(2891)) or (layer4_outputs(1204));
    layer5_outputs(1864) <= layer4_outputs(5400);
    layer5_outputs(1865) <= (layer4_outputs(197)) and not (layer4_outputs(3397));
    layer5_outputs(1866) <= not((layer4_outputs(7052)) xor (layer4_outputs(7492)));
    layer5_outputs(1867) <= not(layer4_outputs(2943));
    layer5_outputs(1868) <= (layer4_outputs(2309)) xor (layer4_outputs(3191));
    layer5_outputs(1869) <= layer4_outputs(2014);
    layer5_outputs(1870) <= (layer4_outputs(2262)) and not (layer4_outputs(25));
    layer5_outputs(1871) <= layer4_outputs(6675);
    layer5_outputs(1872) <= layer4_outputs(7296);
    layer5_outputs(1873) <= (layer4_outputs(265)) xor (layer4_outputs(963));
    layer5_outputs(1874) <= not((layer4_outputs(4374)) and (layer4_outputs(2913)));
    layer5_outputs(1875) <= (layer4_outputs(5251)) and not (layer4_outputs(5998));
    layer5_outputs(1876) <= (layer4_outputs(6339)) or (layer4_outputs(6113));
    layer5_outputs(1877) <= not(layer4_outputs(1982)) or (layer4_outputs(4578));
    layer5_outputs(1878) <= not(layer4_outputs(2862));
    layer5_outputs(1879) <= not((layer4_outputs(6852)) xor (layer4_outputs(2259)));
    layer5_outputs(1880) <= layer4_outputs(2436);
    layer5_outputs(1881) <= not((layer4_outputs(4885)) xor (layer4_outputs(4947)));
    layer5_outputs(1882) <= (layer4_outputs(3820)) or (layer4_outputs(3604));
    layer5_outputs(1883) <= not(layer4_outputs(3162));
    layer5_outputs(1884) <= not(layer4_outputs(6310));
    layer5_outputs(1885) <= (layer4_outputs(2186)) xor (layer4_outputs(5225));
    layer5_outputs(1886) <= layer4_outputs(5254);
    layer5_outputs(1887) <= layer4_outputs(2458);
    layer5_outputs(1888) <= layer4_outputs(7530);
    layer5_outputs(1889) <= '1';
    layer5_outputs(1890) <= (layer4_outputs(6768)) xor (layer4_outputs(6249));
    layer5_outputs(1891) <= not(layer4_outputs(6799)) or (layer4_outputs(1392));
    layer5_outputs(1892) <= not(layer4_outputs(5006));
    layer5_outputs(1893) <= (layer4_outputs(7072)) and not (layer4_outputs(3503));
    layer5_outputs(1894) <= not((layer4_outputs(4559)) xor (layer4_outputs(2282)));
    layer5_outputs(1895) <= layer4_outputs(7401);
    layer5_outputs(1896) <= '0';
    layer5_outputs(1897) <= layer4_outputs(4436);
    layer5_outputs(1898) <= (layer4_outputs(2759)) xor (layer4_outputs(5218));
    layer5_outputs(1899) <= layer4_outputs(6451);
    layer5_outputs(1900) <= not((layer4_outputs(2901)) or (layer4_outputs(4145)));
    layer5_outputs(1901) <= (layer4_outputs(3215)) or (layer4_outputs(4332));
    layer5_outputs(1902) <= '0';
    layer5_outputs(1903) <= layer4_outputs(6582);
    layer5_outputs(1904) <= layer4_outputs(5289);
    layer5_outputs(1905) <= not((layer4_outputs(4995)) or (layer4_outputs(6283)));
    layer5_outputs(1906) <= not(layer4_outputs(4522));
    layer5_outputs(1907) <= layer4_outputs(4623);
    layer5_outputs(1908) <= not(layer4_outputs(1583));
    layer5_outputs(1909) <= not((layer4_outputs(5919)) xor (layer4_outputs(6591)));
    layer5_outputs(1910) <= not((layer4_outputs(7296)) or (layer4_outputs(3813)));
    layer5_outputs(1911) <= not(layer4_outputs(6842));
    layer5_outputs(1912) <= not(layer4_outputs(1469));
    layer5_outputs(1913) <= not((layer4_outputs(907)) or (layer4_outputs(141)));
    layer5_outputs(1914) <= not(layer4_outputs(5638)) or (layer4_outputs(3440));
    layer5_outputs(1915) <= layer4_outputs(5340);
    layer5_outputs(1916) <= layer4_outputs(6957);
    layer5_outputs(1917) <= not((layer4_outputs(4094)) or (layer4_outputs(5246)));
    layer5_outputs(1918) <= not(layer4_outputs(2021));
    layer5_outputs(1919) <= (layer4_outputs(1303)) xor (layer4_outputs(7227));
    layer5_outputs(1920) <= not(layer4_outputs(5621));
    layer5_outputs(1921) <= not((layer4_outputs(5198)) and (layer4_outputs(7668)));
    layer5_outputs(1922) <= (layer4_outputs(7603)) and (layer4_outputs(4202));
    layer5_outputs(1923) <= layer4_outputs(1491);
    layer5_outputs(1924) <= (layer4_outputs(5277)) or (layer4_outputs(2903));
    layer5_outputs(1925) <= '0';
    layer5_outputs(1926) <= layer4_outputs(2475);
    layer5_outputs(1927) <= not(layer4_outputs(989));
    layer5_outputs(1928) <= (layer4_outputs(4426)) xor (layer4_outputs(185));
    layer5_outputs(1929) <= not(layer4_outputs(1286)) or (layer4_outputs(1039));
    layer5_outputs(1930) <= not(layer4_outputs(5549));
    layer5_outputs(1931) <= layer4_outputs(5943);
    layer5_outputs(1932) <= layer4_outputs(5498);
    layer5_outputs(1933) <= (layer4_outputs(6597)) xor (layer4_outputs(4912));
    layer5_outputs(1934) <= not(layer4_outputs(4039));
    layer5_outputs(1935) <= layer4_outputs(4780);
    layer5_outputs(1936) <= not(layer4_outputs(4714)) or (layer4_outputs(161));
    layer5_outputs(1937) <= not((layer4_outputs(2333)) xor (layer4_outputs(2464)));
    layer5_outputs(1938) <= layer4_outputs(6740);
    layer5_outputs(1939) <= not(layer4_outputs(1195));
    layer5_outputs(1940) <= layer4_outputs(6253);
    layer5_outputs(1941) <= not((layer4_outputs(4921)) xor (layer4_outputs(3272)));
    layer5_outputs(1942) <= layer4_outputs(909);
    layer5_outputs(1943) <= layer4_outputs(6308);
    layer5_outputs(1944) <= not((layer4_outputs(3998)) or (layer4_outputs(1573)));
    layer5_outputs(1945) <= (layer4_outputs(4021)) and (layer4_outputs(5644));
    layer5_outputs(1946) <= not(layer4_outputs(7593)) or (layer4_outputs(5940));
    layer5_outputs(1947) <= (layer4_outputs(4223)) and not (layer4_outputs(688));
    layer5_outputs(1948) <= '1';
    layer5_outputs(1949) <= layer4_outputs(2561);
    layer5_outputs(1950) <= not(layer4_outputs(2779));
    layer5_outputs(1951) <= not(layer4_outputs(6070)) or (layer4_outputs(4024));
    layer5_outputs(1952) <= layer4_outputs(554);
    layer5_outputs(1953) <= (layer4_outputs(7353)) and not (layer4_outputs(7280));
    layer5_outputs(1954) <= not(layer4_outputs(3332));
    layer5_outputs(1955) <= not(layer4_outputs(810)) or (layer4_outputs(5009));
    layer5_outputs(1956) <= layer4_outputs(7340);
    layer5_outputs(1957) <= not(layer4_outputs(2195));
    layer5_outputs(1958) <= not(layer4_outputs(73));
    layer5_outputs(1959) <= not(layer4_outputs(6779)) or (layer4_outputs(4350));
    layer5_outputs(1960) <= layer4_outputs(4665);
    layer5_outputs(1961) <= not(layer4_outputs(3481));
    layer5_outputs(1962) <= (layer4_outputs(3624)) xor (layer4_outputs(2235));
    layer5_outputs(1963) <= not(layer4_outputs(5695)) or (layer4_outputs(3616));
    layer5_outputs(1964) <= not((layer4_outputs(3842)) and (layer4_outputs(3791)));
    layer5_outputs(1965) <= (layer4_outputs(1548)) xor (layer4_outputs(3388));
    layer5_outputs(1966) <= not(layer4_outputs(7078));
    layer5_outputs(1967) <= layer4_outputs(6627);
    layer5_outputs(1968) <= layer4_outputs(4340);
    layer5_outputs(1969) <= (layer4_outputs(4026)) and not (layer4_outputs(6523));
    layer5_outputs(1970) <= not(layer4_outputs(7142));
    layer5_outputs(1971) <= (layer4_outputs(2841)) and not (layer4_outputs(2682));
    layer5_outputs(1972) <= not(layer4_outputs(4307));
    layer5_outputs(1973) <= not((layer4_outputs(6529)) xor (layer4_outputs(1292)));
    layer5_outputs(1974) <= layer4_outputs(4807);
    layer5_outputs(1975) <= not(layer4_outputs(362));
    layer5_outputs(1976) <= (layer4_outputs(3719)) xor (layer4_outputs(6034));
    layer5_outputs(1977) <= not(layer4_outputs(6985)) or (layer4_outputs(4910));
    layer5_outputs(1978) <= (layer4_outputs(100)) and (layer4_outputs(5730));
    layer5_outputs(1979) <= (layer4_outputs(871)) and not (layer4_outputs(1661));
    layer5_outputs(1980) <= not(layer4_outputs(6729));
    layer5_outputs(1981) <= (layer4_outputs(7563)) and not (layer4_outputs(2092));
    layer5_outputs(1982) <= (layer4_outputs(249)) and not (layer4_outputs(3255));
    layer5_outputs(1983) <= layer4_outputs(3252);
    layer5_outputs(1984) <= layer4_outputs(1100);
    layer5_outputs(1985) <= not((layer4_outputs(5509)) and (layer4_outputs(3987)));
    layer5_outputs(1986) <= (layer4_outputs(1602)) xor (layer4_outputs(3764));
    layer5_outputs(1987) <= not(layer4_outputs(2841)) or (layer4_outputs(6304));
    layer5_outputs(1988) <= not(layer4_outputs(778));
    layer5_outputs(1989) <= (layer4_outputs(4650)) and (layer4_outputs(3310));
    layer5_outputs(1990) <= '1';
    layer5_outputs(1991) <= not(layer4_outputs(1336));
    layer5_outputs(1992) <= (layer4_outputs(4702)) and (layer4_outputs(7541));
    layer5_outputs(1993) <= not(layer4_outputs(51));
    layer5_outputs(1994) <= (layer4_outputs(5025)) and not (layer4_outputs(1976));
    layer5_outputs(1995) <= not((layer4_outputs(5324)) or (layer4_outputs(2404)));
    layer5_outputs(1996) <= not(layer4_outputs(1625));
    layer5_outputs(1997) <= not(layer4_outputs(6939));
    layer5_outputs(1998) <= (layer4_outputs(5829)) or (layer4_outputs(1964));
    layer5_outputs(1999) <= not((layer4_outputs(5450)) xor (layer4_outputs(6348)));
    layer5_outputs(2000) <= not(layer4_outputs(6070));
    layer5_outputs(2001) <= not((layer4_outputs(7491)) xor (layer4_outputs(5231)));
    layer5_outputs(2002) <= not(layer4_outputs(6401)) or (layer4_outputs(4014));
    layer5_outputs(2003) <= not(layer4_outputs(1888));
    layer5_outputs(2004) <= not(layer4_outputs(2494)) or (layer4_outputs(461));
    layer5_outputs(2005) <= not(layer4_outputs(1455));
    layer5_outputs(2006) <= not((layer4_outputs(4811)) or (layer4_outputs(1332)));
    layer5_outputs(2007) <= layer4_outputs(5366);
    layer5_outputs(2008) <= (layer4_outputs(4350)) and not (layer4_outputs(4703));
    layer5_outputs(2009) <= (layer4_outputs(952)) or (layer4_outputs(6543));
    layer5_outputs(2010) <= (layer4_outputs(214)) or (layer4_outputs(735));
    layer5_outputs(2011) <= not((layer4_outputs(4907)) xor (layer4_outputs(6238)));
    layer5_outputs(2012) <= not(layer4_outputs(2627));
    layer5_outputs(2013) <= layer4_outputs(5502);
    layer5_outputs(2014) <= not(layer4_outputs(1135)) or (layer4_outputs(640));
    layer5_outputs(2015) <= not(layer4_outputs(2396));
    layer5_outputs(2016) <= (layer4_outputs(7643)) or (layer4_outputs(7248));
    layer5_outputs(2017) <= not(layer4_outputs(6714)) or (layer4_outputs(6673));
    layer5_outputs(2018) <= (layer4_outputs(2148)) and (layer4_outputs(3337));
    layer5_outputs(2019) <= layer4_outputs(1078);
    layer5_outputs(2020) <= layer4_outputs(4217);
    layer5_outputs(2021) <= (layer4_outputs(7305)) and (layer4_outputs(621));
    layer5_outputs(2022) <= layer4_outputs(2474);
    layer5_outputs(2023) <= not(layer4_outputs(732));
    layer5_outputs(2024) <= layer4_outputs(93);
    layer5_outputs(2025) <= not(layer4_outputs(3109));
    layer5_outputs(2026) <= (layer4_outputs(413)) or (layer4_outputs(5917));
    layer5_outputs(2027) <= layer4_outputs(6587);
    layer5_outputs(2028) <= not((layer4_outputs(4060)) and (layer4_outputs(1200)));
    layer5_outputs(2029) <= not((layer4_outputs(1864)) or (layer4_outputs(7490)));
    layer5_outputs(2030) <= layer4_outputs(6722);
    layer5_outputs(2031) <= not((layer4_outputs(6076)) xor (layer4_outputs(5937)));
    layer5_outputs(2032) <= not(layer4_outputs(2754));
    layer5_outputs(2033) <= '0';
    layer5_outputs(2034) <= not(layer4_outputs(933)) or (layer4_outputs(1899));
    layer5_outputs(2035) <= not((layer4_outputs(3011)) or (layer4_outputs(6467)));
    layer5_outputs(2036) <= not((layer4_outputs(2305)) xor (layer4_outputs(65)));
    layer5_outputs(2037) <= layer4_outputs(2325);
    layer5_outputs(2038) <= not(layer4_outputs(6596));
    layer5_outputs(2039) <= not((layer4_outputs(1800)) or (layer4_outputs(6466)));
    layer5_outputs(2040) <= (layer4_outputs(2049)) xor (layer4_outputs(2928));
    layer5_outputs(2041) <= not(layer4_outputs(7063));
    layer5_outputs(2042) <= (layer4_outputs(3742)) xor (layer4_outputs(4084));
    layer5_outputs(2043) <= layer4_outputs(4363);
    layer5_outputs(2044) <= '1';
    layer5_outputs(2045) <= not(layer4_outputs(6617));
    layer5_outputs(2046) <= (layer4_outputs(728)) and not (layer4_outputs(377));
    layer5_outputs(2047) <= '1';
    layer5_outputs(2048) <= layer4_outputs(1007);
    layer5_outputs(2049) <= '0';
    layer5_outputs(2050) <= not((layer4_outputs(4958)) or (layer4_outputs(3727)));
    layer5_outputs(2051) <= (layer4_outputs(389)) and not (layer4_outputs(1436));
    layer5_outputs(2052) <= not((layer4_outputs(3053)) xor (layer4_outputs(5081)));
    layer5_outputs(2053) <= layer4_outputs(5635);
    layer5_outputs(2054) <= '0';
    layer5_outputs(2055) <= (layer4_outputs(1368)) xor (layer4_outputs(2930));
    layer5_outputs(2056) <= (layer4_outputs(4663)) or (layer4_outputs(1910));
    layer5_outputs(2057) <= layer4_outputs(6913);
    layer5_outputs(2058) <= (layer4_outputs(6324)) and not (layer4_outputs(695));
    layer5_outputs(2059) <= not(layer4_outputs(2856));
    layer5_outputs(2060) <= (layer4_outputs(72)) and (layer4_outputs(2369));
    layer5_outputs(2061) <= (layer4_outputs(1269)) and not (layer4_outputs(6181));
    layer5_outputs(2062) <= (layer4_outputs(7149)) xor (layer4_outputs(2144));
    layer5_outputs(2063) <= layer4_outputs(5313);
    layer5_outputs(2064) <= '1';
    layer5_outputs(2065) <= not(layer4_outputs(2314));
    layer5_outputs(2066) <= (layer4_outputs(324)) and not (layer4_outputs(2385));
    layer5_outputs(2067) <= layer4_outputs(2936);
    layer5_outputs(2068) <= layer4_outputs(2797);
    layer5_outputs(2069) <= not(layer4_outputs(2722));
    layer5_outputs(2070) <= not((layer4_outputs(3480)) xor (layer4_outputs(5408)));
    layer5_outputs(2071) <= layer4_outputs(2875);
    layer5_outputs(2072) <= (layer4_outputs(7326)) or (layer4_outputs(6286));
    layer5_outputs(2073) <= '0';
    layer5_outputs(2074) <= (layer4_outputs(1386)) and not (layer4_outputs(3430));
    layer5_outputs(2075) <= not((layer4_outputs(1343)) and (layer4_outputs(761)));
    layer5_outputs(2076) <= not(layer4_outputs(7127));
    layer5_outputs(2077) <= layer4_outputs(6035);
    layer5_outputs(2078) <= (layer4_outputs(4133)) and not (layer4_outputs(2508));
    layer5_outputs(2079) <= not(layer4_outputs(4065));
    layer5_outputs(2080) <= not(layer4_outputs(2171));
    layer5_outputs(2081) <= not(layer4_outputs(2895));
    layer5_outputs(2082) <= not(layer4_outputs(4593));
    layer5_outputs(2083) <= not((layer4_outputs(136)) xor (layer4_outputs(7526)));
    layer5_outputs(2084) <= layer4_outputs(1985);
    layer5_outputs(2085) <= layer4_outputs(2318);
    layer5_outputs(2086) <= not(layer4_outputs(149)) or (layer4_outputs(783));
    layer5_outputs(2087) <= not(layer4_outputs(3385));
    layer5_outputs(2088) <= not(layer4_outputs(2665)) or (layer4_outputs(6642));
    layer5_outputs(2089) <= layer4_outputs(2871);
    layer5_outputs(2090) <= (layer4_outputs(1201)) and not (layer4_outputs(7612));
    layer5_outputs(2091) <= (layer4_outputs(4573)) and (layer4_outputs(5586));
    layer5_outputs(2092) <= not(layer4_outputs(3152));
    layer5_outputs(2093) <= not((layer4_outputs(2048)) xor (layer4_outputs(2202)));
    layer5_outputs(2094) <= not(layer4_outputs(3356)) or (layer4_outputs(3320));
    layer5_outputs(2095) <= not(layer4_outputs(2132));
    layer5_outputs(2096) <= (layer4_outputs(5270)) xor (layer4_outputs(948));
    layer5_outputs(2097) <= not(layer4_outputs(4282)) or (layer4_outputs(1321));
    layer5_outputs(2098) <= layer4_outputs(5620);
    layer5_outputs(2099) <= not(layer4_outputs(4170));
    layer5_outputs(2100) <= not(layer4_outputs(2327));
    layer5_outputs(2101) <= not(layer4_outputs(6352)) or (layer4_outputs(2606));
    layer5_outputs(2102) <= not(layer4_outputs(5796));
    layer5_outputs(2103) <= (layer4_outputs(7338)) and not (layer4_outputs(620));
    layer5_outputs(2104) <= layer4_outputs(6507);
    layer5_outputs(2105) <= layer4_outputs(6207);
    layer5_outputs(2106) <= not(layer4_outputs(4429)) or (layer4_outputs(1980));
    layer5_outputs(2107) <= layer4_outputs(5378);
    layer5_outputs(2108) <= '1';
    layer5_outputs(2109) <= (layer4_outputs(3999)) and (layer4_outputs(5120));
    layer5_outputs(2110) <= (layer4_outputs(3934)) or (layer4_outputs(7427));
    layer5_outputs(2111) <= layer4_outputs(4951);
    layer5_outputs(2112) <= not(layer4_outputs(5510));
    layer5_outputs(2113) <= not(layer4_outputs(6033)) or (layer4_outputs(4810));
    layer5_outputs(2114) <= (layer4_outputs(1499)) and not (layer4_outputs(7532));
    layer5_outputs(2115) <= (layer4_outputs(6010)) xor (layer4_outputs(2048));
    layer5_outputs(2116) <= not((layer4_outputs(3513)) xor (layer4_outputs(6254)));
    layer5_outputs(2117) <= (layer4_outputs(5431)) and not (layer4_outputs(3489));
    layer5_outputs(2118) <= (layer4_outputs(2400)) and (layer4_outputs(866));
    layer5_outputs(2119) <= layer4_outputs(5417);
    layer5_outputs(2120) <= layer4_outputs(6422);
    layer5_outputs(2121) <= not(layer4_outputs(318));
    layer5_outputs(2122) <= layer4_outputs(6946);
    layer5_outputs(2123) <= '0';
    layer5_outputs(2124) <= not(layer4_outputs(3439)) or (layer4_outputs(1887));
    layer5_outputs(2125) <= '1';
    layer5_outputs(2126) <= '1';
    layer5_outputs(2127) <= (layer4_outputs(3823)) or (layer4_outputs(1018));
    layer5_outputs(2128) <= layer4_outputs(1456);
    layer5_outputs(2129) <= not(layer4_outputs(4675));
    layer5_outputs(2130) <= not(layer4_outputs(2261));
    layer5_outputs(2131) <= layer4_outputs(1969);
    layer5_outputs(2132) <= not(layer4_outputs(3801));
    layer5_outputs(2133) <= not((layer4_outputs(189)) xor (layer4_outputs(4079)));
    layer5_outputs(2134) <= layer4_outputs(3155);
    layer5_outputs(2135) <= layer4_outputs(4787);
    layer5_outputs(2136) <= (layer4_outputs(6282)) and not (layer4_outputs(7403));
    layer5_outputs(2137) <= not(layer4_outputs(4392));
    layer5_outputs(2138) <= (layer4_outputs(679)) xor (layer4_outputs(1340));
    layer5_outputs(2139) <= (layer4_outputs(2771)) and not (layer4_outputs(7059));
    layer5_outputs(2140) <= layer4_outputs(1217);
    layer5_outputs(2141) <= layer4_outputs(4962);
    layer5_outputs(2142) <= not(layer4_outputs(3632)) or (layer4_outputs(784));
    layer5_outputs(2143) <= layer4_outputs(294);
    layer5_outputs(2144) <= not(layer4_outputs(7019));
    layer5_outputs(2145) <= layer4_outputs(7649);
    layer5_outputs(2146) <= not(layer4_outputs(6015));
    layer5_outputs(2147) <= not((layer4_outputs(490)) xor (layer4_outputs(262)));
    layer5_outputs(2148) <= layer4_outputs(2648);
    layer5_outputs(2149) <= layer4_outputs(4578);
    layer5_outputs(2150) <= not(layer4_outputs(3996));
    layer5_outputs(2151) <= (layer4_outputs(3544)) or (layer4_outputs(6118));
    layer5_outputs(2152) <= layer4_outputs(6231);
    layer5_outputs(2153) <= '0';
    layer5_outputs(2154) <= not(layer4_outputs(6442));
    layer5_outputs(2155) <= (layer4_outputs(4955)) or (layer4_outputs(440));
    layer5_outputs(2156) <= '1';
    layer5_outputs(2157) <= not(layer4_outputs(118)) or (layer4_outputs(4489));
    layer5_outputs(2158) <= not(layer4_outputs(6027)) or (layer4_outputs(328));
    layer5_outputs(2159) <= not(layer4_outputs(1515));
    layer5_outputs(2160) <= (layer4_outputs(6062)) and (layer4_outputs(4667));
    layer5_outputs(2161) <= '1';
    layer5_outputs(2162) <= not(layer4_outputs(2748));
    layer5_outputs(2163) <= not((layer4_outputs(342)) or (layer4_outputs(4227)));
    layer5_outputs(2164) <= not(layer4_outputs(5295)) or (layer4_outputs(5095));
    layer5_outputs(2165) <= layer4_outputs(1103);
    layer5_outputs(2166) <= layer4_outputs(3540);
    layer5_outputs(2167) <= (layer4_outputs(7244)) xor (layer4_outputs(2343));
    layer5_outputs(2168) <= (layer4_outputs(224)) and not (layer4_outputs(5040));
    layer5_outputs(2169) <= (layer4_outputs(7261)) or (layer4_outputs(2137));
    layer5_outputs(2170) <= layer4_outputs(4976);
    layer5_outputs(2171) <= layer4_outputs(1244);
    layer5_outputs(2172) <= (layer4_outputs(2573)) xor (layer4_outputs(6350));
    layer5_outputs(2173) <= layer4_outputs(547);
    layer5_outputs(2174) <= layer4_outputs(6765);
    layer5_outputs(2175) <= not(layer4_outputs(2956));
    layer5_outputs(2176) <= (layer4_outputs(5287)) xor (layer4_outputs(438));
    layer5_outputs(2177) <= not((layer4_outputs(1541)) xor (layer4_outputs(7074)));
    layer5_outputs(2178) <= not(layer4_outputs(3035));
    layer5_outputs(2179) <= not((layer4_outputs(6506)) or (layer4_outputs(7174)));
    layer5_outputs(2180) <= not(layer4_outputs(7562));
    layer5_outputs(2181) <= not((layer4_outputs(6428)) xor (layer4_outputs(7144)));
    layer5_outputs(2182) <= not(layer4_outputs(5544));
    layer5_outputs(2183) <= not(layer4_outputs(122));
    layer5_outputs(2184) <= not(layer4_outputs(5272));
    layer5_outputs(2185) <= layer4_outputs(4927);
    layer5_outputs(2186) <= layer4_outputs(1753);
    layer5_outputs(2187) <= layer4_outputs(788);
    layer5_outputs(2188) <= not(layer4_outputs(1771));
    layer5_outputs(2189) <= not(layer4_outputs(5117));
    layer5_outputs(2190) <= not(layer4_outputs(6755));
    layer5_outputs(2191) <= (layer4_outputs(7075)) and not (layer4_outputs(6390));
    layer5_outputs(2192) <= not(layer4_outputs(6989));
    layer5_outputs(2193) <= layer4_outputs(5198);
    layer5_outputs(2194) <= not((layer4_outputs(3772)) and (layer4_outputs(168)));
    layer5_outputs(2195) <= (layer4_outputs(2642)) and (layer4_outputs(3295));
    layer5_outputs(2196) <= not(layer4_outputs(3941));
    layer5_outputs(2197) <= not(layer4_outputs(1224));
    layer5_outputs(2198) <= not(layer4_outputs(7159)) or (layer4_outputs(6140));
    layer5_outputs(2199) <= layer4_outputs(1483);
    layer5_outputs(2200) <= (layer4_outputs(48)) and not (layer4_outputs(2235));
    layer5_outputs(2201) <= not((layer4_outputs(6871)) or (layer4_outputs(3716)));
    layer5_outputs(2202) <= not(layer4_outputs(3063));
    layer5_outputs(2203) <= not(layer4_outputs(2099)) or (layer4_outputs(949));
    layer5_outputs(2204) <= not(layer4_outputs(7392)) or (layer4_outputs(4518));
    layer5_outputs(2205) <= (layer4_outputs(7619)) xor (layer4_outputs(6781));
    layer5_outputs(2206) <= not(layer4_outputs(7420)) or (layer4_outputs(6450));
    layer5_outputs(2207) <= layer4_outputs(6044);
    layer5_outputs(2208) <= layer4_outputs(5407);
    layer5_outputs(2209) <= not(layer4_outputs(7343));
    layer5_outputs(2210) <= not(layer4_outputs(1838));
    layer5_outputs(2211) <= (layer4_outputs(5346)) xor (layer4_outputs(4645));
    layer5_outputs(2212) <= not((layer4_outputs(3520)) and (layer4_outputs(2384)));
    layer5_outputs(2213) <= not((layer4_outputs(2500)) xor (layer4_outputs(3701)));
    layer5_outputs(2214) <= not((layer4_outputs(5008)) or (layer4_outputs(3822)));
    layer5_outputs(2215) <= not((layer4_outputs(2743)) xor (layer4_outputs(655)));
    layer5_outputs(2216) <= not(layer4_outputs(1785));
    layer5_outputs(2217) <= layer4_outputs(6988);
    layer5_outputs(2218) <= not(layer4_outputs(5301)) or (layer4_outputs(2595));
    layer5_outputs(2219) <= not(layer4_outputs(1546));
    layer5_outputs(2220) <= (layer4_outputs(5738)) and not (layer4_outputs(3161));
    layer5_outputs(2221) <= not((layer4_outputs(3516)) xor (layer4_outputs(4824)));
    layer5_outputs(2222) <= not(layer4_outputs(1617));
    layer5_outputs(2223) <= (layer4_outputs(7574)) and (layer4_outputs(1109));
    layer5_outputs(2224) <= layer4_outputs(467);
    layer5_outputs(2225) <= (layer4_outputs(4165)) xor (layer4_outputs(364));
    layer5_outputs(2226) <= not(layer4_outputs(7368)) or (layer4_outputs(5985));
    layer5_outputs(2227) <= layer4_outputs(6843);
    layer5_outputs(2228) <= '1';
    layer5_outputs(2229) <= not((layer4_outputs(2164)) or (layer4_outputs(4308)));
    layer5_outputs(2230) <= not(layer4_outputs(4179));
    layer5_outputs(2231) <= not(layer4_outputs(6291));
    layer5_outputs(2232) <= layer4_outputs(5988);
    layer5_outputs(2233) <= not(layer4_outputs(5570));
    layer5_outputs(2234) <= (layer4_outputs(5543)) and (layer4_outputs(5640));
    layer5_outputs(2235) <= layer4_outputs(1403);
    layer5_outputs(2236) <= (layer4_outputs(4666)) or (layer4_outputs(11));
    layer5_outputs(2237) <= (layer4_outputs(4852)) or (layer4_outputs(1482));
    layer5_outputs(2238) <= '1';
    layer5_outputs(2239) <= not(layer4_outputs(1165));
    layer5_outputs(2240) <= not(layer4_outputs(912)) or (layer4_outputs(3129));
    layer5_outputs(2241) <= not(layer4_outputs(5939));
    layer5_outputs(2242) <= not(layer4_outputs(7630));
    layer5_outputs(2243) <= layer4_outputs(5605);
    layer5_outputs(2244) <= not((layer4_outputs(939)) and (layer4_outputs(2383)));
    layer5_outputs(2245) <= (layer4_outputs(5850)) and not (layer4_outputs(1213));
    layer5_outputs(2246) <= (layer4_outputs(1628)) and not (layer4_outputs(365));
    layer5_outputs(2247) <= not(layer4_outputs(1486)) or (layer4_outputs(835));
    layer5_outputs(2248) <= (layer4_outputs(7209)) or (layer4_outputs(1635));
    layer5_outputs(2249) <= layer4_outputs(1116);
    layer5_outputs(2250) <= not(layer4_outputs(5170)) or (layer4_outputs(5024));
    layer5_outputs(2251) <= not(layer4_outputs(4977));
    layer5_outputs(2252) <= layer4_outputs(7305);
    layer5_outputs(2253) <= layer4_outputs(2825);
    layer5_outputs(2254) <= layer4_outputs(6770);
    layer5_outputs(2255) <= (layer4_outputs(5362)) and not (layer4_outputs(965));
    layer5_outputs(2256) <= not(layer4_outputs(3513));
    layer5_outputs(2257) <= not(layer4_outputs(2864));
    layer5_outputs(2258) <= not(layer4_outputs(665));
    layer5_outputs(2259) <= not(layer4_outputs(1546));
    layer5_outputs(2260) <= layer4_outputs(2100);
    layer5_outputs(2261) <= not(layer4_outputs(330)) or (layer4_outputs(438));
    layer5_outputs(2262) <= (layer4_outputs(5456)) or (layer4_outputs(1163));
    layer5_outputs(2263) <= not(layer4_outputs(6142)) or (layer4_outputs(103));
    layer5_outputs(2264) <= layer4_outputs(3434);
    layer5_outputs(2265) <= not(layer4_outputs(4027)) or (layer4_outputs(2941));
    layer5_outputs(2266) <= not(layer4_outputs(7234));
    layer5_outputs(2267) <= not(layer4_outputs(4737));
    layer5_outputs(2268) <= layer4_outputs(4733);
    layer5_outputs(2269) <= (layer4_outputs(5579)) and (layer4_outputs(1408));
    layer5_outputs(2270) <= (layer4_outputs(7147)) or (layer4_outputs(6470));
    layer5_outputs(2271) <= not((layer4_outputs(1261)) and (layer4_outputs(2465)));
    layer5_outputs(2272) <= not((layer4_outputs(5156)) and (layer4_outputs(533)));
    layer5_outputs(2273) <= not((layer4_outputs(1046)) or (layer4_outputs(1317)));
    layer5_outputs(2274) <= not(layer4_outputs(3471)) or (layer4_outputs(6272));
    layer5_outputs(2275) <= not(layer4_outputs(3132));
    layer5_outputs(2276) <= '1';
    layer5_outputs(2277) <= not((layer4_outputs(3556)) xor (layer4_outputs(652)));
    layer5_outputs(2278) <= not((layer4_outputs(6863)) or (layer4_outputs(4482)));
    layer5_outputs(2279) <= layer4_outputs(2907);
    layer5_outputs(2280) <= (layer4_outputs(356)) and not (layer4_outputs(2620));
    layer5_outputs(2281) <= (layer4_outputs(7542)) and not (layer4_outputs(7082));
    layer5_outputs(2282) <= not(layer4_outputs(3066));
    layer5_outputs(2283) <= '1';
    layer5_outputs(2284) <= not((layer4_outputs(3642)) xor (layer4_outputs(7016)));
    layer5_outputs(2285) <= layer4_outputs(4041);
    layer5_outputs(2286) <= not(layer4_outputs(6537));
    layer5_outputs(2287) <= not(layer4_outputs(6030));
    layer5_outputs(2288) <= layer4_outputs(3189);
    layer5_outputs(2289) <= not(layer4_outputs(3542)) or (layer4_outputs(3006));
    layer5_outputs(2290) <= not((layer4_outputs(1345)) xor (layer4_outputs(4448)));
    layer5_outputs(2291) <= (layer4_outputs(4460)) and not (layer4_outputs(5353));
    layer5_outputs(2292) <= layer4_outputs(1495);
    layer5_outputs(2293) <= not(layer4_outputs(7056));
    layer5_outputs(2294) <= not((layer4_outputs(5535)) xor (layer4_outputs(6145)));
    layer5_outputs(2295) <= not(layer4_outputs(3172));
    layer5_outputs(2296) <= layer4_outputs(4790);
    layer5_outputs(2297) <= not((layer4_outputs(6054)) and (layer4_outputs(6571)));
    layer5_outputs(2298) <= not((layer4_outputs(7384)) and (layer4_outputs(471)));
    layer5_outputs(2299) <= layer4_outputs(7592);
    layer5_outputs(2300) <= not((layer4_outputs(2283)) or (layer4_outputs(1473)));
    layer5_outputs(2301) <= not(layer4_outputs(7505));
    layer5_outputs(2302) <= not(layer4_outputs(6246));
    layer5_outputs(2303) <= layer4_outputs(6692);
    layer5_outputs(2304) <= layer4_outputs(517);
    layer5_outputs(2305) <= not((layer4_outputs(3399)) and (layer4_outputs(6439)));
    layer5_outputs(2306) <= not((layer4_outputs(5992)) or (layer4_outputs(7517)));
    layer5_outputs(2307) <= not(layer4_outputs(2626));
    layer5_outputs(2308) <= (layer4_outputs(3266)) xor (layer4_outputs(3466));
    layer5_outputs(2309) <= not(layer4_outputs(4172));
    layer5_outputs(2310) <= layer4_outputs(2155);
    layer5_outputs(2311) <= not(layer4_outputs(6982));
    layer5_outputs(2312) <= layer4_outputs(5594);
    layer5_outputs(2313) <= '0';
    layer5_outputs(2314) <= not(layer4_outputs(5839));
    layer5_outputs(2315) <= not(layer4_outputs(4367)) or (layer4_outputs(1138));
    layer5_outputs(2316) <= '1';
    layer5_outputs(2317) <= not((layer4_outputs(7425)) and (layer4_outputs(3722)));
    layer5_outputs(2318) <= layer4_outputs(3351);
    layer5_outputs(2319) <= (layer4_outputs(2563)) and (layer4_outputs(3379));
    layer5_outputs(2320) <= not(layer4_outputs(1645)) or (layer4_outputs(3433));
    layer5_outputs(2321) <= '0';
    layer5_outputs(2322) <= not(layer4_outputs(1873)) or (layer4_outputs(2814));
    layer5_outputs(2323) <= not(layer4_outputs(7101)) or (layer4_outputs(451));
    layer5_outputs(2324) <= not(layer4_outputs(1744)) or (layer4_outputs(6743));
    layer5_outputs(2325) <= (layer4_outputs(6350)) xor (layer4_outputs(3850));
    layer5_outputs(2326) <= layer4_outputs(6521);
    layer5_outputs(2327) <= not((layer4_outputs(3649)) and (layer4_outputs(337)));
    layer5_outputs(2328) <= (layer4_outputs(4338)) and not (layer4_outputs(1152));
    layer5_outputs(2329) <= not((layer4_outputs(2597)) xor (layer4_outputs(3166)));
    layer5_outputs(2330) <= (layer4_outputs(5875)) and not (layer4_outputs(4677));
    layer5_outputs(2331) <= (layer4_outputs(5128)) xor (layer4_outputs(908));
    layer5_outputs(2332) <= layer4_outputs(6963);
    layer5_outputs(2333) <= (layer4_outputs(1982)) xor (layer4_outputs(3831));
    layer5_outputs(2334) <= layer4_outputs(5512);
    layer5_outputs(2335) <= not(layer4_outputs(6002));
    layer5_outputs(2336) <= not((layer4_outputs(6028)) or (layer4_outputs(3994)));
    layer5_outputs(2337) <= not(layer4_outputs(1047));
    layer5_outputs(2338) <= layer4_outputs(6501);
    layer5_outputs(2339) <= (layer4_outputs(6084)) and not (layer4_outputs(2472));
    layer5_outputs(2340) <= '0';
    layer5_outputs(2341) <= not(layer4_outputs(822));
    layer5_outputs(2342) <= not((layer4_outputs(6418)) or (layer4_outputs(7638)));
    layer5_outputs(2343) <= not(layer4_outputs(1996));
    layer5_outputs(2344) <= not((layer4_outputs(4870)) and (layer4_outputs(5938)));
    layer5_outputs(2345) <= not(layer4_outputs(6336));
    layer5_outputs(2346) <= layer4_outputs(4945);
    layer5_outputs(2347) <= not(layer4_outputs(1634));
    layer5_outputs(2348) <= layer4_outputs(4628);
    layer5_outputs(2349) <= not((layer4_outputs(2394)) xor (layer4_outputs(1776)));
    layer5_outputs(2350) <= (layer4_outputs(1746)) and not (layer4_outputs(7004));
    layer5_outputs(2351) <= layer4_outputs(6360);
    layer5_outputs(2352) <= not(layer4_outputs(2511));
    layer5_outputs(2353) <= layer4_outputs(4404);
    layer5_outputs(2354) <= not(layer4_outputs(4050));
    layer5_outputs(2355) <= not((layer4_outputs(6594)) and (layer4_outputs(391)));
    layer5_outputs(2356) <= not(layer4_outputs(6009));
    layer5_outputs(2357) <= layer4_outputs(4412);
    layer5_outputs(2358) <= '0';
    layer5_outputs(2359) <= (layer4_outputs(1537)) and not (layer4_outputs(6379));
    layer5_outputs(2360) <= (layer4_outputs(2459)) or (layer4_outputs(4139));
    layer5_outputs(2361) <= layer4_outputs(5812);
    layer5_outputs(2362) <= not((layer4_outputs(4859)) xor (layer4_outputs(5843)));
    layer5_outputs(2363) <= (layer4_outputs(1050)) and not (layer4_outputs(257));
    layer5_outputs(2364) <= not(layer4_outputs(975));
    layer5_outputs(2365) <= '1';
    layer5_outputs(2366) <= layer4_outputs(4537);
    layer5_outputs(2367) <= not(layer4_outputs(6219));
    layer5_outputs(2368) <= (layer4_outputs(5816)) and not (layer4_outputs(7626));
    layer5_outputs(2369) <= layer4_outputs(5190);
    layer5_outputs(2370) <= '1';
    layer5_outputs(2371) <= layer4_outputs(917);
    layer5_outputs(2372) <= not(layer4_outputs(1351));
    layer5_outputs(2373) <= not(layer4_outputs(3237));
    layer5_outputs(2374) <= not((layer4_outputs(1872)) xor (layer4_outputs(6017)));
    layer5_outputs(2375) <= not(layer4_outputs(2763)) or (layer4_outputs(6329));
    layer5_outputs(2376) <= layer4_outputs(310);
    layer5_outputs(2377) <= (layer4_outputs(420)) or (layer4_outputs(6507));
    layer5_outputs(2378) <= not(layer4_outputs(2992));
    layer5_outputs(2379) <= layer4_outputs(2481);
    layer5_outputs(2380) <= (layer4_outputs(6768)) or (layer4_outputs(3108));
    layer5_outputs(2381) <= layer4_outputs(7403);
    layer5_outputs(2382) <= layer4_outputs(6867);
    layer5_outputs(2383) <= (layer4_outputs(3717)) and not (layer4_outputs(1770));
    layer5_outputs(2384) <= not(layer4_outputs(1183));
    layer5_outputs(2385) <= not(layer4_outputs(5691));
    layer5_outputs(2386) <= not(layer4_outputs(54));
    layer5_outputs(2387) <= layer4_outputs(807);
    layer5_outputs(2388) <= '0';
    layer5_outputs(2389) <= not((layer4_outputs(4809)) and (layer4_outputs(3792)));
    layer5_outputs(2390) <= not(layer4_outputs(6098));
    layer5_outputs(2391) <= layer4_outputs(2230);
    layer5_outputs(2392) <= (layer4_outputs(5842)) and not (layer4_outputs(5696));
    layer5_outputs(2393) <= not(layer4_outputs(6709));
    layer5_outputs(2394) <= not(layer4_outputs(6302));
    layer5_outputs(2395) <= (layer4_outputs(4572)) and not (layer4_outputs(4931));
    layer5_outputs(2396) <= not(layer4_outputs(7213));
    layer5_outputs(2397) <= not((layer4_outputs(5035)) xor (layer4_outputs(1281)));
    layer5_outputs(2398) <= not(layer4_outputs(2295));
    layer5_outputs(2399) <= not(layer4_outputs(429));
    layer5_outputs(2400) <= (layer4_outputs(1075)) and (layer4_outputs(6163));
    layer5_outputs(2401) <= layer4_outputs(5676);
    layer5_outputs(2402) <= not(layer4_outputs(5089));
    layer5_outputs(2403) <= not(layer4_outputs(2493));
    layer5_outputs(2404) <= not(layer4_outputs(2442));
    layer5_outputs(2405) <= (layer4_outputs(7028)) and (layer4_outputs(2449));
    layer5_outputs(2406) <= (layer4_outputs(3838)) and (layer4_outputs(449));
    layer5_outputs(2407) <= not(layer4_outputs(6614));
    layer5_outputs(2408) <= (layer4_outputs(3661)) or (layer4_outputs(3759));
    layer5_outputs(2409) <= (layer4_outputs(4731)) and not (layer4_outputs(4199));
    layer5_outputs(2410) <= not(layer4_outputs(7487));
    layer5_outputs(2411) <= not(layer4_outputs(2459));
    layer5_outputs(2412) <= not((layer4_outputs(4739)) and (layer4_outputs(320)));
    layer5_outputs(2413) <= not(layer4_outputs(374));
    layer5_outputs(2414) <= not((layer4_outputs(4562)) and (layer4_outputs(1501)));
    layer5_outputs(2415) <= not(layer4_outputs(2613));
    layer5_outputs(2416) <= layer4_outputs(902);
    layer5_outputs(2417) <= layer4_outputs(990);
    layer5_outputs(2418) <= not(layer4_outputs(7147));
    layer5_outputs(2419) <= not((layer4_outputs(5953)) xor (layer4_outputs(972)));
    layer5_outputs(2420) <= layer4_outputs(2267);
    layer5_outputs(2421) <= not(layer4_outputs(1656));
    layer5_outputs(2422) <= not(layer4_outputs(5461));
    layer5_outputs(2423) <= not(layer4_outputs(4169));
    layer5_outputs(2424) <= (layer4_outputs(1674)) xor (layer4_outputs(6670));
    layer5_outputs(2425) <= (layer4_outputs(2284)) and not (layer4_outputs(3316));
    layer5_outputs(2426) <= not(layer4_outputs(7477));
    layer5_outputs(2427) <= not(layer4_outputs(1906));
    layer5_outputs(2428) <= (layer4_outputs(7192)) and not (layer4_outputs(1594));
    layer5_outputs(2429) <= not(layer4_outputs(7406));
    layer5_outputs(2430) <= layer4_outputs(3224);
    layer5_outputs(2431) <= (layer4_outputs(6989)) and not (layer4_outputs(1245));
    layer5_outputs(2432) <= layer4_outputs(2256);
    layer5_outputs(2433) <= not((layer4_outputs(2082)) or (layer4_outputs(6976)));
    layer5_outputs(2434) <= not(layer4_outputs(6295)) or (layer4_outputs(502));
    layer5_outputs(2435) <= (layer4_outputs(751)) and (layer4_outputs(248));
    layer5_outputs(2436) <= layer4_outputs(7178);
    layer5_outputs(2437) <= not(layer4_outputs(4029));
    layer5_outputs(2438) <= (layer4_outputs(6146)) and not (layer4_outputs(897));
    layer5_outputs(2439) <= not(layer4_outputs(6180));
    layer5_outputs(2440) <= not(layer4_outputs(7481));
    layer5_outputs(2441) <= not(layer4_outputs(2174));
    layer5_outputs(2442) <= (layer4_outputs(5237)) and (layer4_outputs(2682));
    layer5_outputs(2443) <= not(layer4_outputs(3022)) or (layer4_outputs(3915));
    layer5_outputs(2444) <= (layer4_outputs(1886)) xor (layer4_outputs(1341));
    layer5_outputs(2445) <= not(layer4_outputs(6560));
    layer5_outputs(2446) <= not(layer4_outputs(6413));
    layer5_outputs(2447) <= not(layer4_outputs(6716));
    layer5_outputs(2448) <= layer4_outputs(5984);
    layer5_outputs(2449) <= layer4_outputs(122);
    layer5_outputs(2450) <= not(layer4_outputs(372));
    layer5_outputs(2451) <= layer4_outputs(1958);
    layer5_outputs(2452) <= (layer4_outputs(6373)) xor (layer4_outputs(6106));
    layer5_outputs(2453) <= layer4_outputs(3962);
    layer5_outputs(2454) <= not(layer4_outputs(4378));
    layer5_outputs(2455) <= not(layer4_outputs(4502)) or (layer4_outputs(6496));
    layer5_outputs(2456) <= layer4_outputs(6847);
    layer5_outputs(2457) <= not(layer4_outputs(1781));
    layer5_outputs(2458) <= not(layer4_outputs(3360));
    layer5_outputs(2459) <= (layer4_outputs(3871)) or (layer4_outputs(3060));
    layer5_outputs(2460) <= not((layer4_outputs(3493)) or (layer4_outputs(1844)));
    layer5_outputs(2461) <= not(layer4_outputs(5623)) or (layer4_outputs(2951));
    layer5_outputs(2462) <= layer4_outputs(1076);
    layer5_outputs(2463) <= layer4_outputs(3995);
    layer5_outputs(2464) <= (layer4_outputs(3422)) xor (layer4_outputs(6226));
    layer5_outputs(2465) <= layer4_outputs(1567);
    layer5_outputs(2466) <= (layer4_outputs(4467)) and not (layer4_outputs(1734));
    layer5_outputs(2467) <= layer4_outputs(3078);
    layer5_outputs(2468) <= not((layer4_outputs(1956)) xor (layer4_outputs(7467)));
    layer5_outputs(2469) <= not(layer4_outputs(5554));
    layer5_outputs(2470) <= (layer4_outputs(1218)) and not (layer4_outputs(2328));
    layer5_outputs(2471) <= not(layer4_outputs(314));
    layer5_outputs(2472) <= not(layer4_outputs(5744));
    layer5_outputs(2473) <= not(layer4_outputs(5765));
    layer5_outputs(2474) <= (layer4_outputs(3227)) and (layer4_outputs(2953));
    layer5_outputs(2475) <= (layer4_outputs(5525)) and not (layer4_outputs(6383));
    layer5_outputs(2476) <= (layer4_outputs(4429)) or (layer4_outputs(3669));
    layer5_outputs(2477) <= not(layer4_outputs(4021));
    layer5_outputs(2478) <= not(layer4_outputs(340));
    layer5_outputs(2479) <= layer4_outputs(7585);
    layer5_outputs(2480) <= not((layer4_outputs(207)) or (layer4_outputs(6431)));
    layer5_outputs(2481) <= not(layer4_outputs(6974));
    layer5_outputs(2482) <= layer4_outputs(4286);
    layer5_outputs(2483) <= (layer4_outputs(40)) and not (layer4_outputs(2380));
    layer5_outputs(2484) <= (layer4_outputs(5258)) and (layer4_outputs(1496));
    layer5_outputs(2485) <= (layer4_outputs(4979)) xor (layer4_outputs(5650));
    layer5_outputs(2486) <= not((layer4_outputs(3362)) xor (layer4_outputs(5889)));
    layer5_outputs(2487) <= not(layer4_outputs(3199));
    layer5_outputs(2488) <= layer4_outputs(7329);
    layer5_outputs(2489) <= layer4_outputs(2185);
    layer5_outputs(2490) <= not(layer4_outputs(7322)) or (layer4_outputs(2077));
    layer5_outputs(2491) <= layer4_outputs(6935);
    layer5_outputs(2492) <= not((layer4_outputs(809)) and (layer4_outputs(6645)));
    layer5_outputs(2493) <= not(layer4_outputs(1478));
    layer5_outputs(2494) <= not((layer4_outputs(150)) and (layer4_outputs(1311)));
    layer5_outputs(2495) <= layer4_outputs(5787);
    layer5_outputs(2496) <= layer4_outputs(4401);
    layer5_outputs(2497) <= (layer4_outputs(3878)) and not (layer4_outputs(7143));
    layer5_outputs(2498) <= (layer4_outputs(6865)) or (layer4_outputs(1299));
    layer5_outputs(2499) <= not(layer4_outputs(3306));
    layer5_outputs(2500) <= layer4_outputs(3874);
    layer5_outputs(2501) <= layer4_outputs(2639);
    layer5_outputs(2502) <= not(layer4_outputs(5372));
    layer5_outputs(2503) <= (layer4_outputs(2506)) xor (layer4_outputs(2338));
    layer5_outputs(2504) <= (layer4_outputs(1184)) and not (layer4_outputs(7080));
    layer5_outputs(2505) <= layer4_outputs(4693);
    layer5_outputs(2506) <= layer4_outputs(271);
    layer5_outputs(2507) <= layer4_outputs(4325);
    layer5_outputs(2508) <= not(layer4_outputs(5868)) or (layer4_outputs(3019));
    layer5_outputs(2509) <= layer4_outputs(2091);
    layer5_outputs(2510) <= not((layer4_outputs(308)) and (layer4_outputs(857)));
    layer5_outputs(2511) <= not(layer4_outputs(3225));
    layer5_outputs(2512) <= (layer4_outputs(568)) and not (layer4_outputs(1288));
    layer5_outputs(2513) <= not(layer4_outputs(1468));
    layer5_outputs(2514) <= layer4_outputs(3564);
    layer5_outputs(2515) <= layer4_outputs(4055);
    layer5_outputs(2516) <= (layer4_outputs(5514)) and not (layer4_outputs(5203));
    layer5_outputs(2517) <= layer4_outputs(7155);
    layer5_outputs(2518) <= not(layer4_outputs(2526));
    layer5_outputs(2519) <= not((layer4_outputs(4867)) xor (layer4_outputs(7334)));
    layer5_outputs(2520) <= not(layer4_outputs(4781));
    layer5_outputs(2521) <= layer4_outputs(4708);
    layer5_outputs(2522) <= not(layer4_outputs(3356));
    layer5_outputs(2523) <= not((layer4_outputs(1121)) or (layer4_outputs(4089)));
    layer5_outputs(2524) <= not(layer4_outputs(4042));
    layer5_outputs(2525) <= (layer4_outputs(2990)) or (layer4_outputs(5590));
    layer5_outputs(2526) <= '0';
    layer5_outputs(2527) <= (layer4_outputs(659)) and (layer4_outputs(2528));
    layer5_outputs(2528) <= layer4_outputs(4735);
    layer5_outputs(2529) <= (layer4_outputs(1559)) and not (layer4_outputs(3498));
    layer5_outputs(2530) <= layer4_outputs(5865);
    layer5_outputs(2531) <= (layer4_outputs(6943)) and not (layer4_outputs(6362));
    layer5_outputs(2532) <= layer4_outputs(6353);
    layer5_outputs(2533) <= not(layer4_outputs(5817)) or (layer4_outputs(7271));
    layer5_outputs(2534) <= layer4_outputs(772);
    layer5_outputs(2535) <= layer4_outputs(5152);
    layer5_outputs(2536) <= layer4_outputs(940);
    layer5_outputs(2537) <= (layer4_outputs(4160)) and (layer4_outputs(2468));
    layer5_outputs(2538) <= '1';
    layer5_outputs(2539) <= (layer4_outputs(7163)) or (layer4_outputs(3961));
    layer5_outputs(2540) <= not(layer4_outputs(4191));
    layer5_outputs(2541) <= not(layer4_outputs(2690));
    layer5_outputs(2542) <= not(layer4_outputs(5865));
    layer5_outputs(2543) <= layer4_outputs(673);
    layer5_outputs(2544) <= layer4_outputs(2387);
    layer5_outputs(2545) <= '0';
    layer5_outputs(2546) <= (layer4_outputs(4182)) and not (layer4_outputs(2594));
    layer5_outputs(2547) <= not(layer4_outputs(3478));
    layer5_outputs(2548) <= (layer4_outputs(4579)) and not (layer4_outputs(296));
    layer5_outputs(2549) <= not((layer4_outputs(1176)) xor (layer4_outputs(5289)));
    layer5_outputs(2550) <= (layer4_outputs(2105)) and not (layer4_outputs(282));
    layer5_outputs(2551) <= (layer4_outputs(5915)) and (layer4_outputs(4523));
    layer5_outputs(2552) <= layer4_outputs(6358);
    layer5_outputs(2553) <= not(layer4_outputs(4173));
    layer5_outputs(2554) <= not((layer4_outputs(1704)) xor (layer4_outputs(1258)));
    layer5_outputs(2555) <= not(layer4_outputs(1672)) or (layer4_outputs(4241));
    layer5_outputs(2556) <= layer4_outputs(6954);
    layer5_outputs(2557) <= layer4_outputs(7511);
    layer5_outputs(2558) <= not(layer4_outputs(7379)) or (layer4_outputs(3846));
    layer5_outputs(2559) <= not((layer4_outputs(2835)) and (layer4_outputs(3748)));
    layer5_outputs(2560) <= not((layer4_outputs(2130)) and (layer4_outputs(1140)));
    layer5_outputs(2561) <= layer4_outputs(4713);
    layer5_outputs(2562) <= not(layer4_outputs(766));
    layer5_outputs(2563) <= not(layer4_outputs(5480)) or (layer4_outputs(2350));
    layer5_outputs(2564) <= '0';
    layer5_outputs(2565) <= '0';
    layer5_outputs(2566) <= layer4_outputs(2881);
    layer5_outputs(2567) <= layer4_outputs(2217);
    layer5_outputs(2568) <= not(layer4_outputs(4067));
    layer5_outputs(2569) <= not(layer4_outputs(716)) or (layer4_outputs(5188));
    layer5_outputs(2570) <= (layer4_outputs(2994)) and not (layer4_outputs(5136));
    layer5_outputs(2571) <= not(layer4_outputs(2439));
    layer5_outputs(2572) <= (layer4_outputs(1967)) and not (layer4_outputs(3828));
    layer5_outputs(2573) <= layer4_outputs(2605);
    layer5_outputs(2574) <= layer4_outputs(5281);
    layer5_outputs(2575) <= not(layer4_outputs(2650));
    layer5_outputs(2576) <= (layer4_outputs(860)) and not (layer4_outputs(6482));
    layer5_outputs(2577) <= (layer4_outputs(4411)) xor (layer4_outputs(4152));
    layer5_outputs(2578) <= not((layer4_outputs(4037)) xor (layer4_outputs(5546)));
    layer5_outputs(2579) <= not(layer4_outputs(6059));
    layer5_outputs(2580) <= layer4_outputs(614);
    layer5_outputs(2581) <= (layer4_outputs(889)) and not (layer4_outputs(3481));
    layer5_outputs(2582) <= not(layer4_outputs(6073)) or (layer4_outputs(7084));
    layer5_outputs(2583) <= (layer4_outputs(3015)) and not (layer4_outputs(3415));
    layer5_outputs(2584) <= (layer4_outputs(7469)) and (layer4_outputs(4762));
    layer5_outputs(2585) <= (layer4_outputs(2120)) xor (layer4_outputs(566));
    layer5_outputs(2586) <= layer4_outputs(4493);
    layer5_outputs(2587) <= layer4_outputs(405);
    layer5_outputs(2588) <= not(layer4_outputs(2193));
    layer5_outputs(2589) <= layer4_outputs(1896);
    layer5_outputs(2590) <= layer4_outputs(7434);
    layer5_outputs(2591) <= layer4_outputs(4682);
    layer5_outputs(2592) <= layer4_outputs(3716);
    layer5_outputs(2593) <= (layer4_outputs(1939)) and (layer4_outputs(4216));
    layer5_outputs(2594) <= not(layer4_outputs(309));
    layer5_outputs(2595) <= not((layer4_outputs(1084)) and (layer4_outputs(5895)));
    layer5_outputs(2596) <= not(layer4_outputs(7554)) or (layer4_outputs(1719));
    layer5_outputs(2597) <= layer4_outputs(3604);
    layer5_outputs(2598) <= not(layer4_outputs(6580)) or (layer4_outputs(4574));
    layer5_outputs(2599) <= not(layer4_outputs(6110));
    layer5_outputs(2600) <= (layer4_outputs(2518)) and (layer4_outputs(2749));
    layer5_outputs(2601) <= layer4_outputs(3599);
    layer5_outputs(2602) <= not(layer4_outputs(1277)) or (layer4_outputs(6171));
    layer5_outputs(2603) <= not((layer4_outputs(1186)) or (layer4_outputs(5981)));
    layer5_outputs(2604) <= (layer4_outputs(1741)) xor (layer4_outputs(2363));
    layer5_outputs(2605) <= not(layer4_outputs(7057)) or (layer4_outputs(6503));
    layer5_outputs(2606) <= layer4_outputs(4564);
    layer5_outputs(2607) <= not(layer4_outputs(4857)) or (layer4_outputs(2370));
    layer5_outputs(2608) <= layer4_outputs(1600);
    layer5_outputs(2609) <= (layer4_outputs(6893)) or (layer4_outputs(5093));
    layer5_outputs(2610) <= (layer4_outputs(2599)) or (layer4_outputs(2251));
    layer5_outputs(2611) <= not((layer4_outputs(2696)) or (layer4_outputs(2630)));
    layer5_outputs(2612) <= '0';
    layer5_outputs(2613) <= (layer4_outputs(34)) and (layer4_outputs(4438));
    layer5_outputs(2614) <= (layer4_outputs(7498)) and (layer4_outputs(7132));
    layer5_outputs(2615) <= layer4_outputs(7464);
    layer5_outputs(2616) <= (layer4_outputs(3667)) and (layer4_outputs(4403));
    layer5_outputs(2617) <= layer4_outputs(592);
    layer5_outputs(2618) <= layer4_outputs(6512);
    layer5_outputs(2619) <= not(layer4_outputs(7042));
    layer5_outputs(2620) <= (layer4_outputs(33)) and not (layer4_outputs(4180));
    layer5_outputs(2621) <= (layer4_outputs(7008)) and not (layer4_outputs(2196));
    layer5_outputs(2622) <= (layer4_outputs(5129)) and not (layer4_outputs(1365));
    layer5_outputs(2623) <= not(layer4_outputs(1902));
    layer5_outputs(2624) <= not(layer4_outputs(1670)) or (layer4_outputs(2621));
    layer5_outputs(2625) <= (layer4_outputs(2499)) and not (layer4_outputs(4111));
    layer5_outputs(2626) <= layer4_outputs(6793);
    layer5_outputs(2627) <= not(layer4_outputs(6761));
    layer5_outputs(2628) <= not(layer4_outputs(2429));
    layer5_outputs(2629) <= not(layer4_outputs(916));
    layer5_outputs(2630) <= not(layer4_outputs(6705)) or (layer4_outputs(7517));
    layer5_outputs(2631) <= (layer4_outputs(6934)) and not (layer4_outputs(4001));
    layer5_outputs(2632) <= (layer4_outputs(3137)) and not (layer4_outputs(821));
    layer5_outputs(2633) <= not(layer4_outputs(4402));
    layer5_outputs(2634) <= '0';
    layer5_outputs(2635) <= not(layer4_outputs(1364)) or (layer4_outputs(7146));
    layer5_outputs(2636) <= not((layer4_outputs(5196)) xor (layer4_outputs(5761)));
    layer5_outputs(2637) <= not(layer4_outputs(1702));
    layer5_outputs(2638) <= not(layer4_outputs(135));
    layer5_outputs(2639) <= layer4_outputs(5666);
    layer5_outputs(2640) <= not((layer4_outputs(4457)) xor (layer4_outputs(708)));
    layer5_outputs(2641) <= not(layer4_outputs(2225));
    layer5_outputs(2642) <= not(layer4_outputs(1774));
    layer5_outputs(2643) <= not(layer4_outputs(363));
    layer5_outputs(2644) <= layer4_outputs(204);
    layer5_outputs(2645) <= layer4_outputs(2226);
    layer5_outputs(2646) <= not(layer4_outputs(6831));
    layer5_outputs(2647) <= (layer4_outputs(1646)) and not (layer4_outputs(6039));
    layer5_outputs(2648) <= (layer4_outputs(5468)) xor (layer4_outputs(6125));
    layer5_outputs(2649) <= layer4_outputs(789);
    layer5_outputs(2650) <= layer4_outputs(4862);
    layer5_outputs(2651) <= not(layer4_outputs(5566));
    layer5_outputs(2652) <= not(layer4_outputs(1319));
    layer5_outputs(2653) <= not(layer4_outputs(3837));
    layer5_outputs(2654) <= not(layer4_outputs(1598)) or (layer4_outputs(6898));
    layer5_outputs(2655) <= (layer4_outputs(2424)) xor (layer4_outputs(5875));
    layer5_outputs(2656) <= layer4_outputs(7006);
    layer5_outputs(2657) <= not(layer4_outputs(1694)) or (layer4_outputs(6550));
    layer5_outputs(2658) <= (layer4_outputs(2093)) or (layer4_outputs(2488));
    layer5_outputs(2659) <= not(layer4_outputs(6636));
    layer5_outputs(2660) <= layer4_outputs(3082);
    layer5_outputs(2661) <= not((layer4_outputs(3200)) or (layer4_outputs(7509)));
    layer5_outputs(2662) <= not(layer4_outputs(5423));
    layer5_outputs(2663) <= '0';
    layer5_outputs(2664) <= layer4_outputs(3086);
    layer5_outputs(2665) <= (layer4_outputs(4599)) and not (layer4_outputs(803));
    layer5_outputs(2666) <= not(layer4_outputs(6089));
    layer5_outputs(2667) <= layer4_outputs(5405);
    layer5_outputs(2668) <= not((layer4_outputs(4243)) and (layer4_outputs(2817)));
    layer5_outputs(2669) <= not(layer4_outputs(2253));
    layer5_outputs(2670) <= not((layer4_outputs(1507)) xor (layer4_outputs(3278)));
    layer5_outputs(2671) <= not((layer4_outputs(6072)) or (layer4_outputs(1180)));
    layer5_outputs(2672) <= (layer4_outputs(3260)) xor (layer4_outputs(6621));
    layer5_outputs(2673) <= not(layer4_outputs(1173));
    layer5_outputs(2674) <= (layer4_outputs(7281)) and not (layer4_outputs(5201));
    layer5_outputs(2675) <= not(layer4_outputs(1761));
    layer5_outputs(2676) <= not(layer4_outputs(7076));
    layer5_outputs(2677) <= (layer4_outputs(2278)) and (layer4_outputs(3057));
    layer5_outputs(2678) <= not(layer4_outputs(7494));
    layer5_outputs(2679) <= not(layer4_outputs(2904));
    layer5_outputs(2680) <= layer4_outputs(6479);
    layer5_outputs(2681) <= not(layer4_outputs(4337));
    layer5_outputs(2682) <= (layer4_outputs(2247)) and not (layer4_outputs(954));
    layer5_outputs(2683) <= (layer4_outputs(6223)) or (layer4_outputs(1279));
    layer5_outputs(2684) <= not(layer4_outputs(6855)) or (layer4_outputs(6778));
    layer5_outputs(2685) <= not(layer4_outputs(4818));
    layer5_outputs(2686) <= layer4_outputs(4970);
    layer5_outputs(2687) <= (layer4_outputs(3395)) xor (layer4_outputs(3058));
    layer5_outputs(2688) <= layer4_outputs(2421);
    layer5_outputs(2689) <= (layer4_outputs(6375)) and (layer4_outputs(2292));
    layer5_outputs(2690) <= not((layer4_outputs(2911)) xor (layer4_outputs(1004)));
    layer5_outputs(2691) <= not(layer4_outputs(2619)) or (layer4_outputs(7535));
    layer5_outputs(2692) <= not(layer4_outputs(535));
    layer5_outputs(2693) <= (layer4_outputs(2844)) xor (layer4_outputs(408));
    layer5_outputs(2694) <= layer4_outputs(3976);
    layer5_outputs(2695) <= not(layer4_outputs(7086));
    layer5_outputs(2696) <= (layer4_outputs(6724)) and (layer4_outputs(3104));
    layer5_outputs(2697) <= layer4_outputs(5837);
    layer5_outputs(2698) <= not((layer4_outputs(726)) or (layer4_outputs(1031)));
    layer5_outputs(2699) <= (layer4_outputs(838)) and not (layer4_outputs(1840));
    layer5_outputs(2700) <= layer4_outputs(6022);
    layer5_outputs(2701) <= not(layer4_outputs(7214));
    layer5_outputs(2702) <= '0';
    layer5_outputs(2703) <= not(layer4_outputs(2481));
    layer5_outputs(2704) <= layer4_outputs(3070);
    layer5_outputs(2705) <= (layer4_outputs(2993)) or (layer4_outputs(4854));
    layer5_outputs(2706) <= layer4_outputs(40);
    layer5_outputs(2707) <= not(layer4_outputs(1083));
    layer5_outputs(2708) <= (layer4_outputs(1250)) and (layer4_outputs(3045));
    layer5_outputs(2709) <= layer4_outputs(6586);
    layer5_outputs(2710) <= not(layer4_outputs(2987));
    layer5_outputs(2711) <= (layer4_outputs(2495)) or (layer4_outputs(212));
    layer5_outputs(2712) <= not((layer4_outputs(2138)) xor (layer4_outputs(5834)));
    layer5_outputs(2713) <= not(layer4_outputs(5647));
    layer5_outputs(2714) <= (layer4_outputs(5020)) or (layer4_outputs(5573));
    layer5_outputs(2715) <= layer4_outputs(309);
    layer5_outputs(2716) <= (layer4_outputs(6276)) and (layer4_outputs(4155));
    layer5_outputs(2717) <= not((layer4_outputs(7145)) xor (layer4_outputs(1826)));
    layer5_outputs(2718) <= (layer4_outputs(6808)) xor (layer4_outputs(2086));
    layer5_outputs(2719) <= not(layer4_outputs(5043));
    layer5_outputs(2720) <= layer4_outputs(5145);
    layer5_outputs(2721) <= (layer4_outputs(4828)) and not (layer4_outputs(1301));
    layer5_outputs(2722) <= not((layer4_outputs(867)) and (layer4_outputs(941)));
    layer5_outputs(2723) <= not(layer4_outputs(6131));
    layer5_outputs(2724) <= not(layer4_outputs(2371));
    layer5_outputs(2725) <= layer4_outputs(1474);
    layer5_outputs(2726) <= '1';
    layer5_outputs(2727) <= (layer4_outputs(1384)) and not (layer4_outputs(7672));
    layer5_outputs(2728) <= not(layer4_outputs(1275));
    layer5_outputs(2729) <= not(layer4_outputs(3360));
    layer5_outputs(2730) <= (layer4_outputs(1477)) and not (layer4_outputs(5176));
    layer5_outputs(2731) <= not(layer4_outputs(4825)) or (layer4_outputs(3926));
    layer5_outputs(2732) <= not(layer4_outputs(6747));
    layer5_outputs(2733) <= not((layer4_outputs(1012)) xor (layer4_outputs(5401)));
    layer5_outputs(2734) <= not((layer4_outputs(5312)) xor (layer4_outputs(5726)));
    layer5_outputs(2735) <= not(layer4_outputs(3937));
    layer5_outputs(2736) <= not((layer4_outputs(5381)) and (layer4_outputs(2591)));
    layer5_outputs(2737) <= layer4_outputs(7315);
    layer5_outputs(2738) <= layer4_outputs(5576);
    layer5_outputs(2739) <= layer4_outputs(3293);
    layer5_outputs(2740) <= not((layer4_outputs(1638)) or (layer4_outputs(406)));
    layer5_outputs(2741) <= (layer4_outputs(1865)) or (layer4_outputs(2675));
    layer5_outputs(2742) <= (layer4_outputs(6841)) xor (layer4_outputs(2976));
    layer5_outputs(2743) <= layer4_outputs(6878);
    layer5_outputs(2744) <= layer4_outputs(4780);
    layer5_outputs(2745) <= layer4_outputs(5785);
    layer5_outputs(2746) <= not(layer4_outputs(3284));
    layer5_outputs(2747) <= not(layer4_outputs(2433)) or (layer4_outputs(201));
    layer5_outputs(2748) <= not(layer4_outputs(2668));
    layer5_outputs(2749) <= not(layer4_outputs(326)) or (layer4_outputs(7260));
    layer5_outputs(2750) <= '0';
    layer5_outputs(2751) <= layer4_outputs(3744);
    layer5_outputs(2752) <= not(layer4_outputs(7290)) or (layer4_outputs(951));
    layer5_outputs(2753) <= layer4_outputs(3404);
    layer5_outputs(2754) <= layer4_outputs(2035);
    layer5_outputs(2755) <= (layer4_outputs(2527)) and not (layer4_outputs(1170));
    layer5_outputs(2756) <= layer4_outputs(6638);
    layer5_outputs(2757) <= not(layer4_outputs(7269));
    layer5_outputs(2758) <= not(layer4_outputs(713));
    layer5_outputs(2759) <= (layer4_outputs(4445)) and (layer4_outputs(6838));
    layer5_outputs(2760) <= not(layer4_outputs(5453));
    layer5_outputs(2761) <= not(layer4_outputs(915));
    layer5_outputs(2762) <= (layer4_outputs(1865)) and not (layer4_outputs(1962));
    layer5_outputs(2763) <= not(layer4_outputs(2392)) or (layer4_outputs(4561));
    layer5_outputs(2764) <= not((layer4_outputs(6058)) and (layer4_outputs(1725)));
    layer5_outputs(2765) <= layer4_outputs(3348);
    layer5_outputs(2766) <= layer4_outputs(904);
    layer5_outputs(2767) <= '1';
    layer5_outputs(2768) <= layer4_outputs(3353);
    layer5_outputs(2769) <= not(layer4_outputs(5936)) or (layer4_outputs(3489));
    layer5_outputs(2770) <= (layer4_outputs(1860)) or (layer4_outputs(1510));
    layer5_outputs(2771) <= not(layer4_outputs(3767)) or (layer4_outputs(1249));
    layer5_outputs(2772) <= layer4_outputs(1804);
    layer5_outputs(2773) <= not((layer4_outputs(2886)) xor (layer4_outputs(5951)));
    layer5_outputs(2774) <= (layer4_outputs(2006)) or (layer4_outputs(5365));
    layer5_outputs(2775) <= (layer4_outputs(2343)) xor (layer4_outputs(1338));
    layer5_outputs(2776) <= layer4_outputs(2863);
    layer5_outputs(2777) <= layer4_outputs(5263);
    layer5_outputs(2778) <= (layer4_outputs(1384)) and not (layer4_outputs(2780));
    layer5_outputs(2779) <= not(layer4_outputs(326));
    layer5_outputs(2780) <= (layer4_outputs(6877)) and not (layer4_outputs(950));
    layer5_outputs(2781) <= not(layer4_outputs(6122));
    layer5_outputs(2782) <= not(layer4_outputs(899)) or (layer4_outputs(6029));
    layer5_outputs(2783) <= not(layer4_outputs(4543));
    layer5_outputs(2784) <= not(layer4_outputs(3075));
    layer5_outputs(2785) <= not(layer4_outputs(4306));
    layer5_outputs(2786) <= not(layer4_outputs(3619));
    layer5_outputs(2787) <= not(layer4_outputs(3364));
    layer5_outputs(2788) <= layer4_outputs(6964);
    layer5_outputs(2789) <= not((layer4_outputs(2280)) or (layer4_outputs(3157)));
    layer5_outputs(2790) <= not((layer4_outputs(4200)) and (layer4_outputs(6395)));
    layer5_outputs(2791) <= (layer4_outputs(4638)) or (layer4_outputs(6739));
    layer5_outputs(2792) <= (layer4_outputs(7640)) and not (layer4_outputs(6208));
    layer5_outputs(2793) <= not((layer4_outputs(6885)) and (layer4_outputs(5455)));
    layer5_outputs(2794) <= not(layer4_outputs(1784));
    layer5_outputs(2795) <= not(layer4_outputs(3153));
    layer5_outputs(2796) <= layer4_outputs(6946);
    layer5_outputs(2797) <= not(layer4_outputs(6471));
    layer5_outputs(2798) <= layer4_outputs(7569);
    layer5_outputs(2799) <= not((layer4_outputs(4589)) xor (layer4_outputs(6273)));
    layer5_outputs(2800) <= layer4_outputs(2864);
    layer5_outputs(2801) <= (layer4_outputs(4215)) and (layer4_outputs(5336));
    layer5_outputs(2802) <= layer4_outputs(7064);
    layer5_outputs(2803) <= (layer4_outputs(6694)) and (layer4_outputs(6802));
    layer5_outputs(2804) <= layer4_outputs(4292);
    layer5_outputs(2805) <= not(layer4_outputs(4449));
    layer5_outputs(2806) <= not((layer4_outputs(7191)) and (layer4_outputs(6135)));
    layer5_outputs(2807) <= '1';
    layer5_outputs(2808) <= not(layer4_outputs(1119));
    layer5_outputs(2809) <= layer4_outputs(1139);
    layer5_outputs(2810) <= layer4_outputs(4582);
    layer5_outputs(2811) <= not(layer4_outputs(3388));
    layer5_outputs(2812) <= not(layer4_outputs(1752));
    layer5_outputs(2813) <= layer4_outputs(1766);
    layer5_outputs(2814) <= (layer4_outputs(2017)) xor (layer4_outputs(2583));
    layer5_outputs(2815) <= (layer4_outputs(2656)) or (layer4_outputs(5753));
    layer5_outputs(2816) <= not(layer4_outputs(4408));
    layer5_outputs(2817) <= (layer4_outputs(6037)) and not (layer4_outputs(2805));
    layer5_outputs(2818) <= not(layer4_outputs(3042));
    layer5_outputs(2819) <= (layer4_outputs(5998)) or (layer4_outputs(2460));
    layer5_outputs(2820) <= layer4_outputs(6211);
    layer5_outputs(2821) <= not((layer4_outputs(832)) xor (layer4_outputs(7306)));
    layer5_outputs(2822) <= not(layer4_outputs(266));
    layer5_outputs(2823) <= (layer4_outputs(4520)) xor (layer4_outputs(1530));
    layer5_outputs(2824) <= not((layer4_outputs(7422)) xor (layer4_outputs(3659)));
    layer5_outputs(2825) <= layer4_outputs(1669);
    layer5_outputs(2826) <= layer4_outputs(345);
    layer5_outputs(2827) <= layer4_outputs(4124);
    layer5_outputs(2828) <= (layer4_outputs(1125)) or (layer4_outputs(1668));
    layer5_outputs(2829) <= layer4_outputs(4645);
    layer5_outputs(2830) <= (layer4_outputs(5782)) and not (layer4_outputs(6205));
    layer5_outputs(2831) <= not(layer4_outputs(7196)) or (layer4_outputs(7110));
    layer5_outputs(2832) <= not(layer4_outputs(7114));
    layer5_outputs(2833) <= not(layer4_outputs(5758));
    layer5_outputs(2834) <= not(layer4_outputs(5052));
    layer5_outputs(2835) <= (layer4_outputs(760)) and (layer4_outputs(4028));
    layer5_outputs(2836) <= not((layer4_outputs(4344)) xor (layer4_outputs(1242)));
    layer5_outputs(2837) <= not(layer4_outputs(6073));
    layer5_outputs(2838) <= (layer4_outputs(4555)) and (layer4_outputs(5327));
    layer5_outputs(2839) <= (layer4_outputs(4155)) or (layer4_outputs(6488));
    layer5_outputs(2840) <= layer4_outputs(6902);
    layer5_outputs(2841) <= layer4_outputs(328);
    layer5_outputs(2842) <= (layer4_outputs(317)) xor (layer4_outputs(2649));
    layer5_outputs(2843) <= (layer4_outputs(5154)) and not (layer4_outputs(7001));
    layer5_outputs(2844) <= not((layer4_outputs(884)) or (layer4_outputs(5146)));
    layer5_outputs(2845) <= (layer4_outputs(3457)) or (layer4_outputs(1156));
    layer5_outputs(2846) <= layer4_outputs(1749);
    layer5_outputs(2847) <= layer4_outputs(6414);
    layer5_outputs(2848) <= not(layer4_outputs(5234));
    layer5_outputs(2849) <= layer4_outputs(5321);
    layer5_outputs(2850) <= (layer4_outputs(29)) xor (layer4_outputs(7610));
    layer5_outputs(2851) <= not(layer4_outputs(90)) or (layer4_outputs(7166));
    layer5_outputs(2852) <= layer4_outputs(4442);
    layer5_outputs(2853) <= layer4_outputs(1093);
    layer5_outputs(2854) <= layer4_outputs(3720);
    layer5_outputs(2855) <= not((layer4_outputs(7188)) and (layer4_outputs(696)));
    layer5_outputs(2856) <= layer4_outputs(3443);
    layer5_outputs(2857) <= layer4_outputs(5131);
    layer5_outputs(2858) <= not((layer4_outputs(60)) xor (layer4_outputs(7382)));
    layer5_outputs(2859) <= not(layer4_outputs(312));
    layer5_outputs(2860) <= layer4_outputs(4980);
    layer5_outputs(2861) <= (layer4_outputs(4929)) or (layer4_outputs(7360));
    layer5_outputs(2862) <= layer4_outputs(1306);
    layer5_outputs(2863) <= layer4_outputs(4918);
    layer5_outputs(2864) <= (layer4_outputs(7667)) and (layer4_outputs(4181));
    layer5_outputs(2865) <= not(layer4_outputs(3534));
    layer5_outputs(2866) <= not(layer4_outputs(1487));
    layer5_outputs(2867) <= not(layer4_outputs(3907));
    layer5_outputs(2868) <= layer4_outputs(6650);
    layer5_outputs(2869) <= layer4_outputs(5334);
    layer5_outputs(2870) <= not(layer4_outputs(1080));
    layer5_outputs(2871) <= not((layer4_outputs(2355)) xor (layer4_outputs(5494)));
    layer5_outputs(2872) <= layer4_outputs(7430);
    layer5_outputs(2873) <= (layer4_outputs(1935)) and (layer4_outputs(3980));
    layer5_outputs(2874) <= not((layer4_outputs(723)) or (layer4_outputs(98)));
    layer5_outputs(2875) <= not(layer4_outputs(1485));
    layer5_outputs(2876) <= not(layer4_outputs(6480));
    layer5_outputs(2877) <= (layer4_outputs(7211)) and not (layer4_outputs(4942));
    layer5_outputs(2878) <= not(layer4_outputs(6651));
    layer5_outputs(2879) <= not((layer4_outputs(1704)) or (layer4_outputs(3326)));
    layer5_outputs(2880) <= layer4_outputs(1921);
    layer5_outputs(2881) <= (layer4_outputs(4290)) xor (layer4_outputs(5167));
    layer5_outputs(2882) <= not(layer4_outputs(1867));
    layer5_outputs(2883) <= not((layer4_outputs(305)) xor (layer4_outputs(6870)));
    layer5_outputs(2884) <= (layer4_outputs(3605)) or (layer4_outputs(542));
    layer5_outputs(2885) <= not((layer4_outputs(1006)) and (layer4_outputs(4451)));
    layer5_outputs(2886) <= (layer4_outputs(6654)) and (layer4_outputs(5092));
    layer5_outputs(2887) <= not(layer4_outputs(2849));
    layer5_outputs(2888) <= (layer4_outputs(4465)) xor (layer4_outputs(2294));
    layer5_outputs(2889) <= (layer4_outputs(5971)) or (layer4_outputs(1462));
    layer5_outputs(2890) <= not(layer4_outputs(3662));
    layer5_outputs(2891) <= not((layer4_outputs(6361)) or (layer4_outputs(4046)));
    layer5_outputs(2892) <= (layer4_outputs(2170)) and (layer4_outputs(2187));
    layer5_outputs(2893) <= layer4_outputs(2332);
    layer5_outputs(2894) <= layer4_outputs(6248);
    layer5_outputs(2895) <= not(layer4_outputs(6009));
    layer5_outputs(2896) <= (layer4_outputs(6999)) and not (layer4_outputs(2326));
    layer5_outputs(2897) <= not((layer4_outputs(704)) xor (layer4_outputs(4341)));
    layer5_outputs(2898) <= (layer4_outputs(5386)) xor (layer4_outputs(4930));
    layer5_outputs(2899) <= layer4_outputs(6252);
    layer5_outputs(2900) <= not((layer4_outputs(4136)) or (layer4_outputs(3581)));
    layer5_outputs(2901) <= not(layer4_outputs(6586)) or (layer4_outputs(6377));
    layer5_outputs(2902) <= layer4_outputs(3308);
    layer5_outputs(2903) <= layer4_outputs(2084);
    layer5_outputs(2904) <= not((layer4_outputs(5435)) xor (layer4_outputs(7500)));
    layer5_outputs(2905) <= not((layer4_outputs(3756)) xor (layer4_outputs(7066)));
    layer5_outputs(2906) <= not((layer4_outputs(7333)) and (layer4_outputs(4819)));
    layer5_outputs(2907) <= not(layer4_outputs(6225));
    layer5_outputs(2908) <= not(layer4_outputs(4872));
    layer5_outputs(2909) <= '1';
    layer5_outputs(2910) <= (layer4_outputs(5253)) xor (layer4_outputs(4472));
    layer5_outputs(2911) <= not(layer4_outputs(3127)) or (layer4_outputs(1900));
    layer5_outputs(2912) <= not(layer4_outputs(547));
    layer5_outputs(2913) <= not(layer4_outputs(235));
    layer5_outputs(2914) <= not(layer4_outputs(5383));
    layer5_outputs(2915) <= (layer4_outputs(1145)) and not (layer4_outputs(4984));
    layer5_outputs(2916) <= not(layer4_outputs(6607)) or (layer4_outputs(7363));
    layer5_outputs(2917) <= (layer4_outputs(6279)) and not (layer4_outputs(6992));
    layer5_outputs(2918) <= not((layer4_outputs(57)) and (layer4_outputs(191)));
    layer5_outputs(2919) <= not((layer4_outputs(667)) xor (layer4_outputs(1506)));
    layer5_outputs(2920) <= layer4_outputs(7012);
    layer5_outputs(2921) <= not(layer4_outputs(5955));
    layer5_outputs(2922) <= not(layer4_outputs(5737));
    layer5_outputs(2923) <= not((layer4_outputs(799)) or (layer4_outputs(2466)));
    layer5_outputs(2924) <= layer4_outputs(386);
    layer5_outputs(2925) <= (layer4_outputs(3797)) and (layer4_outputs(985));
    layer5_outputs(2926) <= layer4_outputs(1753);
    layer5_outputs(2927) <= not((layer4_outputs(6406)) or (layer4_outputs(2291)));
    layer5_outputs(2928) <= not(layer4_outputs(3291));
    layer5_outputs(2929) <= not((layer4_outputs(7250)) and (layer4_outputs(2085)));
    layer5_outputs(2930) <= layer4_outputs(3686);
    layer5_outputs(2931) <= not(layer4_outputs(3459));
    layer5_outputs(2932) <= layer4_outputs(6562);
    layer5_outputs(2933) <= (layer4_outputs(4131)) xor (layer4_outputs(6211));
    layer5_outputs(2934) <= (layer4_outputs(123)) or (layer4_outputs(4372));
    layer5_outputs(2935) <= not(layer4_outputs(3188));
    layer5_outputs(2936) <= not(layer4_outputs(4191));
    layer5_outputs(2937) <= layer4_outputs(7388);
    layer5_outputs(2938) <= (layer4_outputs(5316)) or (layer4_outputs(3675));
    layer5_outputs(2939) <= layer4_outputs(4629);
    layer5_outputs(2940) <= (layer4_outputs(1579)) and not (layer4_outputs(3347));
    layer5_outputs(2941) <= not(layer4_outputs(6191));
    layer5_outputs(2942) <= not(layer4_outputs(3787));
    layer5_outputs(2943) <= (layer4_outputs(7416)) and not (layer4_outputs(241));
    layer5_outputs(2944) <= (layer4_outputs(4833)) and not (layer4_outputs(3968));
    layer5_outputs(2945) <= not(layer4_outputs(4362)) or (layer4_outputs(3639));
    layer5_outputs(2946) <= not((layer4_outputs(2842)) or (layer4_outputs(6756)));
    layer5_outputs(2947) <= not(layer4_outputs(3892)) or (layer4_outputs(4446));
    layer5_outputs(2948) <= layer4_outputs(5382);
    layer5_outputs(2949) <= (layer4_outputs(791)) and (layer4_outputs(4632));
    layer5_outputs(2950) <= not(layer4_outputs(1612)) or (layer4_outputs(6496));
    layer5_outputs(2951) <= not((layer4_outputs(4261)) xor (layer4_outputs(1422)));
    layer5_outputs(2952) <= not(layer4_outputs(292));
    layer5_outputs(2953) <= not((layer4_outputs(6316)) or (layer4_outputs(1930)));
    layer5_outputs(2954) <= (layer4_outputs(4162)) and not (layer4_outputs(3986));
    layer5_outputs(2955) <= not(layer4_outputs(2004));
    layer5_outputs(2956) <= not((layer4_outputs(3541)) xor (layer4_outputs(5332)));
    layer5_outputs(2957) <= not(layer4_outputs(565));
    layer5_outputs(2958) <= not(layer4_outputs(3895));
    layer5_outputs(2959) <= (layer4_outputs(2916)) and (layer4_outputs(943));
    layer5_outputs(2960) <= not((layer4_outputs(1331)) xor (layer4_outputs(4752)));
    layer5_outputs(2961) <= not(layer4_outputs(3856));
    layer5_outputs(2962) <= layer4_outputs(3464);
    layer5_outputs(2963) <= layer4_outputs(5559);
    layer5_outputs(2964) <= (layer4_outputs(2851)) and not (layer4_outputs(5094));
    layer5_outputs(2965) <= layer4_outputs(3710);
    layer5_outputs(2966) <= (layer4_outputs(5632)) and not (layer4_outputs(6663));
    layer5_outputs(2967) <= not(layer4_outputs(5960));
    layer5_outputs(2968) <= (layer4_outputs(2462)) xor (layer4_outputs(3742));
    layer5_outputs(2969) <= not(layer4_outputs(5670));
    layer5_outputs(2970) <= not(layer4_outputs(7557));
    layer5_outputs(2971) <= not(layer4_outputs(4072));
    layer5_outputs(2972) <= layer4_outputs(2062);
    layer5_outputs(2973) <= not(layer4_outputs(3265));
    layer5_outputs(2974) <= not(layer4_outputs(3809)) or (layer4_outputs(7099));
    layer5_outputs(2975) <= '1';
    layer5_outputs(2976) <= layer4_outputs(192);
    layer5_outputs(2977) <= not(layer4_outputs(5677)) or (layer4_outputs(2335));
    layer5_outputs(2978) <= not(layer4_outputs(6811));
    layer5_outputs(2979) <= (layer4_outputs(5175)) and not (layer4_outputs(4581));
    layer5_outputs(2980) <= layer4_outputs(2552);
    layer5_outputs(2981) <= not(layer4_outputs(5687));
    layer5_outputs(2982) <= not(layer4_outputs(2127));
    layer5_outputs(2983) <= (layer4_outputs(1929)) and not (layer4_outputs(1020));
    layer5_outputs(2984) <= (layer4_outputs(4551)) and not (layer4_outputs(1049));
    layer5_outputs(2985) <= not((layer4_outputs(5232)) xor (layer4_outputs(246)));
    layer5_outputs(2986) <= (layer4_outputs(2998)) and (layer4_outputs(4151));
    layer5_outputs(2987) <= not(layer4_outputs(2122));
    layer5_outputs(2988) <= not(layer4_outputs(1366));
    layer5_outputs(2989) <= (layer4_outputs(3944)) and (layer4_outputs(4389));
    layer5_outputs(2990) <= (layer4_outputs(4941)) and (layer4_outputs(5308));
    layer5_outputs(2991) <= not(layer4_outputs(5406));
    layer5_outputs(2992) <= not((layer4_outputs(2087)) and (layer4_outputs(1214)));
    layer5_outputs(2993) <= layer4_outputs(5358);
    layer5_outputs(2994) <= not(layer4_outputs(1552));
    layer5_outputs(2995) <= layer4_outputs(6439);
    layer5_outputs(2996) <= layer4_outputs(4051);
    layer5_outputs(2997) <= layer4_outputs(2065);
    layer5_outputs(2998) <= not(layer4_outputs(5338));
    layer5_outputs(2999) <= layer4_outputs(2150);
    layer5_outputs(3000) <= not((layer4_outputs(474)) or (layer4_outputs(3488)));
    layer5_outputs(3001) <= not(layer4_outputs(819)) or (layer4_outputs(4658));
    layer5_outputs(3002) <= not(layer4_outputs(4880));
    layer5_outputs(3003) <= '0';
    layer5_outputs(3004) <= (layer4_outputs(749)) or (layer4_outputs(600));
    layer5_outputs(3005) <= not(layer4_outputs(2318));
    layer5_outputs(3006) <= layer4_outputs(1593);
    layer5_outputs(3007) <= (layer4_outputs(868)) xor (layer4_outputs(5752));
    layer5_outputs(3008) <= not(layer4_outputs(5438));
    layer5_outputs(3009) <= not(layer4_outputs(6879));
    layer5_outputs(3010) <= not(layer4_outputs(6602));
    layer5_outputs(3011) <= not(layer4_outputs(3623));
    layer5_outputs(3012) <= (layer4_outputs(262)) or (layer4_outputs(4020));
    layer5_outputs(3013) <= not((layer4_outputs(55)) xor (layer4_outputs(5734)));
    layer5_outputs(3014) <= not((layer4_outputs(3141)) xor (layer4_outputs(7350)));
    layer5_outputs(3015) <= not(layer4_outputs(2039)) or (layer4_outputs(5615));
    layer5_outputs(3016) <= not(layer4_outputs(7647));
    layer5_outputs(3017) <= not(layer4_outputs(5501)) or (layer4_outputs(2399));
    layer5_outputs(3018) <= '0';
    layer5_outputs(3019) <= (layer4_outputs(67)) and not (layer4_outputs(7346));
    layer5_outputs(3020) <= not(layer4_outputs(1839));
    layer5_outputs(3021) <= not(layer4_outputs(7053));
    layer5_outputs(3022) <= (layer4_outputs(929)) xor (layer4_outputs(7103));
    layer5_outputs(3023) <= layer4_outputs(2302);
    layer5_outputs(3024) <= not(layer4_outputs(6288)) or (layer4_outputs(5407));
    layer5_outputs(3025) <= layer4_outputs(6638);
    layer5_outputs(3026) <= layer4_outputs(3229);
    layer5_outputs(3027) <= not(layer4_outputs(5365));
    layer5_outputs(3028) <= layer4_outputs(6281);
    layer5_outputs(3029) <= not(layer4_outputs(7146));
    layer5_outputs(3030) <= not((layer4_outputs(2650)) and (layer4_outputs(1673)));
    layer5_outputs(3031) <= (layer4_outputs(3844)) xor (layer4_outputs(4483));
    layer5_outputs(3032) <= layer4_outputs(2240);
    layer5_outputs(3033) <= not(layer4_outputs(2676));
    layer5_outputs(3034) <= layer4_outputs(2190);
    layer5_outputs(3035) <= (layer4_outputs(3715)) or (layer4_outputs(7364));
    layer5_outputs(3036) <= not((layer4_outputs(3375)) and (layer4_outputs(4035)));
    layer5_outputs(3037) <= not(layer4_outputs(3311));
    layer5_outputs(3038) <= not(layer4_outputs(942));
    layer5_outputs(3039) <= layer4_outputs(151);
    layer5_outputs(3040) <= layer4_outputs(5120);
    layer5_outputs(3041) <= not(layer4_outputs(5157));
    layer5_outputs(3042) <= not(layer4_outputs(2893));
    layer5_outputs(3043) <= (layer4_outputs(5715)) and (layer4_outputs(4793));
    layer5_outputs(3044) <= layer4_outputs(5229);
    layer5_outputs(3045) <= not(layer4_outputs(1914)) or (layer4_outputs(5063));
    layer5_outputs(3046) <= '0';
    layer5_outputs(3047) <= layer4_outputs(4416);
    layer5_outputs(3048) <= layer4_outputs(7482);
    layer5_outputs(3049) <= not((layer4_outputs(5547)) or (layer4_outputs(3501)));
    layer5_outputs(3050) <= not((layer4_outputs(4072)) or (layer4_outputs(5159)));
    layer5_outputs(3051) <= layer4_outputs(7549);
    layer5_outputs(3052) <= not(layer4_outputs(7489));
    layer5_outputs(3053) <= layer4_outputs(1639);
    layer5_outputs(3054) <= not(layer4_outputs(3672)) or (layer4_outputs(1120));
    layer5_outputs(3055) <= not((layer4_outputs(3537)) and (layer4_outputs(434)));
    layer5_outputs(3056) <= not(layer4_outputs(1335)) or (layer4_outputs(6268));
    layer5_outputs(3057) <= layer4_outputs(922);
    layer5_outputs(3058) <= not(layer4_outputs(4225));
    layer5_outputs(3059) <= not(layer4_outputs(5743)) or (layer4_outputs(2666));
    layer5_outputs(3060) <= (layer4_outputs(1108)) and not (layer4_outputs(4422));
    layer5_outputs(3061) <= not(layer4_outputs(218));
    layer5_outputs(3062) <= not(layer4_outputs(1870));
    layer5_outputs(3063) <= not((layer4_outputs(2088)) xor (layer4_outputs(4988)));
    layer5_outputs(3064) <= (layer4_outputs(2921)) and not (layer4_outputs(6126));
    layer5_outputs(3065) <= not((layer4_outputs(7497)) and (layer4_outputs(5686)));
    layer5_outputs(3066) <= (layer4_outputs(3319)) xor (layer4_outputs(3654));
    layer5_outputs(3067) <= layer4_outputs(1809);
    layer5_outputs(3068) <= layer4_outputs(1271);
    layer5_outputs(3069) <= layer4_outputs(2873);
    layer5_outputs(3070) <= not((layer4_outputs(1484)) and (layer4_outputs(5036)));
    layer5_outputs(3071) <= not(layer4_outputs(1991));
    layer5_outputs(3072) <= not(layer4_outputs(681));
    layer5_outputs(3073) <= not((layer4_outputs(2821)) xor (layer4_outputs(6595)));
    layer5_outputs(3074) <= (layer4_outputs(7580)) and not (layer4_outputs(5274));
    layer5_outputs(3075) <= not(layer4_outputs(4164));
    layer5_outputs(3076) <= (layer4_outputs(3436)) and not (layer4_outputs(6631));
    layer5_outputs(3077) <= not((layer4_outputs(4331)) and (layer4_outputs(722)));
    layer5_outputs(3078) <= layer4_outputs(2631);
    layer5_outputs(3079) <= not((layer4_outputs(3896)) and (layer4_outputs(1425)));
    layer5_outputs(3080) <= layer4_outputs(2228);
    layer5_outputs(3081) <= not(layer4_outputs(2772));
    layer5_outputs(3082) <= not((layer4_outputs(3465)) and (layer4_outputs(2690)));
    layer5_outputs(3083) <= not(layer4_outputs(5266));
    layer5_outputs(3084) <= layer4_outputs(3062);
    layer5_outputs(3085) <= '0';
    layer5_outputs(3086) <= (layer4_outputs(1357)) xor (layer4_outputs(3925));
    layer5_outputs(3087) <= not(layer4_outputs(7038));
    layer5_outputs(3088) <= (layer4_outputs(2929)) and not (layer4_outputs(3175));
    layer5_outputs(3089) <= not((layer4_outputs(2562)) or (layer4_outputs(7242)));
    layer5_outputs(3090) <= (layer4_outputs(1505)) xor (layer4_outputs(7149));
    layer5_outputs(3091) <= (layer4_outputs(7346)) xor (layer4_outputs(4073));
    layer5_outputs(3092) <= not(layer4_outputs(4900));
    layer5_outputs(3093) <= '0';
    layer5_outputs(3094) <= not(layer4_outputs(5306));
    layer5_outputs(3095) <= (layer4_outputs(7476)) and not (layer4_outputs(5661));
    layer5_outputs(3096) <= not(layer4_outputs(5242)) or (layer4_outputs(21));
    layer5_outputs(3097) <= not((layer4_outputs(1082)) and (layer4_outputs(3177)));
    layer5_outputs(3098) <= not(layer4_outputs(1138));
    layer5_outputs(3099) <= not(layer4_outputs(736));
    layer5_outputs(3100) <= not((layer4_outputs(2402)) or (layer4_outputs(1393)));
    layer5_outputs(3101) <= not(layer4_outputs(6713));
    layer5_outputs(3102) <= layer4_outputs(5117);
    layer5_outputs(3103) <= layer4_outputs(1379);
    layer5_outputs(3104) <= (layer4_outputs(1941)) or (layer4_outputs(1490));
    layer5_outputs(3105) <= not(layer4_outputs(7565));
    layer5_outputs(3106) <= not((layer4_outputs(7170)) or (layer4_outputs(5475)));
    layer5_outputs(3107) <= layer4_outputs(892);
    layer5_outputs(3108) <= '0';
    layer5_outputs(3109) <= not(layer4_outputs(2993));
    layer5_outputs(3110) <= '1';
    layer5_outputs(3111) <= not((layer4_outputs(1943)) xor (layer4_outputs(2610)));
    layer5_outputs(3112) <= (layer4_outputs(4989)) and (layer4_outputs(1861));
    layer5_outputs(3113) <= (layer4_outputs(3052)) and not (layer4_outputs(1130));
    layer5_outputs(3114) <= layer4_outputs(1454);
    layer5_outputs(3115) <= not((layer4_outputs(3865)) and (layer4_outputs(186)));
    layer5_outputs(3116) <= (layer4_outputs(1837)) or (layer4_outputs(6919));
    layer5_outputs(3117) <= (layer4_outputs(3179)) and (layer4_outputs(2431));
    layer5_outputs(3118) <= (layer4_outputs(6810)) and not (layer4_outputs(7272));
    layer5_outputs(3119) <= '1';
    layer5_outputs(3120) <= layer4_outputs(4527);
    layer5_outputs(3121) <= layer4_outputs(6588);
    layer5_outputs(3122) <= not((layer4_outputs(5516)) xor (layer4_outputs(1143)));
    layer5_outputs(3123) <= not(layer4_outputs(7226));
    layer5_outputs(3124) <= not((layer4_outputs(501)) and (layer4_outputs(5921)));
    layer5_outputs(3125) <= not(layer4_outputs(2549));
    layer5_outputs(3126) <= layer4_outputs(5837);
    layer5_outputs(3127) <= (layer4_outputs(6948)) and (layer4_outputs(2899));
    layer5_outputs(3128) <= (layer4_outputs(6536)) and (layer4_outputs(855));
    layer5_outputs(3129) <= not(layer4_outputs(1449));
    layer5_outputs(3130) <= not(layer4_outputs(6419)) or (layer4_outputs(4815));
    layer5_outputs(3131) <= (layer4_outputs(6265)) or (layer4_outputs(6622));
    layer5_outputs(3132) <= (layer4_outputs(6942)) or (layer4_outputs(2317));
    layer5_outputs(3133) <= layer4_outputs(6448);
    layer5_outputs(3134) <= layer4_outputs(4103);
    layer5_outputs(3135) <= not(layer4_outputs(2242)) or (layer4_outputs(3782));
    layer5_outputs(3136) <= layer4_outputs(1678);
    layer5_outputs(3137) <= not(layer4_outputs(7417));
    layer5_outputs(3138) <= not((layer4_outputs(666)) and (layer4_outputs(116)));
    layer5_outputs(3139) <= (layer4_outputs(5374)) xor (layer4_outputs(3784));
    layer5_outputs(3140) <= layer4_outputs(4968);
    layer5_outputs(3141) <= not(layer4_outputs(4926));
    layer5_outputs(3142) <= (layer4_outputs(2244)) and not (layer4_outputs(3707));
    layer5_outputs(3143) <= not(layer4_outputs(271));
    layer5_outputs(3144) <= (layer4_outputs(3853)) and not (layer4_outputs(3642));
    layer5_outputs(3145) <= layer4_outputs(6227);
    layer5_outputs(3146) <= not(layer4_outputs(365));
    layer5_outputs(3147) <= not((layer4_outputs(718)) xor (layer4_outputs(1633)));
    layer5_outputs(3148) <= not((layer4_outputs(983)) and (layer4_outputs(6828)));
    layer5_outputs(3149) <= (layer4_outputs(4326)) and not (layer4_outputs(2784));
    layer5_outputs(3150) <= not(layer4_outputs(250)) or (layer4_outputs(446));
    layer5_outputs(3151) <= not(layer4_outputs(5922)) or (layer4_outputs(4096));
    layer5_outputs(3152) <= not(layer4_outputs(5206)) or (layer4_outputs(3094));
    layer5_outputs(3153) <= layer4_outputs(7652);
    layer5_outputs(3154) <= not((layer4_outputs(6716)) xor (layer4_outputs(7445)));
    layer5_outputs(3155) <= not(layer4_outputs(4307));
    layer5_outputs(3156) <= not(layer4_outputs(4565)) or (layer4_outputs(3405));
    layer5_outputs(3157) <= not(layer4_outputs(1260));
    layer5_outputs(3158) <= not(layer4_outputs(5459));
    layer5_outputs(3159) <= layer4_outputs(4425);
    layer5_outputs(3160) <= (layer4_outputs(5322)) and not (layer4_outputs(6022));
    layer5_outputs(3161) <= layer4_outputs(5639);
    layer5_outputs(3162) <= not(layer4_outputs(4217));
    layer5_outputs(3163) <= (layer4_outputs(5517)) xor (layer4_outputs(4975));
    layer5_outputs(3164) <= not((layer4_outputs(7579)) xor (layer4_outputs(4116)));
    layer5_outputs(3165) <= not((layer4_outputs(6572)) and (layer4_outputs(6554)));
    layer5_outputs(3166) <= (layer4_outputs(4171)) or (layer4_outputs(3426));
    layer5_outputs(3167) <= (layer4_outputs(3563)) xor (layer4_outputs(6016));
    layer5_outputs(3168) <= not(layer4_outputs(7275));
    layer5_outputs(3169) <= layer4_outputs(3474);
    layer5_outputs(3170) <= layer4_outputs(5879);
    layer5_outputs(3171) <= not(layer4_outputs(156));
    layer5_outputs(3172) <= not((layer4_outputs(6229)) xor (layer4_outputs(4763)));
    layer5_outputs(3173) <= not(layer4_outputs(7617));
    layer5_outputs(3174) <= not(layer4_outputs(5916));
    layer5_outputs(3175) <= layer4_outputs(5345);
    layer5_outputs(3176) <= layer4_outputs(780);
    layer5_outputs(3177) <= layer4_outputs(3983);
    layer5_outputs(3178) <= layer4_outputs(925);
    layer5_outputs(3179) <= layer4_outputs(6114);
    layer5_outputs(3180) <= (layer4_outputs(5873)) or (layer4_outputs(6794));
    layer5_outputs(3181) <= layer4_outputs(3816);
    layer5_outputs(3182) <= not((layer4_outputs(897)) and (layer4_outputs(4585)));
    layer5_outputs(3183) <= not(layer4_outputs(1401));
    layer5_outputs(3184) <= '1';
    layer5_outputs(3185) <= layer4_outputs(2970);
    layer5_outputs(3186) <= layer4_outputs(4419);
    layer5_outputs(3187) <= not((layer4_outputs(530)) or (layer4_outputs(4866)));
    layer5_outputs(3188) <= not(layer4_outputs(5792));
    layer5_outputs(3189) <= not(layer4_outputs(5974));
    layer5_outputs(3190) <= layer4_outputs(55);
    layer5_outputs(3191) <= layer4_outputs(1278);
    layer5_outputs(3192) <= layer4_outputs(4166);
    layer5_outputs(3193) <= not(layer4_outputs(955));
    layer5_outputs(3194) <= not(layer4_outputs(5422));
    layer5_outputs(3195) <= not(layer4_outputs(1649));
    layer5_outputs(3196) <= (layer4_outputs(1609)) and not (layer4_outputs(6489));
    layer5_outputs(3197) <= not((layer4_outputs(149)) xor (layer4_outputs(521)));
    layer5_outputs(3198) <= not((layer4_outputs(5056)) or (layer4_outputs(5684)));
    layer5_outputs(3199) <= not(layer4_outputs(6772)) or (layer4_outputs(1952));
    layer5_outputs(3200) <= (layer4_outputs(6669)) and not (layer4_outputs(1785));
    layer5_outputs(3201) <= layer4_outputs(6570);
    layer5_outputs(3202) <= not(layer4_outputs(125));
    layer5_outputs(3203) <= not(layer4_outputs(2557));
    layer5_outputs(3204) <= not(layer4_outputs(6311)) or (layer4_outputs(5585));
    layer5_outputs(3205) <= layer4_outputs(1829);
    layer5_outputs(3206) <= not(layer4_outputs(5719));
    layer5_outputs(3207) <= layer4_outputs(5751);
    layer5_outputs(3208) <= layer4_outputs(6102);
    layer5_outputs(3209) <= not((layer4_outputs(1251)) and (layer4_outputs(4056)));
    layer5_outputs(3210) <= (layer4_outputs(558)) and (layer4_outputs(4934));
    layer5_outputs(3211) <= layer4_outputs(3391);
    layer5_outputs(3212) <= not((layer4_outputs(6305)) or (layer4_outputs(5740)));
    layer5_outputs(3213) <= not(layer4_outputs(4511)) or (layer4_outputs(7248));
    layer5_outputs(3214) <= not(layer4_outputs(3872));
    layer5_outputs(3215) <= not(layer4_outputs(1974));
    layer5_outputs(3216) <= (layer4_outputs(4053)) and not (layer4_outputs(4776));
    layer5_outputs(3217) <= not((layer4_outputs(5131)) xor (layer4_outputs(1539)));
    layer5_outputs(3218) <= '1';
    layer5_outputs(3219) <= not(layer4_outputs(894));
    layer5_outputs(3220) <= layer4_outputs(6469);
    layer5_outputs(3221) <= not(layer4_outputs(3140));
    layer5_outputs(3222) <= (layer4_outputs(5148)) xor (layer4_outputs(4614));
    layer5_outputs(3223) <= (layer4_outputs(7343)) and not (layer4_outputs(5656));
    layer5_outputs(3224) <= (layer4_outputs(2013)) xor (layer4_outputs(112));
    layer5_outputs(3225) <= not(layer4_outputs(5784));
    layer5_outputs(3226) <= '1';
    layer5_outputs(3227) <= (layer4_outputs(7127)) and not (layer4_outputs(5463));
    layer5_outputs(3228) <= not(layer4_outputs(4326));
    layer5_outputs(3229) <= not((layer4_outputs(3738)) or (layer4_outputs(2456)));
    layer5_outputs(3230) <= layer4_outputs(1946);
    layer5_outputs(3231) <= not(layer4_outputs(1706));
    layer5_outputs(3232) <= layer4_outputs(59);
    layer5_outputs(3233) <= not(layer4_outputs(1425));
    layer5_outputs(3234) <= layer4_outputs(876);
    layer5_outputs(3235) <= layer4_outputs(5781);
    layer5_outputs(3236) <= '0';
    layer5_outputs(3237) <= not((layer4_outputs(367)) or (layer4_outputs(4916)));
    layer5_outputs(3238) <= not(layer4_outputs(3932));
    layer5_outputs(3239) <= (layer4_outputs(2468)) or (layer4_outputs(5197));
    layer5_outputs(3240) <= layer4_outputs(2755);
    layer5_outputs(3241) <= (layer4_outputs(1479)) and not (layer4_outputs(107));
    layer5_outputs(3242) <= not(layer4_outputs(1238));
    layer5_outputs(3243) <= (layer4_outputs(1733)) xor (layer4_outputs(6138));
    layer5_outputs(3244) <= not(layer4_outputs(3502)) or (layer4_outputs(2054));
    layer5_outputs(3245) <= layer4_outputs(681);
    layer5_outputs(3246) <= not((layer4_outputs(2896)) and (layer4_outputs(3713)));
    layer5_outputs(3247) <= not(layer4_outputs(5425));
    layer5_outputs(3248) <= '1';
    layer5_outputs(3249) <= layer4_outputs(7022);
    layer5_outputs(3250) <= not((layer4_outputs(7040)) or (layer4_outputs(3843)));
    layer5_outputs(3251) <= (layer4_outputs(6683)) and (layer4_outputs(1581));
    layer5_outputs(3252) <= not(layer4_outputs(424));
    layer5_outputs(3253) <= not(layer4_outputs(4992)) or (layer4_outputs(6600));
    layer5_outputs(3254) <= not(layer4_outputs(2623));
    layer5_outputs(3255) <= layer4_outputs(7524);
    layer5_outputs(3256) <= '0';
    layer5_outputs(3257) <= (layer4_outputs(7345)) xor (layer4_outputs(5593));
    layer5_outputs(3258) <= not(layer4_outputs(6801));
    layer5_outputs(3259) <= layer4_outputs(2458);
    layer5_outputs(3260) <= not(layer4_outputs(7162)) or (layer4_outputs(5684));
    layer5_outputs(3261) <= not((layer4_outputs(208)) or (layer4_outputs(6711)));
    layer5_outputs(3262) <= (layer4_outputs(3745)) and not (layer4_outputs(5114));
    layer5_outputs(3263) <= layer4_outputs(5731);
    layer5_outputs(3264) <= (layer4_outputs(1283)) and not (layer4_outputs(4036));
    layer5_outputs(3265) <= (layer4_outputs(3073)) or (layer4_outputs(2662));
    layer5_outputs(3266) <= layer4_outputs(2698);
    layer5_outputs(3267) <= layer4_outputs(6538);
    layer5_outputs(3268) <= not(layer4_outputs(3285));
    layer5_outputs(3269) <= (layer4_outputs(2011)) and not (layer4_outputs(6933));
    layer5_outputs(3270) <= not((layer4_outputs(1219)) or (layer4_outputs(6427)));
    layer5_outputs(3271) <= (layer4_outputs(1650)) and not (layer4_outputs(5609));
    layer5_outputs(3272) <= (layer4_outputs(3352)) and not (layer4_outputs(5114));
    layer5_outputs(3273) <= layer4_outputs(2929);
    layer5_outputs(3274) <= layer4_outputs(1948);
    layer5_outputs(3275) <= layer4_outputs(28);
    layer5_outputs(3276) <= layer4_outputs(6287);
    layer5_outputs(3277) <= not(layer4_outputs(3990)) or (layer4_outputs(4510));
    layer5_outputs(3278) <= not((layer4_outputs(4316)) and (layer4_outputs(3461)));
    layer5_outputs(3279) <= not(layer4_outputs(5414)) or (layer4_outputs(5852));
    layer5_outputs(3280) <= not((layer4_outputs(5159)) or (layer4_outputs(724)));
    layer5_outputs(3281) <= (layer4_outputs(210)) and not (layer4_outputs(6624));
    layer5_outputs(3282) <= not((layer4_outputs(7187)) and (layer4_outputs(4513)));
    layer5_outputs(3283) <= (layer4_outputs(529)) and (layer4_outputs(1817));
    layer5_outputs(3284) <= (layer4_outputs(7215)) and (layer4_outputs(1834));
    layer5_outputs(3285) <= (layer4_outputs(1428)) xor (layer4_outputs(4832));
    layer5_outputs(3286) <= '1';
    layer5_outputs(3287) <= '0';
    layer5_outputs(3288) <= not((layer4_outputs(711)) xor (layer4_outputs(6995)));
    layer5_outputs(3289) <= (layer4_outputs(3426)) or (layer4_outputs(5126));
    layer5_outputs(3290) <= not(layer4_outputs(4406)) or (layer4_outputs(1666));
    layer5_outputs(3291) <= not(layer4_outputs(6996));
    layer5_outputs(3292) <= not(layer4_outputs(6970));
    layer5_outputs(3293) <= not((layer4_outputs(4974)) and (layer4_outputs(6876)));
    layer5_outputs(3294) <= not(layer4_outputs(1498)) or (layer4_outputs(3938));
    layer5_outputs(3295) <= '0';
    layer5_outputs(3296) <= (layer4_outputs(5545)) and not (layer4_outputs(2947));
    layer5_outputs(3297) <= '0';
    layer5_outputs(3298) <= not(layer4_outputs(2518));
    layer5_outputs(3299) <= layer4_outputs(2832);
    layer5_outputs(3300) <= (layer4_outputs(5296)) and (layer4_outputs(2950));
    layer5_outputs(3301) <= (layer4_outputs(4767)) and not (layer4_outputs(30));
    layer5_outputs(3302) <= layer4_outputs(7259);
    layer5_outputs(3303) <= (layer4_outputs(7485)) or (layer4_outputs(4435));
    layer5_outputs(3304) <= not(layer4_outputs(7185));
    layer5_outputs(3305) <= layer4_outputs(6847);
    layer5_outputs(3306) <= layer4_outputs(3330);
    layer5_outputs(3307) <= '0';
    layer5_outputs(3308) <= not(layer4_outputs(6326));
    layer5_outputs(3309) <= (layer4_outputs(2288)) xor (layer4_outputs(5728));
    layer5_outputs(3310) <= (layer4_outputs(6459)) and not (layer4_outputs(1762));
    layer5_outputs(3311) <= (layer4_outputs(4452)) and not (layer4_outputs(1590));
    layer5_outputs(3312) <= not((layer4_outputs(5139)) xor (layer4_outputs(199)));
    layer5_outputs(3313) <= not(layer4_outputs(1375));
    layer5_outputs(3314) <= not((layer4_outputs(3947)) xor (layer4_outputs(1403)));
    layer5_outputs(3315) <= (layer4_outputs(3734)) and not (layer4_outputs(5504));
    layer5_outputs(3316) <= not(layer4_outputs(1135));
    layer5_outputs(3317) <= not(layer4_outputs(2848));
    layer5_outputs(3318) <= not(layer4_outputs(7522)) or (layer4_outputs(4168));
    layer5_outputs(3319) <= layer4_outputs(2544);
    layer5_outputs(3320) <= not((layer4_outputs(6013)) and (layer4_outputs(6385)));
    layer5_outputs(3321) <= layer4_outputs(3394);
    layer5_outputs(3322) <= (layer4_outputs(1203)) and (layer4_outputs(5154));
    layer5_outputs(3323) <= (layer4_outputs(6055)) and not (layer4_outputs(3607));
    layer5_outputs(3324) <= layer4_outputs(6811);
    layer5_outputs(3325) <= (layer4_outputs(1859)) xor (layer4_outputs(569));
    layer5_outputs(3326) <= not(layer4_outputs(6813));
    layer5_outputs(3327) <= (layer4_outputs(3786)) or (layer4_outputs(1861));
    layer5_outputs(3328) <= '0';
    layer5_outputs(3329) <= not(layer4_outputs(2923));
    layer5_outputs(3330) <= not((layer4_outputs(2704)) and (layer4_outputs(1443)));
    layer5_outputs(3331) <= not(layer4_outputs(5261));
    layer5_outputs(3332) <= layer4_outputs(7585);
    layer5_outputs(3333) <= not(layer4_outputs(6774));
    layer5_outputs(3334) <= not(layer4_outputs(6315));
    layer5_outputs(3335) <= not(layer4_outputs(4840)) or (layer4_outputs(2678));
    layer5_outputs(3336) <= not((layer4_outputs(5893)) or (layer4_outputs(39)));
    layer5_outputs(3337) <= layer4_outputs(4804);
    layer5_outputs(3338) <= layer4_outputs(5666);
    layer5_outputs(3339) <= layer4_outputs(5807);
    layer5_outputs(3340) <= not(layer4_outputs(4059));
    layer5_outputs(3341) <= (layer4_outputs(4795)) or (layer4_outputs(7359));
    layer5_outputs(3342) <= not(layer4_outputs(4801));
    layer5_outputs(3343) <= not(layer4_outputs(5459));
    layer5_outputs(3344) <= (layer4_outputs(3760)) and (layer4_outputs(3861));
    layer5_outputs(3345) <= (layer4_outputs(1895)) or (layer4_outputs(1601));
    layer5_outputs(3346) <= not((layer4_outputs(805)) or (layer4_outputs(343)));
    layer5_outputs(3347) <= (layer4_outputs(348)) xor (layer4_outputs(754));
    layer5_outputs(3348) <= not(layer4_outputs(1973));
    layer5_outputs(3349) <= not(layer4_outputs(3053));
    layer5_outputs(3350) <= layer4_outputs(6923);
    layer5_outputs(3351) <= (layer4_outputs(821)) or (layer4_outputs(5339));
    layer5_outputs(3352) <= not((layer4_outputs(2238)) and (layer4_outputs(5578)));
    layer5_outputs(3353) <= layer4_outputs(3739);
    layer5_outputs(3354) <= layer4_outputs(3083);
    layer5_outputs(3355) <= (layer4_outputs(31)) xor (layer4_outputs(4598));
    layer5_outputs(3356) <= not(layer4_outputs(5970)) or (layer4_outputs(6821));
    layer5_outputs(3357) <= layer4_outputs(1954);
    layer5_outputs(3358) <= not(layer4_outputs(6100));
    layer5_outputs(3359) <= not((layer4_outputs(6623)) and (layer4_outputs(5768)));
    layer5_outputs(3360) <= not((layer4_outputs(6789)) and (layer4_outputs(4321)));
    layer5_outputs(3361) <= layer4_outputs(4029);
    layer5_outputs(3362) <= layer4_outputs(4464);
    layer5_outputs(3363) <= (layer4_outputs(2403)) xor (layer4_outputs(689));
    layer5_outputs(3364) <= layer4_outputs(2916);
    layer5_outputs(3365) <= layer4_outputs(7210);
    layer5_outputs(3366) <= not(layer4_outputs(1110));
    layer5_outputs(3367) <= not(layer4_outputs(7503)) or (layer4_outputs(3230));
    layer5_outputs(3368) <= not(layer4_outputs(3124)) or (layer4_outputs(2046));
    layer5_outputs(3369) <= (layer4_outputs(2246)) and not (layer4_outputs(678));
    layer5_outputs(3370) <= not(layer4_outputs(2122)) or (layer4_outputs(5646));
    layer5_outputs(3371) <= not(layer4_outputs(250));
    layer5_outputs(3372) <= not(layer4_outputs(580));
    layer5_outputs(3373) <= (layer4_outputs(2368)) and not (layer4_outputs(5597));
    layer5_outputs(3374) <= not((layer4_outputs(2372)) and (layer4_outputs(6517)));
    layer5_outputs(3375) <= not((layer4_outputs(4100)) xor (layer4_outputs(3143)));
    layer5_outputs(3376) <= not((layer4_outputs(1188)) and (layer4_outputs(4064)));
    layer5_outputs(3377) <= not(layer4_outputs(6064));
    layer5_outputs(3378) <= not(layer4_outputs(798));
    layer5_outputs(3379) <= (layer4_outputs(582)) and not (layer4_outputs(6618));
    layer5_outputs(3380) <= not(layer4_outputs(4396));
    layer5_outputs(3381) <= not((layer4_outputs(240)) xor (layer4_outputs(1308)));
    layer5_outputs(3382) <= not(layer4_outputs(6772));
    layer5_outputs(3383) <= not(layer4_outputs(4972));
    layer5_outputs(3384) <= not(layer4_outputs(7261));
    layer5_outputs(3385) <= not(layer4_outputs(7639)) or (layer4_outputs(7194));
    layer5_outputs(3386) <= layer4_outputs(4265);
    layer5_outputs(3387) <= layer4_outputs(2918);
    layer5_outputs(3388) <= (layer4_outputs(2467)) and not (layer4_outputs(3305));
    layer5_outputs(3389) <= not(layer4_outputs(2487));
    layer5_outputs(3390) <= layer4_outputs(6569);
    layer5_outputs(3391) <= layer4_outputs(5707);
    layer5_outputs(3392) <= layer4_outputs(2560);
    layer5_outputs(3393) <= not((layer4_outputs(1885)) xor (layer4_outputs(3893)));
    layer5_outputs(3394) <= not(layer4_outputs(7654));
    layer5_outputs(3395) <= '1';
    layer5_outputs(3396) <= not(layer4_outputs(228));
    layer5_outputs(3397) <= not((layer4_outputs(2382)) and (layer4_outputs(3118)));
    layer5_outputs(3398) <= layer4_outputs(4966);
    layer5_outputs(3399) <= (layer4_outputs(676)) and not (layer4_outputs(1908));
    layer5_outputs(3400) <= not(layer4_outputs(82)) or (layer4_outputs(2872));
    layer5_outputs(3401) <= not(layer4_outputs(1900));
    layer5_outputs(3402) <= layer4_outputs(2198);
    layer5_outputs(3403) <= (layer4_outputs(6165)) and not (layer4_outputs(3131));
    layer5_outputs(3404) <= (layer4_outputs(1871)) and (layer4_outputs(1460));
    layer5_outputs(3405) <= not(layer4_outputs(4200));
    layer5_outputs(3406) <= not(layer4_outputs(4252));
    layer5_outputs(3407) <= (layer4_outputs(5146)) xor (layer4_outputs(2529));
    layer5_outputs(3408) <= layer4_outputs(6900);
    layer5_outputs(3409) <= (layer4_outputs(6952)) and not (layer4_outputs(1263));
    layer5_outputs(3410) <= (layer4_outputs(2720)) or (layer4_outputs(6749));
    layer5_outputs(3411) <= not(layer4_outputs(5212));
    layer5_outputs(3412) <= not(layer4_outputs(5873));
    layer5_outputs(3413) <= not(layer4_outputs(2396));
    layer5_outputs(3414) <= layer4_outputs(3022);
    layer5_outputs(3415) <= layer4_outputs(6647);
    layer5_outputs(3416) <= layer4_outputs(1409);
    layer5_outputs(3417) <= not((layer4_outputs(5749)) xor (layer4_outputs(900)));
    layer5_outputs(3418) <= not((layer4_outputs(5391)) and (layer4_outputs(2457)));
    layer5_outputs(3419) <= not((layer4_outputs(4483)) xor (layer4_outputs(1874)));
    layer5_outputs(3420) <= not(layer4_outputs(7451));
    layer5_outputs(3421) <= not((layer4_outputs(3866)) xor (layer4_outputs(2762)));
    layer5_outputs(3422) <= not((layer4_outputs(7563)) or (layer4_outputs(3723)));
    layer5_outputs(3423) <= not(layer4_outputs(5811));
    layer5_outputs(3424) <= not(layer4_outputs(1358));
    layer5_outputs(3425) <= not(layer4_outputs(6512)) or (layer4_outputs(2857));
    layer5_outputs(3426) <= layer4_outputs(4361);
    layer5_outputs(3427) <= not(layer4_outputs(6000)) or (layer4_outputs(2463));
    layer5_outputs(3428) <= layer4_outputs(1835);
    layer5_outputs(3429) <= not((layer4_outputs(2376)) and (layer4_outputs(3194)));
    layer5_outputs(3430) <= (layer4_outputs(5041)) xor (layer4_outputs(268));
    layer5_outputs(3431) <= layer4_outputs(5150);
    layer5_outputs(3432) <= not(layer4_outputs(6893));
    layer5_outputs(3433) <= layer4_outputs(6860);
    layer5_outputs(3434) <= not((layer4_outputs(5802)) or (layer4_outputs(5142)));
    layer5_outputs(3435) <= (layer4_outputs(1030)) and (layer4_outputs(1502));
    layer5_outputs(3436) <= (layer4_outputs(1304)) and not (layer4_outputs(4534));
    layer5_outputs(3437) <= (layer4_outputs(1858)) and not (layer4_outputs(6805));
    layer5_outputs(3438) <= (layer4_outputs(546)) and not (layer4_outputs(4671));
    layer5_outputs(3439) <= layer4_outputs(3781);
    layer5_outputs(3440) <= layer4_outputs(5674);
    layer5_outputs(3441) <= not((layer4_outputs(4822)) or (layer4_outputs(5645)));
    layer5_outputs(3442) <= (layer4_outputs(962)) and not (layer4_outputs(3446));
    layer5_outputs(3443) <= (layer4_outputs(14)) and not (layer4_outputs(398));
    layer5_outputs(3444) <= '0';
    layer5_outputs(3445) <= not(layer4_outputs(5705));
    layer5_outputs(3446) <= (layer4_outputs(1670)) and (layer4_outputs(2553));
    layer5_outputs(3447) <= not(layer4_outputs(5090));
    layer5_outputs(3448) <= not(layer4_outputs(3563));
    layer5_outputs(3449) <= not(layer4_outputs(4770));
    layer5_outputs(3450) <= not(layer4_outputs(6130));
    layer5_outputs(3451) <= not(layer4_outputs(2804));
    layer5_outputs(3452) <= layer4_outputs(3086);
    layer5_outputs(3453) <= layer4_outputs(3295);
    layer5_outputs(3454) <= '0';
    layer5_outputs(3455) <= layer4_outputs(5176);
    layer5_outputs(3456) <= not(layer4_outputs(2127));
    layer5_outputs(3457) <= (layer4_outputs(1654)) and not (layer4_outputs(6825));
    layer5_outputs(3458) <= (layer4_outputs(3077)) and not (layer4_outputs(3453));
    layer5_outputs(3459) <= layer4_outputs(4218);
    layer5_outputs(3460) <= not(layer4_outputs(7190)) or (layer4_outputs(1515));
    layer5_outputs(3461) <= layer4_outputs(2113);
    layer5_outputs(3462) <= layer4_outputs(168);
    layer5_outputs(3463) <= (layer4_outputs(1945)) and not (layer4_outputs(5027));
    layer5_outputs(3464) <= '0';
    layer5_outputs(3465) <= not(layer4_outputs(5129)) or (layer4_outputs(2021));
    layer5_outputs(3466) <= not(layer4_outputs(6065));
    layer5_outputs(3467) <= not(layer4_outputs(2145)) or (layer4_outputs(5300));
    layer5_outputs(3468) <= '0';
    layer5_outputs(3469) <= not(layer4_outputs(5928));
    layer5_outputs(3470) <= '0';
    layer5_outputs(3471) <= not(layer4_outputs(6206));
    layer5_outputs(3472) <= not((layer4_outputs(4386)) and (layer4_outputs(5280)));
    layer5_outputs(3473) <= not((layer4_outputs(4841)) xor (layer4_outputs(5829)));
    layer5_outputs(3474) <= not((layer4_outputs(242)) or (layer4_outputs(1912)));
    layer5_outputs(3475) <= layer4_outputs(6856);
    layer5_outputs(3476) <= not((layer4_outputs(2840)) or (layer4_outputs(2268)));
    layer5_outputs(3477) <= layer4_outputs(6556);
    layer5_outputs(3478) <= layer4_outputs(1150);
    layer5_outputs(3479) <= layer4_outputs(3478);
    layer5_outputs(3480) <= layer4_outputs(3232);
    layer5_outputs(3481) <= not(layer4_outputs(3550));
    layer5_outputs(3482) <= layer4_outputs(4270);
    layer5_outputs(3483) <= '1';
    layer5_outputs(3484) <= not((layer4_outputs(4830)) or (layer4_outputs(3541)));
    layer5_outputs(3485) <= layer4_outputs(394);
    layer5_outputs(3486) <= not(layer4_outputs(3076)) or (layer4_outputs(6873));
    layer5_outputs(3487) <= not(layer4_outputs(5811));
    layer5_outputs(3488) <= (layer4_outputs(4977)) xor (layer4_outputs(7326));
    layer5_outputs(3489) <= layer4_outputs(6879);
    layer5_outputs(3490) <= (layer4_outputs(3877)) xor (layer4_outputs(3864));
    layer5_outputs(3491) <= not((layer4_outputs(1747)) and (layer4_outputs(5027)));
    layer5_outputs(3492) <= '0';
    layer5_outputs(3493) <= (layer4_outputs(4544)) and (layer4_outputs(557));
    layer5_outputs(3494) <= (layer4_outputs(1660)) xor (layer4_outputs(3733));
    layer5_outputs(3495) <= not((layer4_outputs(4991)) or (layer4_outputs(2379)));
    layer5_outputs(3496) <= (layer4_outputs(1223)) and (layer4_outputs(1835));
    layer5_outputs(3497) <= not(layer4_outputs(7277));
    layer5_outputs(3498) <= not((layer4_outputs(5392)) xor (layer4_outputs(7646)));
    layer5_outputs(3499) <= not(layer4_outputs(3653));
    layer5_outputs(3500) <= not(layer4_outputs(7614));
    layer5_outputs(3501) <= (layer4_outputs(56)) and not (layer4_outputs(2932));
    layer5_outputs(3502) <= not(layer4_outputs(1038));
    layer5_outputs(3503) <= not((layer4_outputs(3168)) or (layer4_outputs(2836)));
    layer5_outputs(3504) <= (layer4_outputs(5934)) and not (layer4_outputs(6826));
    layer5_outputs(3505) <= not(layer4_outputs(2112));
    layer5_outputs(3506) <= '0';
    layer5_outputs(3507) <= not((layer4_outputs(7598)) xor (layer4_outputs(151)));
    layer5_outputs(3508) <= layer4_outputs(3176);
    layer5_outputs(3509) <= layer4_outputs(7081);
    layer5_outputs(3510) <= layer4_outputs(6065);
    layer5_outputs(3511) <= not(layer4_outputs(6672));
    layer5_outputs(3512) <= layer4_outputs(3522);
    layer5_outputs(3513) <= (layer4_outputs(1274)) xor (layer4_outputs(7218));
    layer5_outputs(3514) <= layer4_outputs(1216);
    layer5_outputs(3515) <= not(layer4_outputs(6573)) or (layer4_outputs(7414));
    layer5_outputs(3516) <= not((layer4_outputs(3704)) xor (layer4_outputs(5245)));
    layer5_outputs(3517) <= not(layer4_outputs(3033));
    layer5_outputs(3518) <= (layer4_outputs(6053)) or (layer4_outputs(6969));
    layer5_outputs(3519) <= not((layer4_outputs(1997)) xor (layer4_outputs(7567)));
    layer5_outputs(3520) <= (layer4_outputs(6565)) or (layer4_outputs(1402));
    layer5_outputs(3521) <= not(layer4_outputs(4474)) or (layer4_outputs(767));
    layer5_outputs(3522) <= layer4_outputs(6437);
    layer5_outputs(3523) <= not(layer4_outputs(6837)) or (layer4_outputs(2738));
    layer5_outputs(3524) <= (layer4_outputs(5521)) xor (layer4_outputs(5353));
    layer5_outputs(3525) <= not(layer4_outputs(7267)) or (layer4_outputs(2978));
    layer5_outputs(3526) <= not(layer4_outputs(5088)) or (layer4_outputs(1023));
    layer5_outputs(3527) <= (layer4_outputs(2220)) and not (layer4_outputs(1363));
    layer5_outputs(3528) <= (layer4_outputs(1481)) xor (layer4_outputs(1141));
    layer5_outputs(3529) <= (layer4_outputs(4314)) and not (layer4_outputs(3383));
    layer5_outputs(3530) <= (layer4_outputs(4461)) and not (layer4_outputs(5770));
    layer5_outputs(3531) <= not(layer4_outputs(2570));
    layer5_outputs(3532) <= (layer4_outputs(5104)) and not (layer4_outputs(5775));
    layer5_outputs(3533) <= (layer4_outputs(6550)) and (layer4_outputs(6597));
    layer5_outputs(3534) <= (layer4_outputs(2268)) or (layer4_outputs(6435));
    layer5_outputs(3535) <= not(layer4_outputs(1948));
    layer5_outputs(3536) <= not((layer4_outputs(1173)) xor (layer4_outputs(1529)));
    layer5_outputs(3537) <= layer4_outputs(4968);
    layer5_outputs(3538) <= '0';
    layer5_outputs(3539) <= layer4_outputs(5892);
    layer5_outputs(3540) <= not(layer4_outputs(6976));
    layer5_outputs(3541) <= not((layer4_outputs(4040)) xor (layer4_outputs(26)));
    layer5_outputs(3542) <= (layer4_outputs(1427)) and not (layer4_outputs(2423));
    layer5_outputs(3543) <= '1';
    layer5_outputs(3544) <= (layer4_outputs(253)) and not (layer4_outputs(4925));
    layer5_outputs(3545) <= (layer4_outputs(2241)) or (layer4_outputs(5466));
    layer5_outputs(3546) <= not(layer4_outputs(5858)) or (layer4_outputs(4409));
    layer5_outputs(3547) <= '1';
    layer5_outputs(3548) <= not(layer4_outputs(4184));
    layer5_outputs(3549) <= (layer4_outputs(4229)) xor (layer4_outputs(3183));
    layer5_outputs(3550) <= layer4_outputs(2559);
    layer5_outputs(3551) <= (layer4_outputs(3158)) xor (layer4_outputs(4159));
    layer5_outputs(3552) <= not((layer4_outputs(2259)) xor (layer4_outputs(6063)));
    layer5_outputs(3553) <= not((layer4_outputs(791)) and (layer4_outputs(345)));
    layer5_outputs(3554) <= (layer4_outputs(5920)) and not (layer4_outputs(1209));
    layer5_outputs(3555) <= not(layer4_outputs(3898));
    layer5_outputs(3556) <= (layer4_outputs(6688)) and (layer4_outputs(2386));
    layer5_outputs(3557) <= '0';
    layer5_outputs(3558) <= (layer4_outputs(2064)) xor (layer4_outputs(4971));
    layer5_outputs(3559) <= not(layer4_outputs(2648));
    layer5_outputs(3560) <= layer4_outputs(6059);
    layer5_outputs(3561) <= layer4_outputs(1156);
    layer5_outputs(3562) <= not((layer4_outputs(6959)) or (layer4_outputs(2078)));
    layer5_outputs(3563) <= layer4_outputs(2342);
    layer5_outputs(3564) <= not(layer4_outputs(5638));
    layer5_outputs(3565) <= (layer4_outputs(4417)) and not (layer4_outputs(1981));
    layer5_outputs(3566) <= not(layer4_outputs(4197));
    layer5_outputs(3567) <= (layer4_outputs(6394)) and (layer4_outputs(3665));
    layer5_outputs(3568) <= not((layer4_outputs(7332)) xor (layer4_outputs(2802)));
    layer5_outputs(3569) <= (layer4_outputs(2638)) and (layer4_outputs(1207));
    layer5_outputs(3570) <= not(layer4_outputs(1494)) or (layer4_outputs(4121));
    layer5_outputs(3571) <= not(layer4_outputs(798));
    layer5_outputs(3572) <= (layer4_outputs(3494)) and not (layer4_outputs(1798));
    layer5_outputs(3573) <= not(layer4_outputs(6279));
    layer5_outputs(3574) <= (layer4_outputs(2887)) and (layer4_outputs(6585));
    layer5_outputs(3575) <= layer4_outputs(1975);
    layer5_outputs(3576) <= not(layer4_outputs(441));
    layer5_outputs(3577) <= (layer4_outputs(2861)) and (layer4_outputs(6373));
    layer5_outputs(3578) <= layer4_outputs(4015);
    layer5_outputs(3579) <= (layer4_outputs(2165)) and not (layer4_outputs(5017));
    layer5_outputs(3580) <= not(layer4_outputs(1117));
    layer5_outputs(3581) <= (layer4_outputs(2843)) and not (layer4_outputs(3676));
    layer5_outputs(3582) <= layer4_outputs(6136);
    layer5_outputs(3583) <= (layer4_outputs(935)) or (layer4_outputs(7598));
    layer5_outputs(3584) <= not((layer4_outputs(7339)) or (layer4_outputs(2684)));
    layer5_outputs(3585) <= not(layer4_outputs(5319)) or (layer4_outputs(964));
    layer5_outputs(3586) <= layer4_outputs(1212);
    layer5_outputs(3587) <= not(layer4_outputs(4122));
    layer5_outputs(3588) <= (layer4_outputs(3100)) xor (layer4_outputs(7303));
    layer5_outputs(3589) <= (layer4_outputs(2284)) and not (layer4_outputs(2229));
    layer5_outputs(3590) <= not(layer4_outputs(3243)) or (layer4_outputs(7641));
    layer5_outputs(3591) <= (layer4_outputs(2694)) or (layer4_outputs(2331));
    layer5_outputs(3592) <= not(layer4_outputs(1092));
    layer5_outputs(3593) <= not(layer4_outputs(4823));
    layer5_outputs(3594) <= not((layer4_outputs(4321)) xor (layer4_outputs(6400)));
    layer5_outputs(3595) <= not(layer4_outputs(95));
    layer5_outputs(3596) <= not(layer4_outputs(1945)) or (layer4_outputs(276));
    layer5_outputs(3597) <= not(layer4_outputs(4576));
    layer5_outputs(3598) <= (layer4_outputs(5526)) xor (layer4_outputs(457));
    layer5_outputs(3599) <= (layer4_outputs(1165)) xor (layer4_outputs(5230));
    layer5_outputs(3600) <= not(layer4_outputs(7409));
    layer5_outputs(3601) <= layer4_outputs(6219);
    layer5_outputs(3602) <= not(layer4_outputs(793));
    layer5_outputs(3603) <= (layer4_outputs(337)) xor (layer4_outputs(4066));
    layer5_outputs(3604) <= layer4_outputs(7131);
    layer5_outputs(3605) <= not((layer4_outputs(2629)) and (layer4_outputs(7459)));
    layer5_outputs(3606) <= not((layer4_outputs(6490)) xor (layer4_outputs(5530)));
    layer5_outputs(3607) <= (layer4_outputs(2435)) and not (layer4_outputs(2444));
    layer5_outputs(3608) <= (layer4_outputs(4776)) and not (layer4_outputs(3393));
    layer5_outputs(3609) <= layer4_outputs(4424);
    layer5_outputs(3610) <= not(layer4_outputs(3182)) or (layer4_outputs(1422));
    layer5_outputs(3611) <= layer4_outputs(4594);
    layer5_outputs(3612) <= not(layer4_outputs(7508)) or (layer4_outputs(6101));
    layer5_outputs(3613) <= layer4_outputs(4173);
    layer5_outputs(3614) <= (layer4_outputs(2430)) and not (layer4_outputs(3191));
    layer5_outputs(3615) <= (layer4_outputs(4783)) xor (layer4_outputs(907));
    layer5_outputs(3616) <= not(layer4_outputs(733));
    layer5_outputs(3617) <= not(layer4_outputs(5486));
    layer5_outputs(3618) <= (layer4_outputs(2917)) or (layer4_outputs(2578));
    layer5_outputs(3619) <= layer4_outputs(6478);
    layer5_outputs(3620) <= not(layer4_outputs(4563));
    layer5_outputs(3621) <= (layer4_outputs(609)) and (layer4_outputs(5138));
    layer5_outputs(3622) <= not(layer4_outputs(2004));
    layer5_outputs(3623) <= (layer4_outputs(3917)) or (layer4_outputs(6723));
    layer5_outputs(3624) <= not((layer4_outputs(1555)) xor (layer4_outputs(2417)));
    layer5_outputs(3625) <= layer4_outputs(6403);
    layer5_outputs(3626) <= (layer4_outputs(6580)) and (layer4_outputs(1696));
    layer5_outputs(3627) <= not(layer4_outputs(1426));
    layer5_outputs(3628) <= layer4_outputs(3246);
    layer5_outputs(3629) <= (layer4_outputs(5786)) and (layer4_outputs(5363));
    layer5_outputs(3630) <= layer4_outputs(6855);
    layer5_outputs(3631) <= not(layer4_outputs(6789));
    layer5_outputs(3632) <= layer4_outputs(6450);
    layer5_outputs(3633) <= not(layer4_outputs(2219));
    layer5_outputs(3634) <= (layer4_outputs(4453)) and (layer4_outputs(1709));
    layer5_outputs(3635) <= not(layer4_outputs(2918));
    layer5_outputs(3636) <= (layer4_outputs(712)) or (layer4_outputs(381));
    layer5_outputs(3637) <= (layer4_outputs(284)) and not (layer4_outputs(6209));
    layer5_outputs(3638) <= layer4_outputs(6231);
    layer5_outputs(3639) <= (layer4_outputs(3419)) and (layer4_outputs(6080));
    layer5_outputs(3640) <= (layer4_outputs(4834)) and not (layer4_outputs(1069));
    layer5_outputs(3641) <= (layer4_outputs(5044)) and not (layer4_outputs(5032));
    layer5_outputs(3642) <= not((layer4_outputs(2140)) xor (layer4_outputs(837)));
    layer5_outputs(3643) <= layer4_outputs(653);
    layer5_outputs(3644) <= (layer4_outputs(4554)) or (layer4_outputs(4641));
    layer5_outputs(3645) <= layer4_outputs(738);
    layer5_outputs(3646) <= not(layer4_outputs(6966));
    layer5_outputs(3647) <= not((layer4_outputs(4937)) or (layer4_outputs(1772)));
    layer5_outputs(3648) <= not(layer4_outputs(1465));
    layer5_outputs(3649) <= not((layer4_outputs(4974)) or (layer4_outputs(396)));
    layer5_outputs(3650) <= not(layer4_outputs(6129)) or (layer4_outputs(3861));
    layer5_outputs(3651) <= (layer4_outputs(5387)) or (layer4_outputs(1655));
    layer5_outputs(3652) <= layer4_outputs(6568);
    layer5_outputs(3653) <= not((layer4_outputs(4636)) or (layer4_outputs(5339)));
    layer5_outputs(3654) <= (layer4_outputs(579)) xor (layer4_outputs(3));
    layer5_outputs(3655) <= layer4_outputs(7389);
    layer5_outputs(3656) <= (layer4_outputs(7549)) and not (layer4_outputs(1695));
    layer5_outputs(3657) <= (layer4_outputs(2333)) or (layer4_outputs(5521));
    layer5_outputs(3658) <= not((layer4_outputs(6505)) or (layer4_outputs(1595)));
    layer5_outputs(3659) <= not(layer4_outputs(6299));
    layer5_outputs(3660) <= not(layer4_outputs(6376));
    layer5_outputs(3661) <= not(layer4_outputs(7360)) or (layer4_outputs(1347));
    layer5_outputs(3662) <= not(layer4_outputs(1087));
    layer5_outputs(3663) <= (layer4_outputs(512)) or (layer4_outputs(407));
    layer5_outputs(3664) <= layer4_outputs(892);
    layer5_outputs(3665) <= not(layer4_outputs(6718));
    layer5_outputs(3666) <= (layer4_outputs(7420)) xor (layer4_outputs(372));
    layer5_outputs(3667) <= (layer4_outputs(5424)) or (layer4_outputs(4238));
    layer5_outputs(3668) <= not(layer4_outputs(885));
    layer5_outputs(3669) <= (layer4_outputs(4761)) xor (layer4_outputs(7566));
    layer5_outputs(3670) <= layer4_outputs(715);
    layer5_outputs(3671) <= not(layer4_outputs(1300));
    layer5_outputs(3672) <= (layer4_outputs(5130)) and not (layer4_outputs(3181));
    layer5_outputs(3673) <= layer4_outputs(4028);
    layer5_outputs(3674) <= layer4_outputs(287);
    layer5_outputs(3675) <= not(layer4_outputs(3640)) or (layer4_outputs(7118));
    layer5_outputs(3676) <= (layer4_outputs(2861)) or (layer4_outputs(3790));
    layer5_outputs(3677) <= not(layer4_outputs(5021));
    layer5_outputs(3678) <= '0';
    layer5_outputs(3679) <= not(layer4_outputs(2782)) or (layer4_outputs(5897));
    layer5_outputs(3680) <= layer4_outputs(4169);
    layer5_outputs(3681) <= not((layer4_outputs(6608)) and (layer4_outputs(6774)));
    layer5_outputs(3682) <= (layer4_outputs(1226)) xor (layer4_outputs(5685));
    layer5_outputs(3683) <= layer4_outputs(2185);
    layer5_outputs(3684) <= (layer4_outputs(2072)) and not (layer4_outputs(7254));
    layer5_outputs(3685) <= (layer4_outputs(2309)) and not (layer4_outputs(4935));
    layer5_outputs(3686) <= not(layer4_outputs(5987)) or (layer4_outputs(3270));
    layer5_outputs(3687) <= layer4_outputs(5997);
    layer5_outputs(3688) <= (layer4_outputs(7273)) or (layer4_outputs(807));
    layer5_outputs(3689) <= not(layer4_outputs(306)) or (layer4_outputs(6714));
    layer5_outputs(3690) <= not(layer4_outputs(6306));
    layer5_outputs(3691) <= layer4_outputs(3119);
    layer5_outputs(3692) <= not((layer4_outputs(4724)) and (layer4_outputs(2938)));
    layer5_outputs(3693) <= not((layer4_outputs(1637)) and (layer4_outputs(3195)));
    layer5_outputs(3694) <= not((layer4_outputs(1857)) or (layer4_outputs(509)));
    layer5_outputs(3695) <= (layer4_outputs(6897)) or (layer4_outputs(610));
    layer5_outputs(3696) <= not(layer4_outputs(5928));
    layer5_outputs(3697) <= layer4_outputs(6425);
    layer5_outputs(3698) <= layer4_outputs(6320);
    layer5_outputs(3699) <= not((layer4_outputs(2371)) or (layer4_outputs(6958)));
    layer5_outputs(3700) <= not(layer4_outputs(4394)) or (layer4_outputs(3891));
    layer5_outputs(3701) <= layer4_outputs(104);
    layer5_outputs(3702) <= not((layer4_outputs(1529)) xor (layer4_outputs(4908)));
    layer5_outputs(3703) <= not((layer4_outputs(648)) xor (layer4_outputs(6571)));
    layer5_outputs(3704) <= not(layer4_outputs(311));
    layer5_outputs(3705) <= (layer4_outputs(1385)) xor (layer4_outputs(3900));
    layer5_outputs(3706) <= (layer4_outputs(1299)) or (layer4_outputs(2814));
    layer5_outputs(3707) <= '1';
    layer5_outputs(3708) <= layer4_outputs(1187);
    layer5_outputs(3709) <= layer4_outputs(5012);
    layer5_outputs(3710) <= layer4_outputs(3455);
    layer5_outputs(3711) <= (layer4_outputs(5516)) and (layer4_outputs(1951));
    layer5_outputs(3712) <= (layer4_outputs(2069)) and not (layer4_outputs(6368));
    layer5_outputs(3713) <= layer4_outputs(6173);
    layer5_outputs(3714) <= not(layer4_outputs(7336));
    layer5_outputs(3715) <= layer4_outputs(5059);
    layer5_outputs(3716) <= not(layer4_outputs(4813));
    layer5_outputs(3717) <= not(layer4_outputs(4299));
    layer5_outputs(3718) <= not(layer4_outputs(7133)) or (layer4_outputs(3496));
    layer5_outputs(3719) <= not(layer4_outputs(538));
    layer5_outputs(3720) <= (layer4_outputs(1203)) and not (layer4_outputs(4303));
    layer5_outputs(3721) <= (layer4_outputs(6764)) and not (layer4_outputs(6074));
    layer5_outputs(3722) <= not((layer4_outputs(3747)) xor (layer4_outputs(462)));
    layer5_outputs(3723) <= not((layer4_outputs(583)) and (layer4_outputs(7012)));
    layer5_outputs(3724) <= (layer4_outputs(3927)) and not (layer4_outputs(6035));
    layer5_outputs(3725) <= not(layer4_outputs(5496));
    layer5_outputs(3726) <= (layer4_outputs(3421)) and (layer4_outputs(3545));
    layer5_outputs(3727) <= not(layer4_outputs(7323));
    layer5_outputs(3728) <= layer4_outputs(3827);
    layer5_outputs(3729) <= not(layer4_outputs(2109));
    layer5_outputs(3730) <= not(layer4_outputs(3664));
    layer5_outputs(3731) <= not(layer4_outputs(6728));
    layer5_outputs(3732) <= layer4_outputs(4574);
    layer5_outputs(3733) <= layer4_outputs(4101);
    layer5_outputs(3734) <= not((layer4_outputs(3264)) xor (layer4_outputs(2251)));
    layer5_outputs(3735) <= layer4_outputs(4077);
    layer5_outputs(3736) <= layer4_outputs(3539);
    layer5_outputs(3737) <= layer4_outputs(2572);
    layer5_outputs(3738) <= not(layer4_outputs(5639));
    layer5_outputs(3739) <= layer4_outputs(7375);
    layer5_outputs(3740) <= (layer4_outputs(4019)) and (layer4_outputs(2160));
    layer5_outputs(3741) <= (layer4_outputs(3003)) and not (layer4_outputs(6647));
    layer5_outputs(3742) <= (layer4_outputs(7216)) and not (layer4_outputs(2347));
    layer5_outputs(3743) <= not(layer4_outputs(4644));
    layer5_outputs(3744) <= not((layer4_outputs(254)) xor (layer4_outputs(882)));
    layer5_outputs(3745) <= (layer4_outputs(4583)) xor (layer4_outputs(7140));
    layer5_outputs(3746) <= not((layer4_outputs(2108)) and (layer4_outputs(5891)));
    layer5_outputs(3747) <= not((layer4_outputs(3181)) xor (layer4_outputs(3226)));
    layer5_outputs(3748) <= layer4_outputs(518);
    layer5_outputs(3749) <= layer4_outputs(298);
    layer5_outputs(3750) <= not((layer4_outputs(3455)) or (layer4_outputs(6687)));
    layer5_outputs(3751) <= layer4_outputs(3797);
    layer5_outputs(3752) <= layer4_outputs(959);
    layer5_outputs(3753) <= layer4_outputs(4473);
    layer5_outputs(3754) <= not((layer4_outputs(4485)) or (layer4_outputs(2779)));
    layer5_outputs(3755) <= not(layer4_outputs(3807));
    layer5_outputs(3756) <= not(layer4_outputs(1880));
    layer5_outputs(3757) <= layer4_outputs(669);
    layer5_outputs(3758) <= layer4_outputs(3342);
    layer5_outputs(3759) <= layer4_outputs(5172);
    layer5_outputs(3760) <= not(layer4_outputs(4749));
    layer5_outputs(3761) <= layer4_outputs(6530);
    layer5_outputs(3762) <= (layer4_outputs(623)) and (layer4_outputs(2192));
    layer5_outputs(3763) <= not(layer4_outputs(4851));
    layer5_outputs(3764) <= layer4_outputs(7484);
    layer5_outputs(3765) <= (layer4_outputs(3410)) xor (layer4_outputs(3129));
    layer5_outputs(3766) <= (layer4_outputs(888)) and not (layer4_outputs(3062));
    layer5_outputs(3767) <= not(layer4_outputs(5792)) or (layer4_outputs(5889));
    layer5_outputs(3768) <= layer4_outputs(6188);
    layer5_outputs(3769) <= not((layer4_outputs(7638)) and (layer4_outputs(3414)));
    layer5_outputs(3770) <= not(layer4_outputs(6389));
    layer5_outputs(3771) <= layer4_outputs(471);
    layer5_outputs(3772) <= not(layer4_outputs(546));
    layer5_outputs(3773) <= layer4_outputs(6777);
    layer5_outputs(3774) <= not(layer4_outputs(5774));
    layer5_outputs(3775) <= not(layer4_outputs(7243)) or (layer4_outputs(3965));
    layer5_outputs(3776) <= (layer4_outputs(1940)) and (layer4_outputs(6982));
    layer5_outputs(3777) <= not(layer4_outputs(630));
    layer5_outputs(3778) <= (layer4_outputs(3975)) or (layer4_outputs(7678));
    layer5_outputs(3779) <= not(layer4_outputs(5561));
    layer5_outputs(3780) <= not(layer4_outputs(7252));
    layer5_outputs(3781) <= not((layer4_outputs(5948)) xor (layer4_outputs(2615)));
    layer5_outputs(3782) <= (layer4_outputs(1915)) and not (layer4_outputs(5137));
    layer5_outputs(3783) <= layer4_outputs(4153);
    layer5_outputs(3784) <= (layer4_outputs(6798)) xor (layer4_outputs(1497));
    layer5_outputs(3785) <= not(layer4_outputs(6822)) or (layer4_outputs(3554));
    layer5_outputs(3786) <= not((layer4_outputs(4178)) xor (layer4_outputs(4959)));
    layer5_outputs(3787) <= '0';
    layer5_outputs(3788) <= not((layer4_outputs(5098)) xor (layer4_outputs(7592)));
    layer5_outputs(3789) <= not(layer4_outputs(6014));
    layer5_outputs(3790) <= not(layer4_outputs(5934));
    layer5_outputs(3791) <= not((layer4_outputs(4512)) and (layer4_outputs(3621)));
    layer5_outputs(3792) <= not(layer4_outputs(4231));
    layer5_outputs(3793) <= layer4_outputs(1393);
    layer5_outputs(3794) <= not(layer4_outputs(4516));
    layer5_outputs(3795) <= not(layer4_outputs(704));
    layer5_outputs(3796) <= not(layer4_outputs(5644));
    layer5_outputs(3797) <= not(layer4_outputs(5836)) or (layer4_outputs(2199));
    layer5_outputs(3798) <= layer4_outputs(6082);
    layer5_outputs(3799) <= not(layer4_outputs(1974));
    layer5_outputs(3800) <= not(layer4_outputs(3001));
    layer5_outputs(3801) <= layer4_outputs(5564);
    layer5_outputs(3802) <= '0';
    layer5_outputs(3803) <= layer4_outputs(5360);
    layer5_outputs(3804) <= not((layer4_outputs(4462)) xor (layer4_outputs(823)));
    layer5_outputs(3805) <= layer4_outputs(3162);
    layer5_outputs(3806) <= not(layer4_outputs(7207));
    layer5_outputs(3807) <= (layer4_outputs(4340)) and not (layer4_outputs(7129));
    layer5_outputs(3808) <= (layer4_outputs(1486)) and not (layer4_outputs(3219));
    layer5_outputs(3809) <= not(layer4_outputs(6653)) or (layer4_outputs(2355));
    layer5_outputs(3810) <= (layer4_outputs(4541)) or (layer4_outputs(1640));
    layer5_outputs(3811) <= (layer4_outputs(269)) or (layer4_outputs(3216));
    layer5_outputs(3812) <= not(layer4_outputs(2331));
    layer5_outputs(3813) <= not(layer4_outputs(4920)) or (layer4_outputs(2211));
    layer5_outputs(3814) <= layer4_outputs(4107);
    layer5_outputs(3815) <= not(layer4_outputs(5362));
    layer5_outputs(3816) <= layer4_outputs(3148);
    layer5_outputs(3817) <= layer4_outputs(1830);
    layer5_outputs(3818) <= (layer4_outputs(5096)) xor (layer4_outputs(7177));
    layer5_outputs(3819) <= not(layer4_outputs(6911)) or (layer4_outputs(2372));
    layer5_outputs(3820) <= not(layer4_outputs(7626));
    layer5_outputs(3821) <= not(layer4_outputs(4230));
    layer5_outputs(3822) <= not((layer4_outputs(3137)) xor (layer4_outputs(2411)));
    layer5_outputs(3823) <= not(layer4_outputs(1525));
    layer5_outputs(3824) <= (layer4_outputs(7316)) xor (layer4_outputs(6667));
    layer5_outputs(3825) <= not((layer4_outputs(5803)) xor (layer4_outputs(1710)));
    layer5_outputs(3826) <= layer4_outputs(3747);
    layer5_outputs(3827) <= not(layer4_outputs(4601));
    layer5_outputs(3828) <= not(layer4_outputs(2047));
    layer5_outputs(3829) <= not((layer4_outputs(3824)) xor (layer4_outputs(4385)));
    layer5_outputs(3830) <= not((layer4_outputs(4990)) and (layer4_outputs(596)));
    layer5_outputs(3831) <= layer4_outputs(5862);
    layer5_outputs(3832) <= layer4_outputs(5161);
    layer5_outputs(3833) <= layer4_outputs(1025);
    layer5_outputs(3834) <= (layer4_outputs(3601)) and not (layer4_outputs(1961));
    layer5_outputs(3835) <= (layer4_outputs(5903)) or (layer4_outputs(7665));
    layer5_outputs(3836) <= '1';
    layer5_outputs(3837) <= (layer4_outputs(6522)) or (layer4_outputs(919));
    layer5_outputs(3838) <= not(layer4_outputs(2345));
    layer5_outputs(3839) <= layer4_outputs(1101);
    layer5_outputs(3840) <= (layer4_outputs(4674)) or (layer4_outputs(1802));
    layer5_outputs(3841) <= not(layer4_outputs(5009)) or (layer4_outputs(693));
    layer5_outputs(3842) <= layer4_outputs(5170);
    layer5_outputs(3843) <= not(layer4_outputs(3220)) or (layer4_outputs(5253));
    layer5_outputs(3844) <= not((layer4_outputs(2075)) xor (layer4_outputs(4140)));
    layer5_outputs(3845) <= not(layer4_outputs(6079)) or (layer4_outputs(208));
    layer5_outputs(3846) <= layer4_outputs(477);
    layer5_outputs(3847) <= not((layer4_outputs(3061)) or (layer4_outputs(3125)));
    layer5_outputs(3848) <= not(layer4_outputs(7314));
    layer5_outputs(3849) <= layer4_outputs(2905);
    layer5_outputs(3850) <= layer4_outputs(4793);
    layer5_outputs(3851) <= not(layer4_outputs(987));
    layer5_outputs(3852) <= not(layer4_outputs(6978));
    layer5_outputs(3853) <= (layer4_outputs(4408)) and not (layer4_outputs(7013));
    layer5_outputs(3854) <= not((layer4_outputs(5943)) xor (layer4_outputs(370)));
    layer5_outputs(3855) <= layer4_outputs(5322);
    layer5_outputs(3856) <= not(layer4_outputs(2443));
    layer5_outputs(3857) <= not((layer4_outputs(577)) or (layer4_outputs(6839)));
    layer5_outputs(3858) <= not(layer4_outputs(6552));
    layer5_outputs(3859) <= not(layer4_outputs(2148));
    layer5_outputs(3860) <= not((layer4_outputs(5054)) or (layer4_outputs(6964)));
    layer5_outputs(3861) <= not((layer4_outputs(3006)) xor (layer4_outputs(6139)));
    layer5_outputs(3862) <= (layer4_outputs(1328)) xor (layer4_outputs(2302));
    layer5_outputs(3863) <= (layer4_outputs(2166)) and not (layer4_outputs(1877));
    layer5_outputs(3864) <= not(layer4_outputs(3453));
    layer5_outputs(3865) <= '0';
    layer5_outputs(3866) <= not(layer4_outputs(6676)) or (layer4_outputs(6929));
    layer5_outputs(3867) <= not(layer4_outputs(3783)) or (layer4_outputs(519));
    layer5_outputs(3868) <= layer4_outputs(2946);
    layer5_outputs(3869) <= not(layer4_outputs(1742));
    layer5_outputs(3870) <= not(layer4_outputs(2077));
    layer5_outputs(3871) <= layer4_outputs(1972);
    layer5_outputs(3872) <= not(layer4_outputs(2718));
    layer5_outputs(3873) <= not(layer4_outputs(5982));
    layer5_outputs(3874) <= (layer4_outputs(5448)) and not (layer4_outputs(7620));
    layer5_outputs(3875) <= (layer4_outputs(5254)) and not (layer4_outputs(2639));
    layer5_outputs(3876) <= not((layer4_outputs(3885)) and (layer4_outputs(6795)));
    layer5_outputs(3877) <= not(layer4_outputs(5986));
    layer5_outputs(3878) <= not(layer4_outputs(6953));
    layer5_outputs(3879) <= '1';
    layer5_outputs(3880) <= (layer4_outputs(3682)) and not (layer4_outputs(2996));
    layer5_outputs(3881) <= (layer4_outputs(5501)) and not (layer4_outputs(4201));
    layer5_outputs(3882) <= (layer4_outputs(4293)) and (layer4_outputs(2019));
    layer5_outputs(3883) <= layer4_outputs(4327);
    layer5_outputs(3884) <= (layer4_outputs(5528)) and not (layer4_outputs(4782));
    layer5_outputs(3885) <= layer4_outputs(605);
    layer5_outputs(3886) <= layer4_outputs(7125);
    layer5_outputs(3887) <= not((layer4_outputs(4150)) and (layer4_outputs(5457)));
    layer5_outputs(3888) <= layer4_outputs(5377);
    layer5_outputs(3889) <= layer4_outputs(3472);
    layer5_outputs(3890) <= (layer4_outputs(3565)) and not (layer4_outputs(573));
    layer5_outputs(3891) <= (layer4_outputs(7525)) or (layer4_outputs(483));
    layer5_outputs(3892) <= not(layer4_outputs(1490));
    layer5_outputs(3893) <= not(layer4_outputs(5860));
    layer5_outputs(3894) <= not((layer4_outputs(4464)) xor (layer4_outputs(1106)));
    layer5_outputs(3895) <= not(layer4_outputs(4546));
    layer5_outputs(3896) <= '0';
    layer5_outputs(3897) <= not((layer4_outputs(18)) xor (layer4_outputs(4858)));
    layer5_outputs(3898) <= not(layer4_outputs(7204)) or (layer4_outputs(6998));
    layer5_outputs(3899) <= not((layer4_outputs(124)) or (layer4_outputs(3937)));
    layer5_outputs(3900) <= (layer4_outputs(654)) or (layer4_outputs(1795));
    layer5_outputs(3901) <= not(layer4_outputs(1764));
    layer5_outputs(3902) <= layer4_outputs(3693);
    layer5_outputs(3903) <= (layer4_outputs(4644)) and not (layer4_outputs(3248));
    layer5_outputs(3904) <= not(layer4_outputs(4937));
    layer5_outputs(3905) <= not((layer4_outputs(5058)) or (layer4_outputs(3361)));
    layer5_outputs(3906) <= layer4_outputs(6696);
    layer5_outputs(3907) <= not(layer4_outputs(2473));
    layer5_outputs(3908) <= (layer4_outputs(5738)) and not (layer4_outputs(109));
    layer5_outputs(3909) <= not(layer4_outputs(7287)) or (layer4_outputs(6979));
    layer5_outputs(3910) <= layer4_outputs(4205);
    layer5_outputs(3911) <= not((layer4_outputs(212)) or (layer4_outputs(4829)));
    layer5_outputs(3912) <= layer4_outputs(656);
    layer5_outputs(3913) <= (layer4_outputs(7621)) and (layer4_outputs(3985));
    layer5_outputs(3914) <= not(layer4_outputs(4194));
    layer5_outputs(3915) <= not(layer4_outputs(4646));
    layer5_outputs(3916) <= layer4_outputs(3559);
    layer5_outputs(3917) <= (layer4_outputs(745)) and (layer4_outputs(2486));
    layer5_outputs(3918) <= (layer4_outputs(1960)) and not (layer4_outputs(7253));
    layer5_outputs(3919) <= not((layer4_outputs(7236)) or (layer4_outputs(3279)));
    layer5_outputs(3920) <= (layer4_outputs(2072)) xor (layer4_outputs(6086));
    layer5_outputs(3921) <= layer4_outputs(4502);
    layer5_outputs(3922) <= (layer4_outputs(1040)) xor (layer4_outputs(6108));
    layer5_outputs(3923) <= not((layer4_outputs(3090)) xor (layer4_outputs(6992)));
    layer5_outputs(3924) <= layer4_outputs(7586);
    layer5_outputs(3925) <= not(layer4_outputs(5584));
    layer5_outputs(3926) <= (layer4_outputs(1444)) xor (layer4_outputs(1431));
    layer5_outputs(3927) <= not((layer4_outputs(371)) xor (layer4_outputs(6195)));
    layer5_outputs(3928) <= not(layer4_outputs(3779));
    layer5_outputs(3929) <= not((layer4_outputs(319)) xor (layer4_outputs(3308)));
    layer5_outputs(3930) <= (layer4_outputs(3016)) and not (layer4_outputs(3666));
    layer5_outputs(3931) <= not((layer4_outputs(7484)) xor (layer4_outputs(4125)));
    layer5_outputs(3932) <= not(layer4_outputs(1405)) or (layer4_outputs(523));
    layer5_outputs(3933) <= (layer4_outputs(3332)) and not (layer4_outputs(2275));
    layer5_outputs(3934) <= not((layer4_outputs(2772)) xor (layer4_outputs(3268)));
    layer5_outputs(3935) <= not(layer4_outputs(1172));
    layer5_outputs(3936) <= layer4_outputs(839);
    layer5_outputs(3937) <= '0';
    layer5_outputs(3938) <= (layer4_outputs(1146)) or (layer4_outputs(4531));
    layer5_outputs(3939) <= not((layer4_outputs(7058)) xor (layer4_outputs(958)));
    layer5_outputs(3940) <= not((layer4_outputs(7244)) or (layer4_outputs(7126)));
    layer5_outputs(3941) <= not(layer4_outputs(5553));
    layer5_outputs(3942) <= layer4_outputs(410);
    layer5_outputs(3943) <= layer4_outputs(5102);
    layer5_outputs(3944) <= (layer4_outputs(5795)) and not (layer4_outputs(541));
    layer5_outputs(3945) <= not((layer4_outputs(6506)) or (layer4_outputs(7672)));
    layer5_outputs(3946) <= not((layer4_outputs(68)) or (layer4_outputs(4381)));
    layer5_outputs(3947) <= not((layer4_outputs(1667)) or (layer4_outputs(1130)));
    layer5_outputs(3948) <= layer4_outputs(4297);
    layer5_outputs(3949) <= layer4_outputs(6890);
    layer5_outputs(3950) <= not((layer4_outputs(1440)) and (layer4_outputs(5771)));
    layer5_outputs(3951) <= (layer4_outputs(5906)) xor (layer4_outputs(4375));
    layer5_outputs(3952) <= not((layer4_outputs(3607)) xor (layer4_outputs(2390)));
    layer5_outputs(3953) <= (layer4_outputs(6492)) and not (layer4_outputs(2894));
    layer5_outputs(3954) <= not(layer4_outputs(1327));
    layer5_outputs(3955) <= (layer4_outputs(2981)) and not (layer4_outputs(2303));
    layer5_outputs(3956) <= not((layer4_outputs(4519)) xor (layer4_outputs(1730)));
    layer5_outputs(3957) <= (layer4_outputs(7151)) and (layer4_outputs(2927));
    layer5_outputs(3958) <= not(layer4_outputs(2761));
    layer5_outputs(3959) <= layer4_outputs(4869);
    layer5_outputs(3960) <= (layer4_outputs(3848)) or (layer4_outputs(1451));
    layer5_outputs(3961) <= (layer4_outputs(5970)) and (layer4_outputs(2034));
    layer5_outputs(3962) <= (layer4_outputs(10)) and (layer4_outputs(2855));
    layer5_outputs(3963) <= not((layer4_outputs(5831)) and (layer4_outputs(6980)));
    layer5_outputs(3964) <= not(layer4_outputs(4160));
    layer5_outputs(3965) <= not(layer4_outputs(1625));
    layer5_outputs(3966) <= not((layer4_outputs(5582)) or (layer4_outputs(5854)));
    layer5_outputs(3967) <= not((layer4_outputs(1675)) or (layer4_outputs(541)));
    layer5_outputs(3968) <= layer4_outputs(6948);
    layer5_outputs(3969) <= not(layer4_outputs(2611));
    layer5_outputs(3970) <= not((layer4_outputs(6370)) xor (layer4_outputs(5977)));
    layer5_outputs(3971) <= '1';
    layer5_outputs(3972) <= '0';
    layer5_outputs(3973) <= layer4_outputs(2823);
    layer5_outputs(3974) <= (layer4_outputs(991)) and not (layer4_outputs(6120));
    layer5_outputs(3975) <= layer4_outputs(5427);
    layer5_outputs(3976) <= layer4_outputs(5443);
    layer5_outputs(3977) <= layer4_outputs(7470);
    layer5_outputs(3978) <= not((layer4_outputs(1354)) xor (layer4_outputs(5010)));
    layer5_outputs(3979) <= not((layer4_outputs(6816)) and (layer4_outputs(6333)));
    layer5_outputs(3980) <= layer4_outputs(7450);
    layer5_outputs(3981) <= (layer4_outputs(5278)) and not (layer4_outputs(3626));
    layer5_outputs(3982) <= (layer4_outputs(7275)) or (layer4_outputs(5389));
    layer5_outputs(3983) <= not(layer4_outputs(5900)) or (layer4_outputs(3829));
    layer5_outputs(3984) <= layer4_outputs(4633);
    layer5_outputs(3985) <= (layer4_outputs(5409)) and not (layer4_outputs(4260));
    layer5_outputs(3986) <= (layer4_outputs(2962)) and not (layer4_outputs(3623));
    layer5_outputs(3987) <= layer4_outputs(3441);
    layer5_outputs(3988) <= layer4_outputs(4834);
    layer5_outputs(3989) <= layer4_outputs(4797);
    layer5_outputs(3990) <= not((layer4_outputs(5565)) xor (layer4_outputs(1558)));
    layer5_outputs(3991) <= '0';
    layer5_outputs(3992) <= '1';
    layer5_outputs(3993) <= not((layer4_outputs(2615)) and (layer4_outputs(7117)));
    layer5_outputs(3994) <= layer4_outputs(5561);
    layer5_outputs(3995) <= layer4_outputs(6693);
    layer5_outputs(3996) <= not(layer4_outputs(312));
    layer5_outputs(3997) <= '1';
    layer5_outputs(3998) <= not(layer4_outputs(2099));
    layer5_outputs(3999) <= layer4_outputs(3645);
    layer5_outputs(4000) <= layer4_outputs(7394);
    layer5_outputs(4001) <= not(layer4_outputs(5201));
    layer5_outputs(4002) <= layer4_outputs(7540);
    layer5_outputs(4003) <= not(layer4_outputs(2036));
    layer5_outputs(4004) <= not(layer4_outputs(5418)) or (layer4_outputs(2959));
    layer5_outputs(4005) <= (layer4_outputs(3110)) and not (layer4_outputs(4083));
    layer5_outputs(4006) <= '1';
    layer5_outputs(4007) <= not((layer4_outputs(1881)) or (layer4_outputs(2729)));
    layer5_outputs(4008) <= layer4_outputs(3425);
    layer5_outputs(4009) <= layer4_outputs(3122);
    layer5_outputs(4010) <= layer4_outputs(5548);
    layer5_outputs(4011) <= layer4_outputs(7618);
    layer5_outputs(4012) <= not((layer4_outputs(5907)) xor (layer4_outputs(4660)));
    layer5_outputs(4013) <= (layer4_outputs(566)) or (layer4_outputs(1309));
    layer5_outputs(4014) <= not(layer4_outputs(4283)) or (layer4_outputs(1992));
    layer5_outputs(4015) <= (layer4_outputs(1770)) and not (layer4_outputs(4883));
    layer5_outputs(4016) <= layer4_outputs(7046);
    layer5_outputs(4017) <= (layer4_outputs(7661)) and (layer4_outputs(3567));
    layer5_outputs(4018) <= (layer4_outputs(4132)) or (layer4_outputs(6947));
    layer5_outputs(4019) <= '0';
    layer5_outputs(4020) <= (layer4_outputs(854)) and not (layer4_outputs(4651));
    layer5_outputs(4021) <= not(layer4_outputs(5628));
    layer5_outputs(4022) <= not(layer4_outputs(6449));
    layer5_outputs(4023) <= (layer4_outputs(4022)) and (layer4_outputs(1027));
    layer5_outputs(4024) <= layer4_outputs(7397);
    layer5_outputs(4025) <= not(layer4_outputs(2644));
    layer5_outputs(4026) <= layer4_outputs(3407);
    layer5_outputs(4027) <= (layer4_outputs(1905)) and not (layer4_outputs(4458));
    layer5_outputs(4028) <= layer4_outputs(5965);
    layer5_outputs(4029) <= layer4_outputs(6696);
    layer5_outputs(4030) <= not(layer4_outputs(7144));
    layer5_outputs(4031) <= layer4_outputs(3175);
    layer5_outputs(4032) <= not((layer4_outputs(6001)) and (layer4_outputs(2129)));
    layer5_outputs(4033) <= not(layer4_outputs(5536)) or (layer4_outputs(4687));
    layer5_outputs(4034) <= not(layer4_outputs(1041));
    layer5_outputs(4035) <= layer4_outputs(2598);
    layer5_outputs(4036) <= not(layer4_outputs(3071));
    layer5_outputs(4037) <= '0';
    layer5_outputs(4038) <= (layer4_outputs(904)) or (layer4_outputs(6611));
    layer5_outputs(4039) <= layer4_outputs(961);
    layer5_outputs(4040) <= not(layer4_outputs(137)) or (layer4_outputs(6561));
    layer5_outputs(4041) <= not(layer4_outputs(3783)) or (layer4_outputs(2660));
    layer5_outputs(4042) <= layer4_outputs(3572);
    layer5_outputs(4043) <= not((layer4_outputs(4035)) xor (layer4_outputs(6542)));
    layer5_outputs(4044) <= (layer4_outputs(3211)) and not (layer4_outputs(194));
    layer5_outputs(4045) <= not((layer4_outputs(2843)) and (layer4_outputs(6620)));
    layer5_outputs(4046) <= layer4_outputs(5583);
    layer5_outputs(4047) <= not((layer4_outputs(4978)) xor (layer4_outputs(1918)));
    layer5_outputs(4048) <= (layer4_outputs(4445)) xor (layer4_outputs(5669));
    layer5_outputs(4049) <= (layer4_outputs(6590)) or (layer4_outputs(7503));
    layer5_outputs(4050) <= (layer4_outputs(5905)) and not (layer4_outputs(3163));
    layer5_outputs(4051) <= (layer4_outputs(7660)) and (layer4_outputs(1854));
    layer5_outputs(4052) <= layer4_outputs(1488);
    layer5_outputs(4053) <= not((layer4_outputs(5916)) or (layer4_outputs(6123)));
    layer5_outputs(4054) <= (layer4_outputs(1381)) and not (layer4_outputs(4503));
    layer5_outputs(4055) <= (layer4_outputs(5394)) and not (layer4_outputs(6673));
    layer5_outputs(4056) <= layer4_outputs(1778);
    layer5_outputs(4057) <= not(layer4_outputs(6240)) or (layer4_outputs(94));
    layer5_outputs(4058) <= layer4_outputs(5284);
    layer5_outputs(4059) <= layer4_outputs(6030);
    layer5_outputs(4060) <= not(layer4_outputs(1573));
    layer5_outputs(4061) <= '1';
    layer5_outputs(4062) <= not(layer4_outputs(1312));
    layer5_outputs(4063) <= layer4_outputs(6335);
    layer5_outputs(4064) <= layer4_outputs(3771);
    layer5_outputs(4065) <= layer4_outputs(7005);
    layer5_outputs(4066) <= (layer4_outputs(6880)) xor (layer4_outputs(1562));
    layer5_outputs(4067) <= not(layer4_outputs(2230)) or (layer4_outputs(246));
    layer5_outputs(4068) <= not(layer4_outputs(4093));
    layer5_outputs(4069) <= (layer4_outputs(3167)) and (layer4_outputs(6484));
    layer5_outputs(4070) <= not(layer4_outputs(3306));
    layer5_outputs(4071) <= (layer4_outputs(1151)) and not (layer4_outputs(721));
    layer5_outputs(4072) <= (layer4_outputs(2931)) xor (layer4_outputs(2147));
    layer5_outputs(4073) <= layer4_outputs(3040);
    layer5_outputs(4074) <= not(layer4_outputs(4809));
    layer5_outputs(4075) <= '0';
    layer5_outputs(4076) <= (layer4_outputs(4715)) and not (layer4_outputs(110));
    layer5_outputs(4077) <= not((layer4_outputs(7571)) xor (layer4_outputs(5700)));
    layer5_outputs(4078) <= not(layer4_outputs(2323)) or (layer4_outputs(611));
    layer5_outputs(4079) <= (layer4_outputs(1746)) or (layer4_outputs(4277));
    layer5_outputs(4080) <= not((layer4_outputs(1275)) and (layer4_outputs(811)));
    layer5_outputs(4081) <= not((layer4_outputs(604)) or (layer4_outputs(7089)));
    layer5_outputs(4082) <= layer4_outputs(1398);
    layer5_outputs(4083) <= not((layer4_outputs(1620)) xor (layer4_outputs(7129)));
    layer5_outputs(4084) <= not((layer4_outputs(7409)) or (layer4_outputs(6327)));
    layer5_outputs(4085) <= (layer4_outputs(3870)) and not (layer4_outputs(5507));
    layer5_outputs(4086) <= not(layer4_outputs(7555));
    layer5_outputs(4087) <= layer4_outputs(3282);
    layer5_outputs(4088) <= (layer4_outputs(533)) xor (layer4_outputs(6503));
    layer5_outputs(4089) <= not(layer4_outputs(3612));
    layer5_outputs(4090) <= not(layer4_outputs(6169));
    layer5_outputs(4091) <= (layer4_outputs(4967)) or (layer4_outputs(5264));
    layer5_outputs(4092) <= not((layer4_outputs(5923)) or (layer4_outputs(4139)));
    layer5_outputs(4093) <= not(layer4_outputs(814)) or (layer4_outputs(7335));
    layer5_outputs(4094) <= (layer4_outputs(6604)) and not (layer4_outputs(6257));
    layer5_outputs(4095) <= not(layer4_outputs(2166));
    layer5_outputs(4096) <= layer4_outputs(3891);
    layer5_outputs(4097) <= not(layer4_outputs(7290));
    layer5_outputs(4098) <= not(layer4_outputs(7457));
    layer5_outputs(4099) <= (layer4_outputs(5823)) xor (layer4_outputs(2831));
    layer5_outputs(4100) <= layer4_outputs(5636);
    layer5_outputs(4101) <= (layer4_outputs(1684)) and not (layer4_outputs(333));
    layer5_outputs(4102) <= not(layer4_outputs(683)) or (layer4_outputs(6130));
    layer5_outputs(4103) <= layer4_outputs(7287);
    layer5_outputs(4104) <= layer4_outputs(2813);
    layer5_outputs(4105) <= layer4_outputs(5039);
    layer5_outputs(4106) <= layer4_outputs(3051);
    layer5_outputs(4107) <= (layer4_outputs(3969)) xor (layer4_outputs(3488));
    layer5_outputs(4108) <= layer4_outputs(6402);
    layer5_outputs(4109) <= not(layer4_outputs(4932));
    layer5_outputs(4110) <= not((layer4_outputs(5125)) xor (layer4_outputs(7443)));
    layer5_outputs(4111) <= not(layer4_outputs(6577));
    layer5_outputs(4112) <= layer4_outputs(2533);
    layer5_outputs(4113) <= layer4_outputs(4299);
    layer5_outputs(4114) <= not(layer4_outputs(2480));
    layer5_outputs(4115) <= not(layer4_outputs(2839));
    layer5_outputs(4116) <= layer4_outputs(5883);
    layer5_outputs(4117) <= (layer4_outputs(6558)) or (layer4_outputs(202));
    layer5_outputs(4118) <= not(layer4_outputs(820));
    layer5_outputs(4119) <= '0';
    layer5_outputs(4120) <= (layer4_outputs(4279)) and (layer4_outputs(2766));
    layer5_outputs(4121) <= (layer4_outputs(6361)) and not (layer4_outputs(2525));
    layer5_outputs(4122) <= (layer4_outputs(1668)) and not (layer4_outputs(6752));
    layer5_outputs(4123) <= not(layer4_outputs(5279));
    layer5_outputs(4124) <= (layer4_outputs(5810)) xor (layer4_outputs(4190));
    layer5_outputs(4125) <= not((layer4_outputs(753)) and (layer4_outputs(7589)));
    layer5_outputs(4126) <= not(layer4_outputs(932));
    layer5_outputs(4127) <= not((layer4_outputs(4835)) xor (layer4_outputs(1627)));
    layer5_outputs(4128) <= not(layer4_outputs(660));
    layer5_outputs(4129) <= (layer4_outputs(3581)) and not (layer4_outputs(4494));
    layer5_outputs(4130) <= '1';
    layer5_outputs(4131) <= not(layer4_outputs(174));
    layer5_outputs(4132) <= not(layer4_outputs(7221));
    layer5_outputs(4133) <= not(layer4_outputs(5326));
    layer5_outputs(4134) <= not((layer4_outputs(1566)) xor (layer4_outputs(2074)));
    layer5_outputs(4135) <= (layer4_outputs(1008)) and not (layer4_outputs(1739));
    layer5_outputs(4136) <= (layer4_outputs(3936)) xor (layer4_outputs(2834));
    layer5_outputs(4137) <= layer4_outputs(1532);
    layer5_outputs(4138) <= layer4_outputs(7155);
    layer5_outputs(4139) <= (layer4_outputs(4199)) and not (layer4_outputs(877));
    layer5_outputs(4140) <= (layer4_outputs(1839)) or (layer4_outputs(6554));
    layer5_outputs(4141) <= not((layer4_outputs(7493)) or (layer4_outputs(1495)));
    layer5_outputs(4142) <= not(layer4_outputs(657));
    layer5_outputs(4143) <= layer4_outputs(1555);
    layer5_outputs(4144) <= layer4_outputs(3281);
    layer5_outputs(4145) <= not((layer4_outputs(898)) and (layer4_outputs(1308)));
    layer5_outputs(4146) <= (layer4_outputs(6834)) and not (layer4_outputs(5857));
    layer5_outputs(4147) <= not(layer4_outputs(7309));
    layer5_outputs(4148) <= not(layer4_outputs(4792)) or (layer4_outputs(6628));
    layer5_outputs(4149) <= not((layer4_outputs(3173)) xor (layer4_outputs(4992)));
    layer5_outputs(4150) <= not(layer4_outputs(2783)) or (layer4_outputs(5245));
    layer5_outputs(4151) <= not(layer4_outputs(134));
    layer5_outputs(4152) <= layer4_outputs(6453);
    layer5_outputs(4153) <= not((layer4_outputs(6404)) or (layer4_outputs(492)));
    layer5_outputs(4154) <= not(layer4_outputs(19));
    layer5_outputs(4155) <= not(layer4_outputs(660));
    layer5_outputs(4156) <= not(layer4_outputs(3375)) or (layer4_outputs(307));
    layer5_outputs(4157) <= '0';
    layer5_outputs(4158) <= not((layer4_outputs(2256)) or (layer4_outputs(3782)));
    layer5_outputs(4159) <= not(layer4_outputs(92));
    layer5_outputs(4160) <= (layer4_outputs(2258)) and not (layer4_outputs(101));
    layer5_outputs(4161) <= not(layer4_outputs(5756));
    layer5_outputs(4162) <= (layer4_outputs(718)) xor (layer4_outputs(2989));
    layer5_outputs(4163) <= not(layer4_outputs(4329)) or (layer4_outputs(2555));
    layer5_outputs(4164) <= layer4_outputs(1240);
    layer5_outputs(4165) <= not(layer4_outputs(2803)) or (layer4_outputs(5099));
    layer5_outputs(4166) <= not(layer4_outputs(5598)) or (layer4_outputs(1913));
    layer5_outputs(4167) <= not(layer4_outputs(2196)) or (layer4_outputs(2869));
    layer5_outputs(4168) <= not(layer4_outputs(5346)) or (layer4_outputs(2870));
    layer5_outputs(4169) <= layer4_outputs(5493);
    layer5_outputs(4170) <= (layer4_outputs(1597)) and not (layer4_outputs(473));
    layer5_outputs(4171) <= layer4_outputs(5515);
    layer5_outputs(4172) <= (layer4_outputs(7389)) and (layer4_outputs(766));
    layer5_outputs(4173) <= layer4_outputs(1935);
    layer5_outputs(4174) <= not(layer4_outputs(7179));
    layer5_outputs(4175) <= '0';
    layer5_outputs(4176) <= not(layer4_outputs(558));
    layer5_outputs(4177) <= not(layer4_outputs(4557));
    layer5_outputs(4178) <= not(layer4_outputs(847));
    layer5_outputs(4179) <= layer4_outputs(3315);
    layer5_outputs(4180) <= layer4_outputs(6106);
    layer5_outputs(4181) <= layer4_outputs(283);
    layer5_outputs(4182) <= layer4_outputs(1136);
    layer5_outputs(4183) <= not(layer4_outputs(3596)) or (layer4_outputs(2237));
    layer5_outputs(4184) <= layer4_outputs(2878);
    layer5_outputs(4185) <= layer4_outputs(2789);
    layer5_outputs(4186) <= not((layer4_outputs(3151)) and (layer4_outputs(7578)));
    layer5_outputs(4187) <= not(layer4_outputs(7088)) or (layer4_outputs(3027));
    layer5_outputs(4188) <= layer4_outputs(7392);
    layer5_outputs(4189) <= layer4_outputs(1794);
    layer5_outputs(4190) <= not((layer4_outputs(2440)) xor (layer4_outputs(201)));
    layer5_outputs(4191) <= layer4_outputs(1737);
    layer5_outputs(4192) <= not(layer4_outputs(7567));
    layer5_outputs(4193) <= not(layer4_outputs(5725));
    layer5_outputs(4194) <= layer4_outputs(5901);
    layer5_outputs(4195) <= not(layer4_outputs(5924));
    layer5_outputs(4196) <= (layer4_outputs(4668)) or (layer4_outputs(3122));
    layer5_outputs(4197) <= layer4_outputs(4397);
    layer5_outputs(4198) <= layer4_outputs(2377);
    layer5_outputs(4199) <= not(layer4_outputs(2920));
    layer5_outputs(4200) <= not((layer4_outputs(457)) and (layer4_outputs(3334)));
    layer5_outputs(4201) <= not(layer4_outputs(1889));
    layer5_outputs(4202) <= not(layer4_outputs(6924));
    layer5_outputs(4203) <= not(layer4_outputs(4142));
    layer5_outputs(4204) <= not(layer4_outputs(5020));
    layer5_outputs(4205) <= not((layer4_outputs(1802)) or (layer4_outputs(2430)));
    layer5_outputs(4206) <= (layer4_outputs(7003)) and (layer4_outputs(6782));
    layer5_outputs(4207) <= not((layer4_outputs(2903)) xor (layer4_outputs(478)));
    layer5_outputs(4208) <= not((layer4_outputs(4507)) xor (layer4_outputs(1294)));
    layer5_outputs(4209) <= layer4_outputs(87);
    layer5_outputs(4210) <= not(layer4_outputs(3208)) or (layer4_outputs(2965));
    layer5_outputs(4211) <= layer4_outputs(3406);
    layer5_outputs(4212) <= layer4_outputs(4587);
    layer5_outputs(4213) <= layer4_outputs(314);
    layer5_outputs(4214) <= layer4_outputs(1613);
    layer5_outputs(4215) <= layer4_outputs(1869);
    layer5_outputs(4216) <= (layer4_outputs(4389)) and not (layer4_outputs(5721));
    layer5_outputs(4217) <= (layer4_outputs(7239)) xor (layer4_outputs(2683));
    layer5_outputs(4218) <= not((layer4_outputs(4662)) xor (layer4_outputs(5128)));
    layer5_outputs(4219) <= '1';
    layer5_outputs(4220) <= layer4_outputs(2906);
    layer5_outputs(4221) <= layer4_outputs(7643);
    layer5_outputs(4222) <= not(layer4_outputs(2605));
    layer5_outputs(4223) <= (layer4_outputs(3968)) and not (layer4_outputs(4735));
    layer5_outputs(4224) <= not(layer4_outputs(6061));
    layer5_outputs(4225) <= (layer4_outputs(1803)) and (layer4_outputs(6355));
    layer5_outputs(4226) <= layer4_outputs(6972);
    layer5_outputs(4227) <= not(layer4_outputs(3731)) or (layer4_outputs(4285));
    layer5_outputs(4228) <= (layer4_outputs(5127)) xor (layer4_outputs(6415));
    layer5_outputs(4229) <= not(layer4_outputs(7429));
    layer5_outputs(4230) <= (layer4_outputs(863)) and not (layer4_outputs(7528));
    layer5_outputs(4231) <= layer4_outputs(5337);
    layer5_outputs(4232) <= not(layer4_outputs(4784));
    layer5_outputs(4233) <= (layer4_outputs(3804)) or (layer4_outputs(5325));
    layer5_outputs(4234) <= not(layer4_outputs(842));
    layer5_outputs(4235) <= not(layer4_outputs(4126));
    layer5_outputs(4236) <= not(layer4_outputs(1229));
    layer5_outputs(4237) <= not(layer4_outputs(6079)) or (layer4_outputs(516));
    layer5_outputs(4238) <= (layer4_outputs(504)) xor (layer4_outputs(4140));
    layer5_outputs(4239) <= layer4_outputs(6343);
    layer5_outputs(4240) <= (layer4_outputs(4045)) and (layer4_outputs(1075));
    layer5_outputs(4241) <= not((layer4_outputs(1773)) and (layer4_outputs(4839)));
    layer5_outputs(4242) <= layer4_outputs(243);
    layer5_outputs(4243) <= not((layer4_outputs(5437)) xor (layer4_outputs(5509)));
    layer5_outputs(4244) <= not(layer4_outputs(4124));
    layer5_outputs(4245) <= not((layer4_outputs(419)) or (layer4_outputs(6085)));
    layer5_outputs(4246) <= layer4_outputs(7353);
    layer5_outputs(4247) <= layer4_outputs(3862);
    layer5_outputs(4248) <= not(layer4_outputs(4336)) or (layer4_outputs(7367));
    layer5_outputs(4249) <= not((layer4_outputs(1822)) or (layer4_outputs(7673)));
    layer5_outputs(4250) <= layer4_outputs(2681);
    layer5_outputs(4251) <= layer4_outputs(6123);
    layer5_outputs(4252) <= (layer4_outputs(2233)) or (layer4_outputs(4183));
    layer5_outputs(4253) <= layer4_outputs(4548);
    layer5_outputs(4254) <= not((layer4_outputs(4617)) xor (layer4_outputs(3789)));
    layer5_outputs(4255) <= layer4_outputs(3045);
    layer5_outputs(4256) <= layer4_outputs(401);
    layer5_outputs(4257) <= (layer4_outputs(2456)) or (layer4_outputs(1689));
    layer5_outputs(4258) <= (layer4_outputs(2663)) and not (layer4_outputs(1295));
    layer5_outputs(4259) <= not(layer4_outputs(1771));
    layer5_outputs(4260) <= not((layer4_outputs(5863)) xor (layer4_outputs(1089)));
    layer5_outputs(4261) <= not(layer4_outputs(621)) or (layer4_outputs(7407));
    layer5_outputs(4262) <= not(layer4_outputs(6633));
    layer5_outputs(4263) <= (layer4_outputs(6593)) and not (layer4_outputs(1305));
    layer5_outputs(4264) <= (layer4_outputs(5736)) xor (layer4_outputs(7256));
    layer5_outputs(4265) <= not(layer4_outputs(976));
    layer5_outputs(4266) <= layer4_outputs(4525);
    layer5_outputs(4267) <= not((layer4_outputs(1005)) and (layer4_outputs(4220)));
    layer5_outputs(4268) <= layer4_outputs(4642);
    layer5_outputs(4269) <= not(layer4_outputs(73));
    layer5_outputs(4270) <= not(layer4_outputs(6429)) or (layer4_outputs(6409));
    layer5_outputs(4271) <= not((layer4_outputs(1388)) xor (layer4_outputs(4995)));
    layer5_outputs(4272) <= (layer4_outputs(7276)) and not (layer4_outputs(3377));
    layer5_outputs(4273) <= not((layer4_outputs(2389)) and (layer4_outputs(5651)));
    layer5_outputs(4274) <= layer4_outputs(5303);
    layer5_outputs(4275) <= not((layer4_outputs(3751)) and (layer4_outputs(7143)));
    layer5_outputs(4276) <= layer4_outputs(164);
    layer5_outputs(4277) <= (layer4_outputs(3286)) xor (layer4_outputs(3984));
    layer5_outputs(4278) <= not(layer4_outputs(378));
    layer5_outputs(4279) <= not((layer4_outputs(2367)) xor (layer4_outputs(3052)));
    layer5_outputs(4280) <= layer4_outputs(7271);
    layer5_outputs(4281) <= layer4_outputs(278);
    layer5_outputs(4282) <= not(layer4_outputs(5370));
    layer5_outputs(4283) <= (layer4_outputs(4355)) and (layer4_outputs(3596));
    layer5_outputs(4284) <= not((layer4_outputs(2733)) or (layer4_outputs(3823)));
    layer5_outputs(4285) <= (layer4_outputs(5211)) and (layer4_outputs(6314));
    layer5_outputs(4286) <= not(layer4_outputs(7268));
    layer5_outputs(4287) <= (layer4_outputs(6041)) and (layer4_outputs(3065));
    layer5_outputs(4288) <= not((layer4_outputs(511)) or (layer4_outputs(7138)));
    layer5_outputs(4289) <= layer4_outputs(7340);
    layer5_outputs(4290) <= layer4_outputs(7268);
    layer5_outputs(4291) <= (layer4_outputs(1501)) and not (layer4_outputs(4740));
    layer5_outputs(4292) <= not(layer4_outputs(6818));
    layer5_outputs(4293) <= (layer4_outputs(5972)) and not (layer4_outputs(2455));
    layer5_outputs(4294) <= not((layer4_outputs(6481)) and (layer4_outputs(4516)));
    layer5_outputs(4295) <= (layer4_outputs(2492)) xor (layer4_outputs(4620));
    layer5_outputs(4296) <= layer4_outputs(2010);
    layer5_outputs(4297) <= (layer4_outputs(5071)) and (layer4_outputs(4222));
    layer5_outputs(4298) <= not(layer4_outputs(3971)) or (layer4_outputs(6213));
    layer5_outputs(4299) <= '0';
    layer5_outputs(4300) <= (layer4_outputs(6462)) xor (layer4_outputs(4400));
    layer5_outputs(4301) <= not((layer4_outputs(2420)) and (layer4_outputs(6399)));
    layer5_outputs(4302) <= not((layer4_outputs(4800)) and (layer4_outputs(5621)));
    layer5_outputs(4303) <= not(layer4_outputs(3303));
    layer5_outputs(4304) <= layer4_outputs(1115);
    layer5_outputs(4305) <= layer4_outputs(5995);
    layer5_outputs(4306) <= (layer4_outputs(3670)) or (layer4_outputs(1949));
    layer5_outputs(4307) <= not(layer4_outputs(6408));
    layer5_outputs(4308) <= not(layer4_outputs(7418));
    layer5_outputs(4309) <= layer4_outputs(6881);
    layer5_outputs(4310) <= layer4_outputs(7375);
    layer5_outputs(4311) <= layer4_outputs(7373);
    layer5_outputs(4312) <= not(layer4_outputs(780));
    layer5_outputs(4313) <= layer4_outputs(4906);
    layer5_outputs(4314) <= not((layer4_outputs(4338)) and (layer4_outputs(5742)));
    layer5_outputs(4315) <= (layer4_outputs(5772)) and (layer4_outputs(4616));
    layer5_outputs(4316) <= layer4_outputs(2963);
    layer5_outputs(4317) <= (layer4_outputs(5166)) and (layer4_outputs(4526));
    layer5_outputs(4318) <= not((layer4_outputs(861)) xor (layer4_outputs(7249)));
    layer5_outputs(4319) <= layer4_outputs(7511);
    layer5_outputs(4320) <= layer4_outputs(374);
    layer5_outputs(4321) <= (layer4_outputs(627)) or (layer4_outputs(2390));
    layer5_outputs(4322) <= layer4_outputs(6502);
    layer5_outputs(4323) <= not(layer4_outputs(5681));
    layer5_outputs(4324) <= layer4_outputs(6221);
    layer5_outputs(4325) <= (layer4_outputs(713)) xor (layer4_outputs(6092));
    layer5_outputs(4326) <= not(layer4_outputs(4170)) or (layer4_outputs(6661));
    layer5_outputs(4327) <= (layer4_outputs(4275)) and (layer4_outputs(6339));
    layer5_outputs(4328) <= not(layer4_outputs(2530));
    layer5_outputs(4329) <= layer4_outputs(175);
    layer5_outputs(4330) <= (layer4_outputs(506)) and not (layer4_outputs(594));
    layer5_outputs(4331) <= not(layer4_outputs(3970)) or (layer4_outputs(6514));
    layer5_outputs(4332) <= (layer4_outputs(3942)) and not (layer4_outputs(6493));
    layer5_outputs(4333) <= not(layer4_outputs(1059));
    layer5_outputs(4334) <= not((layer4_outputs(6645)) and (layer4_outputs(3428)));
    layer5_outputs(4335) <= layer4_outputs(458);
    layer5_outputs(4336) <= not((layer4_outputs(1000)) xor (layer4_outputs(7557)));
    layer5_outputs(4337) <= layer4_outputs(1532);
    layer5_outputs(4338) <= (layer4_outputs(5504)) and not (layer4_outputs(5228));
    layer5_outputs(4339) <= not((layer4_outputs(4057)) xor (layer4_outputs(5214)));
    layer5_outputs(4340) <= '0';
    layer5_outputs(4341) <= not(layer4_outputs(923)) or (layer4_outputs(5840));
    layer5_outputs(4342) <= '1';
    layer5_outputs(4343) <= not((layer4_outputs(4698)) or (layer4_outputs(1933)));
    layer5_outputs(4344) <= layer4_outputs(2880);
    layer5_outputs(4345) <= not((layer4_outputs(3780)) or (layer4_outputs(4238)));
    layer5_outputs(4346) <= (layer4_outputs(477)) and not (layer4_outputs(615));
    layer5_outputs(4347) <= layer4_outputs(4655);
    layer5_outputs(4348) <= layer4_outputs(5890);
    layer5_outputs(4349) <= not((layer4_outputs(7)) and (layer4_outputs(954)));
    layer5_outputs(4350) <= not(layer4_outputs(931));
    layer5_outputs(4351) <= layer4_outputs(6788);
    layer5_outputs(4352) <= not(layer4_outputs(5153));
    layer5_outputs(4353) <= layer4_outputs(4591);
    layer5_outputs(4354) <= (layer4_outputs(662)) and not (layer4_outputs(3092));
    layer5_outputs(4355) <= not((layer4_outputs(3161)) xor (layer4_outputs(4545)));
    layer5_outputs(4356) <= layer4_outputs(5195);
    layer5_outputs(4357) <= not(layer4_outputs(4737)) or (layer4_outputs(3876));
    layer5_outputs(4358) <= (layer4_outputs(7201)) and (layer4_outputs(484));
    layer5_outputs(4359) <= (layer4_outputs(1298)) or (layer4_outputs(2663));
    layer5_outputs(4360) <= not(layer4_outputs(2790));
    layer5_outputs(4361) <= not(layer4_outputs(2024)) or (layer4_outputs(6476));
    layer5_outputs(4362) <= layer4_outputs(4851);
    layer5_outputs(4363) <= not(layer4_outputs(562));
    layer5_outputs(4364) <= (layer4_outputs(6589)) and not (layer4_outputs(5780));
    layer5_outputs(4365) <= layer4_outputs(1636);
    layer5_outputs(4366) <= layer4_outputs(2408);
    layer5_outputs(4367) <= not((layer4_outputs(5704)) or (layer4_outputs(5164)));
    layer5_outputs(4368) <= not(layer4_outputs(2589));
    layer5_outputs(4369) <= (layer4_outputs(1713)) and not (layer4_outputs(624));
    layer5_outputs(4370) <= not(layer4_outputs(3351));
    layer5_outputs(4371) <= layer4_outputs(1072);
    layer5_outputs(4372) <= not((layer4_outputs(6443)) xor (layer4_outputs(63)));
    layer5_outputs(4373) <= layer4_outputs(4214);
    layer5_outputs(4374) <= not((layer4_outputs(4703)) or (layer4_outputs(113)));
    layer5_outputs(4375) <= (layer4_outputs(2279)) and (layer4_outputs(5534));
    layer5_outputs(4376) <= not(layer4_outputs(1359)) or (layer4_outputs(6830));
    layer5_outputs(4377) <= layer4_outputs(1843);
    layer5_outputs(4378) <= (layer4_outputs(4004)) and (layer4_outputs(2336));
    layer5_outputs(4379) <= layer4_outputs(2227);
    layer5_outputs(4380) <= (layer4_outputs(4979)) and not (layer4_outputs(4821));
    layer5_outputs(4381) <= (layer4_outputs(2452)) xor (layer4_outputs(3658));
    layer5_outputs(4382) <= (layer4_outputs(5390)) or (layer4_outputs(6378));
    layer5_outputs(4383) <= not(layer4_outputs(7512)) or (layer4_outputs(7065));
    layer5_outputs(4384) <= not((layer4_outputs(6280)) or (layer4_outputs(7523)));
    layer5_outputs(4385) <= not(layer4_outputs(254));
    layer5_outputs(4386) <= not(layer4_outputs(1789));
    layer5_outputs(4387) <= layer4_outputs(2400);
    layer5_outputs(4388) <= (layer4_outputs(2580)) and not (layer4_outputs(4049));
    layer5_outputs(4389) <= not((layer4_outputs(4557)) or (layer4_outputs(232)));
    layer5_outputs(4390) <= not(layer4_outputs(4410));
    layer5_outputs(4391) <= (layer4_outputs(6216)) and not (layer4_outputs(3618));
    layer5_outputs(4392) <= not(layer4_outputs(1302));
    layer5_outputs(4393) <= layer4_outputs(7318);
    layer5_outputs(4394) <= not(layer4_outputs(4041));
    layer5_outputs(4395) <= not((layer4_outputs(6216)) and (layer4_outputs(674)));
    layer5_outputs(4396) <= not((layer4_outputs(5388)) or (layer4_outputs(1469)));
    layer5_outputs(4397) <= not((layer4_outputs(7214)) or (layer4_outputs(7056)));
    layer5_outputs(4398) <= not((layer4_outputs(6157)) or (layer4_outputs(787)));
    layer5_outputs(4399) <= not(layer4_outputs(3368));
    layer5_outputs(4400) <= not(layer4_outputs(6735));
    layer5_outputs(4401) <= not(layer4_outputs(282));
    layer5_outputs(4402) <= (layer4_outputs(6956)) and not (layer4_outputs(6050));
    layer5_outputs(4403) <= not(layer4_outputs(6311)) or (layer4_outputs(4525));
    layer5_outputs(4404) <= (layer4_outputs(7458)) or (layer4_outputs(2059));
    layer5_outputs(4405) <= layer4_outputs(2171);
    layer5_outputs(4406) <= layer4_outputs(2974);
    layer5_outputs(4407) <= (layer4_outputs(5475)) xor (layer4_outputs(227));
    layer5_outputs(4408) <= not(layer4_outputs(1934));
    layer5_outputs(4409) <= layer4_outputs(6875);
    layer5_outputs(4410) <= (layer4_outputs(5562)) xor (layer4_outputs(4564));
    layer5_outputs(4411) <= (layer4_outputs(603)) or (layer4_outputs(5780));
    layer5_outputs(4412) <= not((layer4_outputs(4686)) xor (layer4_outputs(2391)));
    layer5_outputs(4413) <= not((layer4_outputs(3635)) xor (layer4_outputs(5309)));
    layer5_outputs(4414) <= layer4_outputs(5797);
    layer5_outputs(4415) <= not(layer4_outputs(644));
    layer5_outputs(4416) <= not(layer4_outputs(1881));
    layer5_outputs(4417) <= layer4_outputs(6962);
    layer5_outputs(4418) <= layer4_outputs(3377);
    layer5_outputs(4419) <= not((layer4_outputs(4615)) and (layer4_outputs(5203)));
    layer5_outputs(4420) <= not(layer4_outputs(360));
    layer5_outputs(4421) <= layer4_outputs(3586);
    layer5_outputs(4422) <= not((layer4_outputs(861)) or (layer4_outputs(3665)));
    layer5_outputs(4423) <= (layer4_outputs(5783)) and not (layer4_outputs(700));
    layer5_outputs(4424) <= not(layer4_outputs(5941));
    layer5_outputs(4425) <= not(layer4_outputs(7447)) or (layer4_outputs(5467));
    layer5_outputs(4426) <= not(layer4_outputs(571));
    layer5_outputs(4427) <= (layer4_outputs(263)) and not (layer4_outputs(3696));
    layer5_outputs(4428) <= not(layer4_outputs(3857));
    layer5_outputs(4429) <= not(layer4_outputs(5031));
    layer5_outputs(4430) <= not(layer4_outputs(4300));
    layer5_outputs(4431) <= '1';
    layer5_outputs(4432) <= layer4_outputs(6371);
    layer5_outputs(4433) <= (layer4_outputs(3072)) xor (layer4_outputs(77));
    layer5_outputs(4434) <= (layer4_outputs(3494)) and (layer4_outputs(1894));
    layer5_outputs(4435) <= layer4_outputs(1284);
    layer5_outputs(4436) <= (layer4_outputs(5127)) or (layer4_outputs(6888));
    layer5_outputs(4437) <= not(layer4_outputs(6000));
    layer5_outputs(4438) <= not(layer4_outputs(4864)) or (layer4_outputs(6719));
    layer5_outputs(4439) <= layer4_outputs(169);
    layer5_outputs(4440) <= not((layer4_outputs(4127)) or (layer4_outputs(5464)));
    layer5_outputs(4441) <= not(layer4_outputs(7583));
    layer5_outputs(4442) <= '0';
    layer5_outputs(4443) <= (layer4_outputs(1024)) or (layer4_outputs(6494));
    layer5_outputs(4444) <= layer4_outputs(5963);
    layer5_outputs(4445) <= not(layer4_outputs(4923));
    layer5_outputs(4446) <= layer4_outputs(4187);
    layer5_outputs(4447) <= (layer4_outputs(3465)) or (layer4_outputs(5331));
    layer5_outputs(4448) <= layer4_outputs(1977);
    layer5_outputs(4449) <= not(layer4_outputs(259));
    layer5_outputs(4450) <= layer4_outputs(7425);
    layer5_outputs(4451) <= layer4_outputs(4835);
    layer5_outputs(4452) <= not((layer4_outputs(1290)) and (layer4_outputs(259)));
    layer5_outputs(4453) <= not((layer4_outputs(3639)) xor (layer4_outputs(391)));
    layer5_outputs(4454) <= not(layer4_outputs(834));
    layer5_outputs(4455) <= not(layer4_outputs(2655)) or (layer4_outputs(482));
    layer5_outputs(4456) <= not(layer4_outputs(4223));
    layer5_outputs(4457) <= layer4_outputs(763);
    layer5_outputs(4458) <= not(layer4_outputs(7188));
    layer5_outputs(4459) <= layer4_outputs(2609);
    layer5_outputs(4460) <= '1';
    layer5_outputs(4461) <= layer4_outputs(5078);
    layer5_outputs(4462) <= not(layer4_outputs(3622));
    layer5_outputs(4463) <= layer4_outputs(4739);
    layer5_outputs(4464) <= layer4_outputs(6406);
    layer5_outputs(4465) <= not(layer4_outputs(3087)) or (layer4_outputs(5477));
    layer5_outputs(4466) <= not((layer4_outputs(2227)) xor (layer4_outputs(211)));
    layer5_outputs(4467) <= not(layer4_outputs(7126));
    layer5_outputs(4468) <= not(layer4_outputs(238)) or (layer4_outputs(6186));
    layer5_outputs(4469) <= layer4_outputs(7260);
    layer5_outputs(4470) <= not(layer4_outputs(27));
    layer5_outputs(4471) <= (layer4_outputs(6757)) and (layer4_outputs(520));
    layer5_outputs(4472) <= not(layer4_outputs(937));
    layer5_outputs(4473) <= not(layer4_outputs(6189)) or (layer4_outputs(5246));
    layer5_outputs(4474) <= (layer4_outputs(6072)) or (layer4_outputs(3919));
    layer5_outputs(4475) <= layer4_outputs(5478);
    layer5_outputs(4476) <= (layer4_outputs(1894)) xor (layer4_outputs(5195));
    layer5_outputs(4477) <= layer4_outputs(5336);
    layer5_outputs(4478) <= layer4_outputs(3389);
    layer5_outputs(4479) <= layer4_outputs(2445);
    layer5_outputs(4480) <= not((layer4_outputs(4989)) or (layer4_outputs(3870)));
    layer5_outputs(4481) <= not(layer4_outputs(1958));
    layer5_outputs(4482) <= (layer4_outputs(2454)) xor (layer4_outputs(3839));
    layer5_outputs(4483) <= layer4_outputs(3712);
    layer5_outputs(4484) <= (layer4_outputs(3895)) and (layer4_outputs(2422));
    layer5_outputs(4485) <= not(layer4_outputs(4313));
    layer5_outputs(4486) <= not((layer4_outputs(1689)) and (layer4_outputs(1614)));
    layer5_outputs(4487) <= not(layer4_outputs(459));
    layer5_outputs(4488) <= layer4_outputs(4073);
    layer5_outputs(4489) <= (layer4_outputs(7395)) xor (layer4_outputs(3482));
    layer5_outputs(4490) <= not(layer4_outputs(1334));
    layer5_outputs(4491) <= not(layer4_outputs(6498));
    layer5_outputs(4492) <= layer4_outputs(1233);
    layer5_outputs(4493) <= not(layer4_outputs(7082));
    layer5_outputs(4494) <= not(layer4_outputs(5981));
    layer5_outputs(4495) <= not(layer4_outputs(1342));
    layer5_outputs(4496) <= layer4_outputs(949);
    layer5_outputs(4497) <= layer4_outputs(7470);
    layer5_outputs(4498) <= '0';
    layer5_outputs(4499) <= (layer4_outputs(4356)) or (layer4_outputs(5662));
    layer5_outputs(4500) <= layer4_outputs(6099);
    layer5_outputs(4501) <= not(layer4_outputs(4371));
    layer5_outputs(4502) <= layer4_outputs(6045);
    layer5_outputs(4503) <= layer4_outputs(4491);
    layer5_outputs(4504) <= layer4_outputs(3524);
    layer5_outputs(4505) <= (layer4_outputs(7254)) xor (layer4_outputs(2662));
    layer5_outputs(4506) <= not(layer4_outputs(5702));
    layer5_outputs(4507) <= not(layer4_outputs(6533));
    layer5_outputs(4508) <= not((layer4_outputs(3577)) xor (layer4_outputs(5888)));
    layer5_outputs(4509) <= (layer4_outputs(4189)) and (layer4_outputs(2434));
    layer5_outputs(4510) <= '1';
    layer5_outputs(4511) <= not(layer4_outputs(5191));
    layer5_outputs(4512) <= layer4_outputs(6082);
    layer5_outputs(4513) <= not(layer4_outputs(4487)) or (layer4_outputs(4742));
    layer5_outputs(4514) <= '0';
    layer5_outputs(4515) <= layer4_outputs(6461);
    layer5_outputs(4516) <= layer4_outputs(7606);
    layer5_outputs(4517) <= not((layer4_outputs(3551)) or (layer4_outputs(1310)));
    layer5_outputs(4518) <= layer4_outputs(3487);
    layer5_outputs(4519) <= (layer4_outputs(1257)) and not (layer4_outputs(6906));
    layer5_outputs(4520) <= not((layer4_outputs(5537)) xor (layer4_outputs(598)));
    layer5_outputs(4521) <= not(layer4_outputs(255)) or (layer4_outputs(6197));
    layer5_outputs(4522) <= layer4_outputs(2026);
    layer5_outputs(4523) <= layer4_outputs(7184);
    layer5_outputs(4524) <= not(layer4_outputs(4376));
    layer5_outputs(4525) <= not(layer4_outputs(3222)) or (layer4_outputs(3509));
    layer5_outputs(4526) <= not(layer4_outputs(6441));
    layer5_outputs(4527) <= not(layer4_outputs(5999));
    layer5_outputs(4528) <= not(layer4_outputs(2053));
    layer5_outputs(4529) <= layer4_outputs(3709);
    layer5_outputs(4530) <= (layer4_outputs(4405)) and not (layer4_outputs(3408));
    layer5_outputs(4531) <= not(layer4_outputs(3460));
    layer5_outputs(4532) <= layer4_outputs(1518);
    layer5_outputs(4533) <= (layer4_outputs(6173)) and (layer4_outputs(7109));
    layer5_outputs(4534) <= not((layer4_outputs(3420)) and (layer4_outputs(6874)));
    layer5_outputs(4535) <= not(layer4_outputs(1483));
    layer5_outputs(4536) <= not(layer4_outputs(432));
    layer5_outputs(4537) <= not((layer4_outputs(7061)) or (layer4_outputs(6816)));
    layer5_outputs(4538) <= not(layer4_outputs(5305)) or (layer4_outputs(2447));
    layer5_outputs(4539) <= not(layer4_outputs(1454));
    layer5_outputs(4540) <= not(layer4_outputs(7623));
    layer5_outputs(4541) <= not(layer4_outputs(6967));
    layer5_outputs(4542) <= not(layer4_outputs(7076));
    layer5_outputs(4543) <= layer4_outputs(800);
    layer5_outputs(4544) <= not(layer4_outputs(3672));
    layer5_outputs(4545) <= not(layer4_outputs(5266));
    layer5_outputs(4546) <= layer4_outputs(1767);
    layer5_outputs(4547) <= (layer4_outputs(2208)) xor (layer4_outputs(1867));
    layer5_outputs(4548) <= not(layer4_outputs(4747));
    layer5_outputs(4549) <= not(layer4_outputs(121));
    layer5_outputs(4550) <= layer4_outputs(7378);
    layer5_outputs(4551) <= layer4_outputs(2727);
    layer5_outputs(4552) <= not(layer4_outputs(5307));
    layer5_outputs(4553) <= layer4_outputs(2323);
    layer5_outputs(4554) <= layer4_outputs(2571);
    layer5_outputs(4555) <= layer4_outputs(5301);
    layer5_outputs(4556) <= layer4_outputs(3789);
    layer5_outputs(4557) <= not(layer4_outputs(143)) or (layer4_outputs(5988));
    layer5_outputs(4558) <= layer4_outputs(1683);
    layer5_outputs(4559) <= layer4_outputs(3125);
    layer5_outputs(4560) <= not((layer4_outputs(3384)) and (layer4_outputs(76)));
    layer5_outputs(4561) <= not(layer4_outputs(4883)) or (layer4_outputs(5047));
    layer5_outputs(4562) <= not((layer4_outputs(3275)) and (layer4_outputs(3444)));
    layer5_outputs(4563) <= not(layer4_outputs(5207)) or (layer4_outputs(7400));
    layer5_outputs(4564) <= layer4_outputs(7370);
    layer5_outputs(4565) <= not((layer4_outputs(6048)) and (layer4_outputs(5779)));
    layer5_outputs(4566) <= not((layer4_outputs(3593)) and (layer4_outputs(3599)));
    layer5_outputs(4567) <= (layer4_outputs(4065)) xor (layer4_outputs(3301));
    layer5_outputs(4568) <= (layer4_outputs(400)) and not (layer4_outputs(2509));
    layer5_outputs(4569) <= not(layer4_outputs(167));
    layer5_outputs(4570) <= (layer4_outputs(2192)) and not (layer4_outputs(6455));
    layer5_outputs(4571) <= (layer4_outputs(7474)) xor (layer4_outputs(1176));
    layer5_outputs(4572) <= (layer4_outputs(6473)) and not (layer4_outputs(3196));
    layer5_outputs(4573) <= not((layer4_outputs(4221)) xor (layer4_outputs(4719)));
    layer5_outputs(4574) <= not(layer4_outputs(2608)) or (layer4_outputs(6294));
    layer5_outputs(4575) <= not(layer4_outputs(1177)) or (layer4_outputs(3439));
    layer5_outputs(4576) <= not(layer4_outputs(878));
    layer5_outputs(4577) <= not(layer4_outputs(2742));
    layer5_outputs(4578) <= layer4_outputs(4197);
    layer5_outputs(4579) <= not(layer4_outputs(4943));
    layer5_outputs(4580) <= not((layer4_outputs(6414)) xor (layer4_outputs(7030)));
    layer5_outputs(4581) <= not((layer4_outputs(6883)) and (layer4_outputs(1460)));
    layer5_outputs(4582) <= (layer4_outputs(7419)) and not (layer4_outputs(5396));
    layer5_outputs(4583) <= not(layer4_outputs(6584));
    layer5_outputs(4584) <= not(layer4_outputs(2954)) or (layer4_outputs(4498));
    layer5_outputs(4585) <= (layer4_outputs(5115)) and not (layer4_outputs(608));
    layer5_outputs(4586) <= not(layer4_outputs(3812)) or (layer4_outputs(1387));
    layer5_outputs(4587) <= not(layer4_outputs(4527));
    layer5_outputs(4588) <= layer4_outputs(1984);
    layer5_outputs(4589) <= layer4_outputs(6351);
    layer5_outputs(4590) <= (layer4_outputs(1660)) and not (layer4_outputs(2887));
    layer5_outputs(4591) <= layer4_outputs(2069);
    layer5_outputs(4592) <= layer4_outputs(7551);
    layer5_outputs(4593) <= layer4_outputs(5597);
    layer5_outputs(4594) <= layer4_outputs(180);
    layer5_outputs(4595) <= not(layer4_outputs(6657));
    layer5_outputs(4596) <= layer4_outputs(1177);
    layer5_outputs(4597) <= layer4_outputs(5165);
    layer5_outputs(4598) <= layer4_outputs(3012);
    layer5_outputs(4599) <= not(layer4_outputs(5803));
    layer5_outputs(4600) <= (layer4_outputs(23)) or (layer4_outputs(1310));
    layer5_outputs(4601) <= not((layer4_outputs(3946)) xor (layer4_outputs(4353)));
    layer5_outputs(4602) <= not((layer4_outputs(4239)) or (layer4_outputs(2912)));
    layer5_outputs(4603) <= (layer4_outputs(5603)) and not (layer4_outputs(3982));
    layer5_outputs(4604) <= not((layer4_outputs(3437)) xor (layer4_outputs(1002)));
    layer5_outputs(4605) <= not(layer4_outputs(7160));
    layer5_outputs(4606) <= (layer4_outputs(1062)) or (layer4_outputs(4748));
    layer5_outputs(4607) <= layer4_outputs(4636);
    layer5_outputs(4608) <= layer4_outputs(7454);
    layer5_outputs(4609) <= layer4_outputs(155);
    layer5_outputs(4610) <= (layer4_outputs(2489)) and (layer4_outputs(6440));
    layer5_outputs(4611) <= not(layer4_outputs(4647));
    layer5_outputs(4612) <= (layer4_outputs(3311)) and not (layer4_outputs(525));
    layer5_outputs(4613) <= layer4_outputs(60);
    layer5_outputs(4614) <= (layer4_outputs(4251)) or (layer4_outputs(6938));
    layer5_outputs(4615) <= not(layer4_outputs(2217)) or (layer4_outputs(2391));
    layer5_outputs(4616) <= not(layer4_outputs(2184));
    layer5_outputs(4617) <= not(layer4_outputs(6689));
    layer5_outputs(4618) <= layer4_outputs(3622);
    layer5_outputs(4619) <= layer4_outputs(3794);
    layer5_outputs(4620) <= (layer4_outputs(4477)) and not (layer4_outputs(2487));
    layer5_outputs(4621) <= layer4_outputs(2426);
    layer5_outputs(4622) <= not(layer4_outputs(298));
    layer5_outputs(4623) <= (layer4_outputs(7588)) and not (layer4_outputs(4928));
    layer5_outputs(4624) <= not(layer4_outputs(4133));
    layer5_outputs(4625) <= layer4_outputs(70);
    layer5_outputs(4626) <= not(layer4_outputs(4965));
    layer5_outputs(4627) <= (layer4_outputs(5758)) and (layer4_outputs(5553));
    layer5_outputs(4628) <= layer4_outputs(5589);
    layer5_outputs(4629) <= not(layer4_outputs(3142));
    layer5_outputs(4630) <= layer4_outputs(245);
    layer5_outputs(4631) <= not(layer4_outputs(2467));
    layer5_outputs(4632) <= not(layer4_outputs(4318));
    layer5_outputs(4633) <= layer4_outputs(7580);
    layer5_outputs(4634) <= layer4_outputs(6437);
    layer5_outputs(4635) <= not(layer4_outputs(5052));
    layer5_outputs(4636) <= (layer4_outputs(5118)) and not (layer4_outputs(7534));
    layer5_outputs(4637) <= not(layer4_outputs(5954));
    layer5_outputs(4638) <= layer4_outputs(2061);
    layer5_outputs(4639) <= layer4_outputs(4904);
    layer5_outputs(4640) <= (layer4_outputs(2980)) and (layer4_outputs(313));
    layer5_outputs(4641) <= not(layer4_outputs(7450)) or (layer4_outputs(5118));
    layer5_outputs(4642) <= not((layer4_outputs(7509)) xor (layer4_outputs(3836)));
    layer5_outputs(4643) <= '1';
    layer5_outputs(4644) <= (layer4_outputs(7216)) and (layer4_outputs(1411));
    layer5_outputs(4645) <= not(layer4_outputs(883));
    layer5_outputs(4646) <= not(layer4_outputs(2018)) or (layer4_outputs(6908));
    layer5_outputs(4647) <= (layer4_outputs(561)) or (layer4_outputs(203));
    layer5_outputs(4648) <= layer4_outputs(4670);
    layer5_outputs(4649) <= not((layer4_outputs(3462)) and (layer4_outputs(307)));
    layer5_outputs(4650) <= layer4_outputs(5500);
    layer5_outputs(4651) <= layer4_outputs(5751);
    layer5_outputs(4652) <= layer4_outputs(3731);
    layer5_outputs(4653) <= (layer4_outputs(999)) or (layer4_outputs(683));
    layer5_outputs(4654) <= (layer4_outputs(2909)) xor (layer4_outputs(5710));
    layer5_outputs(4655) <= layer4_outputs(6354);
    layer5_outputs(4656) <= not(layer4_outputs(3240));
    layer5_outputs(4657) <= layer4_outputs(4478);
    layer5_outputs(4658) <= not(layer4_outputs(399));
    layer5_outputs(4659) <= not(layer4_outputs(2700));
    layer5_outputs(4660) <= (layer4_outputs(3721)) and not (layer4_outputs(6901));
    layer5_outputs(4661) <= not(layer4_outputs(2382));
    layer5_outputs(4662) <= not((layer4_outputs(1857)) and (layer4_outputs(787)));
    layer5_outputs(4663) <= not(layer4_outputs(6405));
    layer5_outputs(4664) <= (layer4_outputs(3364)) and not (layer4_outputs(7507));
    layer5_outputs(4665) <= layer4_outputs(5401);
    layer5_outputs(4666) <= layer4_outputs(5102);
    layer5_outputs(4667) <= not(layer4_outputs(6935)) or (layer4_outputs(5347));
    layer5_outputs(4668) <= (layer4_outputs(4397)) or (layer4_outputs(3309));
    layer5_outputs(4669) <= layer4_outputs(2666);
    layer5_outputs(4670) <= not(layer4_outputs(1618));
    layer5_outputs(4671) <= layer4_outputs(6128);
    layer5_outputs(4672) <= (layer4_outputs(5622)) and (layer4_outputs(3950));
    layer5_outputs(4673) <= not(layer4_outputs(6640)) or (layer4_outputs(2152));
    layer5_outputs(4674) <= (layer4_outputs(4044)) and not (layer4_outputs(6200));
    layer5_outputs(4675) <= not((layer4_outputs(5604)) and (layer4_outputs(5456)));
    layer5_outputs(4676) <= not(layer4_outputs(4237));
    layer5_outputs(4677) <= layer4_outputs(3224);
    layer5_outputs(4678) <= layer4_outputs(6942);
    layer5_outputs(4679) <= not((layer4_outputs(6472)) or (layer4_outputs(2991)));
    layer5_outputs(4680) <= not(layer4_outputs(1249)) or (layer4_outputs(3458));
    layer5_outputs(4681) <= layer4_outputs(7602);
    layer5_outputs(4682) <= not(layer4_outputs(6084));
    layer5_outputs(4683) <= not(layer4_outputs(3918)) or (layer4_outputs(6326));
    layer5_outputs(4684) <= '1';
    layer5_outputs(4685) <= layer4_outputs(4888);
    layer5_outputs(4686) <= layer4_outputs(890);
    layer5_outputs(4687) <= (layer4_outputs(5430)) and not (layer4_outputs(7327));
    layer5_outputs(4688) <= not(layer4_outputs(2747));
    layer5_outputs(4689) <= layer4_outputs(1662);
    layer5_outputs(4690) <= not((layer4_outputs(869)) and (layer4_outputs(4315)));
    layer5_outputs(4691) <= not(layer4_outputs(6293));
    layer5_outputs(4692) <= layer4_outputs(3679);
    layer5_outputs(4693) <= layer4_outputs(4227);
    layer5_outputs(4694) <= not((layer4_outputs(1380)) or (layer4_outputs(6316)));
    layer5_outputs(4695) <= (layer4_outputs(6346)) xor (layer4_outputs(2685));
    layer5_outputs(4696) <= not(layer4_outputs(5295));
    layer5_outputs(4697) <= (layer4_outputs(4949)) and not (layer4_outputs(2498));
    layer5_outputs(4698) <= layer4_outputs(7215);
    layer5_outputs(4699) <= not(layer4_outputs(3754));
    layer5_outputs(4700) <= not(layer4_outputs(2291));
    layer5_outputs(4701) <= (layer4_outputs(7513)) xor (layer4_outputs(1494));
    layer5_outputs(4702) <= layer4_outputs(1824);
    layer5_outputs(4703) <= layer4_outputs(3461);
    layer5_outputs(4704) <= '0';
    layer5_outputs(4705) <= '1';
    layer5_outputs(4706) <= layer4_outputs(1889);
    layer5_outputs(4707) <= layer4_outputs(3605);
    layer5_outputs(4708) <= (layer4_outputs(2750)) and (layer4_outputs(5912));
    layer5_outputs(4709) <= layer4_outputs(3458);
    layer5_outputs(4710) <= not(layer4_outputs(2366));
    layer5_outputs(4711) <= layer4_outputs(6853);
    layer5_outputs(4712) <= (layer4_outputs(5177)) xor (layer4_outputs(6729));
    layer5_outputs(4713) <= layer4_outputs(5074);
    layer5_outputs(4714) <= not((layer4_outputs(1761)) or (layer4_outputs(2441)));
    layer5_outputs(4715) <= '1';
    layer5_outputs(4716) <= (layer4_outputs(783)) and (layer4_outputs(131));
    layer5_outputs(4717) <= not(layer4_outputs(4421));
    layer5_outputs(4718) <= (layer4_outputs(6416)) and (layer4_outputs(3038));
    layer5_outputs(4719) <= not(layer4_outputs(4094));
    layer5_outputs(4720) <= layer4_outputs(3290);
    layer5_outputs(4721) <= not(layer4_outputs(2324));
    layer5_outputs(4722) <= layer4_outputs(3833);
    layer5_outputs(4723) <= (layer4_outputs(4312)) and (layer4_outputs(3444));
    layer5_outputs(4724) <= (layer4_outputs(3746)) or (layer4_outputs(6192));
    layer5_outputs(4725) <= (layer4_outputs(1228)) and not (layer4_outputs(2255));
    layer5_outputs(4726) <= not(layer4_outputs(7367));
    layer5_outputs(4727) <= (layer4_outputs(1122)) xor (layer4_outputs(5657));
    layer5_outputs(4728) <= layer4_outputs(6846);
    layer5_outputs(4729) <= not(layer4_outputs(7010));
    layer5_outputs(4730) <= (layer4_outputs(6218)) xor (layer4_outputs(5694));
    layer5_outputs(4731) <= not(layer4_outputs(181)) or (layer4_outputs(5760));
    layer5_outputs(4732) <= not((layer4_outputs(3049)) xor (layer4_outputs(2079)));
    layer5_outputs(4733) <= layer4_outputs(4285);
    layer5_outputs(4734) <= (layer4_outputs(3911)) and not (layer4_outputs(6867));
    layer5_outputs(4735) <= layer4_outputs(7079);
    layer5_outputs(4736) <= not(layer4_outputs(1664));
    layer5_outputs(4737) <= layer4_outputs(3225);
    layer5_outputs(4738) <= not(layer4_outputs(2524));
    layer5_outputs(4739) <= layer4_outputs(2642);
    layer5_outputs(4740) <= (layer4_outputs(4794)) and not (layer4_outputs(3728));
    layer5_outputs(4741) <= not(layer4_outputs(5160));
    layer5_outputs(4742) <= not(layer4_outputs(2071));
    layer5_outputs(4743) <= not(layer4_outputs(5913)) or (layer4_outputs(6970));
    layer5_outputs(4744) <= not(layer4_outputs(6287));
    layer5_outputs(4745) <= not(layer4_outputs(2754));
    layer5_outputs(4746) <= not(layer4_outputs(4440));
    layer5_outputs(4747) <= (layer4_outputs(6475)) or (layer4_outputs(2988));
    layer5_outputs(4748) <= not(layer4_outputs(3867));
    layer5_outputs(4749) <= not(layer4_outputs(1736));
    layer5_outputs(4750) <= not((layer4_outputs(2470)) xor (layer4_outputs(6300)));
    layer5_outputs(4751) <= not(layer4_outputs(6104));
    layer5_outputs(4752) <= (layer4_outputs(2163)) and not (layer4_outputs(442));
    layer5_outputs(4753) <= (layer4_outputs(2711)) or (layer4_outputs(7565));
    layer5_outputs(4754) <= not((layer4_outputs(3619)) and (layer4_outputs(198)));
    layer5_outputs(4755) <= not(layer4_outputs(1954));
    layer5_outputs(4756) <= layer4_outputs(4924);
    layer5_outputs(4757) <= (layer4_outputs(6235)) and (layer4_outputs(2689));
    layer5_outputs(4758) <= not((layer4_outputs(2848)) and (layer4_outputs(3706)));
    layer5_outputs(4759) <= not(layer4_outputs(1830));
    layer5_outputs(4760) <= (layer4_outputs(6109)) and not (layer4_outputs(3973));
    layer5_outputs(4761) <= (layer4_outputs(3456)) and not (layer4_outputs(4894));
    layer5_outputs(4762) <= not((layer4_outputs(2088)) and (layer4_outputs(2583)));
    layer5_outputs(4763) <= not((layer4_outputs(74)) xor (layer4_outputs(7573)));
    layer5_outputs(4764) <= layer4_outputs(7354);
    layer5_outputs(4765) <= layer4_outputs(6469);
    layer5_outputs(4766) <= not((layer4_outputs(5589)) and (layer4_outputs(7180)));
    layer5_outputs(4767) <= layer4_outputs(2827);
    layer5_outputs(4768) <= not(layer4_outputs(4998)) or (layer4_outputs(8));
    layer5_outputs(4769) <= (layer4_outputs(7289)) and (layer4_outputs(7039));
    layer5_outputs(4770) <= not(layer4_outputs(4508));
    layer5_outputs(4771) <= not(layer4_outputs(2667));
    layer5_outputs(4772) <= '1';
    layer5_outputs(4773) <= (layer4_outputs(6274)) and not (layer4_outputs(6783));
    layer5_outputs(4774) <= not((layer4_outputs(4652)) xor (layer4_outputs(7270)));
    layer5_outputs(4775) <= not(layer4_outputs(7213));
    layer5_outputs(4776) <= not(layer4_outputs(540)) or (layer4_outputs(4109));
    layer5_outputs(4777) <= (layer4_outputs(2505)) and not (layer4_outputs(5711));
    layer5_outputs(4778) <= not(layer4_outputs(237)) or (layer4_outputs(5560));
    layer5_outputs(4779) <= not((layer4_outputs(3507)) xor (layer4_outputs(2564)));
    layer5_outputs(4780) <= not(layer4_outputs(3593));
    layer5_outputs(4781) <= layer4_outputs(2984);
    layer5_outputs(4782) <= layer4_outputs(690);
    layer5_outputs(4783) <= not(layer4_outputs(4479)) or (layer4_outputs(6566));
    layer5_outputs(4784) <= (layer4_outputs(2819)) and (layer4_outputs(1109));
    layer5_outputs(4785) <= not(layer4_outputs(5259)) or (layer4_outputs(3512));
    layer5_outputs(4786) <= (layer4_outputs(2581)) and (layer4_outputs(3434));
    layer5_outputs(4787) <= '1';
    layer5_outputs(4788) <= layer4_outputs(5021);
    layer5_outputs(4789) <= '0';
    layer5_outputs(4790) <= not(layer4_outputs(6334));
    layer5_outputs(4791) <= not(layer4_outputs(6682));
    layer5_outputs(4792) <= not((layer4_outputs(5352)) or (layer4_outputs(230)));
    layer5_outputs(4793) <= not(layer4_outputs(976));
    layer5_outputs(4794) <= layer4_outputs(1102);
    layer5_outputs(4795) <= not(layer4_outputs(5678));
    layer5_outputs(4796) <= '1';
    layer5_outputs(4797) <= layer4_outputs(4596);
    layer5_outputs(4798) <= not(layer4_outputs(4115));
    layer5_outputs(4799) <= (layer4_outputs(321)) and not (layer4_outputs(2066));
    layer5_outputs(4800) <= not((layer4_outputs(3254)) xor (layer4_outputs(6341)));
    layer5_outputs(4801) <= not(layer4_outputs(3615));
    layer5_outputs(4802) <= layer4_outputs(7388);
    layer5_outputs(4803) <= layer4_outputs(5932);
    layer5_outputs(4804) <= (layer4_outputs(5978)) and not (layer4_outputs(883));
    layer5_outputs(4805) <= not(layer4_outputs(6610));
    layer5_outputs(4806) <= (layer4_outputs(7060)) or (layer4_outputs(3949));
    layer5_outputs(4807) <= '0';
    layer5_outputs(4808) <= not(layer4_outputs(3908));
    layer5_outputs(4809) <= (layer4_outputs(1509)) and not (layer4_outputs(7150));
    layer5_outputs(4810) <= '1';
    layer5_outputs(4811) <= layer4_outputs(5065);
    layer5_outputs(4812) <= layer4_outputs(1610);
    layer5_outputs(4813) <= not(layer4_outputs(2687)) or (layer4_outputs(222));
    layer5_outputs(4814) <= layer4_outputs(3683);
    layer5_outputs(4815) <= not(layer4_outputs(3072));
    layer5_outputs(4816) <= not(layer4_outputs(3729));
    layer5_outputs(4817) <= not(layer4_outputs(4322));
    layer5_outputs(4818) <= layer4_outputs(4624);
    layer5_outputs(4819) <= (layer4_outputs(2824)) or (layer4_outputs(793));
    layer5_outputs(4820) <= (layer4_outputs(5843)) or (layer4_outputs(652));
    layer5_outputs(4821) <= (layer4_outputs(5517)) and (layer4_outputs(2587));
    layer5_outputs(4822) <= not(layer4_outputs(2731));
    layer5_outputs(4823) <= not((layer4_outputs(2629)) and (layer4_outputs(4550)));
    layer5_outputs(4824) <= not(layer4_outputs(3416));
    layer5_outputs(4825) <= layer4_outputs(4558);
    layer5_outputs(4826) <= (layer4_outputs(7635)) xor (layer4_outputs(7348));
    layer5_outputs(4827) <= not(layer4_outputs(3063));
    layer5_outputs(4828) <= (layer4_outputs(2445)) xor (layer4_outputs(3695));
    layer5_outputs(4829) <= not(layer4_outputs(567));
    layer5_outputs(4830) <= layer4_outputs(1301);
    layer5_outputs(4831) <= layer4_outputs(5221);
    layer5_outputs(4832) <= (layer4_outputs(2121)) and not (layer4_outputs(7376));
    layer5_outputs(4833) <= not(layer4_outputs(4654));
    layer5_outputs(4834) <= not(layer4_outputs(740));
    layer5_outputs(4835) <= layer4_outputs(2730);
    layer5_outputs(4836) <= not(layer4_outputs(2188));
    layer5_outputs(4837) <= not(layer4_outputs(2029));
    layer5_outputs(4838) <= layer4_outputs(1684);
    layer5_outputs(4839) <= not(layer4_outputs(4920));
    layer5_outputs(4840) <= not(layer4_outputs(4263)) or (layer4_outputs(4720));
    layer5_outputs(4841) <= not((layer4_outputs(6003)) xor (layer4_outputs(1315)));
    layer5_outputs(4842) <= '0';
    layer5_outputs(4843) <= (layer4_outputs(4508)) or (layer4_outputs(7446));
    layer5_outputs(4844) <= layer4_outputs(1725);
    layer5_outputs(4845) <= layer4_outputs(6760);
    layer5_outputs(4846) <= layer4_outputs(2736);
    layer5_outputs(4847) <= layer4_outputs(6137);
    layer5_outputs(4848) <= not(layer4_outputs(1586)) or (layer4_outputs(5766));
    layer5_outputs(4849) <= '1';
    layer5_outputs(4850) <= not((layer4_outputs(7081)) or (layer4_outputs(1411)));
    layer5_outputs(4851) <= not((layer4_outputs(3952)) or (layer4_outputs(6182)));
    layer5_outputs(4852) <= not((layer4_outputs(2359)) xor (layer4_outputs(5205)));
    layer5_outputs(4853) <= not((layer4_outputs(6843)) or (layer4_outputs(3044)));
    layer5_outputs(4854) <= not((layer4_outputs(3186)) xor (layer4_outputs(2612)));
    layer5_outputs(4855) <= not(layer4_outputs(5715));
    layer5_outputs(4856) <= layer4_outputs(5444);
    layer5_outputs(4857) <= '0';
    layer5_outputs(4858) <= layer4_outputs(5068);
    layer5_outputs(4859) <= not(layer4_outputs(4522)) or (layer4_outputs(4514));
    layer5_outputs(4860) <= not(layer4_outputs(4795));
    layer5_outputs(4861) <= not(layer4_outputs(6823));
    layer5_outputs(4862) <= layer4_outputs(6973);
    layer5_outputs(4863) <= layer4_outputs(5718);
    layer5_outputs(4864) <= layer4_outputs(1963);
    layer5_outputs(4865) <= (layer4_outputs(3199)) and not (layer4_outputs(2787));
    layer5_outputs(4866) <= (layer4_outputs(2852)) and not (layer4_outputs(3575));
    layer5_outputs(4867) <= not(layer4_outputs(7410)) or (layer4_outputs(129));
    layer5_outputs(4868) <= not(layer4_outputs(425));
    layer5_outputs(4869) <= not(layer4_outputs(2544));
    layer5_outputs(4870) <= '1';
    layer5_outputs(4871) <= not(layer4_outputs(2781));
    layer5_outputs(4872) <= (layer4_outputs(4691)) xor (layer4_outputs(7603));
    layer5_outputs(4873) <= not(layer4_outputs(99));
    layer5_outputs(4874) <= not((layer4_outputs(7054)) or (layer4_outputs(7235)));
    layer5_outputs(4875) <= '0';
    layer5_outputs(4876) <= layer4_outputs(2207);
    layer5_outputs(4877) <= not(layer4_outputs(2334));
    layer5_outputs(4878) <= layer4_outputs(2658);
    layer5_outputs(4879) <= layer4_outputs(1895);
    layer5_outputs(4880) <= not(layer4_outputs(1254));
    layer5_outputs(4881) <= not(layer4_outputs(4387));
    layer5_outputs(4882) <= layer4_outputs(2899);
    layer5_outputs(4883) <= '0';
    layer5_outputs(4884) <= (layer4_outputs(2823)) and not (layer4_outputs(3498));
    layer5_outputs(4885) <= not(layer4_outputs(7070));
    layer5_outputs(4886) <= not(layer4_outputs(1825));
    layer5_outputs(4887) <= not((layer4_outputs(6277)) and (layer4_outputs(4281)));
    layer5_outputs(4888) <= not((layer4_outputs(5285)) or (layer4_outputs(5290)));
    layer5_outputs(4889) <= layer4_outputs(4785);
    layer5_outputs(4890) <= not(layer4_outputs(1211));
    layer5_outputs(4891) <= not((layer4_outputs(4568)) xor (layer4_outputs(4893)));
    layer5_outputs(4892) <= layer4_outputs(1243);
    layer5_outputs(4893) <= layer4_outputs(2783);
    layer5_outputs(4894) <= layer4_outputs(5125);
    layer5_outputs(4895) <= not(layer4_outputs(4721));
    layer5_outputs(4896) <= not(layer4_outputs(1849));
    layer5_outputs(4897) <= layer4_outputs(7007);
    layer5_outputs(4898) <= layer4_outputs(2354);
    layer5_outputs(4899) <= not(layer4_outputs(4005));
    layer5_outputs(4900) <= not((layer4_outputs(162)) and (layer4_outputs(3040)));
    layer5_outputs(4901) <= layer4_outputs(896);
    layer5_outputs(4902) <= (layer4_outputs(4249)) or (layer4_outputs(5438));
    layer5_outputs(4903) <= (layer4_outputs(7114)) and not (layer4_outputs(2986));
    layer5_outputs(4904) <= layer4_outputs(2423);
    layer5_outputs(4905) <= layer4_outputs(3334);
    layer5_outputs(4906) <= not((layer4_outputs(2865)) xor (layer4_outputs(6020)));
    layer5_outputs(4907) <= layer4_outputs(7065);
    layer5_outputs(4908) <= layer4_outputs(7665);
    layer5_outputs(4909) <= not(layer4_outputs(1983)) or (layer4_outputs(668));
    layer5_outputs(4910) <= (layer4_outputs(2028)) or (layer4_outputs(1836));
    layer5_outputs(4911) <= not(layer4_outputs(7486)) or (layer4_outputs(2609));
    layer5_outputs(4912) <= layer4_outputs(591);
    layer5_outputs(4913) <= not((layer4_outputs(4577)) or (layer4_outputs(957)));
    layer5_outputs(4914) <= not(layer4_outputs(4621));
    layer5_outputs(4915) <= layer4_outputs(2539);
    layer5_outputs(4916) <= not(layer4_outputs(283));
    layer5_outputs(4917) <= not((layer4_outputs(2446)) xor (layer4_outputs(7533)));
    layer5_outputs(4918) <= layer4_outputs(1545);
    layer5_outputs(4919) <= not((layer4_outputs(4701)) xor (layer4_outputs(3323)));
    layer5_outputs(4920) <= (layer4_outputs(4717)) or (layer4_outputs(98));
    layer5_outputs(4921) <= not(layer4_outputs(5573));
    layer5_outputs(4922) <= not((layer4_outputs(2204)) xor (layer4_outputs(5657)));
    layer5_outputs(4923) <= (layer4_outputs(7337)) xor (layer4_outputs(5163));
    layer5_outputs(4924) <= not(layer4_outputs(5430));
    layer5_outputs(4925) <= not(layer4_outputs(6567));
    layer5_outputs(4926) <= layer4_outputs(5587);
    layer5_outputs(4927) <= not((layer4_outputs(3126)) and (layer4_outputs(6289)));
    layer5_outputs(4928) <= not(layer4_outputs(3313)) or (layer4_outputs(1587));
    layer5_outputs(4929) <= (layer4_outputs(2239)) and not (layer4_outputs(578));
    layer5_outputs(4930) <= not(layer4_outputs(3399));
    layer5_outputs(4931) <= layer4_outputs(7599);
    layer5_outputs(4932) <= not((layer4_outputs(1036)) xor (layer4_outputs(1756)));
    layer5_outputs(4933) <= not(layer4_outputs(6699));
    layer5_outputs(4934) <= not(layer4_outputs(6792));
    layer5_outputs(4935) <= not(layer4_outputs(6546)) or (layer4_outputs(3491));
    layer5_outputs(4936) <= layer4_outputs(3979);
    layer5_outputs(4937) <= not(layer4_outputs(1408));
    layer5_outputs(4938) <= (layer4_outputs(1686)) or (layer4_outputs(5696));
    layer5_outputs(4939) <= (layer4_outputs(4055)) or (layer4_outputs(5788));
    layer5_outputs(4940) <= layer4_outputs(6078);
    layer5_outputs(4941) <= layer4_outputs(297);
    layer5_outputs(4942) <= '1';
    layer5_outputs(4943) <= (layer4_outputs(4383)) and (layer4_outputs(5169));
    layer5_outputs(4944) <= layer4_outputs(879);
    layer5_outputs(4945) <= layer4_outputs(3763);
    layer5_outputs(4946) <= layer4_outputs(6796);
    layer5_outputs(4947) <= not(layer4_outputs(4668));
    layer5_outputs(4948) <= layer4_outputs(5413);
    layer5_outputs(4949) <= not(layer4_outputs(5538));
    layer5_outputs(4950) <= not((layer4_outputs(3050)) xor (layer4_outputs(2416)));
    layer5_outputs(4951) <= layer4_outputs(4912);
    layer5_outputs(4952) <= layer4_outputs(5334);
    layer5_outputs(4953) <= layer4_outputs(2131);
    layer5_outputs(4954) <= (layer4_outputs(3749)) or (layer4_outputs(6333));
    layer5_outputs(4955) <= layer4_outputs(6416);
    layer5_outputs(4956) <= (layer4_outputs(5282)) or (layer4_outputs(722));
    layer5_outputs(4957) <= layer4_outputs(6281);
    layer5_outputs(4958) <= layer4_outputs(190);
    layer5_outputs(4959) <= not(layer4_outputs(3730));
    layer5_outputs(4960) <= not(layer4_outputs(3132));
    layer5_outputs(4961) <= not((layer4_outputs(2471)) or (layer4_outputs(7449)));
    layer5_outputs(4962) <= (layer4_outputs(6166)) and not (layer4_outputs(1428));
    layer5_outputs(4963) <= not((layer4_outputs(7441)) or (layer4_outputs(3429)));
    layer5_outputs(4964) <= not(layer4_outputs(3710)) or (layer4_outputs(5367));
    layer5_outputs(4965) <= not(layer4_outputs(5016));
    layer5_outputs(4966) <= not(layer4_outputs(2484));
    layer5_outputs(4967) <= (layer4_outputs(7102)) and not (layer4_outputs(663));
    layer5_outputs(4968) <= (layer4_outputs(1510)) xor (layer4_outputs(1315));
    layer5_outputs(4969) <= (layer4_outputs(4783)) or (layer4_outputs(2944));
    layer5_outputs(4970) <= (layer4_outputs(3133)) xor (layer4_outputs(3630));
    layer5_outputs(4971) <= not((layer4_outputs(3595)) or (layer4_outputs(3460)));
    layer5_outputs(4972) <= not(layer4_outputs(1262)) or (layer4_outputs(7458));
    layer5_outputs(4973) <= not(layer4_outputs(7442));
    layer5_outputs(4974) <= not(layer4_outputs(3210)) or (layer4_outputs(257));
    layer5_outputs(4975) <= not(layer4_outputs(7030));
    layer5_outputs(4976) <= not(layer4_outputs(2249));
    layer5_outputs(4977) <= (layer4_outputs(2094)) and (layer4_outputs(5059));
    layer5_outputs(4978) <= not(layer4_outputs(6343));
    layer5_outputs(4979) <= not((layer4_outputs(2979)) and (layer4_outputs(2582)));
    layer5_outputs(4980) <= (layer4_outputs(3796)) and (layer4_outputs(5842));
    layer5_outputs(4981) <= (layer4_outputs(573)) or (layer4_outputs(3904));
    layer5_outputs(4982) <= not(layer4_outputs(5478));
    layer5_outputs(4983) <= not((layer4_outputs(555)) and (layer4_outputs(6677)));
    layer5_outputs(4984) <= not(layer4_outputs(5828));
    layer5_outputs(4985) <= (layer4_outputs(5384)) or (layer4_outputs(6873));
    layer5_outputs(4986) <= (layer4_outputs(4062)) xor (layer4_outputs(3289));
    layer5_outputs(4987) <= not(layer4_outputs(2674));
    layer5_outputs(4988) <= (layer4_outputs(5488)) and not (layer4_outputs(2608));
    layer5_outputs(4989) <= not(layer4_outputs(1506));
    layer5_outputs(4990) <= layer4_outputs(7467);
    layer5_outputs(4991) <= layer4_outputs(5713);
    layer5_outputs(4992) <= (layer4_outputs(852)) and not (layer4_outputs(6260));
    layer5_outputs(4993) <= layer4_outputs(1379);
    layer5_outputs(4994) <= not(layer4_outputs(3921));
    layer5_outputs(4995) <= not(layer4_outputs(5570));
    layer5_outputs(4996) <= not(layer4_outputs(4019)) or (layer4_outputs(1578));
    layer5_outputs(4997) <= not(layer4_outputs(6417));
    layer5_outputs(4998) <= layer4_outputs(352);
    layer5_outputs(4999) <= not((layer4_outputs(5416)) and (layer4_outputs(4838)));
    layer5_outputs(5000) <= not(layer4_outputs(1223));
    layer5_outputs(5001) <= not(layer4_outputs(5701));
    layer5_outputs(5002) <= not(layer4_outputs(5364));
    layer5_outputs(5003) <= not((layer4_outputs(2408)) xor (layer4_outputs(700)));
    layer5_outputs(5004) <= (layer4_outputs(244)) and (layer4_outputs(2169));
    layer5_outputs(5005) <= layer4_outputs(1110);
    layer5_outputs(5006) <= layer4_outputs(2561);
    layer5_outputs(5007) <= not(layer4_outputs(3034)) or (layer4_outputs(801));
    layer5_outputs(5008) <= not(layer4_outputs(268));
    layer5_outputs(5009) <= not(layer4_outputs(3038));
    layer5_outputs(5010) <= not((layer4_outputs(2721)) and (layer4_outputs(6666)));
    layer5_outputs(5011) <= (layer4_outputs(2729)) or (layer4_outputs(2934));
    layer5_outputs(5012) <= not(layer4_outputs(629)) or (layer4_outputs(4915));
    layer5_outputs(5013) <= (layer4_outputs(2399)) or (layer4_outputs(6722));
    layer5_outputs(5014) <= (layer4_outputs(549)) or (layer4_outputs(2626));
    layer5_outputs(5015) <= not((layer4_outputs(5101)) xor (layer4_outputs(7591)));
    layer5_outputs(5016) <= not((layer4_outputs(2263)) or (layer4_outputs(1005)));
    layer5_outputs(5017) <= (layer4_outputs(6819)) and (layer4_outputs(3871));
    layer5_outputs(5018) <= (layer4_outputs(5580)) and (layer4_outputs(321));
    layer5_outputs(5019) <= not(layer4_outputs(5827));
    layer5_outputs(5020) <= layer4_outputs(887);
    layer5_outputs(5021) <= layer4_outputs(118);
    layer5_outputs(5022) <= not(layer4_outputs(2103));
    layer5_outputs(5023) <= not(layer4_outputs(1134));
    layer5_outputs(5024) <= layer4_outputs(4931);
    layer5_outputs(5025) <= layer4_outputs(1376);
    layer5_outputs(5026) <= not((layer4_outputs(3088)) or (layer4_outputs(6132)));
    layer5_outputs(5027) <= layer4_outputs(2232);
    layer5_outputs(5028) <= not(layer4_outputs(3776));
    layer5_outputs(5029) <= not(layer4_outputs(5579));
    layer5_outputs(5030) <= not((layer4_outputs(3953)) and (layer4_outputs(3402)));
    layer5_outputs(5031) <= not(layer4_outputs(1548));
    layer5_outputs(5032) <= (layer4_outputs(6083)) xor (layer4_outputs(1535));
    layer5_outputs(5033) <= (layer4_outputs(3209)) and (layer4_outputs(4519));
    layer5_outputs(5034) <= (layer4_outputs(3678)) and (layer4_outputs(6284));
    layer5_outputs(5035) <= layer4_outputs(6421);
    layer5_outputs(5036) <= not((layer4_outputs(4456)) or (layer4_outputs(1459)));
    layer5_outputs(5037) <= not((layer4_outputs(5030)) xor (layer4_outputs(7026)));
    layer5_outputs(5038) <= '0';
    layer5_outputs(5039) <= layer4_outputs(4841);
    layer5_outputs(5040) <= layer4_outputs(5005);
    layer5_outputs(5041) <= not(layer4_outputs(4003));
    layer5_outputs(5042) <= not(layer4_outputs(59)) or (layer4_outputs(2083));
    layer5_outputs(5043) <= not(layer4_outputs(2922));
    layer5_outputs(5044) <= (layer4_outputs(4182)) xor (layer4_outputs(1616));
    layer5_outputs(5045) <= (layer4_outputs(2364)) xor (layer4_outputs(288));
    layer5_outputs(5046) <= not(layer4_outputs(5771));
    layer5_outputs(5047) <= (layer4_outputs(7045)) xor (layer4_outputs(646));
    layer5_outputs(5048) <= not((layer4_outputs(5741)) and (layer4_outputs(5084)));
    layer5_outputs(5049) <= layer4_outputs(5262);
    layer5_outputs(5050) <= not(layer4_outputs(539));
    layer5_outputs(5051) <= (layer4_outputs(1790)) xor (layer4_outputs(7501));
    layer5_outputs(5052) <= not(layer4_outputs(119));
    layer5_outputs(5053) <= not(layer4_outputs(6820)) or (layer4_outputs(1993));
    layer5_outputs(5054) <= (layer4_outputs(2043)) or (layer4_outputs(4887));
    layer5_outputs(5055) <= not(layer4_outputs(3190)) or (layer4_outputs(3378));
    layer5_outputs(5056) <= not(layer4_outputs(3743));
    layer5_outputs(5057) <= not((layer4_outputs(1239)) xor (layer4_outputs(5298)));
    layer5_outputs(5058) <= (layer4_outputs(880)) or (layer4_outputs(3736));
    layer5_outputs(5059) <= not(layer4_outputs(1286));
    layer5_outputs(5060) <= layer4_outputs(4257);
    layer5_outputs(5061) <= not((layer4_outputs(5137)) xor (layer4_outputs(3779)));
    layer5_outputs(5062) <= not(layer4_outputs(5744));
    layer5_outputs(5063) <= not((layer4_outputs(5799)) or (layer4_outputs(5255)));
    layer5_outputs(5064) <= not((layer4_outputs(3279)) xor (layer4_outputs(3003)));
    layer5_outputs(5065) <= (layer4_outputs(7550)) or (layer4_outputs(1093));
    layer5_outputs(5066) <= not((layer4_outputs(1527)) or (layer4_outputs(3721)));
    layer5_outputs(5067) <= not(layer4_outputs(4002)) or (layer4_outputs(1067));
    layer5_outputs(5068) <= not(layer4_outputs(6945)) or (layer4_outputs(4688));
    layer5_outputs(5069) <= not((layer4_outputs(6467)) and (layer4_outputs(2684)));
    layer5_outputs(5070) <= not(layer4_outputs(2119));
    layer5_outputs(5071) <= layer4_outputs(6277);
    layer5_outputs(5072) <= not(layer4_outputs(6043));
    layer5_outputs(5073) <= not(layer4_outputs(4826));
    layer5_outputs(5074) <= not((layer4_outputs(3762)) and (layer4_outputs(550)));
    layer5_outputs(5075) <= (layer4_outputs(4567)) xor (layer4_outputs(4611));
    layer5_outputs(5076) <= not(layer4_outputs(1545));
    layer5_outputs(5077) <= (layer4_outputs(7572)) and not (layer4_outputs(4874));
    layer5_outputs(5078) <= not(layer4_outputs(1518)) or (layer4_outputs(4105));
    layer5_outputs(5079) <= not(layer4_outputs(2602));
    layer5_outputs(5080) <= not(layer4_outputs(3745));
    layer5_outputs(5081) <= not(layer4_outputs(6472));
    layer5_outputs(5082) <= not(layer4_outputs(1700)) or (layer4_outputs(2435));
    layer5_outputs(5083) <= not((layer4_outputs(3887)) or (layer4_outputs(7128)));
    layer5_outputs(5084) <= (layer4_outputs(3844)) and (layer4_outputs(5075));
    layer5_outputs(5085) <= not((layer4_outputs(5314)) or (layer4_outputs(2346)));
    layer5_outputs(5086) <= layer4_outputs(6143);
    layer5_outputs(5087) <= not(layer4_outputs(2634));
    layer5_outputs(5088) <= layer4_outputs(1698);
    layer5_outputs(5089) <= layer4_outputs(1941);
    layer5_outputs(5090) <= not(layer4_outputs(475));
    layer5_outputs(5091) <= (layer4_outputs(3880)) and not (layer4_outputs(6689));
    layer5_outputs(5092) <= (layer4_outputs(4932)) and not (layer4_outputs(3085));
    layer5_outputs(5093) <= (layer4_outputs(4017)) and (layer4_outputs(6897));
    layer5_outputs(5094) <= (layer4_outputs(4532)) and not (layer4_outputs(4605));
    layer5_outputs(5095) <= (layer4_outputs(664)) xor (layer4_outputs(627));
    layer5_outputs(5096) <= not(layer4_outputs(6865)) or (layer4_outputs(2853));
    layer5_outputs(5097) <= layer4_outputs(1404);
    layer5_outputs(5098) <= (layer4_outputs(6224)) xor (layer4_outputs(2352));
    layer5_outputs(5099) <= layer4_outputs(1327);
    layer5_outputs(5100) <= layer4_outputs(4673);
    layer5_outputs(5101) <= layer4_outputs(6626);
    layer5_outputs(5102) <= not((layer4_outputs(2297)) xor (layer4_outputs(6510)));
    layer5_outputs(5103) <= (layer4_outputs(2856)) xor (layer4_outputs(1014));
    layer5_outputs(5104) <= '1';
    layer5_outputs(5105) <= layer4_outputs(2141);
    layer5_outputs(5106) <= not(layer4_outputs(3247));
    layer5_outputs(5107) <= not((layer4_outputs(4769)) and (layer4_outputs(7050)));
    layer5_outputs(5108) <= not((layer4_outputs(7238)) xor (layer4_outputs(439)));
    layer5_outputs(5109) <= (layer4_outputs(7130)) xor (layer4_outputs(4863));
    layer5_outputs(5110) <= not((layer4_outputs(1870)) or (layer4_outputs(815)));
    layer5_outputs(5111) <= not(layer4_outputs(3080)) or (layer4_outputs(5673));
    layer5_outputs(5112) <= not(layer4_outputs(6008));
    layer5_outputs(5113) <= not(layer4_outputs(5143)) or (layer4_outputs(6327));
    layer5_outputs(5114) <= not((layer4_outputs(4762)) and (layer4_outputs(6668)));
    layer5_outputs(5115) <= not((layer4_outputs(4224)) and (layer4_outputs(4725)));
    layer5_outputs(5116) <= not((layer4_outputs(6664)) and (layer4_outputs(2734)));
    layer5_outputs(5117) <= not(layer4_outputs(4446));
    layer5_outputs(5118) <= layer4_outputs(2741);
    layer5_outputs(5119) <= not(layer4_outputs(6344)) or (layer4_outputs(95));
    layer5_outputs(5120) <= (layer4_outputs(1651)) and (layer4_outputs(3301));
    layer5_outputs(5121) <= (layer4_outputs(7223)) and not (layer4_outputs(4463));
    layer5_outputs(5122) <= '0';
    layer5_outputs(5123) <= (layer4_outputs(3391)) and (layer4_outputs(816));
    layer5_outputs(5124) <= not(layer4_outputs(7274));
    layer5_outputs(5125) <= layer4_outputs(5356);
    layer5_outputs(5126) <= '1';
    layer5_outputs(5127) <= not(layer4_outputs(3028));
    layer5_outputs(5128) <= (layer4_outputs(6910)) xor (layer4_outputs(89));
    layer5_outputs(5129) <= layer4_outputs(7364);
    layer5_outputs(5130) <= layer4_outputs(4971);
    layer5_outputs(5131) <= not((layer4_outputs(5283)) and (layer4_outputs(4727)));
    layer5_outputs(5132) <= (layer4_outputs(2915)) xor (layer4_outputs(3573));
    layer5_outputs(5133) <= (layer4_outputs(2299)) or (layer4_outputs(117));
    layer5_outputs(5134) <= not(layer4_outputs(1105));
    layer5_outputs(5135) <= not(layer4_outputs(3570));
    layer5_outputs(5136) <= not(layer4_outputs(1729));
    layer5_outputs(5137) <= layer4_outputs(7362);
    layer5_outputs(5138) <= not(layer4_outputs(280));
    layer5_outputs(5139) <= layer4_outputs(2688);
    layer5_outputs(5140) <= not(layer4_outputs(6388));
    layer5_outputs(5141) <= not(layer4_outputs(463)) or (layer4_outputs(992));
    layer5_outputs(5142) <= (layer4_outputs(2469)) and not (layer4_outputs(1755));
    layer5_outputs(5143) <= (layer4_outputs(4030)) xor (layer4_outputs(5607));
    layer5_outputs(5144) <= (layer4_outputs(1777)) and not (layer4_outputs(5874));
    layer5_outputs(5145) <= not(layer4_outputs(7024));
    layer5_outputs(5146) <= (layer4_outputs(651)) and (layer4_outputs(3840));
    layer5_outputs(5147) <= not(layer4_outputs(1189));
    layer5_outputs(5148) <= not(layer4_outputs(5067));
    layer5_outputs(5149) <= '1';
    layer5_outputs(5150) <= layer4_outputs(4648);
    layer5_outputs(5151) <= not((layer4_outputs(4614)) xor (layer4_outputs(3452)));
    layer5_outputs(5152) <= not((layer4_outputs(7034)) xor (layer4_outputs(3043)));
    layer5_outputs(5153) <= not((layer4_outputs(3753)) or (layer4_outputs(1196)));
    layer5_outputs(5154) <= (layer4_outputs(3702)) and not (layer4_outputs(2366));
    layer5_outputs(5155) <= not((layer4_outputs(1153)) xor (layer4_outputs(3829)));
    layer5_outputs(5156) <= layer4_outputs(3940);
    layer5_outputs(5157) <= layer4_outputs(6665);
    layer5_outputs(5158) <= (layer4_outputs(1289)) xor (layer4_outputs(806));
    layer5_outputs(5159) <= layer4_outputs(7540);
    layer5_outputs(5160) <= not(layer4_outputs(624));
    layer5_outputs(5161) <= not(layer4_outputs(2098));
    layer5_outputs(5162) <= not((layer4_outputs(5773)) or (layer4_outputs(5389)));
    layer5_outputs(5163) <= not(layer4_outputs(2170));
    layer5_outputs(5164) <= not(layer4_outputs(2811));
    layer5_outputs(5165) <= layer4_outputs(5722);
    layer5_outputs(5166) <= not(layer4_outputs(4830));
    layer5_outputs(5167) <= not(layer4_outputs(2925));
    layer5_outputs(5168) <= not(layer4_outputs(997));
    layer5_outputs(5169) <= (layer4_outputs(1185)) xor (layer4_outputs(2200));
    layer5_outputs(5170) <= not(layer4_outputs(2280));
    layer5_outputs(5171) <= layer4_outputs(1281);
    layer5_outputs(5172) <= layer4_outputs(5406);
    layer5_outputs(5173) <= not(layer4_outputs(2664));
    layer5_outputs(5174) <= not(layer4_outputs(5618));
    layer5_outputs(5175) <= (layer4_outputs(2705)) and not (layer4_outputs(2756));
    layer5_outputs(5176) <= not(layer4_outputs(1737)) or (layer4_outputs(2427));
    layer5_outputs(5177) <= (layer4_outputs(1118)) and not (layer4_outputs(6182));
    layer5_outputs(5178) <= (layer4_outputs(1747)) and not (layer4_outputs(2130));
    layer5_outputs(5179) <= (layer4_outputs(967)) xor (layer4_outputs(7475));
    layer5_outputs(5180) <= not(layer4_outputs(2374));
    layer5_outputs(5181) <= not(layer4_outputs(3641)) or (layer4_outputs(2574));
    layer5_outputs(5182) <= layer4_outputs(1669);
    layer5_outputs(5183) <= not(layer4_outputs(536));
    layer5_outputs(5184) <= not((layer4_outputs(4451)) xor (layer4_outputs(6975)));
    layer5_outputs(5185) <= not(layer4_outputs(6702));
    layer5_outputs(5186) <= (layer4_outputs(3752)) and not (layer4_outputs(6295));
    layer5_outputs(5187) <= not(layer4_outputs(4596));
    layer5_outputs(5188) <= '0';
    layer5_outputs(5189) <= (layer4_outputs(3030)) and not (layer4_outputs(1042));
    layer5_outputs(5190) <= layer4_outputs(5428);
    layer5_outputs(5191) <= not(layer4_outputs(5991));
    layer5_outputs(5192) <= not(layer4_outputs(886));
    layer5_outputs(5193) <= layer4_outputs(7678);
    layer5_outputs(5194) <= not((layer4_outputs(3758)) or (layer4_outputs(4364)));
    layer5_outputs(5195) <= not(layer4_outputs(3854)) or (layer4_outputs(4500));
    layer5_outputs(5196) <= (layer4_outputs(3915)) or (layer4_outputs(4913));
    layer5_outputs(5197) <= not((layer4_outputs(5946)) xor (layer4_outputs(3339)));
    layer5_outputs(5198) <= not(layer4_outputs(5413)) or (layer4_outputs(593));
    layer5_outputs(5199) <= layer4_outputs(4209);
    layer5_outputs(5200) <= (layer4_outputs(2126)) or (layer4_outputs(3369));
    layer5_outputs(5201) <= not(layer4_outputs(5808));
    layer5_outputs(5202) <= not((layer4_outputs(4474)) xor (layer4_outputs(3135)));
    layer5_outputs(5203) <= layer4_outputs(1372);
    layer5_outputs(5204) <= (layer4_outputs(6555)) xor (layer4_outputs(392));
    layer5_outputs(5205) <= layer4_outputs(7164);
    layer5_outputs(5206) <= (layer4_outputs(4004)) and not (layer4_outputs(1160));
    layer5_outputs(5207) <= layer4_outputs(7050);
    layer5_outputs(5208) <= layer4_outputs(153);
    layer5_outputs(5209) <= (layer4_outputs(6633)) and not (layer4_outputs(6861));
    layer5_outputs(5210) <= not(layer4_outputs(4193));
    layer5_outputs(5211) <= '0';
    layer5_outputs(5212) <= not(layer4_outputs(3939));
    layer5_outputs(5213) <= (layer4_outputs(4313)) or (layer4_outputs(3680));
    layer5_outputs(5214) <= not((layer4_outputs(4622)) and (layer4_outputs(4241)));
    layer5_outputs(5215) <= not(layer4_outputs(6588)) or (layer4_outputs(7017));
    layer5_outputs(5216) <= (layer4_outputs(7038)) or (layer4_outputs(6047));
    layer5_outputs(5217) <= layer4_outputs(703);
    layer5_outputs(5218) <= not(layer4_outputs(689)) or (layer4_outputs(1289));
    layer5_outputs(5219) <= not(layer4_outputs(3014));
    layer5_outputs(5220) <= layer4_outputs(720);
    layer5_outputs(5221) <= not(layer4_outputs(2631));
    layer5_outputs(5222) <= not(layer4_outputs(7582));
    layer5_outputs(5223) <= (layer4_outputs(7091)) and not (layer4_outputs(2542));
    layer5_outputs(5224) <= layer4_outputs(7412);
    layer5_outputs(5225) <= layer4_outputs(4652);
    layer5_outputs(5226) <= (layer4_outputs(5600)) xor (layer4_outputs(7177));
    layer5_outputs(5227) <= not((layer4_outputs(1772)) and (layer4_outputs(4627)));
    layer5_outputs(5228) <= not((layer4_outputs(1423)) xor (layer4_outputs(144)));
    layer5_outputs(5229) <= not(layer4_outputs(1439));
    layer5_outputs(5230) <= (layer4_outputs(5140)) and not (layer4_outputs(5953));
    layer5_outputs(5231) <= not(layer4_outputs(775));
    layer5_outputs(5232) <= not((layer4_outputs(4276)) xor (layer4_outputs(1764)));
    layer5_outputs(5233) <= (layer4_outputs(4764)) xor (layer4_outputs(5808));
    layer5_outputs(5234) <= not(layer4_outputs(1756)) or (layer4_outputs(728));
    layer5_outputs(5235) <= not(layer4_outputs(564));
    layer5_outputs(5236) <= not((layer4_outputs(4234)) xor (layer4_outputs(4365)));
    layer5_outputs(5237) <= '1';
    layer5_outputs(5238) <= not(layer4_outputs(1492));
    layer5_outputs(5239) <= (layer4_outputs(4541)) and not (layer4_outputs(16));
    layer5_outputs(5240) <= (layer4_outputs(3771)) and not (layer4_outputs(7575));
    layer5_outputs(5241) <= layer4_outputs(6566);
    layer5_outputs(5242) <= (layer4_outputs(5683)) and not (layer4_outputs(7399));
    layer5_outputs(5243) <= (layer4_outputs(1706)) and not (layer4_outputs(2934));
    layer5_outputs(5244) <= (layer4_outputs(6028)) xor (layer4_outputs(6609));
    layer5_outputs(5245) <= (layer4_outputs(3281)) and not (layer4_outputs(1114));
    layer5_outputs(5246) <= (layer4_outputs(2643)) xor (layer4_outputs(4664));
    layer5_outputs(5247) <= (layer4_outputs(3048)) and not (layer4_outputs(1782));
    layer5_outputs(5248) <= layer4_outputs(5674);
    layer5_outputs(5249) <= layer4_outputs(4981);
    layer5_outputs(5250) <= not((layer4_outputs(2178)) and (layer4_outputs(1741)));
    layer5_outputs(5251) <= layer4_outputs(6950);
    layer5_outputs(5252) <= not(layer4_outputs(2157));
    layer5_outputs(5253) <= (layer4_outputs(3591)) or (layer4_outputs(527));
    layer5_outputs(5254) <= layer4_outputs(7631);
    layer5_outputs(5255) <= not((layer4_outputs(4885)) or (layer4_outputs(1834)));
    layer5_outputs(5256) <= layer4_outputs(4130);
    layer5_outputs(5257) <= layer4_outputs(2596);
    layer5_outputs(5258) <= not(layer4_outputs(2373)) or (layer4_outputs(193));
    layer5_outputs(5259) <= not(layer4_outputs(7476)) or (layer4_outputs(5844));
    layer5_outputs(5260) <= layer4_outputs(1593);
    layer5_outputs(5261) <= not(layer4_outputs(3028));
    layer5_outputs(5262) <= (layer4_outputs(1058)) and (layer4_outputs(5479));
    layer5_outputs(5263) <= layer4_outputs(6162);
    layer5_outputs(5264) <= not(layer4_outputs(6180));
    layer5_outputs(5265) <= not(layer4_outputs(5755));
    layer5_outputs(5266) <= layer4_outputs(6457);
    layer5_outputs(5267) <= layer4_outputs(6092);
    layer5_outputs(5268) <= '0';
    layer5_outputs(5269) <= not((layer4_outputs(5823)) or (layer4_outputs(1019)));
    layer5_outputs(5270) <= layer4_outputs(376);
    layer5_outputs(5271) <= layer4_outputs(5342);
    layer5_outputs(5272) <= (layer4_outputs(6806)) xor (layer4_outputs(4259));
    layer5_outputs(5273) <= layer4_outputs(4008);
    layer5_outputs(5274) <= layer4_outputs(4899);
    layer5_outputs(5275) <= layer4_outputs(3192);
    layer5_outputs(5276) <= not(layer4_outputs(1987));
    layer5_outputs(5277) <= (layer4_outputs(6213)) or (layer4_outputs(357));
    layer5_outputs(5278) <= (layer4_outputs(4521)) xor (layer4_outputs(1046));
    layer5_outputs(5279) <= (layer4_outputs(1943)) and not (layer4_outputs(3027));
    layer5_outputs(5280) <= (layer4_outputs(928)) xor (layer4_outputs(5861));
    layer5_outputs(5281) <= not(layer4_outputs(751));
    layer5_outputs(5282) <= (layer4_outputs(2137)) or (layer4_outputs(107));
    layer5_outputs(5283) <= not(layer4_outputs(6884)) or (layer4_outputs(4294));
    layer5_outputs(5284) <= not(layer4_outputs(2084));
    layer5_outputs(5285) <= not(layer4_outputs(3419));
    layer5_outputs(5286) <= not(layer4_outputs(7663)) or (layer4_outputs(2097));
    layer5_outputs(5287) <= not(layer4_outputs(5683)) or (layer4_outputs(6858));
    layer5_outputs(5288) <= (layer4_outputs(3830)) or (layer4_outputs(1995));
    layer5_outputs(5289) <= not(layer4_outputs(3007));
    layer5_outputs(5290) <= not((layer4_outputs(5474)) or (layer4_outputs(5046)));
    layer5_outputs(5291) <= not(layer4_outputs(6228)) or (layer4_outputs(2022));
    layer5_outputs(5292) <= (layer4_outputs(3677)) and (layer4_outputs(2844));
    layer5_outputs(5293) <= not(layer4_outputs(1252));
    layer5_outputs(5294) <= (layer4_outputs(2491)) and not (layer4_outputs(1449));
    layer5_outputs(5295) <= layer4_outputs(893);
    layer5_outputs(5296) <= layer4_outputs(4328);
    layer5_outputs(5297) <= (layer4_outputs(3941)) and not (layer4_outputs(6008));
    layer5_outputs(5298) <= (layer4_outputs(5872)) and not (layer4_outputs(7530));
    layer5_outputs(5299) <= not(layer4_outputs(5434)) or (layer4_outputs(3350));
    layer5_outputs(5300) <= not(layer4_outputs(5303)) or (layer4_outputs(5255));
    layer5_outputs(5301) <= layer4_outputs(3335);
    layer5_outputs(5302) <= not(layer4_outputs(2210));
    layer5_outputs(5303) <= (layer4_outputs(5724)) xor (layer4_outputs(1126));
    layer5_outputs(5304) <= layer4_outputs(4494);
    layer5_outputs(5305) <= not(layer4_outputs(6928));
    layer5_outputs(5306) <= not((layer4_outputs(1853)) and (layer4_outputs(5714)));
    layer5_outputs(5307) <= layer4_outputs(7237);
    layer5_outputs(5308) <= layer4_outputs(24);
    layer5_outputs(5309) <= not(layer4_outputs(5355));
    layer5_outputs(5310) <= (layer4_outputs(1576)) and not (layer4_outputs(4975));
    layer5_outputs(5311) <= layer4_outputs(4310);
    layer5_outputs(5312) <= (layer4_outputs(1953)) xor (layer4_outputs(4398));
    layer5_outputs(5313) <= layer4_outputs(3322);
    layer5_outputs(5314) <= (layer4_outputs(6784)) xor (layer4_outputs(1798));
    layer5_outputs(5315) <= layer4_outputs(2299);
    layer5_outputs(5316) <= not(layer4_outputs(6757));
    layer5_outputs(5317) <= not(layer4_outputs(6004));
    layer5_outputs(5318) <= (layer4_outputs(5963)) and not (layer4_outputs(4157));
    layer5_outputs(5319) <= (layer4_outputs(5912)) and not (layer4_outputs(4034));
    layer5_outputs(5320) <= not(layer4_outputs(1592)) or (layer4_outputs(5193));
    layer5_outputs(5321) <= (layer4_outputs(2726)) xor (layer4_outputs(2026));
    layer5_outputs(5322) <= not((layer4_outputs(1187)) xor (layer4_outputs(3403)));
    layer5_outputs(5323) <= not(layer4_outputs(7235)) or (layer4_outputs(3170));
    layer5_outputs(5324) <= '1';
    layer5_outputs(5325) <= not(layer4_outputs(5841));
    layer5_outputs(5326) <= layer4_outputs(5549);
    layer5_outputs(5327) <= not((layer4_outputs(0)) and (layer4_outputs(732)));
    layer5_outputs(5328) <= not((layer4_outputs(1185)) xor (layer4_outputs(7197)));
    layer5_outputs(5329) <= (layer4_outputs(4298)) and not (layer4_outputs(3291));
    layer5_outputs(5330) <= not(layer4_outputs(961)) or (layer4_outputs(357));
    layer5_outputs(5331) <= (layer4_outputs(7257)) and not (layer4_outputs(4728));
    layer5_outputs(5332) <= not(layer4_outputs(7043)) or (layer4_outputs(4829));
    layer5_outputs(5333) <= not(layer4_outputs(5767)) or (layer4_outputs(3757));
    layer5_outputs(5334) <= (layer4_outputs(3791)) and not (layer4_outputs(1877));
    layer5_outputs(5335) <= layer4_outputs(3559);
    layer5_outputs(5336) <= layer4_outputs(5379);
    layer5_outputs(5337) <= not(layer4_outputs(2908)) or (layer4_outputs(3634));
    layer5_outputs(5338) <= not((layer4_outputs(2300)) xor (layer4_outputs(2049)));
    layer5_outputs(5339) <= layer4_outputs(5924);
    layer5_outputs(5340) <= not(layer4_outputs(833));
    layer5_outputs(5341) <= not(layer4_outputs(3578));
    layer5_outputs(5342) <= (layer4_outputs(3912)) xor (layer4_outputs(7095));
    layer5_outputs(5343) <= (layer4_outputs(5233)) and not (layer4_outputs(6419));
    layer5_outputs(5344) <= layer4_outputs(7169);
    layer5_outputs(5345) <= layer4_outputs(3617);
    layer5_outputs(5346) <= not((layer4_outputs(2432)) or (layer4_outputs(1927)));
    layer5_outputs(5347) <= (layer4_outputs(114)) and (layer4_outputs(7062));
    layer5_outputs(5348) <= not(layer4_outputs(1280));
    layer5_outputs(5349) <= not(layer4_outputs(1351));
    layer5_outputs(5350) <= not(layer4_outputs(6425)) or (layer4_outputs(6455));
    layer5_outputs(5351) <= not(layer4_outputs(4288));
    layer5_outputs(5352) <= layer4_outputs(3989);
    layer5_outputs(5353) <= not((layer4_outputs(1722)) and (layer4_outputs(4147)));
    layer5_outputs(5354) <= (layer4_outputs(4425)) and (layer4_outputs(4078));
    layer5_outputs(5355) <= not(layer4_outputs(6185));
    layer5_outputs(5356) <= not((layer4_outputs(6050)) and (layer4_outputs(7055)));
    layer5_outputs(5357) <= not(layer4_outputs(7233));
    layer5_outputs(5358) <= layer4_outputs(7105);
    layer5_outputs(5359) <= not((layer4_outputs(5881)) or (layer4_outputs(6366)));
    layer5_outputs(5360) <= (layer4_outputs(6207)) and not (layer4_outputs(2388));
    layer5_outputs(5361) <= (layer4_outputs(6754)) xor (layer4_outputs(5798));
    layer5_outputs(5362) <= (layer4_outputs(28)) or (layer4_outputs(2311));
    layer5_outputs(5363) <= layer4_outputs(3286);
    layer5_outputs(5364) <= not(layer4_outputs(1697));
    layer5_outputs(5365) <= (layer4_outputs(3961)) and not (layer4_outputs(3900));
    layer5_outputs(5366) <= not(layer4_outputs(6690));
    layer5_outputs(5367) <= layer4_outputs(5073);
    layer5_outputs(5368) <= not((layer4_outputs(3962)) or (layer4_outputs(4476)));
    layer5_outputs(5369) <= layer4_outputs(5583);
    layer5_outputs(5370) <= not(layer4_outputs(2928)) or (layer4_outputs(7397));
    layer5_outputs(5371) <= layer4_outputs(7462);
    layer5_outputs(5372) <= (layer4_outputs(5947)) or (layer4_outputs(2958));
    layer5_outputs(5373) <= layer4_outputs(3115);
    layer5_outputs(5374) <= not((layer4_outputs(3202)) or (layer4_outputs(1832)));
    layer5_outputs(5375) <= not(layer4_outputs(3103)) or (layer4_outputs(1891));
    layer5_outputs(5376) <= (layer4_outputs(5)) xor (layer4_outputs(4722));
    layer5_outputs(5377) <= not(layer4_outputs(6615));
    layer5_outputs(5378) <= layer4_outputs(3401);
    layer5_outputs(5379) <= layer4_outputs(206);
    layer5_outputs(5380) <= not((layer4_outputs(1921)) xor (layer4_outputs(4956)));
    layer5_outputs(5381) <= layer4_outputs(5537);
    layer5_outputs(5382) <= '1';
    layer5_outputs(5383) <= (layer4_outputs(2191)) xor (layer4_outputs(7311));
    layer5_outputs(5384) <= layer4_outputs(1701);
    layer5_outputs(5385) <= (layer4_outputs(1318)) xor (layer4_outputs(5664));
    layer5_outputs(5386) <= not(layer4_outputs(3738));
    layer5_outputs(5387) <= (layer4_outputs(6959)) and (layer4_outputs(21));
    layer5_outputs(5388) <= (layer4_outputs(3517)) xor (layer4_outputs(4052));
    layer5_outputs(5389) <= not((layer4_outputs(1556)) xor (layer4_outputs(3903)));
    layer5_outputs(5390) <= not((layer4_outputs(1283)) xor (layer4_outputs(3454)));
    layer5_outputs(5391) <= (layer4_outputs(6029)) or (layer4_outputs(1417));
    layer5_outputs(5392) <= not(layer4_outputs(2328));
    layer5_outputs(5393) <= layer4_outputs(3865);
    layer5_outputs(5394) <= '0';
    layer5_outputs(5395) <= not(layer4_outputs(4371));
    layer5_outputs(5396) <= (layer4_outputs(4942)) and not (layer4_outputs(841));
    layer5_outputs(5397) <= not(layer4_outputs(6198));
    layer5_outputs(5398) <= layer4_outputs(5302);
    layer5_outputs(5399) <= not(layer4_outputs(3171)) or (layer4_outputs(7366));
    layer5_outputs(5400) <= not(layer4_outputs(455));
    layer5_outputs(5401) <= not((layer4_outputs(5896)) xor (layer4_outputs(7124)));
    layer5_outputs(5402) <= not((layer4_outputs(4204)) or (layer4_outputs(4964)));
    layer5_outputs(5403) <= not(layer4_outputs(2735));
    layer5_outputs(5404) <= not(layer4_outputs(560)) or (layer4_outputs(4492));
    layer5_outputs(5405) <= layer4_outputs(2957);
    layer5_outputs(5406) <= layer4_outputs(4671);
    layer5_outputs(5407) <= not((layer4_outputs(551)) or (layer4_outputs(5986)));
    layer5_outputs(5408) <= layer4_outputs(5810);
    layer5_outputs(5409) <= not((layer4_outputs(2275)) xor (layer4_outputs(2866)));
    layer5_outputs(5410) <= layer4_outputs(1054);
    layer5_outputs(5411) <= not(layer4_outputs(616));
    layer5_outputs(5412) <= layer4_outputs(234);
    layer5_outputs(5413) <= not(layer4_outputs(1699));
    layer5_outputs(5414) <= layer4_outputs(7321);
    layer5_outputs(5415) <= (layer4_outputs(2310)) or (layer4_outputs(794));
    layer5_outputs(5416) <= not(layer4_outputs(2813));
    layer5_outputs(5417) <= (layer4_outputs(4385)) or (layer4_outputs(2514));
    layer5_outputs(5418) <= layer4_outputs(6095);
    layer5_outputs(5419) <= layer4_outputs(7334);
    layer5_outputs(5420) <= (layer4_outputs(2643)) or (layer4_outputs(466));
    layer5_outputs(5421) <= layer4_outputs(94);
    layer5_outputs(5422) <= not(layer4_outputs(5883));
    layer5_outputs(5423) <= (layer4_outputs(4906)) or (layer4_outputs(4756));
    layer5_outputs(5424) <= not(layer4_outputs(2788));
    layer5_outputs(5425) <= not(layer4_outputs(5540)) or (layer4_outputs(6530));
    layer5_outputs(5426) <= not((layer4_outputs(3274)) or (layer4_outputs(6426)));
    layer5_outputs(5427) <= layer4_outputs(5408);
    layer5_outputs(5428) <= not((layer4_outputs(6232)) or (layer4_outputs(1065)));
    layer5_outputs(5429) <= (layer4_outputs(2577)) or (layer4_outputs(5783));
    layer5_outputs(5430) <= not((layer4_outputs(6940)) and (layer4_outputs(4709)));
    layer5_outputs(5431) <= layer4_outputs(1744);
    layer5_outputs(5432) <= '0';
    layer5_outputs(5433) <= layer4_outputs(4917);
    layer5_outputs(5434) <= (layer4_outputs(3532)) and not (layer4_outputs(7576));
    layer5_outputs(5435) <= not((layer4_outputs(1528)) or (layer4_outputs(3217)));
    layer5_outputs(5436) <= '0';
    layer5_outputs(5437) <= not(layer4_outputs(1420));
    layer5_outputs(5438) <= (layer4_outputs(4188)) xor (layer4_outputs(7472));
    layer5_outputs(5439) <= not(layer4_outputs(2657));
    layer5_outputs(5440) <= (layer4_outputs(7219)) or (layer4_outputs(1406));
    layer5_outputs(5441) <= layer4_outputs(804);
    layer5_outputs(5442) <= not((layer4_outputs(7508)) and (layer4_outputs(3017)));
    layer5_outputs(5443) <= not(layer4_outputs(5173));
    layer5_outputs(5444) <= not(layer4_outputs(5519));
    layer5_outputs(5445) <= not((layer4_outputs(7314)) and (layer4_outputs(2381)));
    layer5_outputs(5446) <= not(layer4_outputs(4772)) or (layer4_outputs(1513));
    layer5_outputs(5447) <= not(layer4_outputs(411));
    layer5_outputs(5448) <= (layer4_outputs(782)) or (layer4_outputs(2154));
    layer5_outputs(5449) <= (layer4_outputs(5187)) or (layer4_outputs(1280));
    layer5_outputs(5450) <= layer4_outputs(3290);
    layer5_outputs(5451) <= (layer4_outputs(3609)) and not (layer4_outputs(3479));
    layer5_outputs(5452) <= not(layer4_outputs(7153));
    layer5_outputs(5453) <= not(layer4_outputs(229));
    layer5_outputs(5454) <= (layer4_outputs(7300)) and not (layer4_outputs(797));
    layer5_outputs(5455) <= not(layer4_outputs(5995));
    layer5_outputs(5456) <= not(layer4_outputs(6427));
    layer5_outputs(5457) <= not(layer4_outputs(7086));
    layer5_outputs(5458) <= (layer4_outputs(3834)) xor (layer4_outputs(1119));
    layer5_outputs(5459) <= not((layer4_outputs(5251)) xor (layer4_outputs(7113)));
    layer5_outputs(5460) <= layer4_outputs(5956);
    layer5_outputs(5461) <= not(layer4_outputs(4886));
    layer5_outputs(5462) <= layer4_outputs(6184);
    layer5_outputs(5463) <= layer4_outputs(5223);
    layer5_outputs(5464) <= '0';
    layer5_outputs(5465) <= (layer4_outputs(4807)) or (layer4_outputs(6960));
    layer5_outputs(5466) <= layer4_outputs(3450);
    layer5_outputs(5467) <= (layer4_outputs(545)) and (layer4_outputs(5826));
    layer5_outputs(5468) <= layer4_outputs(3652);
    layer5_outputs(5469) <= not(layer4_outputs(5680)) or (layer4_outputs(3610));
    layer5_outputs(5470) <= '1';
    layer5_outputs(5471) <= (layer4_outputs(5239)) xor (layer4_outputs(613));
    layer5_outputs(5472) <= not(layer4_outputs(5005));
    layer5_outputs(5473) <= (layer4_outputs(6291)) and (layer4_outputs(2990));
    layer5_outputs(5474) <= not((layer4_outputs(5566)) and (layer4_outputs(6445)));
    layer5_outputs(5475) <= layer4_outputs(3557);
    layer5_outputs(5476) <= not((layer4_outputs(3568)) and (layer4_outputs(7109)));
    layer5_outputs(5477) <= (layer4_outputs(5672)) and (layer4_outputs(990));
    layer5_outputs(5478) <= layer4_outputs(2943);
    layer5_outputs(5479) <= (layer4_outputs(4306)) xor (layer4_outputs(524));
    layer5_outputs(5480) <= layer4_outputs(7602);
    layer5_outputs(5481) <= layer4_outputs(7527);
    layer5_outputs(5482) <= layer4_outputs(3253);
    layer5_outputs(5483) <= not(layer4_outputs(5971));
    layer5_outputs(5484) <= not((layer4_outputs(7381)) xor (layer4_outputs(2007)));
    layer5_outputs(5485) <= (layer4_outputs(6337)) xor (layer4_outputs(3263));
    layer5_outputs(5486) <= not(layer4_outputs(2570));
    layer5_outputs(5487) <= layer4_outputs(982);
    layer5_outputs(5488) <= not(layer4_outputs(5550));
    layer5_outputs(5489) <= layer4_outputs(6104);
    layer5_outputs(5490) <= not(layer4_outputs(474));
    layer5_outputs(5491) <= (layer4_outputs(6756)) and (layer4_outputs(739));
    layer5_outputs(5492) <= not(layer4_outputs(6087)) or (layer4_outputs(3705));
    layer5_outputs(5493) <= not(layer4_outputs(5902));
    layer5_outputs(5494) <= not((layer4_outputs(1630)) xor (layer4_outputs(5416)));
    layer5_outputs(5495) <= (layer4_outputs(3892)) xor (layer4_outputs(3134));
    layer5_outputs(5496) <= (layer4_outputs(4085)) and not (layer4_outputs(5183));
    layer5_outputs(5497) <= layer4_outputs(1160);
    layer5_outputs(5498) <= not(layer4_outputs(764)) or (layer4_outputs(4040));
    layer5_outputs(5499) <= (layer4_outputs(1882)) and not (layer4_outputs(2109));
    layer5_outputs(5500) <= not(layer4_outputs(1445)) or (layer4_outputs(2028));
    layer5_outputs(5501) <= not((layer4_outputs(3521)) xor (layer4_outputs(2334)));
    layer5_outputs(5502) <= not(layer4_outputs(7311));
    layer5_outputs(5503) <= layer4_outputs(2614);
    layer5_outputs(5504) <= not((layer4_outputs(7100)) and (layer4_outputs(6134)));
    layer5_outputs(5505) <= layer4_outputs(7032);
    layer5_outputs(5506) <= not((layer4_outputs(1481)) or (layer4_outputs(2269)));
    layer5_outputs(5507) <= layer4_outputs(3303);
    layer5_outputs(5508) <= '1';
    layer5_outputs(5509) <= not((layer4_outputs(1212)) or (layer4_outputs(1178)));
    layer5_outputs(5510) <= not(layer4_outputs(2206)) or (layer4_outputs(7395));
    layer5_outputs(5511) <= not(layer4_outputs(3018));
    layer5_outputs(5512) <= not(layer4_outputs(434));
    layer5_outputs(5513) <= layer4_outputs(2281);
    layer5_outputs(5514) <= not(layer4_outputs(964));
    layer5_outputs(5515) <= (layer4_outputs(2540)) or (layer4_outputs(3832));
    layer5_outputs(5516) <= not((layer4_outputs(4694)) or (layer4_outputs(2070)));
    layer5_outputs(5517) <= layer4_outputs(7008);
    layer5_outputs(5518) <= not(layer4_outputs(6237));
    layer5_outputs(5519) <= layer4_outputs(1567);
    layer5_outputs(5520) <= layer4_outputs(3689);
    layer5_outputs(5521) <= not(layer4_outputs(7201));
    layer5_outputs(5522) <= not(layer4_outputs(501));
    layer5_outputs(5523) <= (layer4_outputs(165)) and not (layer4_outputs(4771));
    layer5_outputs(5524) <= layer4_outputs(5343);
    layer5_outputs(5525) <= layer4_outputs(4190);
    layer5_outputs(5526) <= layer4_outputs(2877);
    layer5_outputs(5527) <= (layer4_outputs(3975)) xor (layer4_outputs(5003));
    layer5_outputs(5528) <= '0';
    layer5_outputs(5529) <= not(layer4_outputs(542));
    layer5_outputs(5530) <= layer4_outputs(2357);
    layer5_outputs(5531) <= layer4_outputs(7298);
    layer5_outputs(5532) <= (layer4_outputs(4071)) or (layer4_outputs(5058));
    layer5_outputs(5533) <= not(layer4_outputs(2728)) or (layer4_outputs(5109));
    layer5_outputs(5534) <= (layer4_outputs(6590)) and not (layer4_outputs(4664));
    layer5_outputs(5535) <= layer4_outputs(6593);
    layer5_outputs(5536) <= layer4_outputs(5765);
    layer5_outputs(5537) <= not(layer4_outputs(6803));
    layer5_outputs(5538) <= not(layer4_outputs(3792)) or (layer4_outputs(619));
    layer5_outputs(5539) <= (layer4_outputs(4657)) xor (layer4_outputs(1131));
    layer5_outputs(5540) <= not(layer4_outputs(894));
    layer5_outputs(5541) <= not(layer4_outputs(5343));
    layer5_outputs(5542) <= layer4_outputs(61);
    layer5_outputs(5543) <= layer4_outputs(5640);
    layer5_outputs(5544) <= not((layer4_outputs(6953)) xor (layer4_outputs(4433)));
    layer5_outputs(5545) <= not(layer4_outputs(2977));
    layer5_outputs(5546) <= not((layer4_outputs(2044)) and (layer4_outputs(1504)));
    layer5_outputs(5547) <= not((layer4_outputs(5448)) and (layer4_outputs(2860)));
    layer5_outputs(5548) <= layer4_outputs(233);
    layer5_outputs(5549) <= not((layer4_outputs(5403)) and (layer4_outputs(1528)));
    layer5_outputs(5550) <= layer4_outputs(5479);
    layer5_outputs(5551) <= not(layer4_outputs(4441));
    layer5_outputs(5552) <= not(layer4_outputs(1944));
    layer5_outputs(5553) <= (layer4_outputs(7679)) or (layer4_outputs(5119));
    layer5_outputs(5554) <= not((layer4_outputs(6637)) xor (layer4_outputs(866)));
    layer5_outputs(5555) <= layer4_outputs(1418);
    layer5_outputs(5556) <= not(layer4_outputs(6093));
    layer5_outputs(5557) <= not(layer4_outputs(7433));
    layer5_outputs(5558) <= (layer4_outputs(1159)) and not (layer4_outputs(1942));
    layer5_outputs(5559) <= layer4_outputs(4547);
    layer5_outputs(5560) <= not(layer4_outputs(5418));
    layer5_outputs(5561) <= (layer4_outputs(6445)) xor (layer4_outputs(6269));
    layer5_outputs(5562) <= (layer4_outputs(2867)) and (layer4_outputs(3431));
    layer5_outputs(5563) <= not(layer4_outputs(2670));
    layer5_outputs(5564) <= not(layer4_outputs(3793)) or (layer4_outputs(1860));
    layer5_outputs(5565) <= layer4_outputs(4284);
    layer5_outputs(5566) <= (layer4_outputs(6541)) and not (layer4_outputs(3331));
    layer5_outputs(5567) <= (layer4_outputs(7098)) or (layer4_outputs(7229));
    layer5_outputs(5568) <= (layer4_outputs(6732)) and not (layer4_outputs(784));
    layer5_outputs(5569) <= layer4_outputs(4018);
    layer5_outputs(5570) <= not(layer4_outputs(7412)) or (layer4_outputs(6981));
    layer5_outputs(5571) <= layer4_outputs(6230);
    layer5_outputs(5572) <= not(layer4_outputs(1619));
    layer5_outputs(5573) <= (layer4_outputs(1544)) and not (layer4_outputs(1353));
    layer5_outputs(5574) <= layer4_outputs(1898);
    layer5_outputs(5575) <= layer4_outputs(1325);
    layer5_outputs(5576) <= layer4_outputs(5222);
    layer5_outputs(5577) <= layer4_outputs(1081);
    layer5_outputs(5578) <= not(layer4_outputs(4625));
    layer5_outputs(5579) <= not(layer4_outputs(3830));
    layer5_outputs(5580) <= not((layer4_outputs(6193)) or (layer4_outputs(3145)));
    layer5_outputs(5581) <= layer4_outputs(4440);
    layer5_outputs(5582) <= '1';
    layer5_outputs(5583) <= (layer4_outputs(5331)) and not (layer4_outputs(5135));
    layer5_outputs(5584) <= not(layer4_outputs(2877)) or (layer4_outputs(2842));
    layer5_outputs(5585) <= (layer4_outputs(5642)) and not (layer4_outputs(64));
    layer5_outputs(5586) <= layer4_outputs(2477);
    layer5_outputs(5587) <= not((layer4_outputs(7614)) or (layer4_outputs(147)));
    layer5_outputs(5588) <= not((layer4_outputs(5147)) or (layer4_outputs(6618)));
    layer5_outputs(5589) <= layer4_outputs(4198);
    layer5_outputs(5590) <= not((layer4_outputs(1197)) or (layer4_outputs(2966)));
    layer5_outputs(5591) <= not(layer4_outputs(5647));
    layer5_outputs(5592) <= (layer4_outputs(988)) and not (layer4_outputs(1343));
    layer5_outputs(5593) <= not((layer4_outputs(4096)) or (layer4_outputs(2854)));
    layer5_outputs(5594) <= (layer4_outputs(7431)) xor (layer4_outputs(4998));
    layer5_outputs(5595) <= not(layer4_outputs(3511)) or (layer4_outputs(479));
    layer5_outputs(5596) <= not(layer4_outputs(6551));
    layer5_outputs(5597) <= not(layer4_outputs(2542));
    layer5_outputs(5598) <= not((layer4_outputs(5007)) or (layer4_outputs(4343)));
    layer5_outputs(5599) <= layer4_outputs(1584);
    layer5_outputs(5600) <= '0';
    layer5_outputs(5601) <= layer4_outputs(2111);
    layer5_outputs(5602) <= not(layer4_outputs(4524)) or (layer4_outputs(1918));
    layer5_outputs(5603) <= '1';
    layer5_outputs(5604) <= not((layer4_outputs(1547)) and (layer4_outputs(514)));
    layer5_outputs(5605) <= (layer4_outputs(448)) and not (layer4_outputs(1766));
    layer5_outputs(5606) <= layer4_outputs(6630);
    layer5_outputs(5607) <= not((layer4_outputs(6635)) or (layer4_outputs(7385)));
    layer5_outputs(5608) <= not(layer4_outputs(5769)) or (layer4_outputs(1197));
    layer5_outputs(5609) <= (layer4_outputs(4970)) or (layer4_outputs(2143));
    layer5_outputs(5610) <= not(layer4_outputs(1207));
    layer5_outputs(5611) <= layer4_outputs(3778);
    layer5_outputs(5612) <= '1';
    layer5_outputs(5613) <= (layer4_outputs(1816)) or (layer4_outputs(6011));
    layer5_outputs(5614) <= not(layer4_outputs(4060));
    layer5_outputs(5615) <= not(layer4_outputs(86));
    layer5_outputs(5616) <= not((layer4_outputs(1632)) and (layer4_outputs(6605)));
    layer5_outputs(5617) <= not(layer4_outputs(6424));
    layer5_outputs(5618) <= not(layer4_outputs(585));
    layer5_outputs(5619) <= (layer4_outputs(852)) and (layer4_outputs(2906));
    layer5_outputs(5620) <= layer4_outputs(1724);
    layer5_outputs(5621) <= not(layer4_outputs(1218)) or (layer4_outputs(510));
    layer5_outputs(5622) <= not(layer4_outputs(216));
    layer5_outputs(5623) <= not(layer4_outputs(649)) or (layer4_outputs(2246));
    layer5_outputs(5624) <= not(layer4_outputs(633));
    layer5_outputs(5625) <= not(layer4_outputs(4890));
    layer5_outputs(5626) <= not(layer4_outputs(3529));
    layer5_outputs(5627) <= not((layer4_outputs(5465)) and (layer4_outputs(6160)));
    layer5_outputs(5628) <= (layer4_outputs(7398)) and not (layer4_outputs(5525));
    layer5_outputs(5629) <= layer4_outputs(5578);
    layer5_outputs(5630) <= not((layer4_outputs(7115)) or (layer4_outputs(6829)));
    layer5_outputs(5631) <= not(layer4_outputs(2537));
    layer5_outputs(5632) <= not(layer4_outputs(1740)) or (layer4_outputs(5952));
    layer5_outputs(5633) <= layer4_outputs(2454);
    layer5_outputs(5634) <= not(layer4_outputs(688));
    layer5_outputs(5635) <= not(layer4_outputs(3358)) or (layer4_outputs(4919));
    layer5_outputs(5636) <= not((layer4_outputs(7222)) xor (layer4_outputs(7404)));
    layer5_outputs(5637) <= layer4_outputs(2063);
    layer5_outputs(5638) <= not((layer4_outputs(7317)) xor (layer4_outputs(5712)));
    layer5_outputs(5639) <= not((layer4_outputs(848)) xor (layer4_outputs(3741)));
    layer5_outputs(5640) <= not(layer4_outputs(1820));
    layer5_outputs(5641) <= layer4_outputs(220);
    layer5_outputs(5642) <= layer4_outputs(7313);
    layer5_outputs(5643) <= not(layer4_outputs(3749));
    layer5_outputs(5644) <= (layer4_outputs(6012)) xor (layer4_outputs(2576));
    layer5_outputs(5645) <= not((layer4_outputs(1775)) or (layer4_outputs(3611)));
    layer5_outputs(5646) <= layer4_outputs(323);
    layer5_outputs(5647) <= layer4_outputs(5428);
    layer5_outputs(5648) <= layer4_outputs(4379);
    layer5_outputs(5649) <= not((layer4_outputs(7279)) xor (layer4_outputs(1142)));
    layer5_outputs(5650) <= not(layer4_outputs(485));
    layer5_outputs(5651) <= layer4_outputs(4957);
    layer5_outputs(5652) <= not(layer4_outputs(6790));
    layer5_outputs(5653) <= layer4_outputs(5877);
    layer5_outputs(5654) <= not(layer4_outputs(2270));
    layer5_outputs(5655) <= layer4_outputs(1131);
    layer5_outputs(5656) <= layer4_outputs(7637);
    layer5_outputs(5657) <= not(layer4_outputs(896));
    layer5_outputs(5658) <= (layer4_outputs(2575)) or (layer4_outputs(4103));
    layer5_outputs(5659) <= not(layer4_outputs(1519));
    layer5_outputs(5660) <= not(layer4_outputs(5132));
    layer5_outputs(5661) <= not(layer4_outputs(3008)) or (layer4_outputs(5568));
    layer5_outputs(5662) <= layer4_outputs(7031);
    layer5_outputs(5663) <= not((layer4_outputs(1166)) and (layer4_outputs(1866)));
    layer5_outputs(5664) <= (layer4_outputs(5817)) and (layer4_outputs(4815));
    layer5_outputs(5665) <= '0';
    layer5_outputs(5666) <= not((layer4_outputs(153)) and (layer4_outputs(1695)));
    layer5_outputs(5667) <= (layer4_outputs(455)) and not (layer4_outputs(4651));
    layer5_outputs(5668) <= layer4_outputs(1441);
    layer5_outputs(5669) <= layer4_outputs(2356);
    layer5_outputs(5670) <= (layer4_outputs(380)) xor (layer4_outputs(559));
    layer5_outputs(5671) <= not((layer4_outputs(6369)) and (layer4_outputs(1423)));
    layer5_outputs(5672) <= '0';
    layer5_outputs(5673) <= '1';
    layer5_outputs(5674) <= layer4_outputs(4167);
    layer5_outputs(5675) <= layer4_outputs(6773);
    layer5_outputs(5676) <= not((layer4_outputs(3777)) or (layer4_outputs(1089)));
    layer5_outputs(5677) <= layer4_outputs(2450);
    layer5_outputs(5678) <= (layer4_outputs(731)) and not (layer4_outputs(4368));
    layer5_outputs(5679) <= not((layer4_outputs(6608)) and (layer4_outputs(3688)));
    layer5_outputs(5680) <= '1';
    layer5_outputs(5681) <= not(layer4_outputs(1901));
    layer5_outputs(5682) <= layer4_outputs(4891);
    layer5_outputs(5683) <= (layer4_outputs(673)) and (layer4_outputs(5191));
    layer5_outputs(5684) <= not(layer4_outputs(6703));
    layer5_outputs(5685) <= layer4_outputs(4753);
    layer5_outputs(5686) <= not((layer4_outputs(2507)) xor (layer4_outputs(2336)));
    layer5_outputs(5687) <= layer4_outputs(753);
    layer5_outputs(5688) <= (layer4_outputs(3344)) xor (layer4_outputs(3184));
    layer5_outputs(5689) <= layer4_outputs(221);
    layer5_outputs(5690) <= not((layer4_outputs(1285)) and (layer4_outputs(1720)));
    layer5_outputs(5691) <= not((layer4_outputs(3219)) or (layer4_outputs(1505)));
    layer5_outputs(5692) <= layer4_outputs(3297);
    layer5_outputs(5693) <= not((layer4_outputs(4594)) or (layer4_outputs(2879)));
    layer5_outputs(5694) <= (layer4_outputs(6105)) and not (layer4_outputs(5180));
    layer5_outputs(5695) <= layer4_outputs(2530);
    layer5_outputs(5696) <= not((layer4_outputs(6900)) and (layer4_outputs(2477)));
    layer5_outputs(5697) <= not((layer4_outputs(4756)) or (layer4_outputs(6996)));
    layer5_outputs(5698) <= not((layer4_outputs(4965)) and (layer4_outputs(7590)));
    layer5_outputs(5699) <= not((layer4_outputs(5447)) or (layer4_outputs(4081)));
    layer5_outputs(5700) <= not(layer4_outputs(5135)) or (layer4_outputs(4092));
    layer5_outputs(5701) <= layer4_outputs(2428);
    layer5_outputs(5702) <= (layer4_outputs(2715)) and (layer4_outputs(4439));
    layer5_outputs(5703) <= not((layer4_outputs(4766)) and (layer4_outputs(2566)));
    layer5_outputs(5704) <= not(layer4_outputs(6452));
    layer5_outputs(5705) <= layer4_outputs(5357);
    layer5_outputs(5706) <= (layer4_outputs(1562)) or (layer4_outputs(557));
    layer5_outputs(5707) <= not(layer4_outputs(6749));
    layer5_outputs(5708) <= '1';
    layer5_outputs(5709) <= layer4_outputs(2599);
    layer5_outputs(5710) <= layer4_outputs(7666);
    layer5_outputs(5711) <= (layer4_outputs(7247)) or (layer4_outputs(4304));
    layer5_outputs(5712) <= (layer4_outputs(2656)) and (layer4_outputs(995));
    layer5_outputs(5713) <= not(layer4_outputs(4269));
    layer5_outputs(5714) <= layer4_outputs(7577);
    layer5_outputs(5715) <= not(layer4_outputs(5497));
    layer5_outputs(5716) <= not(layer4_outputs(6367));
    layer5_outputs(5717) <= not((layer4_outputs(6610)) xor (layer4_outputs(3501)));
    layer5_outputs(5718) <= not((layer4_outputs(3989)) xor (layer4_outputs(4956)));
    layer5_outputs(5719) <= (layer4_outputs(966)) or (layer4_outputs(4567));
    layer5_outputs(5720) <= layer4_outputs(2847);
    layer5_outputs(5721) <= (layer4_outputs(6060)) and not (layer4_outputs(3235));
    layer5_outputs(5722) <= not(layer4_outputs(869));
    layer5_outputs(5723) <= not(layer4_outputs(6870));
    layer5_outputs(5724) <= not(layer4_outputs(3680));
    layer5_outputs(5725) <= (layer4_outputs(3855)) and not (layer4_outputs(2821));
    layer5_outputs(5726) <= layer4_outputs(1814);
    layer5_outputs(5727) <= layer4_outputs(2176);
    layer5_outputs(5728) <= (layer4_outputs(1205)) and (layer4_outputs(2722));
    layer5_outputs(5729) <= not(layer4_outputs(655));
    layer5_outputs(5730) <= layer4_outputs(1410);
    layer5_outputs(5731) <= not(layer4_outputs(414)) or (layer4_outputs(5864));
    layer5_outputs(5732) <= layer4_outputs(1001);
    layer5_outputs(5733) <= not(layer4_outputs(2565));
    layer5_outputs(5734) <= layer4_outputs(4893);
    layer5_outputs(5735) <= (layer4_outputs(5347)) and (layer4_outputs(1045));
    layer5_outputs(5736) <= not((layer4_outputs(1268)) xor (layer4_outputs(4000)));
    layer5_outputs(5737) <= not(layer4_outputs(1557));
    layer5_outputs(5738) <= (layer4_outputs(6583)) or (layer4_outputs(3213));
    layer5_outputs(5739) <= layer4_outputs(6829);
    layer5_outputs(5740) <= not(layer4_outputs(6784));
    layer5_outputs(5741) <= layer4_outputs(1519);
    layer5_outputs(5742) <= not(layer4_outputs(3978));
    layer5_outputs(5743) <= layer4_outputs(4558);
    layer5_outputs(5744) <= not(layer4_outputs(2066)) or (layer4_outputs(3658));
    layer5_outputs(5745) <= layer4_outputs(3600);
    layer5_outputs(5746) <= not(layer4_outputs(3409));
    layer5_outputs(5747) <= not((layer4_outputs(5399)) and (layer4_outputs(1965)));
    layer5_outputs(5748) <= layer4_outputs(1032);
    layer5_outputs(5749) <= (layer4_outputs(2376)) or (layer4_outputs(2037));
    layer5_outputs(5750) <= (layer4_outputs(2521)) xor (layer4_outputs(2710));
    layer5_outputs(5751) <= not((layer4_outputs(3735)) or (layer4_outputs(1358)));
    layer5_outputs(5752) <= not(layer4_outputs(5465));
    layer5_outputs(5753) <= '0';
    layer5_outputs(5754) <= layer4_outputs(6721);
    layer5_outputs(5755) <= not(layer4_outputs(1946));
    layer5_outputs(5756) <= '1';
    layer5_outputs(5757) <= not(layer4_outputs(7279));
    layer5_outputs(5758) <= layer4_outputs(6398);
    layer5_outputs(5759) <= not(layer4_outputs(408)) or (layer4_outputs(6785));
    layer5_outputs(5760) <= not((layer4_outputs(6907)) xor (layer4_outputs(4420)));
    layer5_outputs(5761) <= not(layer4_outputs(6905)) or (layer4_outputs(2315));
    layer5_outputs(5762) <= (layer4_outputs(1980)) and not (layer4_outputs(2655));
    layer5_outputs(5763) <= (layer4_outputs(843)) and not (layer4_outputs(3005));
    layer5_outputs(5764) <= not(layer4_outputs(3234));
    layer5_outputs(5765) <= layer4_outputs(680);
    layer5_outputs(5766) <= not((layer4_outputs(2822)) or (layer4_outputs(4210)));
    layer5_outputs(5767) <= (layer4_outputs(714)) or (layer4_outputs(969));
    layer5_outputs(5768) <= layer4_outputs(1025);
    layer5_outputs(5769) <= (layer4_outputs(2015)) and not (layer4_outputs(1582));
    layer5_outputs(5770) <= (layer4_outputs(2941)) xor (layer4_outputs(2146));
    layer5_outputs(5771) <= not(layer4_outputs(2555));
    layer5_outputs(5772) <= (layer4_outputs(6700)) and (layer4_outputs(5152));
    layer5_outputs(5773) <= not(layer4_outputs(1808));
    layer5_outputs(5774) <= (layer4_outputs(3061)) xor (layer4_outputs(7471));
    layer5_outputs(5775) <= (layer4_outputs(677)) or (layer4_outputs(6247));
    layer5_outputs(5776) <= not(layer4_outputs(2271));
    layer5_outputs(5777) <= not(layer4_outputs(5380));
    layer5_outputs(5778) <= layer4_outputs(1714);
    layer5_outputs(5779) <= not(layer4_outputs(3761)) or (layer4_outputs(7284));
    layer5_outputs(5780) <= (layer4_outputs(1897)) and not (layer4_outputs(7192));
    layer5_outputs(5781) <= layer4_outputs(4843);
    layer5_outputs(5782) <= layer4_outputs(7286);
    layer5_outputs(5783) <= (layer4_outputs(915)) and not (layer4_outputs(483));
    layer5_outputs(5784) <= not(layer4_outputs(281));
    layer5_outputs(5785) <= not((layer4_outputs(6005)) xor (layer4_outputs(6851)));
    layer5_outputs(5786) <= not((layer4_outputs(792)) xor (layer4_outputs(3606)));
    layer5_outputs(5787) <= layer4_outputs(7577);
    layer5_outputs(5788) <= (layer4_outputs(473)) and not (layer4_outputs(606));
    layer5_outputs(5789) <= not(layer4_outputs(4503));
    layer5_outputs(5790) <= not(layer4_outputs(1480));
    layer5_outputs(5791) <= (layer4_outputs(1966)) or (layer4_outputs(4747));
    layer5_outputs(5792) <= not(layer4_outputs(6780));
    layer5_outputs(5793) <= not((layer4_outputs(3384)) and (layer4_outputs(2504)));
    layer5_outputs(5794) <= (layer4_outputs(2197)) and (layer4_outputs(818));
    layer5_outputs(5795) <= not(layer4_outputs(4801));
    layer5_outputs(5796) <= not(layer4_outputs(6168));
    layer5_outputs(5797) <= (layer4_outputs(4796)) and (layer4_outputs(5116));
    layer5_outputs(5798) <= not(layer4_outputs(6715));
    layer5_outputs(5799) <= layer4_outputs(6447);
    layer5_outputs(5800) <= '1';
    layer5_outputs(5801) <= not(layer4_outputs(2771));
    layer5_outputs(5802) <= not(layer4_outputs(5126));
    layer5_outputs(5803) <= not((layer4_outputs(1657)) and (layer4_outputs(2424)));
    layer5_outputs(5804) <= not((layer4_outputs(2029)) xor (layer4_outputs(4100)));
    layer5_outputs(5805) <= (layer4_outputs(1311)) xor (layer4_outputs(2151));
    layer5_outputs(5806) <= layer4_outputs(1227);
    layer5_outputs(5807) <= (layer4_outputs(138)) or (layer4_outputs(2278));
    layer5_outputs(5808) <= not(layer4_outputs(5556)) or (layer4_outputs(2229));
    layer5_outputs(5809) <= layer4_outputs(2054);
    layer5_outputs(5810) <= layer4_outputs(7599);
    layer5_outputs(5811) <= (layer4_outputs(5233)) and not (layer4_outputs(4738));
    layer5_outputs(5812) <= layer4_outputs(4454);
    layer5_outputs(5813) <= not(layer4_outputs(7269));
    layer5_outputs(5814) <= layer4_outputs(1198);
    layer5_outputs(5815) <= '1';
    layer5_outputs(5816) <= layer4_outputs(3902);
    layer5_outputs(5817) <= not(layer4_outputs(4757)) or (layer4_outputs(7556));
    layer5_outputs(5818) <= (layer4_outputs(4643)) and not (layer4_outputs(7180));
    layer5_outputs(5819) <= not(layer4_outputs(917)) or (layer4_outputs(6745));
    layer5_outputs(5820) <= not((layer4_outputs(5588)) and (layer4_outputs(7055)));
    layer5_outputs(5821) <= not(layer4_outputs(6534));
    layer5_outputs(5822) <= not(layer4_outputs(3147));
    layer5_outputs(5823) <= (layer4_outputs(3371)) xor (layer4_outputs(671));
    layer5_outputs(5824) <= not(layer4_outputs(425));
    layer5_outputs(5825) <= not(layer4_outputs(562)) or (layer4_outputs(3146));
    layer5_outputs(5826) <= not(layer4_outputs(1521));
    layer5_outputs(5827) <= layer4_outputs(7234);
    layer5_outputs(5828) <= (layer4_outputs(1062)) xor (layer4_outputs(4418));
    layer5_outputs(5829) <= not(layer4_outputs(6601));
    layer5_outputs(5830) <= (layer4_outputs(4653)) and (layer4_outputs(4387));
    layer5_outputs(5831) <= (layer4_outputs(1329)) and (layer4_outputs(2622));
    layer5_outputs(5832) <= not(layer4_outputs(1629)) or (layer4_outputs(4884));
    layer5_outputs(5833) <= layer4_outputs(5714);
    layer5_outputs(5834) <= not(layer4_outputs(6994));
    layer5_outputs(5835) <= layer4_outputs(1252);
    layer5_outputs(5836) <= not((layer4_outputs(6650)) and (layer4_outputs(5667)));
    layer5_outputs(5837) <= not((layer4_outputs(2504)) or (layer4_outputs(3194)));
    layer5_outputs(5838) <= not(layer4_outputs(5794));
    layer5_outputs(5839) <= layer4_outputs(3582);
    layer5_outputs(5840) <= layer4_outputs(6364);
    layer5_outputs(5841) <= not(layer4_outputs(4549));
    layer5_outputs(5842) <= not((layer4_outputs(4254)) or (layer4_outputs(1236)));
    layer5_outputs(5843) <= layer4_outputs(2686);
    layer5_outputs(5844) <= (layer4_outputs(7283)) and not (layer4_outputs(1266));
    layer5_outputs(5845) <= not(layer4_outputs(4997));
    layer5_outputs(5846) <= layer4_outputs(2200);
    layer5_outputs(5847) <= (layer4_outputs(2885)) and not (layer4_outputs(3768));
    layer5_outputs(5848) <= (layer4_outputs(3410)) and not (layer4_outputs(2080));
    layer5_outputs(5849) <= layer4_outputs(6262);
    layer5_outputs(5850) <= (layer4_outputs(4690)) xor (layer4_outputs(6814));
    layer5_outputs(5851) <= not(layer4_outputs(223));
    layer5_outputs(5852) <= layer4_outputs(88);
    layer5_outputs(5853) <= layer4_outputs(1596);
    layer5_outputs(5854) <= layer4_outputs(1467);
    layer5_outputs(5855) <= not(layer4_outputs(1626)) or (layer4_outputs(170));
    layer5_outputs(5856) <= layer4_outputs(2114);
    layer5_outputs(5857) <= not(layer4_outputs(17));
    layer5_outputs(5858) <= layer4_outputs(5047);
    layer5_outputs(5859) <= not((layer4_outputs(1841)) and (layer4_outputs(3553)));
    layer5_outputs(5860) <= not(layer4_outputs(1656));
    layer5_outputs(5861) <= layer4_outputs(2248);
    layer5_outputs(5862) <= layer4_outputs(287);
    layer5_outputs(5863) <= (layer4_outputs(4550)) and (layer4_outputs(5082));
    layer5_outputs(5864) <= not(layer4_outputs(7080));
    layer5_outputs(5865) <= '1';
    layer5_outputs(5866) <= '0';
    layer5_outputs(5867) <= (layer4_outputs(1526)) xor (layer4_outputs(4630));
    layer5_outputs(5868) <= not(layer4_outputs(1400));
    layer5_outputs(5869) <= (layer4_outputs(4962)) or (layer4_outputs(1335));
    layer5_outputs(5870) <= not(layer4_outputs(2714));
    layer5_outputs(5871) <= layer4_outputs(7514);
    layer5_outputs(5872) <= not((layer4_outputs(1415)) and (layer4_outputs(7499)));
    layer5_outputs(5873) <= layer4_outputs(3206);
    layer5_outputs(5874) <= (layer4_outputs(17)) and not (layer4_outputs(6657));
    layer5_outputs(5875) <= (layer4_outputs(7288)) or (layer4_outputs(850));
    layer5_outputs(5876) <= layer4_outputs(2295);
    layer5_outputs(5877) <= not(layer4_outputs(5262)) or (layer4_outputs(2427));
    layer5_outputs(5878) <= layer4_outputs(737);
    layer5_outputs(5879) <= not((layer4_outputs(2620)) and (layer4_outputs(3393)));
    layer5_outputs(5880) <= not(layer4_outputs(5773));
    layer5_outputs(5881) <= not(layer4_outputs(4291));
    layer5_outputs(5882) <= not((layer4_outputs(3499)) or (layer4_outputs(5106)));
    layer5_outputs(5883) <= layer4_outputs(5019);
    layer5_outputs(5884) <= (layer4_outputs(4369)) and not (layer4_outputs(5929));
    layer5_outputs(5885) <= not(layer4_outputs(635));
    layer5_outputs(5886) <= not((layer4_outputs(3590)) or (layer4_outputs(7535)));
    layer5_outputs(5887) <= '1';
    layer5_outputs(5888) <= not(layer4_outputs(6142));
    layer5_outputs(5889) <= (layer4_outputs(2674)) and not (layer4_outputs(4347));
    layer5_outputs(5890) <= not(layer4_outputs(953));
    layer5_outputs(5891) <= layer4_outputs(146);
    layer5_outputs(5892) <= not((layer4_outputs(2123)) or (layer4_outputs(4740)));
    layer5_outputs(5893) <= layer4_outputs(25);
    layer5_outputs(5894) <= not(layer4_outputs(2551));
    layer5_outputs(5895) <= (layer4_outputs(6024)) xor (layer4_outputs(1906));
    layer5_outputs(5896) <= (layer4_outputs(1542)) xor (layer4_outputs(3927));
    layer5_outputs(5897) <= not((layer4_outputs(5884)) xor (layer4_outputs(4063)));
    layer5_outputs(5898) <= (layer4_outputs(2421)) xor (layer4_outputs(638));
    layer5_outputs(5899) <= not((layer4_outputs(2418)) or (layer4_outputs(3115)));
    layer5_outputs(5900) <= not(layer4_outputs(1789));
    layer5_outputs(5901) <= not(layer4_outputs(7642)) or (layer4_outputs(1438));
    layer5_outputs(5902) <= not(layer4_outputs(6578));
    layer5_outputs(5903) <= not(layer4_outputs(3577));
    layer5_outputs(5904) <= not(layer4_outputs(6310));
    layer5_outputs(5905) <= not(layer4_outputs(2875));
    layer5_outputs(5906) <= '1';
    layer5_outputs(5907) <= not(layer4_outputs(6187));
    layer5_outputs(5908) <= not(layer4_outputs(1589));
    layer5_outputs(5909) <= layer4_outputs(1759);
    layer5_outputs(5910) <= layer4_outputs(2793);
    layer5_outputs(5911) <= (layer4_outputs(6741)) and (layer4_outputs(1955));
    layer5_outputs(5912) <= layer4_outputs(6660);
    layer5_outputs(5913) <= not(layer4_outputs(1360));
    layer5_outputs(5914) <= (layer4_outputs(1539)) and (layer4_outputs(5217));
    layer5_outputs(5915) <= not(layer4_outputs(5782));
    layer5_outputs(5916) <= not((layer4_outputs(2917)) xor (layer4_outputs(7379)));
    layer5_outputs(5917) <= not((layer4_outputs(338)) or (layer4_outputs(3217)));
    layer5_outputs(5918) <= not((layer4_outputs(2416)) and (layer4_outputs(1154)));
    layer5_outputs(5919) <= not(layer4_outputs(4080)) or (layer4_outputs(3972));
    layer5_outputs(5920) <= '1';
    layer5_outputs(5921) <= layer4_outputs(7094);
    layer5_outputs(5922) <= layer4_outputs(6234);
    layer5_outputs(5923) <= layer4_outputs(3398);
    layer5_outputs(5924) <= not(layer4_outputs(6662));
    layer5_outputs(5925) <= layer4_outputs(5747);
    layer5_outputs(5926) <= (layer4_outputs(924)) and not (layer4_outputs(1692));
    layer5_outputs(5927) <= not((layer4_outputs(5848)) xor (layer4_outputs(1356)));
    layer5_outputs(5928) <= not(layer4_outputs(6367)) or (layer4_outputs(1846));
    layer5_outputs(5929) <= (layer4_outputs(7200)) and (layer4_outputs(7356));
    layer5_outputs(5930) <= layer4_outputs(7419);
    layer5_outputs(5931) <= not(layer4_outputs(5366));
    layer5_outputs(5932) <= not(layer4_outputs(5944)) or (layer4_outputs(3959));
    layer5_outputs(5933) <= not(layer4_outputs(7605));
    layer5_outputs(5934) <= not(layer4_outputs(4689));
    layer5_outputs(5935) <= not((layer4_outputs(880)) and (layer4_outputs(4666)));
    layer5_outputs(5936) <= not(layer4_outputs(1634));
    layer5_outputs(5937) <= layer4_outputs(1259);
    layer5_outputs(5938) <= not(layer4_outputs(2177)) or (layer4_outputs(7092));
    layer5_outputs(5939) <= layer4_outputs(7000);
    layer5_outputs(5940) <= layer4_outputs(6100);
    layer5_outputs(5941) <= (layer4_outputs(4007)) xor (layer4_outputs(5424));
    layer5_outputs(5942) <= (layer4_outputs(4896)) and (layer4_outputs(4593));
    layer5_outputs(5943) <= layer4_outputs(4710);
    layer5_outputs(5944) <= not(layer4_outputs(5925));
    layer5_outputs(5945) <= not(layer4_outputs(3527)) or (layer4_outputs(6903));
    layer5_outputs(5946) <= layer4_outputs(3910);
    layer5_outputs(5947) <= layer4_outputs(2290);
    layer5_outputs(5948) <= not(layer4_outputs(7341)) or (layer4_outputs(4394));
    layer5_outputs(5949) <= (layer4_outputs(5000)) and not (layer4_outputs(603));
    layer5_outputs(5950) <= not(layer4_outputs(6245));
    layer5_outputs(5951) <= (layer4_outputs(847)) and (layer4_outputs(4786));
    layer5_outputs(5952) <= (layer4_outputs(6032)) and not (layer4_outputs(6087));
    layer5_outputs(5953) <= (layer4_outputs(4944)) and not (layer4_outputs(3558));
    layer5_outputs(5954) <= (layer4_outputs(4415)) and (layer4_outputs(2624));
    layer5_outputs(5955) <= not(layer4_outputs(362));
    layer5_outputs(5956) <= not(layer4_outputs(7546));
    layer5_outputs(5957) <= layer4_outputs(1198);
    layer5_outputs(5958) <= not((layer4_outputs(5112)) or (layer4_outputs(1524)));
    layer5_outputs(5959) <= not(layer4_outputs(4590));
    layer5_outputs(5960) <= layer4_outputs(3452);
    layer5_outputs(5961) <= (layer4_outputs(4604)) or (layer4_outputs(3902));
    layer5_outputs(5962) <= layer4_outputs(6206);
    layer5_outputs(5963) <= not(layer4_outputs(3655));
    layer5_outputs(5964) <= layer4_outputs(6594);
    layer5_outputs(5965) <= (layer4_outputs(7446)) and (layer4_outputs(7020));
    layer5_outputs(5966) <= not(layer4_outputs(143)) or (layer4_outputs(7221));
    layer5_outputs(5967) <= not((layer4_outputs(2874)) or (layer4_outputs(1208)));
    layer5_outputs(5968) <= not(layer4_outputs(7559));
    layer5_outputs(5969) <= not(layer4_outputs(5665));
    layer5_outputs(5970) <= (layer4_outputs(4823)) and not (layer4_outputs(6139));
    layer5_outputs(5971) <= not((layer4_outputs(4842)) xor (layer4_outputs(3256)));
    layer5_outputs(5972) <= '1';
    layer5_outputs(5973) <= not(layer4_outputs(6759));
    layer5_outputs(5974) <= (layer4_outputs(389)) and not (layer4_outputs(6200));
    layer5_outputs(5975) <= not(layer4_outputs(6797));
    layer5_outputs(5976) <= not(layer4_outputs(7222));
    layer5_outputs(5977) <= (layer4_outputs(7455)) xor (layer4_outputs(3490));
    layer5_outputs(5978) <= not((layer4_outputs(5243)) or (layer4_outputs(6787)));
    layer5_outputs(5979) <= '0';
    layer5_outputs(5980) <= layer4_outputs(1391);
    layer5_outputs(5981) <= (layer4_outputs(6178)) or (layer4_outputs(317));
    layer5_outputs(5982) <= (layer4_outputs(3503)) or (layer4_outputs(682));
    layer5_outputs(5983) <= not(layer4_outputs(134));
    layer5_outputs(5984) <= (layer4_outputs(797)) or (layer4_outputs(6836));
    layer5_outputs(5985) <= layer4_outputs(5226);
    layer5_outputs(5986) <= not((layer4_outputs(747)) and (layer4_outputs(4804)));
    layer5_outputs(5987) <= layer4_outputs(332);
    layer5_outputs(5988) <= not(layer4_outputs(1395)) or (layer4_outputs(45));
    layer5_outputs(5989) <= (layer4_outputs(3866)) and not (layer4_outputs(5574));
    layer5_outputs(5990) <= (layer4_outputs(468)) and not (layer4_outputs(1601));
    layer5_outputs(5991) <= (layer4_outputs(1639)) and (layer4_outputs(4637));
    layer5_outputs(5992) <= '1';
    layer5_outputs(5993) <= not(layer4_outputs(6628));
    layer5_outputs(5994) <= '1';
    layer5_outputs(5995) <= not(layer4_outputs(6706));
    layer5_outputs(5996) <= not((layer4_outputs(5500)) and (layer4_outputs(1831)));
    layer5_outputs(5997) <= not((layer4_outputs(6902)) or (layer4_outputs(2924)));
    layer5_outputs(5998) <= not(layer4_outputs(1989));
    layer5_outputs(5999) <= (layer4_outputs(1169)) and (layer4_outputs(3404));
    layer5_outputs(6000) <= '1';
    layer5_outputs(6001) <= (layer4_outputs(6328)) or (layer4_outputs(4207));
    layer5_outputs(6002) <= not(layer4_outputs(2910)) or (layer4_outputs(6760));
    layer5_outputs(6003) <= (layer4_outputs(4879)) or (layer4_outputs(3946));
    layer5_outputs(6004) <= not(layer4_outputs(47));
    layer5_outputs(6005) <= not(layer4_outputs(2752));
    layer5_outputs(6006) <= not((layer4_outputs(4821)) or (layer4_outputs(1057)));
    layer5_outputs(6007) <= not(layer4_outputs(3948));
    layer5_outputs(6008) <= layer4_outputs(698);
    layer5_outputs(6009) <= not(layer4_outputs(7365));
    layer5_outputs(6010) <= '0';
    layer5_outputs(6011) <= layer4_outputs(233);
    layer5_outputs(6012) <= not(layer4_outputs(6895));
    layer5_outputs(6013) <= not(layer4_outputs(6912));
    layer5_outputs(6014) <= layer4_outputs(5216);
    layer5_outputs(6015) <= not(layer4_outputs(1912));
    layer5_outputs(6016) <= layer4_outputs(4433);
    layer5_outputs(6017) <= not(layer4_outputs(2973));
    layer5_outputs(6018) <= not(layer4_outputs(6915));
    layer5_outputs(6019) <= (layer4_outputs(125)) and not (layer4_outputs(1332));
    layer5_outputs(6020) <= not((layer4_outputs(974)) and (layer4_outputs(5420)));
    layer5_outputs(6021) <= (layer4_outputs(6558)) and not (layer4_outputs(1181));
    layer5_outputs(6022) <= (layer4_outputs(3755)) xor (layer4_outputs(5380));
    layer5_outputs(6023) <= layer4_outputs(4084);
    layer5_outputs(6024) <= layer4_outputs(1057);
    layer5_outputs(6025) <= not(layer4_outputs(7306)) or (layer4_outputs(7175));
    layer5_outputs(6026) <= (layer4_outputs(1296)) or (layer4_outputs(6049));
    layer5_outputs(6027) <= not(layer4_outputs(7627));
    layer5_outputs(6028) <= not(layer4_outputs(6223)) or (layer4_outputs(6164));
    layer5_outputs(6029) <= not(layer4_outputs(1735));
    layer5_outputs(6030) <= layer4_outputs(5957);
    layer5_outputs(6031) <= layer4_outputs(277);
    layer5_outputs(6032) <= layer4_outputs(849);
    layer5_outputs(6033) <= layer4_outputs(1104);
    layer5_outputs(6034) <= (layer4_outputs(5252)) xor (layer4_outputs(4430));
    layer5_outputs(6035) <= (layer4_outputs(5939)) xor (layer4_outputs(6740));
    layer5_outputs(6036) <= not(layer4_outputs(2633)) or (layer4_outputs(5012));
    layer5_outputs(6037) <= layer4_outputs(2786);
    layer5_outputs(6038) <= not((layer4_outputs(6047)) xor (layer4_outputs(4913)));
    layer5_outputs(6039) <= (layer4_outputs(7491)) or (layer4_outputs(7167));
    layer5_outputs(6040) <= (layer4_outputs(5080)) and not (layer4_outputs(5160));
    layer5_outputs(6041) <= (layer4_outputs(1644)) or (layer4_outputs(4865));
    layer5_outputs(6042) <= layer4_outputs(3427);
    layer5_outputs(6043) <= (layer4_outputs(5264)) xor (layer4_outputs(7637));
    layer5_outputs(6044) <= not(layer4_outputs(1786));
    layer5_outputs(6045) <= not(layer4_outputs(6098));
    layer5_outputs(6046) <= not(layer4_outputs(1215));
    layer5_outputs(6047) <= not((layer4_outputs(3141)) xor (layer4_outputs(5994)));
    layer5_outputs(6048) <= layer4_outputs(2082);
    layer5_outputs(6049) <= (layer4_outputs(1716)) or (layer4_outputs(3906));
    layer5_outputs(6050) <= (layer4_outputs(4960)) and (layer4_outputs(634));
    layer5_outputs(6051) <= not((layer4_outputs(1097)) xor (layer4_outputs(6067)));
    layer5_outputs(6052) <= not(layer4_outputs(3073));
    layer5_outputs(6053) <= layer4_outputs(2897);
    layer5_outputs(6054) <= not(layer4_outputs(1407));
    layer5_outputs(6055) <= not(layer4_outputs(4296));
    layer5_outputs(6056) <= not(layer4_outputs(226));
    layer5_outputs(6057) <= layer4_outputs(4619);
    layer5_outputs(6058) <= not(layer4_outputs(2080));
    layer5_outputs(6059) <= layer4_outputs(6094);
    layer5_outputs(6060) <= not((layer4_outputs(6157)) xor (layer4_outputs(4046)));
    layer5_outputs(6061) <= (layer4_outputs(4127)) and not (layer4_outputs(2538));
    layer5_outputs(6062) <= not(layer4_outputs(707));
    layer5_outputs(6063) <= not((layer4_outputs(1740)) xor (layer4_outputs(5527)));
    layer5_outputs(6064) <= (layer4_outputs(1511)) and not (layer4_outputs(5341));
    layer5_outputs(6065) <= layer4_outputs(4507);
    layer5_outputs(6066) <= '0';
    layer5_outputs(6067) <= (layer4_outputs(865)) xor (layer4_outputs(3583));
    layer5_outputs(6068) <= layer4_outputs(2579);
    layer5_outputs(6069) <= not((layer4_outputs(5899)) xor (layer4_outputs(46)));
    layer5_outputs(6070) <= layer4_outputs(5008);
    layer5_outputs(6071) <= layer4_outputs(3495);
    layer5_outputs(6072) <= '0';
    layer5_outputs(6073) <= layer4_outputs(3221);
    layer5_outputs(6074) <= not((layer4_outputs(4730)) and (layer4_outputs(3177)));
    layer5_outputs(6075) <= layer4_outputs(2236);
    layer5_outputs(6076) <= not((layer4_outputs(2304)) xor (layer4_outputs(4678)));
    layer5_outputs(6077) <= not(layer4_outputs(4933));
    layer5_outputs(6078) <= layer4_outputs(2303);
    layer5_outputs(6079) <= (layer4_outputs(2223)) and not (layer4_outputs(1352));
    layer5_outputs(6080) <= not((layer4_outputs(984)) or (layer4_outputs(4889)));
    layer5_outputs(6081) <= not(layer4_outputs(1028)) or (layer4_outputs(1922));
    layer5_outputs(6082) <= layer4_outputs(3470);
    layer5_outputs(6083) <= layer4_outputs(2957);
    layer5_outputs(6084) <= (layer4_outputs(2128)) xor (layer4_outputs(1282));
    layer5_outputs(6085) <= (layer4_outputs(4794)) and not (layer4_outputs(1263));
    layer5_outputs(6086) <= (layer4_outputs(52)) xor (layer4_outputs(1715));
    layer5_outputs(6087) <= layer4_outputs(2212);
    layer5_outputs(6088) <= layer4_outputs(5241);
    layer5_outputs(6089) <= layer4_outputs(6844);
    layer5_outputs(6090) <= layer4_outputs(5668);
    layer5_outputs(6091) <= not(layer4_outputs(4329)) or (layer4_outputs(1848));
    layer5_outputs(6092) <= layer4_outputs(2008);
    layer5_outputs(6093) <= not(layer4_outputs(1561));
    layer5_outputs(6094) <= not(layer4_outputs(5104)) or (layer4_outputs(5286));
    layer5_outputs(6095) <= not(layer4_outputs(4356));
    layer5_outputs(6096) <= not(layer4_outputs(6667)) or (layer4_outputs(2377));
    layer5_outputs(6097) <= not(layer4_outputs(1977));
    layer5_outputs(6098) <= not(layer4_outputs(2510));
    layer5_outputs(6099) <= (layer4_outputs(4589)) or (layer4_outputs(2767));
    layer5_outputs(6100) <= (layer4_outputs(97)) and not (layer4_outputs(1225));
    layer5_outputs(6101) <= not((layer4_outputs(163)) xor (layer4_outputs(622)));
    layer5_outputs(6102) <= layer4_outputs(3484);
    layer5_outputs(6103) <= layer4_outputs(7031);
    layer5_outputs(6104) <= not((layer4_outputs(1623)) or (layer4_outputs(1679)));
    layer5_outputs(6105) <= (layer4_outputs(4047)) and not (layer4_outputs(3262));
    layer5_outputs(6106) <= (layer4_outputs(5299)) or (layer4_outputs(5340));
    layer5_outputs(6107) <= not((layer4_outputs(3647)) or (layer4_outputs(413)));
    layer5_outputs(6108) <= layer4_outputs(4236);
    layer5_outputs(6109) <= '0';
    layer5_outputs(6110) <= not((layer4_outputs(726)) xor (layer4_outputs(1635)));
    layer5_outputs(6111) <= (layer4_outputs(5177)) xor (layer4_outputs(293));
    layer5_outputs(6112) <= layer4_outputs(3299);
    layer5_outputs(6113) <= (layer4_outputs(6889)) and (layer4_outputs(4347));
    layer5_outputs(6114) <= layer4_outputs(335);
    layer5_outputs(6115) <= not((layer4_outputs(1743)) and (layer4_outputs(7331)));
    layer5_outputs(6116) <= (layer4_outputs(2672)) xor (layer4_outputs(1282));
    layer5_outputs(6117) <= layer4_outputs(3580);
    layer5_outputs(6118) <= layer4_outputs(1842);
    layer5_outputs(6119) <= not(layer4_outputs(2716));
    layer5_outputs(6120) <= (layer4_outputs(770)) and (layer4_outputs(6271));
    layer5_outputs(6121) <= layer4_outputs(7589);
    layer5_outputs(6122) <= (layer4_outputs(2737)) or (layer4_outputs(5902));
    layer5_outputs(6123) <= (layer4_outputs(256)) and (layer4_outputs(1784));
    layer5_outputs(6124) <= layer4_outputs(7322);
    layer5_outputs(6125) <= not(layer4_outputs(4581)) or (layer4_outputs(3860));
    layer5_outputs(6126) <= layer4_outputs(415);
    layer5_outputs(6127) <= not(layer4_outputs(4018));
    layer5_outputs(6128) <= (layer4_outputs(1647)) and not (layer4_outputs(6951));
    layer5_outputs(6129) <= (layer4_outputs(4520)) and not (layer4_outputs(6229));
    layer5_outputs(6130) <= not(layer4_outputs(5603));
    layer5_outputs(6131) <= not(layer4_outputs(6242));
    layer5_outputs(6132) <= not((layer4_outputs(1250)) xor (layer4_outputs(2961)));
    layer5_outputs(6133) <= (layer4_outputs(4639)) and not (layer4_outputs(6386));
    layer5_outputs(6134) <= not((layer4_outputs(1712)) or (layer4_outputs(1154)));
    layer5_outputs(6135) <= not((layer4_outputs(1925)) xor (layer4_outputs(3423)));
    layer5_outputs(6136) <= layer4_outputs(3146);
    layer5_outputs(6137) <= not(layer4_outputs(2179)) or (layer4_outputs(480));
    layer5_outputs(6138) <= '0';
    layer5_outputs(6139) <= layer4_outputs(5232);
    layer5_outputs(6140) <= layer4_outputs(6369);
    layer5_outputs(6141) <= not((layer4_outputs(3587)) xor (layer4_outputs(5972)));
    layer5_outputs(6142) <= (layer4_outputs(2348)) xor (layer4_outputs(2490));
    layer5_outputs(6143) <= layer4_outputs(759);
    layer5_outputs(6144) <= not((layer4_outputs(6518)) and (layer4_outputs(4864)));
    layer5_outputs(6145) <= layer4_outputs(7659);
    layer5_outputs(6146) <= '0';
    layer5_outputs(6147) <= (layer4_outputs(3235)) and not (layer4_outputs(1031));
    layer5_outputs(6148) <= (layer4_outputs(7152)) and not (layer4_outputs(6846));
    layer5_outputs(6149) <= layer4_outputs(230);
    layer5_outputs(6150) <= not((layer4_outputs(4301)) xor (layer4_outputs(2277)));
    layer5_outputs(6151) <= layer4_outputs(7327);
    layer5_outputs(6152) <= not(layer4_outputs(734));
    layer5_outputs(6153) <= (layer4_outputs(2075)) xor (layer4_outputs(4782));
    layer5_outputs(6154) <= not(layer4_outputs(4768));
    layer5_outputs(6155) <= not(layer4_outputs(3669));
    layer5_outputs(6156) <= not(layer4_outputs(3424));
    layer5_outputs(6157) <= (layer4_outputs(4196)) and (layer4_outputs(4363));
    layer5_outputs(6158) <= not((layer4_outputs(1151)) and (layer4_outputs(2757)));
    layer5_outputs(6159) <= (layer4_outputs(6181)) or (layer4_outputs(4858));
    layer5_outputs(6160) <= not(layer4_outputs(1786));
    layer5_outputs(6161) <= '0';
    layer5_outputs(6162) <= '0';
    layer5_outputs(6163) <= (layer4_outputs(5122)) xor (layer4_outputs(2374));
    layer5_outputs(6164) <= (layer4_outputs(1206)) xor (layer4_outputs(5133));
    layer5_outputs(6165) <= layer4_outputs(6088);
    layer5_outputs(6166) <= (layer4_outputs(2765)) and not (layer4_outputs(6042));
    layer5_outputs(6167) <= (layer4_outputs(3376)) and not (layer4_outputs(1050));
    layer5_outputs(6168) <= (layer4_outputs(5429)) or (layer4_outputs(6161));
    layer5_outputs(6169) <= not((layer4_outputs(6487)) xor (layer4_outputs(5259)));
    layer5_outputs(6170) <= not(layer4_outputs(5055));
    layer5_outputs(6171) <= layer4_outputs(3859);
    layer5_outputs(6172) <= layer4_outputs(7002);
    layer5_outputs(6173) <= (layer4_outputs(1851)) and (layer4_outputs(2363));
    layer5_outputs(6174) <= not((layer4_outputs(7519)) xor (layer4_outputs(2969)));
    layer5_outputs(6175) <= (layer4_outputs(6778)) and (layer4_outputs(3123));
    layer5_outputs(6176) <= not(layer4_outputs(3580));
    layer5_outputs(6177) <= layer4_outputs(4976);
    layer5_outputs(6178) <= (layer4_outputs(2763)) and not (layer4_outputs(1070));
    layer5_outputs(6179) <= not((layer4_outputs(7560)) xor (layer4_outputs(3765)));
    layer5_outputs(6180) <= (layer4_outputs(831)) and (layer4_outputs(6866));
    layer5_outputs(6181) <= not(layer4_outputs(1605));
    layer5_outputs(6182) <= (layer4_outputs(7292)) or (layer4_outputs(5505));
    layer5_outputs(6183) <= not(layer4_outputs(4729));
    layer5_outputs(6184) <= '0';
    layer5_outputs(6185) <= layer4_outputs(3358);
    layer5_outputs(6186) <= (layer4_outputs(277)) and not (layer4_outputs(6312));
    layer5_outputs(6187) <= layer4_outputs(5073);
    layer5_outputs(6188) <= (layer4_outputs(552)) and not (layer4_outputs(5270));
    layer5_outputs(6189) <= (layer4_outputs(855)) or (layer4_outputs(128));
    layer5_outputs(6190) <= not(layer4_outputs(141));
    layer5_outputs(6191) <= not((layer4_outputs(4766)) and (layer4_outputs(6240)));
    layer5_outputs(6192) <= not(layer4_outputs(1188)) or (layer4_outputs(7402));
    layer5_outputs(6193) <= not((layer4_outputs(3571)) xor (layer4_outputs(506)));
    layer5_outputs(6194) <= layer4_outputs(853);
    layer5_outputs(6195) <= not((layer4_outputs(4437)) xor (layer4_outputs(3210)));
    layer5_outputs(6196) <= not((layer4_outputs(1091)) or (layer4_outputs(7239)));
    layer5_outputs(6197) <= (layer4_outputs(3018)) and not (layer4_outputs(7520));
    layer5_outputs(6198) <= (layer4_outputs(953)) or (layer4_outputs(5990));
    layer5_outputs(6199) <= not(layer4_outputs(1292));
    layer5_outputs(6200) <= not((layer4_outputs(922)) and (layer4_outputs(1517)));
    layer5_outputs(6201) <= (layer4_outputs(5113)) xor (layer4_outputs(4088));
    layer5_outputs(6202) <= not(layer4_outputs(3378));
    layer5_outputs(6203) <= layer4_outputs(4354);
    layer5_outputs(6204) <= layer4_outputs(2409);
    layer5_outputs(6205) <= not(layer4_outputs(808));
    layer5_outputs(6206) <= not(layer4_outputs(2594));
    layer5_outputs(6207) <= layer4_outputs(3972);
    layer5_outputs(6208) <= layer4_outputs(3316);
    layer5_outputs(6209) <= layer4_outputs(6709);
    layer5_outputs(6210) <= layer4_outputs(4586);
    layer5_outputs(6211) <= layer4_outputs(181);
    layer5_outputs(6212) <= (layer4_outputs(5552)) and not (layer4_outputs(3486));
    layer5_outputs(6213) <= (layer4_outputs(910)) or (layer4_outputs(4811));
    layer5_outputs(6214) <= not(layer4_outputs(7538)) or (layer4_outputs(4362));
    layer5_outputs(6215) <= layer4_outputs(6256);
    layer5_outputs(6216) <= (layer4_outputs(4426)) xor (layer4_outputs(3775));
    layer5_outputs(6217) <= not(layer4_outputs(2306));
    layer5_outputs(6218) <= (layer4_outputs(5950)) and (layer4_outputs(2677));
    layer5_outputs(6219) <= not((layer4_outputs(5049)) or (layer4_outputs(980)));
    layer5_outputs(6220) <= layer4_outputs(6637);
    layer5_outputs(6221) <= (layer4_outputs(1346)) and (layer4_outputs(6815));
    layer5_outputs(6222) <= not(layer4_outputs(7313));
    layer5_outputs(6223) <= not(layer4_outputs(3379));
    layer5_outputs(6224) <= layer4_outputs(610);
    layer5_outputs(6225) <= not(layer4_outputs(1875));
    layer5_outputs(6226) <= layer4_outputs(1445);
    layer5_outputs(6227) <= not((layer4_outputs(346)) or (layer4_outputs(3634)));
    layer5_outputs(6228) <= not(layer4_outputs(1609)) or (layer4_outputs(4432));
    layer5_outputs(6229) <= not(layer4_outputs(2513));
    layer5_outputs(6230) <= not((layer4_outputs(1917)) or (layer4_outputs(126)));
    layer5_outputs(6231) <= (layer4_outputs(5983)) or (layer4_outputs(3044));
    layer5_outputs(6232) <= not((layer4_outputs(2287)) xor (layer4_outputs(4612)));
    layer5_outputs(6233) <= layer4_outputs(7466);
    layer5_outputs(6234) <= (layer4_outputs(4607)) and not (layer4_outputs(5258));
    layer5_outputs(6235) <= layer4_outputs(803);
    layer5_outputs(6236) <= (layer4_outputs(901)) xor (layer4_outputs(1909));
    layer5_outputs(6237) <= layer4_outputs(3987);
    layer5_outputs(6238) <= (layer4_outputs(2652)) and not (layer4_outputs(996));
    layer5_outputs(6239) <= not((layer4_outputs(2316)) xor (layer4_outputs(3365)));
    layer5_outputs(6240) <= (layer4_outputs(2762)) xor (layer4_outputs(5832));
    layer5_outputs(6241) <= (layer4_outputs(7168)) xor (layer4_outputs(6338));
    layer5_outputs(6242) <= layer4_outputs(4413);
    layer5_outputs(6243) <= not(layer4_outputs(5427));
    layer5_outputs(6244) <= (layer4_outputs(4873)) or (layer4_outputs(5690));
    layer5_outputs(6245) <= layer4_outputs(6850);
    layer5_outputs(6246) <= (layer4_outputs(4358)) and not (layer4_outputs(5288));
    layer5_outputs(6247) <= not(layer4_outputs(7281));
    layer5_outputs(6248) <= not(layer4_outputs(544));
    layer5_outputs(6249) <= not(layer4_outputs(1389));
    layer5_outputs(6250) <= (layer4_outputs(7044)) xor (layer4_outputs(5762));
    layer5_outputs(6251) <= (layer4_outputs(6292)) and not (layer4_outputs(444));
    layer5_outputs(6252) <= layer4_outputs(284);
    layer5_outputs(6253) <= not((layer4_outputs(4732)) xor (layer4_outputs(492)));
    layer5_outputs(6254) <= (layer4_outputs(790)) and not (layer4_outputs(1787));
    layer5_outputs(6255) <= layer4_outputs(6285);
    layer5_outputs(6256) <= (layer4_outputs(5310)) and not (layer4_outputs(6434));
    layer5_outputs(6257) <= layer4_outputs(69);
    layer5_outputs(6258) <= not(layer4_outputs(7356)) or (layer4_outputs(5180));
    layer5_outputs(6259) <= not(layer4_outputs(223));
    layer5_outputs(6260) <= (layer4_outputs(5679)) xor (layer4_outputs(6325));
    layer5_outputs(6261) <= layer4_outputs(6532);
    layer5_outputs(6262) <= (layer4_outputs(6817)) and not (layer4_outputs(7000));
    layer5_outputs(6263) <= not(layer4_outputs(7475));
    layer5_outputs(6264) <= not((layer4_outputs(6844)) and (layer4_outputs(1588)));
    layer5_outputs(6265) <= not(layer4_outputs(7676));
    layer5_outputs(6266) <= not(layer4_outputs(3700));
    layer5_outputs(6267) <= (layer4_outputs(91)) and not (layer4_outputs(2827));
    layer5_outputs(6268) <= not((layer4_outputs(1712)) or (layer4_outputs(1922)));
    layer5_outputs(6269) <= (layer4_outputs(5804)) and not (layer4_outputs(5100));
    layer5_outputs(6270) <= not((layer4_outputs(6838)) xor (layer4_outputs(4843)));
    layer5_outputs(6271) <= not(layer4_outputs(2383));
    layer5_outputs(6272) <= not(layer4_outputs(1476));
    layer5_outputs(6273) <= not((layer4_outputs(5870)) xor (layer4_outputs(7282)));
    layer5_outputs(6274) <= (layer4_outputs(4999)) or (layer4_outputs(3769));
    layer5_outputs(6275) <= layer4_outputs(2023);
    layer5_outputs(6276) <= not(layer4_outputs(2201)) or (layer4_outputs(4280));
    layer5_outputs(6277) <= not(layer4_outputs(1013));
    layer5_outputs(6278) <= not((layer4_outputs(3400)) and (layer4_outputs(3344)));
    layer5_outputs(6279) <= layer4_outputs(920);
    layer5_outputs(6280) <= not(layer4_outputs(7512)) or (layer4_outputs(322));
    layer5_outputs(6281) <= layer4_outputs(2889);
    layer5_outputs(6282) <= layer4_outputs(1253);
    layer5_outputs(6283) <= (layer4_outputs(1497)) or (layer4_outputs(3392));
    layer5_outputs(6284) <= not((layer4_outputs(1202)) and (layer4_outputs(1316)));
    layer5_outputs(6285) <= layer4_outputs(370);
    layer5_outputs(6286) <= (layer4_outputs(882)) xor (layer4_outputs(7660));
    layer5_outputs(6287) <= (layer4_outputs(2520)) and not (layer4_outputs(1412));
    layer5_outputs(6288) <= (layer4_outputs(5386)) xor (layer4_outputs(4120));
    layer5_outputs(6289) <= not((layer4_outputs(288)) xor (layer4_outputs(3477)));
    layer5_outputs(6290) <= not((layer4_outputs(4323)) or (layer4_outputs(3785)));
    layer5_outputs(6291) <= (layer4_outputs(1632)) and not (layer4_outputs(3504));
    layer5_outputs(6292) <= '1';
    layer5_outputs(6293) <= (layer4_outputs(195)) and not (layer4_outputs(5171));
    layer5_outputs(6294) <= not((layer4_outputs(6937)) or (layer4_outputs(6686)));
    layer5_outputs(6295) <= (layer4_outputs(7252)) and not (layer4_outputs(5263));
    layer5_outputs(6296) <= not(layer4_outputs(6433));
    layer5_outputs(6297) <= not(layer4_outputs(1369));
    layer5_outputs(6298) <= (layer4_outputs(2593)) and not (layer4_outputs(3854));
    layer5_outputs(6299) <= not((layer4_outputs(1436)) or (layer4_outputs(2414)));
    layer5_outputs(6300) <= not(layer4_outputs(2022));
    layer5_outputs(6301) <= (layer4_outputs(1808)) xor (layer4_outputs(4193));
    layer5_outputs(6302) <= not(layer4_outputs(6488)) or (layer4_outputs(6874));
    layer5_outputs(6303) <= not(layer4_outputs(1514));
    layer5_outputs(6304) <= not(layer4_outputs(7157)) or (layer4_outputs(1216));
    layer5_outputs(6305) <= not(layer4_outputs(2718));
    layer5_outputs(6306) <= layer4_outputs(2898);
    layer5_outputs(6307) <= not(layer4_outputs(3211));
    layer5_outputs(6308) <= (layer4_outputs(2474)) or (layer4_outputs(2495));
    layer5_outputs(6309) <= not((layer4_outputs(2211)) or (layer4_outputs(5611)));
    layer5_outputs(6310) <= layer4_outputs(5727);
    layer5_outputs(6311) <= layer4_outputs(5219);
    layer5_outputs(6312) <= not(layer4_outputs(1240));
    layer5_outputs(6313) <= not(layer4_outputs(7308));
    layer5_outputs(6314) <= (layer4_outputs(3664)) and not (layer4_outputs(4323));
    layer5_outputs(6315) <= layer4_outputs(5103);
    layer5_outputs(6316) <= (layer4_outputs(2350)) and (layer4_outputs(994));
    layer5_outputs(6317) <= layer4_outputs(6753);
    layer5_outputs(6318) <= not(layer4_outputs(5121));
    layer5_outputs(6319) <= (layer4_outputs(6481)) and not (layer4_outputs(3158));
    layer5_outputs(6320) <= not((layer4_outputs(1320)) xor (layer4_outputs(1174)));
    layer5_outputs(6321) <= layer4_outputs(222);
    layer5_outputs(6322) <= (layer4_outputs(6500)) xor (layer4_outputs(1841));
    layer5_outputs(6323) <= not((layer4_outputs(6446)) xor (layer4_outputs(1570)));
    layer5_outputs(6324) <= not(layer4_outputs(1806));
    layer5_outputs(6325) <= not((layer4_outputs(4317)) and (layer4_outputs(68)));
    layer5_outputs(6326) <= not((layer4_outputs(6939)) or (layer4_outputs(2992)));
    layer5_outputs(6327) <= not((layer4_outputs(7650)) or (layer4_outputs(5870)));
    layer5_outputs(6328) <= not(layer4_outputs(4391));
    layer5_outputs(6329) <= not(layer4_outputs(4899));
    layer5_outputs(6330) <= not(layer4_outputs(4403));
    layer5_outputs(6331) <= not(layer4_outputs(6077));
    layer5_outputs(6332) <= (layer4_outputs(4774)) and not (layer4_outputs(1607));
    layer5_outputs(6333) <= (layer4_outputs(3697)) or (layer4_outputs(2360));
    layer5_outputs(6334) <= layer4_outputs(7354);
    layer5_outputs(6335) <= not((layer4_outputs(50)) or (layer4_outputs(1807)));
    layer5_outputs(6336) <= '0';
    layer5_outputs(6337) <= (layer4_outputs(3058)) and not (layer4_outputs(6264));
    layer5_outputs(6338) <= (layer4_outputs(3525)) and (layer4_outputs(7636));
    layer5_outputs(6339) <= layer4_outputs(7054);
    layer5_outputs(6340) <= not(layer4_outputs(551));
    layer5_outputs(6341) <= (layer4_outputs(1645)) and (layer4_outputs(3120));
    layer5_outputs(6342) <= layer4_outputs(7299);
    layer5_outputs(6343) <= not(layer4_outputs(3324));
    layer5_outputs(6344) <= not(layer4_outputs(5584));
    layer5_outputs(6345) <= layer4_outputs(1048);
    layer5_outputs(6346) <= not((layer4_outputs(4106)) xor (layer4_outputs(996)));
    layer5_outputs(6347) <= layer4_outputs(3953);
    layer5_outputs(6348) <= not(layer4_outputs(4382));
    layer5_outputs(6349) <= not((layer4_outputs(5759)) and (layer4_outputs(2388)));
    layer5_outputs(6350) <= not(layer4_outputs(3031));
    layer5_outputs(6351) <= layer4_outputs(828);
    layer5_outputs(6352) <= (layer4_outputs(1091)) xor (layer4_outputs(423));
    layer5_outputs(6353) <= not(layer4_outputs(7372));
    layer5_outputs(6354) <= not((layer4_outputs(3400)) xor (layer4_outputs(2952)));
    layer5_outputs(6355) <= not(layer4_outputs(1685));
    layer5_outputs(6356) <= not(layer4_outputs(4163));
    layer5_outputs(6357) <= not(layer4_outputs(1592));
    layer5_outputs(6358) <= not(layer4_outputs(1371));
    layer5_outputs(6359) <= layer4_outputs(5822);
    layer5_outputs(6360) <= not(layer4_outputs(6048));
    layer5_outputs(6361) <= (layer4_outputs(3414)) xor (layer4_outputs(5280));
    layer5_outputs(6362) <= (layer4_outputs(535)) and not (layer4_outputs(7096));
    layer5_outputs(6363) <= not((layer4_outputs(5840)) xor (layer4_outputs(2855)));
    layer5_outputs(6364) <= (layer4_outputs(2047)) xor (layer4_outputs(1686));
    layer5_outputs(6365) <= not(layer4_outputs(3602)) or (layer4_outputs(5002));
    layer5_outputs(6366) <= layer4_outputs(3904);
    layer5_outputs(6367) <= not(layer4_outputs(5458)) or (layer4_outputs(101));
    layer5_outputs(6368) <= layer4_outputs(270);
    layer5_outputs(6369) <= layer4_outputs(5886);
    layer5_outputs(6370) <= not(layer4_outputs(4549));
    layer5_outputs(6371) <= not(layer4_outputs(4137));
    layer5_outputs(6372) <= not((layer4_outputs(5350)) and (layer4_outputs(1319)));
    layer5_outputs(6373) <= (layer4_outputs(3564)) and not (layer4_outputs(1224));
    layer5_outputs(6374) <= not(layer4_outputs(1262));
    layer5_outputs(6375) <= layer4_outputs(5179);
    layer5_outputs(6376) <= not((layer4_outputs(7573)) or (layer4_outputs(3085)));
    layer5_outputs(6377) <= not(layer4_outputs(293)) or (layer4_outputs(4935));
    layer5_outputs(6378) <= (layer4_outputs(5961)) or (layer4_outputs(9));
    layer5_outputs(6379) <= (layer4_outputs(49)) and not (layer4_outputs(3057));
    layer5_outputs(6380) <= not((layer4_outputs(5905)) or (layer4_outputs(7650)));
    layer5_outputs(6381) <= not(layer4_outputs(2476)) or (layer4_outputs(6226));
    layer5_outputs(6382) <= not((layer4_outputs(5560)) xor (layer4_outputs(3733)));
    layer5_outputs(6383) <= not(layer4_outputs(7553)) or (layer4_outputs(6148));
    layer5_outputs(6384) <= layer4_outputs(1754);
    layer5_outputs(6385) <= (layer4_outputs(1879)) xor (layer4_outputs(7319));
    layer5_outputs(6386) <= layer4_outputs(5982);
    layer5_outputs(6387) <= (layer4_outputs(53)) and not (layer4_outputs(5612));
    layer5_outputs(6388) <= (layer4_outputs(1707)) and not (layer4_outputs(637));
    layer5_outputs(6389) <= not(layer4_outputs(4592));
    layer5_outputs(6390) <= not(layer4_outputs(7486));
    layer5_outputs(6391) <= (layer4_outputs(3521)) and (layer4_outputs(2710));
    layer5_outputs(6392) <= not(layer4_outputs(1745));
    layer5_outputs(6393) <= (layer4_outputs(5976)) or (layer4_outputs(6598));
    layer5_outputs(6394) <= not(layer4_outputs(5072));
    layer5_outputs(6395) <= layer4_outputs(5807);
    layer5_outputs(6396) <= not((layer4_outputs(1047)) xor (layer4_outputs(3380)));
    layer5_outputs(6397) <= not(layer4_outputs(1333));
    layer5_outputs(6398) <= (layer4_outputs(1763)) xor (layer4_outputs(1727));
    layer5_outputs(6399) <= layer4_outputs(4085);
    layer5_outputs(6400) <= (layer4_outputs(7071)) and not (layer4_outputs(1694));
    layer5_outputs(6401) <= (layer4_outputs(7276)) and not (layer4_outputs(6751));
    layer5_outputs(6402) <= (layer4_outputs(3493)) and not (layer4_outputs(5590));
    layer5_outputs(6403) <= layer4_outputs(5593);
    layer5_outputs(6404) <= layer4_outputs(5658);
    layer5_outputs(6405) <= layer4_outputs(4079);
    layer5_outputs(6406) <= layer4_outputs(1471);
    layer5_outputs(6407) <= '1';
    layer5_outputs(6408) <= not(layer4_outputs(7118)) or (layer4_outputs(3381));
    layer5_outputs(6409) <= (layer4_outputs(1797)) or (layer4_outputs(650));
    layer5_outputs(6410) <= layer4_outputs(5785);
    layer5_outputs(6411) <= layer4_outputs(4963);
    layer5_outputs(6412) <= '0';
    layer5_outputs(6413) <= (layer4_outputs(5234)) and not (layer4_outputs(3608));
    layer5_outputs(6414) <= not((layer4_outputs(3831)) and (layer4_outputs(2111)));
    layer5_outputs(6415) <= not(layer4_outputs(4226));
    layer5_outputs(6416) <= layer4_outputs(1441);
    layer5_outputs(6417) <= (layer4_outputs(334)) or (layer4_outputs(2093));
    layer5_outputs(6418) <= not((layer4_outputs(4746)) and (layer4_outputs(1677)));
    layer5_outputs(6419) <= (layer4_outputs(6669)) or (layer4_outputs(108));
    layer5_outputs(6420) <= not(layer4_outputs(3264));
    layer5_outputs(6421) <= not((layer4_outputs(4076)) or (layer4_outputs(7293)));
    layer5_outputs(6422) <= not((layer4_outputs(2067)) or (layer4_outputs(1730)));
    layer5_outputs(6423) <= layer4_outputs(6127);
    layer5_outputs(6424) <= not(layer4_outputs(1153)) or (layer4_outputs(5442));
    layer5_outputs(6425) <= (layer4_outputs(4099)) or (layer4_outputs(1085));
    layer5_outputs(6426) <= not(layer4_outputs(826)) or (layer4_outputs(6356));
    layer5_outputs(6427) <= not(layer4_outputs(6016));
    layer5_outputs(6428) <= not(layer4_outputs(418));
    layer5_outputs(6429) <= not(layer4_outputs(4626));
    layer5_outputs(6430) <= (layer4_outputs(4141)) or (layer4_outputs(4898));
    layer5_outputs(6431) <= layer4_outputs(6034);
    layer5_outputs(6432) <= (layer4_outputs(6109)) and not (layer4_outputs(1913));
    layer5_outputs(6433) <= not(layer4_outputs(4366)) or (layer4_outputs(479));
    layer5_outputs(6434) <= not(layer4_outputs(3901));
    layer5_outputs(6435) <= layer4_outputs(1406);
    layer5_outputs(6436) <= not(layer4_outputs(5249));
    layer5_outputs(6437) <= layer4_outputs(975);
    layer5_outputs(6438) <= not(layer4_outputs(3632)) or (layer4_outputs(6978));
    layer5_outputs(6439) <= layer4_outputs(3041);
    layer5_outputs(6440) <= layer4_outputs(956);
    layer5_outputs(6441) <= not((layer4_outputs(2361)) xor (layer4_outputs(4185)));
    layer5_outputs(6442) <= (layer4_outputs(7510)) and not (layer4_outputs(5215));
    layer5_outputs(6443) <= not((layer4_outputs(1341)) or (layer4_outputs(4104)));
    layer5_outputs(6444) <= not(layer4_outputs(270)) or (layer4_outputs(2543));
    layer5_outputs(6445) <= layer4_outputs(183);
    layer5_outputs(6446) <= (layer4_outputs(1231)) and not (layer4_outputs(7515));
    layer5_outputs(6447) <= layer4_outputs(6091);
    layer5_outputs(6448) <= not(layer4_outputs(3969));
    layer5_outputs(6449) <= not(layer4_outputs(2272));
    layer5_outputs(6450) <= not((layer4_outputs(3412)) xor (layer4_outputs(138)));
    layer5_outputs(6451) <= (layer4_outputs(4337)) and not (layer4_outputs(7302));
    layer5_outputs(6452) <= not(layer4_outputs(5682));
    layer5_outputs(6453) <= not(layer4_outputs(74));
    layer5_outputs(6454) <= not(layer4_outputs(5513));
    layer5_outputs(6455) <= (layer4_outputs(1998)) and not (layer4_outputs(5838));
    layer5_outputs(6456) <= (layer4_outputs(4042)) xor (layer4_outputs(5690));
    layer5_outputs(6457) <= not(layer4_outputs(1738)) or (layer4_outputs(7651));
    layer5_outputs(6458) <= layer4_outputs(1708);
    layer5_outputs(6459) <= (layer4_outputs(1012)) and not (layer4_outputs(3914));
    layer5_outputs(6460) <= not((layer4_outputs(5595)) xor (layer4_outputs(84)));
    layer5_outputs(6461) <= (layer4_outputs(1386)) and not (layer4_outputs(6313));
    layer5_outputs(6462) <= (layer4_outputs(4010)) and not (layer4_outputs(4774));
    layer5_outputs(6463) <= not((layer4_outputs(1637)) xor (layer4_outputs(5149)));
    layer5_outputs(6464) <= not(layer4_outputs(5627));
    layer5_outputs(6465) <= not(layer4_outputs(350));
    layer5_outputs(6466) <= not(layer4_outputs(3374)) or (layer4_outputs(7117));
    layer5_outputs(6467) <= not(layer4_outputs(2473));
    layer5_outputs(6468) <= layer4_outputs(375);
    layer5_outputs(6469) <= not(layer4_outputs(4184));
    layer5_outputs(6470) <= not((layer4_outputs(2512)) and (layer4_outputs(6308)));
    layer5_outputs(6471) <= not((layer4_outputs(1034)) or (layer4_outputs(6097)));
    layer5_outputs(6472) <= not(layer4_outputs(805));
    layer5_outputs(6473) <= (layer4_outputs(2741)) and not (layer4_outputs(1134));
    layer5_outputs(6474) <= not((layer4_outputs(2969)) or (layer4_outputs(7487)));
    layer5_outputs(6475) <= (layer4_outputs(1588)) or (layer4_outputs(7292));
    layer5_outputs(6476) <= (layer4_outputs(5174)) and not (layer4_outputs(7241));
    layer5_outputs(6477) <= (layer4_outputs(2994)) or (layer4_outputs(4910));
    layer5_outputs(6478) <= (layer4_outputs(4061)) and (layer4_outputs(349));
    layer5_outputs(6479) <= layer4_outputs(84);
    layer5_outputs(6480) <= (layer4_outputs(6012)) xor (layer4_outputs(5224));
    layer5_outputs(6481) <= not(layer4_outputs(3189));
    layer5_outputs(6482) <= not(layer4_outputs(6215));
    layer5_outputs(6483) <= (layer4_outputs(4334)) and not (layer4_outputs(6781));
    layer5_outputs(6484) <= not(layer4_outputs(7152));
    layer5_outputs(6485) <= (layer4_outputs(2228)) and not (layer4_outputs(3805));
    layer5_outputs(6486) <= not((layer4_outputs(5794)) and (layer4_outputs(2218)));
    layer5_outputs(6487) <= not(layer4_outputs(495));
    layer5_outputs(6488) <= (layer4_outputs(4039)) and not (layer4_outputs(234));
    layer5_outputs(6489) <= not(layer4_outputs(5888));
    layer5_outputs(6490) <= not(layer4_outputs(6537));
    layer5_outputs(6491) <= not(layer4_outputs(1083)) or (layer4_outputs(6235));
    layer5_outputs(6492) <= not(layer4_outputs(3327));
    layer5_outputs(6493) <= not((layer4_outputs(4676)) xor (layer4_outputs(4345)));
    layer5_outputs(6494) <= not(layer4_outputs(543));
    layer5_outputs(6495) <= layer4_outputs(4267);
    layer5_outputs(6496) <= not(layer4_outputs(6499));
    layer5_outputs(6497) <= not(layer4_outputs(3663)) or (layer4_outputs(5641));
    layer5_outputs(6498) <= not(layer4_outputs(7071));
    layer5_outputs(6499) <= not(layer4_outputs(5849));
    layer5_outputs(6500) <= layer4_outputs(6242);
    layer5_outputs(6501) <= layer4_outputs(7246);
    layer5_outputs(6502) <= layer4_outputs(2068);
    layer5_outputs(6503) <= not(layer4_outputs(1237));
    layer5_outputs(6504) <= not(layer4_outputs(2274));
    layer5_outputs(6505) <= not(layer4_outputs(4856)) or (layer4_outputs(1571));
    layer5_outputs(6506) <= not(layer4_outputs(4286)) or (layer4_outputs(4432));
    layer5_outputs(6507) <= layer4_outputs(4203);
    layer5_outputs(6508) <= layer4_outputs(4922);
    layer5_outputs(6509) <= not(layer4_outputs(905));
    layer5_outputs(6510) <= layer4_outputs(4909);
    layer5_outputs(6511) <= layer4_outputs(2845);
    layer5_outputs(6512) <= not(layer4_outputs(5109));
    layer5_outputs(6513) <= (layer4_outputs(2735)) and (layer4_outputs(2897));
    layer5_outputs(6514) <= not((layer4_outputs(5622)) or (layer4_outputs(2415)));
    layer5_outputs(6515) <= layer4_outputs(7386);
    layer5_outputs(6516) <= '0';
    layer5_outputs(6517) <= not(layer4_outputs(6217)) or (layer4_outputs(3828));
    layer5_outputs(6518) <= layer4_outputs(3205);
    layer5_outputs(6519) <= not(layer4_outputs(7060));
    layer5_outputs(6520) <= (layer4_outputs(313)) and not (layer4_outputs(841));
    layer5_outputs(6521) <= not(layer4_outputs(3576)) or (layer4_outputs(3223));
    layer5_outputs(6522) <= (layer4_outputs(764)) and not (layer4_outputs(4680));
    layer5_outputs(6523) <= not(layer4_outputs(790));
    layer5_outputs(6524) <= layer4_outputs(6020);
    layer5_outputs(6525) <= (layer4_outputs(4309)) and not (layer4_outputs(6375));
    layer5_outputs(6526) <= layer4_outputs(4860);
    layer5_outputs(6527) <= (layer4_outputs(934)) or (layer4_outputs(5497));
    layer5_outputs(6528) <= not(layer4_outputs(5833)) or (layer4_outputs(5659));
    layer5_outputs(6529) <= layer4_outputs(4138);
    layer5_outputs(6530) <= not(layer4_outputs(7667));
    layer5_outputs(6531) <= layer4_outputs(1782);
    layer5_outputs(6532) <= not(layer4_outputs(5375));
    layer5_outputs(6533) <= layer4_outputs(6371);
    layer5_outputs(6534) <= not(layer4_outputs(2142));
    layer5_outputs(6535) <= not(layer4_outputs(7011)) or (layer4_outputs(1688));
    layer5_outputs(6536) <= (layer4_outputs(2768)) xor (layer4_outputs(4259));
    layer5_outputs(6537) <= (layer4_outputs(2413)) and not (layer4_outputs(6965));
    layer5_outputs(6538) <= not(layer4_outputs(2610));
    layer5_outputs(6539) <= (layer4_outputs(6359)) xor (layer4_outputs(5450));
    layer5_outputs(6540) <= not(layer4_outputs(3656));
    layer5_outputs(6541) <= (layer4_outputs(4216)) and not (layer4_outputs(6576));
    layer5_outputs(6542) <= (layer4_outputs(2189)) and (layer4_outputs(4996));
    layer5_outputs(6543) <= not(layer4_outputs(7495));
    layer5_outputs(6544) <= '0';
    layer5_outputs(6545) <= not(layer4_outputs(4203));
    layer5_outputs(6546) <= not(layer4_outputs(5822));
    layer5_outputs(6547) <= not(layer4_outputs(6055)) or (layer4_outputs(6198));
    layer5_outputs(6548) <= layer4_outputs(5368);
    layer5_outputs(6549) <= not((layer4_outputs(1407)) or (layer4_outputs(5671)));
    layer5_outputs(6550) <= not(layer4_outputs(1009));
    layer5_outputs(6551) <= not(layer4_outputs(7337));
    layer5_outputs(6552) <= (layer4_outputs(523)) or (layer4_outputs(5954));
    layer5_outputs(6553) <= not((layer4_outputs(411)) xor (layer4_outputs(4866)));
    layer5_outputs(6554) <= not(layer4_outputs(7006));
    layer5_outputs(6555) <= (layer4_outputs(4635)) and (layer4_outputs(3373));
    layer5_outputs(6556) <= (layer4_outputs(3300)) and (layer4_outputs(4339));
    layer5_outputs(6557) <= not(layer4_outputs(5879));
    layer5_outputs(6558) <= (layer4_outputs(1410)) and not (layer4_outputs(5745));
    layer5_outputs(6559) <= not(layer4_outputs(6987));
    layer5_outputs(6560) <= not(layer4_outputs(4318)) or (layer4_outputs(1279));
    layer5_outputs(6561) <= (layer4_outputs(3708)) or (layer4_outputs(5608));
    layer5_outputs(6562) <= not(layer4_outputs(6483));
    layer5_outputs(6563) <= not(layer4_outputs(5704));
    layer5_outputs(6564) <= not(layer4_outputs(1801)) or (layer4_outputs(4069));
    layer5_outputs(6565) <= not(layer4_outputs(3114));
    layer5_outputs(6566) <= layer4_outputs(1017);
    layer5_outputs(6567) <= layer4_outputs(6259);
    layer5_outputs(6568) <= not((layer4_outputs(1034)) xor (layer4_outputs(1011)));
    layer5_outputs(6569) <= layer4_outputs(7624);
    layer5_outputs(6570) <= layer4_outputs(4590);
    layer5_outputs(6571) <= (layer4_outputs(3651)) and (layer4_outputs(6679));
    layer5_outputs(6572) <= not(layer4_outputs(7505));
    layer5_outputs(6573) <= not(layer4_outputs(2446)) or (layer4_outputs(2158));
    layer5_outputs(6574) <= not(layer4_outputs(7600));
    layer5_outputs(6575) <= not(layer4_outputs(24));
    layer5_outputs(6576) <= (layer4_outputs(3090)) xor (layer4_outputs(7283));
    layer5_outputs(6577) <= layer4_outputs(1787);
    layer5_outputs(6578) <= not(layer4_outputs(6252));
    layer5_outputs(6579) <= not(layer4_outputs(7514));
    layer5_outputs(6580) <= (layer4_outputs(5973)) and not (layer4_outputs(7506));
    layer5_outputs(6581) <= not(layer4_outputs(4296));
    layer5_outputs(6582) <= layer4_outputs(7502);
    layer5_outputs(6583) <= not((layer4_outputs(856)) or (layer4_outputs(7344)));
    layer5_outputs(6584) <= (layer4_outputs(4472)) and not (layer4_outputs(7297));
    layer5_outputs(6585) <= layer4_outputs(1493);
    layer5_outputs(6586) <= not((layer4_outputs(6250)) and (layer4_outputs(5766)));
    layer5_outputs(6587) <= layer4_outputs(3903);
    layer5_outputs(6588) <= not(layer4_outputs(2721));
    layer5_outputs(6589) <= (layer4_outputs(37)) and (layer4_outputs(4597));
    layer5_outputs(6590) <= layer4_outputs(633);
    layer5_outputs(6591) <= layer4_outputs(2565);
    layer5_outputs(6592) <= not((layer4_outputs(4050)) or (layer4_outputs(1780)));
    layer5_outputs(6593) <= layer4_outputs(1905);
    layer5_outputs(6594) <= (layer4_outputs(2707)) xor (layer4_outputs(3451));
    layer5_outputs(6595) <= (layer4_outputs(7440)) and not (layer4_outputs(6319));
    layer5_outputs(6596) <= layer4_outputs(5046);
    layer5_outputs(6597) <= not(layer4_outputs(3643));
    layer5_outputs(6598) <= layer4_outputs(6412);
    layer5_outputs(6599) <= layer4_outputs(3688);
    layer5_outputs(6600) <= layer4_outputs(1126);
    layer5_outputs(6601) <= '1';
    layer5_outputs(6602) <= not((layer4_outputs(4253)) and (layer4_outputs(7344)));
    layer5_outputs(6603) <= '1';
    layer5_outputs(6604) <= (layer4_outputs(4656)) xor (layer4_outputs(183));
    layer5_outputs(6605) <= layer4_outputs(2770);
    layer5_outputs(6606) <= (layer4_outputs(6175)) or (layer4_outputs(6854));
    layer5_outputs(6607) <= (layer4_outputs(674)) or (layer4_outputs(1063));
    layer5_outputs(6608) <= not(layer4_outputs(4242)) or (layer4_outputs(5451));
    layer5_outputs(6609) <= (layer4_outputs(1696)) xor (layer4_outputs(3398));
    layer5_outputs(6610) <= not(layer4_outputs(4950));
    layer5_outputs(6611) <= not((layer4_outputs(840)) or (layer4_outputs(1320)));
    layer5_outputs(6612) <= (layer4_outputs(1235)) and (layer4_outputs(6254));
    layer5_outputs(6613) <= not(layer4_outputs(100));
    layer5_outputs(6614) <= not((layer4_outputs(530)) or (layer4_outputs(6629)));
    layer5_outputs(6615) <= not(layer4_outputs(1026)) or (layer4_outputs(5222));
    layer5_outputs(6616) <= not((layer4_outputs(7230)) or (layer4_outputs(3586)));
    layer5_outputs(6617) <= not(layer4_outputs(3852));
    layer5_outputs(6618) <= (layer4_outputs(1008)) and not (layer4_outputs(7456));
    layer5_outputs(6619) <= layer4_outputs(5687);
    layer5_outputs(6620) <= layer4_outputs(6553);
    layer5_outputs(6621) <= (layer4_outputs(4015)) or (layer4_outputs(4500));
    layer5_outputs(6622) <= not(layer4_outputs(3335));
    layer5_outputs(6623) <= layer4_outputs(2501);
    layer5_outputs(6624) <= not((layer4_outputs(7546)) or (layer4_outputs(597)));
    layer5_outputs(6625) <= not(layer4_outputs(4785));
    layer5_outputs(6626) <= (layer4_outputs(6387)) and not (layer4_outputs(126));
    layer5_outputs(6627) <= (layer4_outputs(4247)) and not (layer4_outputs(4633));
    layer5_outputs(6628) <= layer4_outputs(2997);
    layer5_outputs(6629) <= not((layer4_outputs(5791)) or (layer4_outputs(2164)));
    layer5_outputs(6630) <= layer4_outputs(925);
    layer5_outputs(6631) <= not(layer4_outputs(7455)) or (layer4_outputs(349));
    layer5_outputs(6632) <= not(layer4_outputs(1412));
    layer5_outputs(6633) <= layer4_outputs(7568);
    layer5_outputs(6634) <= not(layer4_outputs(3964)) or (layer4_outputs(5452));
    layer5_outputs(6635) <= layer4_outputs(2752);
    layer5_outputs(6636) <= not((layer4_outputs(1907)) and (layer4_outputs(4736)));
    layer5_outputs(6637) <= not(layer4_outputs(6318));
    layer5_outputs(6638) <= not(layer4_outputs(6364));
    layer5_outputs(6639) <= not((layer4_outputs(2900)) or (layer4_outputs(7113)));
    layer5_outputs(6640) <= not((layer4_outputs(7604)) or (layer4_outputs(2575)));
    layer5_outputs(6641) <= not((layer4_outputs(1968)) xor (layer4_outputs(1595)));
    layer5_outputs(6642) <= layer4_outputs(3671);
    layer5_outputs(6643) <= not(layer4_outputs(1140));
    layer5_outputs(6644) <= (layer4_outputs(7633)) xor (layer4_outputs(4827));
    layer5_outputs(6645) <= not(layer4_outputs(81));
    layer5_outputs(6646) <= not(layer4_outputs(5830)) or (layer4_outputs(2050));
    layer5_outputs(6647) <= (layer4_outputs(3240)) and (layer4_outputs(1557));
    layer5_outputs(6648) <= layer4_outputs(7304);
    layer5_outputs(6649) <= (layer4_outputs(5736)) and not (layer4_outputs(2898));
    layer5_outputs(6650) <= layer4_outputs(6395);
    layer5_outputs(6651) <= not(layer4_outputs(1803));
    layer5_outputs(6652) <= (layer4_outputs(2810)) xor (layer4_outputs(3882));
    layer5_outputs(6653) <= not((layer4_outputs(6713)) xor (layer4_outputs(2701)));
    layer5_outputs(6654) <= (layer4_outputs(3681)) and (layer4_outputs(7267));
    layer5_outputs(6655) <= not(layer4_outputs(3750));
    layer5_outputs(6656) <= layer4_outputs(7233);
    layer5_outputs(6657) <= layer4_outputs(863);
    layer5_outputs(6658) <= not((layer4_outputs(4044)) and (layer4_outputs(5930)));
    layer5_outputs(6659) <= not((layer4_outputs(1192)) or (layer4_outputs(4481)));
    layer5_outputs(6660) <= (layer4_outputs(3637)) xor (layer4_outputs(708));
    layer5_outputs(6661) <= not(layer4_outputs(6920));
    layer5_outputs(6662) <= layer4_outputs(4258);
    layer5_outputs(6663) <= not(layer4_outputs(1883));
    layer5_outputs(6664) <= not((layer4_outputs(2593)) xor (layer4_outputs(81)));
    layer5_outputs(6665) <= (layer4_outputs(3126)) xor (layer4_outputs(6910));
    layer5_outputs(6666) <= (layer4_outputs(4013)) or (layer4_outputs(7413));
    layer5_outputs(6667) <= layer4_outputs(4538);
    layer5_outputs(6668) <= not(layer4_outputs(1833));
    layer5_outputs(6669) <= not((layer4_outputs(6025)) and (layer4_outputs(4849)));
    layer5_outputs(6670) <= not(layer4_outputs(6892));
    layer5_outputs(6671) <= layer4_outputs(6936);
    layer5_outputs(6672) <= not((layer4_outputs(2678)) or (layer4_outputs(3260)));
    layer5_outputs(6673) <= (layer4_outputs(430)) xor (layer4_outputs(3293));
    layer5_outputs(6674) <= not(layer4_outputs(4876));
    layer5_outputs(6675) <= (layer4_outputs(891)) or (layer4_outputs(6936));
    layer5_outputs(6676) <= layer4_outputs(2181);
    layer5_outputs(6677) <= not(layer4_outputs(6137));
    layer5_outputs(6678) <= layer4_outputs(801);
    layer5_outputs(6679) <= layer4_outputs(526);
    layer5_outputs(6680) <= (layer4_outputs(1973)) and (layer4_outputs(1035));
    layer5_outputs(6681) <= layer4_outputs(4610);
    layer5_outputs(6682) <= (layer4_outputs(1420)) xor (layer4_outputs(3543));
    layer5_outputs(6683) <= not(layer4_outputs(5984));
    layer5_outputs(6684) <= layer4_outputs(3033);
    layer5_outputs(6685) <= (layer4_outputs(493)) xor (layer4_outputs(600));
    layer5_outputs(6686) <= not((layer4_outputs(5866)) xor (layer4_outputs(943)));
    layer5_outputs(6687) <= layer4_outputs(4544);
    layer5_outputs(6688) <= layer4_outputs(78);
    layer5_outputs(6689) <= layer4_outputs(7001);
    layer5_outputs(6690) <= not(layer4_outputs(525));
    layer5_outputs(6691) <= not(layer4_outputs(5220));
    layer5_outputs(6692) <= not(layer4_outputs(7347));
    layer5_outputs(6693) <= layer4_outputs(1985);
    layer5_outputs(6694) <= not((layer4_outputs(5184)) xor (layer4_outputs(5271)));
    layer5_outputs(6695) <= not(layer4_outputs(6516)) or (layer4_outputs(4778));
    layer5_outputs(6696) <= not(layer4_outputs(3087)) or (layer4_outputs(982));
    layer5_outputs(6697) <= (layer4_outputs(1845)) or (layer4_outputs(5804));
    layer5_outputs(6698) <= layer4_outputs(1806);
    layer5_outputs(6699) <= layer4_outputs(196);
    layer5_outputs(6700) <= (layer4_outputs(2616)) and (layer4_outputs(3515));
    layer5_outputs(6701) <= layer4_outputs(7457);
    layer5_outputs(6702) <= layer4_outputs(6492);
    layer5_outputs(6703) <= not(layer4_outputs(7477));
    layer5_outputs(6704) <= (layer4_outputs(6710)) and (layer4_outputs(4444));
    layer5_outputs(6705) <= not(layer4_outputs(7507));
    layer5_outputs(6706) <= not(layer4_outputs(2260));
    layer5_outputs(6707) <= not(layer4_outputs(1613));
    layer5_outputs(6708) <= not(layer4_outputs(2489));
    layer5_outputs(6709) <= layer4_outputs(6337);
    layer5_outputs(6710) <= (layer4_outputs(1551)) and not (layer4_outputs(4112));
    layer5_outputs(6711) <= not((layer4_outputs(4267)) xor (layer4_outputs(5097)));
    layer5_outputs(6712) <= not(layer4_outputs(3317));
    layer5_outputs(6713) <= layer4_outputs(6711);
    layer5_outputs(6714) <= (layer4_outputs(5088)) xor (layer4_outputs(5034));
    layer5_outputs(6715) <= layer4_outputs(1220);
    layer5_outputs(6716) <= not(layer4_outputs(6737));
    layer5_outputs(6717) <= not(layer4_outputs(7462));
    layer5_outputs(6718) <= layer4_outputs(4602);
    layer5_outputs(6719) <= layer4_outputs(6561);
    layer5_outputs(6720) <= not((layer4_outputs(5422)) or (layer4_outputs(2298)));
    layer5_outputs(6721) <= layer4_outputs(3767);
    layer5_outputs(6722) <= (layer4_outputs(7226)) and not (layer4_outputs(5056));
    layer5_outputs(6723) <= (layer4_outputs(3678)) or (layer4_outputs(6880));
    layer5_outputs(6724) <= layer4_outputs(6136);
    layer5_outputs(6725) <= (layer4_outputs(7075)) xor (layer4_outputs(881));
    layer5_outputs(6726) <= (layer4_outputs(2319)) xor (layer4_outputs(2447));
    layer5_outputs(6727) <= not((layer4_outputs(6914)) or (layer4_outputs(1044)));
    layer5_outputs(6728) <= not(layer4_outputs(2276));
    layer5_outputs(6729) <= (layer4_outputs(2788)) or (layer4_outputs(6941));
    layer5_outputs(6730) <= (layer4_outputs(3317)) and not (layer4_outputs(5398));
    layer5_outputs(6731) <= layer4_outputs(5731);
    layer5_outputs(6732) <= not(layer4_outputs(1779));
    layer5_outputs(6733) <= '0';
    layer5_outputs(6734) <= not((layer4_outputs(1191)) or (layer4_outputs(7179)));
    layer5_outputs(6735) <= not((layer4_outputs(537)) or (layer4_outputs(5387)));
    layer5_outputs(6736) <= (layer4_outputs(6260)) xor (layer4_outputs(6592));
    layer5_outputs(6737) <= (layer4_outputs(2102)) xor (layer4_outputs(952));
    layer5_outputs(6738) <= (layer4_outputs(1122)) and not (layer4_outputs(3817));
    layer5_outputs(6739) <= not(layer4_outputs(7193));
    layer5_outputs(6740) <= not(layer4_outputs(3307));
    layer5_outputs(6741) <= layer4_outputs(7659);
    layer5_outputs(6742) <= layer4_outputs(3504);
    layer5_outputs(6743) <= not(layer4_outputs(6205));
    layer5_outputs(6744) <= layer4_outputs(3816);
    layer5_outputs(6745) <= (layer4_outputs(6396)) and not (layer4_outputs(6691));
    layer5_outputs(6746) <= not(layer4_outputs(3714));
    layer5_outputs(6747) <= not((layer4_outputs(3625)) and (layer4_outputs(437)));
    layer5_outputs(6748) <= layer4_outputs(5722);
    layer5_outputs(6749) <= not(layer4_outputs(2556));
    layer5_outputs(6750) <= (layer4_outputs(7613)) and (layer4_outputs(609));
    layer5_outputs(6751) <= not((layer4_outputs(1616)) xor (layer4_outputs(3343)));
    layer5_outputs(6752) <= layer4_outputs(4553);
    layer5_outputs(6753) <= not(layer4_outputs(7209));
    layer5_outputs(6754) <= not(layer4_outputs(7092));
    layer5_outputs(6755) <= '0';
    layer5_outputs(6756) <= not(layer4_outputs(2824)) or (layer4_outputs(5650));
    layer5_outputs(6757) <= not(layer4_outputs(3796));
    layer5_outputs(6758) <= not((layer4_outputs(7153)) and (layer4_outputs(175)));
    layer5_outputs(6759) <= (layer4_outputs(7620)) and not (layer4_outputs(1666));
    layer5_outputs(6760) <= not((layer4_outputs(7463)) xor (layer4_outputs(4255)));
    layer5_outputs(6761) <= layer4_outputs(3197);
    layer5_outputs(6762) <= not(layer4_outputs(4358));
    layer5_outputs(6763) <= (layer4_outputs(1845)) and not (layer4_outputs(3561));
    layer5_outputs(6764) <= layer4_outputs(2133);
    layer5_outputs(6765) <= not((layer4_outputs(6748)) xor (layer4_outputs(6299)));
    layer5_outputs(6766) <= not((layer4_outputs(6832)) and (layer4_outputs(6710)));
    layer5_outputs(6767) <= not((layer4_outputs(727)) xor (layer4_outputs(9)));
    layer5_outputs(6768) <= not(layer4_outputs(2175));
    layer5_outputs(6769) <= not((layer4_outputs(4940)) and (layer4_outputs(2573)));
    layer5_outputs(6770) <= not((layer4_outputs(5555)) xor (layer4_outputs(3744)));
    layer5_outputs(6771) <= layer4_outputs(4346);
    layer5_outputs(6772) <= not((layer4_outputs(6866)) xor (layer4_outputs(6348)));
    layer5_outputs(6773) <= layer4_outputs(6941);
    layer5_outputs(6774) <= '1';
    layer5_outputs(6775) <= (layer4_outputs(1550)) and (layer4_outputs(7625));
    layer5_outputs(6776) <= not(layer4_outputs(4592));
    layer5_outputs(6777) <= not(layer4_outputs(3835));
    layer5_outputs(6778) <= not(layer4_outputs(2290));
    layer5_outputs(6779) <= not(layer4_outputs(2100));
    layer5_outputs(6780) <= not(layer4_outputs(3149));
    layer5_outputs(6781) <= not((layer4_outputs(3537)) and (layer4_outputs(5167)));
    layer5_outputs(6782) <= (layer4_outputs(348)) and not (layer4_outputs(2829));
    layer5_outputs(6783) <= layer4_outputs(5238);
    layer5_outputs(6784) <= '1';
    layer5_outputs(6785) <= (layer4_outputs(1120)) or (layer4_outputs(2761));
    layer5_outputs(6786) <= (layer4_outputs(3069)) or (layer4_outputs(1039));
    layer5_outputs(6787) <= not((layer4_outputs(15)) or (layer4_outputs(4123)));
    layer5_outputs(6788) <= (layer4_outputs(4116)) and not (layer4_outputs(6903));
    layer5_outputs(6789) <= not(layer4_outputs(5559));
    layer5_outputs(6790) <= not(layer4_outputs(6808));
    layer5_outputs(6791) <= not((layer4_outputs(3387)) xor (layer4_outputs(834)));
    layer5_outputs(6792) <= (layer4_outputs(6725)) xor (layer4_outputs(3627));
    layer5_outputs(6793) <= (layer4_outputs(2352)) xor (layer4_outputs(2000));
    layer5_outputs(6794) <= not((layer4_outputs(7426)) or (layer4_outputs(4933)));
    layer5_outputs(6795) <= layer4_outputs(1049);
    layer5_outputs(6796) <= not((layer4_outputs(3021)) and (layer4_outputs(6577)));
    layer5_outputs(6797) <= layer4_outputs(3638);
    layer5_outputs(6798) <= not((layer4_outputs(4535)) or (layer4_outputs(3212)));
    layer5_outputs(6799) <= (layer4_outputs(6824)) and (layer4_outputs(6544));
    layer5_outputs(6800) <= layer4_outputs(1856);
    layer5_outputs(6801) <= layer4_outputs(1524);
    layer5_outputs(6802) <= not(layer4_outputs(5787));
    layer5_outputs(6803) <= '1';
    layer5_outputs(6804) <= (layer4_outputs(2344)) xor (layer4_outputs(400));
    layer5_outputs(6805) <= not(layer4_outputs(7324)) or (layer4_outputs(2997));
    layer5_outputs(6806) <= layer4_outputs(6203);
    layer5_outputs(6807) <= layer4_outputs(3919);
    layer5_outputs(6808) <= not((layer4_outputs(6224)) xor (layer4_outputs(4818)));
    layer5_outputs(6809) <= layer4_outputs(2392);
    layer5_outputs(6810) <= not(layer4_outputs(26));
    layer5_outputs(6811) <= layer4_outputs(2670);
    layer5_outputs(6812) <= not(layer4_outputs(1470));
    layer5_outputs(6813) <= layer4_outputs(7273);
    layer5_outputs(6814) <= not(layer4_outputs(4498));
    layer5_outputs(6815) <= not(layer4_outputs(228));
    layer5_outputs(6816) <= not(layer4_outputs(4459));
    layer5_outputs(6817) <= layer4_outputs(6460);
    layer5_outputs(6818) <= '1';
    layer5_outputs(6819) <= layer4_outputs(4212);
    layer5_outputs(6820) <= not(layer4_outputs(815));
    layer5_outputs(6821) <= layer4_outputs(5410);
    layer5_outputs(6822) <= not(layer4_outputs(6520));
    layer5_outputs(6823) <= not(layer4_outputs(817)) or (layer4_outputs(2933));
    layer5_outputs(6824) <= not(layer4_outputs(4894));
    layer5_outputs(6825) <= layer4_outputs(231);
    layer5_outputs(6826) <= (layer4_outputs(7068)) or (layer4_outputs(96));
    layer5_outputs(6827) <= (layer4_outputs(7175)) and not (layer4_outputs(3059));
    layer5_outputs(6828) <= not(layer4_outputs(5675));
    layer5_outputs(6829) <= not(layer4_outputs(3336));
    layer5_outputs(6830) <= (layer4_outputs(527)) or (layer4_outputs(2554));
    layer5_outputs(6831) <= not(layer4_outputs(4711));
    layer5_outputs(6832) <= (layer4_outputs(2252)) xor (layer4_outputs(5827));
    layer5_outputs(6833) <= (layer4_outputs(373)) and not (layer4_outputs(2630));
    layer5_outputs(6834) <= '1';
    layer5_outputs(6835) <= not((layer4_outputs(330)) xor (layer4_outputs(2673)));
    layer5_outputs(6836) <= not((layer4_outputs(5150)) xor (layer4_outputs(442)));
    layer5_outputs(6837) <= (layer4_outputs(7225)) or (layer4_outputs(5373));
    layer5_outputs(6838) <= not(layer4_outputs(698));
    layer5_outputs(6839) <= layer4_outputs(2007);
    layer5_outputs(6840) <= not(layer4_outputs(2654)) or (layer4_outputs(520));
    layer5_outputs(6841) <= layer4_outputs(5495);
    layer5_outputs(6842) <= layer4_outputs(6883);
    layer5_outputs(6843) <= not(layer4_outputs(341));
    layer5_outputs(6844) <= '1';
    layer5_outputs(6845) <= '0';
    layer5_outputs(6846) <= not(layer4_outputs(2883));
    layer5_outputs(6847) <= not(layer4_outputs(2340));
    layer5_outputs(6848) <= '1';
    layer5_outputs(6849) <= layer4_outputs(3923);
    layer5_outputs(6850) <= layer4_outputs(2652);
    layer5_outputs(6851) <= layer4_outputs(4194);
    layer5_outputs(6852) <= not(layer4_outputs(2023));
    layer5_outputs(6853) <= (layer4_outputs(6916)) and not (layer4_outputs(3944));
    layer5_outputs(6854) <= (layer4_outputs(4434)) or (layer4_outputs(3644));
    layer5_outputs(6855) <= not(layer4_outputs(7594));
    layer5_outputs(6856) <= not(layer4_outputs(3918));
    layer5_outputs(6857) <= layer4_outputs(1297);
    layer5_outputs(6858) <= not(layer4_outputs(1731));
    layer5_outputs(6859) <= layer4_outputs(5864);
    layer5_outputs(6860) <= not(layer4_outputs(2286));
    layer5_outputs(6861) <= not(layer4_outputs(7447));
    layer5_outputs(6862) <= (layer4_outputs(6904)) and not (layer4_outputs(7435));
    layer5_outputs(6863) <= (layer4_outputs(3785)) xor (layer4_outputs(6854));
    layer5_outputs(6864) <= not((layer4_outputs(6332)) xor (layer4_outputs(2912)));
    layer5_outputs(6865) <= not((layer4_outputs(3051)) and (layer4_outputs(6189)));
    layer5_outputs(6866) <= not(layer4_outputs(7545));
    layer5_outputs(6867) <= not(layer4_outputs(6274));
    layer5_outputs(6868) <= not(layer4_outputs(403));
    layer5_outputs(6869) <= not(layer4_outputs(2490));
    layer5_outputs(6870) <= not(layer4_outputs(7542)) or (layer4_outputs(4627));
    layer5_outputs(6871) <= not((layer4_outputs(5996)) or (layer4_outputs(3312)));
    layer5_outputs(6872) <= not(layer4_outputs(7285));
    layer5_outputs(6873) <= layer4_outputs(771);
    layer5_outputs(6874) <= not(layer4_outputs(556));
    layer5_outputs(6875) <= layer4_outputs(7429);
    layer5_outputs(6876) <= layer4_outputs(3608);
    layer5_outputs(6877) <= not(layer4_outputs(7015));
    layer5_outputs(6878) <= (layer4_outputs(2277)) and (layer4_outputs(1397));
    layer5_outputs(6879) <= not(layer4_outputs(2180));
    layer5_outputs(6880) <= layer4_outputs(430);
    layer5_outputs(6881) <= '1';
    layer5_outputs(6882) <= not(layer4_outputs(1884));
    layer5_outputs(6883) <= '0';
    layer5_outputs(6884) <= not(layer4_outputs(2234)) or (layer4_outputs(4902));
    layer5_outputs(6885) <= '1';
    layer5_outputs(6886) <= not(layer4_outputs(4570));
    layer5_outputs(6887) <= not(layer4_outputs(1067));
    layer5_outputs(6888) <= not(layer4_outputs(7183));
    layer5_outputs(6889) <= layer4_outputs(6892);
    layer5_outputs(6890) <= layer4_outputs(6051);
    layer5_outputs(6891) <= (layer4_outputs(7438)) and not (layer4_outputs(6741));
    layer5_outputs(6892) <= layer4_outputs(1400);
    layer5_outputs(6893) <= layer4_outputs(1314);
    layer5_outputs(6894) <= layer4_outputs(20);
    layer5_outputs(6895) <= not(layer4_outputs(6528));
    layer5_outputs(6896) <= layer4_outputs(3128);
    layer5_outputs(6897) <= layer4_outputs(7089);
    layer5_outputs(6898) <= not(layer4_outputs(3995));
    layer5_outputs(6899) <= not(layer4_outputs(5185));
    layer5_outputs(6900) <= layer4_outputs(2051);
    layer5_outputs(6901) <= (layer4_outputs(7303)) and not (layer4_outputs(62));
    layer5_outputs(6902) <= layer4_outputs(2314);
    layer5_outputs(6903) <= (layer4_outputs(3102)) and not (layer4_outputs(132));
    layer5_outputs(6904) <= not(layer4_outputs(6153));
    layer5_outputs(6905) <= (layer4_outputs(329)) and (layer4_outputs(2773));
    layer5_outputs(6906) <= not((layer4_outputs(7358)) or (layer4_outputs(3833)));
    layer5_outputs(6907) <= not(layer4_outputs(3119));
    layer5_outputs(6908) <= not(layer4_outputs(3412));
    layer5_outputs(6909) <= not(layer4_outputs(7150));
    layer5_outputs(6910) <= not(layer4_outputs(1382));
    layer5_outputs(6911) <= layer4_outputs(6712);
    layer5_outputs(6912) <= layer4_outputs(916);
    layer5_outputs(6913) <= not(layer4_outputs(1648));
    layer5_outputs(6914) <= (layer4_outputs(846)) and not (layer4_outputs(383));
    layer5_outputs(6915) <= layer4_outputs(3463);
    layer5_outputs(6916) <= not(layer4_outputs(7134)) or (layer4_outputs(5529));
    layer5_outputs(6917) <= not(layer4_outputs(5277));
    layer5_outputs(6918) <= layer4_outputs(390);
    layer5_outputs(6919) <= layer4_outputs(1166);
    layer5_outputs(6920) <= not(layer4_outputs(1234));
    layer5_outputs(6921) <= layer4_outputs(2955);
    layer5_outputs(6922) <= layer4_outputs(1663);
    layer5_outputs(6923) <= not(layer4_outputs(6415));
    layer5_outputs(6924) <= layer4_outputs(2904);
    layer5_outputs(6925) <= not((layer4_outputs(4673)) or (layer4_outputs(2726)));
    layer5_outputs(6926) <= not(layer4_outputs(5910)) or (layer4_outputs(3881));
    layer5_outputs(6927) <= layer4_outputs(1368);
    layer5_outputs(6928) <= (layer4_outputs(3418)) or (layer4_outputs(2220));
    layer5_outputs(6929) <= not(layer4_outputs(1032));
    layer5_outputs(6930) <= layer4_outputs(4623);
    layer5_outputs(6931) <= (layer4_outputs(6955)) and not (layer4_outputs(5037));
    layer5_outputs(6932) <= (layer4_outputs(1314)) or (layer4_outputs(2135));
    layer5_outputs(6933) <= (layer4_outputs(7341)) or (layer4_outputs(80));
    layer5_outputs(6934) <= (layer4_outputs(6511)) xor (layer4_outputs(3261));
    layer5_outputs(6935) <= not(layer4_outputs(6172));
    layer5_outputs(6936) <= layer4_outputs(7048);
    layer5_outputs(6937) <= layer4_outputs(6539);
    layer5_outputs(6938) <= layer4_outputs(2067);
    layer5_outputs(6939) <= not(layer4_outputs(7618));
    layer5_outputs(6940) <= not((layer4_outputs(2358)) and (layer4_outputs(3562)));
    layer5_outputs(6941) <= (layer4_outputs(4043)) and (layer4_outputs(3492));
    layer5_outputs(6942) <= not(layer4_outputs(4069));
    layer5_outputs(6943) <= not((layer4_outputs(2057)) and (layer4_outputs(4122)));
    layer5_outputs(6944) <= not(layer4_outputs(3250));
    layer5_outputs(6945) <= not((layer4_outputs(4683)) xor (layer4_outputs(1570)));
    layer5_outputs(6946) <= layer4_outputs(3000);
    layer5_outputs(6947) <= not((layer4_outputs(4003)) and (layer4_outputs(5436)));
    layer5_outputs(6948) <= not(layer4_outputs(920));
    layer5_outputs(6949) <= not(layer4_outputs(3251));
    layer5_outputs(6950) <= layer4_outputs(2938);
    layer5_outputs(6951) <= not(layer4_outputs(553)) or (layer4_outputs(6658));
    layer5_outputs(6952) <= not(layer4_outputs(4488));
    layer5_outputs(6953) <= layer4_outputs(4459);
    layer5_outputs(6954) <= (layer4_outputs(4595)) and not (layer4_outputs(3882));
    layer5_outputs(6955) <= layer4_outputs(5536);
    layer5_outputs(6956) <= not(layer4_outputs(5854)) or (layer4_outputs(540));
    layer5_outputs(6957) <= not(layer4_outputs(2219));
    layer5_outputs(6958) <= not(layer4_outputs(1144));
    layer5_outputs(6959) <= not(layer4_outputs(4831));
    layer5_outputs(6960) <= not(layer4_outputs(4290)) or (layer4_outputs(2603));
    layer5_outputs(6961) <= (layer4_outputs(5210)) and not (layer4_outputs(3017));
    layer5_outputs(6962) <= not((layer4_outputs(1129)) xor (layer4_outputs(1959)));
    layer5_outputs(6963) <= not(layer4_outputs(2595)) or (layer4_outputs(707));
    layer5_outputs(6964) <= not(layer4_outputs(6359));
    layer5_outputs(6965) <= not(layer4_outputs(5213)) or (layer4_outputs(3884));
    layer5_outputs(6966) <= not(layer4_outputs(3817)) or (layer4_outputs(154));
    layer5_outputs(6967) <= layer4_outputs(3942);
    layer5_outputs(6968) <= layer4_outputs(2623);
    layer5_outputs(6969) <= (layer4_outputs(662)) or (layer4_outputs(2977));
    layer5_outputs(6970) <= layer4_outputs(7110);
    layer5_outputs(6971) <= (layer4_outputs(1121)) and not (layer4_outputs(7139));
    layer5_outputs(6972) <= not(layer4_outputs(2545));
    layer5_outputs(6973) <= (layer4_outputs(176)) and (layer4_outputs(6525));
    layer5_outputs(6974) <= (layer4_outputs(4817)) xor (layer4_outputs(3685));
    layer5_outputs(6975) <= layer4_outputs(173);
    layer5_outputs(6976) <= not((layer4_outputs(5055)) or (layer4_outputs(591)));
    layer5_outputs(6977) <= layer4_outputs(5169);
    layer5_outputs(6978) <= layer4_outputs(5297);
    layer5_outputs(6979) <= '1';
    layer5_outputs(6980) <= layer4_outputs(513);
    layer5_outputs(6981) <= layer4_outputs(3110);
    layer5_outputs(6982) <= not(layer4_outputs(1847));
    layer5_outputs(6983) <= (layer4_outputs(6151)) xor (layer4_outputs(4825));
    layer5_outputs(6984) <= (layer4_outputs(5287)) and not (layer4_outputs(6564));
    layer5_outputs(6985) <= (layer4_outputs(7212)) xor (layer4_outputs(2695));
    layer5_outputs(6986) <= (layer4_outputs(6502)) and not (layer4_outputs(3774));
    layer5_outputs(6987) <= not((layer4_outputs(4268)) xor (layer4_outputs(6804)));
    layer5_outputs(6988) <= not(layer4_outputs(4799));
    layer5_outputs(6989) <= (layer4_outputs(1979)) xor (layer4_outputs(1643));
    layer5_outputs(6990) <= (layer4_outputs(829)) xor (layer4_outputs(2637));
    layer5_outputs(6991) <= not(layer4_outputs(714)) or (layer4_outputs(3214));
    layer5_outputs(6992) <= not(layer4_outputs(6210)) or (layer4_outputs(2207));
    layer5_outputs(6993) <= (layer4_outputs(4415)) and not (layer4_outputs(7133));
    layer5_outputs(6994) <= (layer4_outputs(184)) or (layer4_outputs(4871));
    layer5_outputs(6995) <= (layer4_outputs(3691)) and not (layer4_outputs(38));
    layer5_outputs(6996) <= not(layer4_outputs(5490));
    layer5_outputs(6997) <= not((layer4_outputs(721)) and (layer4_outputs(3094)));
    layer5_outputs(6998) <= (layer4_outputs(539)) or (layer4_outputs(5635));
    layer5_outputs(6999) <= not(layer4_outputs(258));
    layer5_outputs(7000) <= (layer4_outputs(3868)) and not (layer4_outputs(2658));
    layer5_outputs(7001) <= not((layer4_outputs(4036)) and (layer4_outputs(2828)));
    layer5_outputs(7002) <= not(layer4_outputs(6023));
    layer5_outputs(7003) <= not((layer4_outputs(7493)) xor (layer4_outputs(2828)));
    layer5_outputs(7004) <= (layer4_outputs(5564)) xor (layer4_outputs(6701));
    layer5_outputs(7005) <= (layer4_outputs(4011)) and (layer4_outputs(1983));
    layer5_outputs(7006) <= not(layer4_outputs(5330));
    layer5_outputs(7007) <= '0';
    layer5_outputs(7008) <= (layer4_outputs(4863)) and (layer4_outputs(6464));
    layer5_outputs(7009) <= layer4_outputs(3459);
    layer5_outputs(7010) <= (layer4_outputs(5618)) or (layer4_outputs(6158));
    layer5_outputs(7011) <= not(layer4_outputs(3145));
    layer5_outputs(7012) <= (layer4_outputs(5834)) and not (layer4_outputs(6374));
    layer5_outputs(7013) <= not((layer4_outputs(3156)) and (layer4_outputs(6553)));
    layer5_outputs(7014) <= not(layer4_outputs(7357)) or (layer4_outputs(4665));
    layer5_outputs(7015) <= not(layer4_outputs(864)) or (layer4_outputs(3684));
    layer5_outputs(7016) <= not((layer4_outputs(605)) or (layer4_outputs(1307)));
    layer5_outputs(7017) <= layer4_outputs(3187);
    layer5_outputs(7018) <= not(layer4_outputs(6121));
    layer5_outputs(7019) <= not(layer4_outputs(3659));
    layer5_outputs(7020) <= (layer4_outputs(3140)) and not (layer4_outputs(453));
    layer5_outputs(7021) <= (layer4_outputs(3305)) or (layer4_outputs(7206));
    layer5_outputs(7022) <= (layer4_outputs(1484)) and (layer4_outputs(5763));
    layer5_outputs(7023) <= (layer4_outputs(6385)) xor (layer4_outputs(4528));
    layer5_outputs(7024) <= layer4_outputs(5196);
    layer5_outputs(7025) <= layer4_outputs(5716);
    layer5_outputs(7026) <= (layer4_outputs(6536)) and not (layer4_outputs(7278));
    layer5_outputs(7027) <= (layer4_outputs(2494)) and not (layer4_outputs(2896));
    layer5_outputs(7028) <= layer4_outputs(6671);
    layer5_outputs(7029) <= not(layer4_outputs(6655));
    layer5_outputs(7030) <= layer4_outputs(4308);
    layer5_outputs(7031) <= '0';
    layer5_outputs(7032) <= (layer4_outputs(2522)) and not (layer4_outputs(4758));
    layer5_outputs(7033) <= not(layer4_outputs(3631));
    layer5_outputs(7034) <= (layer4_outputs(4657)) and not (layer4_outputs(3456));
    layer5_outputs(7035) <= not((layer4_outputs(4460)) and (layer4_outputs(468)));
    layer5_outputs(7036) <= (layer4_outputs(1871)) xor (layer4_outputs(130));
    layer5_outputs(7037) <= (layer4_outputs(3355)) and not (layer4_outputs(2978));
    layer5_outputs(7038) <= not((layer4_outputs(6283)) xor (layer4_outputs(242)));
    layer5_outputs(7039) <= not(layer4_outputs(108));
    layer5_outputs(7040) <= (layer4_outputs(6731)) and not (layer4_outputs(7422));
    layer5_outputs(7041) <= not(layer4_outputs(7393));
    layer5_outputs(7042) <= not((layer4_outputs(3530)) or (layer4_outputs(4255)));
    layer5_outputs(7043) <= not(layer4_outputs(3638));
    layer5_outputs(7044) <= not(layer4_outputs(6516));
    layer5_outputs(7045) <= (layer4_outputs(6037)) or (layer4_outputs(2757));
    layer5_outputs(7046) <= not(layer4_outputs(685));
    layer5_outputs(7047) <= layer4_outputs(716);
    layer5_outputs(7048) <= (layer4_outputs(5966)) or (layer4_outputs(4672));
    layer5_outputs(7049) <= not(layer4_outputs(3653)) or (layer4_outputs(6024));
    layer5_outputs(7050) <= layer4_outputs(432);
    layer5_outputs(7051) <= (layer4_outputs(556)) and not (layer4_outputs(1172));
    layer5_outputs(7052) <= (layer4_outputs(1307)) xor (layer4_outputs(4380));
    layer5_outputs(7053) <= (layer4_outputs(4322)) or (layer4_outputs(1117));
    layer5_outputs(7054) <= not(layer4_outputs(1208));
    layer5_outputs(7055) <= not((layer4_outputs(7528)) xor (layer4_outputs(4281)));
    layer5_outputs(7056) <= not(layer4_outputs(5023));
    layer5_outputs(7057) <= not(layer4_outputs(2884));
    layer5_outputs(7058) <= not(layer4_outputs(6546)) or (layer4_outputs(1164));
    layer5_outputs(7059) <= layer4_outputs(2190);
    layer5_outputs(7060) <= (layer4_outputs(5641)) xor (layer4_outputs(2869));
    layer5_outputs(7061) <= not(layer4_outputs(1051));
    layer5_outputs(7062) <= layer4_outputs(1128);
    layer5_outputs(7063) <= not(layer4_outputs(6474)) or (layer4_outputs(5557));
    layer5_outputs(7064) <= not(layer4_outputs(4624));
    layer5_outputs(7065) <= layer4_outputs(4582);
    layer5_outputs(7066) <= not(layer4_outputs(2784));
    layer5_outputs(7067) <= (layer4_outputs(1690)) xor (layer4_outputs(5599));
    layer5_outputs(7068) <= layer4_outputs(570);
    layer5_outputs(7069) <= (layer4_outputs(6805)) xor (layer4_outputs(6990));
    layer5_outputs(7070) <= (layer4_outputs(2826)) and not (layer4_outputs(7531));
    layer5_outputs(7071) <= layer4_outputs(4372);
    layer5_outputs(7072) <= layer4_outputs(3437);
    layer5_outputs(7073) <= not(layer4_outputs(1514));
    layer5_outputs(7074) <= (layer4_outputs(5476)) and (layer4_outputs(356));
    layer5_outputs(7075) <= not(layer4_outputs(5338)) or (layer4_outputs(6147));
    layer5_outputs(7076) <= '1';
    layer5_outputs(7077) <= '1';
    layer5_outputs(7078) <= not(layer4_outputs(5494)) or (layer4_outputs(4013));
    layer5_outputs(7079) <= (layer4_outputs(5721)) and not (layer4_outputs(5249));
    layer5_outputs(7080) <= layer4_outputs(6263);
    layer5_outputs(7081) <= layer4_outputs(3164);
    layer5_outputs(7082) <= not((layer4_outputs(757)) and (layer4_outputs(2547)));
    layer5_outputs(7083) <= layer4_outputs(460);
    layer5_outputs(7084) <= (layer4_outputs(199)) or (layer4_outputs(4609));
    layer5_outputs(7085) <= layer4_outputs(6891);
    layer5_outputs(7086) <= layer4_outputs(5869);
    layer5_outputs(7087) <= (layer4_outputs(5142)) or (layer4_outputs(5576));
    layer5_outputs(7088) <= not(layer4_outputs(1013)) or (layer4_outputs(1708));
    layer5_outputs(7089) <= (layer4_outputs(2106)) xor (layer4_outputs(4820));
    layer5_outputs(7090) <= not(layer4_outputs(6144)) or (layer4_outputs(4985));
    layer5_outputs(7091) <= layer4_outputs(7466);
    layer5_outputs(7092) <= not(layer4_outputs(3201));
    layer5_outputs(7093) <= (layer4_outputs(325)) and (layer4_outputs(1726));
    layer5_outputs(7094) <= not((layer4_outputs(6770)) xor (layer4_outputs(120)));
    layer5_outputs(7095) <= not(layer4_outputs(1488));
    layer5_outputs(7096) <= not(layer4_outputs(1880)) or (layer4_outputs(5660));
    layer5_outputs(7097) <= layer4_outputs(3928);
    layer5_outputs(7098) <= layer4_outputs(4969);
    layer5_outputs(7099) <= not((layer4_outputs(6289)) and (layer4_outputs(7628)));
    layer5_outputs(7100) <= (layer4_outputs(2632)) and not (layer4_outputs(159));
    layer5_outputs(7101) <= layer4_outputs(5325);
    layer5_outputs(7102) <= (layer4_outputs(4816)) or (layer4_outputs(1038));
    layer5_outputs(7103) <= not((layer4_outputs(3912)) and (layer4_outputs(6179)));
    layer5_outputs(7104) <= layer4_outputs(981);
    layer5_outputs(7105) <= (layer4_outputs(6894)) and not (layer4_outputs(5320));
    layer5_outputs(7106) <= '1';
    layer5_outputs(7107) <= (layer4_outputs(7525)) or (layer4_outputs(6513));
    layer5_outputs(7108) <= not(layer4_outputs(4480)) or (layer4_outputs(7330));
    layer5_outputs(7109) <= (layer4_outputs(4156)) and (layer4_outputs(7051));
    layer5_outputs(7110) <= layer4_outputs(6704);
    layer5_outputs(7111) <= layer4_outputs(1171);
    layer5_outputs(7112) <= not(layer4_outputs(2243));
    layer5_outputs(7113) <= (layer4_outputs(4575)) xor (layer4_outputs(2693));
    layer5_outputs(7114) <= layer4_outputs(358);
    layer5_outputs(7115) <= not(layer4_outputs(3277));
    layer5_outputs(7116) <= not(layer4_outputs(6799));
    layer5_outputs(7117) <= (layer4_outputs(6411)) and not (layer4_outputs(2612));
    layer5_outputs(7118) <= not((layer4_outputs(2671)) xor (layer4_outputs(3328)));
    layer5_outputs(7119) <= not(layer4_outputs(2914));
    layer5_outputs(7120) <= layer4_outputs(5757);
    layer5_outputs(7121) <= not(layer4_outputs(6477));
    layer5_outputs(7122) <= '1';
    layer5_outputs(7123) <= not(layer4_outputs(209));
    layer5_outputs(7124) <= (layer4_outputs(6630)) and not (layer4_outputs(1360));
    layer5_outputs(7125) <= not(layer4_outputs(5828));
    layer5_outputs(7126) <= layer4_outputs(1574);
    layer5_outputs(7127) <= not(layer4_outputs(1253));
    layer5_outputs(7128) <= (layer4_outputs(2353)) and not (layer4_outputs(4882));
    layer5_outputs(7129) <= (layer4_outputs(3446)) and not (layer4_outputs(1264));
    layer5_outputs(7130) <= not(layer4_outputs(772));
    layer5_outputs(7131) <= (layer4_outputs(5057)) or (layer4_outputs(1699));
    layer5_outputs(7132) <= (layer4_outputs(2182)) and not (layer4_outputs(7242));
    layer5_outputs(7133) <= not(layer4_outputs(380)) or (layer4_outputs(2775));
    layer5_outputs(7134) <= not((layer4_outputs(3139)) xor (layer4_outputs(7541)));
    layer5_outputs(7135) <= not(layer4_outputs(6360)) or (layer4_outputs(2878));
    layer5_outputs(7136) <= layer4_outputs(4477);
    layer5_outputs(7137) <= not((layer4_outputs(1078)) and (layer4_outputs(1868)));
    layer5_outputs(7138) <= layer4_outputs(5542);
    layer5_outputs(7139) <= (layer4_outputs(2795)) and not (layer4_outputs(4198));
    layer5_outputs(7140) <= layer4_outputs(7526);
    layer5_outputs(7141) <= '1';
    layer5_outputs(7142) <= (layer4_outputs(7225)) and not (layer4_outputs(3445));
    layer5_outputs(7143) <= not((layer4_outputs(176)) xor (layer4_outputs(5543)));
    layer5_outputs(7144) <= (layer4_outputs(5966)) or (layer4_outputs(6159));
    layer5_outputs(7145) <= not((layer4_outputs(6330)) and (layer4_outputs(3333)));
    layer5_outputs(7146) <= layer4_outputs(4504);
    layer5_outputs(7147) <= (layer4_outputs(3727)) and not (layer4_outputs(1799));
    layer5_outputs(7148) <= not((layer4_outputs(6677)) or (layer4_outputs(583)));
    layer5_outputs(7149) <= '1';
    layer5_outputs(7150) <= layer4_outputs(3780);
    layer5_outputs(7151) <= not(layer4_outputs(3180));
    layer5_outputs(7152) <= not(layer4_outputs(2176)) or (layer4_outputs(5466));
    layer5_outputs(7153) <= not((layer4_outputs(2398)) and (layer4_outputs(7405)));
    layer5_outputs(7154) <= not(layer4_outputs(5591));
    layer5_outputs(7155) <= not((layer4_outputs(2135)) and (layer4_outputs(3333)));
    layer5_outputs(7156) <= not(layer4_outputs(3370));
    layer5_outputs(7157) <= not(layer4_outputs(1290)) or (layer4_outputs(3253));
    layer5_outputs(7158) <= not(layer4_outputs(1217));
    layer5_outputs(7159) <= not((layer4_outputs(2413)) and (layer4_outputs(7231)));
    layer5_outputs(7160) <= (layer4_outputs(4987)) and not (layer4_outputs(3819));
    layer5_outputs(7161) <= layer4_outputs(1972);
    layer5_outputs(7162) <= layer4_outputs(723);
    layer5_outputs(7163) <= not(layer4_outputs(2860));
    layer5_outputs(7164) <= not(layer4_outputs(6636));
    layer5_outputs(7165) <= (layer4_outputs(5800)) or (layer4_outputs(3928));
    layer5_outputs(7166) <= not((layer4_outputs(2180)) xor (layer4_outputs(4861)));
    layer5_outputs(7167) <= layer4_outputs(1429);
    layer5_outputs(7168) <= (layer4_outputs(563)) and (layer4_outputs(4047));
    layer5_outputs(7169) <= layer4_outputs(1854);
    layer5_outputs(7170) <= (layer4_outputs(2156)) and not (layer4_outputs(6150));
    layer5_outputs(7171) <= not((layer4_outputs(79)) or (layer4_outputs(6006)));
    layer5_outputs(7172) <= layer4_outputs(857);
    layer5_outputs(7173) <= (layer4_outputs(5261)) and not (layer4_outputs(5898));
    layer5_outputs(7174) <= not(layer4_outputs(6353));
    layer5_outputs(7175) <= (layer4_outputs(4209)) xor (layer4_outputs(4388));
    layer5_outputs(7176) <= layer4_outputs(5472);
    layer5_outputs(7177) <= layer4_outputs(592);
    layer5_outputs(7178) <= not(layer4_outputs(5976));
    layer5_outputs(7179) <= layer4_outputs(1564);
    layer5_outputs(7180) <= layer4_outputs(7036);
    layer5_outputs(7181) <= not((layer4_outputs(3292)) or (layer4_outputs(7632)));
    layer5_outputs(7182) <= (layer4_outputs(2885)) and not (layer4_outputs(705));
    layer5_outputs(7183) <= not(layer4_outputs(6827)) or (layer4_outputs(7278));
    layer5_outputs(7184) <= not(layer4_outputs(253));
    layer5_outputs(7185) <= not(layer4_outputs(5776));
    layer5_outputs(7186) <= not(layer4_outputs(5658));
    layer5_outputs(7187) <= (layer4_outputs(4876)) or (layer4_outputs(6015));
    layer5_outputs(7188) <= (layer4_outputs(6646)) xor (layer4_outputs(4569));
    layer5_outputs(7189) <= not((layer4_outputs(1994)) and (layer4_outputs(7625)));
    layer5_outputs(7190) <= layer4_outputs(1312);
    layer5_outputs(7191) <= '0';
    layer5_outputs(7192) <= not(layer4_outputs(51)) or (layer4_outputs(4881));
    layer5_outputs(7193) <= layer4_outputs(7137);
    layer5_outputs(7194) <= not((layer4_outputs(777)) xor (layer4_outputs(3267)));
    layer5_outputs(7195) <= layer4_outputs(2184);
    layer5_outputs(7196) <= not(layer4_outputs(173));
    layer5_outputs(7197) <= not(layer4_outputs(4172));
    layer5_outputs(7198) <= layer4_outputs(7454);
    layer5_outputs(7199) <= not((layer4_outputs(7387)) and (layer4_outputs(239)));
    layer5_outputs(7200) <= (layer4_outputs(5874)) or (layer4_outputs(5602));
    layer5_outputs(7201) <= not(layer4_outputs(6440)) or (layer4_outputs(5070));
    layer5_outputs(7202) <= (layer4_outputs(5841)) and not (layer4_outputs(3585));
    layer5_outputs(7203) <= (layer4_outputs(5809)) and not (layer4_outputs(5895));
    layer5_outputs(7204) <= not(layer4_outputs(476));
    layer5_outputs(7205) <= (layer4_outputs(4517)) xor (layer4_outputs(6250));
    layer5_outputs(7206) <= not(layer4_outputs(3374)) or (layer4_outputs(5141));
    layer5_outputs(7207) <= not(layer4_outputs(7119));
    layer5_outputs(7208) <= (layer4_outputs(2237)) xor (layer4_outputs(2327));
    layer5_outputs(7209) <= not((layer4_outputs(1748)) or (layer4_outputs(5048)));
    layer5_outputs(7210) <= '1';
    layer5_outputs(7211) <= not(layer4_outputs(1103));
    layer5_outputs(7212) <= (layer4_outputs(578)) xor (layer4_outputs(1687));
    layer5_outputs(7213) <= (layer4_outputs(3468)) and not (layer4_outputs(5158));
    layer5_outputs(7214) <= (layer4_outputs(2613)) and (layer4_outputs(299));
    layer5_outputs(7215) <= not((layer4_outputs(2074)) or (layer4_outputs(4260)));
    layer5_outputs(7216) <= (layer4_outputs(3885)) xor (layer4_outputs(2727));
    layer5_outputs(7217) <= (layer4_outputs(3152)) and (layer4_outputs(2892));
    layer5_outputs(7218) <= layer4_outputs(4946);
    layer5_outputs(7219) <= not(layer4_outputs(7122));
    layer5_outputs(7220) <= layer4_outputs(3314);
    layer5_outputs(7221) <= layer4_outputs(3387);
    layer5_outputs(7222) <= layer4_outputs(221);
    layer5_outputs(7223) <= layer4_outputs(2675);
    layer5_outputs(7224) <= (layer4_outputs(4505)) and not (layer4_outputs(5454));
    layer5_outputs(7225) <= not(layer4_outputs(4682));
    layer5_outputs(7226) <= not(layer4_outputs(2908));
    layer5_outputs(7227) <= layer4_outputs(8);
    layer5_outputs(7228) <= not((layer4_outputs(4409)) xor (layer4_outputs(5592)));
    layer5_outputs(7229) <= layer4_outputs(11);
    layer5_outputs(7230) <= not(layer4_outputs(1098)) or (layer4_outputs(765));
    layer5_outputs(7231) <= layer4_outputs(1471);
    layer5_outputs(7232) <= not((layer4_outputs(6497)) xor (layer4_outputs(849)));
    layer5_outputs(7233) <= not(layer4_outputs(7677));
    layer5_outputs(7234) <= layer4_outputs(1617);
    layer5_outputs(7235) <= not(layer4_outputs(5267)) or (layer4_outputs(1152));
    layer5_outputs(7236) <= layer4_outputs(4530);
    layer5_outputs(7237) <= layer4_outputs(5276);
    layer5_outputs(7238) <= layer4_outputs(6921);
    layer5_outputs(7239) <= not(layer4_outputs(1665));
    layer5_outputs(7240) <= (layer4_outputs(6221)) or (layer4_outputs(2119));
    layer5_outputs(7241) <= layer4_outputs(6932);
    layer5_outputs(7242) <= layer4_outputs(4086);
    layer5_outputs(7243) <= layer4_outputs(2232);
    layer5_outputs(7244) <= not(layer4_outputs(1811)) or (layer4_outputs(7372));
    layer5_outputs(7245) <= not(layer4_outputs(5557)) or (layer4_outputs(5558));
    layer5_outputs(7246) <= not((layer4_outputs(2175)) xor (layer4_outputs(4395)));
    layer5_outputs(7247) <= (layer4_outputs(6086)) and not (layer4_outputs(757));
    layer5_outputs(7248) <= not((layer4_outputs(1847)) and (layer4_outputs(5241)));
    layer5_outputs(7249) <= (layer4_outputs(1432)) and not (layer4_outputs(5948));
    layer5_outputs(7250) <= layer4_outputs(3346);
    layer5_outputs(7251) <= (layer4_outputs(6680)) or (layer4_outputs(172));
    layer5_outputs(7252) <= not(layer4_outputs(7556));
    layer5_outputs(7253) <= layer4_outputs(2239);
    layer5_outputs(7254) <= not(layer4_outputs(6256));
    layer5_outputs(7255) <= not(layer4_outputs(1409));
    layer5_outputs(7256) <= (layer4_outputs(727)) and not (layer4_outputs(4662));
    layer5_outputs(7257) <= layer4_outputs(1330);
    layer5_outputs(7258) <= layer4_outputs(359);
    layer5_outputs(7259) <= not(layer4_outputs(3232));
    layer5_outputs(7260) <= layer4_outputs(4138);
    layer5_outputs(7261) <= layer4_outputs(4262);
    layer5_outputs(7262) <= not((layer4_outputs(444)) and (layer4_outputs(4414)));
    layer5_outputs(7263) <= (layer4_outputs(6904)) xor (layer4_outputs(5702));
    layer5_outputs(7264) <= not(layer4_outputs(5486));
    layer5_outputs(7265) <= layer4_outputs(1849);
    layer5_outputs(7266) <= layer4_outputs(3897);
    layer5_outputs(7267) <= '1';
    layer5_outputs(7268) <= layer4_outputs(368);
    layer5_outputs(7269) <= layer4_outputs(7616);
    layer5_outputs(7270) <= layer4_outputs(1024);
    layer5_outputs(7271) <= layer4_outputs(5789);
    layer5_outputs(7272) <= not(layer4_outputs(2460));
    layer5_outputs(7273) <= not((layer4_outputs(4824)) or (layer4_outputs(2557)));
    layer5_outputs(7274) <= layer4_outputs(5926);
    layer5_outputs(7275) <= layer4_outputs(5240);
    layer5_outputs(7276) <= not(layer4_outputs(1229));
    layer5_outputs(7277) <= layer4_outputs(4927);
    layer5_outputs(7278) <= layer4_outputs(3655);
    layer5_outputs(7279) <= not(layer4_outputs(4890));
    layer5_outputs(7280) <= not((layer4_outputs(3921)) xor (layer4_outputs(6376)));
    layer5_outputs(7281) <= (layer4_outputs(6962)) and (layer4_outputs(3730));
    layer5_outputs(7282) <= layer4_outputs(4575);
    layer5_outputs(7283) <= layer4_outputs(2564);
    layer5_outputs(7284) <= '0';
    layer5_outputs(7285) <= not(layer4_outputs(1602));
    layer5_outputs(7286) <= layer4_outputs(3852);
    layer5_outputs(7287) <= layer4_outputs(4236);
    layer5_outputs(7288) <= not(layer4_outputs(382));
    layer5_outputs(7289) <= not(layer4_outputs(3105));
    layer5_outputs(7290) <= layer4_outputs(4982);
    layer5_outputs(7291) <= (layer4_outputs(4856)) and not (layer4_outputs(6835));
    layer5_outputs(7292) <= (layer4_outputs(6479)) xor (layer4_outputs(5384));
    layer5_outputs(7293) <= (layer4_outputs(7465)) and not (layer4_outputs(347));
    layer5_outputs(7294) <= layer4_outputs(393);
    layer5_outputs(7295) <= layer4_outputs(6487);
    layer5_outputs(7296) <= layer4_outputs(5694);
    layer5_outputs(7297) <= not(layer4_outputs(3936)) or (layer4_outputs(4080));
    layer5_outputs(7298) <= not((layer4_outputs(7519)) or (layer4_outputs(2250)));
    layer5_outputs(7299) <= not(layer4_outputs(6051));
    layer5_outputs(7300) <= not(layer4_outputs(1055));
    layer5_outputs(7301) <= layer4_outputs(4738);
    layer5_outputs(7302) <= (layer4_outputs(3248)) and (layer4_outputs(5877));
    layer5_outputs(7303) <= not(layer4_outputs(3706));
    layer5_outputs(7304) <= not((layer4_outputs(1048)) and (layer4_outputs(386)));
    layer5_outputs(7305) <= not((layer4_outputs(4949)) xor (layer4_outputs(1352)));
    layer5_outputs(7306) <= layer4_outputs(7485);
    layer5_outputs(7307) <= (layer4_outputs(2702)) and (layer4_outputs(54));
    layer5_outputs(7308) <= not(layer4_outputs(1990));
    layer5_outputs(7309) <= layer4_outputs(2422);
    layer5_outputs(7310) <= not((layer4_outputs(361)) xor (layer4_outputs(5463)));
    layer5_outputs(7311) <= layer4_outputs(760);
    layer5_outputs(7312) <= layer4_outputs(7317);
    layer5_outputs(7313) <= not((layer4_outputs(691)) and (layer4_outputs(4487)));
    layer5_outputs(7314) <= not(layer4_outputs(607));
    layer5_outputs(7315) <= not((layer4_outputs(4528)) xor (layer4_outputs(388)));
    layer5_outputs(7316) <= layer4_outputs(382);
    layer5_outputs(7317) <= not((layer4_outputs(2286)) or (layer4_outputs(36)));
    layer5_outputs(7318) <= not((layer4_outputs(5997)) xor (layer4_outputs(1739)));
    layer5_outputs(7319) <= layer4_outputs(3176);
    layer5_outputs(7320) <= (layer4_outputs(3555)) and (layer4_outputs(7576));
    layer5_outputs(7321) <= not(layer4_outputs(3718));
    layer5_outputs(7322) <= layer4_outputs(1757);
    layer5_outputs(7323) <= not(layer4_outputs(6410)) or (layer4_outputs(2815));
    layer5_outputs(7324) <= layer4_outputs(2937);
    layer5_outputs(7325) <= not(layer4_outputs(4707));
    layer5_outputs(7326) <= not(layer4_outputs(1305));
    layer5_outputs(7327) <= not(layer4_outputs(6340)) or (layer4_outputs(3192));
    layer5_outputs(7328) <= not(layer4_outputs(4743));
    layer5_outputs(7329) <= not(layer4_outputs(4727));
    layer5_outputs(7330) <= not(layer4_outputs(2136));
    layer5_outputs(7331) <= (layer4_outputs(5933)) and not (layer4_outputs(1363));
    layer5_outputs(7332) <= layer4_outputs(5213);
    layer5_outputs(7333) <= not(layer4_outputs(4087));
    layer5_outputs(7334) <= not(layer4_outputs(7622));
    layer5_outputs(7335) <= not((layer4_outputs(6666)) or (layer4_outputs(5184)));
    layer5_outputs(7336) <= not(layer4_outputs(2437));
    layer5_outputs(7337) <= '1';
    layer5_outputs(7338) <= layer4_outputs(5967);
    layer5_outputs(7339) <= layer4_outputs(3720);
    layer5_outputs(7340) <= not(layer4_outputs(2886));
    layer5_outputs(7341) <= layer4_outputs(1200);
    layer5_outputs(7342) <= not((layer4_outputs(980)) or (layer4_outputs(5653)));
    layer5_outputs(7343) <= '0';
    layer5_outputs(7344) <= '1';
    layer5_outputs(7345) <= not(layer4_outputs(7515));
    layer5_outputs(7346) <= layer4_outputs(3307);
    layer5_outputs(7347) <= layer4_outputs(5882);
    layer5_outputs(7348) <= layer4_outputs(1902);
    layer5_outputs(7349) <= (layer4_outputs(6426)) and not (layer4_outputs(6352));
    layer5_outputs(7350) <= '1';
    layer5_outputs(7351) <= not(layer4_outputs(6357)) or (layer4_outputs(2838));
    layer5_outputs(7352) <= not(layer4_outputs(6524));
    layer5_outputs(7353) <= layer4_outputs(4772);
    layer5_outputs(7354) <= not((layer4_outputs(4952)) and (layer4_outputs(1453)));
    layer5_outputs(7355) <= (layer4_outputs(4187)) or (layer4_outputs(5980));
    layer5_outputs(7356) <= not((layer4_outputs(1236)) and (layer4_outputs(5959)));
    layer5_outputs(7357) <= not(layer4_outputs(6742));
    layer5_outputs(7358) <= layer4_outputs(3612);
    layer5_outputs(7359) <= (layer4_outputs(879)) xor (layer4_outputs(7265));
    layer5_outputs(7360) <= layer4_outputs(7042);
    layer5_outputs(7361) <= not(layer4_outputs(7622));
    layer5_outputs(7362) <= not(layer4_outputs(4006));
    layer5_outputs(7363) <= layer4_outputs(2965);
    layer5_outputs(7364) <= layer4_outputs(1709);
    layer5_outputs(7365) <= layer4_outputs(846);
    layer5_outputs(7366) <= not((layer4_outputs(5505)) xor (layer4_outputs(2619)));
    layer5_outputs(7367) <= not(layer4_outputs(6267));
    layer5_outputs(7368) <= not(layer4_outputs(6214));
    layer5_outputs(7369) <= not((layer4_outputs(7002)) xor (layer4_outputs(4709)));
    layer5_outputs(7370) <= not((layer4_outputs(5487)) or (layer4_outputs(6753)));
    layer5_outputs(7371) <= '0';
    layer5_outputs(7372) <= layer4_outputs(2979);
    layer5_outputs(7373) <= '0';
    layer5_outputs(7374) <= (layer4_outputs(5812)) and not (layer4_outputs(5626));
    layer5_outputs(7375) <= not(layer4_outputs(2247));
    layer5_outputs(7376) <= not(layer4_outputs(5567));
    layer5_outputs(7377) <= not(layer4_outputs(3533));
    layer5_outputs(7378) <= (layer4_outputs(636)) and not (layer4_outputs(303));
    layer5_outputs(7379) <= not(layer4_outputs(3600));
    layer5_outputs(7380) <= (layer4_outputs(1458)) xor (layer4_outputs(3469));
    layer5_outputs(7381) <= not((layer4_outputs(7652)) and (layer4_outputs(659)));
    layer5_outputs(7382) <= (layer4_outputs(3174)) and (layer4_outputs(5015));
    layer5_outputs(7383) <= layer4_outputs(1688);
    layer5_outputs(7384) <= not((layer4_outputs(7085)) or (layer4_outputs(4529)));
    layer5_outputs(7385) <= not(layer4_outputs(580));
    layer5_outputs(7386) <= layer4_outputs(632);
    layer5_outputs(7387) <= layer4_outputs(2126);
    layer5_outputs(7388) <= layer4_outputs(1720);
    layer5_outputs(7389) <= '0';
    layer5_outputs(7390) <= layer4_outputs(5790);
    layer5_outputs(7391) <= not(layer4_outputs(6907));
    layer5_outputs(7392) <= (layer4_outputs(3777)) and not (layer4_outputs(4556));
    layer5_outputs(7393) <= not(layer4_outputs(522)) or (layer4_outputs(5499));
    layer5_outputs(7394) <= layer4_outputs(4721);
    layer5_outputs(7395) <= (layer4_outputs(3601)) and (layer4_outputs(2955));
    layer5_outputs(7396) <= not((layer4_outputs(1793)) xor (layer4_outputs(5454)));
    layer5_outputs(7397) <= not((layer4_outputs(7439)) xor (layer4_outputs(217)));
    layer5_outputs(7398) <= (layer4_outputs(5909)) or (layer4_outputs(999));
    layer5_outputs(7399) <= not((layer4_outputs(139)) or (layer4_outputs(447)));
    layer5_outputs(7400) <= not(layer4_outputs(4422));
    layer5_outputs(7401) <= not(layer4_outputs(340));
    layer5_outputs(7402) <= (layer4_outputs(3037)) and (layer4_outputs(6255));
    layer5_outputs(7403) <= not(layer4_outputs(5548));
    layer5_outputs(7404) <= layer4_outputs(2097);
    layer5_outputs(7405) <= (layer4_outputs(6856)) and (layer4_outputs(3536));
    layer5_outputs(7406) <= layer4_outputs(5706);
    layer5_outputs(7407) <= not(layer4_outputs(427));
    layer5_outputs(7408) <= (layer4_outputs(3288)) xor (layer4_outputs(4540));
    layer5_outputs(7409) <= not(layer4_outputs(6201));
    layer5_outputs(7410) <= layer4_outputs(2244);
    layer5_outputs(7411) <= layer4_outputs(232);
    layer5_outputs(7412) <= (layer4_outputs(2432)) xor (layer4_outputs(2695));
    layer5_outputs(7413) <= (layer4_outputs(7070)) xor (layer4_outputs(5101));
    layer5_outputs(7414) <= not(layer4_outputs(300)) or (layer4_outputs(1718));
    layer5_outputs(7415) <= not(layer4_outputs(5364));
    layer5_outputs(7416) <= not(layer4_outputs(3198)) or (layer4_outputs(3863));
    layer5_outputs(7417) <= not(layer4_outputs(956));
    layer5_outputs(7418) <= layer4_outputs(3245);
    layer5_outputs(7419) <= not(layer4_outputs(1979));
    layer5_outputs(7420) <= (layer4_outputs(289)) and (layer4_outputs(4790));
    layer5_outputs(7421) <= '1';
    layer5_outputs(7422) <= not(layer4_outputs(3752));
    layer5_outputs(7423) <= layer4_outputs(3908);
    layer5_outputs(7424) <= not(layer4_outputs(6634));
    layer5_outputs(7425) <= not((layer4_outputs(6131)) or (layer4_outputs(4333)));
    layer5_outputs(7426) <= layer4_outputs(7157);
    layer5_outputs(7427) <= not(layer4_outputs(684));
    layer5_outputs(7428) <= not(layer4_outputs(7128));
    layer5_outputs(7429) <= not((layer4_outputs(739)) xor (layer4_outputs(3321)));
    layer5_outputs(7430) <= (layer4_outputs(2614)) and not (layer4_outputs(5820));
    layer5_outputs(7431) <= layer4_outputs(4328);
    layer5_outputs(7432) <= layer4_outputs(5627);
    layer5_outputs(7433) <= layer4_outputs(2711);
    layer5_outputs(7434) <= not(layer4_outputs(7097));
    layer5_outputs(7435) <= layer4_outputs(3402);
    layer5_outputs(7436) <= not(layer4_outputs(3245));
    layer5_outputs(7437) <= layer4_outputs(1503);
    layer5_outputs(7438) <= not((layer4_outputs(1213)) or (layer4_outputs(3049)));
    layer5_outputs(7439) <= (layer4_outputs(6007)) xor (layer4_outputs(5547));
    layer5_outputs(7440) <= not(layer4_outputs(761));
    layer5_outputs(7441) <= (layer4_outputs(1606)) xor (layer4_outputs(1434));
    layer5_outputs(7442) <= layer4_outputs(4106);
    layer5_outputs(7443) <= not(layer4_outputs(7400));
    layer5_outputs(7444) <= (layer4_outputs(6541)) xor (layer4_outputs(2497));
    layer5_outputs(7445) <= layer4_outputs(3511);
    layer5_outputs(7446) <= (layer4_outputs(2701)) and not (layer4_outputs(4755));
    layer5_outputs(7447) <= layer4_outputs(3582);
    layer5_outputs(7448) <= not(layer4_outputs(1100)) or (layer4_outputs(3350));
    layer5_outputs(7449) <= not((layer4_outputs(6053)) or (layer4_outputs(4016)));
    layer5_outputs(7450) <= not(layer4_outputs(6651)) or (layer4_outputs(5532));
    layer5_outputs(7451) <= (layer4_outputs(3542)) and not (layer4_outputs(5431));
    layer5_outputs(7452) <= (layer4_outputs(611)) and not (layer4_outputs(3726));
    layer5_outputs(7453) <= not(layer4_outputs(6019));
    layer5_outputs(7454) <= (layer4_outputs(6068)) and not (layer4_outputs(1936));
    layer5_outputs(7455) <= layer4_outputs(2812);
    layer5_outputs(7456) <= (layer4_outputs(1330)) and not (layer4_outputs(3694));
    layer5_outputs(7457) <= (layer4_outputs(6191)) xor (layer4_outputs(3703));
    layer5_outputs(7458) <= not((layer4_outputs(5186)) xor (layer4_outputs(1339)));
    layer5_outputs(7459) <= (layer4_outputs(2338)) and not (layer4_outputs(3788));
    layer5_outputs(7460) <= not(layer4_outputs(6346));
    layer5_outputs(7461) <= not((layer4_outputs(936)) or (layer4_outputs(3406)));
    layer5_outputs(7462) <= (layer4_outputs(1805)) xor (layer4_outputs(6823));
    layer5_outputs(7463) <= (layer4_outputs(4178)) and not (layer4_outputs(5932));
    layer5_outputs(7464) <= (layer4_outputs(5155)) and not (layer4_outputs(7481));
    layer5_outputs(7465) <= not(layer4_outputs(2945));
    layer5_outputs(7466) <= not(layer4_outputs(4246));
    layer5_outputs(7467) <= not(layer4_outputs(5689));
    layer5_outputs(7468) <= not((layer4_outputs(6994)) xor (layer4_outputs(5656)));
    layer5_outputs(7469) <= not(layer4_outputs(3860)) or (layer4_outputs(3543));
    layer5_outputs(7470) <= (layer4_outputs(6159)) xor (layer4_outputs(1340));
    layer5_outputs(7471) <= (layer4_outputs(5818)) or (layer4_outputs(450));
    layer5_outputs(7472) <= (layer4_outputs(6018)) xor (layer4_outputs(5733));
    layer5_outputs(7473) <= layer4_outputs(876);
    layer5_outputs(7474) <= not(layer4_outputs(630));
    layer5_outputs(7475) <= (layer4_outputs(5419)) or (layer4_outputs(2756));
    layer5_outputs(7476) <= (layer4_outputs(960)) xor (layer4_outputs(6175));
    layer5_outputs(7477) <= layer4_outputs(3098);
    layer5_outputs(7478) <= layer4_outputs(517);
    layer5_outputs(7479) <= (layer4_outputs(7332)) or (layer4_outputs(1272));
    layer5_outputs(7480) <= layer4_outputs(5614);
    layer5_outputs(7481) <= not((layer4_outputs(2546)) and (layer4_outputs(1222)));
    layer5_outputs(7482) <= not(layer4_outputs(7674));
    layer5_outputs(7483) <= not(layer4_outputs(4881));
    layer5_outputs(7484) <= (layer4_outputs(2287)) and not (layer4_outputs(7307));
    layer5_outputs(7485) <= layer4_outputs(6925);
    layer5_outputs(7486) <= layer4_outputs(3267);
    layer5_outputs(7487) <= (layer4_outputs(1056)) and not (layer4_outputs(3428));
    layer5_outputs(7488) <= not(layer4_outputs(938));
    layer5_outputs(7489) <= layer4_outputs(575);
    layer5_outputs(7490) <= layer4_outputs(6662);
    layer5_outputs(7491) <= not(layer4_outputs(626));
    layer5_outputs(7492) <= layer4_outputs(5307);
    layer5_outputs(7493) <= layer4_outputs(7309);
    layer5_outputs(7494) <= not((layer4_outputs(4311)) or (layer4_outputs(2952)));
    layer5_outputs(7495) <= not(layer4_outputs(1498));
    layer5_outputs(7496) <= layer4_outputs(1585);
    layer5_outputs(7497) <= '1';
    layer5_outputs(7498) <= (layer4_outputs(4591)) and (layer4_outputs(4718));
    layer5_outputs(7499) <= (layer4_outputs(1419)) and not (layer4_outputs(5958));
    layer5_outputs(7500) <= layer4_outputs(7324);
    layer5_outputs(7501) <= not(layer4_outputs(2922)) or (layer4_outputs(6911));
    layer5_outputs(7502) <= not(layer4_outputs(4247));
    layer5_outputs(7503) <= not(layer4_outputs(1998)) or (layer4_outputs(2720));
    layer5_outputs(7504) <= not(layer4_outputs(5119)) or (layer4_outputs(3239));
    layer5_outputs(7505) <= layer4_outputs(5790);
    layer5_outputs(7506) <= not(layer4_outputs(6567));
    layer5_outputs(7507) <= (layer4_outputs(5062)) and not (layer4_outputs(4489));
    layer5_outputs(7508) <= (layer4_outputs(6840)) xor (layer4_outputs(6116));
    layer5_outputs(7509) <= not(layer4_outputs(3084));
    layer5_outputs(7510) <= layer4_outputs(7445);
    layer5_outputs(7511) <= not(layer4_outputs(5495));
    layer5_outputs(7512) <= (layer4_outputs(5026)) and (layer4_outputs(486));
    layer5_outputs(7513) <= not(layer4_outputs(2847));
    layer5_outputs(7514) <= not(layer4_outputs(4631));
    layer5_outputs(7515) <= (layer4_outputs(6255)) and not (layer4_outputs(7207));
    layer5_outputs(7516) <= layer4_outputs(2349);
    layer5_outputs(7517) <= not(layer4_outputs(4948));
    layer5_outputs(7518) <= layer4_outputs(1326);
    layer5_outputs(7519) <= not((layer4_outputs(3297)) and (layer4_outputs(608)));
    layer5_outputs(7520) <= (layer4_outputs(534)) xor (layer4_outputs(5231));
    layer5_outputs(7521) <= not(layer4_outputs(6622));
    layer5_outputs(7522) <= layer4_outputs(225);
    layer5_outputs(7523) <= not(layer4_outputs(2519)) or (layer4_outputs(7391));
    layer5_outputs(7524) <= not((layer4_outputs(2709)) xor (layer4_outputs(2851)));
    layer5_outputs(7525) <= layer4_outputs(6381);
    layer5_outputs(7526) <= layer4_outputs(2515);
    layer5_outputs(7527) <= not(layer4_outputs(4125));
    layer5_outputs(7528) <= not(layer4_outputs(2537));
    layer5_outputs(7529) <= layer4_outputs(5813);
    layer5_outputs(7530) <= (layer4_outputs(3929)) and not (layer4_outputs(1300));
    layer5_outputs(7531) <= not(layer4_outputs(2981)) or (layer4_outputs(7669));
    layer5_outputs(7532) <= (layer4_outputs(4268)) and not (layer4_outputs(6036));
    layer5_outputs(7533) <= not((layer4_outputs(7423)) and (layer4_outputs(2625)));
    layer5_outputs(7534) <= not(layer4_outputs(7195)) or (layer4_outputs(5076));
    layer5_outputs(7535) <= layer4_outputs(5229);
    layer5_outputs(7536) <= layer4_outputs(6928);
    layer5_outputs(7537) <= (layer4_outputs(3464)) and not (layer4_outputs(4366));
    layer5_outputs(7538) <= not(layer4_outputs(3784));
    layer5_outputs(7539) <= (layer4_outputs(4741)) and (layer4_outputs(6114));
    layer5_outputs(7540) <= not(layer4_outputs(5946));
    layer5_outputs(7541) <= not((layer4_outputs(5623)) xor (layer4_outputs(7186)));
    layer5_outputs(7542) <= not(layer4_outputs(4658));
    layer5_outputs(7543) <= not((layer4_outputs(5452)) xor (layer4_outputs(5311)));
    layer5_outputs(7544) <= (layer4_outputs(2293)) or (layer4_outputs(1371));
    layer5_outputs(7545) <= layer4_outputs(6563);
    layer5_outputs(7546) <= not((layer4_outputs(5273)) and (layer4_outputs(5945)));
    layer5_outputs(7547) <= layer4_outputs(2087);
    layer5_outputs(7548) <= not(layer4_outputs(5753)) or (layer4_outputs(6551));
    layer5_outputs(7549) <= not(layer4_outputs(433));
    layer5_outputs(7550) <= layer4_outputs(1124);
    layer5_outputs(7551) <= (layer4_outputs(165)) and not (layer4_outputs(7263));
    layer5_outputs(7552) <= not(layer4_outputs(2859)) or (layer4_outputs(2551));
    layer5_outputs(7553) <= layer4_outputs(5795);
    layer5_outputs(7554) <= not(layer4_outputs(5707));
    layer5_outputs(7555) <= not(layer4_outputs(1377));
    layer5_outputs(7556) <= not(layer4_outputs(4731)) or (layer4_outputs(5518));
    layer5_outputs(7557) <= not(layer4_outputs(5596));
    layer5_outputs(7558) <= not((layer4_outputs(7648)) and (layer4_outputs(1757)));
    layer5_outputs(7559) <= '1';
    layer5_outputs(7560) <= layer4_outputs(2132);
    layer5_outputs(7561) <= (layer4_outputs(3164)) and not (layer4_outputs(3628));
    layer5_outputs(7562) <= not(layer4_outputs(2749)) or (layer4_outputs(4784));
    layer5_outputs(7563) <= layer4_outputs(2443);
    layer5_outputs(7564) <= not(layer4_outputs(7607)) or (layer4_outputs(7029));
    layer5_outputs(7565) <= (layer4_outputs(2725)) and not (layer4_outputs(429));
    layer5_outputs(7566) <= not(layer4_outputs(6918));
    layer5_outputs(7567) <= not(layer4_outputs(5050));
    layer5_outputs(7568) <= '0';
    layer5_outputs(7569) <= not(layer4_outputs(4246)) or (layer4_outputs(2640));
    layer5_outputs(7570) <= layer4_outputs(6321);
    layer5_outputs(7571) <= (layer4_outputs(2070)) or (layer4_outputs(587));
    layer5_outputs(7572) <= (layer4_outputs(494)) or (layer4_outputs(4518));
    layer5_outputs(7573) <= layer4_outputs(2448);
    layer5_outputs(7574) <= layer4_outputs(4744);
    layer5_outputs(7575) <= layer4_outputs(4799);
    layer5_outputs(7576) <= not((layer4_outputs(1313)) or (layer4_outputs(205)));
    layer5_outputs(7577) <= layer4_outputs(665);
    layer5_outputs(7578) <= not(layer4_outputs(6297)) or (layer4_outputs(6701));
    layer5_outputs(7579) <= (layer4_outputs(2304)) and not (layer4_outputs(7545));
    layer5_outputs(7580) <= (layer4_outputs(3002)) xor (layer4_outputs(5359));
    layer5_outputs(7581) <= not(layer4_outputs(3352)) or (layer4_outputs(3552));
    layer5_outputs(7582) <= not(layer4_outputs(5784)) or (layer4_outputs(3100));
    layer5_outputs(7583) <= (layer4_outputs(1999)) and (layer4_outputs(5514));
    layer5_outputs(7584) <= (layer4_outputs(2932)) and (layer4_outputs(2167));
    layer5_outputs(7585) <= not(layer4_outputs(3030));
    layer5_outputs(7586) <= layer4_outputs(3905);
    layer5_outputs(7587) <= layer4_outputs(5445);
    layer5_outputs(7588) <= not(layer4_outputs(3967));
    layer5_outputs(7589) <= not(layer4_outputs(3933));
    layer5_outputs(7590) <= not(layer4_outputs(3500));
    layer5_outputs(7591) <= layer4_outputs(1820);
    layer5_outputs(7592) <= (layer4_outputs(482)) and not (layer4_outputs(2558));
    layer5_outputs(7593) <= not((layer4_outputs(840)) or (layer4_outputs(4232)));
    layer5_outputs(7594) <= layer4_outputs(4233);
    layer5_outputs(7595) <= '1';
    layer5_outputs(7596) <= layer4_outputs(3497);
    layer5_outputs(7597) <= (layer4_outputs(512)) or (layer4_outputs(2873));
    layer5_outputs(7598) <= not(layer4_outputs(7448));
    layer5_outputs(7599) <= not(layer4_outputs(179));
    layer5_outputs(7600) <= not((layer4_outputs(7595)) xor (layer4_outputs(3878)));
    layer5_outputs(7601) <= not(layer4_outputs(1294));
    layer5_outputs(7602) <= not((layer4_outputs(7608)) xor (layer4_outputs(2362)));
    layer5_outputs(7603) <= layer4_outputs(967);
    layer5_outputs(7604) <= (layer4_outputs(4486)) xor (layer4_outputs(1750));
    layer5_outputs(7605) <= not(layer4_outputs(1080)) or (layer4_outputs(3383));
    layer5_outputs(7606) <= (layer4_outputs(7091)) and (layer4_outputs(2665));
    layer5_outputs(7607) <= (layer4_outputs(6603)) or (layer4_outputs(2210));
    layer5_outputs(7608) <= (layer4_outputs(6776)) and (layer4_outputs(2688));
    layer5_outputs(7609) <= not(layer4_outputs(364)) or (layer4_outputs(5571));
    layer5_outputs(7610) <= not(layer4_outputs(4231)) or (layer4_outputs(719));
    layer5_outputs(7611) <= not(layer4_outputs(4090));
    layer5_outputs(7612) <= not((layer4_outputs(7523)) or (layer4_outputs(3405)));
    layer5_outputs(7613) <= '1';
    layer5_outputs(7614) <= layer4_outputs(3084);
    layer5_outputs(7615) <= (layer4_outputs(2902)) or (layer4_outputs(7424));
    layer5_outputs(7616) <= not(layer4_outputs(2113));
    layer5_outputs(7617) <= not(layer4_outputs(146));
    layer5_outputs(7618) <= not(layer4_outputs(162));
    layer5_outputs(7619) <= (layer4_outputs(4393)) and not (layer4_outputs(5022));
    layer5_outputs(7620) <= (layer4_outputs(6563)) and not (layer4_outputs(5194));
    layer5_outputs(7621) <= (layer4_outputs(1002)) xor (layer4_outputs(1929));
    layer5_outputs(7622) <= not(layer4_outputs(2791)) or (layer4_outputs(6629));
    layer5_outputs(7623) <= not(layer4_outputs(4006));
    layer5_outputs(7624) <= not(layer4_outputs(2935)) or (layer4_outputs(15));
    layer5_outputs(7625) <= layer4_outputs(13);
    layer5_outputs(7626) <= not(layer4_outputs(2131));
    layer5_outputs(7627) <= layer4_outputs(5139);
    layer5_outputs(7628) <= not(layer4_outputs(1232));
    layer5_outputs(7629) <= layer4_outputs(3178);
    layer5_outputs(7630) <= (layer4_outputs(3447)) and (layer4_outputs(6750));
    layer5_outputs(7631) <= not(layer4_outputs(210));
    layer5_outputs(7632) <= '1';
    layer5_outputs(7633) <= not(layer4_outputs(1731));
    layer5_outputs(7634) <= not((layer4_outputs(1260)) or (layer4_outputs(6398)));
    layer5_outputs(7635) <= (layer4_outputs(5244)) and not (layer4_outputs(6052));
    layer5_outputs(7636) <= layer4_outputs(3021);
    layer5_outputs(7637) <= not((layer4_outputs(7138)) or (layer4_outputs(3617)));
    layer5_outputs(7638) <= layer4_outputs(5091);
    layer5_outputs(7639) <= layer4_outputs(2289);
    layer5_outputs(7640) <= not(layer4_outputs(2552));
    layer5_outputs(7641) <= not(layer4_outputs(5228));
    layer5_outputs(7642) <= not((layer4_outputs(2406)) xor (layer4_outputs(7256)));
    layer5_outputs(7643) <= not(layer4_outputs(6932));
    layer5_outputs(7644) <= (layer4_outputs(6835)) and not (layer4_outputs(297));
    layer5_outputs(7645) <= not(layer4_outputs(6809));
    layer5_outputs(7646) <= not(layer4_outputs(6328));
    layer5_outputs(7647) <= layer4_outputs(3249);
    layer5_outputs(7648) <= not(layer4_outputs(1534));
    layer5_outputs(7649) <= not(layer4_outputs(6730));
    layer5_outputs(7650) <= layer4_outputs(4749);
    layer5_outputs(7651) <= not(layer4_outputs(4493));
    layer5_outputs(7652) <= not(layer4_outputs(6314));
    layer5_outputs(7653) <= (layer4_outputs(3077)) xor (layer4_outputs(5240));
    layer5_outputs(7654) <= layer4_outputs(4569);
    layer5_outputs(7655) <= not((layer4_outputs(2125)) or (layer4_outputs(7301)));
    layer5_outputs(7656) <= not(layer4_outputs(5697));
    layer5_outputs(7657) <= not(layer4_outputs(3381));
    layer5_outputs(7658) <= not(layer4_outputs(2820));
    layer5_outputs(7659) <= layer4_outputs(5608);
    layer5_outputs(7660) <= layer4_outputs(6971);
    layer5_outputs(7661) <= not(layer4_outputs(161)) or (layer4_outputs(6362));
    layer5_outputs(7662) <= not((layer4_outputs(1440)) xor (layer4_outputs(1137)));
    layer5_outputs(7663) <= not(layer4_outputs(669));
    layer5_outputs(7664) <= not(layer4_outputs(2836));
    layer5_outputs(7665) <= layer4_outputs(7636);
    layer5_outputs(7666) <= not((layer4_outputs(5850)) and (layer4_outputs(6307)));
    layer5_outputs(7667) <= layer4_outputs(6848);
    layer5_outputs(7668) <= (layer4_outputs(2967)) and (layer4_outputs(7255));
    layer5_outputs(7669) <= layer4_outputs(758);
    layer5_outputs(7670) <= (layer4_outputs(5926)) xor (layer4_outputs(6209));
    layer5_outputs(7671) <= layer4_outputs(2012);
    layer5_outputs(7672) <= not(layer4_outputs(1447));
    layer5_outputs(7673) <= (layer4_outputs(3956)) and (layer4_outputs(4353));
    layer5_outputs(7674) <= not((layer4_outputs(6806)) and (layer4_outputs(7266)));
    layer5_outputs(7675) <= (layer4_outputs(7182)) and not (layer4_outputs(3651));
    layer5_outputs(7676) <= layer4_outputs(4580);
    layer5_outputs(7677) <= (layer4_outputs(7250)) and not (layer4_outputs(6961));
    layer5_outputs(7678) <= not(layer4_outputs(1321));
    layer5_outputs(7679) <= (layer4_outputs(2914)) or (layer4_outputs(3636));
    layer6_outputs(0) <= (layer5_outputs(3788)) and (layer5_outputs(1764));
    layer6_outputs(1) <= layer5_outputs(6707);
    layer6_outputs(2) <= not((layer5_outputs(7529)) or (layer5_outputs(69)));
    layer6_outputs(3) <= (layer5_outputs(4627)) xor (layer5_outputs(6624));
    layer6_outputs(4) <= layer5_outputs(4460);
    layer6_outputs(5) <= not((layer5_outputs(1995)) xor (layer5_outputs(4584)));
    layer6_outputs(6) <= (layer5_outputs(5834)) and not (layer5_outputs(5365));
    layer6_outputs(7) <= not(layer5_outputs(400));
    layer6_outputs(8) <= layer5_outputs(5841);
    layer6_outputs(9) <= not(layer5_outputs(3630));
    layer6_outputs(10) <= not((layer5_outputs(4673)) xor (layer5_outputs(406)));
    layer6_outputs(11) <= (layer5_outputs(7523)) and not (layer5_outputs(3692));
    layer6_outputs(12) <= (layer5_outputs(6768)) or (layer5_outputs(6716));
    layer6_outputs(13) <= not(layer5_outputs(3895)) or (layer5_outputs(5342));
    layer6_outputs(14) <= not((layer5_outputs(102)) or (layer5_outputs(71)));
    layer6_outputs(15) <= not(layer5_outputs(4769));
    layer6_outputs(16) <= not(layer5_outputs(7450));
    layer6_outputs(17) <= (layer5_outputs(4387)) or (layer5_outputs(6730));
    layer6_outputs(18) <= (layer5_outputs(547)) and not (layer5_outputs(7316));
    layer6_outputs(19) <= not((layer5_outputs(5094)) xor (layer5_outputs(7221)));
    layer6_outputs(20) <= not(layer5_outputs(5226));
    layer6_outputs(21) <= not((layer5_outputs(3789)) xor (layer5_outputs(5533)));
    layer6_outputs(22) <= '1';
    layer6_outputs(23) <= (layer5_outputs(5242)) xor (layer5_outputs(2));
    layer6_outputs(24) <= layer5_outputs(998);
    layer6_outputs(25) <= not(layer5_outputs(3398));
    layer6_outputs(26) <= (layer5_outputs(6221)) or (layer5_outputs(920));
    layer6_outputs(27) <= not((layer5_outputs(4977)) and (layer5_outputs(7166)));
    layer6_outputs(28) <= '0';
    layer6_outputs(29) <= layer5_outputs(1630);
    layer6_outputs(30) <= not((layer5_outputs(5298)) or (layer5_outputs(943)));
    layer6_outputs(31) <= (layer5_outputs(6400)) and not (layer5_outputs(4849));
    layer6_outputs(32) <= layer5_outputs(3327);
    layer6_outputs(33) <= (layer5_outputs(1991)) or (layer5_outputs(7487));
    layer6_outputs(34) <= not(layer5_outputs(910));
    layer6_outputs(35) <= not(layer5_outputs(1997));
    layer6_outputs(36) <= not(layer5_outputs(5178));
    layer6_outputs(37) <= layer5_outputs(4387);
    layer6_outputs(38) <= not(layer5_outputs(5299)) or (layer5_outputs(5483));
    layer6_outputs(39) <= not(layer5_outputs(3594)) or (layer5_outputs(6287));
    layer6_outputs(40) <= (layer5_outputs(7382)) xor (layer5_outputs(2868));
    layer6_outputs(41) <= not((layer5_outputs(5922)) xor (layer5_outputs(623)));
    layer6_outputs(42) <= layer5_outputs(3892);
    layer6_outputs(43) <= (layer5_outputs(5407)) xor (layer5_outputs(2442));
    layer6_outputs(44) <= (layer5_outputs(1140)) and (layer5_outputs(6437));
    layer6_outputs(45) <= layer5_outputs(6744);
    layer6_outputs(46) <= not(layer5_outputs(1497));
    layer6_outputs(47) <= not(layer5_outputs(5142));
    layer6_outputs(48) <= not((layer5_outputs(5434)) or (layer5_outputs(694)));
    layer6_outputs(49) <= (layer5_outputs(2716)) and not (layer5_outputs(3520));
    layer6_outputs(50) <= not((layer5_outputs(7601)) or (layer5_outputs(6380)));
    layer6_outputs(51) <= layer5_outputs(2016);
    layer6_outputs(52) <= not(layer5_outputs(3274));
    layer6_outputs(53) <= (layer5_outputs(1951)) and not (layer5_outputs(4253));
    layer6_outputs(54) <= layer5_outputs(4160);
    layer6_outputs(55) <= not(layer5_outputs(2263));
    layer6_outputs(56) <= not((layer5_outputs(4068)) xor (layer5_outputs(2740)));
    layer6_outputs(57) <= layer5_outputs(7258);
    layer6_outputs(58) <= (layer5_outputs(3627)) and (layer5_outputs(3047));
    layer6_outputs(59) <= layer5_outputs(3309);
    layer6_outputs(60) <= not(layer5_outputs(2465));
    layer6_outputs(61) <= not((layer5_outputs(668)) xor (layer5_outputs(5187)));
    layer6_outputs(62) <= layer5_outputs(359);
    layer6_outputs(63) <= layer5_outputs(1402);
    layer6_outputs(64) <= not((layer5_outputs(5380)) or (layer5_outputs(4529)));
    layer6_outputs(65) <= (layer5_outputs(3322)) and not (layer5_outputs(3557));
    layer6_outputs(66) <= not(layer5_outputs(4572));
    layer6_outputs(67) <= not(layer5_outputs(6912));
    layer6_outputs(68) <= not(layer5_outputs(505));
    layer6_outputs(69) <= layer5_outputs(6992);
    layer6_outputs(70) <= not((layer5_outputs(2969)) xor (layer5_outputs(7313)));
    layer6_outputs(71) <= not(layer5_outputs(5983));
    layer6_outputs(72) <= layer5_outputs(2397);
    layer6_outputs(73) <= layer5_outputs(1025);
    layer6_outputs(74) <= layer5_outputs(1797);
    layer6_outputs(75) <= not((layer5_outputs(4899)) and (layer5_outputs(3182)));
    layer6_outputs(76) <= layer5_outputs(604);
    layer6_outputs(77) <= '0';
    layer6_outputs(78) <= (layer5_outputs(4593)) and not (layer5_outputs(4781));
    layer6_outputs(79) <= (layer5_outputs(271)) xor (layer5_outputs(5966));
    layer6_outputs(80) <= not(layer5_outputs(1737));
    layer6_outputs(81) <= not(layer5_outputs(3369));
    layer6_outputs(82) <= not(layer5_outputs(630));
    layer6_outputs(83) <= not(layer5_outputs(5654)) or (layer5_outputs(6331));
    layer6_outputs(84) <= not(layer5_outputs(5598));
    layer6_outputs(85) <= not(layer5_outputs(2014));
    layer6_outputs(86) <= not(layer5_outputs(2784)) or (layer5_outputs(964));
    layer6_outputs(87) <= layer5_outputs(7365);
    layer6_outputs(88) <= not(layer5_outputs(3488)) or (layer5_outputs(2060));
    layer6_outputs(89) <= not(layer5_outputs(2494));
    layer6_outputs(90) <= not(layer5_outputs(5476)) or (layer5_outputs(3654));
    layer6_outputs(91) <= not(layer5_outputs(4907));
    layer6_outputs(92) <= layer5_outputs(3246);
    layer6_outputs(93) <= (layer5_outputs(4174)) xor (layer5_outputs(6022));
    layer6_outputs(94) <= (layer5_outputs(1247)) and not (layer5_outputs(6004));
    layer6_outputs(95) <= not(layer5_outputs(616));
    layer6_outputs(96) <= not(layer5_outputs(1494));
    layer6_outputs(97) <= (layer5_outputs(95)) xor (layer5_outputs(4369));
    layer6_outputs(98) <= layer5_outputs(4325);
    layer6_outputs(99) <= not(layer5_outputs(1650)) or (layer5_outputs(2793));
    layer6_outputs(100) <= (layer5_outputs(1791)) and (layer5_outputs(5772));
    layer6_outputs(101) <= (layer5_outputs(7267)) and not (layer5_outputs(377));
    layer6_outputs(102) <= layer5_outputs(5732);
    layer6_outputs(103) <= layer5_outputs(2617);
    layer6_outputs(104) <= not(layer5_outputs(953));
    layer6_outputs(105) <= not(layer5_outputs(5702)) or (layer5_outputs(4958));
    layer6_outputs(106) <= not(layer5_outputs(4414)) or (layer5_outputs(5948));
    layer6_outputs(107) <= (layer5_outputs(875)) or (layer5_outputs(7286));
    layer6_outputs(108) <= not(layer5_outputs(3072)) or (layer5_outputs(7013));
    layer6_outputs(109) <= not(layer5_outputs(4635));
    layer6_outputs(110) <= (layer5_outputs(6636)) or (layer5_outputs(5968));
    layer6_outputs(111) <= not((layer5_outputs(1567)) and (layer5_outputs(2410)));
    layer6_outputs(112) <= layer5_outputs(3353);
    layer6_outputs(113) <= layer5_outputs(2968);
    layer6_outputs(114) <= (layer5_outputs(3956)) and not (layer5_outputs(7265));
    layer6_outputs(115) <= layer5_outputs(6684);
    layer6_outputs(116) <= (layer5_outputs(1641)) or (layer5_outputs(1366));
    layer6_outputs(117) <= layer5_outputs(5552);
    layer6_outputs(118) <= not(layer5_outputs(5048)) or (layer5_outputs(1807));
    layer6_outputs(119) <= not(layer5_outputs(3835)) or (layer5_outputs(5257));
    layer6_outputs(120) <= (layer5_outputs(3150)) and (layer5_outputs(3500));
    layer6_outputs(121) <= layer5_outputs(6554);
    layer6_outputs(122) <= not(layer5_outputs(2002));
    layer6_outputs(123) <= not(layer5_outputs(2306));
    layer6_outputs(124) <= layer5_outputs(7528);
    layer6_outputs(125) <= layer5_outputs(219);
    layer6_outputs(126) <= not((layer5_outputs(7134)) xor (layer5_outputs(7187)));
    layer6_outputs(127) <= (layer5_outputs(190)) xor (layer5_outputs(838));
    layer6_outputs(128) <= not(layer5_outputs(342));
    layer6_outputs(129) <= not(layer5_outputs(7311));
    layer6_outputs(130) <= layer5_outputs(1830);
    layer6_outputs(131) <= not(layer5_outputs(7130));
    layer6_outputs(132) <= layer5_outputs(6715);
    layer6_outputs(133) <= not(layer5_outputs(3904));
    layer6_outputs(134) <= (layer5_outputs(6041)) and not (layer5_outputs(2331));
    layer6_outputs(135) <= not(layer5_outputs(2288));
    layer6_outputs(136) <= '0';
    layer6_outputs(137) <= not(layer5_outputs(6602));
    layer6_outputs(138) <= (layer5_outputs(7155)) or (layer5_outputs(5212));
    layer6_outputs(139) <= layer5_outputs(646);
    layer6_outputs(140) <= not((layer5_outputs(467)) xor (layer5_outputs(7157)));
    layer6_outputs(141) <= (layer5_outputs(6088)) xor (layer5_outputs(6266));
    layer6_outputs(142) <= not(layer5_outputs(557));
    layer6_outputs(143) <= layer5_outputs(1478);
    layer6_outputs(144) <= not(layer5_outputs(7448));
    layer6_outputs(145) <= (layer5_outputs(3265)) xor (layer5_outputs(110));
    layer6_outputs(146) <= (layer5_outputs(6796)) or (layer5_outputs(3493));
    layer6_outputs(147) <= layer5_outputs(1093);
    layer6_outputs(148) <= layer5_outputs(3718);
    layer6_outputs(149) <= (layer5_outputs(3040)) xor (layer5_outputs(2585));
    layer6_outputs(150) <= not(layer5_outputs(3871));
    layer6_outputs(151) <= not((layer5_outputs(2074)) or (layer5_outputs(1874)));
    layer6_outputs(152) <= not(layer5_outputs(7219)) or (layer5_outputs(1279));
    layer6_outputs(153) <= not(layer5_outputs(4470));
    layer6_outputs(154) <= layer5_outputs(6713);
    layer6_outputs(155) <= not(layer5_outputs(3484));
    layer6_outputs(156) <= (layer5_outputs(3223)) and not (layer5_outputs(1155));
    layer6_outputs(157) <= layer5_outputs(2006);
    layer6_outputs(158) <= layer5_outputs(5912);
    layer6_outputs(159) <= not((layer5_outputs(6846)) xor (layer5_outputs(2100)));
    layer6_outputs(160) <= not((layer5_outputs(2649)) and (layer5_outputs(5395)));
    layer6_outputs(161) <= not(layer5_outputs(122));
    layer6_outputs(162) <= layer5_outputs(7380);
    layer6_outputs(163) <= not(layer5_outputs(3045));
    layer6_outputs(164) <= not(layer5_outputs(3366));
    layer6_outputs(165) <= (layer5_outputs(515)) and not (layer5_outputs(2833));
    layer6_outputs(166) <= not((layer5_outputs(3080)) or (layer5_outputs(1448)));
    layer6_outputs(167) <= (layer5_outputs(2059)) and not (layer5_outputs(529));
    layer6_outputs(168) <= not((layer5_outputs(414)) xor (layer5_outputs(6311)));
    layer6_outputs(169) <= (layer5_outputs(1241)) and (layer5_outputs(5897));
    layer6_outputs(170) <= not(layer5_outputs(5091)) or (layer5_outputs(5206));
    layer6_outputs(171) <= not((layer5_outputs(7162)) xor (layer5_outputs(1695)));
    layer6_outputs(172) <= not(layer5_outputs(908)) or (layer5_outputs(1955));
    layer6_outputs(173) <= layer5_outputs(1749);
    layer6_outputs(174) <= not(layer5_outputs(1771));
    layer6_outputs(175) <= (layer5_outputs(5221)) and not (layer5_outputs(6516));
    layer6_outputs(176) <= (layer5_outputs(5384)) and not (layer5_outputs(3393));
    layer6_outputs(177) <= layer5_outputs(4894);
    layer6_outputs(178) <= not(layer5_outputs(5038));
    layer6_outputs(179) <= not(layer5_outputs(201)) or (layer5_outputs(2521));
    layer6_outputs(180) <= (layer5_outputs(4662)) and not (layer5_outputs(3593));
    layer6_outputs(181) <= layer5_outputs(7436);
    layer6_outputs(182) <= not(layer5_outputs(1669));
    layer6_outputs(183) <= not((layer5_outputs(6078)) xor (layer5_outputs(7536)));
    layer6_outputs(184) <= not(layer5_outputs(2870));
    layer6_outputs(185) <= layer5_outputs(3332);
    layer6_outputs(186) <= (layer5_outputs(3433)) and not (layer5_outputs(3786));
    layer6_outputs(187) <= layer5_outputs(7546);
    layer6_outputs(188) <= not(layer5_outputs(2168));
    layer6_outputs(189) <= not(layer5_outputs(5387));
    layer6_outputs(190) <= (layer5_outputs(6628)) or (layer5_outputs(1153));
    layer6_outputs(191) <= (layer5_outputs(6727)) and (layer5_outputs(5747));
    layer6_outputs(192) <= not(layer5_outputs(4512));
    layer6_outputs(193) <= (layer5_outputs(6896)) and not (layer5_outputs(3733));
    layer6_outputs(194) <= not((layer5_outputs(3955)) and (layer5_outputs(828)));
    layer6_outputs(195) <= not(layer5_outputs(5977));
    layer6_outputs(196) <= (layer5_outputs(3913)) xor (layer5_outputs(4537));
    layer6_outputs(197) <= (layer5_outputs(1781)) and not (layer5_outputs(2367));
    layer6_outputs(198) <= layer5_outputs(7562);
    layer6_outputs(199) <= (layer5_outputs(7169)) xor (layer5_outputs(1056));
    layer6_outputs(200) <= layer5_outputs(4612);
    layer6_outputs(201) <= layer5_outputs(176);
    layer6_outputs(202) <= layer5_outputs(854);
    layer6_outputs(203) <= (layer5_outputs(3154)) xor (layer5_outputs(6624));
    layer6_outputs(204) <= not((layer5_outputs(2871)) and (layer5_outputs(4454)));
    layer6_outputs(205) <= not(layer5_outputs(4359)) or (layer5_outputs(7173));
    layer6_outputs(206) <= (layer5_outputs(6050)) xor (layer5_outputs(1834));
    layer6_outputs(207) <= layer5_outputs(926);
    layer6_outputs(208) <= not(layer5_outputs(5720));
    layer6_outputs(209) <= layer5_outputs(891);
    layer6_outputs(210) <= not(layer5_outputs(6753));
    layer6_outputs(211) <= layer5_outputs(4970);
    layer6_outputs(212) <= not((layer5_outputs(2151)) xor (layer5_outputs(4009)));
    layer6_outputs(213) <= not(layer5_outputs(3009));
    layer6_outputs(214) <= (layer5_outputs(2515)) or (layer5_outputs(5909));
    layer6_outputs(215) <= (layer5_outputs(3830)) and (layer5_outputs(1064));
    layer6_outputs(216) <= (layer5_outputs(2629)) and not (layer5_outputs(840));
    layer6_outputs(217) <= not(layer5_outputs(178));
    layer6_outputs(218) <= (layer5_outputs(6628)) and not (layer5_outputs(7114));
    layer6_outputs(219) <= not(layer5_outputs(778));
    layer6_outputs(220) <= not(layer5_outputs(2235));
    layer6_outputs(221) <= (layer5_outputs(4499)) and (layer5_outputs(2871));
    layer6_outputs(222) <= not(layer5_outputs(4777));
    layer6_outputs(223) <= layer5_outputs(7558);
    layer6_outputs(224) <= not((layer5_outputs(5702)) and (layer5_outputs(4424)));
    layer6_outputs(225) <= (layer5_outputs(3477)) and not (layer5_outputs(2945));
    layer6_outputs(226) <= layer5_outputs(848);
    layer6_outputs(227) <= not(layer5_outputs(7537));
    layer6_outputs(228) <= layer5_outputs(4263);
    layer6_outputs(229) <= not(layer5_outputs(885));
    layer6_outputs(230) <= not((layer5_outputs(7660)) xor (layer5_outputs(3273)));
    layer6_outputs(231) <= (layer5_outputs(6284)) and (layer5_outputs(4337));
    layer6_outputs(232) <= not(layer5_outputs(1909));
    layer6_outputs(233) <= not((layer5_outputs(2395)) and (layer5_outputs(800)));
    layer6_outputs(234) <= (layer5_outputs(7055)) and (layer5_outputs(3179));
    layer6_outputs(235) <= layer5_outputs(4201);
    layer6_outputs(236) <= not((layer5_outputs(2570)) and (layer5_outputs(6431)));
    layer6_outputs(237) <= not(layer5_outputs(4816));
    layer6_outputs(238) <= (layer5_outputs(3565)) and not (layer5_outputs(3868));
    layer6_outputs(239) <= not((layer5_outputs(7099)) xor (layer5_outputs(3790)));
    layer6_outputs(240) <= not(layer5_outputs(6577));
    layer6_outputs(241) <= (layer5_outputs(2084)) or (layer5_outputs(7500));
    layer6_outputs(242) <= not((layer5_outputs(4639)) or (layer5_outputs(1060)));
    layer6_outputs(243) <= not((layer5_outputs(5931)) or (layer5_outputs(6660)));
    layer6_outputs(244) <= layer5_outputs(7319);
    layer6_outputs(245) <= not(layer5_outputs(7252));
    layer6_outputs(246) <= not(layer5_outputs(7125));
    layer6_outputs(247) <= not(layer5_outputs(6279));
    layer6_outputs(248) <= (layer5_outputs(7521)) or (layer5_outputs(1384));
    layer6_outputs(249) <= (layer5_outputs(5173)) and not (layer5_outputs(1015));
    layer6_outputs(250) <= not(layer5_outputs(5578)) or (layer5_outputs(7313));
    layer6_outputs(251) <= (layer5_outputs(6378)) and (layer5_outputs(761));
    layer6_outputs(252) <= (layer5_outputs(2939)) and not (layer5_outputs(7579));
    layer6_outputs(253) <= layer5_outputs(1369);
    layer6_outputs(254) <= not((layer5_outputs(2424)) xor (layer5_outputs(2076)));
    layer6_outputs(255) <= layer5_outputs(4775);
    layer6_outputs(256) <= not((layer5_outputs(7087)) and (layer5_outputs(6192)));
    layer6_outputs(257) <= not(layer5_outputs(2515)) or (layer5_outputs(5156));
    layer6_outputs(258) <= not(layer5_outputs(6867)) or (layer5_outputs(5608));
    layer6_outputs(259) <= layer5_outputs(3642);
    layer6_outputs(260) <= not(layer5_outputs(1924)) or (layer5_outputs(6320));
    layer6_outputs(261) <= not(layer5_outputs(6804));
    layer6_outputs(262) <= not(layer5_outputs(3073));
    layer6_outputs(263) <= not(layer5_outputs(6012)) or (layer5_outputs(687));
    layer6_outputs(264) <= (layer5_outputs(6973)) or (layer5_outputs(4883));
    layer6_outputs(265) <= layer5_outputs(2277);
    layer6_outputs(266) <= not(layer5_outputs(4123)) or (layer5_outputs(6470));
    layer6_outputs(267) <= not(layer5_outputs(2746));
    layer6_outputs(268) <= (layer5_outputs(7254)) xor (layer5_outputs(928));
    layer6_outputs(269) <= not(layer5_outputs(1573)) or (layer5_outputs(605));
    layer6_outputs(270) <= not(layer5_outputs(573));
    layer6_outputs(271) <= layer5_outputs(1826);
    layer6_outputs(272) <= not(layer5_outputs(2640));
    layer6_outputs(273) <= not(layer5_outputs(6659));
    layer6_outputs(274) <= (layer5_outputs(3562)) or (layer5_outputs(3633));
    layer6_outputs(275) <= not(layer5_outputs(1866));
    layer6_outputs(276) <= (layer5_outputs(1574)) or (layer5_outputs(2773));
    layer6_outputs(277) <= not(layer5_outputs(6934));
    layer6_outputs(278) <= not(layer5_outputs(7628));
    layer6_outputs(279) <= not(layer5_outputs(1526)) or (layer5_outputs(6953));
    layer6_outputs(280) <= not(layer5_outputs(7189));
    layer6_outputs(281) <= not(layer5_outputs(1965));
    layer6_outputs(282) <= not(layer5_outputs(5159)) or (layer5_outputs(1226));
    layer6_outputs(283) <= not(layer5_outputs(7624)) or (layer5_outputs(1441));
    layer6_outputs(284) <= (layer5_outputs(1671)) or (layer5_outputs(1487));
    layer6_outputs(285) <= (layer5_outputs(4)) and not (layer5_outputs(2992));
    layer6_outputs(286) <= not(layer5_outputs(7020));
    layer6_outputs(287) <= (layer5_outputs(4542)) and (layer5_outputs(3829));
    layer6_outputs(288) <= not(layer5_outputs(2451)) or (layer5_outputs(1946));
    layer6_outputs(289) <= (layer5_outputs(483)) and not (layer5_outputs(1857));
    layer6_outputs(290) <= not((layer5_outputs(5189)) and (layer5_outputs(1721)));
    layer6_outputs(291) <= layer5_outputs(4759);
    layer6_outputs(292) <= layer5_outputs(3637);
    layer6_outputs(293) <= (layer5_outputs(3836)) and not (layer5_outputs(3964));
    layer6_outputs(294) <= layer5_outputs(7653);
    layer6_outputs(295) <= (layer5_outputs(6423)) and not (layer5_outputs(4630));
    layer6_outputs(296) <= not(layer5_outputs(3624));
    layer6_outputs(297) <= not((layer5_outputs(5363)) xor (layer5_outputs(5599)));
    layer6_outputs(298) <= not(layer5_outputs(19)) or (layer5_outputs(7435));
    layer6_outputs(299) <= layer5_outputs(2149);
    layer6_outputs(300) <= not(layer5_outputs(965));
    layer6_outputs(301) <= not(layer5_outputs(4349));
    layer6_outputs(302) <= layer5_outputs(4755);
    layer6_outputs(303) <= not(layer5_outputs(4818));
    layer6_outputs(304) <= not(layer5_outputs(6598)) or (layer5_outputs(6347));
    layer6_outputs(305) <= (layer5_outputs(4242)) xor (layer5_outputs(1283));
    layer6_outputs(306) <= (layer5_outputs(6402)) or (layer5_outputs(6785));
    layer6_outputs(307) <= (layer5_outputs(2627)) xor (layer5_outputs(888));
    layer6_outputs(308) <= not((layer5_outputs(2405)) xor (layer5_outputs(1003)));
    layer6_outputs(309) <= layer5_outputs(2003);
    layer6_outputs(310) <= layer5_outputs(4211);
    layer6_outputs(311) <= (layer5_outputs(214)) xor (layer5_outputs(5111));
    layer6_outputs(312) <= (layer5_outputs(1964)) xor (layer5_outputs(266));
    layer6_outputs(313) <= not((layer5_outputs(6379)) or (layer5_outputs(6539)));
    layer6_outputs(314) <= not((layer5_outputs(465)) or (layer5_outputs(6538)));
    layer6_outputs(315) <= not(layer5_outputs(6409));
    layer6_outputs(316) <= not((layer5_outputs(6498)) xor (layer5_outputs(1774)));
    layer6_outputs(317) <= not((layer5_outputs(5759)) and (layer5_outputs(1794)));
    layer6_outputs(318) <= '1';
    layer6_outputs(319) <= (layer5_outputs(3842)) and not (layer5_outputs(1909));
    layer6_outputs(320) <= not((layer5_outputs(6180)) or (layer5_outputs(2601)));
    layer6_outputs(321) <= layer5_outputs(897);
    layer6_outputs(322) <= layer5_outputs(4135);
    layer6_outputs(323) <= not(layer5_outputs(4213));
    layer6_outputs(324) <= (layer5_outputs(3005)) or (layer5_outputs(360));
    layer6_outputs(325) <= not(layer5_outputs(5366)) or (layer5_outputs(4083));
    layer6_outputs(326) <= layer5_outputs(6685);
    layer6_outputs(327) <= not((layer5_outputs(5806)) and (layer5_outputs(92)));
    layer6_outputs(328) <= (layer5_outputs(6738)) and not (layer5_outputs(3649));
    layer6_outputs(329) <= (layer5_outputs(7198)) and (layer5_outputs(4478));
    layer6_outputs(330) <= layer5_outputs(5881);
    layer6_outputs(331) <= (layer5_outputs(3638)) xor (layer5_outputs(6616));
    layer6_outputs(332) <= (layer5_outputs(2639)) and not (layer5_outputs(6799));
    layer6_outputs(333) <= layer5_outputs(2244);
    layer6_outputs(334) <= not(layer5_outputs(2308));
    layer6_outputs(335) <= layer5_outputs(2174);
    layer6_outputs(336) <= layer5_outputs(2296);
    layer6_outputs(337) <= (layer5_outputs(5544)) or (layer5_outputs(1660));
    layer6_outputs(338) <= (layer5_outputs(4491)) xor (layer5_outputs(5237));
    layer6_outputs(339) <= not(layer5_outputs(4333));
    layer6_outputs(340) <= not((layer5_outputs(4677)) xor (layer5_outputs(2624)));
    layer6_outputs(341) <= not(layer5_outputs(512)) or (layer5_outputs(5383));
    layer6_outputs(342) <= (layer5_outputs(4888)) xor (layer5_outputs(5680));
    layer6_outputs(343) <= (layer5_outputs(6466)) or (layer5_outputs(4029));
    layer6_outputs(344) <= not((layer5_outputs(160)) and (layer5_outputs(1467)));
    layer6_outputs(345) <= (layer5_outputs(465)) xor (layer5_outputs(5071));
    layer6_outputs(346) <= not(layer5_outputs(4502)) or (layer5_outputs(5288));
    layer6_outputs(347) <= (layer5_outputs(517)) xor (layer5_outputs(1248));
    layer6_outputs(348) <= not((layer5_outputs(970)) xor (layer5_outputs(3190)));
    layer6_outputs(349) <= layer5_outputs(4463);
    layer6_outputs(350) <= not(layer5_outputs(2116));
    layer6_outputs(351) <= not(layer5_outputs(3164));
    layer6_outputs(352) <= (layer5_outputs(7061)) and not (layer5_outputs(2756));
    layer6_outputs(353) <= not((layer5_outputs(7371)) and (layer5_outputs(3142)));
    layer6_outputs(354) <= layer5_outputs(3137);
    layer6_outputs(355) <= (layer5_outputs(2827)) and not (layer5_outputs(2423));
    layer6_outputs(356) <= not(layer5_outputs(2821));
    layer6_outputs(357) <= (layer5_outputs(2279)) and not (layer5_outputs(2430));
    layer6_outputs(358) <= (layer5_outputs(7221)) xor (layer5_outputs(7068));
    layer6_outputs(359) <= not((layer5_outputs(2616)) xor (layer5_outputs(2535)));
    layer6_outputs(360) <= (layer5_outputs(732)) and not (layer5_outputs(5893));
    layer6_outputs(361) <= (layer5_outputs(6545)) or (layer5_outputs(6481));
    layer6_outputs(362) <= not((layer5_outputs(3714)) or (layer5_outputs(3881)));
    layer6_outputs(363) <= not(layer5_outputs(7214)) or (layer5_outputs(5808));
    layer6_outputs(364) <= layer5_outputs(2825);
    layer6_outputs(365) <= layer5_outputs(4319);
    layer6_outputs(366) <= (layer5_outputs(647)) or (layer5_outputs(6868));
    layer6_outputs(367) <= not(layer5_outputs(4332));
    layer6_outputs(368) <= not(layer5_outputs(6113)) or (layer5_outputs(371));
    layer6_outputs(369) <= layer5_outputs(4583);
    layer6_outputs(370) <= layer5_outputs(2889);
    layer6_outputs(371) <= not(layer5_outputs(1618));
    layer6_outputs(372) <= layer5_outputs(4294);
    layer6_outputs(373) <= (layer5_outputs(7093)) and (layer5_outputs(4035));
    layer6_outputs(374) <= layer5_outputs(993);
    layer6_outputs(375) <= not(layer5_outputs(3350));
    layer6_outputs(376) <= layer5_outputs(2210);
    layer6_outputs(377) <= (layer5_outputs(3699)) xor (layer5_outputs(7424));
    layer6_outputs(378) <= layer5_outputs(6513);
    layer6_outputs(379) <= not((layer5_outputs(3557)) xor (layer5_outputs(250)));
    layer6_outputs(380) <= (layer5_outputs(3134)) and not (layer5_outputs(2940));
    layer6_outputs(381) <= (layer5_outputs(1988)) or (layer5_outputs(2493));
    layer6_outputs(382) <= not(layer5_outputs(4928));
    layer6_outputs(383) <= layer5_outputs(2808);
    layer6_outputs(384) <= (layer5_outputs(6146)) xor (layer5_outputs(6484));
    layer6_outputs(385) <= (layer5_outputs(6194)) xor (layer5_outputs(1994));
    layer6_outputs(386) <= layer5_outputs(1607);
    layer6_outputs(387) <= (layer5_outputs(6313)) xor (layer5_outputs(4366));
    layer6_outputs(388) <= not(layer5_outputs(4391));
    layer6_outputs(389) <= (layer5_outputs(6781)) xor (layer5_outputs(6900));
    layer6_outputs(390) <= (layer5_outputs(6448)) and not (layer5_outputs(2497));
    layer6_outputs(391) <= layer5_outputs(3277);
    layer6_outputs(392) <= not(layer5_outputs(653)) or (layer5_outputs(6828));
    layer6_outputs(393) <= (layer5_outputs(5541)) xor (layer5_outputs(1868));
    layer6_outputs(394) <= not(layer5_outputs(5215)) or (layer5_outputs(2956));
    layer6_outputs(395) <= layer5_outputs(6325);
    layer6_outputs(396) <= layer5_outputs(4106);
    layer6_outputs(397) <= (layer5_outputs(585)) or (layer5_outputs(5754));
    layer6_outputs(398) <= not(layer5_outputs(3684)) or (layer5_outputs(129));
    layer6_outputs(399) <= not(layer5_outputs(867));
    layer6_outputs(400) <= layer5_outputs(1385);
    layer6_outputs(401) <= not(layer5_outputs(2303));
    layer6_outputs(402) <= not(layer5_outputs(1628));
    layer6_outputs(403) <= not(layer5_outputs(2800));
    layer6_outputs(404) <= not(layer5_outputs(5277));
    layer6_outputs(405) <= not((layer5_outputs(5810)) xor (layer5_outputs(1873)));
    layer6_outputs(406) <= not((layer5_outputs(4756)) xor (layer5_outputs(7486)));
    layer6_outputs(407) <= not((layer5_outputs(5723)) xor (layer5_outputs(7104)));
    layer6_outputs(408) <= layer5_outputs(588);
    layer6_outputs(409) <= (layer5_outputs(717)) xor (layer5_outputs(4711));
    layer6_outputs(410) <= (layer5_outputs(7584)) xor (layer5_outputs(5052));
    layer6_outputs(411) <= not(layer5_outputs(3375));
    layer6_outputs(412) <= not(layer5_outputs(5287));
    layer6_outputs(413) <= not(layer5_outputs(646));
    layer6_outputs(414) <= layer5_outputs(596);
    layer6_outputs(415) <= layer5_outputs(5115);
    layer6_outputs(416) <= layer5_outputs(5533);
    layer6_outputs(417) <= layer5_outputs(7016);
    layer6_outputs(418) <= (layer5_outputs(5268)) xor (layer5_outputs(621));
    layer6_outputs(419) <= not(layer5_outputs(3839));
    layer6_outputs(420) <= not(layer5_outputs(6736));
    layer6_outputs(421) <= not((layer5_outputs(1904)) and (layer5_outputs(4840)));
    layer6_outputs(422) <= layer5_outputs(2495);
    layer6_outputs(423) <= not(layer5_outputs(7305));
    layer6_outputs(424) <= not(layer5_outputs(5984)) or (layer5_outputs(2984));
    layer6_outputs(425) <= not(layer5_outputs(1319));
    layer6_outputs(426) <= layer5_outputs(7623);
    layer6_outputs(427) <= layer5_outputs(157);
    layer6_outputs(428) <= layer5_outputs(619);
    layer6_outputs(429) <= not((layer5_outputs(3531)) xor (layer5_outputs(4442)));
    layer6_outputs(430) <= not(layer5_outputs(2462)) or (layer5_outputs(6831));
    layer6_outputs(431) <= (layer5_outputs(2486)) or (layer5_outputs(7209));
    layer6_outputs(432) <= not(layer5_outputs(3442));
    layer6_outputs(433) <= not(layer5_outputs(2253));
    layer6_outputs(434) <= not((layer5_outputs(4394)) and (layer5_outputs(5988)));
    layer6_outputs(435) <= not((layer5_outputs(3765)) xor (layer5_outputs(1395)));
    layer6_outputs(436) <= layer5_outputs(7066);
    layer6_outputs(437) <= not((layer5_outputs(449)) xor (layer5_outputs(4838)));
    layer6_outputs(438) <= layer5_outputs(3977);
    layer6_outputs(439) <= (layer5_outputs(1122)) and not (layer5_outputs(135));
    layer6_outputs(440) <= (layer5_outputs(4724)) or (layer5_outputs(5991));
    layer6_outputs(441) <= not(layer5_outputs(4280));
    layer6_outputs(442) <= not(layer5_outputs(6030));
    layer6_outputs(443) <= layer5_outputs(2566);
    layer6_outputs(444) <= (layer5_outputs(7227)) xor (layer5_outputs(2710));
    layer6_outputs(445) <= (layer5_outputs(6316)) or (layer5_outputs(6476));
    layer6_outputs(446) <= (layer5_outputs(3026)) xor (layer5_outputs(1031));
    layer6_outputs(447) <= (layer5_outputs(6336)) and (layer5_outputs(4314));
    layer6_outputs(448) <= not((layer5_outputs(1301)) xor (layer5_outputs(6546)));
    layer6_outputs(449) <= not(layer5_outputs(3743));
    layer6_outputs(450) <= not(layer5_outputs(5854));
    layer6_outputs(451) <= not(layer5_outputs(2913));
    layer6_outputs(452) <= layer5_outputs(5293);
    layer6_outputs(453) <= (layer5_outputs(4333)) and (layer5_outputs(2556));
    layer6_outputs(454) <= not(layer5_outputs(935));
    layer6_outputs(455) <= layer5_outputs(4878);
    layer6_outputs(456) <= (layer5_outputs(2505)) xor (layer5_outputs(3657));
    layer6_outputs(457) <= (layer5_outputs(2751)) and (layer5_outputs(2769));
    layer6_outputs(458) <= not((layer5_outputs(5290)) or (layer5_outputs(3436)));
    layer6_outputs(459) <= layer5_outputs(4836);
    layer6_outputs(460) <= not(layer5_outputs(1681));
    layer6_outputs(461) <= (layer5_outputs(3166)) and (layer5_outputs(3096));
    layer6_outputs(462) <= layer5_outputs(6522);
    layer6_outputs(463) <= not(layer5_outputs(1001));
    layer6_outputs(464) <= not(layer5_outputs(6172));
    layer6_outputs(465) <= (layer5_outputs(2312)) or (layer5_outputs(6818));
    layer6_outputs(466) <= (layer5_outputs(6917)) and (layer5_outputs(5353));
    layer6_outputs(467) <= not(layer5_outputs(5822));
    layer6_outputs(468) <= not((layer5_outputs(1675)) and (layer5_outputs(5041)));
    layer6_outputs(469) <= not((layer5_outputs(7418)) or (layer5_outputs(6665)));
    layer6_outputs(470) <= (layer5_outputs(216)) and not (layer5_outputs(7063));
    layer6_outputs(471) <= not(layer5_outputs(1583)) or (layer5_outputs(2755));
    layer6_outputs(472) <= (layer5_outputs(596)) and not (layer5_outputs(4079));
    layer6_outputs(473) <= not(layer5_outputs(3595));
    layer6_outputs(474) <= layer5_outputs(5835);
    layer6_outputs(475) <= not(layer5_outputs(4120));
    layer6_outputs(476) <= layer5_outputs(2302);
    layer6_outputs(477) <= not((layer5_outputs(3579)) and (layer5_outputs(1602)));
    layer6_outputs(478) <= not(layer5_outputs(6849)) or (layer5_outputs(6863));
    layer6_outputs(479) <= layer5_outputs(5216);
    layer6_outputs(480) <= layer5_outputs(3758);
    layer6_outputs(481) <= not(layer5_outputs(4059));
    layer6_outputs(482) <= layer5_outputs(2552);
    layer6_outputs(483) <= not((layer5_outputs(4992)) xor (layer5_outputs(1906)));
    layer6_outputs(484) <= '0';
    layer6_outputs(485) <= not(layer5_outputs(5542)) or (layer5_outputs(4591));
    layer6_outputs(486) <= not(layer5_outputs(1093));
    layer6_outputs(487) <= layer5_outputs(6332);
    layer6_outputs(488) <= (layer5_outputs(976)) xor (layer5_outputs(6834));
    layer6_outputs(489) <= layer5_outputs(629);
    layer6_outputs(490) <= not((layer5_outputs(1214)) xor (layer5_outputs(1841)));
    layer6_outputs(491) <= not((layer5_outputs(1320)) xor (layer5_outputs(3562)));
    layer6_outputs(492) <= (layer5_outputs(4862)) and not (layer5_outputs(4031));
    layer6_outputs(493) <= (layer5_outputs(1059)) and not (layer5_outputs(7332));
    layer6_outputs(494) <= (layer5_outputs(4063)) xor (layer5_outputs(4342));
    layer6_outputs(495) <= (layer5_outputs(5313)) xor (layer5_outputs(5666));
    layer6_outputs(496) <= layer5_outputs(4097);
    layer6_outputs(497) <= not((layer5_outputs(2563)) xor (layer5_outputs(4703)));
    layer6_outputs(498) <= (layer5_outputs(4505)) and (layer5_outputs(4924));
    layer6_outputs(499) <= layer5_outputs(7287);
    layer6_outputs(500) <= layer5_outputs(2483);
    layer6_outputs(501) <= (layer5_outputs(1799)) and not (layer5_outputs(326));
    layer6_outputs(502) <= '0';
    layer6_outputs(503) <= not((layer5_outputs(1061)) xor (layer5_outputs(3931)));
    layer6_outputs(504) <= layer5_outputs(1042);
    layer6_outputs(505) <= not(layer5_outputs(785)) or (layer5_outputs(2509));
    layer6_outputs(506) <= not(layer5_outputs(2903));
    layer6_outputs(507) <= not(layer5_outputs(1239));
    layer6_outputs(508) <= not(layer5_outputs(746));
    layer6_outputs(509) <= layer5_outputs(7465);
    layer6_outputs(510) <= not((layer5_outputs(7318)) xor (layer5_outputs(575)));
    layer6_outputs(511) <= not((layer5_outputs(1455)) xor (layer5_outputs(4656)));
    layer6_outputs(512) <= (layer5_outputs(4997)) xor (layer5_outputs(6596));
    layer6_outputs(513) <= layer5_outputs(6784);
    layer6_outputs(514) <= (layer5_outputs(5552)) and not (layer5_outputs(1105));
    layer6_outputs(515) <= (layer5_outputs(2769)) xor (layer5_outputs(7330));
    layer6_outputs(516) <= not(layer5_outputs(5438)) or (layer5_outputs(5385));
    layer6_outputs(517) <= not(layer5_outputs(2853));
    layer6_outputs(518) <= (layer5_outputs(5535)) xor (layer5_outputs(1543));
    layer6_outputs(519) <= not(layer5_outputs(979));
    layer6_outputs(520) <= not(layer5_outputs(3952));
    layer6_outputs(521) <= not((layer5_outputs(5511)) xor (layer5_outputs(7497)));
    layer6_outputs(522) <= not(layer5_outputs(3998));
    layer6_outputs(523) <= layer5_outputs(6606);
    layer6_outputs(524) <= layer5_outputs(6463);
    layer6_outputs(525) <= not((layer5_outputs(3704)) xor (layer5_outputs(3731)));
    layer6_outputs(526) <= layer5_outputs(314);
    layer6_outputs(527) <= layer5_outputs(1309);
    layer6_outputs(528) <= not(layer5_outputs(4660));
    layer6_outputs(529) <= not(layer5_outputs(4052)) or (layer5_outputs(6245));
    layer6_outputs(530) <= not(layer5_outputs(1547)) or (layer5_outputs(5454));
    layer6_outputs(531) <= layer5_outputs(884);
    layer6_outputs(532) <= not(layer5_outputs(3803));
    layer6_outputs(533) <= layer5_outputs(1256);
    layer6_outputs(534) <= not(layer5_outputs(986));
    layer6_outputs(535) <= not(layer5_outputs(2831));
    layer6_outputs(536) <= not(layer5_outputs(1091));
    layer6_outputs(537) <= not(layer5_outputs(6404));
    layer6_outputs(538) <= layer5_outputs(2877);
    layer6_outputs(539) <= (layer5_outputs(959)) or (layer5_outputs(734));
    layer6_outputs(540) <= not((layer5_outputs(2494)) and (layer5_outputs(2592)));
    layer6_outputs(541) <= not((layer5_outputs(1336)) or (layer5_outputs(7401)));
    layer6_outputs(542) <= (layer5_outputs(3672)) and (layer5_outputs(6420));
    layer6_outputs(543) <= not((layer5_outputs(2530)) xor (layer5_outputs(5305)));
    layer6_outputs(544) <= layer5_outputs(1835);
    layer6_outputs(545) <= not(layer5_outputs(6727)) or (layer5_outputs(1350));
    layer6_outputs(546) <= not((layer5_outputs(2417)) or (layer5_outputs(5970)));
    layer6_outputs(547) <= layer5_outputs(1736);
    layer6_outputs(548) <= (layer5_outputs(2105)) or (layer5_outputs(6978));
    layer6_outputs(549) <= (layer5_outputs(5669)) and not (layer5_outputs(767));
    layer6_outputs(550) <= (layer5_outputs(4144)) and not (layer5_outputs(6479));
    layer6_outputs(551) <= not(layer5_outputs(7564)) or (layer5_outputs(2021));
    layer6_outputs(552) <= (layer5_outputs(4188)) and not (layer5_outputs(2714));
    layer6_outputs(553) <= layer5_outputs(6093);
    layer6_outputs(554) <= not(layer5_outputs(4822)) or (layer5_outputs(7377));
    layer6_outputs(555) <= not(layer5_outputs(6677));
    layer6_outputs(556) <= (layer5_outputs(3858)) xor (layer5_outputs(2112));
    layer6_outputs(557) <= (layer5_outputs(6752)) or (layer5_outputs(5614));
    layer6_outputs(558) <= not(layer5_outputs(1341));
    layer6_outputs(559) <= not(layer5_outputs(4549));
    layer6_outputs(560) <= not(layer5_outputs(3346));
    layer6_outputs(561) <= not(layer5_outputs(6215)) or (layer5_outputs(713));
    layer6_outputs(562) <= layer5_outputs(3052);
    layer6_outputs(563) <= not((layer5_outputs(3609)) and (layer5_outputs(4261)));
    layer6_outputs(564) <= (layer5_outputs(311)) xor (layer5_outputs(6485));
    layer6_outputs(565) <= not(layer5_outputs(6180));
    layer6_outputs(566) <= layer5_outputs(7072);
    layer6_outputs(567) <= not(layer5_outputs(6950));
    layer6_outputs(568) <= not(layer5_outputs(6279));
    layer6_outputs(569) <= not(layer5_outputs(6438)) or (layer5_outputs(7269));
    layer6_outputs(570) <= (layer5_outputs(2420)) xor (layer5_outputs(2206));
    layer6_outputs(571) <= not(layer5_outputs(6956));
    layer6_outputs(572) <= layer5_outputs(7110);
    layer6_outputs(573) <= (layer5_outputs(5492)) xor (layer5_outputs(5764));
    layer6_outputs(574) <= not(layer5_outputs(2844)) or (layer5_outputs(3811));
    layer6_outputs(575) <= not((layer5_outputs(4368)) and (layer5_outputs(5002)));
    layer6_outputs(576) <= '0';
    layer6_outputs(577) <= not(layer5_outputs(4111));
    layer6_outputs(578) <= not(layer5_outputs(3491));
    layer6_outputs(579) <= layer5_outputs(6983);
    layer6_outputs(580) <= layer5_outputs(3652);
    layer6_outputs(581) <= not(layer5_outputs(183));
    layer6_outputs(582) <= layer5_outputs(2310);
    layer6_outputs(583) <= (layer5_outputs(4218)) xor (layer5_outputs(3396));
    layer6_outputs(584) <= layer5_outputs(847);
    layer6_outputs(585) <= layer5_outputs(4886);
    layer6_outputs(586) <= not((layer5_outputs(6428)) and (layer5_outputs(6520)));
    layer6_outputs(587) <= layer5_outputs(3382);
    layer6_outputs(588) <= layer5_outputs(3226);
    layer6_outputs(589) <= not((layer5_outputs(6372)) or (layer5_outputs(5207)));
    layer6_outputs(590) <= layer5_outputs(7625);
    layer6_outputs(591) <= layer5_outputs(3724);
    layer6_outputs(592) <= not(layer5_outputs(4304));
    layer6_outputs(593) <= not((layer5_outputs(3891)) or (layer5_outputs(2212)));
    layer6_outputs(594) <= not(layer5_outputs(7671));
    layer6_outputs(595) <= layer5_outputs(6640);
    layer6_outputs(596) <= (layer5_outputs(779)) and (layer5_outputs(4566));
    layer6_outputs(597) <= not(layer5_outputs(931));
    layer6_outputs(598) <= layer5_outputs(1996);
    layer6_outputs(599) <= layer5_outputs(4243);
    layer6_outputs(600) <= (layer5_outputs(1850)) or (layer5_outputs(6081));
    layer6_outputs(601) <= (layer5_outputs(5681)) or (layer5_outputs(7591));
    layer6_outputs(602) <= not(layer5_outputs(6189));
    layer6_outputs(603) <= (layer5_outputs(4155)) xor (layer5_outputs(6667));
    layer6_outputs(604) <= layer5_outputs(7588);
    layer6_outputs(605) <= not((layer5_outputs(4425)) or (layer5_outputs(790)));
    layer6_outputs(606) <= (layer5_outputs(4163)) xor (layer5_outputs(7481));
    layer6_outputs(607) <= not((layer5_outputs(5780)) or (layer5_outputs(2387)));
    layer6_outputs(608) <= (layer5_outputs(2509)) xor (layer5_outputs(6547));
    layer6_outputs(609) <= not(layer5_outputs(3070));
    layer6_outputs(610) <= (layer5_outputs(7661)) and not (layer5_outputs(3918));
    layer6_outputs(611) <= layer5_outputs(5526);
    layer6_outputs(612) <= not(layer5_outputs(2744));
    layer6_outputs(613) <= layer5_outputs(7346);
    layer6_outputs(614) <= not(layer5_outputs(868));
    layer6_outputs(615) <= (layer5_outputs(4933)) xor (layer5_outputs(124));
    layer6_outputs(616) <= (layer5_outputs(2113)) xor (layer5_outputs(3472));
    layer6_outputs(617) <= layer5_outputs(6759);
    layer6_outputs(618) <= (layer5_outputs(6807)) xor (layer5_outputs(4740));
    layer6_outputs(619) <= not(layer5_outputs(4831));
    layer6_outputs(620) <= (layer5_outputs(4946)) and not (layer5_outputs(3295));
    layer6_outputs(621) <= not((layer5_outputs(1)) or (layer5_outputs(5602)));
    layer6_outputs(622) <= not((layer5_outputs(6787)) and (layer5_outputs(5421)));
    layer6_outputs(623) <= not(layer5_outputs(7028));
    layer6_outputs(624) <= (layer5_outputs(3722)) xor (layer5_outputs(7124));
    layer6_outputs(625) <= not(layer5_outputs(6419));
    layer6_outputs(626) <= not((layer5_outputs(4938)) and (layer5_outputs(7502)));
    layer6_outputs(627) <= (layer5_outputs(6906)) or (layer5_outputs(6302));
    layer6_outputs(628) <= not(layer5_outputs(5532));
    layer6_outputs(629) <= layer5_outputs(4890);
    layer6_outputs(630) <= not((layer5_outputs(1957)) or (layer5_outputs(4898)));
    layer6_outputs(631) <= (layer5_outputs(6498)) or (layer5_outputs(2748));
    layer6_outputs(632) <= layer5_outputs(1159);
    layer6_outputs(633) <= not(layer5_outputs(1865));
    layer6_outputs(634) <= not(layer5_outputs(3322));
    layer6_outputs(635) <= not(layer5_outputs(7510)) or (layer5_outputs(2763));
    layer6_outputs(636) <= not((layer5_outputs(4867)) xor (layer5_outputs(3588)));
    layer6_outputs(637) <= not((layer5_outputs(5300)) xor (layer5_outputs(4690)));
    layer6_outputs(638) <= '0';
    layer6_outputs(639) <= not(layer5_outputs(2598));
    layer6_outputs(640) <= not(layer5_outputs(6769));
    layer6_outputs(641) <= not(layer5_outputs(1432));
    layer6_outputs(642) <= not((layer5_outputs(3016)) xor (layer5_outputs(2466)));
    layer6_outputs(643) <= layer5_outputs(7283);
    layer6_outputs(644) <= layer5_outputs(4302);
    layer6_outputs(645) <= (layer5_outputs(699)) or (layer5_outputs(6910));
    layer6_outputs(646) <= not(layer5_outputs(1976));
    layer6_outputs(647) <= layer5_outputs(5017);
    layer6_outputs(648) <= not(layer5_outputs(6145));
    layer6_outputs(649) <= layer5_outputs(2548);
    layer6_outputs(650) <= not(layer5_outputs(2197));
    layer6_outputs(651) <= layer5_outputs(1753);
    layer6_outputs(652) <= (layer5_outputs(5962)) and not (layer5_outputs(6173));
    layer6_outputs(653) <= not(layer5_outputs(784));
    layer6_outputs(654) <= layer5_outputs(3137);
    layer6_outputs(655) <= layer5_outputs(7585);
    layer6_outputs(656) <= (layer5_outputs(5467)) and (layer5_outputs(4618));
    layer6_outputs(657) <= layer5_outputs(5403);
    layer6_outputs(658) <= layer5_outputs(7393);
    layer6_outputs(659) <= layer5_outputs(5979);
    layer6_outputs(660) <= not(layer5_outputs(5575)) or (layer5_outputs(5219));
    layer6_outputs(661) <= not((layer5_outputs(2469)) and (layer5_outputs(2595)));
    layer6_outputs(662) <= (layer5_outputs(5024)) and not (layer5_outputs(7148));
    layer6_outputs(663) <= layer5_outputs(2914);
    layer6_outputs(664) <= layer5_outputs(6697);
    layer6_outputs(665) <= not(layer5_outputs(2810));
    layer6_outputs(666) <= layer5_outputs(7367);
    layer6_outputs(667) <= not(layer5_outputs(2135));
    layer6_outputs(668) <= not((layer5_outputs(2369)) xor (layer5_outputs(6754)));
    layer6_outputs(669) <= not(layer5_outputs(681)) or (layer5_outputs(5316));
    layer6_outputs(670) <= (layer5_outputs(5377)) and not (layer5_outputs(151));
    layer6_outputs(671) <= not(layer5_outputs(15));
    layer6_outputs(672) <= not(layer5_outputs(6581));
    layer6_outputs(673) <= not((layer5_outputs(7193)) or (layer5_outputs(5992)));
    layer6_outputs(674) <= not(layer5_outputs(3228));
    layer6_outputs(675) <= not((layer5_outputs(6286)) or (layer5_outputs(1725)));
    layer6_outputs(676) <= layer5_outputs(3028);
    layer6_outputs(677) <= not((layer5_outputs(1303)) xor (layer5_outputs(5540)));
    layer6_outputs(678) <= layer5_outputs(736);
    layer6_outputs(679) <= layer5_outputs(7043);
    layer6_outputs(680) <= layer5_outputs(5147);
    layer6_outputs(681) <= not((layer5_outputs(4377)) xor (layer5_outputs(917)));
    layer6_outputs(682) <= not((layer5_outputs(599)) xor (layer5_outputs(231)));
    layer6_outputs(683) <= layer5_outputs(1258);
    layer6_outputs(684) <= not(layer5_outputs(5171));
    layer6_outputs(685) <= (layer5_outputs(5489)) xor (layer5_outputs(285));
    layer6_outputs(686) <= layer5_outputs(7290);
    layer6_outputs(687) <= layer5_outputs(7599);
    layer6_outputs(688) <= layer5_outputs(5826);
    layer6_outputs(689) <= not(layer5_outputs(5897));
    layer6_outputs(690) <= not((layer5_outputs(7658)) or (layer5_outputs(666)));
    layer6_outputs(691) <= layer5_outputs(3625);
    layer6_outputs(692) <= (layer5_outputs(2113)) and not (layer5_outputs(6008));
    layer6_outputs(693) <= not(layer5_outputs(1981));
    layer6_outputs(694) <= not((layer5_outputs(3453)) and (layer5_outputs(7098)));
    layer6_outputs(695) <= (layer5_outputs(1340)) and (layer5_outputs(298));
    layer6_outputs(696) <= not((layer5_outputs(6155)) or (layer5_outputs(4019)));
    layer6_outputs(697) <= not(layer5_outputs(6913));
    layer6_outputs(698) <= not(layer5_outputs(1095));
    layer6_outputs(699) <= layer5_outputs(3781);
    layer6_outputs(700) <= not(layer5_outputs(2490));
    layer6_outputs(701) <= not((layer5_outputs(7637)) xor (layer5_outputs(3820)));
    layer6_outputs(702) <= not(layer5_outputs(5796)) or (layer5_outputs(2006));
    layer6_outputs(703) <= not((layer5_outputs(4537)) or (layer5_outputs(6492)));
    layer6_outputs(704) <= layer5_outputs(3231);
    layer6_outputs(705) <= (layer5_outputs(4468)) and (layer5_outputs(3507));
    layer6_outputs(706) <= not(layer5_outputs(1321));
    layer6_outputs(707) <= not(layer5_outputs(1157)) or (layer5_outputs(5500));
    layer6_outputs(708) <= (layer5_outputs(5573)) xor (layer5_outputs(3877));
    layer6_outputs(709) <= not(layer5_outputs(3431));
    layer6_outputs(710) <= (layer5_outputs(3595)) and not (layer5_outputs(5904));
    layer6_outputs(711) <= layer5_outputs(1570);
    layer6_outputs(712) <= layer5_outputs(6288);
    layer6_outputs(713) <= layer5_outputs(41);
    layer6_outputs(714) <= layer5_outputs(7570);
    layer6_outputs(715) <= not(layer5_outputs(2894));
    layer6_outputs(716) <= '0';
    layer6_outputs(717) <= not(layer5_outputs(7205));
    layer6_outputs(718) <= not(layer5_outputs(4335)) or (layer5_outputs(3078));
    layer6_outputs(719) <= layer5_outputs(1740);
    layer6_outputs(720) <= not(layer5_outputs(611));
    layer6_outputs(721) <= not(layer5_outputs(1178));
    layer6_outputs(722) <= not(layer5_outputs(656));
    layer6_outputs(723) <= not(layer5_outputs(6399));
    layer6_outputs(724) <= not((layer5_outputs(4880)) xor (layer5_outputs(2290)));
    layer6_outputs(725) <= layer5_outputs(3357);
    layer6_outputs(726) <= layer5_outputs(3904);
    layer6_outputs(727) <= layer5_outputs(5755);
    layer6_outputs(728) <= not((layer5_outputs(5609)) and (layer5_outputs(310)));
    layer6_outputs(729) <= not(layer5_outputs(3262));
    layer6_outputs(730) <= not(layer5_outputs(2552)) or (layer5_outputs(1919));
    layer6_outputs(731) <= layer5_outputs(5024);
    layer6_outputs(732) <= not((layer5_outputs(3607)) xor (layer5_outputs(634)));
    layer6_outputs(733) <= layer5_outputs(7492);
    layer6_outputs(734) <= (layer5_outputs(1751)) and (layer5_outputs(6234));
    layer6_outputs(735) <= not((layer5_outputs(3923)) xor (layer5_outputs(3474)));
    layer6_outputs(736) <= not(layer5_outputs(5374));
    layer6_outputs(737) <= layer5_outputs(2765);
    layer6_outputs(738) <= layer5_outputs(3131);
    layer6_outputs(739) <= layer5_outputs(728);
    layer6_outputs(740) <= layer5_outputs(3281);
    layer6_outputs(741) <= not((layer5_outputs(3057)) xor (layer5_outputs(2215)));
    layer6_outputs(742) <= not(layer5_outputs(3221));
    layer6_outputs(743) <= not(layer5_outputs(4981)) or (layer5_outputs(1144));
    layer6_outputs(744) <= not(layer5_outputs(267)) or (layer5_outputs(3999));
    layer6_outputs(745) <= not(layer5_outputs(6064)) or (layer5_outputs(5896));
    layer6_outputs(746) <= not((layer5_outputs(4936)) or (layer5_outputs(183)));
    layer6_outputs(747) <= not(layer5_outputs(5472));
    layer6_outputs(748) <= (layer5_outputs(2852)) or (layer5_outputs(3408));
    layer6_outputs(749) <= (layer5_outputs(3164)) and not (layer5_outputs(430));
    layer6_outputs(750) <= (layer5_outputs(5211)) and not (layer5_outputs(5318));
    layer6_outputs(751) <= layer5_outputs(3863);
    layer6_outputs(752) <= not(layer5_outputs(7664));
    layer6_outputs(753) <= not(layer5_outputs(6903));
    layer6_outputs(754) <= layer5_outputs(2605);
    layer6_outputs(755) <= not(layer5_outputs(6717));
    layer6_outputs(756) <= not(layer5_outputs(856));
    layer6_outputs(757) <= not(layer5_outputs(3234));
    layer6_outputs(758) <= not(layer5_outputs(1233));
    layer6_outputs(759) <= layer5_outputs(13);
    layer6_outputs(760) <= not(layer5_outputs(5601)) or (layer5_outputs(6928));
    layer6_outputs(761) <= (layer5_outputs(7531)) and not (layer5_outputs(4181));
    layer6_outputs(762) <= not(layer5_outputs(3101));
    layer6_outputs(763) <= (layer5_outputs(5090)) xor (layer5_outputs(4855));
    layer6_outputs(764) <= layer5_outputs(3537);
    layer6_outputs(765) <= (layer5_outputs(4708)) and (layer5_outputs(5538));
    layer6_outputs(766) <= not(layer5_outputs(619));
    layer6_outputs(767) <= not(layer5_outputs(3756));
    layer6_outputs(768) <= not(layer5_outputs(6352));
    layer6_outputs(769) <= not(layer5_outputs(4887));
    layer6_outputs(770) <= not(layer5_outputs(649));
    layer6_outputs(771) <= (layer5_outputs(5623)) and (layer5_outputs(2886));
    layer6_outputs(772) <= (layer5_outputs(6937)) and not (layer5_outputs(2841));
    layer6_outputs(773) <= (layer5_outputs(1333)) and (layer5_outputs(7518));
    layer6_outputs(774) <= (layer5_outputs(2347)) and not (layer5_outputs(2679));
    layer6_outputs(775) <= layer5_outputs(3648);
    layer6_outputs(776) <= not((layer5_outputs(5784)) or (layer5_outputs(6675)));
    layer6_outputs(777) <= layer5_outputs(6593);
    layer6_outputs(778) <= not(layer5_outputs(4308));
    layer6_outputs(779) <= not(layer5_outputs(6934));
    layer6_outputs(780) <= (layer5_outputs(5407)) and not (layer5_outputs(2481));
    layer6_outputs(781) <= layer5_outputs(2287);
    layer6_outputs(782) <= (layer5_outputs(6997)) and (layer5_outputs(5042));
    layer6_outputs(783) <= not((layer5_outputs(5495)) and (layer5_outputs(6484)));
    layer6_outputs(784) <= not((layer5_outputs(98)) or (layer5_outputs(3056)));
    layer6_outputs(785) <= not(layer5_outputs(426));
    layer6_outputs(786) <= not(layer5_outputs(6905));
    layer6_outputs(787) <= (layer5_outputs(5256)) and not (layer5_outputs(5535));
    layer6_outputs(788) <= layer5_outputs(3885);
    layer6_outputs(789) <= layer5_outputs(3415);
    layer6_outputs(790) <= not((layer5_outputs(2220)) and (layer5_outputs(7370)));
    layer6_outputs(791) <= (layer5_outputs(7495)) and not (layer5_outputs(5471));
    layer6_outputs(792) <= not(layer5_outputs(4326));
    layer6_outputs(793) <= not(layer5_outputs(5707));
    layer6_outputs(794) <= not((layer5_outputs(6460)) and (layer5_outputs(5526)));
    layer6_outputs(795) <= layer5_outputs(4273);
    layer6_outputs(796) <= not((layer5_outputs(5427)) xor (layer5_outputs(7240)));
    layer6_outputs(797) <= not((layer5_outputs(3866)) xor (layer5_outputs(85)));
    layer6_outputs(798) <= (layer5_outputs(4306)) and (layer5_outputs(6625));
    layer6_outputs(799) <= not(layer5_outputs(1697)) or (layer5_outputs(1872));
    layer6_outputs(800) <= '0';
    layer6_outputs(801) <= not((layer5_outputs(744)) xor (layer5_outputs(1774)));
    layer6_outputs(802) <= layer5_outputs(983);
    layer6_outputs(803) <= layer5_outputs(586);
    layer6_outputs(804) <= not(layer5_outputs(101)) or (layer5_outputs(107));
    layer6_outputs(805) <= layer5_outputs(1617);
    layer6_outputs(806) <= not((layer5_outputs(2474)) xor (layer5_outputs(4991)));
    layer6_outputs(807) <= layer5_outputs(6963);
    layer6_outputs(808) <= not((layer5_outputs(90)) xor (layer5_outputs(1042)));
    layer6_outputs(809) <= not(layer5_outputs(963)) or (layer5_outputs(4620));
    layer6_outputs(810) <= layer5_outputs(457);
    layer6_outputs(811) <= not(layer5_outputs(7089)) or (layer5_outputs(1950));
    layer6_outputs(812) <= not(layer5_outputs(4841));
    layer6_outputs(813) <= not((layer5_outputs(5680)) xor (layer5_outputs(2890)));
    layer6_outputs(814) <= not(layer5_outputs(655)) or (layer5_outputs(5032));
    layer6_outputs(815) <= layer5_outputs(7306);
    layer6_outputs(816) <= layer5_outputs(7076);
    layer6_outputs(817) <= layer5_outputs(384);
    layer6_outputs(818) <= not((layer5_outputs(292)) xor (layer5_outputs(4989)));
    layer6_outputs(819) <= not(layer5_outputs(3618));
    layer6_outputs(820) <= layer5_outputs(4960);
    layer6_outputs(821) <= not((layer5_outputs(1072)) and (layer5_outputs(4510)));
    layer6_outputs(822) <= (layer5_outputs(1407)) xor (layer5_outputs(4700));
    layer6_outputs(823) <= layer5_outputs(1597);
    layer6_outputs(824) <= not(layer5_outputs(1044));
    layer6_outputs(825) <= not(layer5_outputs(2615));
    layer6_outputs(826) <= not(layer5_outputs(1039));
    layer6_outputs(827) <= not(layer5_outputs(868));
    layer6_outputs(828) <= not(layer5_outputs(4713)) or (layer5_outputs(1337));
    layer6_outputs(829) <= layer5_outputs(3449);
    layer6_outputs(830) <= layer5_outputs(4684);
    layer6_outputs(831) <= (layer5_outputs(7559)) xor (layer5_outputs(5166));
    layer6_outputs(832) <= (layer5_outputs(2575)) and not (layer5_outputs(6778));
    layer6_outputs(833) <= not(layer5_outputs(6020)) or (layer5_outputs(1524));
    layer6_outputs(834) <= layer5_outputs(4162);
    layer6_outputs(835) <= (layer5_outputs(952)) xor (layer5_outputs(3925));
    layer6_outputs(836) <= layer5_outputs(3038);
    layer6_outputs(837) <= not(layer5_outputs(7290)) or (layer5_outputs(1848));
    layer6_outputs(838) <= not(layer5_outputs(5861));
    layer6_outputs(839) <= layer5_outputs(3318);
    layer6_outputs(840) <= not(layer5_outputs(1606));
    layer6_outputs(841) <= not(layer5_outputs(5961));
    layer6_outputs(842) <= not(layer5_outputs(4860));
    layer6_outputs(843) <= (layer5_outputs(2659)) or (layer5_outputs(6327));
    layer6_outputs(844) <= not((layer5_outputs(1956)) and (layer5_outputs(5987)));
    layer6_outputs(845) <= layer5_outputs(2422);
    layer6_outputs(846) <= not((layer5_outputs(1474)) or (layer5_outputs(716)));
    layer6_outputs(847) <= not((layer5_outputs(493)) xor (layer5_outputs(4119)));
    layer6_outputs(848) <= not((layer5_outputs(2897)) xor (layer5_outputs(1411)));
    layer6_outputs(849) <= not((layer5_outputs(5743)) or (layer5_outputs(1091)));
    layer6_outputs(850) <= (layer5_outputs(1486)) and not (layer5_outputs(5315));
    layer6_outputs(851) <= (layer5_outputs(3408)) and not (layer5_outputs(2512));
    layer6_outputs(852) <= not((layer5_outputs(1552)) and (layer5_outputs(250)));
    layer6_outputs(853) <= layer5_outputs(7247);
    layer6_outputs(854) <= not((layer5_outputs(6869)) xor (layer5_outputs(2641)));
    layer6_outputs(855) <= layer5_outputs(5954);
    layer6_outputs(856) <= layer5_outputs(2528);
    layer6_outputs(857) <= (layer5_outputs(6384)) and not (layer5_outputs(2362));
    layer6_outputs(858) <= (layer5_outputs(258)) xor (layer5_outputs(7204));
    layer6_outputs(859) <= layer5_outputs(5609);
    layer6_outputs(860) <= not(layer5_outputs(840));
    layer6_outputs(861) <= not((layer5_outputs(1732)) xor (layer5_outputs(5067)));
    layer6_outputs(862) <= (layer5_outputs(7250)) and not (layer5_outputs(5694));
    layer6_outputs(863) <= (layer5_outputs(2644)) xor (layer5_outputs(7448));
    layer6_outputs(864) <= not((layer5_outputs(1422)) or (layer5_outputs(7361)));
    layer6_outputs(865) <= not(layer5_outputs(7540));
    layer6_outputs(866) <= not(layer5_outputs(1137));
    layer6_outputs(867) <= not(layer5_outputs(5483));
    layer6_outputs(868) <= not(layer5_outputs(6509));
    layer6_outputs(869) <= (layer5_outputs(7308)) and not (layer5_outputs(870));
    layer6_outputs(870) <= not(layer5_outputs(6745));
    layer6_outputs(871) <= layer5_outputs(1556);
    layer6_outputs(872) <= layer5_outputs(5392);
    layer6_outputs(873) <= not((layer5_outputs(407)) xor (layer5_outputs(4556)));
    layer6_outputs(874) <= (layer5_outputs(175)) and not (layer5_outputs(4908));
    layer6_outputs(875) <= not((layer5_outputs(6108)) or (layer5_outputs(7423)));
    layer6_outputs(876) <= (layer5_outputs(204)) and not (layer5_outputs(7655));
    layer6_outputs(877) <= not(layer5_outputs(2412)) or (layer5_outputs(5697));
    layer6_outputs(878) <= (layer5_outputs(707)) and not (layer5_outputs(6132));
    layer6_outputs(879) <= (layer5_outputs(4619)) or (layer5_outputs(2188));
    layer6_outputs(880) <= (layer5_outputs(7039)) and not (layer5_outputs(1571));
    layer6_outputs(881) <= layer5_outputs(1048);
    layer6_outputs(882) <= not(layer5_outputs(1498));
    layer6_outputs(883) <= layer5_outputs(1076);
    layer6_outputs(884) <= (layer5_outputs(7623)) and not (layer5_outputs(1719));
    layer6_outputs(885) <= not(layer5_outputs(7263));
    layer6_outputs(886) <= (layer5_outputs(1034)) xor (layer5_outputs(5301));
    layer6_outputs(887) <= not((layer5_outputs(4504)) xor (layer5_outputs(7423)));
    layer6_outputs(888) <= (layer5_outputs(4250)) and not (layer5_outputs(1342));
    layer6_outputs(889) <= layer5_outputs(1019);
    layer6_outputs(890) <= not(layer5_outputs(1070));
    layer6_outputs(891) <= not((layer5_outputs(3519)) xor (layer5_outputs(2652)));
    layer6_outputs(892) <= not(layer5_outputs(7294)) or (layer5_outputs(4316));
    layer6_outputs(893) <= not(layer5_outputs(5106)) or (layer5_outputs(1006));
    layer6_outputs(894) <= not(layer5_outputs(3423));
    layer6_outputs(895) <= not(layer5_outputs(1101)) or (layer5_outputs(5443));
    layer6_outputs(896) <= not((layer5_outputs(61)) or (layer5_outputs(3157)));
    layer6_outputs(897) <= (layer5_outputs(6333)) and not (layer5_outputs(2185));
    layer6_outputs(898) <= '1';
    layer6_outputs(899) <= not(layer5_outputs(7394));
    layer6_outputs(900) <= not((layer5_outputs(6270)) and (layer5_outputs(1431)));
    layer6_outputs(901) <= not(layer5_outputs(6356));
    layer6_outputs(902) <= layer5_outputs(4409);
    layer6_outputs(903) <= not(layer5_outputs(7140)) or (layer5_outputs(2347));
    layer6_outputs(904) <= (layer5_outputs(7647)) or (layer5_outputs(2797));
    layer6_outputs(905) <= not(layer5_outputs(7324));
    layer6_outputs(906) <= (layer5_outputs(3400)) and (layer5_outputs(4101));
    layer6_outputs(907) <= not((layer5_outputs(3344)) xor (layer5_outputs(2724)));
    layer6_outputs(908) <= (layer5_outputs(5712)) and (layer5_outputs(6290));
    layer6_outputs(909) <= not(layer5_outputs(1750));
    layer6_outputs(910) <= layer5_outputs(2786);
    layer6_outputs(911) <= not((layer5_outputs(5356)) and (layer5_outputs(2011)));
    layer6_outputs(912) <= layer5_outputs(4906);
    layer6_outputs(913) <= (layer5_outputs(5226)) and not (layer5_outputs(6999));
    layer6_outputs(914) <= not(layer5_outputs(3315));
    layer6_outputs(915) <= not(layer5_outputs(5627));
    layer6_outputs(916) <= layer5_outputs(1652);
    layer6_outputs(917) <= (layer5_outputs(5678)) or (layer5_outputs(2707));
    layer6_outputs(918) <= not(layer5_outputs(1675)) or (layer5_outputs(1635));
    layer6_outputs(919) <= not((layer5_outputs(7475)) xor (layer5_outputs(5727)));
    layer6_outputs(920) <= layer5_outputs(3040);
    layer6_outputs(921) <= layer5_outputs(2933);
    layer6_outputs(922) <= layer5_outputs(1813);
    layer6_outputs(923) <= (layer5_outputs(4000)) or (layer5_outputs(4272));
    layer6_outputs(924) <= (layer5_outputs(3587)) and not (layer5_outputs(1451));
    layer6_outputs(925) <= not(layer5_outputs(5393));
    layer6_outputs(926) <= not((layer5_outputs(7625)) xor (layer5_outputs(6343)));
    layer6_outputs(927) <= not(layer5_outputs(4712));
    layer6_outputs(928) <= not((layer5_outputs(253)) xor (layer5_outputs(2761)));
    layer6_outputs(929) <= layer5_outputs(1826);
    layer6_outputs(930) <= (layer5_outputs(3621)) and (layer5_outputs(7063));
    layer6_outputs(931) <= not(layer5_outputs(4546));
    layer6_outputs(932) <= not(layer5_outputs(901)) or (layer5_outputs(2512));
    layer6_outputs(933) <= not(layer5_outputs(5596));
    layer6_outputs(934) <= not((layer5_outputs(6450)) xor (layer5_outputs(7434)));
    layer6_outputs(935) <= layer5_outputs(850);
    layer6_outputs(936) <= not(layer5_outputs(7029));
    layer6_outputs(937) <= not(layer5_outputs(5691));
    layer6_outputs(938) <= layer5_outputs(7412);
    layer6_outputs(939) <= (layer5_outputs(50)) and not (layer5_outputs(1677));
    layer6_outputs(940) <= not((layer5_outputs(1818)) and (layer5_outputs(2503)));
    layer6_outputs(941) <= (layer5_outputs(4795)) or (layer5_outputs(3795));
    layer6_outputs(942) <= not((layer5_outputs(1517)) xor (layer5_outputs(2020)));
    layer6_outputs(943) <= (layer5_outputs(5462)) xor (layer5_outputs(6197));
    layer6_outputs(944) <= not(layer5_outputs(2267)) or (layer5_outputs(4320));
    layer6_outputs(945) <= (layer5_outputs(7453)) or (layer5_outputs(5540));
    layer6_outputs(946) <= (layer5_outputs(4026)) or (layer5_outputs(6386));
    layer6_outputs(947) <= (layer5_outputs(6204)) or (layer5_outputs(594));
    layer6_outputs(948) <= not(layer5_outputs(774));
    layer6_outputs(949) <= not(layer5_outputs(7432));
    layer6_outputs(950) <= not((layer5_outputs(890)) xor (layer5_outputs(6652)));
    layer6_outputs(951) <= not(layer5_outputs(7105));
    layer6_outputs(952) <= layer5_outputs(6903);
    layer6_outputs(953) <= layer5_outputs(4622);
    layer6_outputs(954) <= not((layer5_outputs(1668)) and (layer5_outputs(1862)));
    layer6_outputs(955) <= not((layer5_outputs(4628)) xor (layer5_outputs(669)));
    layer6_outputs(956) <= layer5_outputs(7094);
    layer6_outputs(957) <= '0';
    layer6_outputs(958) <= not(layer5_outputs(1090));
    layer6_outputs(959) <= layer5_outputs(399);
    layer6_outputs(960) <= layer5_outputs(576);
    layer6_outputs(961) <= (layer5_outputs(6639)) xor (layer5_outputs(2450));
    layer6_outputs(962) <= not(layer5_outputs(5367));
    layer6_outputs(963) <= (layer5_outputs(374)) or (layer5_outputs(7265));
    layer6_outputs(964) <= (layer5_outputs(2392)) or (layer5_outputs(7408));
    layer6_outputs(965) <= not(layer5_outputs(3824));
    layer6_outputs(966) <= not((layer5_outputs(5458)) or (layer5_outputs(3621)));
    layer6_outputs(967) <= not(layer5_outputs(3909));
    layer6_outputs(968) <= (layer5_outputs(3626)) or (layer5_outputs(6505));
    layer6_outputs(969) <= (layer5_outputs(398)) xor (layer5_outputs(3342));
    layer6_outputs(970) <= (layer5_outputs(536)) and not (layer5_outputs(7463));
    layer6_outputs(971) <= not((layer5_outputs(7646)) xor (layer5_outputs(5688)));
    layer6_outputs(972) <= not(layer5_outputs(5404));
    layer6_outputs(973) <= not(layer5_outputs(887));
    layer6_outputs(974) <= not((layer5_outputs(389)) xor (layer5_outputs(841)));
    layer6_outputs(975) <= not(layer5_outputs(3616));
    layer6_outputs(976) <= layer5_outputs(7217);
    layer6_outputs(977) <= not((layer5_outputs(979)) xor (layer5_outputs(5979)));
    layer6_outputs(978) <= (layer5_outputs(6781)) and (layer5_outputs(2634));
    layer6_outputs(979) <= (layer5_outputs(7478)) or (layer5_outputs(5617));
    layer6_outputs(980) <= not(layer5_outputs(6837));
    layer6_outputs(981) <= not((layer5_outputs(5776)) or (layer5_outputs(5790)));
    layer6_outputs(982) <= not((layer5_outputs(1669)) xor (layer5_outputs(7172)));
    layer6_outputs(983) <= layer5_outputs(3784);
    layer6_outputs(984) <= not(layer5_outputs(4543)) or (layer5_outputs(5752));
    layer6_outputs(985) <= not(layer5_outputs(2569)) or (layer5_outputs(5902));
    layer6_outputs(986) <= (layer5_outputs(5666)) xor (layer5_outputs(366));
    layer6_outputs(987) <= layer5_outputs(5393);
    layer6_outputs(988) <= not(layer5_outputs(700));
    layer6_outputs(989) <= layer5_outputs(5989);
    layer6_outputs(990) <= (layer5_outputs(1109)) and not (layer5_outputs(1202));
    layer6_outputs(991) <= not((layer5_outputs(6183)) or (layer5_outputs(662)));
    layer6_outputs(992) <= not(layer5_outputs(4178));
    layer6_outputs(993) <= not(layer5_outputs(2743));
    layer6_outputs(994) <= layer5_outputs(2788);
    layer6_outputs(995) <= not(layer5_outputs(5377));
    layer6_outputs(996) <= not(layer5_outputs(79));
    layer6_outputs(997) <= (layer5_outputs(36)) and not (layer5_outputs(922));
    layer6_outputs(998) <= layer5_outputs(1051);
    layer6_outputs(999) <= layer5_outputs(3127);
    layer6_outputs(1000) <= (layer5_outputs(1354)) and not (layer5_outputs(2270));
    layer6_outputs(1001) <= not((layer5_outputs(6689)) and (layer5_outputs(877)));
    layer6_outputs(1002) <= not((layer5_outputs(3357)) xor (layer5_outputs(6276)));
    layer6_outputs(1003) <= layer5_outputs(4815);
    layer6_outputs(1004) <= (layer5_outputs(2308)) and not (layer5_outputs(7302));
    layer6_outputs(1005) <= not(layer5_outputs(1797)) or (layer5_outputs(5287));
    layer6_outputs(1006) <= not(layer5_outputs(5697));
    layer6_outputs(1007) <= (layer5_outputs(6027)) and not (layer5_outputs(5304));
    layer6_outputs(1008) <= not((layer5_outputs(6100)) xor (layer5_outputs(4893)));
    layer6_outputs(1009) <= not(layer5_outputs(5958));
    layer6_outputs(1010) <= (layer5_outputs(6208)) xor (layer5_outputs(5271));
    layer6_outputs(1011) <= (layer5_outputs(1454)) and not (layer5_outputs(1000));
    layer6_outputs(1012) <= not(layer5_outputs(6978));
    layer6_outputs(1013) <= not(layer5_outputs(855));
    layer6_outputs(1014) <= not((layer5_outputs(5853)) and (layer5_outputs(5795)));
    layer6_outputs(1015) <= not(layer5_outputs(4339));
    layer6_outputs(1016) <= layer5_outputs(5510);
    layer6_outputs(1017) <= not(layer5_outputs(2385));
    layer6_outputs(1018) <= (layer5_outputs(5150)) and not (layer5_outputs(1110));
    layer6_outputs(1019) <= (layer5_outputs(3768)) and not (layer5_outputs(1608));
    layer6_outputs(1020) <= not(layer5_outputs(5217));
    layer6_outputs(1021) <= layer5_outputs(59);
    layer6_outputs(1022) <= not((layer5_outputs(6220)) or (layer5_outputs(2558)));
    layer6_outputs(1023) <= layer5_outputs(933);
    layer6_outputs(1024) <= (layer5_outputs(1073)) and not (layer5_outputs(3629));
    layer6_outputs(1025) <= layer5_outputs(7519);
    layer6_outputs(1026) <= not(layer5_outputs(7274)) or (layer5_outputs(214));
    layer6_outputs(1027) <= layer5_outputs(4803);
    layer6_outputs(1028) <= layer5_outputs(7026);
    layer6_outputs(1029) <= (layer5_outputs(281)) and not (layer5_outputs(4429));
    layer6_outputs(1030) <= not(layer5_outputs(4088)) or (layer5_outputs(4791));
    layer6_outputs(1031) <= layer5_outputs(7495);
    layer6_outputs(1032) <= (layer5_outputs(6136)) and not (layer5_outputs(7261));
    layer6_outputs(1033) <= not(layer5_outputs(2976));
    layer6_outputs(1034) <= layer5_outputs(6186);
    layer6_outputs(1035) <= (layer5_outputs(4668)) xor (layer5_outputs(5270));
    layer6_outputs(1036) <= (layer5_outputs(6840)) or (layer5_outputs(6235));
    layer6_outputs(1037) <= not(layer5_outputs(1780));
    layer6_outputs(1038) <= not(layer5_outputs(3042));
    layer6_outputs(1039) <= not(layer5_outputs(6478));
    layer6_outputs(1040) <= not(layer5_outputs(1869)) or (layer5_outputs(7539));
    layer6_outputs(1041) <= not((layer5_outputs(4758)) xor (layer5_outputs(3589)));
    layer6_outputs(1042) <= layer5_outputs(2812);
    layer6_outputs(1043) <= not(layer5_outputs(1739));
    layer6_outputs(1044) <= (layer5_outputs(4983)) xor (layer5_outputs(742));
    layer6_outputs(1045) <= (layer5_outputs(1644)) xor (layer5_outputs(2106));
    layer6_outputs(1046) <= not(layer5_outputs(317));
    layer6_outputs(1047) <= not(layer5_outputs(537));
    layer6_outputs(1048) <= not((layer5_outputs(4954)) or (layer5_outputs(3880)));
    layer6_outputs(1049) <= (layer5_outputs(7664)) and (layer5_outputs(7090));
    layer6_outputs(1050) <= layer5_outputs(2215);
    layer6_outputs(1051) <= not((layer5_outputs(2480)) or (layer5_outputs(3793)));
    layer6_outputs(1052) <= not(layer5_outputs(561));
    layer6_outputs(1053) <= layer5_outputs(4876);
    layer6_outputs(1054) <= not((layer5_outputs(3532)) and (layer5_outputs(6902)));
    layer6_outputs(1055) <= (layer5_outputs(490)) or (layer5_outputs(2069));
    layer6_outputs(1056) <= not(layer5_outputs(5548));
    layer6_outputs(1057) <= not(layer5_outputs(2335));
    layer6_outputs(1058) <= not((layer5_outputs(4606)) xor (layer5_outputs(1094)));
    layer6_outputs(1059) <= not((layer5_outputs(698)) and (layer5_outputs(7482)));
    layer6_outputs(1060) <= (layer5_outputs(545)) and not (layer5_outputs(5352));
    layer6_outputs(1061) <= (layer5_outputs(1257)) or (layer5_outputs(772));
    layer6_outputs(1062) <= not(layer5_outputs(1108));
    layer6_outputs(1063) <= (layer5_outputs(3851)) and not (layer5_outputs(7119));
    layer6_outputs(1064) <= (layer5_outputs(2045)) and (layer5_outputs(4604));
    layer6_outputs(1065) <= layer5_outputs(5098);
    layer6_outputs(1066) <= layer5_outputs(3103);
    layer6_outputs(1067) <= not(layer5_outputs(6096)) or (layer5_outputs(2641));
    layer6_outputs(1068) <= not((layer5_outputs(3761)) and (layer5_outputs(7588)));
    layer6_outputs(1069) <= not(layer5_outputs(5128));
    layer6_outputs(1070) <= (layer5_outputs(5208)) xor (layer5_outputs(337));
    layer6_outputs(1071) <= (layer5_outputs(1949)) or (layer5_outputs(7088));
    layer6_outputs(1072) <= layer5_outputs(1097);
    layer6_outputs(1073) <= (layer5_outputs(5712)) or (layer5_outputs(5132));
    layer6_outputs(1074) <= not(layer5_outputs(2039));
    layer6_outputs(1075) <= layer5_outputs(3872);
    layer6_outputs(1076) <= layer5_outputs(387);
    layer6_outputs(1077) <= (layer5_outputs(6690)) and (layer5_outputs(6839));
    layer6_outputs(1078) <= layer5_outputs(5043);
    layer6_outputs(1079) <= layer5_outputs(495);
    layer6_outputs(1080) <= (layer5_outputs(2377)) and (layer5_outputs(1426));
    layer6_outputs(1081) <= (layer5_outputs(974)) and not (layer5_outputs(4905));
    layer6_outputs(1082) <= layer5_outputs(3585);
    layer6_outputs(1083) <= not(layer5_outputs(7228));
    layer6_outputs(1084) <= not((layer5_outputs(4207)) xor (layer5_outputs(5819)));
    layer6_outputs(1085) <= (layer5_outputs(4585)) and not (layer5_outputs(331));
    layer6_outputs(1086) <= not(layer5_outputs(7281));
    layer6_outputs(1087) <= (layer5_outputs(3703)) or (layer5_outputs(7400));
    layer6_outputs(1088) <= layer5_outputs(2357);
    layer6_outputs(1089) <= not(layer5_outputs(4515)) or (layer5_outputs(5486));
    layer6_outputs(1090) <= not(layer5_outputs(5755));
    layer6_outputs(1091) <= layer5_outputs(6722);
    layer6_outputs(1092) <= (layer5_outputs(6650)) and not (layer5_outputs(4027));
    layer6_outputs(1093) <= not((layer5_outputs(582)) or (layer5_outputs(760)));
    layer6_outputs(1094) <= layer5_outputs(4358);
    layer6_outputs(1095) <= layer5_outputs(4566);
    layer6_outputs(1096) <= layer5_outputs(6627);
    layer6_outputs(1097) <= (layer5_outputs(2935)) or (layer5_outputs(4365));
    layer6_outputs(1098) <= (layer5_outputs(1977)) xor (layer5_outputs(1918));
    layer6_outputs(1099) <= layer5_outputs(4187);
    layer6_outputs(1100) <= not(layer5_outputs(1568));
    layer6_outputs(1101) <= layer5_outputs(4433);
    layer6_outputs(1102) <= not((layer5_outputs(3369)) or (layer5_outputs(7122)));
    layer6_outputs(1103) <= layer5_outputs(4900);
    layer6_outputs(1104) <= not(layer5_outputs(5253));
    layer6_outputs(1105) <= layer5_outputs(6179);
    layer6_outputs(1106) <= (layer5_outputs(7292)) xor (layer5_outputs(2012));
    layer6_outputs(1107) <= (layer5_outputs(6917)) and not (layer5_outputs(584));
    layer6_outputs(1108) <= layer5_outputs(5141);
    layer6_outputs(1109) <= not(layer5_outputs(6944)) or (layer5_outputs(6370));
    layer6_outputs(1110) <= not(layer5_outputs(2230));
    layer6_outputs(1111) <= (layer5_outputs(2829)) xor (layer5_outputs(994));
    layer6_outputs(1112) <= layer5_outputs(787);
    layer6_outputs(1113) <= not(layer5_outputs(296));
    layer6_outputs(1114) <= not(layer5_outputs(6867));
    layer6_outputs(1115) <= not(layer5_outputs(1162));
    layer6_outputs(1116) <= not((layer5_outputs(6458)) or (layer5_outputs(6825)));
    layer6_outputs(1117) <= layer5_outputs(109);
    layer6_outputs(1118) <= (layer5_outputs(5077)) xor (layer5_outputs(5046));
    layer6_outputs(1119) <= (layer5_outputs(2361)) and not (layer5_outputs(4301));
    layer6_outputs(1120) <= layer5_outputs(6599);
    layer6_outputs(1121) <= (layer5_outputs(4568)) and (layer5_outputs(3958));
    layer6_outputs(1122) <= layer5_outputs(7420);
    layer6_outputs(1123) <= (layer5_outputs(732)) and not (layer5_outputs(6731));
    layer6_outputs(1124) <= not(layer5_outputs(5700));
    layer6_outputs(1125) <= not(layer5_outputs(6970)) or (layer5_outputs(2054));
    layer6_outputs(1126) <= layer5_outputs(6036);
    layer6_outputs(1127) <= not(layer5_outputs(466));
    layer6_outputs(1128) <= layer5_outputs(5081);
    layer6_outputs(1129) <= not(layer5_outputs(4226));
    layer6_outputs(1130) <= layer5_outputs(6632);
    layer6_outputs(1131) <= not(layer5_outputs(508)) or (layer5_outputs(3612));
    layer6_outputs(1132) <= layer5_outputs(1807);
    layer6_outputs(1133) <= (layer5_outputs(356)) xor (layer5_outputs(6149));
    layer6_outputs(1134) <= layer5_outputs(7548);
    layer6_outputs(1135) <= not(layer5_outputs(7216));
    layer6_outputs(1136) <= layer5_outputs(4641);
    layer6_outputs(1137) <= not(layer5_outputs(5522));
    layer6_outputs(1138) <= '0';
    layer6_outputs(1139) <= not((layer5_outputs(2667)) and (layer5_outputs(7545)));
    layer6_outputs(1140) <= layer5_outputs(6036);
    layer6_outputs(1141) <= layer5_outputs(2129);
    layer6_outputs(1142) <= layer5_outputs(2783);
    layer6_outputs(1143) <= layer5_outputs(3435);
    layer6_outputs(1144) <= not(layer5_outputs(501));
    layer6_outputs(1145) <= (layer5_outputs(3207)) xor (layer5_outputs(5567));
    layer6_outputs(1146) <= not(layer5_outputs(5667));
    layer6_outputs(1147) <= not(layer5_outputs(2335));
    layer6_outputs(1148) <= layer5_outputs(1484);
    layer6_outputs(1149) <= (layer5_outputs(1753)) and not (layer5_outputs(3940));
    layer6_outputs(1150) <= layer5_outputs(1023);
    layer6_outputs(1151) <= not(layer5_outputs(2454));
    layer6_outputs(1152) <= not(layer5_outputs(0));
    layer6_outputs(1153) <= not((layer5_outputs(4956)) xor (layer5_outputs(2110)));
    layer6_outputs(1154) <= not((layer5_outputs(7667)) xor (layer5_outputs(5119)));
    layer6_outputs(1155) <= (layer5_outputs(3191)) or (layer5_outputs(3388));
    layer6_outputs(1156) <= (layer5_outputs(6019)) or (layer5_outputs(6466));
    layer6_outputs(1157) <= not(layer5_outputs(2390));
    layer6_outputs(1158) <= not((layer5_outputs(565)) and (layer5_outputs(6663)));
    layer6_outputs(1159) <= not(layer5_outputs(1022));
    layer6_outputs(1160) <= layer5_outputs(1141);
    layer6_outputs(1161) <= layer5_outputs(5127);
    layer6_outputs(1162) <= not((layer5_outputs(4146)) and (layer5_outputs(7149)));
    layer6_outputs(1163) <= (layer5_outputs(4108)) and (layer5_outputs(4445));
    layer6_outputs(1164) <= (layer5_outputs(2518)) and not (layer5_outputs(5933));
    layer6_outputs(1165) <= not(layer5_outputs(4142)) or (layer5_outputs(3857));
    layer6_outputs(1166) <= not(layer5_outputs(2225));
    layer6_outputs(1167) <= not(layer5_outputs(2426));
    layer6_outputs(1168) <= not((layer5_outputs(6521)) or (layer5_outputs(6010)));
    layer6_outputs(1169) <= not(layer5_outputs(6859));
    layer6_outputs(1170) <= layer5_outputs(6872);
    layer6_outputs(1171) <= (layer5_outputs(6912)) xor (layer5_outputs(7392));
    layer6_outputs(1172) <= (layer5_outputs(715)) and not (layer5_outputs(5479));
    layer6_outputs(1173) <= not((layer5_outputs(6318)) xor (layer5_outputs(3650)));
    layer6_outputs(1174) <= (layer5_outputs(664)) xor (layer5_outputs(2565));
    layer6_outputs(1175) <= layer5_outputs(5963);
    layer6_outputs(1176) <= not((layer5_outputs(288)) and (layer5_outputs(5844)));
    layer6_outputs(1177) <= layer5_outputs(1572);
    layer6_outputs(1178) <= (layer5_outputs(5381)) xor (layer5_outputs(4856));
    layer6_outputs(1179) <= (layer5_outputs(109)) and not (layer5_outputs(7576));
    layer6_outputs(1180) <= not((layer5_outputs(6949)) xor (layer5_outputs(7170)));
    layer6_outputs(1181) <= layer5_outputs(750);
    layer6_outputs(1182) <= not(layer5_outputs(1347));
    layer6_outputs(1183) <= layer5_outputs(5340);
    layer6_outputs(1184) <= layer5_outputs(7644);
    layer6_outputs(1185) <= not((layer5_outputs(2822)) or (layer5_outputs(5574)));
    layer6_outputs(1186) <= not((layer5_outputs(5809)) xor (layer5_outputs(6035)));
    layer6_outputs(1187) <= not(layer5_outputs(6270)) or (layer5_outputs(1772));
    layer6_outputs(1188) <= not(layer5_outputs(1592));
    layer6_outputs(1189) <= (layer5_outputs(1119)) xor (layer5_outputs(2593));
    layer6_outputs(1190) <= not(layer5_outputs(4905)) or (layer5_outputs(6014));
    layer6_outputs(1191) <= not(layer5_outputs(1892));
    layer6_outputs(1192) <= layer5_outputs(676);
    layer6_outputs(1193) <= not(layer5_outputs(789));
    layer6_outputs(1194) <= (layer5_outputs(677)) xor (layer5_outputs(4920));
    layer6_outputs(1195) <= layer5_outputs(5765);
    layer6_outputs(1196) <= layer5_outputs(7561);
    layer6_outputs(1197) <= not((layer5_outputs(4322)) and (layer5_outputs(4092)));
    layer6_outputs(1198) <= not(layer5_outputs(6267)) or (layer5_outputs(2633));
    layer6_outputs(1199) <= not((layer5_outputs(2441)) or (layer5_outputs(6604)));
    layer6_outputs(1200) <= (layer5_outputs(1545)) and (layer5_outputs(3003));
    layer6_outputs(1201) <= not((layer5_outputs(717)) xor (layer5_outputs(5025)));
    layer6_outputs(1202) <= not((layer5_outputs(7334)) xor (layer5_outputs(3501)));
    layer6_outputs(1203) <= not((layer5_outputs(1182)) xor (layer5_outputs(2972)));
    layer6_outputs(1204) <= not(layer5_outputs(1814)) or (layer5_outputs(3712));
    layer6_outputs(1205) <= not((layer5_outputs(2703)) or (layer5_outputs(286)));
    layer6_outputs(1206) <= layer5_outputs(2024);
    layer6_outputs(1207) <= layer5_outputs(366);
    layer6_outputs(1208) <= layer5_outputs(6280);
    layer6_outputs(1209) <= not(layer5_outputs(6623));
    layer6_outputs(1210) <= layer5_outputs(3706);
    layer6_outputs(1211) <= not(layer5_outputs(370));
    layer6_outputs(1212) <= not(layer5_outputs(531));
    layer6_outputs(1213) <= not(layer5_outputs(4940));
    layer6_outputs(1214) <= not(layer5_outputs(2685));
    layer6_outputs(1215) <= not(layer5_outputs(485));
    layer6_outputs(1216) <= layer5_outputs(4592);
    layer6_outputs(1217) <= (layer5_outputs(1842)) and (layer5_outputs(710));
    layer6_outputs(1218) <= not(layer5_outputs(7078));
    layer6_outputs(1219) <= layer5_outputs(6418);
    layer6_outputs(1220) <= not(layer5_outputs(5615));
    layer6_outputs(1221) <= (layer5_outputs(6894)) and not (layer5_outputs(7566));
    layer6_outputs(1222) <= not((layer5_outputs(1765)) xor (layer5_outputs(4395)));
    layer6_outputs(1223) <= not((layer5_outputs(6280)) xor (layer5_outputs(4544)));
    layer6_outputs(1224) <= layer5_outputs(335);
    layer6_outputs(1225) <= (layer5_outputs(1473)) xor (layer5_outputs(2239));
    layer6_outputs(1226) <= layer5_outputs(1490);
    layer6_outputs(1227) <= not(layer5_outputs(7249));
    layer6_outputs(1228) <= layer5_outputs(1171);
    layer6_outputs(1229) <= not(layer5_outputs(3849)) or (layer5_outputs(5214));
    layer6_outputs(1230) <= not(layer5_outputs(5827));
    layer6_outputs(1231) <= not(layer5_outputs(4483));
    layer6_outputs(1232) <= (layer5_outputs(5060)) xor (layer5_outputs(4929));
    layer6_outputs(1233) <= not((layer5_outputs(4256)) xor (layer5_outputs(1707)));
    layer6_outputs(1234) <= not(layer5_outputs(6173));
    layer6_outputs(1235) <= layer5_outputs(6226);
    layer6_outputs(1236) <= (layer5_outputs(2632)) xor (layer5_outputs(2262));
    layer6_outputs(1237) <= layer5_outputs(4249);
    layer6_outputs(1238) <= not(layer5_outputs(2004));
    layer6_outputs(1239) <= not(layer5_outputs(5905));
    layer6_outputs(1240) <= (layer5_outputs(4737)) and not (layer5_outputs(3635));
    layer6_outputs(1241) <= layer5_outputs(1244);
    layer6_outputs(1242) <= not((layer5_outputs(7579)) and (layer5_outputs(4575)));
    layer6_outputs(1243) <= not(layer5_outputs(5598)) or (layer5_outputs(277));
    layer6_outputs(1244) <= not(layer5_outputs(3339));
    layer6_outputs(1245) <= (layer5_outputs(1608)) or (layer5_outputs(2166));
    layer6_outputs(1246) <= not(layer5_outputs(2988));
    layer6_outputs(1247) <= (layer5_outputs(4570)) xor (layer5_outputs(3984));
    layer6_outputs(1248) <= layer5_outputs(2376);
    layer6_outputs(1249) <= not(layer5_outputs(4706));
    layer6_outputs(1250) <= not(layer5_outputs(5515)) or (layer5_outputs(4251));
    layer6_outputs(1251) <= not((layer5_outputs(5789)) xor (layer5_outputs(1637)));
    layer6_outputs(1252) <= (layer5_outputs(6666)) xor (layer5_outputs(2625));
    layer6_outputs(1253) <= (layer5_outputs(1209)) xor (layer5_outputs(115));
    layer6_outputs(1254) <= layer5_outputs(4577);
    layer6_outputs(1255) <= not(layer5_outputs(3965));
    layer6_outputs(1256) <= layer5_outputs(5036);
    layer6_outputs(1257) <= not(layer5_outputs(6789)) or (layer5_outputs(1581));
    layer6_outputs(1258) <= layer5_outputs(3147);
    layer6_outputs(1259) <= (layer5_outputs(3533)) xor (layer5_outputs(5708));
    layer6_outputs(1260) <= (layer5_outputs(4582)) xor (layer5_outputs(5706));
    layer6_outputs(1261) <= not(layer5_outputs(2278));
    layer6_outputs(1262) <= layer5_outputs(5551);
    layer6_outputs(1263) <= (layer5_outputs(6342)) xor (layer5_outputs(1536));
    layer6_outputs(1264) <= layer5_outputs(7617);
    layer6_outputs(1265) <= not(layer5_outputs(626));
    layer6_outputs(1266) <= (layer5_outputs(3155)) and (layer5_outputs(4942));
    layer6_outputs(1267) <= layer5_outputs(5291);
    layer6_outputs(1268) <= not(layer5_outputs(1724)) or (layer5_outputs(4550));
    layer6_outputs(1269) <= (layer5_outputs(4644)) or (layer5_outputs(5297));
    layer6_outputs(1270) <= layer5_outputs(2599);
    layer6_outputs(1271) <= layer5_outputs(6513);
    layer6_outputs(1272) <= layer5_outputs(4211);
    layer6_outputs(1273) <= not(layer5_outputs(2848));
    layer6_outputs(1274) <= not(layer5_outputs(4104));
    layer6_outputs(1275) <= (layer5_outputs(6447)) xor (layer5_outputs(4491));
    layer6_outputs(1276) <= (layer5_outputs(946)) and (layer5_outputs(5317));
    layer6_outputs(1277) <= (layer5_outputs(896)) xor (layer5_outputs(4615));
    layer6_outputs(1278) <= (layer5_outputs(1260)) xor (layer5_outputs(2986));
    layer6_outputs(1279) <= (layer5_outputs(5151)) and not (layer5_outputs(6207));
    layer6_outputs(1280) <= (layer5_outputs(3580)) and (layer5_outputs(819));
    layer6_outputs(1281) <= not((layer5_outputs(2882)) or (layer5_outputs(5592)));
    layer6_outputs(1282) <= layer5_outputs(5103);
    layer6_outputs(1283) <= '0';
    layer6_outputs(1284) <= not(layer5_outputs(1993));
    layer6_outputs(1285) <= layer5_outputs(3325);
    layer6_outputs(1286) <= not(layer5_outputs(5777));
    layer6_outputs(1287) <= not(layer5_outputs(5184));
    layer6_outputs(1288) <= layer5_outputs(6701);
    layer6_outputs(1289) <= not(layer5_outputs(5931));
    layer6_outputs(1290) <= layer5_outputs(2468);
    layer6_outputs(1291) <= not(layer5_outputs(5711)) or (layer5_outputs(255));
    layer6_outputs(1292) <= not(layer5_outputs(7059));
    layer6_outputs(1293) <= layer5_outputs(4655);
    layer6_outputs(1294) <= layer5_outputs(4324);
    layer6_outputs(1295) <= not(layer5_outputs(1288));
    layer6_outputs(1296) <= (layer5_outputs(4567)) xor (layer5_outputs(7614));
    layer6_outputs(1297) <= layer5_outputs(2009);
    layer6_outputs(1298) <= not(layer5_outputs(4581)) or (layer5_outputs(94));
    layer6_outputs(1299) <= layer5_outputs(1539);
    layer6_outputs(1300) <= not(layer5_outputs(2199));
    layer6_outputs(1301) <= layer5_outputs(3976);
    layer6_outputs(1302) <= not((layer5_outputs(1279)) or (layer5_outputs(3254)));
    layer6_outputs(1303) <= '1';
    layer6_outputs(1304) <= not(layer5_outputs(6961));
    layer6_outputs(1305) <= layer5_outputs(2194);
    layer6_outputs(1306) <= not(layer5_outputs(3586));
    layer6_outputs(1307) <= layer5_outputs(2709);
    layer6_outputs(1308) <= not(layer5_outputs(4927)) or (layer5_outputs(173));
    layer6_outputs(1309) <= (layer5_outputs(3230)) xor (layer5_outputs(2082));
    layer6_outputs(1310) <= not((layer5_outputs(5364)) and (layer5_outputs(4854)));
    layer6_outputs(1311) <= layer5_outputs(5520);
    layer6_outputs(1312) <= not((layer5_outputs(3238)) or (layer5_outputs(4923)));
    layer6_outputs(1313) <= (layer5_outputs(4706)) or (layer5_outputs(1136));
    layer6_outputs(1314) <= (layer5_outputs(3746)) and not (layer5_outputs(2245));
    layer6_outputs(1315) <= not(layer5_outputs(6786));
    layer6_outputs(1316) <= not(layer5_outputs(7237));
    layer6_outputs(1317) <= (layer5_outputs(287)) and (layer5_outputs(6561));
    layer6_outputs(1318) <= layer5_outputs(1998);
    layer6_outputs(1319) <= layer5_outputs(2800);
    layer6_outputs(1320) <= not(layer5_outputs(5120));
    layer6_outputs(1321) <= not(layer5_outputs(3862));
    layer6_outputs(1322) <= layer5_outputs(4745);
    layer6_outputs(1323) <= not(layer5_outputs(6887));
    layer6_outputs(1324) <= not(layer5_outputs(6125)) or (layer5_outputs(1817));
    layer6_outputs(1325) <= not(layer5_outputs(2698));
    layer6_outputs(1326) <= not(layer5_outputs(460));
    layer6_outputs(1327) <= not((layer5_outputs(51)) or (layer5_outputs(2077)));
    layer6_outputs(1328) <= layer5_outputs(4362);
    layer6_outputs(1329) <= not(layer5_outputs(2999));
    layer6_outputs(1330) <= layer5_outputs(1537);
    layer6_outputs(1331) <= not(layer5_outputs(1800));
    layer6_outputs(1332) <= not((layer5_outputs(2590)) and (layer5_outputs(3418)));
    layer6_outputs(1333) <= layer5_outputs(3447);
    layer6_outputs(1334) <= not(layer5_outputs(4188));
    layer6_outputs(1335) <= layer5_outputs(3085);
    layer6_outputs(1336) <= not((layer5_outputs(6415)) xor (layer5_outputs(2718)));
    layer6_outputs(1337) <= not((layer5_outputs(5664)) and (layer5_outputs(3188)));
    layer6_outputs(1338) <= not(layer5_outputs(3747)) or (layer5_outputs(3539));
    layer6_outputs(1339) <= layer5_outputs(4866);
    layer6_outputs(1340) <= not((layer5_outputs(3008)) xor (layer5_outputs(3572)));
    layer6_outputs(1341) <= layer5_outputs(5286);
    layer6_outputs(1342) <= not(layer5_outputs(4954));
    layer6_outputs(1343) <= layer5_outputs(6580);
    layer6_outputs(1344) <= layer5_outputs(6523);
    layer6_outputs(1345) <= not((layer5_outputs(7303)) and (layer5_outputs(2112)));
    layer6_outputs(1346) <= layer5_outputs(1132);
    layer6_outputs(1347) <= not((layer5_outputs(1577)) xor (layer5_outputs(693)));
    layer6_outputs(1348) <= not((layer5_outputs(2732)) or (layer5_outputs(2651)));
    layer6_outputs(1349) <= not(layer5_outputs(6707));
    layer6_outputs(1350) <= layer5_outputs(4109);
    layer6_outputs(1351) <= not((layer5_outputs(558)) xor (layer5_outputs(3993)));
    layer6_outputs(1352) <= layer5_outputs(2910);
    layer6_outputs(1353) <= (layer5_outputs(6618)) xor (layer5_outputs(1483));
    layer6_outputs(1354) <= not(layer5_outputs(2152));
    layer6_outputs(1355) <= layer5_outputs(2704);
    layer6_outputs(1356) <= not(layer5_outputs(2774));
    layer6_outputs(1357) <= layer5_outputs(2121);
    layer6_outputs(1358) <= not(layer5_outputs(2531));
    layer6_outputs(1359) <= not(layer5_outputs(1016));
    layer6_outputs(1360) <= not((layer5_outputs(1695)) xor (layer5_outputs(1593)));
    layer6_outputs(1361) <= not(layer5_outputs(1500));
    layer6_outputs(1362) <= layer5_outputs(289);
    layer6_outputs(1363) <= layer5_outputs(3548);
    layer6_outputs(1364) <= not(layer5_outputs(94)) or (layer5_outputs(4618));
    layer6_outputs(1365) <= not(layer5_outputs(6217)) or (layer5_outputs(2745));
    layer6_outputs(1366) <= layer5_outputs(3345);
    layer6_outputs(1367) <= layer5_outputs(6277);
    layer6_outputs(1368) <= layer5_outputs(5508);
    layer6_outputs(1369) <= (layer5_outputs(4446)) xor (layer5_outputs(658));
    layer6_outputs(1370) <= not(layer5_outputs(4306));
    layer6_outputs(1371) <= (layer5_outputs(1890)) xor (layer5_outputs(3927));
    layer6_outputs(1372) <= layer5_outputs(6678);
    layer6_outputs(1373) <= not((layer5_outputs(1003)) or (layer5_outputs(5012)));
    layer6_outputs(1374) <= not(layer5_outputs(2058)) or (layer5_outputs(5307));
    layer6_outputs(1375) <= (layer5_outputs(715)) xor (layer5_outputs(5236));
    layer6_outputs(1376) <= (layer5_outputs(1318)) and (layer5_outputs(4159));
    layer6_outputs(1377) <= '1';
    layer6_outputs(1378) <= not(layer5_outputs(5264));
    layer6_outputs(1379) <= layer5_outputs(3884);
    layer6_outputs(1380) <= not(layer5_outputs(1389));
    layer6_outputs(1381) <= layer5_outputs(2554);
    layer6_outputs(1382) <= layer5_outputs(6739);
    layer6_outputs(1383) <= not((layer5_outputs(1300)) xor (layer5_outputs(2399)));
    layer6_outputs(1384) <= not(layer5_outputs(3487));
    layer6_outputs(1385) <= not(layer5_outputs(1192));
    layer6_outputs(1386) <= layer5_outputs(4071);
    layer6_outputs(1387) <= not((layer5_outputs(5523)) and (layer5_outputs(5929)));
    layer6_outputs(1388) <= (layer5_outputs(3235)) and (layer5_outputs(1234));
    layer6_outputs(1389) <= not(layer5_outputs(4617)) or (layer5_outputs(2625));
    layer6_outputs(1390) <= not(layer5_outputs(1941));
    layer6_outputs(1391) <= not((layer5_outputs(4085)) or (layer5_outputs(3882)));
    layer6_outputs(1392) <= not((layer5_outputs(4008)) xor (layer5_outputs(2081)));
    layer6_outputs(1393) <= not(layer5_outputs(2795)) or (layer5_outputs(2449));
    layer6_outputs(1394) <= not(layer5_outputs(2522));
    layer6_outputs(1395) <= layer5_outputs(2759);
    layer6_outputs(1396) <= (layer5_outputs(6916)) or (layer5_outputs(4683));
    layer6_outputs(1397) <= layer5_outputs(1424);
    layer6_outputs(1398) <= not((layer5_outputs(4939)) xor (layer5_outputs(3853)));
    layer6_outputs(1399) <= layer5_outputs(2118);
    layer6_outputs(1400) <= not((layer5_outputs(6614)) xor (layer5_outputs(226)));
    layer6_outputs(1401) <= not(layer5_outputs(638));
    layer6_outputs(1402) <= not(layer5_outputs(13));
    layer6_outputs(1403) <= (layer5_outputs(2811)) and (layer5_outputs(7614));
    layer6_outputs(1404) <= not((layer5_outputs(6998)) xor (layer5_outputs(2224)));
    layer6_outputs(1405) <= not(layer5_outputs(5453));
    layer6_outputs(1406) <= not(layer5_outputs(7246));
    layer6_outputs(1407) <= layer5_outputs(1360);
    layer6_outputs(1408) <= not(layer5_outputs(6076)) or (layer5_outputs(6159));
    layer6_outputs(1409) <= not((layer5_outputs(5983)) xor (layer5_outputs(188)));
    layer6_outputs(1410) <= layer5_outputs(2594);
    layer6_outputs(1411) <= (layer5_outputs(5423)) xor (layer5_outputs(346));
    layer6_outputs(1412) <= layer5_outputs(5416);
    layer6_outputs(1413) <= not((layer5_outputs(2676)) xor (layer5_outputs(1445)));
    layer6_outputs(1414) <= not((layer5_outputs(1699)) xor (layer5_outputs(3511)));
    layer6_outputs(1415) <= not(layer5_outputs(2885));
    layer6_outputs(1416) <= layer5_outputs(2463);
    layer6_outputs(1417) <= layer5_outputs(6247);
    layer6_outputs(1418) <= not(layer5_outputs(5493));
    layer6_outputs(1419) <= layer5_outputs(6788);
    layer6_outputs(1420) <= not((layer5_outputs(7605)) and (layer5_outputs(229)));
    layer6_outputs(1421) <= not(layer5_outputs(7561));
    layer6_outputs(1422) <= layer5_outputs(3998);
    layer6_outputs(1423) <= not(layer5_outputs(3360));
    layer6_outputs(1424) <= not(layer5_outputs(1743));
    layer6_outputs(1425) <= not(layer5_outputs(6499)) or (layer5_outputs(3951));
    layer6_outputs(1426) <= not(layer5_outputs(4772)) or (layer5_outputs(3189));
    layer6_outputs(1427) <= not(layer5_outputs(3971));
    layer6_outputs(1428) <= (layer5_outputs(4808)) xor (layer5_outputs(2182));
    layer6_outputs(1429) <= not((layer5_outputs(5515)) xor (layer5_outputs(2951)));
    layer6_outputs(1430) <= layer5_outputs(7428);
    layer6_outputs(1431) <= layer5_outputs(7460);
    layer6_outputs(1432) <= not(layer5_outputs(3411));
    layer6_outputs(1433) <= not((layer5_outputs(5578)) xor (layer5_outputs(3130)));
    layer6_outputs(1434) <= not(layer5_outputs(4279));
    layer6_outputs(1435) <= layer5_outputs(3237);
    layer6_outputs(1436) <= not((layer5_outputs(1822)) xor (layer5_outputs(4982)));
    layer6_outputs(1437) <= layer5_outputs(777);
    layer6_outputs(1438) <= not(layer5_outputs(3603));
    layer6_outputs(1439) <= layer5_outputs(6597);
    layer6_outputs(1440) <= layer5_outputs(1359);
    layer6_outputs(1441) <= not(layer5_outputs(4916));
    layer6_outputs(1442) <= not(layer5_outputs(3578));
    layer6_outputs(1443) <= layer5_outputs(4082);
    layer6_outputs(1444) <= '0';
    layer6_outputs(1445) <= (layer5_outputs(3279)) xor (layer5_outputs(1733));
    layer6_outputs(1446) <= layer5_outputs(5706);
    layer6_outputs(1447) <= (layer5_outputs(3210)) xor (layer5_outputs(3897));
    layer6_outputs(1448) <= layer5_outputs(1894);
    layer6_outputs(1449) <= not(layer5_outputs(7148));
    layer6_outputs(1450) <= not((layer5_outputs(1847)) and (layer5_outputs(943)));
    layer6_outputs(1451) <= not((layer5_outputs(2437)) xor (layer5_outputs(4834)));
    layer6_outputs(1452) <= layer5_outputs(7273);
    layer6_outputs(1453) <= not(layer5_outputs(7651));
    layer6_outputs(1454) <= layer5_outputs(3622);
    layer6_outputs(1455) <= not((layer5_outputs(5796)) and (layer5_outputs(237)));
    layer6_outputs(1456) <= layer5_outputs(3343);
    layer6_outputs(1457) <= not(layer5_outputs(4629));
    layer6_outputs(1458) <= layer5_outputs(2795);
    layer6_outputs(1459) <= not(layer5_outputs(1377));
    layer6_outputs(1460) <= not((layer5_outputs(5822)) xor (layer5_outputs(1246)));
    layer6_outputs(1461) <= not(layer5_outputs(5563));
    layer6_outputs(1462) <= layer5_outputs(6188);
    layer6_outputs(1463) <= not((layer5_outputs(7366)) xor (layer5_outputs(937)));
    layer6_outputs(1464) <= layer5_outputs(6059);
    layer6_outputs(1465) <= (layer5_outputs(4137)) xor (layer5_outputs(2117));
    layer6_outputs(1466) <= not(layer5_outputs(6202)) or (layer5_outputs(3306));
    layer6_outputs(1467) <= not((layer5_outputs(6467)) xor (layer5_outputs(3828)));
    layer6_outputs(1468) <= (layer5_outputs(6127)) xor (layer5_outputs(2788));
    layer6_outputs(1469) <= layer5_outputs(3223);
    layer6_outputs(1470) <= layer5_outputs(176);
    layer6_outputs(1471) <= layer5_outputs(3042);
    layer6_outputs(1472) <= not(layer5_outputs(1164));
    layer6_outputs(1473) <= layer5_outputs(2846);
    layer6_outputs(1474) <= not((layer5_outputs(7171)) and (layer5_outputs(3194)));
    layer6_outputs(1475) <= (layer5_outputs(2638)) and not (layer5_outputs(931));
    layer6_outputs(1476) <= not(layer5_outputs(4136)) or (layer5_outputs(1478));
    layer6_outputs(1477) <= (layer5_outputs(6827)) xor (layer5_outputs(2386));
    layer6_outputs(1478) <= (layer5_outputs(6163)) or (layer5_outputs(3591));
    layer6_outputs(1479) <= not(layer5_outputs(2090)) or (layer5_outputs(2725));
    layer6_outputs(1480) <= (layer5_outputs(2485)) and not (layer5_outputs(2608));
    layer6_outputs(1481) <= (layer5_outputs(5013)) and (layer5_outputs(7096));
    layer6_outputs(1482) <= not(layer5_outputs(2213));
    layer6_outputs(1483) <= not(layer5_outputs(6222));
    layer6_outputs(1484) <= layer5_outputs(3831);
    layer6_outputs(1485) <= not(layer5_outputs(339));
    layer6_outputs(1486) <= not(layer5_outputs(947));
    layer6_outputs(1487) <= not(layer5_outputs(6385));
    layer6_outputs(1488) <= layer5_outputs(1382);
    layer6_outputs(1489) <= (layer5_outputs(2863)) xor (layer5_outputs(725));
    layer6_outputs(1490) <= (layer5_outputs(6642)) or (layer5_outputs(4423));
    layer6_outputs(1491) <= layer5_outputs(6421);
    layer6_outputs(1492) <= layer5_outputs(7444);
    layer6_outputs(1493) <= not(layer5_outputs(890));
    layer6_outputs(1494) <= (layer5_outputs(2923)) or (layer5_outputs(2557));
    layer6_outputs(1495) <= not(layer5_outputs(1143));
    layer6_outputs(1496) <= layer5_outputs(4692);
    layer6_outputs(1497) <= not(layer5_outputs(6719));
    layer6_outputs(1498) <= not(layer5_outputs(4358));
    layer6_outputs(1499) <= layer5_outputs(7489);
    layer6_outputs(1500) <= layer5_outputs(4328);
    layer6_outputs(1501) <= not(layer5_outputs(5479));
    layer6_outputs(1502) <= layer5_outputs(5310);
    layer6_outputs(1503) <= not(layer5_outputs(3154));
    layer6_outputs(1504) <= not((layer5_outputs(3710)) or (layer5_outputs(6982)));
    layer6_outputs(1505) <= (layer5_outputs(5205)) xor (layer5_outputs(2046));
    layer6_outputs(1506) <= (layer5_outputs(289)) and (layer5_outputs(6783));
    layer6_outputs(1507) <= not(layer5_outputs(6301)) or (layer5_outputs(6546));
    layer6_outputs(1508) <= layer5_outputs(3335);
    layer6_outputs(1509) <= not(layer5_outputs(3109));
    layer6_outputs(1510) <= layer5_outputs(2706);
    layer6_outputs(1511) <= not(layer5_outputs(687));
    layer6_outputs(1512) <= (layer5_outputs(3845)) and not (layer5_outputs(4524));
    layer6_outputs(1513) <= (layer5_outputs(3701)) or (layer5_outputs(2038));
    layer6_outputs(1514) <= not((layer5_outputs(3577)) xor (layer5_outputs(3801)));
    layer6_outputs(1515) <= not((layer5_outputs(3064)) or (layer5_outputs(1102)));
    layer6_outputs(1516) <= layer5_outputs(4780);
    layer6_outputs(1517) <= (layer5_outputs(1511)) or (layer5_outputs(949));
    layer6_outputs(1518) <= not((layer5_outputs(546)) xor (layer5_outputs(1644)));
    layer6_outputs(1519) <= not(layer5_outputs(736)) or (layer5_outputs(5967));
    layer6_outputs(1520) <= (layer5_outputs(4761)) and not (layer5_outputs(3000));
    layer6_outputs(1521) <= not(layer5_outputs(6729));
    layer6_outputs(1522) <= (layer5_outputs(1329)) or (layer5_outputs(5312));
    layer6_outputs(1523) <= not(layer5_outputs(1751));
    layer6_outputs(1524) <= not(layer5_outputs(221)) or (layer5_outputs(1290));
    layer6_outputs(1525) <= not(layer5_outputs(1126)) or (layer5_outputs(3721));
    layer6_outputs(1526) <= not((layer5_outputs(647)) xor (layer5_outputs(3407)));
    layer6_outputs(1527) <= not(layer5_outputs(1373));
    layer6_outputs(1528) <= not(layer5_outputs(6481));
    layer6_outputs(1529) <= not(layer5_outputs(3367)) or (layer5_outputs(6291));
    layer6_outputs(1530) <= (layer5_outputs(4697)) or (layer5_outputs(1551));
    layer6_outputs(1531) <= (layer5_outputs(1924)) and not (layer5_outputs(1825));
    layer6_outputs(1532) <= layer5_outputs(4889);
    layer6_outputs(1533) <= not(layer5_outputs(2408));
    layer6_outputs(1534) <= not(layer5_outputs(1713));
    layer6_outputs(1535) <= layer5_outputs(720);
    layer6_outputs(1536) <= (layer5_outputs(5085)) and not (layer5_outputs(3444));
    layer6_outputs(1537) <= layer5_outputs(6603);
    layer6_outputs(1538) <= layer5_outputs(3785);
    layer6_outputs(1539) <= not((layer5_outputs(3821)) xor (layer5_outputs(7093)));
    layer6_outputs(1540) <= (layer5_outputs(1938)) and not (layer5_outputs(1648));
    layer6_outputs(1541) <= not(layer5_outputs(3293));
    layer6_outputs(1542) <= (layer5_outputs(2200)) or (layer5_outputs(1150));
    layer6_outputs(1543) <= not((layer5_outputs(6123)) xor (layer5_outputs(2889)));
    layer6_outputs(1544) <= not(layer5_outputs(4196)) or (layer5_outputs(5046));
    layer6_outputs(1545) <= not(layer5_outputs(7009));
    layer6_outputs(1546) <= layer5_outputs(5277);
    layer6_outputs(1547) <= not(layer5_outputs(3650));
    layer6_outputs(1548) <= not(layer5_outputs(5049));
    layer6_outputs(1549) <= not(layer5_outputs(7363));
    layer6_outputs(1550) <= layer5_outputs(772);
    layer6_outputs(1551) <= layer5_outputs(2301);
    layer6_outputs(1552) <= not((layer5_outputs(4538)) and (layer5_outputs(2660)));
    layer6_outputs(1553) <= layer5_outputs(1115);
    layer6_outputs(1554) <= not((layer5_outputs(622)) xor (layer5_outputs(2266)));
    layer6_outputs(1555) <= layer5_outputs(6257);
    layer6_outputs(1556) <= layer5_outputs(1544);
    layer6_outputs(1557) <= layer5_outputs(3470);
    layer6_outputs(1558) <= not((layer5_outputs(4240)) xor (layer5_outputs(6001)));
    layer6_outputs(1559) <= layer5_outputs(6575);
    layer6_outputs(1560) <= not(layer5_outputs(306));
    layer6_outputs(1561) <= layer5_outputs(966);
    layer6_outputs(1562) <= not(layer5_outputs(169));
    layer6_outputs(1563) <= layer5_outputs(1274);
    layer6_outputs(1564) <= not(layer5_outputs(7524));
    layer6_outputs(1565) <= (layer5_outputs(4690)) and not (layer5_outputs(7650));
    layer6_outputs(1566) <= (layer5_outputs(3930)) xor (layer5_outputs(3916));
    layer6_outputs(1567) <= not(layer5_outputs(4480));
    layer6_outputs(1568) <= layer5_outputs(6111);
    layer6_outputs(1569) <= layer5_outputs(5467);
    layer6_outputs(1570) <= layer5_outputs(242);
    layer6_outputs(1571) <= not(layer5_outputs(3461));
    layer6_outputs(1572) <= layer5_outputs(4531);
    layer6_outputs(1573) <= not(layer5_outputs(4021));
    layer6_outputs(1574) <= not((layer5_outputs(7636)) or (layer5_outputs(3568)));
    layer6_outputs(1575) <= not(layer5_outputs(5418));
    layer6_outputs(1576) <= layer5_outputs(2692);
    layer6_outputs(1577) <= layer5_outputs(1708);
    layer6_outputs(1578) <= (layer5_outputs(4743)) xor (layer5_outputs(6354));
    layer6_outputs(1579) <= not(layer5_outputs(7606));
    layer6_outputs(1580) <= not((layer5_outputs(6771)) xor (layer5_outputs(1028)));
    layer6_outputs(1581) <= (layer5_outputs(6657)) xor (layer5_outputs(4324));
    layer6_outputs(1582) <= not(layer5_outputs(4935));
    layer6_outputs(1583) <= not(layer5_outputs(3421));
    layer6_outputs(1584) <= not(layer5_outputs(1148));
    layer6_outputs(1585) <= not((layer5_outputs(1492)) xor (layer5_outputs(4084)));
    layer6_outputs(1586) <= not((layer5_outputs(5657)) xor (layer5_outputs(202)));
    layer6_outputs(1587) <= not((layer5_outputs(5484)) xor (layer5_outputs(2150)));
    layer6_outputs(1588) <= not((layer5_outputs(4191)) xor (layer5_outputs(4420)));
    layer6_outputs(1589) <= not((layer5_outputs(6495)) xor (layer5_outputs(1779)));
    layer6_outputs(1590) <= not((layer5_outputs(5417)) xor (layer5_outputs(5655)));
    layer6_outputs(1591) <= layer5_outputs(7144);
    layer6_outputs(1592) <= not(layer5_outputs(4884));
    layer6_outputs(1593) <= not(layer5_outputs(4151));
    layer6_outputs(1594) <= not(layer5_outputs(1340)) or (layer5_outputs(886));
    layer6_outputs(1595) <= not(layer5_outputs(6391));
    layer6_outputs(1596) <= layer5_outputs(6306);
    layer6_outputs(1597) <= (layer5_outputs(6294)) xor (layer5_outputs(552));
    layer6_outputs(1598) <= layer5_outputs(845);
    layer6_outputs(1599) <= layer5_outputs(2356);
    layer6_outputs(1600) <= layer5_outputs(3451);
    layer6_outputs(1601) <= layer5_outputs(5658);
    layer6_outputs(1602) <= layer5_outputs(2707);
    layer6_outputs(1603) <= layer5_outputs(4972);
    layer6_outputs(1604) <= (layer5_outputs(556)) and (layer5_outputs(4235));
    layer6_outputs(1605) <= layer5_outputs(6696);
    layer6_outputs(1606) <= (layer5_outputs(6070)) and not (layer5_outputs(5401));
    layer6_outputs(1607) <= not(layer5_outputs(6687)) or (layer5_outputs(6898));
    layer6_outputs(1608) <= (layer5_outputs(7048)) and not (layer5_outputs(3947));
    layer6_outputs(1609) <= not((layer5_outputs(3669)) xor (layer5_outputs(1821)));
    layer6_outputs(1610) <= (layer5_outputs(7135)) and not (layer5_outputs(1013));
    layer6_outputs(1611) <= not(layer5_outputs(6303));
    layer6_outputs(1612) <= layer5_outputs(3769);
    layer6_outputs(1613) <= (layer5_outputs(3539)) and not (layer5_outputs(5596));
    layer6_outputs(1614) <= layer5_outputs(3215);
    layer6_outputs(1615) <= not(layer5_outputs(6913)) or (layer5_outputs(2723));
    layer6_outputs(1616) <= layer5_outputs(5022);
    layer6_outputs(1617) <= not(layer5_outputs(1118));
    layer6_outputs(1618) <= not(layer5_outputs(5261)) or (layer5_outputs(3203));
    layer6_outputs(1619) <= (layer5_outputs(3034)) xor (layer5_outputs(636));
    layer6_outputs(1620) <= (layer5_outputs(1169)) xor (layer5_outputs(2155));
    layer6_outputs(1621) <= not(layer5_outputs(4449)) or (layer5_outputs(770));
    layer6_outputs(1622) <= (layer5_outputs(5386)) xor (layer5_outputs(6374));
    layer6_outputs(1623) <= layer5_outputs(3617);
    layer6_outputs(1624) <= not(layer5_outputs(5757));
    layer6_outputs(1625) <= (layer5_outputs(479)) and not (layer5_outputs(1653));
    layer6_outputs(1626) <= not((layer5_outputs(6183)) xor (layer5_outputs(591)));
    layer6_outputs(1627) <= not(layer5_outputs(2434));
    layer6_outputs(1628) <= (layer5_outputs(5195)) xor (layer5_outputs(637));
    layer6_outputs(1629) <= not(layer5_outputs(6045));
    layer6_outputs(1630) <= not(layer5_outputs(1327));
    layer6_outputs(1631) <= not(layer5_outputs(3708)) or (layer5_outputs(2247));
    layer6_outputs(1632) <= (layer5_outputs(1757)) and not (layer5_outputs(3481));
    layer6_outputs(1633) <= (layer5_outputs(297)) and not (layer5_outputs(7366));
    layer6_outputs(1634) <= not(layer5_outputs(2902));
    layer6_outputs(1635) <= not((layer5_outputs(3312)) or (layer5_outputs(6635)));
    layer6_outputs(1636) <= layer5_outputs(3722);
    layer6_outputs(1637) <= (layer5_outputs(6763)) and not (layer5_outputs(5395));
    layer6_outputs(1638) <= layer5_outputs(3628);
    layer6_outputs(1639) <= not((layer5_outputs(5188)) xor (layer5_outputs(4168)));
    layer6_outputs(1640) <= layer5_outputs(5577);
    layer6_outputs(1641) <= not((layer5_outputs(431)) or (layer5_outputs(3422)));
    layer6_outputs(1642) <= not(layer5_outputs(3061));
    layer6_outputs(1643) <= (layer5_outputs(2205)) and not (layer5_outputs(1498));
    layer6_outputs(1644) <= not(layer5_outputs(5453));
    layer6_outputs(1645) <= not(layer5_outputs(1496));
    layer6_outputs(1646) <= layer5_outputs(1948);
    layer6_outputs(1647) <= not(layer5_outputs(5485));
    layer6_outputs(1648) <= (layer5_outputs(1429)) xor (layer5_outputs(5341));
    layer6_outputs(1649) <= not(layer5_outputs(2436));
    layer6_outputs(1650) <= (layer5_outputs(1879)) xor (layer5_outputs(5136));
    layer6_outputs(1651) <= not(layer5_outputs(6557)) or (layer5_outputs(3752));
    layer6_outputs(1652) <= layer5_outputs(3792);
    layer6_outputs(1653) <= '1';
    layer6_outputs(1654) <= layer5_outputs(5307);
    layer6_outputs(1655) <= not(layer5_outputs(2471));
    layer6_outputs(1656) <= not(layer5_outputs(7279));
    layer6_outputs(1657) <= not(layer5_outputs(2326));
    layer6_outputs(1658) <= (layer5_outputs(3552)) xor (layer5_outputs(4779));
    layer6_outputs(1659) <= layer5_outputs(7487);
    layer6_outputs(1660) <= '1';
    layer6_outputs(1661) <= not(layer5_outputs(4704)) or (layer5_outputs(575));
    layer6_outputs(1662) <= (layer5_outputs(4434)) and not (layer5_outputs(4307));
    layer6_outputs(1663) <= (layer5_outputs(5392)) and (layer5_outputs(1251));
    layer6_outputs(1664) <= layer5_outputs(208);
    layer6_outputs(1665) <= not(layer5_outputs(1552));
    layer6_outputs(1666) <= layer5_outputs(4871);
    layer6_outputs(1667) <= not(layer5_outputs(2511));
    layer6_outputs(1668) <= not(layer5_outputs(1559));
    layer6_outputs(1669) <= layer5_outputs(5717);
    layer6_outputs(1670) <= not(layer5_outputs(5888));
    layer6_outputs(1671) <= not((layer5_outputs(2114)) xor (layer5_outputs(2480)));
    layer6_outputs(1672) <= layer5_outputs(1272);
    layer6_outputs(1673) <= not((layer5_outputs(1921)) xor (layer5_outputs(344)));
    layer6_outputs(1674) <= layer5_outputs(3347);
    layer6_outputs(1675) <= layer5_outputs(5070);
    layer6_outputs(1676) <= not(layer5_outputs(5504)) or (layer5_outputs(3986));
    layer6_outputs(1677) <= layer5_outputs(1581);
    layer6_outputs(1678) <= layer5_outputs(6996);
    layer6_outputs(1679) <= (layer5_outputs(3146)) and not (layer5_outputs(5371));
    layer6_outputs(1680) <= not((layer5_outputs(1858)) and (layer5_outputs(904)));
    layer6_outputs(1681) <= layer5_outputs(7295);
    layer6_outputs(1682) <= not(layer5_outputs(3263));
    layer6_outputs(1683) <= not((layer5_outputs(3327)) or (layer5_outputs(3717)));
    layer6_outputs(1684) <= '0';
    layer6_outputs(1685) <= not(layer5_outputs(6753));
    layer6_outputs(1686) <= not((layer5_outputs(3449)) xor (layer5_outputs(4234)));
    layer6_outputs(1687) <= layer5_outputs(2031);
    layer6_outputs(1688) <= layer5_outputs(6745);
    layer6_outputs(1689) <= layer5_outputs(4135);
    layer6_outputs(1690) <= not(layer5_outputs(1548));
    layer6_outputs(1691) <= layer5_outputs(5032);
    layer6_outputs(1692) <= not(layer5_outputs(1285));
    layer6_outputs(1693) <= not(layer5_outputs(7504));
    layer6_outputs(1694) <= (layer5_outputs(5788)) or (layer5_outputs(5058));
    layer6_outputs(1695) <= not(layer5_outputs(5576)) or (layer5_outputs(4057));
    layer6_outputs(1696) <= not((layer5_outputs(6957)) xor (layer5_outputs(7303)));
    layer6_outputs(1697) <= (layer5_outputs(6890)) and not (layer5_outputs(4409));
    layer6_outputs(1698) <= not(layer5_outputs(3588));
    layer6_outputs(1699) <= not((layer5_outputs(525)) xor (layer5_outputs(1779)));
    layer6_outputs(1700) <= layer5_outputs(2646);
    layer6_outputs(1701) <= (layer5_outputs(1172)) and not (layer5_outputs(3800));
    layer6_outputs(1702) <= not(layer5_outputs(4336));
    layer6_outputs(1703) <= (layer5_outputs(3779)) and not (layer5_outputs(5123));
    layer6_outputs(1704) <= not((layer5_outputs(2849)) xor (layer5_outputs(1415)));
    layer6_outputs(1705) <= layer5_outputs(6140);
    layer6_outputs(1706) <= not(layer5_outputs(4498));
    layer6_outputs(1707) <= not(layer5_outputs(5632));
    layer6_outputs(1708) <= not(layer5_outputs(5951));
    layer6_outputs(1709) <= not(layer5_outputs(6503));
    layer6_outputs(1710) <= not(layer5_outputs(3245));
    layer6_outputs(1711) <= not(layer5_outputs(4197));
    layer6_outputs(1712) <= (layer5_outputs(1642)) xor (layer5_outputs(4479));
    layer6_outputs(1713) <= layer5_outputs(744);
    layer6_outputs(1714) <= (layer5_outputs(305)) or (layer5_outputs(894));
    layer6_outputs(1715) <= not(layer5_outputs(4813)) or (layer5_outputs(4730));
    layer6_outputs(1716) <= not(layer5_outputs(2980));
    layer6_outputs(1717) <= layer5_outputs(1887);
    layer6_outputs(1718) <= (layer5_outputs(4195)) xor (layer5_outputs(7488));
    layer6_outputs(1719) <= not((layer5_outputs(249)) and (layer5_outputs(3162)));
    layer6_outputs(1720) <= not(layer5_outputs(697));
    layer6_outputs(1721) <= (layer5_outputs(5859)) xor (layer5_outputs(4617));
    layer6_outputs(1722) <= (layer5_outputs(4370)) and (layer5_outputs(1337));
    layer6_outputs(1723) <= (layer5_outputs(4435)) and not (layer5_outputs(3613));
    layer6_outputs(1724) <= not(layer5_outputs(5468));
    layer6_outputs(1725) <= layer5_outputs(2730);
    layer6_outputs(1726) <= layer5_outputs(426);
    layer6_outputs(1727) <= not(layer5_outputs(6578));
    layer6_outputs(1728) <= layer5_outputs(1115);
    layer6_outputs(1729) <= not(layer5_outputs(1898));
    layer6_outputs(1730) <= not(layer5_outputs(4383)) or (layer5_outputs(5705));
    layer6_outputs(1731) <= not(layer5_outputs(1152));
    layer6_outputs(1732) <= not((layer5_outputs(4050)) xor (layer5_outputs(6674)));
    layer6_outputs(1733) <= not(layer5_outputs(3320));
    layer6_outputs(1734) <= not(layer5_outputs(5223));
    layer6_outputs(1735) <= not(layer5_outputs(1560)) or (layer5_outputs(3913));
    layer6_outputs(1736) <= layer5_outputs(3220);
    layer6_outputs(1737) <= not((layer5_outputs(447)) and (layer5_outputs(1121)));
    layer6_outputs(1738) <= layer5_outputs(4089);
    layer6_outputs(1739) <= not((layer5_outputs(7315)) and (layer5_outputs(2317)));
    layer6_outputs(1740) <= '1';
    layer6_outputs(1741) <= not(layer5_outputs(6919));
    layer6_outputs(1742) <= not(layer5_outputs(2482));
    layer6_outputs(1743) <= layer5_outputs(5985);
    layer6_outputs(1744) <= (layer5_outputs(7671)) and not (layer5_outputs(3553));
    layer6_outputs(1745) <= not((layer5_outputs(3647)) or (layer5_outputs(1933)));
    layer6_outputs(1746) <= layer5_outputs(5653);
    layer6_outputs(1747) <= (layer5_outputs(203)) xor (layer5_outputs(1082));
    layer6_outputs(1748) <= (layer5_outputs(6979)) and not (layer5_outputs(247));
    layer6_outputs(1749) <= (layer5_outputs(1089)) xor (layer5_outputs(2755));
    layer6_outputs(1750) <= not(layer5_outputs(5027));
    layer6_outputs(1751) <= not(layer5_outputs(3748)) or (layer5_outputs(4472));
    layer6_outputs(1752) <= (layer5_outputs(2189)) or (layer5_outputs(5342));
    layer6_outputs(1753) <= not(layer5_outputs(1339));
    layer6_outputs(1754) <= layer5_outputs(180);
    layer6_outputs(1755) <= not((layer5_outputs(5432)) xor (layer5_outputs(6451)));
    layer6_outputs(1756) <= not(layer5_outputs(3250)) or (layer5_outputs(26));
    layer6_outputs(1757) <= not((layer5_outputs(5325)) and (layer5_outputs(7626)));
    layer6_outputs(1758) <= (layer5_outputs(1216)) xor (layer5_outputs(3776));
    layer6_outputs(1759) <= layer5_outputs(3524);
    layer6_outputs(1760) <= not(layer5_outputs(4426)) or (layer5_outputs(6259));
    layer6_outputs(1761) <= (layer5_outputs(1103)) xor (layer5_outputs(1847));
    layer6_outputs(1762) <= layer5_outputs(7618);
    layer6_outputs(1763) <= layer5_outputs(7616);
    layer6_outputs(1764) <= (layer5_outputs(1588)) and (layer5_outputs(3188));
    layer6_outputs(1765) <= layer5_outputs(475);
    layer6_outputs(1766) <= (layer5_outputs(89)) and not (layer5_outputs(3336));
    layer6_outputs(1767) <= layer5_outputs(5138);
    layer6_outputs(1768) <= (layer5_outputs(5606)) and (layer5_outputs(1173));
    layer6_outputs(1769) <= layer5_outputs(1107);
    layer6_outputs(1770) <= not(layer5_outputs(3307));
    layer6_outputs(1771) <= not(layer5_outputs(5323));
    layer6_outputs(1772) <= not(layer5_outputs(4225));
    layer6_outputs(1773) <= (layer5_outputs(2913)) and not (layer5_outputs(2694));
    layer6_outputs(1774) <= not((layer5_outputs(5838)) xor (layer5_outputs(6306)));
    layer6_outputs(1775) <= (layer5_outputs(3301)) or (layer5_outputs(3157));
    layer6_outputs(1776) <= not(layer5_outputs(2791)) or (layer5_outputs(5101));
    layer6_outputs(1777) <= not(layer5_outputs(1129));
    layer6_outputs(1778) <= layer5_outputs(1787);
    layer6_outputs(1779) <= (layer5_outputs(5536)) xor (layer5_outputs(3324));
    layer6_outputs(1780) <= (layer5_outputs(5390)) and not (layer5_outputs(3459));
    layer6_outputs(1781) <= not(layer5_outputs(3729)) or (layer5_outputs(3762));
    layer6_outputs(1782) <= not(layer5_outputs(5070)) or (layer5_outputs(1876));
    layer6_outputs(1783) <= not(layer5_outputs(2177));
    layer6_outputs(1784) <= (layer5_outputs(5247)) xor (layer5_outputs(1885));
    layer6_outputs(1785) <= layer5_outputs(5907);
    layer6_outputs(1786) <= not((layer5_outputs(4193)) xor (layer5_outputs(2563)));
    layer6_outputs(1787) <= not(layer5_outputs(1113));
    layer6_outputs(1788) <= not(layer5_outputs(4786));
    layer6_outputs(1789) <= (layer5_outputs(4641)) or (layer5_outputs(3455));
    layer6_outputs(1790) <= layer5_outputs(5590);
    layer6_outputs(1791) <= layer5_outputs(1798);
    layer6_outputs(1792) <= layer5_outputs(4380);
    layer6_outputs(1793) <= not(layer5_outputs(1583));
    layer6_outputs(1794) <= not((layer5_outputs(2220)) or (layer5_outputs(1837)));
    layer6_outputs(1795) <= not((layer5_outputs(1098)) or (layer5_outputs(6315)));
    layer6_outputs(1796) <= (layer5_outputs(1715)) xor (layer5_outputs(2634));
    layer6_outputs(1797) <= not(layer5_outputs(618)) or (layer5_outputs(5619));
    layer6_outputs(1798) <= not(layer5_outputs(5360)) or (layer5_outputs(4015));
    layer6_outputs(1799) <= layer5_outputs(459);
    layer6_outputs(1800) <= (layer5_outputs(1634)) xor (layer5_outputs(5923));
    layer6_outputs(1801) <= layer5_outputs(2536);
    layer6_outputs(1802) <= not(layer5_outputs(5595));
    layer6_outputs(1803) <= (layer5_outputs(3392)) and not (layer5_outputs(5175));
    layer6_outputs(1804) <= layer5_outputs(3351);
    layer6_outputs(1805) <= layer5_outputs(705);
    layer6_outputs(1806) <= (layer5_outputs(3202)) and (layer5_outputs(1190));
    layer6_outputs(1807) <= not(layer5_outputs(954)) or (layer5_outputs(2460));
    layer6_outputs(1808) <= not((layer5_outputs(4839)) and (layer5_outputs(5327)));
    layer6_outputs(1809) <= (layer5_outputs(3641)) or (layer5_outputs(2211));
    layer6_outputs(1810) <= (layer5_outputs(5119)) and not (layer5_outputs(7031));
    layer6_outputs(1811) <= layer5_outputs(199);
    layer6_outputs(1812) <= (layer5_outputs(7109)) and not (layer5_outputs(81));
    layer6_outputs(1813) <= not(layer5_outputs(2159));
    layer6_outputs(1814) <= layer5_outputs(5477);
    layer6_outputs(1815) <= not((layer5_outputs(2674)) and (layer5_outputs(3826)));
    layer6_outputs(1816) <= layer5_outputs(4236);
    layer6_outputs(1817) <= layer5_outputs(2275);
    layer6_outputs(1818) <= (layer5_outputs(3391)) and not (layer5_outputs(6190));
    layer6_outputs(1819) <= not(layer5_outputs(3337));
    layer6_outputs(1820) <= (layer5_outputs(1784)) and not (layer5_outputs(5825));
    layer6_outputs(1821) <= not((layer5_outputs(4590)) xor (layer5_outputs(3721)));
    layer6_outputs(1822) <= not(layer5_outputs(7446));
    layer6_outputs(1823) <= not(layer5_outputs(7017));
    layer6_outputs(1824) <= '1';
    layer6_outputs(1825) <= layer5_outputs(4412);
    layer6_outputs(1826) <= layer5_outputs(2890);
    layer6_outputs(1827) <= (layer5_outputs(6457)) and not (layer5_outputs(6201));
    layer6_outputs(1828) <= not(layer5_outputs(963)) or (layer5_outputs(1506));
    layer6_outputs(1829) <= not(layer5_outputs(7053));
    layer6_outputs(1830) <= not(layer5_outputs(3372));
    layer6_outputs(1831) <= not(layer5_outputs(6851));
    layer6_outputs(1832) <= layer5_outputs(7047);
    layer6_outputs(1833) <= layer5_outputs(2462);
    layer6_outputs(1834) <= layer5_outputs(4012);
    layer6_outputs(1835) <= not(layer5_outputs(1376));
    layer6_outputs(1836) <= '1';
    layer6_outputs(1837) <= not(layer5_outputs(5380)) or (layer5_outputs(1848));
    layer6_outputs(1838) <= not((layer5_outputs(2090)) xor (layer5_outputs(4378)));
    layer6_outputs(1839) <= layer5_outputs(7193);
    layer6_outputs(1840) <= layer5_outputs(1745);
    layer6_outputs(1841) <= not(layer5_outputs(5095)) or (layer5_outputs(3856));
    layer6_outputs(1842) <= layer5_outputs(2535);
    layer6_outputs(1843) <= (layer5_outputs(2772)) and not (layer5_outputs(6400));
    layer6_outputs(1844) <= not(layer5_outputs(4356)) or (layer5_outputs(957));
    layer6_outputs(1845) <= not(layer5_outputs(4833));
    layer6_outputs(1846) <= layer5_outputs(4226);
    layer6_outputs(1847) <= (layer5_outputs(7322)) and (layer5_outputs(635));
    layer6_outputs(1848) <= not(layer5_outputs(7143)) or (layer5_outputs(4258));
    layer6_outputs(1849) <= layer5_outputs(3974);
    layer6_outputs(1850) <= layer5_outputs(1480);
    layer6_outputs(1851) <= not(layer5_outputs(5921));
    layer6_outputs(1852) <= not((layer5_outputs(7577)) or (layer5_outputs(5567)));
    layer6_outputs(1853) <= not(layer5_outputs(6435)) or (layer5_outputs(294));
    layer6_outputs(1854) <= not((layer5_outputs(5582)) xor (layer5_outputs(4749)));
    layer6_outputs(1855) <= not((layer5_outputs(7173)) xor (layer5_outputs(6065)));
    layer6_outputs(1856) <= (layer5_outputs(2443)) xor (layer5_outputs(1776));
    layer6_outputs(1857) <= not((layer5_outputs(5656)) and (layer5_outputs(421)));
    layer6_outputs(1858) <= not((layer5_outputs(467)) or (layer5_outputs(3921)));
    layer6_outputs(1859) <= (layer5_outputs(6817)) or (layer5_outputs(2783));
    layer6_outputs(1860) <= not(layer5_outputs(3462));
    layer6_outputs(1861) <= not((layer5_outputs(505)) or (layer5_outputs(4754)));
    layer6_outputs(1862) <= not(layer5_outputs(1829));
    layer6_outputs(1863) <= layer5_outputs(7603);
    layer6_outputs(1864) <= (layer5_outputs(4813)) and not (layer5_outputs(2353));
    layer6_outputs(1865) <= not(layer5_outputs(7672));
    layer6_outputs(1866) <= not(layer5_outputs(6654));
    layer6_outputs(1867) <= not((layer5_outputs(921)) and (layer5_outputs(3679)));
    layer6_outputs(1868) <= layer5_outputs(3052);
    layer6_outputs(1869) <= not(layer5_outputs(3352)) or (layer5_outputs(4081));
    layer6_outputs(1870) <= layer5_outputs(7437);
    layer6_outputs(1871) <= (layer5_outputs(6213)) and not (layer5_outputs(7273));
    layer6_outputs(1872) <= (layer5_outputs(5554)) and (layer5_outputs(2580));
    layer6_outputs(1873) <= not((layer5_outputs(4286)) or (layer5_outputs(6295)));
    layer6_outputs(1874) <= layer5_outputs(2577);
    layer6_outputs(1875) <= (layer5_outputs(5041)) xor (layer5_outputs(3816));
    layer6_outputs(1876) <= layer5_outputs(6811);
    layer6_outputs(1877) <= (layer5_outputs(2699)) and not (layer5_outputs(6755));
    layer6_outputs(1878) <= (layer5_outputs(6532)) and not (layer5_outputs(4171));
    layer6_outputs(1879) <= not(layer5_outputs(1456)) or (layer5_outputs(4455));
    layer6_outputs(1880) <= (layer5_outputs(1019)) and (layer5_outputs(3099));
    layer6_outputs(1881) <= (layer5_outputs(2016)) and not (layer5_outputs(7369));
    layer6_outputs(1882) <= not((layer5_outputs(5953)) or (layer5_outputs(3911)));
    layer6_outputs(1883) <= (layer5_outputs(6398)) and not (layer5_outputs(3521));
    layer6_outputs(1884) <= (layer5_outputs(802)) xor (layer5_outputs(503));
    layer6_outputs(1885) <= not(layer5_outputs(4250));
    layer6_outputs(1886) <= layer5_outputs(483);
    layer6_outputs(1887) <= not(layer5_outputs(5664));
    layer6_outputs(1888) <= layer5_outputs(7196);
    layer6_outputs(1889) <= not((layer5_outputs(4801)) and (layer5_outputs(6589)));
    layer6_outputs(1890) <= not((layer5_outputs(1235)) or (layer5_outputs(7177)));
    layer6_outputs(1891) <= not(layer5_outputs(6068));
    layer6_outputs(1892) <= layer5_outputs(1444);
    layer6_outputs(1893) <= not(layer5_outputs(1759));
    layer6_outputs(1894) <= layer5_outputs(5080);
    layer6_outputs(1895) <= (layer5_outputs(1716)) and (layer5_outputs(1103));
    layer6_outputs(1896) <= not(layer5_outputs(197)) or (layer5_outputs(6747));
    layer6_outputs(1897) <= layer5_outputs(2962);
    layer6_outputs(1898) <= not(layer5_outputs(3757)) or (layer5_outputs(7334));
    layer6_outputs(1899) <= not(layer5_outputs(4824));
    layer6_outputs(1900) <= not(layer5_outputs(5109)) or (layer5_outputs(5409));
    layer6_outputs(1901) <= not((layer5_outputs(2704)) or (layer5_outputs(1700)));
    layer6_outputs(1902) <= layer5_outputs(3993);
    layer6_outputs(1903) <= not((layer5_outputs(4592)) xor (layer5_outputs(5616)));
    layer6_outputs(1904) <= layer5_outputs(2265);
    layer6_outputs(1905) <= layer5_outputs(7407);
    layer6_outputs(1906) <= not(layer5_outputs(4111));
    layer6_outputs(1907) <= layer5_outputs(5700);
    layer6_outputs(1908) <= (layer5_outputs(1465)) and not (layer5_outputs(7526));
    layer6_outputs(1909) <= layer5_outputs(5062);
    layer6_outputs(1910) <= (layer5_outputs(4733)) xor (layer5_outputs(678));
    layer6_outputs(1911) <= not((layer5_outputs(4628)) xor (layer5_outputs(3373)));
    layer6_outputs(1912) <= not(layer5_outputs(4364));
    layer6_outputs(1913) <= not(layer5_outputs(7066));
    layer6_outputs(1914) <= not(layer5_outputs(7602));
    layer6_outputs(1915) <= not(layer5_outputs(3121));
    layer6_outputs(1916) <= not(layer5_outputs(6122)) or (layer5_outputs(563));
    layer6_outputs(1917) <= not((layer5_outputs(6273)) or (layer5_outputs(1554)));
    layer6_outputs(1918) <= layer5_outputs(2447);
    layer6_outputs(1919) <= layer5_outputs(7482);
    layer6_outputs(1920) <= (layer5_outputs(486)) xor (layer5_outputs(5520));
    layer6_outputs(1921) <= not((layer5_outputs(6815)) xor (layer5_outputs(1288)));
    layer6_outputs(1922) <= (layer5_outputs(7402)) xor (layer5_outputs(4702));
    layer6_outputs(1923) <= layer5_outputs(5028);
    layer6_outputs(1924) <= layer5_outputs(311);
    layer6_outputs(1925) <= layer5_outputs(7413);
    layer6_outputs(1926) <= not(layer5_outputs(6018));
    layer6_outputs(1927) <= layer5_outputs(3424);
    layer6_outputs(1928) <= layer5_outputs(1173);
    layer6_outputs(1929) <= not((layer5_outputs(6128)) or (layer5_outputs(5258)));
    layer6_outputs(1930) <= not(layer5_outputs(5244));
    layer6_outputs(1931) <= not((layer5_outputs(1643)) or (layer5_outputs(7235)));
    layer6_outputs(1932) <= layer5_outputs(7202);
    layer6_outputs(1933) <= layer5_outputs(4930);
    layer6_outputs(1934) <= not((layer5_outputs(4156)) and (layer5_outputs(1497)));
    layer6_outputs(1935) <= (layer5_outputs(5426)) xor (layer5_outputs(5386));
    layer6_outputs(1936) <= not((layer5_outputs(6828)) xor (layer5_outputs(7570)));
    layer6_outputs(1937) <= layer5_outputs(3678);
    layer6_outputs(1938) <= not((layer5_outputs(1701)) xor (layer5_outputs(3691)));
    layer6_outputs(1939) <= layer5_outputs(2511);
    layer6_outputs(1940) <= not((layer5_outputs(2510)) and (layer5_outputs(5309)));
    layer6_outputs(1941) <= not(layer5_outputs(1768)) or (layer5_outputs(1129));
    layer6_outputs(1942) <= not((layer5_outputs(7060)) xor (layer5_outputs(2919)));
    layer6_outputs(1943) <= not(layer5_outputs(6821));
    layer6_outputs(1944) <= not(layer5_outputs(709));
    layer6_outputs(1945) <= (layer5_outputs(1804)) and (layer5_outputs(1990));
    layer6_outputs(1946) <= layer5_outputs(6869);
    layer6_outputs(1947) <= not(layer5_outputs(466));
    layer6_outputs(1948) <= not(layer5_outputs(4847));
    layer6_outputs(1949) <= layer5_outputs(1679);
    layer6_outputs(1950) <= (layer5_outputs(1636)) xor (layer5_outputs(3521));
    layer6_outputs(1951) <= not((layer5_outputs(4262)) xor (layer5_outputs(1296)));
    layer6_outputs(1952) <= (layer5_outputs(4476)) and not (layer5_outputs(7317));
    layer6_outputs(1953) <= (layer5_outputs(7393)) and (layer5_outputs(4351));
    layer6_outputs(1954) <= (layer5_outputs(1282)) or (layer5_outputs(2292));
    layer6_outputs(1955) <= layer5_outputs(532);
    layer6_outputs(1956) <= not((layer5_outputs(5852)) or (layer5_outputs(1811)));
    layer6_outputs(1957) <= (layer5_outputs(29)) and (layer5_outputs(7395));
    layer6_outputs(1958) <= (layer5_outputs(3933)) and not (layer5_outputs(1846));
    layer6_outputs(1959) <= not((layer5_outputs(6461)) xor (layer5_outputs(6576)));
    layer6_outputs(1960) <= layer5_outputs(524);
    layer6_outputs(1961) <= not(layer5_outputs(2744));
    layer6_outputs(1962) <= layer5_outputs(615);
    layer6_outputs(1963) <= not(layer5_outputs(984));
    layer6_outputs(1964) <= layer5_outputs(6841);
    layer6_outputs(1965) <= not((layer5_outputs(3073)) and (layer5_outputs(3859)));
    layer6_outputs(1966) <= (layer5_outputs(4783)) xor (layer5_outputs(2977));
    layer6_outputs(1967) <= not(layer5_outputs(4818));
    layer6_outputs(1968) <= layer5_outputs(6611);
    layer6_outputs(1969) <= layer5_outputs(5917);
    layer6_outputs(1970) <= not((layer5_outputs(703)) and (layer5_outputs(2097)));
    layer6_outputs(1971) <= layer5_outputs(10);
    layer6_outputs(1972) <= not(layer5_outputs(66));
    layer6_outputs(1973) <= not(layer5_outputs(5590));
    layer6_outputs(1974) <= layer5_outputs(507);
    layer6_outputs(1975) <= (layer5_outputs(4598)) and not (layer5_outputs(5396));
    layer6_outputs(1976) <= (layer5_outputs(4259)) and (layer5_outputs(3643));
    layer6_outputs(1977) <= not(layer5_outputs(3880));
    layer6_outputs(1978) <= not((layer5_outputs(7097)) and (layer5_outputs(4963)));
    layer6_outputs(1979) <= (layer5_outputs(4237)) or (layer5_outputs(514));
    layer6_outputs(1980) <= layer5_outputs(2741);
    layer6_outputs(1981) <= not((layer5_outputs(864)) xor (layer5_outputs(5496)));
    layer6_outputs(1982) <= (layer5_outputs(5186)) xor (layer5_outputs(3639));
    layer6_outputs(1983) <= layer5_outputs(7597);
    layer6_outputs(1984) <= not((layer5_outputs(3375)) and (layer5_outputs(4134)));
    layer6_outputs(1985) <= layer5_outputs(5204);
    layer6_outputs(1986) <= layer5_outputs(1624);
    layer6_outputs(1987) <= not(layer5_outputs(3466)) or (layer5_outputs(5271));
    layer6_outputs(1988) <= not((layer5_outputs(5198)) xor (layer5_outputs(4651)));
    layer6_outputs(1989) <= (layer5_outputs(4268)) xor (layer5_outputs(706));
    layer6_outputs(1990) <= not(layer5_outputs(514));
    layer6_outputs(1991) <= not(layer5_outputs(5250)) or (layer5_outputs(2167));
    layer6_outputs(1992) <= (layer5_outputs(4321)) or (layer5_outputs(4607));
    layer6_outputs(1993) <= layer5_outputs(521);
    layer6_outputs(1994) <= (layer5_outputs(5073)) xor (layer5_outputs(4444));
    layer6_outputs(1995) <= not(layer5_outputs(3931));
    layer6_outputs(1996) <= (layer5_outputs(4530)) or (layer5_outputs(3224));
    layer6_outputs(1997) <= (layer5_outputs(1252)) and not (layer5_outputs(7135));
    layer6_outputs(1998) <= not(layer5_outputs(657));
    layer6_outputs(1999) <= not(layer5_outputs(2085)) or (layer5_outputs(5264));
    layer6_outputs(2000) <= layer5_outputs(1568);
    layer6_outputs(2001) <= (layer5_outputs(6738)) xor (layer5_outputs(2328));
    layer6_outputs(2002) <= not((layer5_outputs(6996)) or (layer5_outputs(3317)));
    layer6_outputs(2003) <= not((layer5_outputs(6422)) or (layer5_outputs(105)));
    layer6_outputs(2004) <= layer5_outputs(6929);
    layer6_outputs(2005) <= (layer5_outputs(1966)) and (layer5_outputs(5811));
    layer6_outputs(2006) <= layer5_outputs(1025);
    layer6_outputs(2007) <= not(layer5_outputs(4374));
    layer6_outputs(2008) <= (layer5_outputs(6440)) and not (layer5_outputs(3922));
    layer6_outputs(2009) <= not(layer5_outputs(1703));
    layer6_outputs(2010) <= not(layer5_outputs(3497));
    layer6_outputs(2011) <= layer5_outputs(1832);
    layer6_outputs(2012) <= (layer5_outputs(7121)) or (layer5_outputs(4004));
    layer6_outputs(2013) <= not(layer5_outputs(7578));
    layer6_outputs(2014) <= not(layer5_outputs(6860));
    layer6_outputs(2015) <= not(layer5_outputs(2141));
    layer6_outputs(2016) <= (layer5_outputs(2226)) or (layer5_outputs(5847));
    layer6_outputs(2017) <= not(layer5_outputs(1686));
    layer6_outputs(2018) <= not(layer5_outputs(4671));
    layer6_outputs(2019) <= not(layer5_outputs(6748));
    layer6_outputs(2020) <= layer5_outputs(1600);
    layer6_outputs(2021) <= not((layer5_outputs(7659)) and (layer5_outputs(3499)));
    layer6_outputs(2022) <= not(layer5_outputs(1308));
    layer6_outputs(2023) <= not(layer5_outputs(4689));
    layer6_outputs(2024) <= not(layer5_outputs(3690));
    layer6_outputs(2025) <= (layer5_outputs(5197)) and (layer5_outputs(116));
    layer6_outputs(2026) <= not(layer5_outputs(5327));
    layer6_outputs(2027) <= not(layer5_outputs(2906));
    layer6_outputs(2028) <= layer5_outputs(162);
    layer6_outputs(2029) <= layer5_outputs(3445);
    layer6_outputs(2030) <= not((layer5_outputs(6446)) xor (layer5_outputs(3846)));
    layer6_outputs(2031) <= not((layer5_outputs(6167)) or (layer5_outputs(5787)));
    layer6_outputs(2032) <= not(layer5_outputs(5007));
    layer6_outputs(2033) <= not(layer5_outputs(3215));
    layer6_outputs(2034) <= not(layer5_outputs(4987));
    layer6_outputs(2035) <= not(layer5_outputs(5583));
    layer6_outputs(2036) <= not(layer5_outputs(5894));
    layer6_outputs(2037) <= (layer5_outputs(6263)) and not (layer5_outputs(1466));
    layer6_outputs(2038) <= not(layer5_outputs(711));
    layer6_outputs(2039) <= (layer5_outputs(4595)) and not (layer5_outputs(7479));
    layer6_outputs(2040) <= not((layer5_outputs(4834)) and (layer5_outputs(3143)));
    layer6_outputs(2041) <= not(layer5_outputs(4626));
    layer6_outputs(2042) <= layer5_outputs(4839);
    layer6_outputs(2043) <= not(layer5_outputs(3181)) or (layer5_outputs(7254));
    layer6_outputs(2044) <= layer5_outputs(901);
    layer6_outputs(2045) <= not((layer5_outputs(835)) xor (layer5_outputs(4805)));
    layer6_outputs(2046) <= layer5_outputs(3458);
    layer6_outputs(2047) <= not(layer5_outputs(6638));
    layer6_outputs(2048) <= not(layer5_outputs(5415));
    layer6_outputs(2049) <= (layer5_outputs(4577)) and not (layer5_outputs(3082));
    layer6_outputs(2050) <= not(layer5_outputs(833));
    layer6_outputs(2051) <= (layer5_outputs(4001)) and not (layer5_outputs(2043));
    layer6_outputs(2052) <= not(layer5_outputs(6312));
    layer6_outputs(2053) <= not(layer5_outputs(7367));
    layer6_outputs(2054) <= not(layer5_outputs(2562));
    layer6_outputs(2055) <= not(layer5_outputs(6617));
    layer6_outputs(2056) <= not((layer5_outputs(6153)) or (layer5_outputs(3032)));
    layer6_outputs(2057) <= not(layer5_outputs(3689));
    layer6_outputs(2058) <= not(layer5_outputs(4561)) or (layer5_outputs(1335));
    layer6_outputs(2059) <= not(layer5_outputs(4419)) or (layer5_outputs(7132));
    layer6_outputs(2060) <= layer5_outputs(1504);
    layer6_outputs(2061) <= (layer5_outputs(2295)) and not (layer5_outputs(5521));
    layer6_outputs(2062) <= layer5_outputs(3780);
    layer6_outputs(2063) <= not(layer5_outputs(5160)) or (layer5_outputs(3573));
    layer6_outputs(2064) <= (layer5_outputs(4408)) xor (layer5_outputs(6384));
    layer6_outputs(2065) <= (layer5_outputs(5300)) and not (layer5_outputs(3911));
    layer6_outputs(2066) <= not(layer5_outputs(226)) or (layer5_outputs(5944));
    layer6_outputs(2067) <= not(layer5_outputs(5877));
    layer6_outputs(2068) <= not((layer5_outputs(4580)) or (layer5_outputs(174)));
    layer6_outputs(2069) <= layer5_outputs(1150);
    layer6_outputs(2070) <= not((layer5_outputs(239)) xor (layer5_outputs(1459)));
    layer6_outputs(2071) <= layer5_outputs(4750);
    layer6_outputs(2072) <= not((layer5_outputs(7262)) and (layer5_outputs(7022)));
    layer6_outputs(2073) <= not((layer5_outputs(5030)) xor (layer5_outputs(6763)));
    layer6_outputs(2074) <= layer5_outputs(470);
    layer6_outputs(2075) <= not((layer5_outputs(325)) and (layer5_outputs(4826)));
    layer6_outputs(2076) <= (layer5_outputs(6637)) and not (layer5_outputs(4128));
    layer6_outputs(2077) <= not(layer5_outputs(1016));
    layer6_outputs(2078) <= (layer5_outputs(1897)) xor (layer5_outputs(7550));
    layer6_outputs(2079) <= (layer5_outputs(713)) and (layer5_outputs(2303));
    layer6_outputs(2080) <= layer5_outputs(275);
    layer6_outputs(2081) <= not((layer5_outputs(2867)) and (layer5_outputs(4658)));
    layer6_outputs(2082) <= not(layer5_outputs(3382));
    layer6_outputs(2083) <= not(layer5_outputs(906));
    layer6_outputs(2084) <= layer5_outputs(5524);
    layer6_outputs(2085) <= layer5_outputs(6741);
    layer6_outputs(2086) <= layer5_outputs(5472);
    layer6_outputs(2087) <= layer5_outputs(7288);
    layer6_outputs(2088) <= layer5_outputs(5406);
    layer6_outputs(2089) <= layer5_outputs(1046);
    layer6_outputs(2090) <= not(layer5_outputs(3502));
    layer6_outputs(2091) <= layer5_outputs(2541);
    layer6_outputs(2092) <= not((layer5_outputs(1094)) and (layer5_outputs(5770)));
    layer6_outputs(2093) <= (layer5_outputs(944)) xor (layer5_outputs(329));
    layer6_outputs(2094) <= layer5_outputs(4417);
    layer6_outputs(2095) <= not((layer5_outputs(7402)) xor (layer5_outputs(4360)));
    layer6_outputs(2096) <= layer5_outputs(5116);
    layer6_outputs(2097) <= (layer5_outputs(118)) or (layer5_outputs(4353));
    layer6_outputs(2098) <= layer5_outputs(4156);
    layer6_outputs(2099) <= not((layer5_outputs(3018)) or (layer5_outputs(2752)));
    layer6_outputs(2100) <= layer5_outputs(817);
    layer6_outputs(2101) <= not(layer5_outputs(2782));
    layer6_outputs(2102) <= (layer5_outputs(1114)) xor (layer5_outputs(4527));
    layer6_outputs(2103) <= (layer5_outputs(143)) xor (layer5_outputs(4028));
    layer6_outputs(2104) <= layer5_outputs(2487);
    layer6_outputs(2105) <= (layer5_outputs(2357)) and not (layer5_outputs(2165));
    layer6_outputs(2106) <= not(layer5_outputs(3012));
    layer6_outputs(2107) <= (layer5_outputs(2933)) and not (layer5_outputs(4167));
    layer6_outputs(2108) <= layer5_outputs(3561);
    layer6_outputs(2109) <= layer5_outputs(4830);
    layer6_outputs(2110) <= layer5_outputs(2392);
    layer6_outputs(2111) <= not(layer5_outputs(4430)) or (layer5_outputs(358));
    layer6_outputs(2112) <= not(layer5_outputs(3720));
    layer6_outputs(2113) <= not((layer5_outputs(7660)) xor (layer5_outputs(5688)));
    layer6_outputs(2114) <= layer5_outputs(5870);
    layer6_outputs(2115) <= not(layer5_outputs(4043));
    layer6_outputs(2116) <= (layer5_outputs(3048)) and not (layer5_outputs(2391));
    layer6_outputs(2117) <= layer5_outputs(3437);
    layer6_outputs(2118) <= (layer5_outputs(697)) xor (layer5_outputs(6533));
    layer6_outputs(2119) <= (layer5_outputs(7427)) and (layer5_outputs(1584));
    layer6_outputs(2120) <= (layer5_outputs(6804)) xor (layer5_outputs(1535));
    layer6_outputs(2121) <= layer5_outputs(1286);
    layer6_outputs(2122) <= layer5_outputs(5095);
    layer6_outputs(2123) <= not(layer5_outputs(1621));
    layer6_outputs(2124) <= not(layer5_outputs(4323));
    layer6_outputs(2125) <= not(layer5_outputs(4995));
    layer6_outputs(2126) <= layer5_outputs(7269);
    layer6_outputs(2127) <= (layer5_outputs(1061)) xor (layer5_outputs(3089));
    layer6_outputs(2128) <= layer5_outputs(7168);
    layer6_outputs(2129) <= (layer5_outputs(4124)) and not (layer5_outputs(4811));
    layer6_outputs(2130) <= not(layer5_outputs(5201));
    layer6_outputs(2131) <= not(layer5_outputs(2758));
    layer6_outputs(2132) <= not((layer5_outputs(849)) or (layer5_outputs(3529)));
    layer6_outputs(2133) <= not(layer5_outputs(1334)) or (layer5_outputs(2735));
    layer6_outputs(2134) <= not(layer5_outputs(5035));
    layer6_outputs(2135) <= not(layer5_outputs(6452));
    layer6_outputs(2136) <= not((layer5_outputs(3359)) xor (layer5_outputs(2224)));
    layer6_outputs(2137) <= not(layer5_outputs(5269));
    layer6_outputs(2138) <= not((layer5_outputs(738)) xor (layer5_outputs(2958)));
    layer6_outputs(2139) <= not(layer5_outputs(6456));
    layer6_outputs(2140) <= layer5_outputs(609);
    layer6_outputs(2141) <= (layer5_outputs(5260)) xor (layer5_outputs(473));
    layer6_outputs(2142) <= layer5_outputs(2458);
    layer6_outputs(2143) <= '0';
    layer6_outputs(2144) <= (layer5_outputs(4403)) and (layer5_outputs(3122));
    layer6_outputs(2145) <= not((layer5_outputs(6836)) xor (layer5_outputs(5689)));
    layer6_outputs(2146) <= (layer5_outputs(1725)) and not (layer5_outputs(6166));
    layer6_outputs(2147) <= not(layer5_outputs(265)) or (layer5_outputs(866));
    layer6_outputs(2148) <= (layer5_outputs(6026)) xor (layer5_outputs(5965));
    layer6_outputs(2149) <= not(layer5_outputs(2418));
    layer6_outputs(2150) <= not(layer5_outputs(2237));
    layer6_outputs(2151) <= layer5_outputs(5192);
    layer6_outputs(2152) <= layer5_outputs(1027);
    layer6_outputs(2153) <= not(layer5_outputs(4980));
    layer6_outputs(2154) <= not(layer5_outputs(6307));
    layer6_outputs(2155) <= not(layer5_outputs(4202));
    layer6_outputs(2156) <= not((layer5_outputs(1437)) or (layer5_outputs(3749)));
    layer6_outputs(2157) <= not(layer5_outputs(6854));
    layer6_outputs(2158) <= not(layer5_outputs(3624));
    layer6_outputs(2159) <= (layer5_outputs(3196)) and not (layer5_outputs(2131));
    layer6_outputs(2160) <= (layer5_outputs(3310)) xor (layer5_outputs(2125));
    layer6_outputs(2161) <= not((layer5_outputs(5718)) xor (layer5_outputs(1781)));
    layer6_outputs(2162) <= layer5_outputs(1157);
    layer6_outputs(2163) <= (layer5_outputs(4009)) and not (layer5_outputs(3445));
    layer6_outputs(2164) <= (layer5_outputs(1657)) and not (layer5_outputs(4507));
    layer6_outputs(2165) <= not(layer5_outputs(2120));
    layer6_outputs(2166) <= not(layer5_outputs(3814));
    layer6_outputs(2167) <= (layer5_outputs(7266)) xor (layer5_outputs(6629));
    layer6_outputs(2168) <= layer5_outputs(436);
    layer6_outputs(2169) <= layer5_outputs(5643);
    layer6_outputs(2170) <= not((layer5_outputs(5660)) xor (layer5_outputs(7251)));
    layer6_outputs(2171) <= not(layer5_outputs(6823));
    layer6_outputs(2172) <= not((layer5_outputs(5106)) xor (layer5_outputs(6560)));
    layer6_outputs(2173) <= not(layer5_outputs(6677)) or (layer5_outputs(4809));
    layer6_outputs(2174) <= layer5_outputs(685);
    layer6_outputs(2175) <= layer5_outputs(7414);
    layer6_outputs(2176) <= not(layer5_outputs(1665));
    layer6_outputs(2177) <= not(layer5_outputs(820));
    layer6_outputs(2178) <= (layer5_outputs(7593)) and not (layer5_outputs(1381));
    layer6_outputs(2179) <= not(layer5_outputs(7018));
    layer6_outputs(2180) <= (layer5_outputs(4204)) xor (layer5_outputs(5174));
    layer6_outputs(2181) <= not(layer5_outputs(2109));
    layer6_outputs(2182) <= not(layer5_outputs(1264));
    layer6_outputs(2183) <= not(layer5_outputs(909)) or (layer5_outputs(3028));
    layer6_outputs(2184) <= not(layer5_outputs(1336));
    layer6_outputs(2185) <= layer5_outputs(6285);
    layer6_outputs(2186) <= layer5_outputs(6369);
    layer6_outputs(2187) <= (layer5_outputs(1270)) and (layer5_outputs(2376));
    layer6_outputs(2188) <= layer5_outputs(3368);
    layer6_outputs(2189) <= not(layer5_outputs(1641));
    layer6_outputs(2190) <= not(layer5_outputs(6855));
    layer6_outputs(2191) <= (layer5_outputs(5353)) and (layer5_outputs(2666));
    layer6_outputs(2192) <= layer5_outputs(6110);
    layer6_outputs(2193) <= not(layer5_outputs(5281));
    layer6_outputs(2194) <= (layer5_outputs(5369)) and not (layer5_outputs(6691));
    layer6_outputs(2195) <= layer5_outputs(7347);
    layer6_outputs(2196) <= not(layer5_outputs(4033)) or (layer5_outputs(2471));
    layer6_outputs(2197) <= not(layer5_outputs(7229));
    layer6_outputs(2198) <= not((layer5_outputs(3456)) xor (layer5_outputs(1836)));
    layer6_outputs(2199) <= not(layer5_outputs(3174));
    layer6_outputs(2200) <= not((layer5_outputs(7071)) and (layer5_outputs(7509)));
    layer6_outputs(2201) <= not((layer5_outputs(7452)) or (layer5_outputs(7538)));
    layer6_outputs(2202) <= layer5_outputs(6539);
    layer6_outputs(2203) <= layer5_outputs(1052);
    layer6_outputs(2204) <= not((layer5_outputs(5557)) xor (layer5_outputs(6307)));
    layer6_outputs(2205) <= not(layer5_outputs(3407));
    layer6_outputs(2206) <= (layer5_outputs(6210)) and (layer5_outputs(2533));
    layer6_outputs(2207) <= layer5_outputs(1528);
    layer6_outputs(2208) <= not(layer5_outputs(4602)) or (layer5_outputs(3544));
    layer6_outputs(2209) <= layer5_outputs(1984);
    layer6_outputs(2210) <= not(layer5_outputs(2294));
    layer6_outputs(2211) <= not(layer5_outputs(727));
    layer6_outputs(2212) <= not(layer5_outputs(5498)) or (layer5_outputs(4895));
    layer6_outputs(2213) <= layer5_outputs(6237);
    layer6_outputs(2214) <= layer5_outputs(5308);
    layer6_outputs(2215) <= not(layer5_outputs(7045)) or (layer5_outputs(6496));
    layer6_outputs(2216) <= not(layer5_outputs(1365));
    layer6_outputs(2217) <= not(layer5_outputs(961)) or (layer5_outputs(2619));
    layer6_outputs(2218) <= '1';
    layer6_outputs(2219) <= not(layer5_outputs(2259));
    layer6_outputs(2220) <= (layer5_outputs(6922)) xor (layer5_outputs(600));
    layer6_outputs(2221) <= not(layer5_outputs(1959)) or (layer5_outputs(3371));
    layer6_outputs(2222) <= layer5_outputs(5255);
    layer6_outputs(2223) <= (layer5_outputs(313)) and not (layer5_outputs(4624));
    layer6_outputs(2224) <= not(layer5_outputs(2612));
    layer6_outputs(2225) <= not(layer5_outputs(7019));
    layer6_outputs(2226) <= not(layer5_outputs(4767));
    layer6_outputs(2227) <= not(layer5_outputs(1503)) or (layer5_outputs(2597));
    layer6_outputs(2228) <= layer5_outputs(7115);
    layer6_outputs(2229) <= layer5_outputs(779);
    layer6_outputs(2230) <= layer5_outputs(621);
    layer6_outputs(2231) <= (layer5_outputs(7514)) xor (layer5_outputs(285));
    layer6_outputs(2232) <= not((layer5_outputs(4666)) or (layer5_outputs(612)));
    layer6_outputs(2233) <= not(layer5_outputs(1904));
    layer6_outputs(2234) <= layer5_outputs(3160);
    layer6_outputs(2235) <= not(layer5_outputs(6339));
    layer6_outputs(2236) <= not((layer5_outputs(4653)) xor (layer5_outputs(3695)));
    layer6_outputs(2237) <= layer5_outputs(5317);
    layer6_outputs(2238) <= not(layer5_outputs(2431));
    layer6_outputs(2239) <= (layer5_outputs(332)) and not (layer5_outputs(5883));
    layer6_outputs(2240) <= not(layer5_outputs(3118)) or (layer5_outputs(7352));
    layer6_outputs(2241) <= layer5_outputs(973);
    layer6_outputs(2242) <= (layer5_outputs(492)) and not (layer5_outputs(4980));
    layer6_outputs(2243) <= layer5_outputs(2049);
    layer6_outputs(2244) <= not((layer5_outputs(2916)) xor (layer5_outputs(1075)));
    layer6_outputs(2245) <= not((layer5_outputs(3272)) xor (layer5_outputs(6243)));
    layer6_outputs(2246) <= (layer5_outputs(1877)) and not (layer5_outputs(5870));
    layer6_outputs(2247) <= not(layer5_outputs(1928));
    layer6_outputs(2248) <= not(layer5_outputs(6847));
    layer6_outputs(2249) <= (layer5_outputs(335)) xor (layer5_outputs(5828));
    layer6_outputs(2250) <= not(layer5_outputs(1582));
    layer6_outputs(2251) <= layer5_outputs(2973);
    layer6_outputs(2252) <= not(layer5_outputs(5180)) or (layer5_outputs(6570));
    layer6_outputs(2253) <= not(layer5_outputs(7161));
    layer6_outputs(2254) <= layer5_outputs(1859);
    layer6_outputs(2255) <= layer5_outputs(3661);
    layer6_outputs(2256) <= not(layer5_outputs(6709)) or (layer5_outputs(2466));
    layer6_outputs(2257) <= layer5_outputs(1175);
    layer6_outputs(2258) <= not(layer5_outputs(939));
    layer6_outputs(2259) <= not(layer5_outputs(201));
    layer6_outputs(2260) <= layer5_outputs(3653);
    layer6_outputs(2261) <= layer5_outputs(6633);
    layer6_outputs(2262) <= (layer5_outputs(6196)) and (layer5_outputs(4429));
    layer6_outputs(2263) <= not((layer5_outputs(7155)) xor (layer5_outputs(6761)));
    layer6_outputs(2264) <= layer5_outputs(7416);
    layer6_outputs(2265) <= not(layer5_outputs(532));
    layer6_outputs(2266) <= layer5_outputs(2604);
    layer6_outputs(2267) <= layer5_outputs(3817);
    layer6_outputs(2268) <= not(layer5_outputs(6592));
    layer6_outputs(2269) <= not((layer5_outputs(2966)) or (layer5_outputs(2644)));
    layer6_outputs(2270) <= not(layer5_outputs(881)) or (layer5_outputs(3545));
    layer6_outputs(2271) <= (layer5_outputs(3139)) xor (layer5_outputs(571));
    layer6_outputs(2272) <= not(layer5_outputs(2866)) or (layer5_outputs(2581));
    layer6_outputs(2273) <= not(layer5_outputs(888)) or (layer5_outputs(4703));
    layer6_outputs(2274) <= not(layer5_outputs(3590));
    layer6_outputs(2275) <= not((layer5_outputs(1765)) xor (layer5_outputs(5803)));
    layer6_outputs(2276) <= not(layer5_outputs(6076));
    layer6_outputs(2277) <= not(layer5_outputs(6198));
    layer6_outputs(2278) <= layer5_outputs(3497);
    layer6_outputs(2279) <= not(layer5_outputs(5767));
    layer6_outputs(2280) <= not(layer5_outputs(4645));
    layer6_outputs(2281) <= layer5_outputs(7359);
    layer6_outputs(2282) <= (layer5_outputs(2532)) and not (layer5_outputs(295));
    layer6_outputs(2283) <= layer5_outputs(6464);
    layer6_outputs(2284) <= layer5_outputs(2217);
    layer6_outputs(2285) <= not(layer5_outputs(4389));
    layer6_outputs(2286) <= layer5_outputs(6341);
    layer6_outputs(2287) <= not(layer5_outputs(6919)) or (layer5_outputs(3894));
    layer6_outputs(2288) <= (layer5_outputs(159)) and not (layer5_outputs(120));
    layer6_outputs(2289) <= (layer5_outputs(257)) xor (layer5_outputs(2437));
    layer6_outputs(2290) <= layer5_outputs(3854);
    layer6_outputs(2291) <= not(layer5_outputs(1915));
    layer6_outputs(2292) <= not(layer5_outputs(1897));
    layer6_outputs(2293) <= not(layer5_outputs(7348));
    layer6_outputs(2294) <= layer5_outputs(5388);
    layer6_outputs(2295) <= not((layer5_outputs(1955)) xor (layer5_outputs(5794)));
    layer6_outputs(2296) <= (layer5_outputs(2808)) and not (layer5_outputs(4734));
    layer6_outputs(2297) <= layer5_outputs(3990);
    layer6_outputs(2298) <= (layer5_outputs(1080)) and (layer5_outputs(5337));
    layer6_outputs(2299) <= (layer5_outputs(5735)) xor (layer5_outputs(5538));
    layer6_outputs(2300) <= not((layer5_outputs(6257)) xor (layer5_outputs(3256)));
    layer6_outputs(2301) <= layer5_outputs(5293);
    layer6_outputs(2302) <= (layer5_outputs(5072)) or (layer5_outputs(1145));
    layer6_outputs(2303) <= layer5_outputs(3113);
    layer6_outputs(2304) <= not((layer5_outputs(2618)) xor (layer5_outputs(3674)));
    layer6_outputs(2305) <= layer5_outputs(3430);
    layer6_outputs(2306) <= (layer5_outputs(6231)) xor (layer5_outputs(5245));
    layer6_outputs(2307) <= layer5_outputs(7526);
    layer6_outputs(2308) <= not((layer5_outputs(3086)) xor (layer5_outputs(6656)));
    layer6_outputs(2309) <= not(layer5_outputs(1756));
    layer6_outputs(2310) <= layer5_outputs(3652);
    layer6_outputs(2311) <= not(layer5_outputs(6820));
    layer6_outputs(2312) <= layer5_outputs(3748);
    layer6_outputs(2313) <= not(layer5_outputs(3657));
    layer6_outputs(2314) <= layer5_outputs(7353);
    layer6_outputs(2315) <= not((layer5_outputs(5671)) and (layer5_outputs(474)));
    layer6_outputs(2316) <= layer5_outputs(4177);
    layer6_outputs(2317) <= not(layer5_outputs(1989));
    layer6_outputs(2318) <= not((layer5_outputs(1545)) and (layer5_outputs(7080)));
    layer6_outputs(2319) <= not(layer5_outputs(4670));
    layer6_outputs(2320) <= layer5_outputs(6346);
    layer6_outputs(2321) <= not(layer5_outputs(4516)) or (layer5_outputs(4896));
    layer6_outputs(2322) <= '1';
    layer6_outputs(2323) <= not((layer5_outputs(3962)) or (layer5_outputs(2263)));
    layer6_outputs(2324) <= not(layer5_outputs(6985)) or (layer5_outputs(2079));
    layer6_outputs(2325) <= (layer5_outputs(3117)) and not (layer5_outputs(1505));
    layer6_outputs(2326) <= (layer5_outputs(7594)) and (layer5_outputs(5047));
    layer6_outputs(2327) <= layer5_outputs(6);
    layer6_outputs(2328) <= not((layer5_outputs(2990)) xor (layer5_outputs(5200)));
    layer6_outputs(2329) <= '0';
    layer6_outputs(2330) <= (layer5_outputs(2964)) and (layer5_outputs(385));
    layer6_outputs(2331) <= not(layer5_outputs(4916));
    layer6_outputs(2332) <= not(layer5_outputs(534));
    layer6_outputs(2333) <= (layer5_outputs(3596)) or (layer5_outputs(519));
    layer6_outputs(2334) <= not(layer5_outputs(3141)) or (layer5_outputs(5534));
    layer6_outputs(2335) <= (layer5_outputs(7505)) xor (layer5_outputs(3850));
    layer6_outputs(2336) <= layer5_outputs(2159);
    layer6_outputs(2337) <= layer5_outputs(5685);
    layer6_outputs(2338) <= (layer5_outputs(799)) and (layer5_outputs(6404));
    layer6_outputs(2339) <= (layer5_outputs(4735)) and not (layer5_outputs(3756));
    layer6_outputs(2340) <= not(layer5_outputs(2448));
    layer6_outputs(2341) <= not(layer5_outputs(259));
    layer6_outputs(2342) <= not(layer5_outputs(2022)) or (layer5_outputs(2070));
    layer6_outputs(2343) <= not(layer5_outputs(6668)) or (layer5_outputs(3217));
    layer6_outputs(2344) <= not((layer5_outputs(5553)) xor (layer5_outputs(5659)));
    layer6_outputs(2345) <= not(layer5_outputs(1227)) or (layer5_outputs(7464));
    layer6_outputs(2346) <= layer5_outputs(3888);
    layer6_outputs(2347) <= not(layer5_outputs(1576));
    layer6_outputs(2348) <= not(layer5_outputs(4503));
    layer6_outputs(2349) <= not((layer5_outputs(6357)) or (layer5_outputs(4346)));
    layer6_outputs(2350) <= (layer5_outputs(7045)) xor (layer5_outputs(7204));
    layer6_outputs(2351) <= not((layer5_outputs(540)) xor (layer5_outputs(7409)));
    layer6_outputs(2352) <= (layer5_outputs(4099)) or (layer5_outputs(5403));
    layer6_outputs(2353) <= layer5_outputs(4929);
    layer6_outputs(2354) <= not(layer5_outputs(5669));
    layer6_outputs(2355) <= not((layer5_outputs(5069)) xor (layer5_outputs(1098)));
    layer6_outputs(2356) <= not(layer5_outputs(7053)) or (layer5_outputs(6757));
    layer6_outputs(2357) <= layer5_outputs(2917);
    layer6_outputs(2358) <= (layer5_outputs(2360)) and not (layer5_outputs(4737));
    layer6_outputs(2359) <= not((layer5_outputs(7513)) and (layer5_outputs(5417)));
    layer6_outputs(2360) <= layer5_outputs(1509);
    layer6_outputs(2361) <= not(layer5_outputs(5731));
    layer6_outputs(2362) <= not((layer5_outputs(343)) xor (layer5_outputs(3036)));
    layer6_outputs(2363) <= layer5_outputs(1033);
    layer6_outputs(2364) <= not(layer5_outputs(1120));
    layer6_outputs(2365) <= not((layer5_outputs(6382)) or (layer5_outputs(878)));
    layer6_outputs(2366) <= layer5_outputs(6099);
    layer6_outputs(2367) <= (layer5_outputs(1967)) and (layer5_outputs(3175));
    layer6_outputs(2368) <= not(layer5_outputs(1392)) or (layer5_outputs(7453));
    layer6_outputs(2369) <= layer5_outputs(755);
    layer6_outputs(2370) <= not(layer5_outputs(4694));
    layer6_outputs(2371) <= layer5_outputs(2728);
    layer6_outputs(2372) <= not(layer5_outputs(7112));
    layer6_outputs(2373) <= layer5_outputs(130);
    layer6_outputs(2374) <= (layer5_outputs(2757)) and (layer5_outputs(2481));
    layer6_outputs(2375) <= not(layer5_outputs(5424)) or (layer5_outputs(2927));
    layer6_outputs(2376) <= not(layer5_outputs(3682));
    layer6_outputs(2377) <= layer5_outputs(5757);
    layer6_outputs(2378) <= (layer5_outputs(6575)) and not (layer5_outputs(5135));
    layer6_outputs(2379) <= layer5_outputs(5587);
    layer6_outputs(2380) <= not(layer5_outputs(5204));
    layer6_outputs(2381) <= layer5_outputs(3645);
    layer6_outputs(2382) <= not(layer5_outputs(4944));
    layer6_outputs(2383) <= layer5_outputs(423);
    layer6_outputs(2384) <= not(layer5_outputs(1933));
    layer6_outputs(2385) <= not(layer5_outputs(261));
    layer6_outputs(2386) <= not(layer5_outputs(5668));
    layer6_outputs(2387) <= not(layer5_outputs(6502));
    layer6_outputs(2388) <= not(layer5_outputs(589));
    layer6_outputs(2389) <= not(layer5_outputs(1674)) or (layer5_outputs(5121));
    layer6_outputs(2390) <= layer5_outputs(5159);
    layer6_outputs(2391) <= layer5_outputs(6536);
    layer6_outputs(2392) <= layer5_outputs(2760);
    layer6_outputs(2393) <= (layer5_outputs(3751)) and not (layer5_outputs(1565));
    layer6_outputs(2394) <= layer5_outputs(4590);
    layer6_outputs(2395) <= not((layer5_outputs(1621)) xor (layer5_outputs(6944)));
    layer6_outputs(2396) <= not(layer5_outputs(4113));
    layer6_outputs(2397) <= not(layer5_outputs(7381));
    layer6_outputs(2398) <= not((layer5_outputs(6803)) xor (layer5_outputs(5134)));
    layer6_outputs(2399) <= not((layer5_outputs(2216)) xor (layer5_outputs(25)));
    layer6_outputs(2400) <= not(layer5_outputs(2805));
    layer6_outputs(2401) <= layer5_outputs(4486);
    layer6_outputs(2402) <= not((layer5_outputs(4386)) or (layer5_outputs(7282)));
    layer6_outputs(2403) <= layer5_outputs(1595);
    layer6_outputs(2404) <= layer5_outputs(5857);
    layer6_outputs(2405) <= (layer5_outputs(6403)) and not (layer5_outputs(7652));
    layer6_outputs(2406) <= not((layer5_outputs(3412)) or (layer5_outputs(5566)));
    layer6_outputs(2407) <= not(layer5_outputs(3946));
    layer6_outputs(2408) <= layer5_outputs(1350);
    layer6_outputs(2409) <= not(layer5_outputs(4644));
    layer6_outputs(2410) <= not(layer5_outputs(1883));
    layer6_outputs(2411) <= layer5_outputs(2028);
    layer6_outputs(2412) <= (layer5_outputs(3966)) xor (layer5_outputs(880));
    layer6_outputs(2413) <= not((layer5_outputs(1596)) and (layer5_outputs(2673)));
    layer6_outputs(2414) <= layer5_outputs(5345);
    layer6_outputs(2415) <= layer5_outputs(5855);
    layer6_outputs(2416) <= layer5_outputs(3009);
    layer6_outputs(2417) <= layer5_outputs(601);
    layer6_outputs(2418) <= (layer5_outputs(3924)) and not (layer5_outputs(5693));
    layer6_outputs(2419) <= not(layer5_outputs(633));
    layer6_outputs(2420) <= not(layer5_outputs(131)) or (layer5_outputs(7256));
    layer6_outputs(2421) <= not((layer5_outputs(4989)) or (layer5_outputs(1454)));
    layer6_outputs(2422) <= layer5_outputs(5186);
    layer6_outputs(2423) <= (layer5_outputs(451)) xor (layer5_outputs(6443));
    layer6_outputs(2424) <= layer5_outputs(1939);
    layer6_outputs(2425) <= not((layer5_outputs(5628)) xor (layer5_outputs(5102)));
    layer6_outputs(2426) <= (layer5_outputs(2300)) or (layer5_outputs(6644));
    layer6_outputs(2427) <= not(layer5_outputs(3874));
    layer6_outputs(2428) <= layer5_outputs(893);
    layer6_outputs(2429) <= not(layer5_outputs(4078));
    layer6_outputs(2430) <= (layer5_outputs(7399)) xor (layer5_outputs(836));
    layer6_outputs(2431) <= not(layer5_outputs(248));
    layer6_outputs(2432) <= not((layer5_outputs(6084)) or (layer5_outputs(2643)));
    layer6_outputs(2433) <= not((layer5_outputs(3735)) and (layer5_outputs(169)));
    layer6_outputs(2434) <= layer5_outputs(7535);
    layer6_outputs(2435) <= not((layer5_outputs(3297)) or (layer5_outputs(2478)));
    layer6_outputs(2436) <= layer5_outputs(602);
    layer6_outputs(2437) <= not(layer5_outputs(2921));
    layer6_outputs(2438) <= not(layer5_outputs(4276));
    layer6_outputs(2439) <= (layer5_outputs(6289)) or (layer5_outputs(2586));
    layer6_outputs(2440) <= not((layer5_outputs(1182)) xor (layer5_outputs(5676)));
    layer6_outputs(2441) <= not(layer5_outputs(5233));
    layer6_outputs(2442) <= not(layer5_outputs(6282));
    layer6_outputs(2443) <= (layer5_outputs(6508)) and not (layer5_outputs(7280));
    layer6_outputs(2444) <= layer5_outputs(5408);
    layer6_outputs(2445) <= not((layer5_outputs(1744)) xor (layer5_outputs(4754)));
    layer6_outputs(2446) <= '1';
    layer6_outputs(2447) <= not((layer5_outputs(4184)) xor (layer5_outputs(4651)));
    layer6_outputs(2448) <= layer5_outputs(2399);
    layer6_outputs(2449) <= not((layer5_outputs(1218)) xor (layer5_outputs(5170)));
    layer6_outputs(2450) <= (layer5_outputs(4861)) xor (layer5_outputs(3592));
    layer6_outputs(2451) <= layer5_outputs(2396);
    layer6_outputs(2452) <= layer5_outputs(4229);
    layer6_outputs(2453) <= layer5_outputs(2642);
    layer6_outputs(2454) <= layer5_outputs(2350);
    layer6_outputs(2455) <= not(layer5_outputs(7046));
    layer6_outputs(2456) <= (layer5_outputs(6664)) and not (layer5_outputs(3151));
    layer6_outputs(2457) <= not((layer5_outputs(2824)) or (layer5_outputs(2632)));
    layer6_outputs(2458) <= layer5_outputs(1858);
    layer6_outputs(2459) <= not(layer5_outputs(1799));
    layer6_outputs(2460) <= not(layer5_outputs(2316)) or (layer5_outputs(24));
    layer6_outputs(2461) <= (layer5_outputs(2517)) and not (layer5_outputs(1896));
    layer6_outputs(2462) <= not(layer5_outputs(1064));
    layer6_outputs(2463) <= (layer5_outputs(1837)) xor (layer5_outputs(7288));
    layer6_outputs(2464) <= layer5_outputs(6954);
    layer6_outputs(2465) <= not((layer5_outputs(3838)) and (layer5_outputs(4571)));
    layer6_outputs(2466) <= not(layer5_outputs(839)) or (layer5_outputs(6954));
    layer6_outputs(2467) <= not(layer5_outputs(4759));
    layer6_outputs(2468) <= (layer5_outputs(6366)) xor (layer5_outputs(2181));
    layer6_outputs(2469) <= layer5_outputs(7384);
    layer6_outputs(2470) <= (layer5_outputs(3696)) and not (layer5_outputs(899));
    layer6_outputs(2471) <= layer5_outputs(5310);
    layer6_outputs(2472) <= (layer5_outputs(3102)) xor (layer5_outputs(2051));
    layer6_outputs(2473) <= not(layer5_outputs(1142));
    layer6_outputs(2474) <= (layer5_outputs(587)) xor (layer5_outputs(4757));
    layer6_outputs(2475) <= layer5_outputs(1794);
    layer6_outputs(2476) <= not(layer5_outputs(1819));
    layer6_outputs(2477) <= not(layer5_outputs(2473));
    layer6_outputs(2478) <= (layer5_outputs(924)) or (layer5_outputs(4263));
    layer6_outputs(2479) <= (layer5_outputs(1907)) and not (layer5_outputs(5239));
    layer6_outputs(2480) <= '1';
    layer6_outputs(2481) <= layer5_outputs(641);
    layer6_outputs(2482) <= layer5_outputs(6212);
    layer6_outputs(2483) <= not((layer5_outputs(696)) xor (layer5_outputs(2419)));
    layer6_outputs(2484) <= layer5_outputs(5387);
    layer6_outputs(2485) <= layer5_outputs(6212);
    layer6_outputs(2486) <= not((layer5_outputs(2794)) xor (layer5_outputs(2143)));
    layer6_outputs(2487) <= (layer5_outputs(5889)) or (layer5_outputs(7208));
    layer6_outputs(2488) <= layer5_outputs(517);
    layer6_outputs(2489) <= not(layer5_outputs(1719));
    layer6_outputs(2490) <= not(layer5_outputs(4166));
    layer6_outputs(2491) <= (layer5_outputs(5722)) xor (layer5_outputs(3543));
    layer6_outputs(2492) <= (layer5_outputs(5412)) and (layer5_outputs(563));
    layer6_outputs(2493) <= not(layer5_outputs(2032)) or (layer5_outputs(6535));
    layer6_outputs(2494) <= layer5_outputs(7628);
    layer6_outputs(2495) <= not(layer5_outputs(3004)) or (layer5_outputs(1647));
    layer6_outputs(2496) <= (layer5_outputs(6527)) xor (layer5_outputs(4799));
    layer6_outputs(2497) <= not(layer5_outputs(2708));
    layer6_outputs(2498) <= not(layer5_outputs(2681));
    layer6_outputs(2499) <= not(layer5_outputs(3540));
    layer6_outputs(2500) <= layer5_outputs(4751);
    layer6_outputs(2501) <= not((layer5_outputs(4994)) or (layer5_outputs(3917)));
    layer6_outputs(2502) <= layer5_outputs(3049);
    layer6_outputs(2503) <= not(layer5_outputs(3402));
    layer6_outputs(2504) <= not(layer5_outputs(5261));
    layer6_outputs(2505) <= not(layer5_outputs(108));
    layer6_outputs(2506) <= not((layer5_outputs(674)) xor (layer5_outputs(4971)));
    layer6_outputs(2507) <= (layer5_outputs(3512)) and not (layer5_outputs(3245));
    layer6_outputs(2508) <= not((layer5_outputs(2372)) or (layer5_outputs(7218)));
    layer6_outputs(2509) <= not(layer5_outputs(2099));
    layer6_outputs(2510) <= not(layer5_outputs(6563));
    layer6_outputs(2511) <= not(layer5_outputs(7030));
    layer6_outputs(2512) <= (layer5_outputs(5238)) or (layer5_outputs(31));
    layer6_outputs(2513) <= layer5_outputs(4406);
    layer6_outputs(2514) <= not(layer5_outputs(1353));
    layer6_outputs(2515) <= not((layer5_outputs(4231)) or (layer5_outputs(7413)));
    layer6_outputs(2516) <= layer5_outputs(7666);
    layer6_outputs(2517) <= (layer5_outputs(5374)) xor (layer5_outputs(5802));
    layer6_outputs(2518) <= not((layer5_outputs(6454)) xor (layer5_outputs(6230)));
    layer6_outputs(2519) <= layer5_outputs(6142);
    layer6_outputs(2520) <= (layer5_outputs(5315)) and (layer5_outputs(2594));
    layer6_outputs(2521) <= not((layer5_outputs(1327)) xor (layer5_outputs(6560)));
    layer6_outputs(2522) <= layer5_outputs(4518);
    layer6_outputs(2523) <= (layer5_outputs(6144)) and not (layer5_outputs(644));
    layer6_outputs(2524) <= layer5_outputs(5910);
    layer6_outputs(2525) <= not(layer5_outputs(5781));
    layer6_outputs(2526) <= not(layer5_outputs(2695));
    layer6_outputs(2527) <= (layer5_outputs(4236)) and not (layer5_outputs(5568));
    layer6_outputs(2528) <= not((layer5_outputs(5985)) xor (layer5_outputs(4796)));
    layer6_outputs(2529) <= not(layer5_outputs(3421));
    layer6_outputs(2530) <= layer5_outputs(6857);
    layer6_outputs(2531) <= not(layer5_outputs(5905));
    layer6_outputs(2532) <= (layer5_outputs(2609)) xor (layer5_outputs(812));
    layer6_outputs(2533) <= not((layer5_outputs(3718)) xor (layer5_outputs(576)));
    layer6_outputs(2534) <= layer5_outputs(7422);
    layer6_outputs(2535) <= layer5_outputs(2684);
    layer6_outputs(2536) <= not((layer5_outputs(2675)) xor (layer5_outputs(1134)));
    layer6_outputs(2537) <= not(layer5_outputs(3819)) or (layer5_outputs(1043));
    layer6_outputs(2538) <= not(layer5_outputs(4285));
    layer6_outputs(2539) <= layer5_outputs(1645);
    layer6_outputs(2540) <= not(layer5_outputs(7234));
    layer6_outputs(2541) <= layer5_outputs(2087);
    layer6_outputs(2542) <= not(layer5_outputs(4312));
    layer6_outputs(2543) <= not((layer5_outputs(5522)) and (layer5_outputs(1018)));
    layer6_outputs(2544) <= layer5_outputs(1224);
    layer6_outputs(2545) <= (layer5_outputs(1690)) xor (layer5_outputs(4382));
    layer6_outputs(2546) <= not((layer5_outputs(6530)) or (layer5_outputs(6132)));
    layer6_outputs(2547) <= not(layer5_outputs(1133));
    layer6_outputs(2548) <= (layer5_outputs(6492)) or (layer5_outputs(3726));
    layer6_outputs(2549) <= not(layer5_outputs(3579));
    layer6_outputs(2550) <= not(layer5_outputs(4166)) or (layer5_outputs(3314));
    layer6_outputs(2551) <= layer5_outputs(1100);
    layer6_outputs(2552) <= (layer5_outputs(4845)) or (layer5_outputs(1666));
    layer6_outputs(2553) <= not((layer5_outputs(4557)) and (layer5_outputs(7201)));
    layer6_outputs(2554) <= layer5_outputs(446);
    layer6_outputs(2555) <= layer5_outputs(150);
    layer6_outputs(2556) <= not(layer5_outputs(895));
    layer6_outputs(2557) <= layer5_outputs(7475);
    layer6_outputs(2558) <= not(layer5_outputs(6011));
    layer6_outputs(2559) <= not(layer5_outputs(6900)) or (layer5_outputs(6429));
    layer6_outputs(2560) <= (layer5_outputs(5554)) xor (layer5_outputs(1044));
    layer6_outputs(2561) <= not(layer5_outputs(733));
    layer6_outputs(2562) <= layer5_outputs(4832);
    layer6_outputs(2563) <= not((layer5_outputs(832)) and (layer5_outputs(3879)));
    layer6_outputs(2564) <= not(layer5_outputs(6228));
    layer6_outputs(2565) <= not((layer5_outputs(1946)) xor (layer5_outputs(2126)));
    layer6_outputs(2566) <= (layer5_outputs(5687)) and not (layer5_outputs(3617));
    layer6_outputs(2567) <= not(layer5_outputs(2393));
    layer6_outputs(2568) <= not(layer5_outputs(637)) or (layer5_outputs(3532));
    layer6_outputs(2569) <= not(layer5_outputs(1405)) or (layer5_outputs(112));
    layer6_outputs(2570) <= not((layer5_outputs(6123)) xor (layer5_outputs(606)));
    layer6_outputs(2571) <= layer5_outputs(2807);
    layer6_outputs(2572) <= (layer5_outputs(7619)) xor (layer5_outputs(824));
    layer6_outputs(2573) <= not(layer5_outputs(89));
    layer6_outputs(2574) <= (layer5_outputs(4978)) and (layer5_outputs(3091));
    layer6_outputs(2575) <= layer5_outputs(1784);
    layer6_outputs(2576) <= not((layer5_outputs(987)) or (layer5_outputs(207)));
    layer6_outputs(2577) <= layer5_outputs(437);
    layer6_outputs(2578) <= (layer5_outputs(6687)) xor (layer5_outputs(7113));
    layer6_outputs(2579) <= not(layer5_outputs(3961));
    layer6_outputs(2580) <= layer5_outputs(6852);
    layer6_outputs(2581) <= layer5_outputs(2425);
    layer6_outputs(2582) <= (layer5_outputs(2631)) and not (layer5_outputs(1723));
    layer6_outputs(2583) <= not(layer5_outputs(5232));
    layer6_outputs(2584) <= not((layer5_outputs(1331)) xor (layer5_outputs(5884)));
    layer6_outputs(2585) <= not(layer5_outputs(4269));
    layer6_outputs(2586) <= not((layer5_outputs(1944)) xor (layer5_outputs(1423)));
    layer6_outputs(2587) <= (layer5_outputs(1062)) or (layer5_outputs(6686));
    layer6_outputs(2588) <= layer5_outputs(4533);
    layer6_outputs(2589) <= not(layer5_outputs(4185));
    layer6_outputs(2590) <= (layer5_outputs(3128)) xor (layer5_outputs(6324));
    layer6_outputs(2591) <= '0';
    layer6_outputs(2592) <= not(layer5_outputs(2926));
    layer6_outputs(2593) <= not(layer5_outputs(2477));
    layer6_outputs(2594) <= layer5_outputs(5636);
    layer6_outputs(2595) <= not(layer5_outputs(2448));
    layer6_outputs(2596) <= not(layer5_outputs(3467));
    layer6_outputs(2597) <= layer5_outputs(482);
    layer6_outputs(2598) <= not(layer5_outputs(4110));
    layer6_outputs(2599) <= not(layer5_outputs(7040)) or (layer5_outputs(831));
    layer6_outputs(2600) <= (layer5_outputs(7226)) xor (layer5_outputs(3152));
    layer6_outputs(2601) <= (layer5_outputs(7461)) xor (layer5_outputs(2028));
    layer6_outputs(2602) <= not(layer5_outputs(5934));
    layer6_outputs(2603) <= not(layer5_outputs(6043));
    layer6_outputs(2604) <= not((layer5_outputs(2596)) and (layer5_outputs(6836)));
    layer6_outputs(2605) <= (layer5_outputs(11)) xor (layer5_outputs(2389));
    layer6_outputs(2606) <= (layer5_outputs(258)) and not (layer5_outputs(5603));
    layer6_outputs(2607) <= (layer5_outputs(5548)) xor (layer5_outputs(7525));
    layer6_outputs(2608) <= (layer5_outputs(222)) xor (layer5_outputs(3782));
    layer6_outputs(2609) <= not((layer5_outputs(5846)) xor (layer5_outputs(1923)));
    layer6_outputs(2610) <= not(layer5_outputs(2194));
    layer6_outputs(2611) <= (layer5_outputs(4631)) xor (layer5_outputs(2021));
    layer6_outputs(2612) <= '0';
    layer6_outputs(2613) <= not((layer5_outputs(5009)) or (layer5_outputs(1197)));
    layer6_outputs(2614) <= layer5_outputs(1849);
    layer6_outputs(2615) <= not((layer5_outputs(7485)) xor (layer5_outputs(3309)));
    layer6_outputs(2616) <= layer5_outputs(4453);
    layer6_outputs(2617) <= '1';
    layer6_outputs(2618) <= not(layer5_outputs(1280));
    layer6_outputs(2619) <= not(layer5_outputs(2025));
    layer6_outputs(2620) <= not(layer5_outputs(6160));
    layer6_outputs(2621) <= (layer5_outputs(5476)) xor (layer5_outputs(6052));
    layer6_outputs(2622) <= layer5_outputs(4271);
    layer6_outputs(2623) <= not((layer5_outputs(4406)) and (layer5_outputs(2086)));
    layer6_outputs(2624) <= not((layer5_outputs(7491)) and (layer5_outputs(4967)));
    layer6_outputs(2625) <= not(layer5_outputs(6613));
    layer6_outputs(2626) <= not(layer5_outputs(2453));
    layer6_outputs(2627) <= not((layer5_outputs(2456)) xor (layer5_outputs(4545)));
    layer6_outputs(2628) <= not((layer5_outputs(1255)) xor (layer5_outputs(6299)));
    layer6_outputs(2629) <= not(layer5_outputs(1856));
    layer6_outputs(2630) <= (layer5_outputs(3969)) and not (layer5_outputs(4458));
    layer6_outputs(2631) <= not(layer5_outputs(4312));
    layer6_outputs(2632) <= not(layer5_outputs(5433));
    layer6_outputs(2633) <= not((layer5_outputs(3985)) xor (layer5_outputs(6423)));
    layer6_outputs(2634) <= (layer5_outputs(218)) and (layer5_outputs(4073));
    layer6_outputs(2635) <= not(layer5_outputs(2948));
    layer6_outputs(2636) <= (layer5_outputs(6928)) and (layer5_outputs(1370));
    layer6_outputs(2637) <= not(layer5_outputs(3012)) or (layer5_outputs(4800));
    layer6_outputs(2638) <= not(layer5_outputs(6089));
    layer6_outputs(2639) <= layer5_outputs(1081);
    layer6_outputs(2640) <= layer5_outputs(2962);
    layer6_outputs(2641) <= not((layer5_outputs(6604)) or (layer5_outputs(3093)));
    layer6_outputs(2642) <= layer5_outputs(6482);
    layer6_outputs(2643) <= not(layer5_outputs(2866));
    layer6_outputs(2644) <= not(layer5_outputs(3995));
    layer6_outputs(2645) <= layer5_outputs(3829);
    layer6_outputs(2646) <= (layer5_outputs(1664)) xor (layer5_outputs(2525));
    layer6_outputs(2647) <= not(layer5_outputs(1491));
    layer6_outputs(2648) <= layer5_outputs(6006);
    layer6_outputs(2649) <= layer5_outputs(762);
    layer6_outputs(2650) <= not(layer5_outputs(6495)) or (layer5_outputs(7633));
    layer6_outputs(2651) <= not(layer5_outputs(1383));
    layer6_outputs(2652) <= layer5_outputs(7305);
    layer6_outputs(2653) <= not((layer5_outputs(1662)) xor (layer5_outputs(1895)));
    layer6_outputs(2654) <= not(layer5_outputs(3247));
    layer6_outputs(2655) <= (layer5_outputs(5763)) and not (layer5_outputs(4943));
    layer6_outputs(2656) <= not(layer5_outputs(2302));
    layer6_outputs(2657) <= not(layer5_outputs(2418));
    layer6_outputs(2658) <= (layer5_outputs(362)) xor (layer5_outputs(4047));
    layer6_outputs(2659) <= (layer5_outputs(5854)) xor (layer5_outputs(3422));
    layer6_outputs(2660) <= not(layer5_outputs(5560)) or (layer5_outputs(5183));
    layer6_outputs(2661) <= not(layer5_outputs(3331)) or (layer5_outputs(245));
    layer6_outputs(2662) <= not(layer5_outputs(3391));
    layer6_outputs(2663) <= not((layer5_outputs(4018)) xor (layer5_outputs(4450)));
    layer6_outputs(2664) <= not(layer5_outputs(3900));
    layer6_outputs(2665) <= layer5_outputs(5360);
    layer6_outputs(2666) <= not(layer5_outputs(6553));
    layer6_outputs(2667) <= not(layer5_outputs(4072));
    layer6_outputs(2668) <= layer5_outputs(7014);
    layer6_outputs(2669) <= not((layer5_outputs(5840)) and (layer5_outputs(2351)));
    layer6_outputs(2670) <= (layer5_outputs(6891)) and not (layer5_outputs(2331));
    layer6_outputs(2671) <= not(layer5_outputs(5758));
    layer6_outputs(2672) <= not(layer5_outputs(4164));
    layer6_outputs(2673) <= not(layer5_outputs(4215));
    layer6_outputs(2674) <= not(layer5_outputs(6533));
    layer6_outputs(2675) <= not(layer5_outputs(5879));
    layer6_outputs(2676) <= (layer5_outputs(6918)) and (layer5_outputs(4017));
    layer6_outputs(2677) <= (layer5_outputs(4867)) and not (layer5_outputs(4474));
    layer6_outputs(2678) <= not((layer5_outputs(4451)) xor (layer5_outputs(4912)));
    layer6_outputs(2679) <= not((layer5_outputs(2653)) xor (layer5_outputs(1834)));
    layer6_outputs(2680) <= not((layer5_outputs(4007)) xor (layer5_outputs(3656)));
    layer6_outputs(2681) <= (layer5_outputs(3516)) and not (layer5_outputs(1676));
    layer6_outputs(2682) <= not((layer5_outputs(6473)) and (layer5_outputs(6385)));
    layer6_outputs(2683) <= not(layer5_outputs(3370));
    layer6_outputs(2684) <= layer5_outputs(2432);
    layer6_outputs(2685) <= not(layer5_outputs(948));
    layer6_outputs(2686) <= (layer5_outputs(5543)) and (layer5_outputs(5252));
    layer6_outputs(2687) <= layer5_outputs(5750);
    layer6_outputs(2688) <= layer5_outputs(2289);
    layer6_outputs(2689) <= (layer5_outputs(1566)) and not (layer5_outputs(6990));
    layer6_outputs(2690) <= layer5_outputs(1202);
    layer6_outputs(2691) <= layer5_outputs(2273);
    layer6_outputs(2692) <= not(layer5_outputs(368));
    layer6_outputs(2693) <= layer5_outputs(7333);
    layer6_outputs(2694) <= (layer5_outputs(2111)) xor (layer5_outputs(6608));
    layer6_outputs(2695) <= layer5_outputs(5896);
    layer6_outputs(2696) <= not(layer5_outputs(2953));
    layer6_outputs(2697) <= not(layer5_outputs(3304)) or (layer5_outputs(3608));
    layer6_outputs(2698) <= layer5_outputs(2768);
    layer6_outputs(2699) <= layer5_outputs(726);
    layer6_outputs(2700) <= layer5_outputs(392);
    layer6_outputs(2701) <= not((layer5_outputs(1932)) xor (layer5_outputs(4175)));
    layer6_outputs(2702) <= layer5_outputs(833);
    layer6_outputs(2703) <= (layer5_outputs(622)) or (layer5_outputs(7158));
    layer6_outputs(2704) <= (layer5_outputs(1123)) and (layer5_outputs(6047));
    layer6_outputs(2705) <= not(layer5_outputs(5113)) or (layer5_outputs(4593));
    layer6_outputs(2706) <= not(layer5_outputs(971));
    layer6_outputs(2707) <= (layer5_outputs(2652)) and not (layer5_outputs(6204));
    layer6_outputs(2708) <= not(layer5_outputs(4676));
    layer6_outputs(2709) <= (layer5_outputs(3252)) and (layer5_outputs(1258));
    layer6_outputs(2710) <= not(layer5_outputs(2428));
    layer6_outputs(2711) <= layer5_outputs(3611);
    layer6_outputs(2712) <= layer5_outputs(5841);
    layer6_outputs(2713) <= layer5_outputs(3742);
    layer6_outputs(2714) <= (layer5_outputs(839)) or (layer5_outputs(2269));
    layer6_outputs(2715) <= not(layer5_outputs(4262));
    layer6_outputs(2716) <= not(layer5_outputs(6507));
    layer6_outputs(2717) <= not((layer5_outputs(5545)) xor (layer5_outputs(992)));
    layer6_outputs(2718) <= not(layer5_outputs(6300));
    layer6_outputs(2719) <= not((layer5_outputs(3660)) or (layer5_outputs(2569)));
    layer6_outputs(2720) <= layer5_outputs(1480);
    layer6_outputs(2721) <= (layer5_outputs(7103)) xor (layer5_outputs(4287));
    layer6_outputs(2722) <= layer5_outputs(4353);
    layer6_outputs(2723) <= layer5_outputs(484);
    layer6_outputs(2724) <= layer5_outputs(1199);
    layer6_outputs(2725) <= not(layer5_outputs(3694));
    layer6_outputs(2726) <= not((layer5_outputs(2510)) xor (layer5_outputs(1271)));
    layer6_outputs(2727) <= (layer5_outputs(187)) and (layer5_outputs(630));
    layer6_outputs(2728) <= not(layer5_outputs(6650));
    layer6_outputs(2729) <= not(layer5_outputs(5882)) or (layer5_outputs(7432));
    layer6_outputs(2730) <= not((layer5_outputs(4810)) xor (layer5_outputs(7104)));
    layer6_outputs(2731) <= layer5_outputs(7520);
    layer6_outputs(2732) <= not((layer5_outputs(1865)) or (layer5_outputs(6801)));
    layer6_outputs(2733) <= not(layer5_outputs(2942));
    layer6_outputs(2734) <= not(layer5_outputs(7143));
    layer6_outputs(2735) <= layer5_outputs(783);
    layer6_outputs(2736) <= not(layer5_outputs(5684)) or (layer5_outputs(535));
    layer6_outputs(2737) <= (layer5_outputs(7474)) and not (layer5_outputs(3503));
    layer6_outputs(2738) <= not(layer5_outputs(1181));
    layer6_outputs(2739) <= layer5_outputs(7414);
    layer6_outputs(2740) <= layer5_outputs(2290);
    layer6_outputs(2741) <= not(layer5_outputs(2268));
    layer6_outputs(2742) <= not(layer5_outputs(758));
    layer6_outputs(2743) <= layer5_outputs(6407);
    layer6_outputs(2744) <= layer5_outputs(7460);
    layer6_outputs(2745) <= not(layer5_outputs(5001));
    layer6_outputs(2746) <= (layer5_outputs(1161)) xor (layer5_outputs(3340));
    layer6_outputs(2747) <= (layer5_outputs(3525)) and not (layer5_outputs(7109));
    layer6_outputs(2748) <= (layer5_outputs(1224)) and not (layer5_outputs(5411));
    layer6_outputs(2749) <= not(layer5_outputs(3092));
    layer6_outputs(2750) <= (layer5_outputs(1764)) xor (layer5_outputs(7222));
    layer6_outputs(2751) <= layer5_outputs(3867);
    layer6_outputs(2752) <= (layer5_outputs(5805)) and (layer5_outputs(7050));
    layer6_outputs(2753) <= not((layer5_outputs(4424)) xor (layer5_outputs(1604)));
    layer6_outputs(2754) <= not(layer5_outputs(1018));
    layer6_outputs(2755) <= not((layer5_outputs(5195)) and (layer5_outputs(3861)));
    layer6_outputs(2756) <= not(layer5_outputs(296)) or (layer5_outputs(6728));
    layer6_outputs(2757) <= not((layer5_outputs(5705)) and (layer5_outputs(3493)));
    layer6_outputs(2758) <= (layer5_outputs(6405)) or (layer5_outputs(7215));
    layer6_outputs(2759) <= layer5_outputs(4109);
    layer6_outputs(2760) <= not(layer5_outputs(3222)) or (layer5_outputs(4220));
    layer6_outputs(2761) <= not(layer5_outputs(2847));
    layer6_outputs(2762) <= layer5_outputs(5066);
    layer6_outputs(2763) <= (layer5_outputs(7027)) xor (layer5_outputs(4903));
    layer6_outputs(2764) <= layer5_outputs(6865);
    layer6_outputs(2765) <= layer5_outputs(7326);
    layer6_outputs(2766) <= not(layer5_outputs(2074)) or (layer5_outputs(115));
    layer6_outputs(2767) <= not(layer5_outputs(938));
    layer6_outputs(2768) <= layer5_outputs(818);
    layer6_outputs(2769) <= '1';
    layer6_outputs(2770) <= layer5_outputs(2193);
    layer6_outputs(2771) <= (layer5_outputs(1181)) xor (layer5_outputs(2911));
    layer6_outputs(2772) <= (layer5_outputs(1490)) and not (layer5_outputs(456));
    layer6_outputs(2773) <= not(layer5_outputs(5976)) or (layer5_outputs(6464));
    layer6_outputs(2774) <= layer5_outputs(5750);
    layer6_outputs(2775) <= not(layer5_outputs(3479));
    layer6_outputs(2776) <= layer5_outputs(4791);
    layer6_outputs(2777) <= not(layer5_outputs(2825));
    layer6_outputs(2778) <= (layer5_outputs(4313)) or (layer5_outputs(3085));
    layer6_outputs(2779) <= not(layer5_outputs(799));
    layer6_outputs(2780) <= layer5_outputs(2432);
    layer6_outputs(2781) <= layer5_outputs(1540);
    layer6_outputs(2782) <= layer5_outputs(7195);
    layer6_outputs(2783) <= not(layer5_outputs(7294));
    layer6_outputs(2784) <= (layer5_outputs(5358)) and not (layer5_outputs(4727));
    layer6_outputs(2785) <= (layer5_outputs(6952)) xor (layer5_outputs(2038));
    layer6_outputs(2786) <= not(layer5_outputs(3158));
    layer6_outputs(2787) <= not(layer5_outputs(2762));
    layer6_outputs(2788) <= not(layer5_outputs(7065));
    layer6_outputs(2789) <= (layer5_outputs(3794)) and (layer5_outputs(3840));
    layer6_outputs(2790) <= (layer5_outputs(503)) xor (layer5_outputs(7516));
    layer6_outputs(2791) <= layer5_outputs(3044);
    layer6_outputs(2792) <= not(layer5_outputs(6075)) or (layer5_outputs(5333));
    layer6_outputs(2793) <= layer5_outputs(7297);
    layer6_outputs(2794) <= not((layer5_outputs(7403)) xor (layer5_outputs(782)));
    layer6_outputs(2795) <= layer5_outputs(4906);
    layer6_outputs(2796) <= not((layer5_outputs(7318)) xor (layer5_outputs(4069)));
    layer6_outputs(2797) <= not((layer5_outputs(6830)) xor (layer5_outputs(6596)));
    layer6_outputs(2798) <= not((layer5_outputs(2030)) xor (layer5_outputs(5193)));
    layer6_outputs(2799) <= not(layer5_outputs(5441));
    layer6_outputs(2800) <= layer5_outputs(5958);
    layer6_outputs(2801) <= not((layer5_outputs(5045)) or (layer5_outputs(3186)));
    layer6_outputs(2802) <= not(layer5_outputs(6316));
    layer6_outputs(2803) <= (layer5_outputs(4821)) and not (layer5_outputs(546));
    layer6_outputs(2804) <= not(layer5_outputs(6630));
    layer6_outputs(2805) <= not(layer5_outputs(631));
    layer6_outputs(2806) <= layer5_outputs(1613);
    layer6_outputs(2807) <= not(layer5_outputs(1775)) or (layer5_outputs(5491));
    layer6_outputs(2808) <= (layer5_outputs(6703)) and not (layer5_outputs(7483));
    layer6_outputs(2809) <= (layer5_outputs(5148)) and not (layer5_outputs(42));
    layer6_outputs(2810) <= (layer5_outputs(5137)) xor (layer5_outputs(4079));
    layer6_outputs(2811) <= layer5_outputs(2101);
    layer6_outputs(2812) <= not(layer5_outputs(4597));
    layer6_outputs(2813) <= not((layer5_outputs(4161)) xor (layer5_outputs(1186)));
    layer6_outputs(2814) <= not(layer5_outputs(4077));
    layer6_outputs(2815) <= not(layer5_outputs(1558));
    layer6_outputs(2816) <= layer5_outputs(1917);
    layer6_outputs(2817) <= (layer5_outputs(5027)) and not (layer5_outputs(6095));
    layer6_outputs(2818) <= layer5_outputs(7426);
    layer6_outputs(2819) <= not((layer5_outputs(3742)) or (layer5_outputs(3601)));
    layer6_outputs(2820) <= layer5_outputs(1213);
    layer6_outputs(2821) <= not((layer5_outputs(516)) xor (layer5_outputs(1083)));
    layer6_outputs(2822) <= not(layer5_outputs(886));
    layer6_outputs(2823) <= not(layer5_outputs(7346));
    layer6_outputs(2824) <= not(layer5_outputs(220));
    layer6_outputs(2825) <= (layer5_outputs(6401)) and (layer5_outputs(6915));
    layer6_outputs(2826) <= layer5_outputs(3143);
    layer6_outputs(2827) <= layer5_outputs(6534);
    layer6_outputs(2828) <= (layer5_outputs(7117)) and (layer5_outputs(4157));
    layer6_outputs(2829) <= not((layer5_outputs(6371)) and (layer5_outputs(1268)));
    layer6_outputs(2830) <= not(layer5_outputs(4609));
    layer6_outputs(2831) <= layer5_outputs(1989);
    layer6_outputs(2832) <= (layer5_outputs(2958)) and not (layer5_outputs(3974));
    layer6_outputs(2833) <= not(layer5_outputs(5152));
    layer6_outputs(2834) <= '1';
    layer6_outputs(2835) <= not((layer5_outputs(4461)) xor (layer5_outputs(3981)));
    layer6_outputs(2836) <= not(layer5_outputs(3603));
    layer6_outputs(2837) <= not((layer5_outputs(5932)) xor (layer5_outputs(4024)));
    layer6_outputs(2838) <= layer5_outputs(5647);
    layer6_outputs(2839) <= not((layer5_outputs(4634)) xor (layer5_outputs(2007)));
    layer6_outputs(2840) <= not(layer5_outputs(6946));
    layer6_outputs(2841) <= not((layer5_outputs(3872)) or (layer5_outputs(1401)));
    layer6_outputs(2842) <= layer5_outputs(439);
    layer6_outputs(2843) <= '1';
    layer6_outputs(2844) <= not(layer5_outputs(5701));
    layer6_outputs(2845) <= (layer5_outputs(4778)) xor (layer5_outputs(3985));
    layer6_outputs(2846) <= (layer5_outputs(6469)) xor (layer5_outputs(947));
    layer6_outputs(2847) <= not((layer5_outputs(6821)) or (layer5_outputs(3049)));
    layer6_outputs(2848) <= layer5_outputs(6557);
    layer6_outputs(2849) <= (layer5_outputs(4107)) and (layer5_outputs(2162));
    layer6_outputs(2850) <= (layer5_outputs(6548)) and not (layer5_outputs(2849));
    layer6_outputs(2851) <= not(layer5_outputs(6350));
    layer6_outputs(2852) <= (layer5_outputs(7086)) and not (layer5_outputs(5430));
    layer6_outputs(2853) <= not(layer5_outputs(2976));
    layer6_outputs(2854) <= (layer5_outputs(3797)) xor (layer5_outputs(4743));
    layer6_outputs(2855) <= layer5_outputs(848);
    layer6_outputs(2856) <= '0';
    layer6_outputs(2857) <= layer5_outputs(2176);
    layer6_outputs(2858) <= not(layer5_outputs(2492));
    layer6_outputs(2859) <= not(layer5_outputs(6565));
    layer6_outputs(2860) <= layer5_outputs(5227);
    layer6_outputs(2861) <= not(layer5_outputs(7130));
    layer6_outputs(2862) <= not(layer5_outputs(6561));
    layer6_outputs(2863) <= layer5_outputs(4277);
    layer6_outputs(2864) <= (layer5_outputs(2440)) xor (layer5_outputs(3705));
    layer6_outputs(2865) <= layer5_outputs(6621);
    layer6_outputs(2866) <= not((layer5_outputs(5254)) or (layer5_outputs(56)));
    layer6_outputs(2867) <= not(layer5_outputs(217));
    layer6_outputs(2868) <= layer5_outputs(597);
    layer6_outputs(2869) <= not(layer5_outputs(6880));
    layer6_outputs(2870) <= layer5_outputs(193);
    layer6_outputs(2871) <= not(layer5_outputs(6337));
    layer6_outputs(2872) <= layer5_outputs(6169);
    layer6_outputs(2873) <= (layer5_outputs(7563)) and not (layer5_outputs(1875));
    layer6_outputs(2874) <= not((layer5_outputs(6208)) xor (layer5_outputs(5592)));
    layer6_outputs(2875) <= not(layer5_outputs(142));
    layer6_outputs(2876) <= '1';
    layer6_outputs(2877) <= not(layer5_outputs(3982));
    layer6_outputs(2878) <= '1';
    layer6_outputs(2879) <= (layer5_outputs(1166)) xor (layer5_outputs(911));
    layer6_outputs(2880) <= (layer5_outputs(2198)) and not (layer5_outputs(1932));
    layer6_outputs(2881) <= layer5_outputs(1864);
    layer6_outputs(2882) <= layer5_outputs(4497);
    layer6_outputs(2883) <= (layer5_outputs(6564)) or (layer5_outputs(4854));
    layer6_outputs(2884) <= layer5_outputs(2398);
    layer6_outputs(2885) <= not(layer5_outputs(7142));
    layer6_outputs(2886) <= not(layer5_outputs(2754)) or (layer5_outputs(6013));
    layer6_outputs(2887) <= not(layer5_outputs(5208));
    layer6_outputs(2888) <= layer5_outputs(3419);
    layer6_outputs(2889) <= not(layer5_outputs(6610));
    layer6_outputs(2890) <= not((layer5_outputs(7005)) xor (layer5_outputs(2026)));
    layer6_outputs(2891) <= not(layer5_outputs(2055));
    layer6_outputs(2892) <= not(layer5_outputs(3438));
    layer6_outputs(2893) <= layer5_outputs(9);
    layer6_outputs(2894) <= not(layer5_outputs(1540));
    layer6_outputs(2895) <= not((layer5_outputs(6739)) and (layer5_outputs(6296)));
    layer6_outputs(2896) <= not(layer5_outputs(1254)) or (layer5_outputs(4172));
    layer6_outputs(2897) <= (layer5_outputs(6269)) and not (layer5_outputs(6888));
    layer6_outputs(2898) <= layer5_outputs(6793);
    layer6_outputs(2899) <= (layer5_outputs(1419)) and (layer5_outputs(1918));
    layer6_outputs(2900) <= not(layer5_outputs(3446));
    layer6_outputs(2901) <= not(layer5_outputs(2479));
    layer6_outputs(2902) <= (layer5_outputs(3425)) and not (layer5_outputs(2506));
    layer6_outputs(2903) <= not(layer5_outputs(5450));
    layer6_outputs(2904) <= layer5_outputs(7405);
    layer6_outputs(2905) <= not(layer5_outputs(3275)) or (layer5_outputs(1699));
    layer6_outputs(2906) <= (layer5_outputs(2877)) xor (layer5_outputs(2223));
    layer6_outputs(2907) <= layer5_outputs(4623);
    layer6_outputs(2908) <= layer5_outputs(2171);
    layer6_outputs(2909) <= not(layer5_outputs(6373));
    layer6_outputs(2910) <= not(layer5_outputs(178));
    layer6_outputs(2911) <= (layer5_outputs(4911)) and not (layer5_outputs(491));
    layer6_outputs(2912) <= layer5_outputs(1782);
    layer6_outputs(2913) <= layer5_outputs(1033);
    layer6_outputs(2914) <= layer5_outputs(4998);
    layer6_outputs(2915) <= not(layer5_outputs(5735));
    layer6_outputs(2916) <= not((layer5_outputs(6765)) or (layer5_outputs(5824)));
    layer6_outputs(2917) <= layer5_outputs(7309);
    layer6_outputs(2918) <= not(layer5_outputs(4895));
    layer6_outputs(2919) <= '0';
    layer6_outputs(2920) <= layer5_outputs(683);
    layer6_outputs(2921) <= '0';
    layer6_outputs(2922) <= layer5_outputs(6277);
    layer6_outputs(2923) <= not(layer5_outputs(7119));
    layer6_outputs(2924) <= layer5_outputs(3736);
    layer6_outputs(2925) <= (layer5_outputs(2027)) and (layer5_outputs(509));
    layer6_outputs(2926) <= not(layer5_outputs(6948));
    layer6_outputs(2927) <= layer5_outputs(4304);
    layer6_outputs(2928) <= (layer5_outputs(4354)) xor (layer5_outputs(4746));
    layer6_outputs(2929) <= (layer5_outputs(3936)) xor (layer5_outputs(4084));
    layer6_outputs(2930) <= not(layer5_outputs(288));
    layer6_outputs(2931) <= (layer5_outputs(3236)) or (layer5_outputs(241));
    layer6_outputs(2932) <= not(layer5_outputs(3901)) or (layer5_outputs(5957));
    layer6_outputs(2933) <= not(layer5_outputs(4436));
    layer6_outputs(2934) <= layer5_outputs(2957);
    layer6_outputs(2935) <= not(layer5_outputs(7511));
    layer6_outputs(2936) <= layer5_outputs(4730);
    layer6_outputs(2937) <= (layer5_outputs(7615)) xor (layer5_outputs(2665));
    layer6_outputs(2938) <= (layer5_outputs(7245)) xor (layer5_outputs(6232));
    layer6_outputs(2939) <= '0';
    layer6_outputs(2940) <= not(layer5_outputs(4198));
    layer6_outputs(2941) <= not(layer5_outputs(77)) or (layer5_outputs(6865));
    layer6_outputs(2942) <= layer5_outputs(752);
    layer6_outputs(2943) <= (layer5_outputs(6696)) and not (layer5_outputs(6653));
    layer6_outputs(2944) <= not(layer5_outputs(1246));
    layer6_outputs(2945) <= (layer5_outputs(3644)) xor (layer5_outputs(1049));
    layer6_outputs(2946) <= not(layer5_outputs(2367));
    layer6_outputs(2947) <= layer5_outputs(7118);
    layer6_outputs(2948) <= not(layer5_outputs(1284));
    layer6_outputs(2949) <= (layer5_outputs(3631)) xor (layer5_outputs(6609));
    layer6_outputs(2950) <= not(layer5_outputs(47));
    layer6_outputs(2951) <= (layer5_outputs(5122)) and not (layer5_outputs(494));
    layer6_outputs(2952) <= layer5_outputs(4576);
    layer6_outputs(2953) <= not(layer5_outputs(1921));
    layer6_outputs(2954) <= not(layer5_outputs(4017)) or (layer5_outputs(321));
    layer6_outputs(2955) <= layer5_outputs(3924);
    layer6_outputs(2956) <= layer5_outputs(3677);
    layer6_outputs(2957) <= not(layer5_outputs(415));
    layer6_outputs(2958) <= (layer5_outputs(6310)) and (layer5_outputs(6024));
    layer6_outputs(2959) <= (layer5_outputs(2128)) and not (layer5_outputs(6505));
    layer6_outputs(2960) <= not(layer5_outputs(2779)) or (layer5_outputs(7363));
    layer6_outputs(2961) <= (layer5_outputs(2656)) and (layer5_outputs(4094));
    layer6_outputs(2962) <= not(layer5_outputs(857));
    layer6_outputs(2963) <= not(layer5_outputs(1646));
    layer6_outputs(2964) <= not(layer5_outputs(4093));
    layer6_outputs(2965) <= (layer5_outputs(1013)) and not (layer5_outputs(673));
    layer6_outputs(2966) <= not(layer5_outputs(1311)) or (layer5_outputs(4581));
    layer6_outputs(2967) <= not((layer5_outputs(7675)) or (layer5_outputs(6888)));
    layer6_outputs(2968) <= not(layer5_outputs(1519)) or (layer5_outputs(3115));
    layer6_outputs(2969) <= layer5_outputs(1249);
    layer6_outputs(2970) <= not(layer5_outputs(5221));
    layer6_outputs(2971) <= not(layer5_outputs(4039));
    layer6_outputs(2972) <= not(layer5_outputs(5089));
    layer6_outputs(2973) <= layer5_outputs(213);
    layer6_outputs(2974) <= not(layer5_outputs(3968));
    layer6_outputs(2975) <= layer5_outputs(4550);
    layer6_outputs(2976) <= (layer5_outputs(4710)) and not (layer5_outputs(6963));
    layer6_outputs(2977) <= not((layer5_outputs(6224)) xor (layer5_outputs(3261)));
    layer6_outputs(2978) <= not((layer5_outputs(86)) and (layer5_outputs(5010)));
    layer6_outputs(2979) <= (layer5_outputs(4734)) and (layer5_outputs(6942));
    layer6_outputs(2980) <= not((layer5_outputs(5149)) xor (layer5_outputs(1840)));
    layer6_outputs(2981) <= (layer5_outputs(755)) and not (layer5_outputs(549));
    layer6_outputs(2982) <= (layer5_outputs(7129)) or (layer5_outputs(4150));
    layer6_outputs(2983) <= '0';
    layer6_outputs(2984) <= not((layer5_outputs(5167)) xor (layer5_outputs(2427)));
    layer6_outputs(2985) <= not(layer5_outputs(5748));
    layer6_outputs(2986) <= not((layer5_outputs(4732)) or (layer5_outputs(5328)));
    layer6_outputs(2987) <= layer5_outputs(6430);
    layer6_outputs(2988) <= not((layer5_outputs(2565)) xor (layer5_outputs(3687)));
    layer6_outputs(2989) <= not(layer5_outputs(4606));
    layer6_outputs(2990) <= layer5_outputs(3087);
    layer6_outputs(2991) <= layer5_outputs(2095);
    layer6_outputs(2992) <= not(layer5_outputs(2589));
    layer6_outputs(2993) <= (layer5_outputs(895)) and not (layer5_outputs(3633));
    layer6_outputs(2994) <= not((layer5_outputs(5685)) and (layer5_outputs(2266)));
    layer6_outputs(2995) <= (layer5_outputs(4021)) or (layer5_outputs(7484));
    layer6_outputs(2996) <= not(layer5_outputs(3288));
    layer6_outputs(2997) <= (layer5_outputs(2620)) and not (layer5_outputs(1458));
    layer6_outputs(2998) <= not(layer5_outputs(6293));
    layer6_outputs(2999) <= not(layer5_outputs(3560));
    layer6_outputs(3000) <= layer5_outputs(7276);
    layer6_outputs(3001) <= not(layer5_outputs(3549)) or (layer5_outputs(7365));
    layer6_outputs(3002) <= layer5_outputs(425);
    layer6_outputs(3003) <= layer5_outputs(2896);
    layer6_outputs(3004) <= not(layer5_outputs(511));
    layer6_outputs(3005) <= not(layer5_outputs(2369));
    layer6_outputs(3006) <= not(layer5_outputs(3478)) or (layer5_outputs(7164));
    layer6_outputs(3007) <= not(layer5_outputs(3156));
    layer6_outputs(3008) <= not((layer5_outputs(1529)) and (layer5_outputs(4104)));
    layer6_outputs(3009) <= (layer5_outputs(5062)) and not (layer5_outputs(4044));
    layer6_outputs(3010) <= layer5_outputs(1065);
    layer6_outputs(3011) <= not(layer5_outputs(4278));
    layer6_outputs(3012) <= layer5_outputs(805);
    layer6_outputs(3013) <= not(layer5_outputs(4014));
    layer6_outputs(3014) <= (layer5_outputs(6375)) and not (layer5_outputs(3805));
    layer6_outputs(3015) <= layer5_outputs(314);
    layer6_outputs(3016) <= not(layer5_outputs(6389));
    layer6_outputs(3017) <= (layer5_outputs(4410)) and (layer5_outputs(2988));
    layer6_outputs(3018) <= (layer5_outputs(1349)) or (layer5_outputs(119));
    layer6_outputs(3019) <= layer5_outputs(2905);
    layer6_outputs(3020) <= layer5_outputs(2183);
    layer6_outputs(3021) <= not((layer5_outputs(5065)) xor (layer5_outputs(5302)));
    layer6_outputs(3022) <= not(layer5_outputs(882)) or (layer5_outputs(7396));
    layer6_outputs(3023) <= layer5_outputs(3268);
    layer6_outputs(3024) <= layer5_outputs(3600);
    layer6_outputs(3025) <= not((layer5_outputs(2336)) xor (layer5_outputs(7211)));
    layer6_outputs(3026) <= not(layer5_outputs(5874));
    layer6_outputs(3027) <= not(layer5_outputs(4923));
    layer6_outputs(3028) <= layer5_outputs(7000);
    layer6_outputs(3029) <= not(layer5_outputs(3663)) or (layer5_outputs(2719));
    layer6_outputs(3030) <= not((layer5_outputs(6322)) xor (layer5_outputs(7419)));
    layer6_outputs(3031) <= not((layer5_outputs(5096)) xor (layer5_outputs(3496)));
    layer6_outputs(3032) <= not((layer5_outputs(100)) or (layer5_outputs(7539)));
    layer6_outputs(3033) <= not(layer5_outputs(6149)) or (layer5_outputs(2803));
    layer6_outputs(3034) <= (layer5_outputs(1812)) and (layer5_outputs(1450));
    layer6_outputs(3035) <= layer5_outputs(3171);
    layer6_outputs(3036) <= not(layer5_outputs(1495));
    layer6_outputs(3037) <= layer5_outputs(4966);
    layer6_outputs(3038) <= not((layer5_outputs(7344)) xor (layer5_outputs(1292)));
    layer6_outputs(3039) <= not((layer5_outputs(4653)) xor (layer5_outputs(2285)));
    layer6_outputs(3040) <= (layer5_outputs(2461)) and not (layer5_outputs(929));
    layer6_outputs(3041) <= (layer5_outputs(3193)) and not (layer5_outputs(5851));
    layer6_outputs(3042) <= (layer5_outputs(2379)) and not (layer5_outputs(1935));
    layer6_outputs(3043) <= not(layer5_outputs(1938));
    layer6_outputs(3044) <= not(layer5_outputs(5508)) or (layer5_outputs(211));
    layer6_outputs(3045) <= (layer5_outputs(424)) and not (layer5_outputs(2827));
    layer6_outputs(3046) <= not((layer5_outputs(2154)) xor (layer5_outputs(93)));
    layer6_outputs(3047) <= not(layer5_outputs(5113)) or (layer5_outputs(1055));
    layer6_outputs(3048) <= not(layer5_outputs(6719));
    layer6_outputs(3049) <= layer5_outputs(7437);
    layer6_outputs(3050) <= not(layer5_outputs(823));
    layer6_outputs(3051) <= (layer5_outputs(6386)) xor (layer5_outputs(6442));
    layer6_outputs(3052) <= layer5_outputs(5350);
    layer6_outputs(3053) <= (layer5_outputs(6621)) and (layer5_outputs(427));
    layer6_outputs(3054) <= (layer5_outputs(6117)) and (layer5_outputs(7425));
    layer6_outputs(3055) <= not(layer5_outputs(3410));
    layer6_outputs(3056) <= not(layer5_outputs(4820)) or (layer5_outputs(6999));
    layer6_outputs(3057) <= not((layer5_outputs(4707)) xor (layer5_outputs(6749)));
    layer6_outputs(3058) <= not(layer5_outputs(6882));
    layer6_outputs(3059) <= (layer5_outputs(2832)) and not (layer5_outputs(5714));
    layer6_outputs(3060) <= not(layer5_outputs(572));
    layer6_outputs(3061) <= layer5_outputs(4437);
    layer6_outputs(3062) <= layer5_outputs(7456);
    layer6_outputs(3063) <= layer5_outputs(524);
    layer6_outputs(3064) <= layer5_outputs(2523);
    layer6_outputs(3065) <= layer5_outputs(1352);
    layer6_outputs(3066) <= not(layer5_outputs(1446)) or (layer5_outputs(3266));
    layer6_outputs(3067) <= not(layer5_outputs(1065));
    layer6_outputs(3068) <= layer5_outputs(6473);
    layer6_outputs(3069) <= not((layer5_outputs(1057)) and (layer5_outputs(3713)));
    layer6_outputs(3070) <= (layer5_outputs(6643)) or (layer5_outputs(217));
    layer6_outputs(3071) <= not(layer5_outputs(2606));
    layer6_outputs(3072) <= (layer5_outputs(5993)) or (layer5_outputs(652));
    layer6_outputs(3073) <= layer5_outputs(1899);
    layer6_outputs(3074) <= not((layer5_outputs(3333)) or (layer5_outputs(1236)));
    layer6_outputs(3075) <= not(layer5_outputs(6107));
    layer6_outputs(3076) <= layer5_outputs(1136);
    layer6_outputs(3077) <= not((layer5_outputs(3005)) or (layer5_outputs(6449)));
    layer6_outputs(3078) <= (layer5_outputs(1445)) and not (layer5_outputs(215));
    layer6_outputs(3079) <= not(layer5_outputs(7036)) or (layer5_outputs(3432));
    layer6_outputs(3080) <= (layer5_outputs(7248)) and not (layer5_outputs(17));
    layer6_outputs(3081) <= '1';
    layer6_outputs(3082) <= layer5_outputs(4127);
    layer6_outputs(3083) <= layer5_outputs(2902);
    layer6_outputs(3084) <= layer5_outputs(7219);
    layer6_outputs(3085) <= layer5_outputs(2394);
    layer6_outputs(3086) <= not((layer5_outputs(1913)) or (layer5_outputs(6363)));
    layer6_outputs(3087) <= not((layer5_outputs(7137)) xor (layer5_outputs(3761)));
    layer6_outputs(3088) <= (layer5_outputs(5051)) or (layer5_outputs(2434));
    layer6_outputs(3089) <= layer5_outputs(3843);
    layer6_outputs(3090) <= layer5_outputs(3197);
    layer6_outputs(3091) <= not(layer5_outputs(4635));
    layer6_outputs(3092) <= not(layer5_outputs(3901)) or (layer5_outputs(6194));
    layer6_outputs(3093) <= not(layer5_outputs(5716)) or (layer5_outputs(6679));
    layer6_outputs(3094) <= not((layer5_outputs(4231)) xor (layer5_outputs(2406)));
    layer6_outputs(3095) <= layer5_outputs(2633);
    layer6_outputs(3096) <= layer5_outputs(817);
    layer6_outputs(3097) <= not(layer5_outputs(2943));
    layer6_outputs(3098) <= layer5_outputs(5172);
    layer6_outputs(3099) <= (layer5_outputs(454)) and not (layer5_outputs(6647));
    layer6_outputs(3100) <= not(layer5_outputs(1657));
    layer6_outputs(3101) <= layer5_outputs(6955);
    layer6_outputs(3102) <= not(layer5_outputs(1502));
    layer6_outputs(3103) <= (layer5_outputs(541)) and not (layer5_outputs(5673));
    layer6_outputs(3104) <= (layer5_outputs(3697)) xor (layer5_outputs(1916));
    layer6_outputs(3105) <= not(layer5_outputs(1443)) or (layer5_outputs(2142));
    layer6_outputs(3106) <= not((layer5_outputs(1526)) xor (layer5_outputs(5767)));
    layer6_outputs(3107) <= not((layer5_outputs(520)) and (layer5_outputs(2011)));
    layer6_outputs(3108) <= layer5_outputs(3437);
    layer6_outputs(3109) <= not(layer5_outputs(5007));
    layer6_outputs(3110) <= not(layer5_outputs(5187));
    layer6_outputs(3111) <= layer5_outputs(4971);
    layer6_outputs(3112) <= (layer5_outputs(1267)) and not (layer5_outputs(5199));
    layer6_outputs(3113) <= layer5_outputs(2982);
    layer6_outputs(3114) <= '0';
    layer6_outputs(3115) <= not(layer5_outputs(3639));
    layer6_outputs(3116) <= (layer5_outputs(1378)) and (layer5_outputs(3201));
    layer6_outputs(3117) <= not(layer5_outputs(5413));
    layer6_outputs(3118) <= not(layer5_outputs(5281));
    layer6_outputs(3119) <= layer5_outputs(1880);
    layer6_outputs(3120) <= (layer5_outputs(4484)) xor (layer5_outputs(5862));
    layer6_outputs(3121) <= not(layer5_outputs(754));
    layer6_outputs(3122) <= (layer5_outputs(4203)) xor (layer5_outputs(4886));
    layer6_outputs(3123) <= layer5_outputs(5273);
    layer6_outputs(3124) <= not(layer5_outputs(1092));
    layer6_outputs(3125) <= not((layer5_outputs(5100)) xor (layer5_outputs(1720)));
    layer6_outputs(3126) <= not(layer5_outputs(1838));
    layer6_outputs(3127) <= not((layer5_outputs(5738)) xor (layer5_outputs(4149)));
    layer6_outputs(3128) <= not(layer5_outputs(5513));
    layer6_outputs(3129) <= not(layer5_outputs(5611)) or (layer5_outputs(3295));
    layer6_outputs(3130) <= layer5_outputs(4944);
    layer6_outputs(3131) <= not(layer5_outputs(977)) or (layer5_outputs(6490));
    layer6_outputs(3132) <= layer5_outputs(6079);
    layer6_outputs(3133) <= (layer5_outputs(1971)) or (layer5_outputs(433));
    layer6_outputs(3134) <= layer5_outputs(2839);
    layer6_outputs(3135) <= (layer5_outputs(5708)) and not (layer5_outputs(1134));
    layer6_outputs(3136) <= not(layer5_outputs(2762));
    layer6_outputs(3137) <= (layer5_outputs(2614)) or (layer5_outputs(6490));
    layer6_outputs(3138) <= not(layer5_outputs(852));
    layer6_outputs(3139) <= (layer5_outputs(526)) or (layer5_outputs(4238));
    layer6_outputs(3140) <= (layer5_outputs(6118)) and (layer5_outputs(974));
    layer6_outputs(3141) <= layer5_outputs(3676);
    layer6_outputs(3142) <= layer5_outputs(973);
    layer6_outputs(3143) <= not(layer5_outputs(4245));
    layer6_outputs(3144) <= not(layer5_outputs(6102));
    layer6_outputs(3145) <= not(layer5_outputs(6862)) or (layer5_outputs(3041));
    layer6_outputs(3146) <= not((layer5_outputs(4257)) xor (layer5_outputs(4040)));
    layer6_outputs(3147) <= not(layer5_outputs(5678));
    layer6_outputs(3148) <= (layer5_outputs(4122)) and not (layer5_outputs(1859));
    layer6_outputs(3149) <= not((layer5_outputs(5279)) or (layer5_outputs(1449)));
    layer6_outputs(3150) <= layer5_outputs(6051);
    layer6_outputs(3151) <= not(layer5_outputs(574));
    layer6_outputs(3152) <= (layer5_outputs(5180)) xor (layer5_outputs(4910));
    layer6_outputs(3153) <= not(layer5_outputs(450));
    layer6_outputs(3154) <= not(layer5_outputs(2364));
    layer6_outputs(3155) <= (layer5_outputs(6673)) xor (layer5_outputs(7552));
    layer6_outputs(3156) <= not((layer5_outputs(2990)) xor (layer5_outputs(5524)));
    layer6_outputs(3157) <= not((layer5_outputs(375)) xor (layer5_outputs(5285)));
    layer6_outputs(3158) <= '0';
    layer6_outputs(3159) <= layer5_outputs(6907);
    layer6_outputs(3160) <= (layer5_outputs(5017)) and not (layer5_outputs(5817));
    layer6_outputs(3161) <= not(layer5_outputs(7312));
    layer6_outputs(3162) <= not(layer5_outputs(6326));
    layer6_outputs(3163) <= not(layer5_outputs(6715));
    layer6_outputs(3164) <= layer5_outputs(7079);
    layer6_outputs(3165) <= (layer5_outputs(3364)) xor (layer5_outputs(4244));
    layer6_outputs(3166) <= not((layer5_outputs(2897)) and (layer5_outputs(4418)));
    layer6_outputs(3167) <= (layer5_outputs(6217)) xor (layer5_outputs(823));
    layer6_outputs(3168) <= not(layer5_outputs(1408));
    layer6_outputs(3169) <= not(layer5_outputs(6623)) or (layer5_outputs(6147));
    layer6_outputs(3170) <= not(layer5_outputs(44));
    layer6_outputs(3171) <= (layer5_outputs(3989)) or (layer5_outputs(5792));
    layer6_outputs(3172) <= layer5_outputs(2204);
    layer6_outputs(3173) <= layer5_outputs(3031);
    layer6_outputs(3174) <= layer5_outputs(3316);
    layer6_outputs(3175) <= '0';
    layer6_outputs(3176) <= (layer5_outputs(123)) and not (layer5_outputs(2042));
    layer6_outputs(3177) <= not(layer5_outputs(1809));
    layer6_outputs(3178) <= layer5_outputs(1021);
    layer6_outputs(3179) <= not(layer5_outputs(1245)) or (layer5_outputs(4639));
    layer6_outputs(3180) <= layer5_outputs(6474);
    layer6_outputs(3181) <= layer5_outputs(2017);
    layer6_outputs(3182) <= layer5_outputs(2354);
    layer6_outputs(3183) <= layer5_outputs(788);
    layer6_outputs(3184) <= not(layer5_outputs(3973));
    layer6_outputs(3185) <= '1';
    layer6_outputs(3186) <= layer5_outputs(2089);
    layer6_outputs(3187) <= not(layer5_outputs(6994));
    layer6_outputs(3188) <= layer5_outputs(188);
    layer6_outputs(3189) <= not(layer5_outputs(1656));
    layer6_outputs(3190) <= not((layer5_outputs(438)) xor (layer5_outputs(1527)));
    layer6_outputs(3191) <= layer5_outputs(2429);
    layer6_outputs(3192) <= layer5_outputs(2377);
    layer6_outputs(3193) <= (layer5_outputs(2309)) or (layer5_outputs(5176));
    layer6_outputs(3194) <= not((layer5_outputs(4097)) and (layer5_outputs(7088)));
    layer6_outputs(3195) <= not(layer5_outputs(424));
    layer6_outputs(3196) <= not(layer5_outputs(4070)) or (layer5_outputs(5724));
    layer6_outputs(3197) <= not(layer5_outputs(6572)) or (layer5_outputs(2409));
    layer6_outputs(3198) <= layer5_outputs(4679);
    layer6_outputs(3199) <= layer5_outputs(3219);
    layer6_outputs(3200) <= layer5_outputs(5402);
    layer6_outputs(3201) <= layer5_outputs(7087);
    layer6_outputs(3202) <= not(layer5_outputs(6487));
    layer6_outputs(3203) <= layer5_outputs(3220);
    layer6_outputs(3204) <= not((layer5_outputs(1523)) or (layer5_outputs(3038)));
    layer6_outputs(3205) <= not(layer5_outputs(1743));
    layer6_outputs(3206) <= not(layer5_outputs(7673));
    layer6_outputs(3207) <= layer5_outputs(5224);
    layer6_outputs(3208) <= layer5_outputs(2333);
    layer6_outputs(3209) <= (layer5_outputs(5379)) or (layer5_outputs(4363));
    layer6_outputs(3210) <= (layer5_outputs(2816)) and not (layer5_outputs(6253));
    layer6_outputs(3211) <= layer5_outputs(1587);
    layer6_outputs(3212) <= (layer5_outputs(2135)) xor (layer5_outputs(2258));
    layer6_outputs(3213) <= not(layer5_outputs(3409)) or (layer5_outputs(7476));
    layer6_outputs(3214) <= (layer5_outputs(6216)) xor (layer5_outputs(284));
    layer6_outputs(3215) <= not(layer5_outputs(3116)) or (layer5_outputs(5282));
    layer6_outputs(3216) <= not((layer5_outputs(2119)) or (layer5_outputs(3646)));
    layer6_outputs(3217) <= not((layer5_outputs(2963)) xor (layer5_outputs(965)));
    layer6_outputs(3218) <= (layer5_outputs(6020)) and not (layer5_outputs(7490));
    layer6_outputs(3219) <= not((layer5_outputs(5125)) xor (layer5_outputs(4952)));
    layer6_outputs(3220) <= not((layer5_outputs(7298)) or (layer5_outputs(3728)));
    layer6_outputs(3221) <= '0';
    layer6_outputs(3222) <= layer5_outputs(6746);
    layer6_outputs(3223) <= not((layer5_outputs(5501)) or (layer5_outputs(3332)));
    layer6_outputs(3224) <= not(layer5_outputs(6876)) or (layer5_outputs(2978));
    layer6_outputs(3225) <= (layer5_outputs(7506)) and not (layer5_outputs(3723));
    layer6_outputs(3226) <= not(layer5_outputs(3060));
    layer6_outputs(3227) <= not(layer5_outputs(44));
    layer6_outputs(3228) <= not(layer5_outputs(1259));
    layer6_outputs(3229) <= (layer5_outputs(1132)) and (layer5_outputs(3394));
    layer6_outputs(3230) <= (layer5_outputs(3783)) and not (layer5_outputs(6556));
    layer6_outputs(3231) <= not((layer5_outputs(7633)) or (layer5_outputs(2759)));
    layer6_outputs(3232) <= layer5_outputs(3211);
    layer6_outputs(3233) <= layer5_outputs(3611);
    layer6_outputs(3234) <= not(layer5_outputs(345));
    layer6_outputs(3235) <= not((layer5_outputs(3951)) xor (layer5_outputs(280)));
    layer6_outputs(3236) <= layer5_outputs(6472);
    layer6_outputs(3237) <= (layer5_outputs(7510)) and not (layer5_outputs(1885));
    layer6_outputs(3238) <= not((layer5_outputs(595)) or (layer5_outputs(4176)));
    layer6_outputs(3239) <= not(layer5_outputs(1894)) or (layer5_outputs(7224));
    layer6_outputs(3240) <= (layer5_outputs(4049)) and not (layer5_outputs(3115));
    layer6_outputs(3241) <= (layer5_outputs(4140)) and not (layer5_outputs(2710));
    layer6_outputs(3242) <= not(layer5_outputs(3651));
    layer6_outputs(3243) <= (layer5_outputs(7396)) and not (layer5_outputs(6885));
    layer6_outputs(3244) <= '1';
    layer6_outputs(3245) <= not(layer5_outputs(3044));
    layer6_outputs(3246) <= not(layer5_outputs(2770));
    layer6_outputs(3247) <= layer5_outputs(1126);
    layer6_outputs(3248) <= (layer5_outputs(2276)) and (layer5_outputs(6125));
    layer6_outputs(3249) <= not(layer5_outputs(4190));
    layer6_outputs(3250) <= not((layer5_outputs(1262)) xor (layer5_outputs(3918)));
    layer6_outputs(3251) <= layer5_outputs(6625);
    layer6_outputs(3252) <= (layer5_outputs(938)) and (layer5_outputs(3979));
    layer6_outputs(3253) <= not(layer5_outputs(2072));
    layer6_outputs(3254) <= layer5_outputs(328);
    layer6_outputs(3255) <= not(layer5_outputs(2761));
    layer6_outputs(3256) <= not(layer5_outputs(2739));
    layer6_outputs(3257) <= not(layer5_outputs(5650));
    layer6_outputs(3258) <= not(layer5_outputs(4608));
    layer6_outputs(3259) <= not(layer5_outputs(5324)) or (layer5_outputs(7237));
    layer6_outputs(3260) <= not((layer5_outputs(1322)) xor (layer5_outputs(3177)));
    layer6_outputs(3261) <= (layer5_outputs(4744)) and not (layer5_outputs(88));
    layer6_outputs(3262) <= layer5_outputs(5913);
    layer6_outputs(3263) <= (layer5_outputs(5878)) and not (layer5_outputs(6015));
    layer6_outputs(3264) <= not((layer5_outputs(5646)) and (layer5_outputs(3627)));
    layer6_outputs(3265) <= not(layer5_outputs(2285));
    layer6_outputs(3266) <= (layer5_outputs(5255)) or (layer5_outputs(1259));
    layer6_outputs(3267) <= not(layer5_outputs(1338));
    layer6_outputs(3268) <= not(layer5_outputs(2674));
    layer6_outputs(3269) <= not((layer5_outputs(373)) or (layer5_outputs(4827)));
    layer6_outputs(3270) <= not(layer5_outputs(4825));
    layer6_outputs(3271) <= layer5_outputs(4046);
    layer6_outputs(3272) <= layer5_outputs(2520);
    layer6_outputs(3273) <= layer5_outputs(5031);
    layer6_outputs(3274) <= not((layer5_outputs(5311)) or (layer5_outputs(2170)));
    layer6_outputs(3275) <= not((layer5_outputs(4053)) xor (layer5_outputs(5532)));
    layer6_outputs(3276) <= (layer5_outputs(6547)) xor (layer5_outputs(6267));
    layer6_outputs(3277) <= (layer5_outputs(2182)) and not (layer5_outputs(2484));
    layer6_outputs(3278) <= layer5_outputs(4371);
    layer6_outputs(3279) <= not(layer5_outputs(4029));
    layer6_outputs(3280) <= layer5_outputs(435);
    layer6_outputs(3281) <= not(layer5_outputs(7568)) or (layer5_outputs(2414));
    layer6_outputs(3282) <= layer5_outputs(4482);
    layer6_outputs(3283) <= not(layer5_outputs(5049));
    layer6_outputs(3284) <= not(layer5_outputs(2405));
    layer6_outputs(3285) <= not(layer5_outputs(4372));
    layer6_outputs(3286) <= not(layer5_outputs(342));
    layer6_outputs(3287) <= layer5_outputs(2037);
    layer6_outputs(3288) <= layer5_outputs(3129);
    layer6_outputs(3289) <= (layer5_outputs(5254)) and not (layer5_outputs(6818));
    layer6_outputs(3290) <= not((layer5_outputs(4275)) xor (layer5_outputs(4161)));
    layer6_outputs(3291) <= (layer5_outputs(7519)) xor (layer5_outputs(1005));
    layer6_outputs(3292) <= not(layer5_outputs(2568));
    layer6_outputs(3293) <= not((layer5_outputs(2052)) xor (layer5_outputs(1952)));
    layer6_outputs(3294) <= not(layer5_outputs(2091)) or (layer5_outputs(5546));
    layer6_outputs(3295) <= (layer5_outputs(1750)) and not (layer5_outputs(3202));
    layer6_outputs(3296) <= layer5_outputs(3370);
    layer6_outputs(3297) <= not((layer5_outputs(2610)) or (layer5_outputs(1457)));
    layer6_outputs(3298) <= not(layer5_outputs(2106));
    layer6_outputs(3299) <= (layer5_outputs(418)) and not (layer5_outputs(6503));
    layer6_outputs(3300) <= layer5_outputs(6708);
    layer6_outputs(3301) <= not(layer5_outputs(6886));
    layer6_outputs(3302) <= not(layer5_outputs(241)) or (layer5_outputs(1004));
    layer6_outputs(3303) <= not(layer5_outputs(240));
    layer6_outputs(3304) <= not(layer5_outputs(4797)) or (layer5_outputs(4904));
    layer6_outputs(3305) <= '0';
    layer6_outputs(3306) <= not(layer5_outputs(4345));
    layer6_outputs(3307) <= not(layer5_outputs(5954));
    layer6_outputs(3308) <= not(layer5_outputs(1985));
    layer6_outputs(3309) <= (layer5_outputs(1961)) and not (layer5_outputs(4336));
    layer6_outputs(3310) <= (layer5_outputs(3555)) xor (layer5_outputs(5238));
    layer6_outputs(3311) <= not(layer5_outputs(58)) or (layer5_outputs(5814));
    layer6_outputs(3312) <= layer5_outputs(1521);
    layer6_outputs(3313) <= not((layer5_outputs(2901)) xor (layer5_outputs(1531)));
    layer6_outputs(3314) <= (layer5_outputs(194)) and not (layer5_outputs(5973));
    layer6_outputs(3315) <= layer5_outputs(7678);
    layer6_outputs(3316) <= layer5_outputs(5361);
    layer6_outputs(3317) <= not(layer5_outputs(3316));
    layer6_outputs(3318) <= layer5_outputs(1785);
    layer6_outputs(3319) <= (layer5_outputs(4176)) xor (layer5_outputs(1277));
    layer6_outputs(3320) <= layer5_outputs(7300);
    layer6_outputs(3321) <= layer5_outputs(4678);
    layer6_outputs(3322) <= (layer5_outputs(6537)) xor (layer5_outputs(658));
    layer6_outputs(3323) <= layer5_outputs(5643);
    layer6_outputs(3324) <= (layer5_outputs(1599)) xor (layer5_outputs(3175));
    layer6_outputs(3325) <= layer5_outputs(6512);
    layer6_outputs(3326) <= layer5_outputs(3498);
    layer6_outputs(3327) <= layer5_outputs(6835);
    layer6_outputs(3328) <= not((layer5_outputs(3330)) xor (layer5_outputs(5130)));
    layer6_outputs(3329) <= layer5_outputs(4995);
    layer6_outputs(3330) <= layer5_outputs(4138);
    layer6_outputs(3331) <= (layer5_outputs(2196)) xor (layer5_outputs(6413));
    layer6_outputs(3332) <= not((layer5_outputs(2426)) or (layer5_outputs(437)));
    layer6_outputs(3333) <= not((layer5_outputs(3249)) xor (layer5_outputs(702)));
    layer6_outputs(3334) <= not(layer5_outputs(2065));
    layer6_outputs(3335) <= not(layer5_outputs(4458));
    layer6_outputs(3336) <= not((layer5_outputs(4331)) or (layer5_outputs(1603)));
    layer6_outputs(3337) <= not(layer5_outputs(2700));
    layer6_outputs(3338) <= not(layer5_outputs(3167)) or (layer5_outputs(4765));
    layer6_outputs(3339) <= (layer5_outputs(1425)) and not (layer5_outputs(7344));
    layer6_outputs(3340) <= not(layer5_outputs(1748));
    layer6_outputs(3341) <= not(layer5_outputs(1200));
    layer6_outputs(3342) <= not(layer5_outputs(4950));
    layer6_outputs(3343) <= (layer5_outputs(7457)) and (layer5_outputs(4148));
    layer6_outputs(3344) <= not((layer5_outputs(6692)) xor (layer5_outputs(7634)));
    layer6_outputs(3345) <= layer5_outputs(4383);
    layer6_outputs(3346) <= not((layer5_outputs(6085)) xor (layer5_outputs(659)));
    layer6_outputs(3347) <= not(layer5_outputs(182));
    layer6_outputs(3348) <= layer5_outputs(1673);
    layer6_outputs(3349) <= not(layer5_outputs(2048)) or (layer5_outputs(3525));
    layer6_outputs(3350) <= (layer5_outputs(2893)) and not (layer5_outputs(5842));
    layer6_outputs(3351) <= layer5_outputs(4775);
    layer6_outputs(3352) <= layer5_outputs(6034);
    layer6_outputs(3353) <= not(layer5_outputs(6670)) or (layer5_outputs(6506));
    layer6_outputs(3354) <= not(layer5_outputs(7218));
    layer6_outputs(3355) <= layer5_outputs(2203);
    layer6_outputs(3356) <= not(layer5_outputs(1957));
    layer6_outputs(3357) <= (layer5_outputs(5205)) xor (layer5_outputs(491));
    layer6_outputs(3358) <= (layer5_outputs(5584)) xor (layer5_outputs(7477));
    layer6_outputs(3359) <= not(layer5_outputs(1777));
    layer6_outputs(3360) <= layer5_outputs(360);
    layer6_outputs(3361) <= not((layer5_outputs(3152)) xor (layer5_outputs(4762)));
    layer6_outputs(3362) <= (layer5_outputs(2499)) xor (layer5_outputs(1219));
    layer6_outputs(3363) <= (layer5_outputs(7507)) xor (layer5_outputs(2799));
    layer6_outputs(3364) <= layer5_outputs(3533);
    layer6_outputs(3365) <= not(layer5_outputs(7386));
    layer6_outputs(3366) <= not(layer5_outputs(4794));
    layer6_outputs(3367) <= layer5_outputs(757);
    layer6_outputs(3368) <= not((layer5_outputs(2772)) or (layer5_outputs(283)));
    layer6_outputs(3369) <= (layer5_outputs(6478)) or (layer5_outputs(189));
    layer6_outputs(3370) <= not(layer5_outputs(6822));
    layer6_outputs(3371) <= not(layer5_outputs(1748)) or (layer5_outputs(4961));
    layer6_outputs(3372) <= (layer5_outputs(2314)) xor (layer5_outputs(4964));
    layer6_outputs(3373) <= layer5_outputs(4751);
    layer6_outputs(3374) <= not((layer5_outputs(2421)) and (layer5_outputs(2773)));
    layer6_outputs(3375) <= not((layer5_outputs(1284)) xor (layer5_outputs(3329)));
    layer6_outputs(3376) <= not(layer5_outputs(5354));
    layer6_outputs(3377) <= (layer5_outputs(3758)) xor (layer5_outputs(2869));
    layer6_outputs(3378) <= not((layer5_outputs(2359)) xor (layer5_outputs(5442)));
    layer6_outputs(3379) <= not(layer5_outputs(1884));
    layer6_outputs(3380) <= layer5_outputs(2351);
    layer6_outputs(3381) <= layer5_outputs(5179);
    layer6_outputs(3382) <= not(layer5_outputs(2272));
    layer6_outputs(3383) <= not(layer5_outputs(5182)) or (layer5_outputs(6192));
    layer6_outputs(3384) <= (layer5_outputs(402)) xor (layer5_outputs(7399));
    layer6_outputs(3385) <= layer5_outputs(5677);
    layer6_outputs(3386) <= not(layer5_outputs(6383));
    layer6_outputs(3387) <= not(layer5_outputs(7629));
    layer6_outputs(3388) <= layer5_outputs(2430);
    layer6_outputs(3389) <= layer5_outputs(4742);
    layer6_outputs(3390) <= (layer5_outputs(3893)) xor (layer5_outputs(3686));
    layer6_outputs(3391) <= layer5_outputs(6445);
    layer6_outputs(3392) <= not(layer5_outputs(2184)) or (layer5_outputs(5243));
    layer6_outputs(3393) <= (layer5_outputs(4499)) and not (layer5_outputs(2527));
    layer6_outputs(3394) <= not(layer5_outputs(1469));
    layer6_outputs(3395) <= (layer5_outputs(4148)) and not (layer5_outputs(1701));
    layer6_outputs(3396) <= not(layer5_outputs(3088));
    layer6_outputs(3397) <= layer5_outputs(4065);
    layer6_outputs(3398) <= not(layer5_outputs(2884));
    layer6_outputs(3399) <= not((layer5_outputs(6356)) and (layer5_outputs(3671)));
    layer6_outputs(3400) <= (layer5_outputs(1516)) and not (layer5_outputs(5148));
    layer6_outputs(3401) <= layer5_outputs(5704);
    layer6_outputs(3402) <= layer5_outputs(7580);
    layer6_outputs(3403) <= (layer5_outputs(6502)) and not (layer5_outputs(6177));
    layer6_outputs(3404) <= not((layer5_outputs(4311)) xor (layer5_outputs(6162)));
    layer6_outputs(3405) <= layer5_outputs(276);
    layer6_outputs(3406) <= not(layer5_outputs(4394)) or (layer5_outputs(4177));
    layer6_outputs(3407) <= not(layer5_outputs(3450));
    layer6_outputs(3408) <= layer5_outputs(498);
    layer6_outputs(3409) <= layer5_outputs(627);
    layer6_outputs(3410) <= (layer5_outputs(2764)) and not (layer5_outputs(3420));
    layer6_outputs(3411) <= not(layer5_outputs(5160));
    layer6_outputs(3412) <= not(layer5_outputs(2055)) or (layer5_outputs(1692));
    layer6_outputs(3413) <= not(layer5_outputs(5465));
    layer6_outputs(3414) <= layer5_outputs(6667);
    layer6_outputs(3415) <= layer5_outputs(2587);
    layer6_outputs(3416) <= (layer5_outputs(3023)) xor (layer5_outputs(6966));
    layer6_outputs(3417) <= layer5_outputs(7509);
    layer6_outputs(3418) <= layer5_outputs(4384);
    layer6_outputs(3419) <= layer5_outputs(2542);
    layer6_outputs(3420) <= (layer5_outputs(3287)) xor (layer5_outputs(1640));
    layer6_outputs(3421) <= not(layer5_outputs(2162));
    layer6_outputs(3422) <= layer5_outputs(5434);
    layer6_outputs(3423) <= layer5_outputs(1406);
    layer6_outputs(3424) <= layer5_outputs(4788);
    layer6_outputs(3425) <= layer5_outputs(3947);
    layer6_outputs(3426) <= (layer5_outputs(501)) xor (layer5_outputs(3155));
    layer6_outputs(3427) <= (layer5_outputs(1770)) and not (layer5_outputs(2734));
    layer6_outputs(3428) <= not(layer5_outputs(5653));
    layer6_outputs(3429) <= layer5_outputs(7401);
    layer6_outputs(3430) <= not(layer5_outputs(7372));
    layer6_outputs(3431) <= not((layer5_outputs(4825)) and (layer5_outputs(5336)));
    layer6_outputs(3432) <= (layer5_outputs(997)) xor (layer5_outputs(2802));
    layer6_outputs(3433) <= not(layer5_outputs(3105));
    layer6_outputs(3434) <= not((layer5_outputs(4738)) xor (layer5_outputs(1428)));
    layer6_outputs(3435) <= not(layer5_outputs(2504));
    layer6_outputs(3436) <= not(layer5_outputs(2857)) or (layer5_outputs(200));
    layer6_outputs(3437) <= not(layer5_outputs(2077));
    layer6_outputs(3438) <= (layer5_outputs(7165)) and not (layer5_outputs(4622));
    layer6_outputs(3439) <= not(layer5_outputs(7604)) or (layer5_outputs(1328));
    layer6_outputs(3440) <= not(layer5_outputs(4200)) or (layer5_outputs(5835));
    layer6_outputs(3441) <= not((layer5_outputs(5719)) xor (layer5_outputs(269)));
    layer6_outputs(3442) <= not(layer5_outputs(2550));
    layer6_outputs(3443) <= layer5_outputs(4400);
    layer6_outputs(3444) <= not(layer5_outputs(1163));
    layer6_outputs(3445) <= layer5_outputs(1154);
    layer6_outputs(3446) <= not(layer5_outputs(1958));
    layer6_outputs(3447) <= not(layer5_outputs(3279));
    layer6_outputs(3448) <= (layer5_outputs(4576)) xor (layer5_outputs(4367));
    layer6_outputs(3449) <= not((layer5_outputs(5918)) xor (layer5_outputs(2041)));
    layer6_outputs(3450) <= not(layer5_outputs(481));
    layer6_outputs(3451) <= (layer5_outputs(3590)) and (layer5_outputs(4116));
    layer6_outputs(3452) <= not(layer5_outputs(1520)) or (layer5_outputs(196));
    layer6_outputs(3453) <= not((layer5_outputs(3140)) xor (layer5_outputs(7355)));
    layer6_outputs(3454) <= layer5_outputs(5026);
    layer6_outputs(3455) <= not((layer5_outputs(235)) xor (layer5_outputs(1104)));
    layer6_outputs(3456) <= layer5_outputs(2932);
    layer6_outputs(3457) <= (layer5_outputs(509)) and (layer5_outputs(2815));
    layer6_outputs(3458) <= layer5_outputs(604);
    layer6_outputs(3459) <= layer5_outputs(6711);
    layer6_outputs(3460) <= not(layer5_outputs(4728)) or (layer5_outputs(869));
    layer6_outputs(3461) <= not((layer5_outputs(7312)) or (layer5_outputs(2765)));
    layer6_outputs(3462) <= layer5_outputs(5378);
    layer6_outputs(3463) <= not((layer5_outputs(4646)) xor (layer5_outputs(5518)));
    layer6_outputs(3464) <= layer5_outputs(3233);
    layer6_outputs(3465) <= not(layer5_outputs(2679));
    layer6_outputs(3466) <= not(layer5_outputs(4432)) or (layer5_outputs(6798));
    layer6_outputs(3467) <= not(layer5_outputs(6779)) or (layer5_outputs(6285));
    layer6_outputs(3468) <= not(layer5_outputs(6082)) or (layer5_outputs(6589));
    layer6_outputs(3469) <= layer5_outputs(396);
    layer6_outputs(3470) <= (layer5_outputs(2813)) and (layer5_outputs(2598));
    layer6_outputs(3471) <= layer5_outputs(2413);
    layer6_outputs(3472) <= layer5_outputs(471);
    layer6_outputs(3473) <= (layer5_outputs(638)) or (layer5_outputs(167));
    layer6_outputs(3474) <= not((layer5_outputs(4665)) and (layer5_outputs(180)));
    layer6_outputs(3475) <= layer5_outputs(472);
    layer6_outputs(3476) <= (layer5_outputs(6417)) xor (layer5_outputs(686));
    layer6_outputs(3477) <= not((layer5_outputs(6926)) xor (layer5_outputs(5960)));
    layer6_outputs(3478) <= not((layer5_outputs(4852)) or (layer5_outputs(7577)));
    layer6_outputs(3479) <= not(layer5_outputs(3887));
    layer6_outputs(3480) <= not(layer5_outputs(6345));
    layer6_outputs(3481) <= (layer5_outputs(7378)) or (layer5_outputs(2341));
    layer6_outputs(3482) <= (layer5_outputs(1162)) and not (layer5_outputs(5340));
    layer6_outputs(3483) <= (layer5_outputs(1620)) and (layer5_outputs(1020));
    layer6_outputs(3484) <= layer5_outputs(4246);
    layer6_outputs(3485) <= (layer5_outputs(4902)) and (layer5_outputs(4605));
    layer6_outputs(3486) <= (layer5_outputs(3136)) xor (layer5_outputs(5214));
    layer6_outputs(3487) <= not((layer5_outputs(4132)) xor (layer5_outputs(7212)));
    layer6_outputs(3488) <= not(layer5_outputs(6343));
    layer6_outputs(3489) <= not(layer5_outputs(4275));
    layer6_outputs(3490) <= not(layer5_outputs(7544));
    layer6_outputs(3491) <= not((layer5_outputs(4194)) and (layer5_outputs(59)));
    layer6_outputs(3492) <= not(layer5_outputs(3772));
    layer6_outputs(3493) <= not(layer5_outputs(1451));
    layer6_outputs(3494) <= (layer5_outputs(5610)) xor (layer5_outputs(6168));
    layer6_outputs(3495) <= not((layer5_outputs(488)) xor (layer5_outputs(2514)));
    layer6_outputs(3496) <= layer5_outputs(5521);
    layer6_outputs(3497) <= not(layer5_outputs(4598)) or (layer5_outputs(4385));
    layer6_outputs(3498) <= not(layer5_outputs(1438));
    layer6_outputs(3499) <= (layer5_outputs(572)) or (layer5_outputs(1295));
    layer6_outputs(3500) <= not(layer5_outputs(5500));
    layer6_outputs(3501) <= layer5_outputs(3549);
    layer6_outputs(3502) <= (layer5_outputs(5203)) and (layer5_outputs(5641));
    layer6_outputs(3503) <= not(layer5_outputs(7255));
    layer6_outputs(3504) <= not(layer5_outputs(4240));
    layer6_outputs(3505) <= (layer5_outputs(6655)) xor (layer5_outputs(5338));
    layer6_outputs(3506) <= (layer5_outputs(6809)) or (layer5_outputs(2628));
    layer6_outputs(3507) <= layer5_outputs(1315);
    layer6_outputs(3508) <= layer5_outputs(2204);
    layer6_outputs(3509) <= (layer5_outputs(274)) xor (layer5_outputs(5245));
    layer6_outputs(3510) <= not(layer5_outputs(896));
    layer6_outputs(3511) <= not(layer5_outputs(5948));
    layer6_outputs(3512) <= (layer5_outputs(1542)) or (layer5_outputs(6170));
    layer6_outputs(3513) <= not(layer5_outputs(1824));
    layer6_outputs(3514) <= not((layer5_outputs(4490)) and (layer5_outputs(4846)));
    layer6_outputs(3515) <= not((layer5_outputs(4005)) or (layer5_outputs(3959)));
    layer6_outputs(3516) <= (layer5_outputs(5591)) xor (layer5_outputs(2164));
    layer6_outputs(3517) <= not((layer5_outputs(6152)) and (layer5_outputs(7603)));
    layer6_outputs(3518) <= not(layer5_outputs(580));
    layer6_outputs(3519) <= (layer5_outputs(7229)) and not (layer5_outputs(6148));
    layer6_outputs(3520) <= (layer5_outputs(6648)) and not (layer5_outputs(6462));
    layer6_outputs(3521) <= layer5_outputs(4329);
    layer6_outputs(3522) <= (layer5_outputs(6701)) or (layer5_outputs(381));
    layer6_outputs(3523) <= not(layer5_outputs(5925));
    layer6_outputs(3524) <= not(layer5_outputs(1252));
    layer6_outputs(3525) <= not(layer5_outputs(7029));
    layer6_outputs(3526) <= layer5_outputs(2818);
    layer6_outputs(3527) <= not(layer5_outputs(4887));
    layer6_outputs(3528) <= not(layer5_outputs(3877));
    layer6_outputs(3529) <= (layer5_outputs(7339)) or (layer5_outputs(1536));
    layer6_outputs(3530) <= not(layer5_outputs(2275));
    layer6_outputs(3531) <= not(layer5_outputs(6364));
    layer6_outputs(3532) <= layer5_outputs(5568);
    layer6_outputs(3533) <= (layer5_outputs(3439)) and (layer5_outputs(7242));
    layer6_outputs(3534) <= not(layer5_outputs(3986)) or (layer5_outputs(3699));
    layer6_outputs(3535) <= (layer5_outputs(1674)) xor (layer5_outputs(6255));
    layer6_outputs(3536) <= '0';
    layer6_outputs(3537) <= (layer5_outputs(125)) and not (layer5_outputs(1014));
    layer6_outputs(3538) <= layer5_outputs(4837);
    layer6_outputs(3539) <= (layer5_outputs(5915)) xor (layer5_outputs(2449));
    layer6_outputs(3540) <= (layer5_outputs(4368)) xor (layer5_outputs(6308));
    layer6_outputs(3541) <= layer5_outputs(3401);
    layer6_outputs(3542) <= not((layer5_outputs(5799)) and (layer5_outputs(2879)));
    layer6_outputs(3543) <= layer5_outputs(1537);
    layer6_outputs(3544) <= layer5_outputs(3011);
    layer6_outputs(3545) <= not(layer5_outputs(4248));
    layer6_outputs(3546) <= not(layer5_outputs(4664));
    layer6_outputs(3547) <= layer5_outputs(4117);
    layer6_outputs(3548) <= (layer5_outputs(2545)) xor (layer5_outputs(3991));
    layer6_outputs(3549) <= (layer5_outputs(5851)) xor (layer5_outputs(415));
    layer6_outputs(3550) <= not(layer5_outputs(143));
    layer6_outputs(3551) <= (layer5_outputs(5451)) or (layer5_outputs(4022));
    layer6_outputs(3552) <= layer5_outputs(6712);
    layer6_outputs(3553) <= not(layer5_outputs(4239));
    layer6_outputs(3554) <= not(layer5_outputs(5930));
    layer6_outputs(3555) <= layer5_outputs(4551);
    layer6_outputs(3556) <= layer5_outputs(2164);
    layer6_outputs(3557) <= not((layer5_outputs(1398)) or (layer5_outputs(5443)));
    layer6_outputs(3558) <= layer5_outputs(4087);
    layer6_outputs(3559) <= (layer5_outputs(5901)) xor (layer5_outputs(4721));
    layer6_outputs(3560) <= layer5_outputs(6526);
    layer6_outputs(3561) <= (layer5_outputs(6969)) and (layer5_outputs(1228));
    layer6_outputs(3562) <= not(layer5_outputs(2939)) or (layer5_outputs(305));
    layer6_outputs(3563) <= layer5_outputs(6632);
    layer6_outputs(3564) <= layer5_outputs(439);
    layer6_outputs(3565) <= not(layer5_outputs(1097));
    layer6_outputs(3566) <= layer5_outputs(7138);
    layer6_outputs(3567) <= layer5_outputs(1899);
    layer6_outputs(3568) <= layer5_outputs(2094);
    layer6_outputs(3569) <= not(layer5_outputs(2955));
    layer6_outputs(3570) <= not((layer5_outputs(6885)) and (layer5_outputs(3745)));
    layer6_outputs(3571) <= layer5_outputs(3659);
    layer6_outputs(3572) <= not(layer5_outputs(1846));
    layer6_outputs(3573) <= layer5_outputs(4555);
    layer6_outputs(3574) <= (layer5_outputs(4228)) xor (layer5_outputs(3350));
    layer6_outputs(3575) <= (layer5_outputs(5134)) or (layer5_outputs(7052));
    layer6_outputs(3576) <= not(layer5_outputs(1205)) or (layer5_outputs(4238));
    layer6_outputs(3577) <= (layer5_outputs(3508)) or (layer5_outputs(1419));
    layer6_outputs(3578) <= not(layer5_outputs(4232));
    layer6_outputs(3579) <= not(layer5_outputs(4579)) or (layer5_outputs(6832));
    layer6_outputs(3580) <= not(layer5_outputs(5812));
    layer6_outputs(3581) <= not(layer5_outputs(7073));
    layer6_outputs(3582) <= layer5_outputs(4300);
    layer6_outputs(3583) <= not((layer5_outputs(1291)) and (layer5_outputs(1054)));
    layer6_outputs(3584) <= (layer5_outputs(2489)) xor (layer5_outputs(3970));
    layer6_outputs(3585) <= not(layer5_outputs(2325));
    layer6_outputs(3586) <= not(layer5_outputs(7563));
    layer6_outputs(3587) <= (layer5_outputs(7394)) xor (layer5_outputs(4668));
    layer6_outputs(3588) <= not(layer5_outputs(2235));
    layer6_outputs(3589) <= not(layer5_outputs(1305));
    layer6_outputs(3590) <= not((layer5_outputs(506)) xor (layer5_outputs(225)));
    layer6_outputs(3591) <= not((layer5_outputs(3282)) xor (layer5_outputs(2035)));
    layer6_outputs(3592) <= layer5_outputs(1591);
    layer6_outputs(3593) <= (layer5_outputs(5762)) and not (layer5_outputs(3802));
    layer6_outputs(3594) <= not(layer5_outputs(7481));
    layer6_outputs(3595) <= layer5_outputs(2946);
    layer6_outputs(3596) <= not((layer5_outputs(83)) or (layer5_outputs(93)));
    layer6_outputs(3597) <= layer5_outputs(6931);
    layer6_outputs(3598) <= not(layer5_outputs(205));
    layer6_outputs(3599) <= not(layer5_outputs(4501));
    layer6_outputs(3600) <= not((layer5_outputs(4380)) or (layer5_outputs(1482)));
    layer6_outputs(3601) <= not(layer5_outputs(3266));
    layer6_outputs(3602) <= (layer5_outputs(106)) xor (layer5_outputs(2476));
    layer6_outputs(3603) <= (layer5_outputs(2495)) and not (layer5_outputs(3640));
    layer6_outputs(3604) <= not(layer5_outputs(7356)) or (layer5_outputs(1283));
    layer6_outputs(3605) <= not(layer5_outputs(1945));
    layer6_outputs(3606) <= (layer5_outputs(3563)) or (layer5_outputs(4535));
    layer6_outputs(3607) <= (layer5_outputs(7328)) and (layer5_outputs(242));
    layer6_outputs(3608) <= (layer5_outputs(4559)) and not (layer5_outputs(7102));
    layer6_outputs(3609) <= not(layer5_outputs(933));
    layer6_outputs(3610) <= not((layer5_outputs(1352)) xor (layer5_outputs(3193)));
    layer6_outputs(3611) <= not((layer5_outputs(5938)) or (layer5_outputs(2172)));
    layer6_outputs(3612) <= not(layer5_outputs(1718));
    layer6_outputs(3613) <= '0';
    layer6_outputs(3614) <= not(layer5_outputs(3263));
    layer6_outputs(3615) <= not((layer5_outputs(6520)) xor (layer5_outputs(3251)));
    layer6_outputs(3616) <= layer5_outputs(684);
    layer6_outputs(3617) <= (layer5_outputs(7455)) or (layer5_outputs(5128));
    layer6_outputs(3618) <= not(layer5_outputs(1786)) or (layer5_outputs(7654));
    layer6_outputs(3619) <= not(layer5_outputs(5785));
    layer6_outputs(3620) <= not(layer5_outputs(1822));
    layer6_outputs(3621) <= (layer5_outputs(164)) and (layer5_outputs(4157));
    layer6_outputs(3622) <= (layer5_outputs(3656)) and not (layer5_outputs(2572));
    layer6_outputs(3623) <= not(layer5_outputs(4034));
    layer6_outputs(3624) <= not(layer5_outputs(5546));
    layer6_outputs(3625) <= (layer5_outputs(4064)) and not (layer5_outputs(7502));
    layer6_outputs(3626) <= layer5_outputs(1810);
    layer6_outputs(3627) <= layer5_outputs(2034);
    layer6_outputs(3628) <= (layer5_outputs(6295)) and not (layer5_outputs(156));
    layer6_outputs(3629) <= (layer5_outputs(2918)) or (layer5_outputs(3534));
    layer6_outputs(3630) <= not(layer5_outputs(4072));
    layer6_outputs(3631) <= (layer5_outputs(248)) and not (layer5_outputs(6584));
    layer6_outputs(3632) <= not(layer5_outputs(1789));
    layer6_outputs(3633) <= (layer5_outputs(3715)) xor (layer5_outputs(1476));
    layer6_outputs(3634) <= layer5_outputs(5726);
    layer6_outputs(3635) <= (layer5_outputs(819)) xor (layer5_outputs(3767));
    layer6_outputs(3636) <= (layer5_outputs(7417)) xor (layer5_outputs(1604));
    layer6_outputs(3637) <= not((layer5_outputs(5622)) or (layer5_outputs(1569)));
    layer6_outputs(3638) <= not(layer5_outputs(2221));
    layer6_outputs(3639) <= not(layer5_outputs(6866));
    layer6_outputs(3640) <= layer5_outputs(1678);
    layer6_outputs(3641) <= (layer5_outputs(6898)) and not (layer5_outputs(2411));
    layer6_outputs(3642) <= layer5_outputs(6564);
    layer6_outputs(3643) <= not((layer5_outputs(5655)) xor (layer5_outputs(4138)));
    layer6_outputs(3644) <= layer5_outputs(5241);
    layer6_outputs(3645) <= (layer5_outputs(2186)) xor (layer5_outputs(2830));
    layer6_outputs(3646) <= not((layer5_outputs(3864)) and (layer5_outputs(6237)));
    layer6_outputs(3647) <= not((layer5_outputs(7051)) xor (layer5_outputs(4560)));
    layer6_outputs(3648) <= not((layer5_outputs(1514)) and (layer5_outputs(3268)));
    layer6_outputs(3649) <= not(layer5_outputs(634));
    layer6_outputs(3650) <= not(layer5_outputs(899));
    layer6_outputs(3651) <= not(layer5_outputs(6262));
    layer6_outputs(3652) <= not(layer5_outputs(338));
    layer6_outputs(3653) <= (layer5_outputs(4765)) xor (layer5_outputs(1529));
    layer6_outputs(3654) <= not(layer5_outputs(257));
    layer6_outputs(3655) <= not(layer5_outputs(3239)) or (layer5_outputs(578));
    layer6_outputs(3656) <= not(layer5_outputs(1855));
    layer6_outputs(3657) <= not(layer5_outputs(2453));
    layer6_outputs(3658) <= not(layer5_outputs(7123));
    layer6_outputs(3659) <= layer5_outputs(2954);
    layer6_outputs(3660) <= layer5_outputs(15);
    layer6_outputs(3661) <= not((layer5_outputs(2687)) and (layer5_outputs(1845)));
    layer6_outputs(3662) <= (layer5_outputs(324)) xor (layer5_outputs(4059));
    layer6_outputs(3663) <= not(layer5_outputs(6248));
    layer6_outputs(3664) <= layer5_outputs(3921);
    layer6_outputs(3665) <= not(layer5_outputs(5127));
    layer6_outputs(3666) <= not((layer5_outputs(3252)) xor (layer5_outputs(4481)));
    layer6_outputs(3667) <= not(layer5_outputs(1066));
    layer6_outputs(3668) <= not(layer5_outputs(4812));
    layer6_outputs(3669) <= (layer5_outputs(3884)) or (layer5_outputs(4382));
    layer6_outputs(3670) <= layer5_outputs(6360);
    layer6_outputs(3671) <= (layer5_outputs(777)) and not (layer5_outputs(7275));
    layer6_outputs(3672) <= not(layer5_outputs(3781));
    layer6_outputs(3673) <= not(layer5_outputs(7043));
    layer6_outputs(3674) <= not(layer5_outputs(6392));
    layer6_outputs(3675) <= not(layer5_outputs(2689));
    layer6_outputs(3676) <= layer5_outputs(3238);
    layer6_outputs(3677) <= not((layer5_outputs(4540)) and (layer5_outputs(2475)));
    layer6_outputs(3678) <= (layer5_outputs(6997)) and not (layer5_outputs(4208));
    layer6_outputs(3679) <= not(layer5_outputs(2623));
    layer6_outputs(3680) <= not((layer5_outputs(6921)) xor (layer5_outputs(2942)));
    layer6_outputs(3681) <= layer5_outputs(2541);
    layer6_outputs(3682) <= layer5_outputs(43);
    layer6_outputs(3683) <= (layer5_outputs(4621)) and (layer5_outputs(7060));
    layer6_outputs(3684) <= not(layer5_outputs(1053));
    layer6_outputs(3685) <= not(layer5_outputs(1230));
    layer6_outputs(3686) <= not((layer5_outputs(3537)) and (layer5_outputs(5284)));
    layer6_outputs(3687) <= not(layer5_outputs(1543));
    layer6_outputs(3688) <= layer5_outputs(3296);
    layer6_outputs(3689) <= not(layer5_outputs(3414)) or (layer5_outputs(7375));
    layer6_outputs(3690) <= not(layer5_outputs(758));
    layer6_outputs(3691) <= layer5_outputs(1809);
    layer6_outputs(3692) <= not(layer5_outputs(2673));
    layer6_outputs(3693) <= layer5_outputs(181);
    layer6_outputs(3694) <= not((layer5_outputs(7055)) xor (layer5_outputs(2160)));
    layer6_outputs(3695) <= not(layer5_outputs(1768));
    layer6_outputs(3696) <= not((layer5_outputs(2703)) and (layer5_outputs(5174)));
    layer6_outputs(3697) <= layer5_outputs(4580);
    layer6_outputs(3698) <= not(layer5_outputs(4214));
    layer6_outputs(3699) <= not(layer5_outputs(3509));
    layer6_outputs(3700) <= not(layer5_outputs(6092));
    layer6_outputs(3701) <= not((layer5_outputs(264)) and (layer5_outputs(2380)));
    layer6_outputs(3702) <= '1';
    layer6_outputs(3703) <= not((layer5_outputs(6572)) xor (layer5_outputs(1927)));
    layer6_outputs(3704) <= (layer5_outputs(3474)) or (layer5_outputs(1024));
    layer6_outputs(3705) <= '0';
    layer6_outputs(3706) <= not((layer5_outputs(5181)) xor (layer5_outputs(813)));
    layer6_outputs(3707) <= layer5_outputs(7327);
    layer6_outputs(3708) <= layer5_outputs(2705);
    layer6_outputs(3709) <= layer5_outputs(7216);
    layer6_outputs(3710) <= '1';
    layer6_outputs(3711) <= '0';
    layer6_outputs(3712) <= not((layer5_outputs(6549)) and (layer5_outputs(8)));
    layer6_outputs(3713) <= (layer5_outputs(6427)) and not (layer5_outputs(6789));
    layer6_outputs(3714) <= not(layer5_outputs(4902));
    layer6_outputs(3715) <= layer5_outputs(3851);
    layer6_outputs(3716) <= layer5_outputs(4943);
    layer6_outputs(3717) <= layer5_outputs(7256);
    layer6_outputs(3718) <= layer5_outputs(26);
    layer6_outputs(3719) <= (layer5_outputs(3738)) and not (layer5_outputs(3399));
    layer6_outputs(3720) <= layer5_outputs(2239);
    layer6_outputs(3721) <= layer5_outputs(2190);
    layer6_outputs(3722) <= not(layer5_outputs(3698));
    layer6_outputs(3723) <= layer5_outputs(5791);
    layer6_outputs(3724) <= not(layer5_outputs(5853)) or (layer5_outputs(5766));
    layer6_outputs(3725) <= not((layer5_outputs(3083)) xor (layer5_outputs(7600)));
    layer6_outputs(3726) <= layer5_outputs(6839);
    layer6_outputs(3727) <= layer5_outputs(4347);
    layer6_outputs(3728) <= not(layer5_outputs(56));
    layer6_outputs(3729) <= (layer5_outputs(4071)) and (layer5_outputs(5599));
    layer6_outputs(3730) <= not(layer5_outputs(2969)) or (layer5_outputs(5528));
    layer6_outputs(3731) <= layer5_outputs(5659);
    layer6_outputs(3732) <= not(layer5_outputs(3077));
    layer6_outputs(3733) <= layer5_outputs(528);
    layer6_outputs(3734) <= (layer5_outputs(2867)) and not (layer5_outputs(2572));
    layer6_outputs(3735) <= layer5_outputs(262);
    layer6_outputs(3736) <= not(layer5_outputs(397)) or (layer5_outputs(3530));
    layer6_outputs(3737) <= not(layer5_outputs(4108)) or (layer5_outputs(3209));
    layer6_outputs(3738) <= layer5_outputs(4223);
    layer6_outputs(3739) <= not(layer5_outputs(1193));
    layer6_outputs(3740) <= not(layer5_outputs(5862));
    layer6_outputs(3741) <= not((layer5_outputs(1710)) xor (layer5_outputs(2340)));
    layer6_outputs(3742) <= not((layer5_outputs(1801)) or (layer5_outputs(2533)));
    layer6_outputs(3743) <= not(layer5_outputs(1410)) or (layer5_outputs(6987));
    layer6_outputs(3744) <= not((layer5_outputs(3962)) and (layer5_outputs(1980)));
    layer6_outputs(3745) <= not((layer5_outputs(377)) xor (layer5_outputs(464)));
    layer6_outputs(3746) <= (layer5_outputs(3531)) and not (layer5_outputs(677));
    layer6_outputs(3747) <= not(layer5_outputs(885)) or (layer5_outputs(6938));
    layer6_outputs(3748) <= layer5_outputs(2387);
    layer6_outputs(3749) <= (layer5_outputs(7670)) xor (layer5_outputs(539));
    layer6_outputs(3750) <= (layer5_outputs(2097)) and not (layer5_outputs(7341));
    layer6_outputs(3751) <= layer5_outputs(4189);
    layer6_outputs(3752) <= not((layer5_outputs(527)) xor (layer5_outputs(4525)));
    layer6_outputs(3753) <= layer5_outputs(150);
    layer6_outputs(3754) <= layer5_outputs(5947);
    layer6_outputs(3755) <= layer5_outputs(513);
    layer6_outputs(3756) <= not(layer5_outputs(6896));
    layer6_outputs(3757) <= not((layer5_outputs(2484)) xor (layer5_outputs(2063)));
    layer6_outputs(3758) <= (layer5_outputs(7074)) xor (layer5_outputs(3572));
    layer6_outputs(3759) <= not(layer5_outputs(4141));
    layer6_outputs(3760) <= layer5_outputs(809);
    layer6_outputs(3761) <= not(layer5_outputs(971));
    layer6_outputs(3762) <= (layer5_outputs(1735)) or (layer5_outputs(645));
    layer6_outputs(3763) <= not((layer5_outputs(4219)) and (layer5_outputs(7484)));
    layer6_outputs(3764) <= layer5_outputs(1638);
    layer6_outputs(3765) <= not(layer5_outputs(624));
    layer6_outputs(3766) <= not(layer5_outputs(2896));
    layer6_outputs(3767) <= not((layer5_outputs(1931)) or (layer5_outputs(3151)));
    layer6_outputs(3768) <= (layer5_outputs(2604)) and not (layer5_outputs(7123));
    layer6_outputs(3769) <= not((layer5_outputs(1057)) or (layer5_outputs(5200)));
    layer6_outputs(3770) <= (layer5_outputs(583)) and not (layer5_outputs(3431));
    layer6_outputs(3771) <= not(layer5_outputs(3527));
    layer6_outputs(3772) <= (layer5_outputs(3959)) and not (layer5_outputs(781));
    layer6_outputs(3773) <= layer5_outputs(4154);
    layer6_outputs(3774) <= not(layer5_outputs(616));
    layer6_outputs(3775) <= layer5_outputs(1836);
    layer6_outputs(3776) <= layer5_outputs(6846);
    layer6_outputs(3777) <= (layer5_outputs(5743)) and not (layer5_outputs(2834));
    layer6_outputs(3778) <= layer5_outputs(3949);
    layer6_outputs(3779) <= (layer5_outputs(5170)) and (layer5_outputs(789));
    layer6_outputs(3780) <= layer5_outputs(287);
    layer6_outputs(3781) <= not(layer5_outputs(4959));
    layer6_outputs(3782) <= layer5_outputs(4688);
    layer6_outputs(3783) <= (layer5_outputs(433)) and not (layer5_outputs(6370));
    layer6_outputs(3784) <= not(layer5_outputs(7097)) or (layer5_outputs(695));
    layer6_outputs(3785) <= layer5_outputs(2996);
    layer6_outputs(3786) <= (layer5_outputs(1310)) and not (layer5_outputs(5087));
    layer6_outputs(3787) <= layer5_outputs(1345);
    layer6_outputs(3788) <= not(layer5_outputs(4766));
    layer6_outputs(3789) <= not((layer5_outputs(3400)) xor (layer5_outputs(3845)));
    layer6_outputs(3790) <= (layer5_outputs(6483)) or (layer5_outputs(4508));
    layer6_outputs(3791) <= layer5_outputs(6793);
    layer6_outputs(3792) <= (layer5_outputs(3135)) or (layer5_outputs(2218));
    layer6_outputs(3793) <= layer5_outputs(7243);
    layer6_outputs(3794) <= layer5_outputs(6358);
    layer6_outputs(3795) <= not(layer5_outputs(398));
    layer6_outputs(3796) <= layer5_outputs(2000);
    layer6_outputs(3797) <= (layer5_outputs(4315)) xor (layer5_outputs(6908));
    layer6_outputs(3798) <= (layer5_outputs(4968)) xor (layer5_outputs(3807));
    layer6_outputs(3799) <= not((layer5_outputs(255)) xor (layer5_outputs(2856)));
    layer6_outputs(3800) <= not(layer5_outputs(6203));
    layer6_outputs(3801) <= not(layer5_outputs(49));
    layer6_outputs(3802) <= not((layer5_outputs(6393)) and (layer5_outputs(1499)));
    layer6_outputs(3803) <= not(layer5_outputs(1723));
    layer6_outputs(3804) <= not(layer5_outputs(5169));
    layer6_outputs(3805) <= not((layer5_outputs(1749)) xor (layer5_outputs(1325)));
    layer6_outputs(3806) <= not(layer5_outputs(3681));
    layer6_outputs(3807) <= not(layer5_outputs(7499));
    layer6_outputs(3808) <= not((layer5_outputs(6964)) or (layer5_outputs(5023)));
    layer6_outputs(3809) <= not(layer5_outputs(6351));
    layer6_outputs(3810) <= (layer5_outputs(2539)) and (layer5_outputs(3668));
    layer6_outputs(3811) <= layer5_outputs(162);
    layer6_outputs(3812) <= not((layer5_outputs(5482)) xor (layer5_outputs(4552)));
    layer6_outputs(3813) <= not(layer5_outputs(2311));
    layer6_outputs(3814) <= not(layer5_outputs(6299));
    layer6_outputs(3815) <= (layer5_outputs(6615)) and not (layer5_outputs(6271));
    layer6_outputs(3816) <= not((layer5_outputs(233)) and (layer5_outputs(3168)));
    layer6_outputs(3817) <= not(layer5_outputs(3671)) or (layer5_outputs(2127));
    layer6_outputs(3818) <= not(layer5_outputs(737));
    layer6_outputs(3819) <= not((layer5_outputs(3282)) xor (layer5_outputs(4296)));
    layer6_outputs(3820) <= layer5_outputs(2953);
    layer6_outputs(3821) <= not((layer5_outputs(4522)) and (layer5_outputs(811)));
    layer6_outputs(3822) <= (layer5_outputs(2550)) xor (layer5_outputs(5079));
    layer6_outputs(3823) <= not((layer5_outputs(5741)) xor (layer5_outputs(1684)));
    layer6_outputs(3824) <= not((layer5_outputs(5047)) and (layer5_outputs(7584)));
    layer6_outputs(3825) <= not(layer5_outputs(3599));
    layer6_outputs(3826) <= not(layer5_outputs(450));
    layer6_outputs(3827) <= (layer5_outputs(2010)) and not (layer5_outputs(1623));
    layer6_outputs(3828) <= not(layer5_outputs(2900)) or (layer5_outputs(7375));
    layer6_outputs(3829) <= not((layer5_outputs(6176)) xor (layer5_outputs(741)));
    layer6_outputs(3830) <= not(layer5_outputs(2517)) or (layer5_outputs(3821));
    layer6_outputs(3831) <= layer5_outputs(4812);
    layer6_outputs(3832) <= layer5_outputs(5435);
    layer6_outputs(3833) <= layer5_outputs(668);
    layer6_outputs(3834) <= (layer5_outputs(6071)) and not (layer5_outputs(1965));
    layer6_outputs(3835) <= (layer5_outputs(2763)) or (layer5_outputs(518));
    layer6_outputs(3836) <= not(layer5_outputs(395));
    layer6_outputs(3837) <= (layer5_outputs(6050)) or (layer5_outputs(7332));
    layer6_outputs(3838) <= not(layer5_outputs(2582));
    layer6_outputs(3839) <= not(layer5_outputs(4334));
    layer6_outputs(3840) <= layer5_outputs(1733);
    layer6_outputs(3841) <= layer5_outputs(3112);
    layer6_outputs(3842) <= (layer5_outputs(3515)) xor (layer5_outputs(5389));
    layer6_outputs(3843) <= not(layer5_outputs(352)) or (layer5_outputs(1149));
    layer6_outputs(3844) <= (layer5_outputs(5165)) and not (layer5_outputs(1579));
    layer6_outputs(3845) <= not(layer5_outputs(7310));
    layer6_outputs(3846) <= layer5_outputs(1607);
    layer6_outputs(3847) <= layer5_outputs(6698);
    layer6_outputs(3848) <= layer5_outputs(3527);
    layer6_outputs(3849) <= not(layer5_outputs(6330));
    layer6_outputs(3850) <= layer5_outputs(4974);
    layer6_outputs(3851) <= '0';
    layer6_outputs(3852) <= not(layer5_outputs(3809));
    layer6_outputs(3853) <= not((layer5_outputs(3425)) xor (layer5_outputs(6028)));
    layer6_outputs(3854) <= layer5_outputs(4151);
    layer6_outputs(3855) <= not(layer5_outputs(2787));
    layer6_outputs(3856) <= not(layer5_outputs(2315));
    layer6_outputs(3857) <= (layer5_outputs(5633)) and (layer5_outputs(2116));
    layer6_outputs(3858) <= (layer5_outputs(4863)) and (layer5_outputs(4664));
    layer6_outputs(3859) <= layer5_outputs(2360);
    layer6_outputs(3860) <= not((layer5_outputs(34)) xor (layer5_outputs(3374)));
    layer6_outputs(3861) <= (layer5_outputs(6901)) xor (layer5_outputs(5252));
    layer6_outputs(3862) <= not((layer5_outputs(4797)) and (layer5_outputs(2416)));
    layer6_outputs(3863) <= not(layer5_outputs(3349));
    layer6_outputs(3864) <= not(layer5_outputs(4663)) or (layer5_outputs(1002));
    layer6_outputs(3865) <= not(layer5_outputs(6304)) or (layer5_outputs(152));
    layer6_outputs(3866) <= layer5_outputs(1558);
    layer6_outputs(3867) <= (layer5_outputs(7530)) xor (layer5_outputs(533));
    layer6_outputs(3868) <= not(layer5_outputs(5375));
    layer6_outputs(3869) <= not((layer5_outputs(5893)) or (layer5_outputs(5085)));
    layer6_outputs(3870) <= layer5_outputs(3623);
    layer6_outputs(3871) <= layer5_outputs(1242);
    layer6_outputs(3872) <= (layer5_outputs(3585)) and (layer5_outputs(5111));
    layer6_outputs(3873) <= (layer5_outputs(3014)) and not (layer5_outputs(2209));
    layer6_outputs(3874) <= not(layer5_outputs(6844));
    layer6_outputs(3875) <= (layer5_outputs(7003)) xor (layer5_outputs(7052));
    layer6_outputs(3876) <= not(layer5_outputs(6486));
    layer6_outputs(3877) <= (layer5_outputs(842)) xor (layer5_outputs(1443));
    layer6_outputs(3878) <= layer5_outputs(269);
    layer6_outputs(3879) <= not((layer5_outputs(7245)) and (layer5_outputs(1037)));
    layer6_outputs(3880) <= not((layer5_outputs(1286)) and (layer5_outputs(275)));
    layer6_outputs(3881) <= (layer5_outputs(5444)) and (layer5_outputs(25));
    layer6_outputs(3882) <= not(layer5_outputs(1139)) or (layer5_outputs(3653));
    layer6_outputs(3883) <= not(layer5_outputs(941));
    layer6_outputs(3884) <= (layer5_outputs(6083)) or (layer5_outputs(806));
    layer6_outputs(3885) <= (layer5_outputs(2872)) xor (layer5_outputs(548));
    layer6_outputs(3886) <= not(layer5_outputs(4055)) or (layer5_outputs(5242));
    layer6_outputs(3887) <= not((layer5_outputs(6098)) xor (layer5_outputs(7282)));
    layer6_outputs(3888) <= not(layer5_outputs(3494));
    layer6_outputs(3889) <= '0';
    layer6_outputs(3890) <= layer5_outputs(2636);
    layer6_outputs(3891) <= layer5_outputs(2374);
    layer6_outputs(3892) <= not(layer5_outputs(3906)) or (layer5_outputs(7389));
    layer6_outputs(3893) <= layer5_outputs(1179);
    layer6_outputs(3894) <= layer5_outputs(1465);
    layer6_outputs(3895) <= layer5_outputs(5713);
    layer6_outputs(3896) <= layer5_outputs(4257);
    layer6_outputs(3897) <= not(layer5_outputs(4425));
    layer6_outputs(3898) <= layer5_outputs(2506);
    layer6_outputs(3899) <= not((layer5_outputs(1125)) xor (layer5_outputs(6721)));
    layer6_outputs(3900) <= (layer5_outputs(2738)) or (layer5_outputs(4056));
    layer6_outputs(3901) <= layer5_outputs(4515);
    layer6_outputs(3902) <= not((layer5_outputs(5379)) and (layer5_outputs(5970)));
    layer6_outputs(3903) <= (layer5_outputs(23)) xor (layer5_outputs(5634));
    layer6_outputs(3904) <= not(layer5_outputs(6320));
    layer6_outputs(3905) <= not(layer5_outputs(2371));
    layer6_outputs(3906) <= layer5_outputs(2407);
    layer6_outputs(3907) <= layer5_outputs(2611);
    layer6_outputs(3908) <= not(layer5_outputs(825));
    layer6_outputs(3909) <= not(layer5_outputs(2309));
    layer6_outputs(3910) <= (layer5_outputs(3305)) and not (layer5_outputs(3329));
    layer6_outputs(3911) <= (layer5_outputs(2582)) and not (layer5_outputs(3072));
    layer6_outputs(3912) <= not(layer5_outputs(6998));
    layer6_outputs(3913) <= (layer5_outputs(1114)) xor (layer5_outputs(5249));
    layer6_outputs(3914) <= not(layer5_outputs(3560));
    layer6_outputs(3915) <= (layer5_outputs(5635)) xor (layer5_outputs(6410));
    layer6_outputs(3916) <= not(layer5_outputs(5054));
    layer6_outputs(3917) <= layer5_outputs(5259);
    layer6_outputs(3918) <= (layer5_outputs(2175)) and not (layer5_outputs(1596));
    layer6_outputs(3919) <= not(layer5_outputs(2555)) or (layer5_outputs(3221));
    layer6_outputs(3920) <= layer5_outputs(2439);
    layer6_outputs(3921) <= (layer5_outputs(2088)) and (layer5_outputs(3853));
    layer6_outputs(3922) <= not(layer5_outputs(3310));
    layer6_outputs(3923) <= layer5_outputs(5439);
    layer6_outputs(3924) <= layer5_outputs(4039);
    layer6_outputs(3925) <= not(layer5_outputs(7091));
    layer6_outputs(3926) <= not(layer5_outputs(6910));
    layer6_outputs(3927) <= (layer5_outputs(4180)) xor (layer5_outputs(6673));
    layer6_outputs(3928) <= (layer5_outputs(6488)) xor (layer5_outputs(244));
    layer6_outputs(3929) <= not(layer5_outputs(409));
    layer6_outputs(3930) <= layer5_outputs(5450);
    layer6_outputs(3931) <= not(layer5_outputs(6959));
    layer6_outputs(3932) <= not(layer5_outputs(7435));
    layer6_outputs(3933) <= not(layer5_outputs(6786));
    layer6_outputs(3934) <= layer5_outputs(441);
    layer6_outputs(3935) <= layer5_outputs(2752);
    layer6_outputs(3936) <= (layer5_outputs(6175)) xor (layer5_outputs(4198));
    layer6_outputs(3937) <= layer5_outputs(4520);
    layer6_outputs(3938) <= '1';
    layer6_outputs(3939) <= (layer5_outputs(5018)) or (layer5_outputs(4987));
    layer6_outputs(3940) <= layer5_outputs(7581);
    layer6_outputs(3941) <= layer5_outputs(4351);
    layer6_outputs(3942) <= not(layer5_outputs(4137));
    layer6_outputs(3943) <= (layer5_outputs(6499)) and (layer5_outputs(1469));
    layer6_outputs(3944) <= not(layer5_outputs(2465));
    layer6_outputs(3945) <= layer5_outputs(1211);
    layer6_outputs(3946) <= layer5_outputs(2628);
    layer6_outputs(3947) <= not(layer5_outputs(408));
    layer6_outputs(3948) <= not((layer5_outputs(6119)) and (layer5_outputs(74)));
    layer6_outputs(3949) <= not(layer5_outputs(7291));
    layer6_outputs(3950) <= layer5_outputs(7263);
    layer6_outputs(3951) <= layer5_outputs(3948);
    layer6_outputs(3952) <= not((layer5_outputs(3556)) xor (layer5_outputs(383)));
    layer6_outputs(3953) <= (layer5_outputs(7542)) xor (layer5_outputs(7069));
    layer6_outputs(3954) <= layer5_outputs(6162);
    layer6_outputs(3955) <= not(layer5_outputs(5509));
    layer6_outputs(3956) <= (layer5_outputs(4390)) xor (layer5_outputs(1702));
    layer6_outputs(3957) <= not((layer5_outputs(861)) xor (layer5_outputs(3145)));
    layer6_outputs(3958) <= not((layer5_outputs(3483)) xor (layer5_outputs(3584)));
    layer6_outputs(3959) <= (layer5_outputs(1934)) or (layer5_outputs(6315));
    layer6_outputs(3960) <= not(layer5_outputs(6046)) or (layer5_outputs(2281));
    layer6_outputs(3961) <= not(layer5_outputs(6631));
    layer6_outputs(3962) <= '0';
    layer6_outputs(3963) <= not((layer5_outputs(2209)) or (layer5_outputs(1820)));
    layer6_outputs(3964) <= not(layer5_outputs(5008));
    layer6_outputs(3965) <= not(layer5_outputs(4323));
    layer6_outputs(3966) <= not((layer5_outputs(7007)) xor (layer5_outputs(83)));
    layer6_outputs(3967) <= (layer5_outputs(1553)) and not (layer5_outputs(5842));
    layer6_outputs(3968) <= not((layer5_outputs(628)) xor (layer5_outputs(3328)));
    layer6_outputs(3969) <= (layer5_outputs(2156)) and not (layer5_outputs(768));
    layer6_outputs(3970) <= not(layer5_outputs(6236));
    layer6_outputs(3971) <= not(layer5_outputs(6057));
    layer6_outputs(3972) <= layer5_outputs(3869);
    layer6_outputs(3973) <= layer5_outputs(2210);
    layer6_outputs(3974) <= '1';
    layer6_outputs(3975) <= not(layer5_outputs(4052));
    layer6_outputs(3976) <= not(layer5_outputs(5898));
    layer6_outputs(3977) <= not((layer5_outputs(4897)) and (layer5_outputs(5274)));
    layer6_outputs(3978) <= not(layer5_outputs(3875));
    layer6_outputs(3979) <= not(layer5_outputs(4165));
    layer6_outputs(3980) <= (layer5_outputs(3976)) and not (layer5_outputs(6567));
    layer6_outputs(3981) <= not(layer5_outputs(3673));
    layer6_outputs(3982) <= layer5_outputs(1713);
    layer6_outputs(3983) <= not((layer5_outputs(5656)) xor (layer5_outputs(6472)));
    layer6_outputs(3984) <= (layer5_outputs(1368)) xor (layer5_outputs(3033));
    layer6_outputs(3985) <= layer5_outputs(5751);
    layer6_outputs(3986) <= layer5_outputs(2722);
    layer6_outputs(3987) <= not(layer5_outputs(1612));
    layer6_outputs(3988) <= not((layer5_outputs(3729)) xor (layer5_outputs(2051)));
    layer6_outputs(3989) <= layer5_outputs(5638);
    layer6_outputs(3990) <= not(layer5_outputs(384));
    layer6_outputs(3991) <= (layer5_outputs(5332)) xor (layer5_outputs(6834));
    layer6_outputs(3992) <= (layer5_outputs(597)) and not (layer5_outputs(1646));
    layer6_outputs(3993) <= not(layer5_outputs(4689));
    layer6_outputs(3994) <= layer5_outputs(5507);
    layer6_outputs(3995) <= (layer5_outputs(981)) or (layer5_outputs(5478));
    layer6_outputs(3996) <= layer5_outputs(2019);
    layer6_outputs(3997) <= not(layer5_outputs(7473));
    layer6_outputs(3998) <= not(layer5_outputs(6567));
    layer6_outputs(3999) <= (layer5_outputs(2000)) xor (layer5_outputs(1092));
    layer6_outputs(4000) <= (layer5_outputs(3479)) xor (layer5_outputs(5832));
    layer6_outputs(4001) <= (layer5_outputs(3195)) xor (layer5_outputs(3345));
    layer6_outputs(4002) <= layer5_outputs(4633);
    layer6_outputs(4003) <= (layer5_outputs(2497)) xor (layer5_outputs(2764));
    layer6_outputs(4004) <= layer5_outputs(6436);
    layer6_outputs(4005) <= (layer5_outputs(7627)) or (layer5_outputs(2403));
    layer6_outputs(4006) <= not(layer5_outputs(6951));
    layer6_outputs(4007) <= not(layer5_outputs(4976));
    layer6_outputs(4008) <= layer5_outputs(1734);
    layer6_outputs(4009) <= not(layer5_outputs(7234));
    layer6_outputs(4010) <= not(layer5_outputs(7129));
    layer6_outputs(4011) <= (layer5_outputs(3270)) or (layer5_outputs(4239));
    layer6_outputs(4012) <= (layer5_outputs(190)) and not (layer5_outputs(129));
    layer6_outputs(4013) <= not(layer5_outputs(4656)) or (layer5_outputs(4857));
    layer6_outputs(4014) <= layer5_outputs(7368);
    layer6_outputs(4015) <= (layer5_outputs(6694)) and not (layer5_outputs(2954));
    layer6_outputs(4016) <= layer5_outputs(1328);
    layer6_outputs(4017) <= (layer5_outputs(2393)) or (layer5_outputs(6875));
    layer6_outputs(4018) <= not((layer5_outputs(4412)) xor (layer5_outputs(4343)));
    layer6_outputs(4019) <= not((layer5_outputs(571)) xor (layer5_outputs(177)));
    layer6_outputs(4020) <= not((layer5_outputs(7008)) xor (layer5_outputs(6640)));
    layer6_outputs(4021) <= not((layer5_outputs(7284)) or (layer5_outputs(294)));
    layer6_outputs(4022) <= not(layer5_outputs(4126));
    layer6_outputs(4023) <= not(layer5_outputs(980));
    layer6_outputs(4024) <= layer5_outputs(6282);
    layer6_outputs(4025) <= not(layer5_outputs(554));
    layer6_outputs(4026) <= (layer5_outputs(2910)) or (layer5_outputs(4714));
    layer6_outputs(4027) <= (layer5_outputs(2602)) and not (layer5_outputs(6712));
    layer6_outputs(4028) <= not((layer5_outputs(3658)) and (layer5_outputs(1835)));
    layer6_outputs(4029) <= (layer5_outputs(6028)) and not (layer5_outputs(5543));
    layer6_outputs(4030) <= not(layer5_outputs(6939)) or (layer5_outputs(2817));
    layer6_outputs(4031) <= (layer5_outputs(35)) xor (layer5_outputs(2199));
    layer6_outputs(4032) <= not(layer5_outputs(4784));
    layer6_outputs(4033) <= not(layer5_outputs(6406)) or (layer5_outputs(2757));
    layer6_outputs(4034) <= not((layer5_outputs(2170)) xor (layer5_outputs(6364)));
    layer6_outputs(4035) <= not((layer5_outputs(5764)) and (layer5_outputs(7527)));
    layer6_outputs(4036) <= (layer5_outputs(3393)) xor (layer5_outputs(2181));
    layer6_outputs(4037) <= not((layer5_outputs(6819)) xor (layer5_outputs(802)));
    layer6_outputs(4038) <= layer5_outputs(425);
    layer6_outputs(4039) <= (layer5_outputs(2683)) xor (layer5_outputs(4467));
    layer6_outputs(4040) <= not(layer5_outputs(3894));
    layer6_outputs(4041) <= layer5_outputs(316);
    layer6_outputs(4042) <= not(layer5_outputs(1736));
    layer6_outputs(4043) <= (layer5_outputs(6130)) and (layer5_outputs(4543));
    layer6_outputs(4044) <= not(layer5_outputs(2264));
    layer6_outputs(4045) <= (layer5_outputs(2680)) or (layer5_outputs(3122));
    layer6_outputs(4046) <= not(layer5_outputs(2440));
    layer6_outputs(4047) <= not((layer5_outputs(5559)) and (layer5_outputs(5593)));
    layer6_outputs(4048) <= not(layer5_outputs(7186)) or (layer5_outputs(4168));
    layer6_outputs(4049) <= not(layer5_outputs(4292));
    layer6_outputs(4050) <= (layer5_outputs(1692)) and not (layer5_outputs(2949));
    layer6_outputs(4051) <= not((layer5_outputs(5651)) xor (layer5_outputs(5457)));
    layer6_outputs(4052) <= layer5_outputs(1983);
    layer6_outputs(4053) <= not(layer5_outputs(5989));
    layer6_outputs(4054) <= (layer5_outputs(298)) and not (layer5_outputs(4343));
    layer6_outputs(4055) <= (layer5_outputs(1149)) and (layer5_outputs(474));
    layer6_outputs(4056) <= (layer5_outputs(4258)) and (layer5_outputs(7512));
    layer6_outputs(4057) <= not((layer5_outputs(5376)) xor (layer5_outputs(267)));
    layer6_outputs(4058) <= layer5_outputs(4728);
    layer6_outputs(4059) <= not(layer5_outputs(5514));
    layer6_outputs(4060) <= (layer5_outputs(1759)) xor (layer5_outputs(2280));
    layer6_outputs(4061) <= (layer5_outputs(4482)) and not (layer5_outputs(4410));
    layer6_outputs(4062) <= layer5_outputs(2232);
    layer6_outputs(4063) <= layer5_outputs(4061);
    layer6_outputs(4064) <= layer5_outputs(6408);
    layer6_outputs(4065) <= layer5_outputs(320);
    layer6_outputs(4066) <= not((layer5_outputs(1864)) or (layer5_outputs(1495)));
    layer6_outputs(4067) <= layer5_outputs(1706);
    layer6_outputs(4068) <= not((layer5_outputs(7121)) or (layer5_outputs(5781)));
    layer6_outputs(4069) <= not((layer5_outputs(6655)) or (layer5_outputs(6633)));
    layer6_outputs(4070) <= not((layer5_outputs(4030)) xor (layer5_outputs(5114)));
    layer6_outputs(4071) <= layer5_outputs(6970);
    layer6_outputs(4072) <= layer5_outputs(3286);
    layer6_outputs(4073) <= not(layer5_outputs(4604));
    layer6_outputs(4074) <= layer5_outputs(1481);
    layer6_outputs(4075) <= (layer5_outputs(5196)) and not (layer5_outputs(3240));
    layer6_outputs(4076) <= layer5_outputs(4103);
    layer6_outputs(4077) <= not(layer5_outputs(3634));
    layer6_outputs(4078) <= '0';
    layer6_outputs(4079) <= layer5_outputs(7677);
    layer6_outputs(4080) <= (layer5_outputs(3104)) and not (layer5_outputs(610));
    layer6_outputs(4081) <= not((layer5_outputs(6856)) xor (layer5_outputs(5528)));
    layer6_outputs(4082) <= not(layer5_outputs(997));
    layer6_outputs(4083) <= (layer5_outputs(800)) and not (layer5_outputs(5265));
    layer6_outputs(4084) <= (layer5_outputs(3361)) and not (layer5_outputs(3514));
    layer6_outputs(4085) <= layer5_outputs(2787);
    layer6_outputs(4086) <= layer5_outputs(428);
    layer6_outputs(4087) <= not(layer5_outputs(2193));
    layer6_outputs(4088) <= not(layer5_outputs(6538));
    layer6_outputs(4089) <= not(layer5_outputs(3476));
    layer6_outputs(4090) <= (layer5_outputs(4616)) xor (layer5_outputs(3670));
    layer6_outputs(4091) <= not((layer5_outputs(6570)) xor (layer5_outputs(5621)));
    layer6_outputs(4092) <= layer5_outputs(4023);
    layer6_outputs(4093) <= layer5_outputs(7065);
    layer6_outputs(4094) <= not((layer5_outputs(1275)) and (layer5_outputs(4293)));
    layer6_outputs(4095) <= not(layer5_outputs(7259));
    layer6_outputs(4096) <= (layer5_outputs(7111)) and (layer5_outputs(54));
    layer6_outputs(4097) <= not(layer5_outputs(3573));
    layer6_outputs(4098) <= not(layer5_outputs(6814));
    layer6_outputs(4099) <= layer5_outputs(5787);
    layer6_outputs(4100) <= not(layer5_outputs(2638));
    layer6_outputs(4101) <= not(layer5_outputs(7154));
    layer6_outputs(4102) <= layer5_outputs(7483);
    layer6_outputs(4103) <= (layer5_outputs(5343)) xor (layer5_outputs(693));
    layer6_outputs(4104) <= not((layer5_outputs(3714)) xor (layer5_outputs(3681)));
    layer6_outputs(4105) <= not((layer5_outputs(5381)) and (layer5_outputs(2455)));
    layer6_outputs(4106) <= layer5_outputs(2989);
    layer6_outputs(4107) <= (layer5_outputs(4832)) xor (layer5_outputs(6369));
    layer6_outputs(4108) <= not(layer5_outputs(6362));
    layer6_outputs(4109) <= layer5_outputs(6334);
    layer6_outputs(4110) <= (layer5_outputs(2)) and (layer5_outputs(2898));
    layer6_outputs(4111) <= not(layer5_outputs(7668)) or (layer5_outputs(6938));
    layer6_outputs(4112) <= not(layer5_outputs(1861));
    layer6_outputs(4113) <= layer5_outputs(1205);
    layer6_outputs(4114) <= layer5_outputs(3102);
    layer6_outputs(4115) <= (layer5_outputs(631)) and not (layer5_outputs(4700));
    layer6_outputs(4116) <= (layer5_outputs(5901)) xor (layer5_outputs(4297));
    layer6_outputs(4117) <= not(layer5_outputs(5269));
    layer6_outputs(4118) <= (layer5_outputs(3185)) and not (layer5_outputs(3286));
    layer6_outputs(4119) <= layer5_outputs(659);
    layer6_outputs(4120) <= (layer5_outputs(6737)) xor (layer5_outputs(679));
    layer6_outputs(4121) <= not((layer5_outputs(1524)) or (layer5_outputs(4955)));
    layer6_outputs(4122) <= not(layer5_outputs(6357));
    layer6_outputs(4123) <= layer5_outputs(4965);
    layer6_outputs(4124) <= layer5_outputs(1131);
    layer6_outputs(4125) <= (layer5_outputs(435)) xor (layer5_outputs(3255));
    layer6_outputs(4126) <= layer5_outputs(7054);
    layer6_outputs(4127) <= not((layer5_outputs(7304)) and (layer5_outputs(2078)));
    layer6_outputs(4128) <= '0';
    layer6_outputs(4129) <= (layer5_outputs(6433)) and not (layer5_outputs(3229));
    layer6_outputs(4130) <= layer5_outputs(1999);
    layer6_outputs(4131) <= not(layer5_outputs(1179));
    layer6_outputs(4132) <= not((layer5_outputs(2865)) xor (layer5_outputs(1325)));
    layer6_outputs(4133) <= not((layer5_outputs(2254)) and (layer5_outputs(4510)));
    layer6_outputs(4134) <= not((layer5_outputs(3100)) xor (layer5_outputs(3365)));
    layer6_outputs(4135) <= (layer5_outputs(4277)) or (layer5_outputs(1177));
    layer6_outputs(4136) <= not((layer5_outputs(6514)) or (layer5_outputs(4402)));
    layer6_outputs(4137) <= not(layer5_outputs(7176));
    layer6_outputs(4138) <= layer5_outputs(493);
    layer6_outputs(4139) <= not(layer5_outputs(5776)) or (layer5_outputs(3596));
    layer6_outputs(4140) <= not(layer5_outputs(5692));
    layer6_outputs(4141) <= not((layer5_outputs(3418)) or (layer5_outputs(2697)));
    layer6_outputs(4142) <= not((layer5_outputs(2797)) or (layer5_outputs(2943)));
    layer6_outputs(4143) <= not(layer5_outputs(608)) or (layer5_outputs(696));
    layer6_outputs(4144) <= layer5_outputs(7151);
    layer6_outputs(4145) <= layer5_outputs(5092);
    layer6_outputs(4146) <= (layer5_outputs(5455)) or (layer5_outputs(4010));
    layer6_outputs(4147) <= not(layer5_outputs(6622));
    layer6_outputs(4148) <= (layer5_outputs(420)) or (layer5_outputs(7565));
    layer6_outputs(4149) <= (layer5_outputs(4023)) xor (layer5_outputs(5686));
    layer6_outputs(4150) <= '0';
    layer6_outputs(4151) <= not(layer5_outputs(7606)) or (layer5_outputs(4480));
    layer6_outputs(4152) <= layer5_outputs(3209);
    layer6_outputs(4153) <= not((layer5_outputs(1281)) and (layer5_outputs(4885)));
    layer6_outputs(4154) <= not(layer5_outputs(1503)) or (layer5_outputs(5813));
    layer6_outputs(4155) <= not(layer5_outputs(7572)) or (layer5_outputs(7192));
    layer6_outputs(4156) <= layer5_outputs(6253);
    layer6_outputs(4157) <= (layer5_outputs(2850)) and not (layer5_outputs(3126));
    layer6_outputs(4158) <= not(layer5_outputs(999));
    layer6_outputs(4159) <= not(layer5_outputs(2786));
    layer6_outputs(4160) <= not(layer5_outputs(640));
    layer6_outputs(4161) <= (layer5_outputs(7410)) xor (layer5_outputs(349));
    layer6_outputs(4162) <= (layer5_outputs(5981)) and not (layer5_outputs(6268));
    layer6_outputs(4163) <= not((layer5_outputs(3338)) xor (layer5_outputs(1234)));
    layer6_outputs(4164) <= not(layer5_outputs(7112)) or (layer5_outputs(312));
    layer6_outputs(4165) <= not((layer5_outputs(7589)) and (layer5_outputs(1078)));
    layer6_outputs(4166) <= not(layer5_outputs(3296));
    layer6_outputs(4167) <= layer5_outputs(1308);
    layer6_outputs(4168) <= not(layer5_outputs(4774));
    layer6_outputs(4169) <= not(layer5_outputs(1882));
    layer6_outputs(4170) <= layer5_outputs(6971);
    layer6_outputs(4171) <= (layer5_outputs(3844)) and not (layer5_outputs(2879));
    layer6_outputs(4172) <= not(layer5_outputs(3083)) or (layer5_outputs(2297));
    layer6_outputs(4173) <= (layer5_outputs(3107)) and not (layer5_outputs(4076));
    layer6_outputs(4174) <= layer5_outputs(3126);
    layer6_outputs(4175) <= not(layer5_outputs(2695));
    layer6_outputs(4176) <= (layer5_outputs(1302)) xor (layer5_outputs(836));
    layer6_outputs(4177) <= '1';
    layer6_outputs(4178) <= not(layer5_outputs(1688));
    layer6_outputs(4179) <= not(layer5_outputs(2779));
    layer6_outputs(4180) <= not((layer5_outputs(626)) or (layer5_outputs(4523)));
    layer6_outputs(4181) <= layer5_outputs(7206);
    layer6_outputs(4182) <= (layer5_outputs(3138)) xor (layer5_outputs(976));
    layer6_outputs(4183) <= (layer5_outputs(5833)) and not (layer5_outputs(4150));
    layer6_outputs(4184) <= layer5_outputs(6511);
    layer6_outputs(4185) <= not(layer5_outputs(5194));
    layer6_outputs(4186) <= (layer5_outputs(2702)) and (layer5_outputs(2328));
    layer6_outputs(4187) <= not(layer5_outputs(1349));
    layer6_outputs(4188) <= not(layer5_outputs(2188));
    layer6_outputs(4189) <= not(layer5_outputs(1099));
    layer6_outputs(4190) <= layer5_outputs(4850);
    layer6_outputs(4191) <= layer5_outputs(1113);
    layer6_outputs(4192) <= '1';
    layer6_outputs(4193) <= (layer5_outputs(4783)) or (layer5_outputs(6691));
    layer6_outputs(4194) <= not((layer5_outputs(4911)) xor (layer5_outputs(202)));
    layer6_outputs(4195) <= '1';
    layer6_outputs(4196) <= not((layer5_outputs(3204)) xor (layer5_outputs(1521)));
    layer6_outputs(4197) <= layer5_outputs(1612);
    layer6_outputs(4198) <= not(layer5_outputs(6992));
    layer6_outputs(4199) <= not((layer5_outputs(1853)) xor (layer5_outputs(200)));
    layer6_outputs(4200) <= not((layer5_outputs(5813)) and (layer5_outputs(1256)));
    layer6_outputs(4201) <= not(layer5_outputs(5064));
    layer6_outputs(4202) <= not(layer5_outputs(4298));
    layer6_outputs(4203) <= layer5_outputs(2747);
    layer6_outputs(4204) <= (layer5_outputs(4891)) xor (layer5_outputs(7070));
    layer6_outputs(4205) <= layer5_outputs(2189);
    layer6_outputs(4206) <= not(layer5_outputs(5262));
    layer6_outputs(4207) <= (layer5_outputs(2255)) or (layer5_outputs(5331));
    layer6_outputs(4208) <= not(layer5_outputs(7336));
    layer6_outputs(4209) <= not(layer5_outputs(5818));
    layer6_outputs(4210) <= layer5_outputs(7612);
    layer6_outputs(4211) <= (layer5_outputs(5754)) and (layer5_outputs(5042));
    layer6_outputs(4212) <= layer5_outputs(1546);
    layer6_outputs(4213) <= (layer5_outputs(3057)) or (layer5_outputs(240));
    layer6_outputs(4214) <= (layer5_outputs(5660)) and (layer5_outputs(2067));
    layer6_outputs(4215) <= not(layer5_outputs(3253)) or (layer5_outputs(4848));
    layer6_outputs(4216) <= not(layer5_outputs(7556));
    layer6_outputs(4217) <= layer5_outputs(2107);
    layer6_outputs(4218) <= layer5_outputs(728);
    layer6_outputs(4219) <= layer5_outputs(29);
    layer6_outputs(4220) <= not(layer5_outputs(6304));
    layer6_outputs(4221) <= layer5_outputs(681);
    layer6_outputs(4222) <= not(layer5_outputs(829));
    layer6_outputs(4223) <= (layer5_outputs(5982)) and (layer5_outputs(5614));
    layer6_outputs(4224) <= (layer5_outputs(6281)) xor (layer5_outputs(2793));
    layer6_outputs(4225) <= not(layer5_outputs(5662));
    layer6_outputs(4226) <= (layer5_outputs(3810)) and not (layer5_outputs(1373));
    layer6_outputs(4227) <= layer5_outputs(2963);
    layer6_outputs(4228) <= (layer5_outputs(1867)) and not (layer5_outputs(4133));
    layer6_outputs(4229) <= not((layer5_outputs(594)) xor (layer5_outputs(4993)));
    layer6_outputs(4230) <= not((layer5_outputs(3939)) and (layer5_outputs(2845)));
    layer6_outputs(4231) <= not((layer5_outputs(727)) xor (layer5_outputs(2015)));
    layer6_outputs(4232) <= not(layer5_outputs(5067));
    layer6_outputs(4233) <= not(layer5_outputs(780));
    layer6_outputs(4234) <= layer5_outputs(6167);
    layer6_outputs(4235) <= not(layer5_outputs(4996)) or (layer5_outputs(4249));
    layer6_outputs(4236) <= not(layer5_outputs(6953));
    layer6_outputs(4237) <= (layer5_outputs(1289)) xor (layer5_outputs(7421));
    layer6_outputs(4238) <= not(layer5_outputs(2589));
    layer6_outputs(4239) <= not(layer5_outputs(1811)) or (layer5_outputs(6077));
    layer6_outputs(4240) <= (layer5_outputs(6805)) and not (layer5_outputs(1575));
    layer6_outputs(4241) <= (layer5_outputs(110)) and (layer5_outputs(618));
    layer6_outputs(4242) <= not(layer5_outputs(6363)) or (layer5_outputs(2938));
    layer6_outputs(4243) <= (layer5_outputs(6124)) and not (layer5_outputs(4913));
    layer6_outputs(4244) <= not((layer5_outputs(2806)) or (layer5_outputs(232)));
    layer6_outputs(4245) <= not(layer5_outputs(5572));
    layer6_outputs(4246) <= layer5_outputs(2179);
    layer6_outputs(4247) <= not(layer5_outputs(4024));
    layer6_outputs(4248) <= not(layer5_outputs(998));
    layer6_outputs(4249) <= (layer5_outputs(35)) and (layer5_outputs(2431));
    layer6_outputs(4250) <= layer5_outputs(702);
    layer6_outputs(4251) <= layer5_outputs(4637);
    layer6_outputs(4252) <= (layer5_outputs(1261)) and (layer5_outputs(4875));
    layer6_outputs(4253) <= not(layer5_outputs(3515));
    layer6_outputs(4254) <= layer5_outputs(6932);
    layer6_outputs(4255) <= not(layer5_outputs(5298));
    layer6_outputs(4256) <= (layer5_outputs(1194)) or (layer5_outputs(368));
    layer6_outputs(4257) <= (layer5_outputs(776)) and not (layer5_outputs(1546));
    layer6_outputs(4258) <= not(layer5_outputs(605));
    layer6_outputs(4259) <= not(layer5_outputs(6005));
    layer6_outputs(4260) <= (layer5_outputs(5419)) and (layer5_outputs(2476));
    layer6_outputs(4261) <= not(layer5_outputs(7631));
    layer6_outputs(4262) <= not((layer5_outputs(6555)) xor (layer5_outputs(5964)));
    layer6_outputs(4263) <= layer5_outputs(5372);
    layer6_outputs(4264) <= layer5_outputs(137);
    layer6_outputs(4265) <= not((layer5_outputs(7278)) xor (layer5_outputs(3301)));
    layer6_outputs(4266) <= (layer5_outputs(682)) or (layer5_outputs(5339));
    layer6_outputs(4267) <= (layer5_outputs(4501)) or (layer5_outputs(5405));
    layer6_outputs(4268) <= (layer5_outputs(5419)) and (layer5_outputs(7522));
    layer6_outputs(4269) <= not(layer5_outputs(543));
    layer6_outputs(4270) <= not(layer5_outputs(4909));
    layer6_outputs(4271) <= not(layer5_outputs(7662));
    layer6_outputs(4272) <= (layer5_outputs(1606)) and (layer5_outputs(6426));
    layer6_outputs(4273) <= (layer5_outputs(6844)) and not (layer5_outputs(6723));
    layer6_outputs(4274) <= (layer5_outputs(5424)) or (layer5_outputs(330));
    layer6_outputs(4275) <= not((layer5_outputs(1384)) and (layer5_outputs(2155)));
    layer6_outputs(4276) <= not((layer5_outputs(5328)) and (layer5_outputs(5742)));
    layer6_outputs(4277) <= not(layer5_outputs(4473));
    layer6_outputs(4278) <= (layer5_outputs(419)) xor (layer5_outputs(3035));
    layer6_outputs(4279) <= not(layer5_outputs(4528));
    layer6_outputs(4280) <= not(layer5_outputs(3128));
    layer6_outputs(4281) <= '1';
    layer6_outputs(4282) <= not(layer5_outputs(2892));
    layer6_outputs(4283) <= layer5_outputs(72);
    layer6_outputs(4284) <= '0';
    layer6_outputs(4285) <= not((layer5_outputs(3726)) xor (layer5_outputs(2356)));
    layer6_outputs(4286) <= not(layer5_outputs(2502));
    layer6_outputs(4287) <= layer5_outputs(6471);
    layer6_outputs(4288) <= (layer5_outputs(4568)) and (layer5_outputs(3808));
    layer6_outputs(4289) <= not(layer5_outputs(1130));
    layer6_outputs(4290) <= not(layer5_outputs(7617));
    layer6_outputs(4291) <= (layer5_outputs(3948)) and not (layer5_outputs(7501));
    layer6_outputs(4292) <= not(layer5_outputs(5566));
    layer6_outputs(4293) <= not((layer5_outputs(1430)) xor (layer5_outputs(4794)));
    layer6_outputs(4294) <= not(layer5_outputs(5953));
    layer6_outputs(4295) <= not(layer5_outputs(141));
    layer6_outputs(4296) <= layer5_outputs(198);
    layer6_outputs(4297) <= not((layer5_outputs(6335)) or (layer5_outputs(5768)));
    layer6_outputs(4298) <= not((layer5_outputs(4318)) or (layer5_outputs(2661)));
    layer6_outputs(4299) <= not(layer5_outputs(2202));
    layer6_outputs(4300) <= not(layer5_outputs(7430));
    layer6_outputs(4301) <= not((layer5_outputs(7249)) xor (layer5_outputs(3725)));
    layer6_outputs(4302) <= layer5_outputs(7192);
    layer6_outputs(4303) <= layer5_outputs(1767);
    layer6_outputs(4304) <= layer5_outputs(614);
    layer6_outputs(4305) <= (layer5_outputs(5943)) and not (layer5_outputs(2397));
    layer6_outputs(4306) <= not(layer5_outputs(4164));
    layer6_outputs(4307) <= not((layer5_outputs(7635)) xor (layer5_outputs(6039)));
    layer6_outputs(4308) <= '1';
    layer6_outputs(4309) <= layer5_outputs(5135);
    layer6_outputs(4310) <= layer5_outputs(4673);
    layer6_outputs(4311) <= layer5_outputs(5496);
    layer6_outputs(4312) <= not(layer5_outputs(2831));
    layer6_outputs(4313) <= layer5_outputs(5076);
    layer6_outputs(4314) <= (layer5_outputs(6613)) or (layer5_outputs(1615));
    layer6_outputs(4315) <= not((layer5_outputs(6767)) xor (layer5_outputs(1752)));
    layer6_outputs(4316) <= layer5_outputs(6619);
    layer6_outputs(4317) <= (layer5_outputs(1812)) and not (layer5_outputs(607));
    layer6_outputs(4318) <= layer5_outputs(3140);
    layer6_outputs(4319) <= not(layer5_outputs(2345));
    layer6_outputs(4320) <= (layer5_outputs(2004)) and not (layer5_outputs(4399));
    layer6_outputs(4321) <= (layer5_outputs(6897)) xor (layer5_outputs(1603));
    layer6_outputs(4322) <= (layer5_outputs(5924)) and (layer5_outputs(6195));
    layer6_outputs(4323) <= (layer5_outputs(1875)) xor (layer5_outputs(5569));
    layer6_outputs(4324) <= not(layer5_outputs(2587));
    layer6_outputs(4325) <= not(layer5_outputs(4027));
    layer6_outputs(4326) <= not(layer5_outputs(7560));
    layer6_outputs(4327) <= not(layer5_outputs(5076)) or (layer5_outputs(6501));
    layer6_outputs(4328) <= not((layer5_outputs(5995)) or (layer5_outputs(6968)));
    layer6_outputs(4329) <= not(layer5_outputs(1342));
    layer6_outputs(4330) <= layer5_outputs(1789);
    layer6_outputs(4331) <= layer5_outputs(7020);
    layer6_outputs(4332) <= not(layer5_outputs(731));
    layer6_outputs(4333) <= layer5_outputs(388);
    layer6_outputs(4334) <= layer5_outputs(1559);
    layer6_outputs(4335) <= layer5_outputs(1348);
    layer6_outputs(4336) <= (layer5_outputs(7458)) and not (layer5_outputs(5838));
    layer6_outputs(4337) <= (layer5_outputs(4405)) xor (layer5_outputs(6936));
    layer6_outputs(4338) <= (layer5_outputs(4859)) and not (layer5_outputs(1877));
    layer6_outputs(4339) <= layer5_outputs(731);
    layer6_outputs(4340) <= not((layer5_outputs(5280)) and (layer5_outputs(5308)));
    layer6_outputs(4341) <= (layer5_outputs(4033)) and not (layer5_outputs(2454));
    layer6_outputs(4342) <= (layer5_outputs(688)) xor (layer5_outputs(3241));
    layer6_outputs(4343) <= not(layer5_outputs(7468));
    layer6_outputs(4344) <= layer5_outputs(4237);
    layer6_outputs(4345) <= (layer5_outputs(5904)) xor (layer5_outputs(5385));
    layer6_outputs(4346) <= layer5_outputs(1530);
    layer6_outputs(4347) <= not(layer5_outputs(2599));
    layer6_outputs(4348) <= (layer5_outputs(2975)) or (layer5_outputs(3090));
    layer6_outputs(4349) <= layer5_outputs(2032);
    layer6_outputs(4350) <= not(layer5_outputs(1289)) or (layer5_outputs(1513));
    layer6_outputs(4351) <= not(layer5_outputs(370));
    layer6_outputs(4352) <= (layer5_outputs(5241)) and not (layer5_outputs(4005));
    layer6_outputs(4353) <= '0';
    layer6_outputs(4354) <= layer5_outputs(2904);
    layer6_outputs(4355) <= not(layer5_outputs(6686));
    layer6_outputs(4356) <= layer5_outputs(4056);
    layer6_outputs(4357) <= not((layer5_outputs(613)) and (layer5_outputs(3788)));
    layer6_outputs(4358) <= not((layer5_outputs(6514)) xor (layer5_outputs(6743)));
    layer6_outputs(4359) <= (layer5_outputs(20)) and (layer5_outputs(884));
    layer6_outputs(4360) <= (layer5_outputs(2250)) and not (layer5_outputs(3733));
    layer6_outputs(4361) <= layer5_outputs(3688);
    layer6_outputs(4362) <= (layer5_outputs(653)) or (layer5_outputs(1793));
    layer6_outputs(4363) <= not(layer5_outputs(448));
    layer6_outputs(4364) <= (layer5_outputs(1648)) xor (layer5_outputs(7639));
    layer6_outputs(4365) <= not(layer5_outputs(2402));
    layer6_outputs(4366) <= layer5_outputs(1802);
    layer6_outputs(4367) <= layer5_outputs(4422);
    layer6_outputs(4368) <= not(layer5_outputs(1362));
    layer6_outputs(4369) <= layer5_outputs(4869);
    layer6_outputs(4370) <= layer5_outputs(2681);
    layer6_outputs(4371) <= (layer5_outputs(6206)) xor (layer5_outputs(4732));
    layer6_outputs(4372) <= layer5_outputs(2244);
    layer6_outputs(4373) <= not(layer5_outputs(3358));
    layer6_outputs(4374) <= not(layer5_outputs(5087));
    layer6_outputs(4375) <= not(layer5_outputs(5235));
    layer6_outputs(4376) <= (layer5_outputs(6322)) xor (layer5_outputs(5814));
    layer6_outputs(4377) <= (layer5_outputs(390)) xor (layer5_outputs(2061));
    layer6_outputs(4378) <= not(layer5_outputs(1786));
    layer6_outputs(4379) <= not(layer5_outputs(2592));
    layer6_outputs(4380) <= layer5_outputs(3033);
    layer6_outputs(4381) <= not(layer5_outputs(444));
    layer6_outputs(4382) <= not(layer5_outputs(2820));
    layer6_outputs(4383) <= (layer5_outputs(1483)) xor (layer5_outputs(1217));
    layer6_outputs(4384) <= (layer5_outputs(5772)) or (layer5_outputs(3046));
    layer6_outputs(4385) <= layer5_outputs(6822);
    layer6_outputs(4386) <= layer5_outputs(1452);
    layer6_outputs(4387) <= not((layer5_outputs(4807)) xor (layer5_outputs(6091)));
    layer6_outputs(4388) <= not((layer5_outputs(5820)) xor (layer5_outputs(5203)));
    layer6_outputs(4389) <= not(layer5_outputs(5758));
    layer6_outputs(4390) <= layer5_outputs(407);
    layer6_outputs(4391) <= layer5_outputs(3637);
    layer6_outputs(4392) <= not(layer5_outputs(6233));
    layer6_outputs(4393) <= layer5_outputs(1979);
    layer6_outputs(4394) <= not((layer5_outputs(4692)) xor (layer5_outputs(7011)));
    layer6_outputs(4395) <= not(layer5_outputs(967));
    layer6_outputs(4396) <= layer5_outputs(2901);
    layer6_outputs(4397) <= layer5_outputs(3571);
    layer6_outputs(4398) <= not((layer5_outputs(2539)) or (layer5_outputs(5390)));
    layer6_outputs(4399) <= layer5_outputs(1048);
    layer6_outputs(4400) <= not((layer5_outputs(1722)) or (layer5_outputs(1961)));
    layer6_outputs(4401) <= not(layer5_outputs(5661)) or (layer5_outputs(4172));
    layer6_outputs(4402) <= layer5_outputs(161);
    layer6_outputs(4403) <= layer5_outputs(2518);
    layer6_outputs(4404) <= not(layer5_outputs(4305));
    layer6_outputs(4405) <= not(layer5_outputs(2274));
    layer6_outputs(4406) <= not((layer5_outputs(853)) xor (layer5_outputs(355)));
    layer6_outputs(4407) <= not(layer5_outputs(5278));
    layer6_outputs(4408) <= layer5_outputs(3113);
    layer6_outputs(4409) <= not((layer5_outputs(6743)) and (layer5_outputs(6897)));
    layer6_outputs(4410) <= (layer5_outputs(1051)) and not (layer5_outputs(7532));
    layer6_outputs(4411) <= not(layer5_outputs(1874));
    layer6_outputs(4412) <= (layer5_outputs(3542)) and not (layer5_outputs(7583));
    layer6_outputs(4413) <= (layer5_outputs(1984)) and not (layer5_outputs(2728));
    layer6_outputs(4414) <= not(layer5_outputs(7558));
    layer6_outputs(4415) <= not(layer5_outputs(5414));
    layer6_outputs(4416) <= not(layer5_outputs(3058));
    layer6_outputs(4417) <= layer5_outputs(186);
    layer6_outputs(4418) <= not(layer5_outputs(3096));
    layer6_outputs(4419) <= layer5_outputs(3094);
    layer6_outputs(4420) <= layer5_outputs(380);
    layer6_outputs(4421) <= not((layer5_outputs(2887)) and (layer5_outputs(1783)));
    layer6_outputs(4422) <= not((layer5_outputs(4785)) and (layer5_outputs(5663)));
    layer6_outputs(4423) <= not(layer5_outputs(1412));
    layer6_outputs(4424) <= not((layer5_outputs(5924)) and (layer5_outputs(4163)));
    layer6_outputs(4425) <= (layer5_outputs(688)) and not (layer5_outputs(5730));
    layer6_outputs(4426) <= (layer5_outputs(4570)) and not (layer5_outputs(7559));
    layer6_outputs(4427) <= layer5_outputs(6242);
    layer6_outputs(4428) <= layer5_outputs(6703);
    layer6_outputs(4429) <= not((layer5_outputs(1795)) and (layer5_outputs(3734)));
    layer6_outputs(4430) <= not(layer5_outputs(5213));
    layer6_outputs(4431) <= not((layer5_outputs(2893)) and (layer5_outputs(1187)));
    layer6_outputs(4432) <= not((layer5_outputs(2853)) xor (layer5_outputs(1344)));
    layer6_outputs(4433) <= not(layer5_outputs(832));
    layer6_outputs(4434) <= layer5_outputs(2196);
    layer6_outputs(4435) <= (layer5_outputs(3208)) or (layer5_outputs(2924));
    layer6_outputs(4436) <= not(layer5_outputs(6441));
    layer6_outputs(4437) <= layer5_outputs(5858);
    layer6_outputs(4438) <= layer5_outputs(4320);
    layer6_outputs(4439) <= layer5_outputs(4488);
    layer6_outputs(4440) <= not((layer5_outputs(7649)) xor (layer5_outputs(1029)));
    layer6_outputs(4441) <= (layer5_outputs(7005)) xor (layer5_outputs(7146));
    layer6_outputs(4442) <= (layer5_outputs(5864)) and (layer5_outputs(1856));
    layer6_outputs(4443) <= layer5_outputs(648);
    layer6_outputs(4444) <= not((layer5_outputs(3859)) xor (layer5_outputs(1275)));
    layer6_outputs(4445) <= not(layer5_outputs(661));
    layer6_outputs(4446) <= layer5_outputs(7232);
    layer6_outputs(4447) <= (layer5_outputs(1319)) and not (layer5_outputs(3625));
    layer6_outputs(4448) <= (layer5_outputs(3961)) and not (layer5_outputs(4504));
    layer6_outputs(4449) <= (layer5_outputs(1704)) and not (layer5_outputs(2606));
    layer6_outputs(4450) <= not(layer5_outputs(3092));
    layer6_outputs(4451) <= not(layer5_outputs(4790));
    layer6_outputs(4452) <= not((layer5_outputs(5946)) xor (layer5_outputs(2071)));
    layer6_outputs(4453) <= not(layer5_outputs(1271));
    layer6_outputs(4454) <= (layer5_outputs(4246)) and not (layer5_outputs(2630));
    layer6_outputs(4455) <= (layer5_outputs(1035)) xor (layer5_outputs(768));
    layer6_outputs(4456) <= not(layer5_outputs(7064));
    layer6_outputs(4457) <= layer5_outputs(6199);
    layer6_outputs(4458) <= (layer5_outputs(4447)) and not (layer5_outputs(2819));
    layer6_outputs(4459) <= layer5_outputs(7654);
    layer6_outputs(4460) <= not((layer5_outputs(3299)) xor (layer5_outputs(6227)));
    layer6_outputs(4461) <= layer5_outputs(7085);
    layer6_outputs(4462) <= not(layer5_outputs(5883));
    layer6_outputs(4463) <= not((layer5_outputs(3618)) xor (layer5_outputs(4981)));
    layer6_outputs(4464) <= not(layer5_outputs(4307));
    layer6_outputs(4465) <= layer5_outputs(6275);
    layer6_outputs(4466) <= not((layer5_outputs(4047)) xor (layer5_outputs(980)));
    layer6_outputs(4467) <= (layer5_outputs(511)) and (layer5_outputs(1655));
    layer6_outputs(4468) <= (layer5_outputs(1050)) xor (layer5_outputs(765));
    layer6_outputs(4469) <= not(layer5_outputs(1513));
    layer6_outputs(4470) <= (layer5_outputs(7376)) and (layer5_outputs(2522));
    layer6_outputs(4471) <= (layer5_outputs(740)) and not (layer5_outputs(1665));
    layer6_outputs(4472) <= layer5_outputs(6651);
    layer6_outputs(4473) <= not(layer5_outputs(6528));
    layer6_outputs(4474) <= (layer5_outputs(353)) and not (layer5_outputs(5941));
    layer6_outputs(4475) <= not(layer5_outputs(6035));
    layer6_outputs(4476) <= layer5_outputs(1007);
    layer6_outputs(4477) <= layer5_outputs(5000);
    layer6_outputs(4478) <= not(layer5_outputs(3313));
    layer6_outputs(4479) <= layer5_outputs(7059);
    layer6_outputs(4480) <= layer5_outputs(2998);
    layer6_outputs(4481) <= (layer5_outputs(2373)) or (layer5_outputs(6465));
    layer6_outputs(4482) <= layer5_outputs(3439);
    layer6_outputs(4483) <= (layer5_outputs(6576)) xor (layer5_outputs(5876));
    layer6_outputs(4484) <= layer5_outputs(2256);
    layer6_outputs(4485) <= layer5_outputs(5829);
    layer6_outputs(4486) <= layer5_outputs(2750);
    layer6_outputs(4487) <= layer5_outputs(847);
    layer6_outputs(4488) <= not(layer5_outputs(996));
    layer6_outputs(4489) <= (layer5_outputs(6029)) xor (layer5_outputs(7554));
    layer6_outputs(4490) <= not(layer5_outputs(1270));
    layer6_outputs(4491) <= (layer5_outputs(3755)) and not (layer5_outputs(482));
    layer6_outputs(4492) <= not(layer5_outputs(4298));
    layer6_outputs(4493) <= (layer5_outputs(5890)) and not (layer5_outputs(7272));
    layer6_outputs(4494) <= layer5_outputs(3480);
    layer6_outputs(4495) <= not(layer5_outputs(3039));
    layer6_outputs(4496) <= layer5_outputs(1079);
    layer6_outputs(4497) <= (layer5_outputs(1922)) and not (layer5_outputs(5437));
    layer6_outputs(4498) <= (layer5_outputs(5477)) and (layer5_outputs(5196));
    layer6_outputs(4499) <= (layer5_outputs(3763)) and not (layer5_outputs(1523));
    layer6_outputs(4500) <= (layer5_outputs(347)) xor (layer5_outputs(4961));
    layer6_outputs(4501) <= (layer5_outputs(5547)) xor (layer5_outputs(5052));
    layer6_outputs(4502) <= not(layer5_outputs(5292));
    layer6_outputs(4503) <= not((layer5_outputs(181)) and (layer5_outputs(4579)));
    layer6_outputs(4504) <= not(layer5_outputs(1578)) or (layer5_outputs(3552));
    layer6_outputs(4505) <= layer5_outputs(2132);
    layer6_outputs(4506) <= layer5_outputs(3559);
    layer6_outputs(4507) <= not((layer5_outputs(172)) or (layer5_outputs(837)));
    layer6_outputs(4508) <= not(layer5_outputs(4048)) or (layer5_outputs(540));
    layer6_outputs(4509) <= not(layer5_outputs(7562));
    layer6_outputs(4510) <= (layer5_outputs(5389)) xor (layer5_outputs(5016));
    layer6_outputs(4511) <= (layer5_outputs(6264)) and not (layer5_outputs(5235));
    layer6_outputs(4512) <= not(layer5_outputs(4448));
    layer6_outputs(4513) <= (layer5_outputs(2898)) xor (layer5_outputs(4910));
    layer6_outputs(4514) <= not((layer5_outputs(555)) or (layer5_outputs(1479)));
    layer6_outputs(4515) <= (layer5_outputs(7156)) xor (layer5_outputs(3022));
    layer6_outputs(4516) <= not(layer5_outputs(1154));
    layer6_outputs(4517) <= not(layer5_outputs(2046));
    layer6_outputs(4518) <= (layer5_outputs(5928)) or (layer5_outputs(5740));
    layer6_outputs(4519) <= not(layer5_outputs(774));
    layer6_outputs(4520) <= layer5_outputs(3365);
    layer6_outputs(4521) <= not((layer5_outputs(1501)) xor (layer5_outputs(3705)));
    layer6_outputs(4522) <= not(layer5_outputs(2846));
    layer6_outputs(4523) <= not((layer5_outputs(2102)) or (layer5_outputs(5178)));
    layer6_outputs(4524) <= not(layer5_outputs(2738));
    layer6_outputs(4525) <= layer5_outputs(5410);
    layer6_outputs(4526) <= not(layer5_outputs(5917));
    layer6_outputs(4527) <= (layer5_outputs(4793)) or (layer5_outputs(3178));
    layer6_outputs(4528) <= (layer5_outputs(6118)) and not (layer5_outputs(2549));
    layer6_outputs(4529) <= not(layer5_outputs(5625));
    layer6_outputs(4530) <= not(layer5_outputs(4002));
    layer6_outputs(4531) <= (layer5_outputs(4549)) xor (layer5_outputs(459));
    layer6_outputs(4532) <= not(layer5_outputs(6859));
    layer6_outputs(4533) <= not((layer5_outputs(3011)) xor (layer5_outputs(4016)));
    layer6_outputs(4534) <= not(layer5_outputs(2374));
    layer6_outputs(4535) <= layer5_outputs(4492);
    layer6_outputs(4536) <= layer5_outputs(593);
    layer6_outputs(4537) <= (layer5_outputs(6568)) and not (layer5_outputs(6480));
    layer6_outputs(4538) <= (layer5_outputs(5145)) and not (layer5_outputs(3708));
    layer6_outputs(4539) <= (layer5_outputs(5558)) xor (layer5_outputs(5066));
    layer6_outputs(4540) <= (layer5_outputs(157)) and not (layer5_outputs(3265));
    layer6_outputs(4541) <= not(layer5_outputs(5121));
    layer6_outputs(4542) <= layer5_outputs(3757);
    layer6_outputs(4543) <= (layer5_outputs(80)) and not (layer5_outputs(4413));
    layer6_outputs(4544) <= not(layer5_outputs(1908));
    layer6_outputs(4545) <= not(layer5_outputs(7572)) or (layer5_outputs(4869));
    layer6_outputs(4546) <= not(layer5_outputs(6777));
    layer6_outputs(4547) <= not(layer5_outputs(367));
    layer6_outputs(4548) <= not((layer5_outputs(2529)) xor (layer5_outputs(103)));
    layer6_outputs(4549) <= not(layer5_outputs(741));
    layer6_outputs(4550) <= layer5_outputs(6283);
    layer6_outputs(4551) <= not(layer5_outputs(5679));
    layer6_outputs(4552) <= not(layer5_outputs(4196));
    layer6_outputs(4553) <= not(layer5_outputs(2499));
    layer6_outputs(4554) <= not((layer5_outputs(623)) xor (layer5_outputs(71)));
    layer6_outputs(4555) <= not((layer5_outputs(4647)) and (layer5_outputs(4747)));
    layer6_outputs(4556) <= not((layer5_outputs(1978)) or (layer5_outputs(4629)));
    layer6_outputs(4557) <= not(layer5_outputs(3285));
    layer6_outputs(4558) <= (layer5_outputs(2860)) or (layer5_outputs(2294));
    layer6_outputs(4559) <= (layer5_outputs(985)) xor (layer5_outputs(2646));
    layer6_outputs(4560) <= layer5_outputs(1484);
    layer6_outputs(4561) <= layer5_outputs(1975);
    layer6_outputs(4562) <= not((layer5_outputs(1201)) xor (layer5_outputs(5285)));
    layer6_outputs(4563) <= not(layer5_outputs(3546)) or (layer5_outputs(2968));
    layer6_outputs(4564) <= layer5_outputs(4475);
    layer6_outputs(4565) <= (layer5_outputs(4633)) xor (layer5_outputs(1579));
    layer6_outputs(4566) <= not(layer5_outputs(5068));
    layer6_outputs(4567) <= layer5_outputs(2403);
    layer6_outputs(4568) <= not(layer5_outputs(3594));
    layer6_outputs(4569) <= not((layer5_outputs(7170)) or (layer5_outputs(1078)));
    layer6_outputs(4570) <= layer5_outputs(7039);
    layer6_outputs(4571) <= not(layer5_outputs(862));
    layer6_outputs(4572) <= not(layer5_outputs(3300));
    layer6_outputs(4573) <= (layer5_outputs(665)) and not (layer5_outputs(2504));
    layer6_outputs(4574) <= not((layer5_outputs(4284)) xor (layer5_outputs(6857)));
    layer6_outputs(4575) <= not((layer5_outputs(3558)) and (layer5_outputs(5149)));
    layer6_outputs(4576) <= not(layer5_outputs(5460)) or (layer5_outputs(4709));
    layer6_outputs(4577) <= (layer5_outputs(7485)) and not (layer5_outputs(1982));
    layer6_outputs(4578) <= (layer5_outputs(6195)) xor (layer5_outputs(1320));
    layer6_outputs(4579) <= (layer5_outputs(582)) and not (layer5_outputs(1331));
    layer6_outputs(4580) <= not(layer5_outputs(6074)) or (layer5_outputs(3660));
    layer6_outputs(4581) <= not((layer5_outputs(6136)) and (layer5_outputs(3006)));
    layer6_outputs(4582) <= (layer5_outputs(1714)) xor (layer5_outputs(3641));
    layer6_outputs(4583) <= not(layer5_outputs(2591)) or (layer5_outputs(2931));
    layer6_outputs(4584) <= not(layer5_outputs(4748));
    layer6_outputs(4585) <= layer5_outputs(5461);
    layer6_outputs(4586) <= not((layer5_outputs(430)) xor (layer5_outputs(4715)));
    layer6_outputs(4587) <= layer5_outputs(716);
    layer6_outputs(4588) <= not(layer5_outputs(2946)) or (layer5_outputs(5220));
    layer6_outputs(4589) <= not((layer5_outputs(1089)) xor (layer5_outputs(7280)));
    layer6_outputs(4590) <= not(layer5_outputs(7548));
    layer6_outputs(4591) <= (layer5_outputs(881)) xor (layer5_outputs(761));
    layer6_outputs(4592) <= layer5_outputs(2218);
    layer6_outputs(4593) <= not(layer5_outputs(4756));
    layer6_outputs(4594) <= layer5_outputs(6353);
    layer6_outputs(4595) <= not((layer5_outputs(19)) xor (layer5_outputs(1405)));
    layer6_outputs(4596) <= (layer5_outputs(5362)) xor (layer5_outputs(951));
    layer6_outputs(4597) <= layer5_outputs(2911);
    layer6_outputs(4598) <= not(layer5_outputs(4113));
    layer6_outputs(4599) <= not(layer5_outputs(5428)) or (layer5_outputs(4857));
    layer6_outputs(4600) <= (layer5_outputs(7472)) and not (layer5_outputs(690));
    layer6_outputs(4601) <= (layer5_outputs(5153)) or (layer5_outputs(6273));
    layer6_outputs(4602) <= (layer5_outputs(6858)) and (layer5_outputs(5939));
    layer6_outputs(4603) <= (layer5_outputs(4132)) xor (layer5_outputs(3935));
    layer6_outputs(4604) <= not(layer5_outputs(7302));
    layer6_outputs(4605) <= not(layer5_outputs(5692)) or (layer5_outputs(3029));
    layer6_outputs(4606) <= (layer5_outputs(1312)) xor (layer5_outputs(3125));
    layer6_outputs(4607) <= not(layer5_outputs(590));
    layer6_outputs(4608) <= not(layer5_outputs(6374));
    layer6_outputs(4609) <= not((layer5_outputs(2122)) xor (layer5_outputs(1943)));
    layer6_outputs(4610) <= (layer5_outputs(1001)) xor (layer5_outputs(5606));
    layer6_outputs(4611) <= layer5_outputs(2605);
    layer6_outputs(4612) <= layer5_outputs(1444);
    layer6_outputs(4613) <= not((layer5_outputs(4809)) and (layer5_outputs(2241)));
    layer6_outputs(4614) <= not(layer5_outputs(7179));
    layer6_outputs(4615) <= (layer5_outputs(4764)) and (layer5_outputs(4696));
    layer6_outputs(4616) <= not(layer5_outputs(513));
    layer6_outputs(4617) <= not(layer5_outputs(2354));
    layer6_outputs(4618) <= layer5_outputs(2214);
    layer6_outputs(4619) <= layer5_outputs(2672);
    layer6_outputs(4620) <= not(layer5_outputs(628)) or (layer5_outputs(1215));
    layer6_outputs(4621) <= not((layer5_outputs(6792)) xor (layer5_outputs(5934)));
    layer6_outputs(4622) <= (layer5_outputs(4376)) xor (layer5_outputs(2903));
    layer6_outputs(4623) <= layer5_outputs(205);
    layer6_outputs(4624) <= (layer5_outputs(730)) xor (layer5_outputs(6252));
    layer6_outputs(4625) <= (layer5_outputs(7409)) or (layer5_outputs(3615));
    layer6_outputs(4626) <= layer5_outputs(5165);
    layer6_outputs(4627) <= (layer5_outputs(5030)) xor (layer5_outputs(6166));
    layer6_outputs(4628) <= (layer5_outputs(6241)) xor (layer5_outputs(1399));
    layer6_outputs(4629) <= (layer5_outputs(1128)) xor (layer5_outputs(2513));
    layer6_outputs(4630) <= (layer5_outputs(168)) xor (layer5_outputs(2712));
    layer6_outputs(4631) <= not(layer5_outputs(6652)) or (layer5_outputs(743));
    layer6_outputs(4632) <= layer5_outputs(5471);
    layer6_outputs(4633) <= (layer5_outputs(804)) and not (layer5_outputs(6855));
    layer6_outputs(4634) <= layer5_outputs(3739);
    layer6_outputs(4635) <= not((layer5_outputs(7605)) and (layer5_outputs(5845)));
    layer6_outputs(4636) <= not(layer5_outputs(5894)) or (layer5_outputs(5260));
    layer6_outputs(4637) <= not(layer5_outputs(1758)) or (layer5_outputs(3198));
    layer6_outputs(4638) <= not((layer5_outputs(3022)) xor (layer5_outputs(3389)));
    layer6_outputs(4639) <= not((layer5_outputs(7248)) and (layer5_outputs(6108)));
    layer6_outputs(4640) <= not(layer5_outputs(1586));
    layer6_outputs(4641) <= not((layer5_outputs(5763)) xor (layer5_outputs(5910)));
    layer6_outputs(4642) <= '0';
    layer6_outputs(4643) <= not((layer5_outputs(3454)) and (layer5_outputs(1306)));
    layer6_outputs(4644) <= layer5_outputs(2467);
    layer6_outputs(4645) <= layer5_outputs(5240);
    layer6_outputs(4646) <= (layer5_outputs(7160)) and not (layer5_outputs(4367));
    layer6_outputs(4647) <= not(layer5_outputs(7527));
    layer6_outputs(4648) <= not((layer5_outputs(7239)) xor (layer5_outputs(4018)));
    layer6_outputs(4649) <= (layer5_outputs(391)) xor (layer5_outputs(1111));
    layer6_outputs(4650) <= (layer5_outputs(2740)) xor (layer5_outputs(5850));
    layer6_outputs(4651) <= not((layer5_outputs(3451)) xor (layer5_outputs(5454)));
    layer6_outputs(4652) <= not(layer5_outputs(2251));
    layer6_outputs(4653) <= not(layer5_outputs(5519));
    layer6_outputs(4654) <= layer5_outputs(1548);
    layer6_outputs(4655) <= not(layer5_outputs(2884));
    layer6_outputs(4656) <= layer5_outputs(3406);
    layer6_outputs(4657) <= not(layer5_outputs(3388)) or (layer5_outputs(7002));
    layer6_outputs(4658) <= not(layer5_outputs(1538));
    layer6_outputs(4659) <= layer5_outputs(4492);
    layer6_outputs(4660) <= layer5_outputs(3242);
    layer6_outputs(4661) <= not(layer5_outputs(6816));
    layer6_outputs(4662) <= layer5_outputs(5721);
    layer6_outputs(4663) <= not((layer5_outputs(6742)) xor (layer5_outputs(694)));
    layer6_outputs(4664) <= layer5_outputs(6872);
    layer6_outputs(4665) <= layer5_outputs(7522);
    layer6_outputs(4666) <= layer5_outputs(272);
    layer6_outputs(4667) <= not(layer5_outputs(5441)) or (layer5_outputs(3457));
    layer6_outputs(4668) <= (layer5_outputs(701)) and not (layer5_outputs(6058));
    layer6_outputs(4669) <= layer5_outputs(2172);
    layer6_outputs(4670) <= layer5_outputs(76);
    layer6_outputs(4671) <= not((layer5_outputs(4567)) xor (layer5_outputs(4091)));
    layer6_outputs(4672) <= (layer5_outputs(2001)) and not (layer5_outputs(6221));
    layer6_outputs(4673) <= not(layer5_outputs(962)) or (layer5_outputs(4105));
    layer6_outputs(4674) <= (layer5_outputs(6962)) and not (layer5_outputs(2895));
    layer6_outputs(4675) <= (layer5_outputs(489)) and not (layer5_outputs(4054));
    layer6_outputs(4676) <= layer5_outputs(6428);
    layer6_outputs(4677) <= (layer5_outputs(153)) and (layer5_outputs(3070));
    layer6_outputs(4678) <= (layer5_outputs(2144)) xor (layer5_outputs(2597));
    layer6_outputs(4679) <= not(layer5_outputs(4154));
    layer6_outputs(4680) <= layer5_outputs(6416);
    layer6_outputs(4681) <= not(layer5_outputs(7640));
    layer6_outputs(4682) <= layer5_outputs(6190);
    layer6_outputs(4683) <= (layer5_outputs(3305)) and not (layer5_outputs(1481));
    layer6_outputs(4684) <= not(layer5_outputs(4215));
    layer6_outputs(4685) <= layer5_outputs(645);
    layer6_outputs(4686) <= not((layer5_outputs(4787)) and (layer5_outputs(3670)));
    layer6_outputs(4687) <= not(layer5_outputs(1199));
    layer6_outputs(4688) <= '0';
    layer6_outputs(4689) <= not(layer5_outputs(3024));
    layer6_outputs(4690) <= not((layer5_outputs(7534)) and (layer5_outputs(7339)));
    layer6_outputs(4691) <= not(layer5_outputs(6232));
    layer6_outputs(4692) <= layer5_outputs(6146);
    layer6_outputs(4693) <= layer5_outputs(5556);
    layer6_outputs(4694) <= layer5_outputs(5107);
    layer6_outputs(4695) <= not(layer5_outputs(5322)) or (layer5_outputs(651));
    layer6_outputs(4696) <= not(layer5_outputs(6797));
    layer6_outputs(4697) <= (layer5_outputs(551)) xor (layer5_outputs(7007));
    layer6_outputs(4698) <= (layer5_outputs(4083)) xor (layer5_outputs(5218));
    layer6_outputs(4699) <= not(layer5_outputs(6158)) or (layer5_outputs(4746));
    layer6_outputs(4700) <= not(layer5_outputs(7616));
    layer6_outputs(4701) <= (layer5_outputs(7220)) xor (layer5_outputs(3438));
    layer6_outputs(4702) <= layer5_outputs(4488);
    layer6_outputs(4703) <= not(layer5_outputs(4720)) or (layer5_outputs(6254));
    layer6_outputs(4704) <= not((layer5_outputs(6785)) and (layer5_outputs(1165)));
    layer6_outputs(4705) <= layer5_outputs(2888);
    layer6_outputs(4706) <= not((layer5_outputs(6584)) xor (layer5_outputs(3977)));
    layer6_outputs(4707) <= not(layer5_outputs(3424));
    layer6_outputs(4708) <= (layer5_outputs(1886)) and (layer5_outputs(5759));
    layer6_outputs(4709) <= not(layer5_outputs(4496));
    layer6_outputs(4710) <= not(layer5_outputs(6437));
    layer6_outputs(4711) <= layer5_outputs(332);
    layer6_outputs(4712) <= not(layer5_outputs(6930));
    layer6_outputs(4713) <= (layer5_outputs(1633)) xor (layer5_outputs(3259));
    layer6_outputs(4714) <= not(layer5_outputs(7600)) or (layer5_outputs(1464));
    layer6_outputs(4715) <= not(layer5_outputs(5289));
    layer6_outputs(4716) <= layer5_outputs(6689);
    layer6_outputs(4717) <= (layer5_outputs(461)) or (layer5_outputs(7663));
    layer6_outputs(4718) <= (layer5_outputs(3435)) or (layer5_outputs(1172));
    layer6_outputs(4719) <= not(layer5_outputs(7333));
    layer6_outputs(4720) <= layer5_outputs(1510);
    layer6_outputs(4721) <= (layer5_outputs(950)) xor (layer5_outputs(2435));
    layer6_outputs(4722) <= '1';
    layer6_outputs(4723) <= layer5_outputs(4074);
    layer6_outputs(4724) <= layer5_outputs(6746);
    layer6_outputs(4725) <= not((layer5_outputs(822)) and (layer5_outputs(3513)));
    layer6_outputs(4726) <= not(layer5_outputs(7014));
    layer6_outputs(4727) <= layer5_outputs(6457);
    layer6_outputs(4728) <= layer5_outputs(2395);
    layer6_outputs(4729) <= not(layer5_outputs(1590)) or (layer5_outputs(4217));
    layer6_outputs(4730) <= not((layer5_outputs(3505)) or (layer5_outputs(4772)));
    layer6_outputs(4731) <= layer5_outputs(5311);
    layer6_outputs(4732) <= not((layer5_outputs(5303)) and (layer5_outputs(1963)));
    layer6_outputs(4733) <= not((layer5_outputs(2658)) xor (layer5_outputs(2191)));
    layer6_outputs(4734) <= layer5_outputs(4286);
    layer6_outputs(4735) <= (layer5_outputs(1482)) or (layer5_outputs(4269));
    layer6_outputs(4736) <= not((layer5_outputs(6735)) xor (layer5_outputs(7340)));
    layer6_outputs(4737) <= not(layer5_outputs(6211));
    layer6_outputs(4738) <= layer5_outputs(7325);
    layer6_outputs(4739) <= layer5_outputs(5777);
    layer6_outputs(4740) <= not(layer5_outputs(2995));
    layer6_outputs(4741) <= (layer5_outputs(4645)) xor (layer5_outputs(2075));
    layer6_outputs(4742) <= (layer5_outputs(5798)) and (layer5_outputs(7674));
    layer6_outputs(4743) <= layer5_outputs(871);
    layer6_outputs(4744) <= not(layer5_outputs(4947));
    layer6_outputs(4745) <= not((layer5_outputs(6784)) xor (layer5_outputs(3081)));
    layer6_outputs(4746) <= not((layer5_outputs(4179)) or (layer5_outputs(5722)));
    layer6_outputs(4747) <= not(layer5_outputs(915));
    layer6_outputs(4748) <= layer5_outputs(4907);
    layer6_outputs(4749) <= (layer5_outputs(6797)) or (layer5_outputs(4310));
    layer6_outputs(4750) <= not(layer5_outputs(4366));
    layer6_outputs(4751) <= not(layer5_outputs(5806)) or (layer5_outputs(1447));
    layer6_outputs(4752) <= layer5_outputs(620);
    layer6_outputs(4753) <= not(layer5_outputs(6355));
    layer6_outputs(4754) <= not(layer5_outputs(2324));
    layer6_outputs(4755) <= layer5_outputs(6353);
    layer6_outputs(4756) <= (layer5_outputs(463)) and (layer5_outputs(6240));
    layer6_outputs(4757) <= not(layer5_outputs(206));
    layer6_outputs(4758) <= not((layer5_outputs(3124)) or (layer5_outputs(2214)));
    layer6_outputs(4759) <= layer5_outputs(3026);
    layer6_outputs(4760) <= not(layer5_outputs(2654));
    layer6_outputs(4761) <= not((layer5_outputs(5956)) xor (layer5_outputs(5826)));
    layer6_outputs(4762) <= (layer5_outputs(5695)) xor (layer5_outputs(3619));
    layer6_outputs(4763) <= not((layer5_outputs(6305)) xor (layer5_outputs(5290)));
    layer6_outputs(4764) <= not(layer5_outputs(3604));
    layer6_outputs(4765) <= layer5_outputs(6198);
    layer6_outputs(4766) <= layer5_outputs(4838);
    layer6_outputs(4767) <= layer5_outputs(6710);
    layer6_outputs(4768) <= not((layer5_outputs(640)) and (layer5_outputs(7073)));
    layer6_outputs(4769) <= not(layer5_outputs(2994));
    layer6_outputs(4770) <= layer5_outputs(6339);
    layer6_outputs(4771) <= layer5_outputs(4191);
    layer6_outputs(4772) <= not(layer5_outputs(6507));
    layer6_outputs(4773) <= (layer5_outputs(209)) and not (layer5_outputs(745));
    layer6_outputs(4774) <= not((layer5_outputs(978)) xor (layer5_outputs(6972)));
    layer6_outputs(4775) <= (layer5_outputs(6529)) xor (layer5_outputs(3753));
    layer6_outputs(4776) <= (layer5_outputs(2029)) and (layer5_outputs(3210));
    layer6_outputs(4777) <= not(layer5_outputs(6425)) or (layer5_outputs(5031));
    layer6_outputs(4778) <= not((layer5_outputs(5570)) xor (layer5_outputs(1580)));
    layer6_outputs(4779) <= not(layer5_outputs(5026));
    layer6_outputs(4780) <= not(layer5_outputs(6245));
    layer6_outputs(4781) <= not(layer5_outputs(2542));
    layer6_outputs(4782) <= not((layer5_outputs(6766)) xor (layer5_outputs(2467)));
    layer6_outputs(4783) <= layer5_outputs(2301);
    layer6_outputs(4784) <= not(layer5_outputs(6309));
    layer6_outputs(4785) <= layer5_outputs(5890);
    layer6_outputs(4786) <= not(layer5_outputs(7677));
    layer6_outputs(4787) <= layer5_outputs(5671);
    layer6_outputs(4788) <= not(layer5_outputs(3065));
    layer6_outputs(4789) <= layer5_outputs(2071);
    layer6_outputs(4790) <= (layer5_outputs(4671)) and not (layer5_outputs(7034));
    layer6_outputs(4791) <= not(layer5_outputs(930));
    layer6_outputs(4792) <= not((layer5_outputs(6301)) and (layer5_outputs(2916)));
    layer6_outputs(4793) <= (layer5_outputs(5686)) or (layer5_outputs(1919));
    layer6_outputs(4794) <= (layer5_outputs(4643)) and not (layer5_outputs(2820));
    layer6_outputs(4795) <= layer5_outputs(4031);
    layer6_outputs(4796) <= not((layer5_outputs(4124)) xor (layer5_outputs(6483)));
    layer6_outputs(4797) <= (layer5_outputs(6695)) or (layer5_outputs(771));
    layer6_outputs(4798) <= not(layer5_outputs(3808));
    layer6_outputs(4799) <= (layer5_outputs(3080)) and not (layer5_outputs(4901));
    layer6_outputs(4800) <= not((layer5_outputs(2349)) xor (layer5_outputs(7551)));
    layer6_outputs(4801) <= (layer5_outputs(3741)) or (layer5_outputs(5171));
    layer6_outputs(4802) <= (layer5_outputs(7567)) and (layer5_outputs(2874));
    layer6_outputs(4803) <= not(layer5_outputs(4317));
    layer6_outputs(4804) <= not((layer5_outputs(3734)) xor (layer5_outputs(1658)));
    layer6_outputs(4805) <= not((layer5_outputs(797)) or (layer5_outputs(5638)));
    layer6_outputs(4806) <= layer5_outputs(2447);
    layer6_outputs(4807) <= (layer5_outputs(2961)) and not (layer5_outputs(6684));
    layer6_outputs(4808) <= layer5_outputs(6671);
    layer6_outputs(4809) <= layer5_outputs(6774);
    layer6_outputs(4810) <= (layer5_outputs(1557)) and not (layer5_outputs(7321));
    layer6_outputs(4811) <= not(layer5_outputs(3176));
    layer6_outputs(4812) <= not(layer5_outputs(4152)) or (layer5_outputs(234));
    layer6_outputs(4813) <= layer5_outputs(3195);
    layer6_outputs(4814) <= not(layer5_outputs(661));
    layer6_outputs(4815) <= not(layer5_outputs(2332)) or (layer5_outputs(4741));
    layer6_outputs(4816) <= not((layer5_outputs(101)) xor (layer5_outputs(3526)));
    layer6_outputs(4817) <= not(layer5_outputs(3319));
    layer6_outputs(4818) <= layer5_outputs(6974);
    layer6_outputs(4819) <= not((layer5_outputs(3719)) xor (layer5_outputs(6914)));
    layer6_outputs(4820) <= (layer5_outputs(1843)) and not (layer5_outputs(951));
    layer6_outputs(4821) <= not(layer5_outputs(5635));
    layer6_outputs(4822) <= layer5_outputs(6319);
    layer6_outputs(4823) <= not(layer5_outputs(6271));
    layer6_outputs(4824) <= not(layer5_outputs(1068));
    layer6_outputs(4825) <= (layer5_outputs(6558)) and (layer5_outputs(7608));
    layer6_outputs(4826) <= not(layer5_outputs(5843)) or (layer5_outputs(683));
    layer6_outputs(4827) <= layer5_outputs(4090);
    layer6_outputs(4828) <= not(layer5_outputs(1276));
    layer6_outputs(4829) <= not(layer5_outputs(2811));
    layer6_outputs(4830) <= not(layer5_outputs(317));
    layer6_outputs(4831) <= (layer5_outputs(3192)) xor (layer5_outputs(4541));
    layer6_outputs(4832) <= (layer5_outputs(6151)) or (layer5_outputs(792));
    layer6_outputs(4833) <= layer5_outputs(1067);
    layer6_outputs(4834) <= not((layer5_outputs(6278)) xor (layer5_outputs(4948)));
    layer6_outputs(4835) <= layer5_outputs(7357);
    layer6_outputs(4836) <= layer5_outputs(5939);
    layer6_outputs(4837) <= not(layer5_outputs(2531));
    layer6_outputs(4838) <= not(layer5_outputs(1506)) or (layer5_outputs(146));
    layer6_outputs(4839) <= (layer5_outputs(4051)) or (layer5_outputs(3416));
    layer6_outputs(4840) <= layer5_outputs(6704);
    layer6_outputs(4841) <= layer5_outputs(5233);
    layer6_outputs(4842) <= not((layer5_outputs(304)) xor (layer5_outputs(502)));
    layer6_outputs(4843) <= not((layer5_outputs(6397)) xor (layer5_outputs(2383)));
    layer6_outputs(4844) <= (layer5_outputs(4972)) xor (layer5_outputs(2100));
    layer6_outputs(4845) <= (layer5_outputs(1791)) and (layer5_outputs(4517));
    layer6_outputs(4846) <= layer5_outputs(4352);
    layer6_outputs(4847) <= not(layer5_outputs(2050));
    layer6_outputs(4848) <= not((layer5_outputs(1222)) xor (layer5_outputs(4411)));
    layer6_outputs(4849) <= not(layer5_outputs(844));
    layer6_outputs(4850) <= not(layer5_outputs(1741)) or (layer5_outputs(140));
    layer6_outputs(4851) <= not(layer5_outputs(3540)) or (layer5_outputs(2380));
    layer6_outputs(4852) <= layer5_outputs(6805);
    layer6_outputs(4853) <= (layer5_outputs(413)) xor (layer5_outputs(5969));
    layer6_outputs(4854) <= layer5_outputs(4375);
    layer6_outputs(4855) <= (layer5_outputs(3968)) or (layer5_outputs(3267));
    layer6_outputs(4856) <= layer5_outputs(2547);
    layer6_outputs(4857) <= not(layer5_outputs(874));
    layer6_outputs(4858) <= layer5_outputs(560);
    layer6_outputs(4859) <= not(layer5_outputs(1494));
    layer6_outputs(4860) <= (layer5_outputs(3001)) and not (layer5_outputs(3326));
    layer6_outputs(4861) <= (layer5_outputs(5491)) and not (layer5_outputs(2600));
    layer6_outputs(4862) <= layer5_outputs(120);
    layer6_outputs(4863) <= (layer5_outputs(1507)) and not (layer5_outputs(2766));
    layer6_outputs(4864) <= (layer5_outputs(4448)) and not (layer5_outputs(6995));
    layer6_outputs(4865) <= not(layer5_outputs(2519));
    layer6_outputs(4866) <= (layer5_outputs(3450)) and (layer5_outputs(1077));
    layer6_outputs(4867) <= not(layer5_outputs(6155));
    layer6_outputs(4868) <= not(layer5_outputs(5779)) or (layer5_outputs(3766));
    layer6_outputs(4869) <= not((layer5_outputs(7593)) or (layer5_outputs(5463)));
    layer6_outputs(4870) <= not(layer5_outputs(6718));
    layer6_outputs(4871) <= layer5_outputs(1378);
    layer6_outputs(4872) <= not(layer5_outputs(6471));
    layer6_outputs(4873) <= (layer5_outputs(1767)) or (layer5_outputs(2843));
    layer6_outputs(4874) <= not(layer5_outputs(2137));
    layer6_outputs(4875) <= not(layer5_outputs(2802));
    layer6_outputs(4876) <= layer5_outputs(336);
    layer6_outputs(4877) <= (layer5_outputs(6540)) xor (layer5_outputs(807));
    layer6_outputs(4878) <= (layer5_outputs(7520)) xor (layer5_outputs(5231));
    layer6_outputs(4879) <= '1';
    layer6_outputs(4880) <= layer5_outputs(1986);
    layer6_outputs(4881) <= not(layer5_outputs(4189));
    layer6_outputs(4882) <= not(layer5_outputs(1467));
    layer6_outputs(4883) <= (layer5_outputs(2022)) and not (layer5_outputs(5732));
    layer6_outputs(4884) <= (layer5_outputs(6948)) or (layer5_outputs(1175));
    layer6_outputs(4885) <= layer5_outputs(7388);
    layer6_outputs(4886) <= not(layer5_outputs(4850));
    layer6_outputs(4887) <= layer5_outputs(5493);
    layer6_outputs(4888) <= (layer5_outputs(189)) and not (layer5_outputs(5556));
    layer6_outputs(4889) <= not(layer5_outputs(4095));
    layer6_outputs(4890) <= layer5_outputs(3355);
    layer6_outputs(4891) <= not(layer5_outputs(3371));
    layer6_outputs(4892) <= not(layer5_outputs(7106)) or (layer5_outputs(2741));
    layer6_outputs(4893) <= (layer5_outputs(3138)) xor (layer5_outputs(1250));
    layer6_outputs(4894) <= layer5_outputs(5825);
    layer6_outputs(4895) <= (layer5_outputs(3071)) or (layer5_outputs(1881));
    layer6_outputs(4896) <= not((layer5_outputs(5994)) xor (layer5_outputs(270)));
    layer6_outputs(4897) <= not(layer5_outputs(7278));
    layer6_outputs(4898) <= layer5_outputs(6619);
    layer6_outputs(4899) <= layer5_outputs(2997);
    layer6_outputs(4900) <= not(layer5_outputs(6565));
    layer6_outputs(4901) <= not(layer5_outputs(5726)) or (layer5_outputs(5603));
    layer6_outputs(4902) <= not(layer5_outputs(3112));
    layer6_outputs(4903) <= not(layer5_outputs(5164));
    layer6_outputs(4904) <= not(layer5_outputs(4982));
    layer6_outputs(4905) <= (layer5_outputs(591)) and (layer5_outputs(1407));
    layer6_outputs(4906) <= layer5_outputs(764);
    layer6_outputs(4907) <= (layer5_outputs(233)) and not (layer5_outputs(4300));
    layer6_outputs(4908) <= not(layer5_outputs(4804));
    layer6_outputs(4909) <= not((layer5_outputs(7188)) xor (layer5_outputs(6477)));
    layer6_outputs(4910) <= not((layer5_outputs(4147)) xor (layer5_outputs(3779)));
    layer6_outputs(4911) <= not(layer5_outputs(4483));
    layer6_outputs(4912) <= (layer5_outputs(2857)) or (layer5_outputs(3975));
    layer6_outputs(4913) <= layer5_outputs(948);
    layer6_outputs(4914) <= (layer5_outputs(698)) xor (layer5_outputs(3487));
    layer6_outputs(4915) <= not(layer5_outputs(2390));
    layer6_outputs(4916) <= (layer5_outputs(5857)) and not (layer5_outputs(4008));
    layer6_outputs(4917) <= (layer5_outputs(1183)) xor (layer5_outputs(7586));
    layer6_outputs(4918) <= not(layer5_outputs(5799));
    layer6_outputs(4919) <= layer5_outputs(7438);
    layer6_outputs(4920) <= layer5_outputs(4393);
    layer6_outputs(4921) <= layer5_outputs(4748);
    layer6_outputs(4922) <= (layer5_outputs(5601)) and (layer5_outputs(2621));
    layer6_outputs(4923) <= not(layer5_outputs(7503));
    layer6_outputs(4924) <= layer5_outputs(3023);
    layer6_outputs(4925) <= not((layer5_outputs(3907)) and (layer5_outputs(5421)));
    layer6_outputs(4926) <= (layer5_outputs(1898)) or (layer5_outputs(2398));
    layer6_outputs(4927) <= (layer5_outputs(7587)) or (layer5_outputs(1032));
    layer6_outputs(4928) <= layer5_outputs(3317);
    layer6_outputs(4929) <= not((layer5_outputs(323)) xor (layer5_outputs(5336)));
    layer6_outputs(4930) <= not(layer5_outputs(6065));
    layer6_outputs(4931) <= not(layer5_outputs(5652));
    layer6_outputs(4932) <= not((layer5_outputs(519)) or (layer5_outputs(2441)));
    layer6_outputs(4933) <= not((layer5_outputs(912)) or (layer5_outputs(1022)));
    layer6_outputs(4934) <= not((layer5_outputs(6044)) or (layer5_outputs(4998)));
    layer6_outputs(4935) <= layer5_outputs(45);
    layer6_outputs(4936) <= (layer5_outputs(7205)) and not (layer5_outputs(2019));
    layer6_outputs(4937) <= not(layer5_outputs(2134));
    layer6_outputs(4938) <= not(layer5_outputs(7488));
    layer6_outputs(4939) <= not((layer5_outputs(5115)) or (layer5_outputs(3798)));
    layer6_outputs(4940) <= (layer5_outputs(3581)) xor (layer5_outputs(7598));
    layer6_outputs(4941) <= layer5_outputs(3021);
    layer6_outputs(4942) <= (layer5_outputs(1109)) xor (layer5_outputs(4118));
    layer6_outputs(4943) <= layer5_outputs(78);
    layer6_outputs(4944) <= not(layer5_outputs(5610));
    layer6_outputs(4945) <= not(layer5_outputs(5234));
    layer6_outputs(4946) <= not((layer5_outputs(4957)) and (layer5_outputs(4864)));
    layer6_outputs(4947) <= not(layer5_outputs(565));
    layer6_outputs(4948) <= not((layer5_outputs(2803)) xor (layer5_outputs(6485)));
    layer6_outputs(4949) <= (layer5_outputs(2929)) and (layer5_outputs(916));
    layer6_outputs(4950) <= (layer5_outputs(2662)) or (layer5_outputs(5202));
    layer6_outputs(4951) <= not((layer5_outputs(6890)) xor (layer5_outputs(4381)));
    layer6_outputs(4952) <= layer5_outputs(714);
    layer6_outputs(4953) <= layer5_outputs(7425);
    layer6_outputs(4954) <= not((layer5_outputs(3362)) xor (layer5_outputs(7665)));
    layer6_outputs(4955) <= layer5_outputs(6968);
    layer6_outputs(4956) <= not(layer5_outputs(570)) or (layer5_outputs(7289));
    layer6_outputs(4957) <= not(layer5_outputs(2362));
    layer6_outputs(4958) <= layer5_outputs(7131);
    layer6_outputs(4959) <= (layer5_outputs(3910)) xor (layer5_outputs(1085));
    layer6_outputs(4960) <= not((layer5_outputs(3818)) xor (layer5_outputs(2125)));
    layer6_outputs(4961) <= not(layer5_outputs(5634));
    layer6_outputs(4962) <= (layer5_outputs(2878)) and not (layer5_outputs(2874));
    layer6_outputs(4963) <= (layer5_outputs(1402)) xor (layer5_outputs(1253));
    layer6_outputs(4964) <= (layer5_outputs(6087)) and (layer5_outputs(550));
    layer6_outputs(4965) <= not(layer5_outputs(2061));
    layer6_outputs(4966) <= layer5_outputs(2982);
    layer6_outputs(4967) <= layer5_outputs(2269);
    layer6_outputs(4968) <= (layer5_outputs(1967)) and not (layer5_outputs(4630));
    layer6_outputs(4969) <= layer5_outputs(2078);
    layer6_outputs(4970) <= not((layer5_outputs(4519)) or (layer5_outputs(4979)));
    layer6_outputs(4971) <= (layer5_outputs(6734)) or (layer5_outputs(1687));
    layer6_outputs(4972) <= not((layer5_outputs(1170)) and (layer5_outputs(2543)));
    layer6_outputs(4973) <= not(layer5_outputs(349));
    layer6_outputs(4974) <= not(layer5_outputs(5928));
    layer6_outputs(4975) <= not(layer5_outputs(598)) or (layer5_outputs(1533));
    layer6_outputs(4976) <= not(layer5_outputs(1854));
    layer6_outputs(4977) <= not((layer5_outputs(4585)) xor (layer5_outputs(4632)));
    layer6_outputs(4978) <= not((layer5_outputs(2492)) and (layer5_outputs(4594)));
    layer6_outputs(4979) <= layer5_outputs(4502);
    layer6_outputs(4980) <= (layer5_outputs(2107)) xor (layer5_outputs(729));
    layer6_outputs(4981) <= '1';
    layer6_outputs(4982) <= layer5_outputs(5436);
    layer6_outputs(4983) <= (layer5_outputs(1307)) xor (layer5_outputs(389));
    layer6_outputs(4984) <= not(layer5_outputs(5559));
    layer6_outputs(4985) <= layer5_outputs(1017);
    layer6_outputs(4986) <= not(layer5_outputs(2283)) or (layer5_outputs(7185));
    layer6_outputs(4987) <= (layer5_outputs(172)) and not (layer5_outputs(972));
    layer6_outputs(4988) <= (layer5_outputs(7620)) or (layer5_outputs(5908));
    layer6_outputs(4989) <= layer5_outputs(3468);
    layer6_outputs(4990) <= not((layer5_outputs(494)) xor (layer5_outputs(2066)));
    layer6_outputs(4991) <= not((layer5_outputs(617)) and (layer5_outputs(856)));
    layer6_outputs(4992) <= (layer5_outputs(6129)) xor (layer5_outputs(28));
    layer6_outputs(4993) <= (layer5_outputs(1082)) and not (layer5_outputs(6682));
    layer6_outputs(4994) <= not(layer5_outputs(7114));
    layer6_outputs(4995) <= (layer5_outputs(4963)) xor (layer5_outputs(2063));
    layer6_outputs(4996) <= layer5_outputs(5273);
    layer6_outputs(4997) <= not(layer5_outputs(4181));
    layer6_outputs(4998) <= layer5_outputs(6790);
    layer6_outputs(4999) <= (layer5_outputs(3336)) and (layer5_outputs(2460));
    layer6_outputs(5000) <= not(layer5_outputs(2058)) or (layer5_outputs(63));
    layer6_outputs(5001) <= not(layer5_outputs(5827));
    layer6_outputs(5002) <= not((layer5_outputs(2527)) or (layer5_outputs(6848)));
    layer6_outputs(5003) <= not((layer5_outputs(4267)) xor (layer5_outputs(3840)));
    layer6_outputs(5004) <= not(layer5_outputs(7372));
    layer6_outputs(5005) <= layer5_outputs(3343);
    layer6_outputs(5006) <= (layer5_outputs(5914)) xor (layer5_outputs(3666));
    layer6_outputs(5007) <= not(layer5_outputs(4687));
    layer6_outputs(5008) <= layer5_outputs(2688);
    layer6_outputs(5009) <= (layer5_outputs(4938)) or (layer5_outputs(6761));
    layer6_outputs(5010) <= not(layer5_outputs(1131));
    layer6_outputs(5011) <= not(layer5_outputs(1084)) or (layer5_outputs(7574));
    layer6_outputs(5012) <= layer5_outputs(4272);
    layer6_outputs(5013) <= (layer5_outputs(236)) and not (layer5_outputs(3614));
    layer6_outputs(5014) <= layer5_outputs(4462);
    layer6_outputs(5015) <= (layer5_outputs(7213)) and (layer5_outputs(6419));
    layer6_outputs(5016) <= not(layer5_outputs(4270));
    layer6_outputs(5017) <= (layer5_outputs(1550)) and not (layer5_outputs(30));
    layer6_outputs(5018) <= layer5_outputs(6147);
    layer6_outputs(5019) <= not((layer5_outputs(2246)) xor (layer5_outputs(4881)));
    layer6_outputs(5020) <= not(layer5_outputs(7127));
    layer6_outputs(5021) <= not((layer5_outputs(5497)) xor (layer5_outputs(5015)));
    layer6_outputs(5022) <= (layer5_outputs(6117)) and not (layer5_outputs(3908));
    layer6_outputs(5023) <= layer5_outputs(319);
    layer6_outputs(5024) <= (layer5_outputs(4660)) xor (layer5_outputs(5131));
    layer6_outputs(5025) <= not(layer5_outputs(6517));
    layer6_outputs(5026) <= not((layer5_outputs(3535)) xor (layer5_outputs(2818)));
    layer6_outputs(5027) <= not((layer5_outputs(1994)) and (layer5_outputs(7018)));
    layer6_outputs(5028) <= not((layer5_outputs(6311)) xor (layer5_outputs(5422)));
    layer6_outputs(5029) <= not(layer5_outputs(6070));
    layer6_outputs(5030) <= not(layer5_outputs(5579)) or (layer5_outputs(639));
    layer6_outputs(5031) <= not((layer5_outputs(4139)) or (layer5_outputs(6874)));
    layer6_outputs(5032) <= not((layer5_outputs(5152)) xor (layer5_outputs(7534)));
    layer6_outputs(5033) <= not(layer5_outputs(2855));
    layer6_outputs(5034) <= not((layer5_outputs(1207)) xor (layer5_outputs(7242)));
    layer6_outputs(5035) <= not((layer5_outputs(4723)) xor (layer5_outputs(4682)));
    layer6_outputs(5036) <= layer5_outputs(2796);
    layer6_outputs(5037) <= not((layer5_outputs(462)) and (layer5_outputs(2184)));
    layer6_outputs(5038) <= layer5_outputs(7199);
    layer6_outputs(5039) <= '1';
    layer6_outputs(5040) <= not(layer5_outputs(4407));
    layer6_outputs(5041) <= layer5_outputs(4816);
    layer6_outputs(5042) <= not((layer5_outputs(194)) or (layer5_outputs(4090)));
    layer6_outputs(5043) <= (layer5_outputs(4114)) xor (layer5_outputs(5039));
    layer6_outputs(5044) <= layer5_outputs(264);
    layer6_outputs(5045) <= (layer5_outputs(5673)) and not (layer5_outputs(926));
    layer6_outputs(5046) <= (layer5_outputs(4614)) and not (layer5_outputs(7494));
    layer6_outputs(5047) <= (layer5_outputs(2891)) xor (layer5_outputs(6626));
    layer6_outputs(5048) <= not((layer5_outputs(4958)) or (layer5_outputs(355)));
    layer6_outputs(5049) <= not(layer5_outputs(4356)) or (layer5_outputs(5734));
    layer6_outputs(5050) <= not(layer5_outputs(4360));
    layer6_outputs(5051) <= not(layer5_outputs(4843)) or (layer5_outputs(5582));
    layer6_outputs(5052) <= not(layer5_outputs(6881)) or (layer5_outputs(4070));
    layer6_outputs(5053) <= (layer5_outputs(4893)) xor (layer5_outputs(515));
    layer6_outputs(5054) <= layer5_outputs(1318);
    layer6_outputs(5055) <= not(layer5_outputs(1374));
    layer6_outputs(5056) <= (layer5_outputs(6760)) and not (layer5_outputs(6825));
    layer6_outputs(5057) <= not(layer5_outputs(6115));
    layer6_outputs(5058) <= (layer5_outputs(3517)) and not (layer5_outputs(5332));
    layer6_outputs(5059) <= (layer5_outputs(7467)) and not (layer5_outputs(6796));
    layer6_outputs(5060) <= not(layer5_outputs(273));
    layer6_outputs(5061) <= layer5_outputs(3915);
    layer6_outputs(5062) <= not(layer5_outputs(5576));
    layer6_outputs(5063) <= layer5_outputs(5021);
    layer6_outputs(5064) <= not((layer5_outputs(3020)) and (layer5_outputs(2098)));
    layer6_outputs(5065) <= not((layer5_outputs(7010)) and (layer5_outputs(1666)));
    layer6_outputs(5066) <= (layer5_outputs(5551)) and not (layer5_outputs(6395));
    layer6_outputs(5067) <= (layer5_outputs(1863)) xor (layer5_outputs(1076));
    layer6_outputs(5068) <= not(layer5_outputs(3837)) or (layer5_outputs(1027));
    layer6_outputs(5069) <= not(layer5_outputs(3218)) or (layer5_outputs(5696));
    layer6_outputs(5070) <= not(layer5_outputs(5123));
    layer6_outputs(5071) <= not(layer5_outputs(6348)) or (layer5_outputs(6407));
    layer6_outputs(5072) <= not(layer5_outputs(5745));
    layer6_outputs(5073) <= layer5_outputs(2293);
    layer6_outputs(5074) <= not(layer5_outputs(4718));
    layer6_outputs(5075) <= layer5_outputs(1587);
    layer6_outputs(5076) <= layer5_outputs(4032);
    layer6_outputs(5077) <= not((layer5_outputs(6980)) and (layer5_outputs(1080)));
    layer6_outputs(5078) <= (layer5_outputs(1493)) xor (layer5_outputs(5002));
    layer6_outputs(5079) <= not(layer5_outputs(3039));
    layer6_outputs(5080) <= (layer5_outputs(141)) and not (layer5_outputs(7174));
    layer6_outputs(5081) <= layer5_outputs(1722);
    layer6_outputs(5082) <= not(layer5_outputs(7328)) or (layer5_outputs(1200));
    layer6_outputs(5083) <= not(layer5_outputs(4100));
    layer6_outputs(5084) <= not(layer5_outputs(432));
    layer6_outputs(5085) <= (layer5_outputs(4588)) xor (layer5_outputs(2321));
    layer6_outputs(5086) <= not(layer5_outputs(4685));
    layer6_outputs(5087) <= layer5_outputs(5682);
    layer6_outputs(5088) <= not(layer5_outputs(588)) or (layer5_outputs(1432));
    layer6_outputs(5089) <= layer5_outputs(2053);
    layer6_outputs(5090) <= not(layer5_outputs(4247)) or (layer5_outputs(945));
    layer6_outputs(5091) <= layer5_outputs(1705);
    layer6_outputs(5092) <= '1';
    layer6_outputs(5093) <= not(layer5_outputs(2585));
    layer6_outputs(5094) <= not((layer5_outputs(341)) xor (layer5_outputs(2297)));
    layer6_outputs(5095) <= not((layer5_outputs(1802)) xor (layer5_outputs(2507)));
    layer6_outputs(5096) <= (layer5_outputs(5209)) and (layer5_outputs(4934));
    layer6_outputs(5097) <= layer5_outputs(6840);
    layer6_outputs(5098) <= not((layer5_outputs(40)) or (layer5_outputs(1406)));
    layer6_outputs(5099) <= not(layer5_outputs(7231));
    layer6_outputs(5100) <= not(layer5_outputs(4302));
    layer6_outputs(5101) <= not((layer5_outputs(1323)) and (layer5_outputs(3187)));
    layer6_outputs(5102) <= not((layer5_outputs(3898)) and (layer5_outputs(3111)));
    layer6_outputs(5103) <= not(layer5_outputs(2813));
    layer6_outputs(5104) <= layer5_outputs(4260);
    layer6_outputs(5105) <= not(layer5_outputs(2907));
    layer6_outputs(5106) <= not(layer5_outputs(5459)) or (layer5_outputs(1508));
    layer6_outputs(5107) <= not(layer5_outputs(6868));
    layer6_outputs(5108) <= not(layer5_outputs(6375)) or (layer5_outputs(1213));
    layer6_outputs(5109) <= (layer5_outputs(2178)) and (layer5_outputs(5475));
    layer6_outputs(5110) <= not(layer5_outputs(953));
    layer6_outputs(5111) <= not(layer5_outputs(6145));
    layer6_outputs(5112) <= not((layer5_outputs(1664)) and (layer5_outputs(5844)));
    layer6_outputs(5113) <= not(layer5_outputs(1309));
    layer6_outputs(5114) <= not(layer5_outputs(1611)) or (layer5_outputs(1952));
    layer6_outputs(5115) <= not(layer5_outputs(7629));
    layer6_outputs(5116) <= (layer5_outputs(6936)) xor (layer5_outputs(3825));
    layer6_outputs(5117) <= (layer5_outputs(6185)) xor (layer5_outputs(2930));
    layer6_outputs(5118) <= '1';
    layer6_outputs(5119) <= not(layer5_outputs(4511));
    layer6_outputs(5120) <= not(layer5_outputs(2863));
    layer6_outputs(5121) <= not(layer5_outputs(4197));
    layer6_outputs(5122) <= (layer5_outputs(2749)) and not (layer5_outputs(6408));
    layer6_outputs(5123) <= not(layer5_outputs(2671));
    layer6_outputs(5124) <= not(layer5_outputs(6062));
    layer6_outputs(5125) <= not((layer5_outputs(6046)) xor (layer5_outputs(445)));
    layer6_outputs(5126) <= not(layer5_outputs(9));
    layer6_outputs(5127) <= layer5_outputs(6067);
    layer6_outputs(5128) <= not((layer5_outputs(497)) and (layer5_outputs(1693)));
    layer6_outputs(5129) <= not((layer5_outputs(6061)) xor (layer5_outputs(3063)));
    layer6_outputs(5130) <= layer5_outputs(3061);
    layer6_outputs(5131) <= not((layer5_outputs(2993)) or (layer5_outputs(1672)));
    layer6_outputs(5132) <= layer5_outputs(1055);
    layer6_outputs(5133) <= '1';
    layer6_outputs(5134) <= not((layer5_outputs(5097)) xor (layer5_outputs(5969)));
    layer6_outputs(5135) <= (layer5_outputs(4278)) xor (layer5_outputs(97));
    layer6_outputs(5136) <= not((layer5_outputs(7408)) xor (layer5_outputs(6645)));
    layer6_outputs(5137) <= layer5_outputs(1832);
    layer6_outputs(5138) <= not((layer5_outputs(603)) xor (layer5_outputs(6747)));
    layer6_outputs(5139) <= not(layer5_outputs(6642));
    layer6_outputs(5140) <= layer5_outputs(5089);
    layer6_outputs(5141) <= layer5_outputs(5812);
    layer6_outputs(5142) <= not((layer5_outputs(4778)) or (layer5_outputs(3244)));
    layer6_outputs(5143) <= (layer5_outputs(2433)) or (layer5_outputs(2895));
    layer6_outputs(5144) <= not(layer5_outputs(2147));
    layer6_outputs(5145) <= layer5_outputs(2295);
    layer6_outputs(5146) <= not((layer5_outputs(1651)) and (layer5_outputs(3452)));
    layer6_outputs(5147) <= not((layer5_outputs(1541)) xor (layer5_outputs(7390)));
    layer6_outputs(5148) <= not((layer5_outputs(7276)) and (layer5_outputs(6813)));
    layer6_outputs(5149) <= not((layer5_outputs(1842)) or (layer5_outputs(3776)));
    layer6_outputs(5150) <= not(layer5_outputs(6009));
    layer6_outputs(5151) <= not(layer5_outputs(3822));
    layer6_outputs(5152) <= not((layer5_outputs(5774)) xor (layer5_outputs(1773)));
    layer6_outputs(5153) <= not(layer5_outputs(291)) or (layer5_outputs(6200));
    layer6_outputs(5154) <= not(layer5_outputs(5155));
    layer6_outputs(5155) <= (layer5_outputs(4554)) and not (layer5_outputs(959));
    layer6_outputs(5156) <= '1';
    layer6_outputs(5157) <= not(layer5_outputs(4774));
    layer6_outputs(5158) <= layer5_outputs(4348);
    layer6_outputs(5159) <= not(layer5_outputs(7364)) or (layer5_outputs(704));
    layer6_outputs(5160) <= not((layer5_outputs(2750)) xor (layer5_outputs(2766)));
    layer6_outputs(5161) <= not(layer5_outputs(6909));
    layer6_outputs(5162) <= (layer5_outputs(2886)) xor (layer5_outputs(1853));
    layer6_outputs(5163) <= (layer5_outputs(3410)) or (layer5_outputs(4427));
    layer6_outputs(5164) <= layer5_outputs(3351);
    layer6_outputs(5165) <= not(layer5_outputs(4362));
    layer6_outputs(5166) <= layer5_outputs(6829);
    layer6_outputs(5167) <= layer5_outputs(3952);
    layer6_outputs(5168) <= layer5_outputs(5253);
    layer6_outputs(5169) <= layer5_outputs(2323);
    layer6_outputs(5170) <= layer5_outputs(5404);
    layer6_outputs(5171) <= not((layer5_outputs(5334)) xor (layer5_outputs(4808)));
    layer6_outputs(5172) <= not(layer5_outputs(3737));
    layer6_outputs(5173) <= not(layer5_outputs(5510)) or (layer5_outputs(3303));
    layer6_outputs(5174) <= not(layer5_outputs(6798));
    layer6_outputs(5175) <= layer5_outputs(4974);
    layer6_outputs(5176) <= not(layer5_outputs(4877));
    layer6_outputs(5177) <= not(layer5_outputs(1418));
    layer6_outputs(5178) <= (layer5_outputs(5723)) and not (layer5_outputs(2286));
    layer6_outputs(5179) <= not(layer5_outputs(7103)) or (layer5_outputs(5676));
    layer6_outputs(5180) <= (layer5_outputs(1058)) or (layer5_outputs(5348));
    layer6_outputs(5181) <= not((layer5_outputs(4500)) xor (layer5_outputs(2610)));
    layer6_outputs(5182) <= not((layer5_outputs(1616)) or (layer5_outputs(4594)));
    layer6_outputs(5183) <= (layer5_outputs(91)) and not (layer5_outputs(5801));
    layer6_outputs(5184) <= not(layer5_outputs(1040));
    layer6_outputs(5185) <= not((layer5_outputs(3127)) xor (layer5_outputs(6724)));
    layer6_outputs(5186) <= layer5_outputs(2551);
    layer6_outputs(5187) <= not(layer5_outputs(3728));
    layer6_outputs(5188) <= not((layer5_outputs(5338)) or (layer5_outputs(2578)));
    layer6_outputs(5189) <= not(layer5_outputs(3356));
    layer6_outputs(5190) <= not(layer5_outputs(4498));
    layer6_outputs(5191) <= not(layer5_outputs(978));
    layer6_outputs(5192) <= layer5_outputs(2568);
    layer6_outputs(5193) <= not(layer5_outputs(3257));
    layer6_outputs(5194) <= not((layer5_outputs(2555)) and (layer5_outputs(553)));
    layer6_outputs(5195) <= not(layer5_outputs(5818));
    layer6_outputs(5196) <= (layer5_outputs(6100)) xor (layer5_outputs(3771));
    layer6_outputs(5197) <= not((layer5_outputs(1620)) and (layer5_outputs(794)));
    layer6_outputs(5198) <= layer5_outputs(7183);
    layer6_outputs(5199) <= layer5_outputs(193);
    layer6_outputs(5200) <= layer5_outputs(2984);
    layer6_outputs(5201) <= not(layer5_outputs(7492));
    layer6_outputs(5202) <= not(layer5_outputs(3891)) or (layer5_outputs(598));
    layer6_outputs(5203) <= not((layer5_outputs(5627)) and (layer5_outputs(3994)));
    layer6_outputs(5204) <= not((layer5_outputs(2977)) xor (layer5_outputs(5681)));
    layer6_outputs(5205) <= not(layer5_outputs(3548));
    layer6_outputs(5206) <= not(layer5_outputs(5048)) or (layer5_outputs(7196));
    layer6_outputs(5207) <= layer5_outputs(7042);
    layer6_outputs(5208) <= not(layer5_outputs(7439));
    layer6_outputs(5209) <= not((layer5_outputs(2452)) xor (layer5_outputs(3852)));
    layer6_outputs(5210) <= '1';
    layer6_outputs(5211) <= not(layer5_outputs(1379));
    layer6_outputs(5212) <= layer5_outputs(3511);
    layer6_outputs(5213) <= not(layer5_outputs(4337));
    layer6_outputs(5214) <= not(layer5_outputs(3234));
    layer6_outputs(5215) <= not(layer5_outputs(766));
    layer6_outputs(5216) <= not((layer5_outputs(6776)) xor (layer5_outputs(4648)));
    layer6_outputs(5217) <= layer5_outputs(5306);
    layer6_outputs(5218) <= not(layer5_outputs(4344));
    layer6_outputs(5219) <= not(layer5_outputs(327));
    layer6_outputs(5220) <= not(layer5_outputs(510)) or (layer5_outputs(712));
    layer6_outputs(5221) <= not(layer5_outputs(3118));
    layer6_outputs(5222) <= (layer5_outputs(2658)) and (layer5_outputs(5240));
    layer6_outputs(5223) <= (layer5_outputs(403)) and not (layer5_outputs(2478));
    layer6_outputs(5224) <= not((layer5_outputs(3069)) xor (layer5_outputs(1827)));
    layer6_outputs(5225) <= not(layer5_outputs(4736)) or (layer5_outputs(1343));
    layer6_outputs(5226) <= not(layer5_outputs(7538));
    layer6_outputs(5227) <= not((layer5_outputs(4020)) and (layer5_outputs(4733)));
    layer6_outputs(5228) <= layer5_outputs(3411);
    layer6_outputs(5229) <= (layer5_outputs(3568)) or (layer5_outputs(6017));
    layer6_outputs(5230) <= not(layer5_outputs(3434));
    layer6_outputs(5231) <= not(layer5_outputs(6254));
    layer6_outputs(5232) <= layer5_outputs(7243);
    layer6_outputs(5233) <= not((layer5_outputs(218)) xor (layer5_outputs(4006)));
    layer6_outputs(5234) <= (layer5_outputs(3545)) xor (layer5_outputs(6074));
    layer6_outputs(5235) <= not((layer5_outputs(6042)) and (layer5_outputs(2284)));
    layer6_outputs(5236) <= (layer5_outputs(1330)) xor (layer5_outputs(1515));
    layer6_outputs(5237) <= not((layer5_outputs(5915)) xor (layer5_outputs(5011)));
    layer6_outputs(5238) <= not(layer5_outputs(5704));
    layer6_outputs(5239) <= layer5_outputs(11);
    layer6_outputs(5240) <= (layer5_outputs(6177)) and not (layer5_outputs(989));
    layer6_outputs(5241) <= (layer5_outputs(3468)) xor (layer5_outputs(1518));
    layer6_outputs(5242) <= not(layer5_outputs(352));
    layer6_outputs(5243) <= layer5_outputs(5412);
    layer6_outputs(5244) <= layer5_outputs(1782);
    layer6_outputs(5245) <= not((layer5_outputs(2929)) or (layer5_outputs(863)));
    layer6_outputs(5246) <= layer5_outputs(1470);
    layer6_outputs(5247) <= not((layer5_outputs(7330)) and (layer5_outputs(6073)));
    layer6_outputs(5248) <= not(layer5_outputs(369));
    layer6_outputs(5249) <= not(layer5_outputs(3027));
    layer6_outputs(5250) <= not(layer5_outputs(3321));
    layer6_outputs(5251) <= layer5_outputs(382);
    layer6_outputs(5252) <= not(layer5_outputs(6007));
    layer6_outputs(5253) <= (layer5_outputs(2525)) or (layer5_outputs(3576));
    layer6_outputs(5254) <= not(layer5_outputs(820));
    layer6_outputs(5255) <= (layer5_outputs(2656)) and not (layer5_outputs(3811));
    layer6_outputs(5256) <= (layer5_outputs(1599)) xor (layer5_outputs(6509));
    layer6_outputs(5257) <= layer5_outputs(5013);
    layer6_outputs(5258) <= layer5_outputs(1947);
    layer6_outputs(5259) <= not(layer5_outputs(6455));
    layer6_outputs(5260) <= not(layer5_outputs(3610)) or (layer5_outputs(3819));
    layer6_outputs(5261) <= not(layer5_outputs(2908));
    layer6_outputs(5262) <= not(layer5_outputs(2394));
    layer6_outputs(5263) <= not((layer5_outputs(5839)) or (layer5_outputs(2456)));
    layer6_outputs(5264) <= (layer5_outputs(5975)) xor (layer5_outputs(4643));
    layer6_outputs(5265) <= (layer5_outputs(7264)) and not (layer5_outputs(4463));
    layer6_outputs(5266) <= layer5_outputs(5320);
    layer6_outputs(5267) <= layer5_outputs(4547);
    layer6_outputs(5268) <= not(layer5_outputs(1732)) or (layer5_outputs(3902));
    layer6_outputs(5269) <= not(layer5_outputs(2493));
    layer6_outputs(5270) <= layer5_outputs(6115);
    layer6_outputs(5271) <= not(layer5_outputs(4414));
    layer6_outputs(5272) <= not((layer5_outputs(2721)) and (layer5_outputs(2143)));
    layer6_outputs(5273) <= layer5_outputs(7001);
    layer6_outputs(5274) <= not((layer5_outputs(7340)) xor (layer5_outputs(1066)));
    layer6_outputs(5275) <= layer5_outputs(4222);
    layer6_outputs(5276) <= layer5_outputs(128);
    layer6_outputs(5277) <= (layer5_outputs(798)) and (layer5_outputs(964));
    layer6_outputs(5278) <= layer5_outputs(4638);
    layer6_outputs(5279) <= not((layer5_outputs(632)) xor (layer5_outputs(3396)));
    layer6_outputs(5280) <= not((layer5_outputs(1313)) and (layer5_outputs(6819)));
    layer6_outputs(5281) <= layer5_outputs(725);
    layer6_outputs(5282) <= not(layer5_outputs(268));
    layer6_outputs(5283) <= layer5_outputs(613);
    layer6_outputs(5284) <= not((layer5_outputs(119)) xor (layer5_outputs(2781)));
    layer6_outputs(5285) <= not(layer5_outputs(2677));
    layer6_outputs(5286) <= (layer5_outputs(10)) xor (layer5_outputs(1512));
    layer6_outputs(5287) <= layer5_outputs(2789);
    layer6_outputs(5288) <= layer5_outputs(6931);
    layer6_outputs(5289) <= not(layer5_outputs(2892));
    layer6_outputs(5290) <= (layer5_outputs(5662)) xor (layer5_outputs(1609));
    layer6_outputs(5291) <= (layer5_outputs(4217)) xor (layer5_outputs(7427));
    layer6_outputs(5292) <= (layer5_outputs(7076)) xor (layer5_outputs(6591));
    layer6_outputs(5293) <= layer5_outputs(5422);
    layer6_outputs(5294) <= (layer5_outputs(5949)) xor (layer5_outputs(6246));
    layer6_outputs(5295) <= layer5_outputs(6421);
    layer6_outputs(5296) <= (layer5_outputs(3994)) and (layer5_outputs(1247));
    layer6_outputs(5297) <= layer5_outputs(3982);
    layer6_outputs(5298) <= layer5_outputs(1643);
    layer6_outputs(5299) <= (layer5_outputs(2470)) or (layer5_outputs(5612));
    layer6_outputs(5300) <= layer5_outputs(6401);
    layer6_outputs(5301) <= not((layer5_outputs(909)) xor (layer5_outputs(5875)));
    layer6_outputs(5302) <= not(layer5_outputs(1896));
    layer6_outputs(5303) <= not(layer5_outputs(70));
    layer6_outputs(5304) <= layer5_outputs(2187);
    layer6_outputs(5305) <= not(layer5_outputs(6396));
    layer6_outputs(5306) <= layer5_outputs(5624);
    layer6_outputs(5307) <= (layer5_outputs(473)) and not (layer5_outputs(1140));
    layer6_outputs(5308) <= not(layer5_outputs(4649));
    layer6_outputs(5309) <= not(layer5_outputs(2917)) or (layer5_outputs(1528));
    layer6_outputs(5310) <= not((layer5_outputs(2666)) xor (layer5_outputs(6700)));
    layer6_outputs(5311) <= not((layer5_outputs(3455)) xor (layer5_outputs(3432)));
    layer6_outputs(5312) <= (layer5_outputs(4976)) and not (layer5_outputs(2928));
    layer6_outputs(5313) <= (layer5_outputs(5006)) and not (layer5_outputs(6054));
    layer6_outputs(5314) <= not((layer5_outputs(5889)) or (layer5_outputs(1501)));
    layer6_outputs(5315) <= not((layer5_outputs(6947)) or (layer5_outputs(4266)));
    layer6_outputs(5316) <= (layer5_outputs(5952)) or (layer5_outputs(2919));
    layer6_outputs(5317) <= not(layer5_outputs(568));
    layer6_outputs(5318) <= layer5_outputs(5347);
    layer6_outputs(5319) <= not(layer5_outputs(5537));
    layer6_outputs(5320) <= (layer5_outputs(905)) xor (layer5_outputs(2643));
    layer6_outputs(5321) <= (layer5_outputs(3050)) and (layer5_outputs(4199));
    layer6_outputs(5322) <= not(layer5_outputs(6905));
    layer6_outputs(5323) <= not((layer5_outputs(3702)) xor (layer5_outputs(1217)));
    layer6_outputs(5324) <= layer5_outputs(3196);
    layer6_outputs(5325) <= not(layer5_outputs(3419));
    layer6_outputs(5326) <= not(layer5_outputs(2298));
    layer6_outputs(5327) <= layer5_outputs(3094);
    layer6_outputs(5328) <= layer5_outputs(2286);
    layer6_outputs(5329) <= layer5_outputs(7202);
    layer6_outputs(5330) <= not((layer5_outputs(7227)) xor (layer5_outputs(955)));
    layer6_outputs(5331) <= layer5_outputs(5435);
    layer6_outputs(5332) <= not(layer5_outputs(6653));
    layer6_outputs(5333) <= not((layer5_outputs(6688)) xor (layer5_outputs(907)));
    layer6_outputs(5334) <= not(layer5_outputs(4405));
    layer6_outputs(5335) <= not(layer5_outputs(5197));
    layer6_outputs(5336) <= (layer5_outputs(2630)) or (layer5_outputs(2685));
    layer6_outputs(5337) <= not((layer5_outputs(2408)) and (layer5_outputs(1474)));
    layer6_outputs(5338) <= not(layer5_outputs(1037));
    layer6_outputs(5339) <= (layer5_outputs(238)) or (layer5_outputs(7225));
    layer6_outputs(5340) <= layer5_outputs(2756);
    layer6_outputs(5341) <= layer5_outputs(2171);
    layer6_outputs(5342) <= not(layer5_outputs(6140));
    layer6_outputs(5343) <= not((layer5_outputs(6018)) xor (layer5_outputs(4290)));
    layer6_outputs(5344) <= not(layer5_outputs(3683)) or (layer5_outputs(3106));
    layer6_outputs(5345) <= layer5_outputs(1250);
    layer6_outputs(5346) <= not((layer5_outputs(2092)) and (layer5_outputs(3483)));
    layer6_outputs(5347) <= not((layer5_outputs(3706)) xor (layer5_outputs(4625)));
    layer6_outputs(5348) <= not(layer5_outputs(3171));
    layer6_outputs(5349) <= layer5_outputs(3569);
    layer6_outputs(5350) <= layer5_outputs(7207);
    layer6_outputs(5351) <= not(layer5_outputs(3008)) or (layer5_outputs(2576));
    layer6_outputs(5352) <= not(layer5_outputs(1364)) or (layer5_outputs(5280));
    layer6_outputs(5353) <= (layer5_outputs(6549)) or (layer5_outputs(4860));
    layer6_outputs(5354) <= not((layer5_outputs(1520)) or (layer5_outputs(730)));
    layer6_outputs(5355) <= not(layer5_outputs(3704));
    layer6_outputs(5356) <= (layer5_outputs(6179)) or (layer5_outputs(2279));
    layer6_outputs(5357) <= layer5_outputs(6876);
    layer6_outputs(5358) <= not((layer5_outputs(5587)) or (layer5_outputs(7187)));
    layer6_outputs(5359) <= not(layer5_outputs(158));
    layer6_outputs(5360) <= not(layer5_outputs(6780));
    layer6_outputs(5361) <= not(layer5_outputs(6711));
    layer6_outputs(5362) <= layer5_outputs(5229);
    layer6_outputs(5363) <= (layer5_outputs(6646)) xor (layer5_outputs(4127));
    layer6_outputs(5364) <= not(layer5_outputs(2876));
    layer6_outputs(5365) <= layer5_outputs(4837);
    layer6_outputs(5366) <= (layer5_outputs(5803)) and not (layer5_outputs(3489));
    layer6_outputs(5367) <= (layer5_outputs(7001)) xor (layer5_outputs(5804));
    layer6_outputs(5368) <= not(layer5_outputs(5313));
    layer6_outputs(5369) <= layer5_outputs(3672);
    layer6_outputs(5370) <= layer5_outputs(6111);
    layer6_outputs(5371) <= not((layer5_outputs(6501)) and (layer5_outputs(1911)));
    layer6_outputs(5372) <= not(layer5_outputs(2299)) or (layer5_outputs(4471));
    layer6_outputs(5373) <= not(layer5_outputs(569));
    layer6_outputs(5374) <= layer5_outputs(4749);
    layer6_outputs(5375) <= not(layer5_outputs(1805));
    layer6_outputs(5376) <= not(layer5_outputs(4489));
    layer6_outputs(5377) <= not((layer5_outputs(5562)) and (layer5_outputs(6191)));
    layer6_outputs(5378) <= not((layer5_outputs(914)) xor (layer5_outputs(6924)));
    layer6_outputs(5379) <= (layer5_outputs(469)) and not (layer5_outputs(3024));
    layer6_outputs(5380) <= not((layer5_outputs(6672)) and (layer5_outputs(5438)));
    layer6_outputs(5381) <= '0';
    layer6_outputs(5382) <= layer5_outputs(6250);
    layer6_outputs(5383) <= layer5_outputs(2237);
    layer6_outputs(5384) <= not((layer5_outputs(810)) and (layer5_outputs(6239)));
    layer6_outputs(5385) <= not(layer5_outputs(1164));
    layer6_outputs(5386) <= (layer5_outputs(6833)) or (layer5_outputs(3000));
    layer6_outputs(5387) <= not(layer5_outputs(809));
    layer6_outputs(5388) <= not(layer5_outputs(438));
    layer6_outputs(5389) <= layer5_outputs(2686);
    layer6_outputs(5390) <= not(layer5_outputs(2417));
    layer6_outputs(5391) <= not(layer5_outputs(3730));
    layer6_outputs(5392) <= (layer5_outputs(2724)) and (layer5_outputs(5999));
    layer6_outputs(5393) <= layer5_outputs(3988);
    layer6_outputs(5394) <= not((layer5_outputs(1367)) xor (layer5_outputs(4856)));
    layer6_outputs(5395) <= layer5_outputs(6097);
    layer6_outputs(5396) <= '1';
    layer6_outputs(5397) <= layer5_outputs(499);
    layer6_outputs(5398) <= layer5_outputs(586);
    layer6_outputs(5399) <= layer5_outputs(2758);
    layer6_outputs(5400) <= not(layer5_outputs(3416));
    layer6_outputs(5401) <= not((layer5_outputs(4789)) and (layer5_outputs(1086)));
    layer6_outputs(5402) <= not(layer5_outputs(5283)) or (layer5_outputs(405));
    layer6_outputs(5403) <= not((layer5_outputs(6551)) or (layer5_outputs(2690)));
    layer6_outputs(5404) <= layer5_outputs(5455);
    layer6_outputs(5405) <= not((layer5_outputs(3168)) and (layer5_outputs(3916)));
    layer6_outputs(5406) <= (layer5_outputs(3554)) and not (layer5_outputs(1214));
    layer6_outputs(5407) <= (layer5_outputs(6063)) and not (layer5_outputs(3564));
    layer6_outputs(5408) <= (layer5_outputs(6361)) and (layer5_outputs(42));
    layer6_outputs(5409) <= (layer5_outputs(1087)) and not (layer5_outputs(6665));
    layer6_outputs(5410) <= not((layer5_outputs(4925)) or (layer5_outputs(3543)));
    layer6_outputs(5411) <= layer5_outputs(6629);
    layer6_outputs(5412) <= layer5_outputs(4204);
    layer6_outputs(5413) <= not((layer5_outputs(5444)) xor (layer5_outputs(3185)));
    layer6_outputs(5414) <= not(layer5_outputs(2250)) or (layer5_outputs(6366));
    layer6_outputs(5415) <= not(layer5_outputs(2415)) or (layer5_outputs(5335));
    layer6_outputs(5416) <= not((layer5_outputs(1005)) or (layer5_outputs(1293)));
    layer6_outputs(5417) <= not(layer5_outputs(6360));
    layer6_outputs(5418) <= not(layer5_outputs(2842));
    layer6_outputs(5419) <= not(layer5_outputs(5630));
    layer6_outputs(5420) <= not(layer5_outputs(6159)) or (layer5_outputs(1628));
    layer6_outputs(5421) <= not((layer5_outputs(5122)) xor (layer5_outputs(7618)));
    layer6_outputs(5422) <= layer5_outputs(2837);
    layer6_outputs(5423) <= not((layer5_outputs(6956)) and (layer5_outputs(6187)));
    layer6_outputs(5424) <= not(layer5_outputs(7067));
    layer6_outputs(5425) <= layer5_outputs(4376);
    layer6_outputs(5426) <= not((layer5_outputs(5903)) and (layer5_outputs(5425)));
    layer6_outputs(5427) <= (layer5_outputs(4335)) and not (layer5_outputs(2557));
    layer6_outputs(5428) <= not((layer5_outputs(5999)) or (layer5_outputs(826)));
    layer6_outputs(5429) <= (layer5_outputs(4725)) and not (layer5_outputs(5701));
    layer6_outputs(5430) <= not(layer5_outputs(3067)) or (layer5_outputs(1861));
    layer6_outputs(5431) <= layer5_outputs(7341);
    layer6_outputs(5432) <= layer5_outputs(2925);
    layer6_outputs(5433) <= not(layer5_outputs(3257));
    layer6_outputs(5434) <= not(layer5_outputs(6627));
    layer6_outputs(5435) <= layer5_outputs(6114);
    layer6_outputs(5436) <= (layer5_outputs(3941)) and not (layer5_outputs(1849));
    layer6_outputs(5437) <= (layer5_outputs(3833)) and (layer5_outputs(1038));
    layer6_outputs(5438) <= layer5_outputs(2036);
    layer6_outputs(5439) <= not((layer5_outputs(431)) and (layer5_outputs(2526)));
    layer6_outputs(5440) <= (layer5_outputs(1912)) and not (layer5_outputs(3645));
    layer6_outputs(5441) <= not(layer5_outputs(4235));
    layer6_outputs(5442) <= layer5_outputs(6216);
    layer6_outputs(5443) <= not(layer5_outputs(1011));
    layer6_outputs(5444) <= not(layer5_outputs(7343));
    layer6_outputs(5445) <= not(layer5_outputs(4182));
    layer6_outputs(5446) <= not(layer5_outputs(496));
    layer6_outputs(5447) <= not((layer5_outputs(4565)) or (layer5_outputs(5909)));
    layer6_outputs(5448) <= (layer5_outputs(7480)) xor (layer5_outputs(934));
    layer6_outputs(5449) <= layer5_outputs(2039);
    layer6_outputs(5450) <= layer5_outputs(2131);
    layer6_outputs(5451) <= not((layer5_outputs(1962)) and (layer5_outputs(3144)));
    layer6_outputs(5452) <= not(layer5_outputs(3253));
    layer6_outputs(5453) <= layer5_outputs(1099);
    layer6_outputs(5454) <= not(layer5_outputs(2366));
    layer6_outputs(5455) <= layer5_outputs(1744);
    layer6_outputs(5456) <= layer5_outputs(6445);
    layer6_outputs(5457) <= not(layer5_outputs(1104));
    layer6_outputs(5458) <= (layer5_outputs(1207)) and not (layer5_outputs(6453));
    layer6_outputs(5459) <= not(layer5_outputs(1036));
    layer6_outputs(5460) <= layer5_outputs(4350);
    layer6_outputs(5461) <= layer5_outputs(3240);
    layer6_outputs(5462) <= (layer5_outputs(3775)) or (layer5_outputs(7674));
    layer6_outputs(5463) <= layer5_outputs(7258);
    layer6_outputs(5464) <= not((layer5_outputs(2261)) or (layer5_outputs(1564)));
    layer6_outputs(5465) <= not(layer5_outputs(3111)) or (layer5_outputs(2280));
    layer6_outputs(5466) <= not(layer5_outputs(4384));
    layer6_outputs(5467) <= not(layer5_outputs(6351));
    layer6_outputs(5468) <= not((layer5_outputs(889)) xor (layer5_outputs(2805)));
    layer6_outputs(5469) <= not((layer5_outputs(6154)) or (layer5_outputs(6571)));
    layer6_outputs(5470) <= layer5_outputs(7016);
    layer6_outputs(5471) <= (layer5_outputs(4348)) and not (layer5_outputs(2381));
    layer6_outputs(5472) <= not((layer5_outputs(4932)) xor (layer5_outputs(6573)));
    layer6_outputs(5473) <= (layer5_outputs(277)) and (layer5_outputs(2842));
    layer6_outputs(5474) <= not(layer5_outputs(247)) or (layer5_outputs(5224));
    layer6_outputs(5475) <= not((layer5_outputs(4540)) xor (layer5_outputs(1116)));
    layer6_outputs(5476) <= not(layer5_outputs(5319)) or (layer5_outputs(5231));
    layer6_outputs(5477) <= not(layer5_outputs(3276));
    layer6_outputs(5478) <= layer5_outputs(4386);
    layer6_outputs(5479) <= layer5_outputs(6399);
    layer6_outputs(5480) <= (layer5_outputs(3276)) and (layer5_outputs(2433));
    layer6_outputs(5481) <= (layer5_outputs(2352)) xor (layer5_outputs(5955));
    layer6_outputs(5482) <= layer5_outputs(6056);
    layer6_outputs(5483) <= not(layer5_outputs(531));
    layer6_outputs(5484) <= not((layer5_outputs(6772)) and (layer5_outputs(2299)));
    layer6_outputs(5485) <= not(layer5_outputs(2579));
    layer6_outputs(5486) <= layer5_outputs(1740);
    layer6_outputs(5487) <= not(layer5_outputs(446)) or (layer5_outputs(3043));
    layer6_outputs(5488) <= not(layer5_outputs(3636)) or (layer5_outputs(4589));
    layer6_outputs(5489) <= not(layer5_outputs(1455));
    layer6_outputs(5490) <= layer5_outputs(2965);
    layer6_outputs(5491) <= not(layer5_outputs(2966));
    layer6_outputs(5492) <= (layer5_outputs(955)) and (layer5_outputs(4925));
    layer6_outputs(5493) <= not(layer5_outputs(1060)) or (layer5_outputs(7320));
    layer6_outputs(5494) <= not(layer5_outputs(1201));
    layer6_outputs(5495) <= '1';
    layer6_outputs(5496) <= not((layer5_outputs(4439)) or (layer5_outputs(3448)));
    layer6_outputs(5497) <= layer5_outputs(3231);
    layer6_outputs(5498) <= layer5_outputs(1726);
    layer6_outputs(5499) <= layer5_outputs(750);
    layer6_outputs(5500) <= not(layer5_outputs(6816));
    layer6_outputs(5501) <= not(layer5_outputs(724)) or (layer5_outputs(5699));
    layer6_outputs(5502) <= (layer5_outputs(2010)) and not (layer5_outputs(3124));
    layer6_outputs(5503) <= not(layer5_outputs(1424));
    layer6_outputs(5504) <= not(layer5_outputs(1108)) or (layer5_outputs(2151));
    layer6_outputs(5505) <= not((layer5_outputs(5775)) xor (layer5_outputs(3773)));
    layer6_outputs(5506) <= not(layer5_outputs(4377)) or (layer5_outputs(476));
    layer6_outputs(5507) <= (layer5_outputs(116)) and not (layer5_outputs(6518));
    layer6_outputs(5508) <= (layer5_outputs(5333)) xor (layer5_outputs(6372));
    layer6_outputs(5509) <= (layer5_outputs(6730)) or (layer5_outputs(3377));
    layer6_outputs(5510) <= layer5_outputs(3724);
    layer6_outputs(5511) <= not(layer5_outputs(5101));
    layer6_outputs(5512) <= not(layer5_outputs(4559)) or (layer5_outputs(1670));
    layer6_outputs(5513) <= not(layer5_outputs(930));
    layer6_outputs(5514) <= not((layer5_outputs(1054)) or (layer5_outputs(7163)));
    layer6_outputs(5515) <= not(layer5_outputs(4398));
    layer6_outputs(5516) <= layer5_outputs(942);
    layer6_outputs(5517) <= layer5_outputs(564);
    layer6_outputs(5518) <= not(layer5_outputs(5084));
    layer6_outputs(5519) <= layer5_outputs(5366);
    layer6_outputs(5520) <= layer5_outputs(5354);
    layer6_outputs(5521) <= (layer5_outputs(4486)) or (layer5_outputs(5155));
    layer6_outputs(5522) <= layer5_outputs(3010);
    layer6_outputs(5523) <= layer5_outputs(1913);
    layer6_outputs(5524) <= not(layer5_outputs(3622)) or (layer5_outputs(903));
    layer6_outputs(5525) <= (layer5_outputs(5324)) and not (layer5_outputs(4471));
    layer6_outputs(5526) <= layer5_outputs(4701);
    layer6_outputs(5527) <= layer5_outputs(12);
    layer6_outputs(5528) <= not(layer5_outputs(1059));
    layer6_outputs(5529) <= not(layer5_outputs(3717));
    layer6_outputs(5530) <= not(layer5_outputs(3523)) or (layer5_outputs(3441));
    layer6_outputs(5531) <= not(layer5_outputs(804)) or (layer5_outputs(3069));
    layer6_outputs(5532) <= not((layer5_outputs(6926)) and (layer5_outputs(764)));
    layer6_outputs(5533) <= not(layer5_outputs(6801));
    layer6_outputs(5534) <= layer5_outputs(2338);
    layer6_outputs(5535) <= not((layer5_outputs(2508)) xor (layer5_outputs(672)));
    layer6_outputs(5536) <= layer5_outputs(2883);
    layer6_outputs(5537) <= layer5_outputs(6991);
    layer6_outputs(5538) <= not(layer5_outputs(7159));
    layer6_outputs(5539) <= not(layer5_outputs(173)) or (layer5_outputs(5771));
    layer6_outputs(5540) <= (layer5_outputs(4036)) or (layer5_outputs(6522));
    layer6_outputs(5541) <= (layer5_outputs(7146)) xor (layer5_outputs(3860));
    layer6_outputs(5542) <= (layer5_outputs(5209)) or (layer5_outputs(1372));
    layer6_outputs(5543) <= not(layer5_outputs(1637));
    layer6_outputs(5544) <= not(layer5_outputs(2799)) or (layer5_outputs(5018));
    layer6_outputs(5545) <= not((layer5_outputs(7377)) xor (layer5_outputs(2538)));
    layer6_outputs(5546) <= not(layer5_outputs(1244));
    layer6_outputs(5547) <= not((layer5_outputs(737)) xor (layer5_outputs(4301)));
    layer6_outputs(5548) <= not((layer5_outputs(6368)) and (layer5_outputs(4740)));
    layer6_outputs(5549) <= layer5_outputs(2422);
    layer6_outputs(5550) <= not(layer5_outputs(2013)) or (layer5_outputs(43));
    layer6_outputs(5551) <= (layer5_outputs(4767)) and not (layer5_outputs(6993));
    layer6_outputs(5552) <= not(layer5_outputs(1204));
    layer6_outputs(5553) <= not(layer5_outputs(4776));
    layer6_outputs(5554) <= not((layer5_outputs(4314)) xor (layer5_outputs(5654)));
    layer6_outputs(5555) <= not(layer5_outputs(7575));
    layer6_outputs(5556) <= layer5_outputs(6659);
    layer6_outputs(5557) <= not(layer5_outputs(5769));
    layer6_outputs(5558) <= not(layer5_outputs(4956));
    layer6_outputs(5559) <= not((layer5_outputs(4803)) xor (layer5_outputs(6544)));
    layer6_outputs(5560) <= not(layer5_outputs(6973));
    layer6_outputs(5561) <= not((layer5_outputs(4455)) xor (layer5_outputs(7667)));
    layer6_outputs(5562) <= not((layer5_outputs(7455)) xor (layer5_outputs(1420)));
    layer6_outputs(5563) <= (layer5_outputs(7384)) and (layer5_outputs(3278));
    layer6_outputs(5564) <= not(layer5_outputs(577));
    layer6_outputs(5565) <= not((layer5_outputs(7033)) xor (layer5_outputs(4251)));
    layer6_outputs(5566) <= (layer5_outputs(7150)) and (layer5_outputs(5266));
    layer6_outputs(5567) <= layer5_outputs(3892);
    layer6_outputs(5568) <= layer5_outputs(3664);
    layer6_outputs(5569) <= (layer5_outputs(7335)) xor (layer5_outputs(811));
    layer6_outputs(5570) <= not(layer5_outputs(354));
    layer6_outputs(5571) <= (layer5_outputs(4186)) or (layer5_outputs(6864));
    layer6_outputs(5572) <= not(layer5_outputs(612)) or (layer5_outputs(3577));
    layer6_outputs(5573) <= not(layer5_outputs(7368));
    layer6_outputs(5574) <= layer5_outputs(7180);
    layer6_outputs(5575) <= (layer5_outputs(6964)) and not (layer5_outputs(5143));
    layer6_outputs(5576) <= not(layer5_outputs(3926));
    layer6_outputs(5577) <= (layer5_outputs(2023)) xor (layer5_outputs(6089));
    layer6_outputs(5578) <= (layer5_outputs(2133)) and not (layer5_outputs(136));
    layer6_outputs(5579) <= layer5_outputs(3059);
    layer6_outputs(5580) <= not(layer5_outputs(2794));
    layer6_outputs(5581) <= not(layer5_outputs(1229));
    layer6_outputs(5582) <= (layer5_outputs(4451)) xor (layer5_outputs(7068));
    layer6_outputs(5583) <= not(layer5_outputs(6620)) or (layer5_outputs(569));
    layer6_outputs(5584) <= (layer5_outputs(3136)) xor (layer5_outputs(154));
    layer6_outputs(5585) <= not(layer5_outputs(961));
    layer6_outputs(5586) <= not(layer5_outputs(2053));
    layer6_outputs(5587) <= (layer5_outputs(4719)) and (layer5_outputs(7308));
    layer6_outputs(5588) <= not(layer5_outputs(751));
    layer6_outputs(5589) <= not(layer5_outputs(5378));
    layer6_outputs(5590) <= layer5_outputs(3716);
    layer6_outputs(5591) <= layer5_outputs(70);
    layer6_outputs(5592) <= (layer5_outputs(5234)) and not (layer5_outputs(7356));
    layer6_outputs(5593) <= not((layer5_outputs(6824)) xor (layer5_outputs(7547)));
    layer6_outputs(5594) <= not(layer5_outputs(357));
    layer6_outputs(5595) <= (layer5_outputs(6096)) xor (layer5_outputs(3751));
    layer6_outputs(5596) <= not((layer5_outputs(5695)) and (layer5_outputs(4012)));
    layer6_outputs(5597) <= not(layer5_outputs(6988)) or (layer5_outputs(5798));
    layer6_outputs(5598) <= not(layer5_outputs(6114));
    layer6_outputs(5599) <= layer5_outputs(3732);
    layer6_outputs(5600) <= (layer5_outputs(6002)) and not (layer5_outputs(3401));
    layer6_outputs(5601) <= (layer5_outputs(2065)) or (layer5_outputs(3148));
    layer6_outputs(5602) <= not(layer5_outputs(6907));
    layer6_outputs(5603) <= not((layer5_outputs(1694)) xor (layer5_outputs(1285)));
    layer6_outputs(5604) <= layer5_outputs(4283);
    layer6_outputs(5605) <= layer5_outputs(1910);
    layer6_outputs(5606) <= layer5_outputs(2987);
    layer6_outputs(5607) <= not((layer5_outputs(6571)) xor (layer5_outputs(3581)));
    layer6_outputs(5608) <= not((layer5_outputs(4973)) xor (layer5_outputs(55)));
    layer6_outputs(5609) <= not(layer5_outputs(6995)) or (layer5_outputs(5084));
    layer6_outputs(5610) <= not(layer5_outputs(5773));
    layer6_outputs(5611) <= layer5_outputs(5016);
    layer6_outputs(5612) <= layer5_outputs(3101);
    layer6_outputs(5613) <= not(layer5_outputs(5452));
    layer6_outputs(5614) <= not(layer5_outputs(1034));
    layer6_outputs(5615) <= not(layer5_outputs(319)) or (layer5_outputs(2844));
    layer6_outputs(5616) <= not((layer5_outputs(3886)) xor (layer5_outputs(1360)));
    layer6_outputs(5617) <= not(layer5_outputs(3203));
    layer6_outputs(5618) <= not(layer5_outputs(2770));
    layer6_outputs(5619) <= layer5_outputs(4960);
    layer6_outputs(5620) <= not(layer5_outputs(7657));
    layer6_outputs(5621) <= (layer5_outputs(3526)) and (layer5_outputs(3007));
    layer6_outputs(5622) <= (layer5_outputs(5370)) xor (layer5_outputs(7343));
    layer6_outputs(5623) <= (layer5_outputs(7607)) or (layer5_outputs(722));
    layer6_outputs(5624) <= layer5_outputs(1863);
    layer6_outputs(5625) <= not((layer5_outputs(1726)) or (layer5_outputs(210)));
    layer6_outputs(5626) <= not(layer5_outputs(5807)) or (layer5_outputs(252));
    layer6_outputs(5627) <= not(layer5_outputs(126));
    layer6_outputs(5628) <= (layer5_outputs(21)) xor (layer5_outputs(7038));
    layer6_outputs(5629) <= not((layer5_outputs(3598)) xor (layer5_outputs(228)));
    layer6_outputs(5630) <= layer5_outputs(3065);
    layer6_outputs(5631) <= not(layer5_outputs(3360));
    layer6_outputs(5632) <= layer5_outputs(4000);
    layer6_outputs(5633) <= (layer5_outputs(670)) and not (layer5_outputs(4558));
    layer6_outputs(5634) <= not(layer5_outputs(7665));
    layer6_outputs(5635) <= not(layer5_outputs(2701));
    layer6_outputs(5636) <= '1';
    layer6_outputs(5637) <= not(layer5_outputs(5093));
    layer6_outputs(5638) <= not(layer5_outputs(6436));
    layer6_outputs(5639) <= (layer5_outputs(872)) and not (layer5_outputs(6184));
    layer6_outputs(5640) <= not(layer5_outputs(3091));
    layer6_outputs(5641) <= layer5_outputs(2045);
    layer6_outputs(5642) <= not(layer5_outputs(4518));
    layer6_outputs(5643) <= layer5_outputs(3789);
    layer6_outputs(5644) <= layer5_outputs(2822);
    layer6_outputs(5645) <= (layer5_outputs(4762)) and not (layer5_outputs(5534));
    layer6_outputs(5646) <= layer5_outputs(1945);
    layer6_outputs(5647) <= layer5_outputs(6178);
    layer6_outputs(5648) <= '0';
    layer6_outputs(5649) <= layer5_outputs(3875);
    layer6_outputs(5650) <= (layer5_outputs(3963)) xor (layer5_outputs(6732));
    layer6_outputs(5651) <= layer5_outputs(3274);
    layer6_outputs(5652) <= layer5_outputs(6946);
    layer6_outputs(5653) <= layer5_outputs(3804);
    layer6_outputs(5654) <= not(layer5_outputs(3943));
    layer6_outputs(5655) <= layer5_outputs(112);
    layer6_outputs(5656) <= not(layer5_outputs(4296));
    layer6_outputs(5657) <= not((layer5_outputs(2178)) or (layer5_outputs(2134)));
    layer6_outputs(5658) <= (layer5_outputs(5090)) and not (layer5_outputs(6590));
    layer6_outputs(5659) <= not(layer5_outputs(5346));
    layer6_outputs(5660) <= layer5_outputs(6443);
    layer6_outputs(5661) <= not(layer5_outputs(2446));
    layer6_outputs(5662) <= not(layer5_outputs(2826));
    layer6_outputs(5663) <= not(layer5_outputs(6972)) or (layer5_outputs(4990));
    layer6_outputs(5664) <= layer5_outputs(2498);
    layer6_outputs(5665) <= not(layer5_outputs(5529));
    layer6_outputs(5666) <= not((layer5_outputs(3104)) xor (layer5_outputs(2736)));
    layer6_outputs(5667) <= not(layer5_outputs(2023)) or (layer5_outputs(6858));
    layer6_outputs(5668) <= not(layer5_outputs(2008));
    layer6_outputs(5669) <= (layer5_outputs(4940)) xor (layer5_outputs(7325));
    layer6_outputs(5670) <= not(layer5_outputs(6430));
    layer6_outputs(5671) <= not(layer5_outputs(6831)) or (layer5_outputs(5836));
    layer6_outputs(5672) <= not((layer5_outputs(4986)) xor (layer5_outputs(975)));
    layer6_outputs(5673) <= not(layer5_outputs(456));
    layer6_outputs(5674) <= (layer5_outputs(2915)) and not (layer5_outputs(615));
    layer6_outputs(5675) <= not(layer5_outputs(3882));
    layer6_outputs(5676) <= not(layer5_outputs(1187));
    layer6_outputs(5677) <= layer5_outputs(4871);
    layer6_outputs(5678) <= layer5_outputs(5304);
    layer6_outputs(5679) <= layer5_outputs(2981);
    layer6_outputs(5680) <= layer5_outputs(132);
    layer6_outputs(5681) <= layer5_outputs(1884);
    layer6_outputs(5682) <= (layer5_outputs(6252)) and (layer5_outputs(4192));
    layer6_outputs(5683) <= layer5_outputs(3774);
    layer6_outputs(5684) <= (layer5_outputs(5088)) xor (layer5_outputs(5950));
    layer6_outputs(5685) <= layer5_outputs(137);
    layer6_outputs(5686) <= not(layer5_outputs(2166));
    layer6_outputs(5687) <= layer5_outputs(2140);
    layer6_outputs(5688) <= not((layer5_outputs(893)) xor (layer5_outputs(5368)));
    layer6_outputs(5689) <= layer5_outputs(5077);
    layer6_outputs(5690) <= not(layer5_outputs(2639)) or (layer5_outputs(464));
    layer6_outputs(5691) <= not((layer5_outputs(2945)) xor (layer5_outputs(7169)));
    layer6_outputs(5692) <= (layer5_outputs(104)) xor (layer5_outputs(7064));
    layer6_outputs(5693) <= (layer5_outputs(265)) xor (layer5_outputs(5225));
    layer6_outputs(5694) <= layer5_outputs(721);
    layer6_outputs(5695) <= (layer5_outputs(6206)) and not (layer5_outputs(6845));
    layer6_outputs(5696) <= not((layer5_outputs(4229)) xor (layer5_outputs(1636)));
    layer6_outputs(5697) <= not(layer5_outputs(358)) or (layer5_outputs(5875));
    layer6_outputs(5698) <= not(layer5_outputs(707)) or (layer5_outputs(1542));
    layer6_outputs(5699) <= layer5_outputs(2293);
    layer6_outputs(5700) <= (layer5_outputs(1485)) and not (layer5_outputs(5219));
    layer6_outputs(5701) <= not(layer5_outputs(5620));
    layer6_outputs(5702) <= not(layer5_outputs(5133));
    layer6_outputs(5703) <= layer5_outputs(4587);
    layer6_outputs(5704) <= layer5_outputs(1981);
    layer6_outputs(5705) <= not((layer5_outputs(3133)) and (layer5_outputs(1803)));
    layer6_outputs(5706) <= layer5_outputs(1911);
    layer6_outputs(5707) <= not(layer5_outputs(4565));
    layer6_outputs(5708) <= not(layer5_outputs(195));
    layer6_outputs(5709) <= layer5_outputs(408);
    layer6_outputs(5710) <= layer5_outputs(7050);
    layer6_outputs(5711) <= not(layer5_outputs(4255)) or (layer5_outputs(4654));
    layer6_outputs(5712) <= (layer5_outputs(6205)) and not (layer5_outputs(6989));
    layer6_outputs(5713) <= not((layer5_outputs(3794)) or (layer5_outputs(6861)));
    layer6_outputs(5714) <= (layer5_outputs(1840)) and not (layer5_outputs(2272));
    layer6_outputs(5715) <= layer5_outputs(3132);
    layer6_outputs(5716) <= not(layer5_outputs(5718));
    layer6_outputs(5717) <= not(layer5_outputs(2697));
    layer6_outputs(5718) <= not(layer5_outputs(5906));
    layer6_outputs(5719) <= layer5_outputs(7102);
    layer6_outputs(5720) <= (layer5_outputs(2607)) and not (layer5_outputs(6373));
    layer6_outputs(5721) <= (layer5_outputs(5736)) and not (layer5_outputs(801));
    layer6_outputs(5722) <= (layer5_outputs(1697)) xor (layer5_outputs(5296));
    layer6_outputs(5723) <= not(layer5_outputs(5840));
    layer6_outputs(5724) <= layer5_outputs(67);
    layer6_outputs(5725) <= not((layer5_outputs(2536)) and (layer5_outputs(1222)));
    layer6_outputs(5726) <= layer5_outputs(3427);
    layer6_outputs(5727) <= layer5_outputs(5683);
    layer6_outputs(5728) <= not(layer5_outputs(3423)) or (layer5_outputs(3709));
    layer6_outputs(5729) <= not((layer5_outputs(1563)) xor (layer5_outputs(4408)));
    layer6_outputs(5730) <= not(layer5_outputs(3321));
    layer6_outputs(5731) <= not((layer5_outputs(4992)) and (layer5_outputs(1174)));
    layer6_outputs(5732) <= (layer5_outputs(5367)) and not (layer5_outputs(4662));
    layer6_outputs(5733) <= not(layer5_outputs(6152));
    layer6_outputs(5734) <= layer5_outputs(1185);
    layer6_outputs(5735) <= layer5_outputs(2705);
    layer6_outputs(5736) <= layer5_outputs(5661);
    layer6_outputs(5737) <= layer5_outputs(50);
    layer6_outputs(5738) <= layer5_outputs(3803);
    layer6_outputs(5739) <= layer5_outputs(2202);
    layer6_outputs(5740) <= not(layer5_outputs(2931));
    layer6_outputs(5741) <= not(layer5_outputs(5144));
    layer6_outputs(5742) <= not(layer5_outputs(7307));
    layer6_outputs(5743) <= (layer5_outputs(6337)) and not (layer5_outputs(6367));
    layer6_outputs(5744) <= not((layer5_outputs(5072)) or (layer5_outputs(7551)));
    layer6_outputs(5745) <= layer5_outputs(6676);
    layer6_outputs(5746) <= layer5_outputs(3098);
    layer6_outputs(5747) <= not(layer5_outputs(7025));
    layer6_outputs(5748) <= (layer5_outputs(5793)) and not (layer5_outputs(7416));
    layer6_outputs(5749) <= not(layer5_outputs(7582));
    layer6_outputs(5750) <= not((layer5_outputs(1390)) xor (layer5_outputs(1632)));
    layer6_outputs(5751) <= (layer5_outputs(5168)) and not (layer5_outputs(4858));
    layer6_outputs(5752) <= (layer5_outputs(336)) and not (layer5_outputs(3883));
    layer6_outputs(5753) <= (layer5_outputs(6614)) and (layer5_outputs(6044));
    layer6_outputs(5754) <= not(layer5_outputs(5397)) or (layer5_outputs(3687));
    layer6_outputs(5755) <= not((layer5_outputs(1824)) or (layer5_outputs(5)));
    layer6_outputs(5756) <= (layer5_outputs(2834)) and not (layer5_outputs(2091));
    layer6_outputs(5757) <= layer5_outputs(62);
    layer6_outputs(5758) <= not(layer5_outputs(3413));
    layer6_outputs(5759) <= not(layer5_outputs(1917));
    layer6_outputs(5760) <= layer5_outputs(5431);
    layer6_outputs(5761) <= not(layer5_outputs(5081));
    layer6_outputs(5762) <= layer5_outputs(6251);
    layer6_outputs(5763) <= (layer5_outputs(2668)) and (layer5_outputs(5891));
    layer6_outputs(5764) <= not(layer5_outputs(6062));
    layer6_outputs(5765) <= not((layer5_outputs(1752)) xor (layer5_outputs(4259)));
    layer6_outputs(5766) <= not((layer5_outputs(2955)) or (layer5_outputs(318)));
    layer6_outputs(5767) <= not(layer5_outputs(862)) or (layer5_outputs(6782));
    layer6_outputs(5768) <= not((layer5_outputs(6154)) and (layer5_outputs(2236)));
    layer6_outputs(5769) <= (layer5_outputs(7556)) xor (layer5_outputs(3632));
    layer6_outputs(5770) <= (layer5_outputs(453)) and not (layer5_outputs(5154));
    layer6_outputs(5771) <= layer5_outputs(685);
    layer6_outputs(5772) <= layer5_outputs(7549);
    layer6_outputs(5773) <= not((layer5_outputs(6080)) xor (layer5_outputs(5145)));
    layer6_outputs(5774) <= (layer5_outputs(1385)) xor (layer5_outputs(4634));
    layer6_outputs(5775) <= not(layer5_outputs(3161));
    layer6_outputs(5776) <= '0';
    layer6_outputs(5777) <= layer5_outputs(2158);
    layer6_outputs(5778) <= not(layer5_outputs(4947));
    layer6_outputs(5779) <= layer5_outputs(3574);
    layer6_outputs(5780) <= layer5_outputs(333);
    layer6_outputs(5781) <= not((layer5_outputs(5808)) xor (layer5_outputs(1696)));
    layer6_outputs(5782) <= '1';
    layer6_outputs(5783) <= (layer5_outputs(6405)) xor (layer5_outputs(416));
    layer6_outputs(5784) <= not((layer5_outputs(397)) xor (layer5_outputs(1310)));
    layer6_outputs(5785) <= layer5_outputs(898);
    layer6_outputs(5786) <= (layer5_outputs(7008)) or (layer5_outputs(4994));
    layer6_outputs(5787) <= (layer5_outputs(2070)) xor (layer5_outputs(3841));
    layer6_outputs(5788) <= layer5_outputs(3381);
    layer6_outputs(5789) <= (layer5_outputs(7190)) xor (layer5_outputs(4855));
    layer6_outputs(5790) <= not(layer5_outputs(4125));
    layer6_outputs(5791) <= not(layer5_outputs(2439));
    layer6_outputs(5792) <= layer5_outputs(5710);
    layer6_outputs(5793) <= not((layer5_outputs(6875)) xor (layer5_outputs(5248)));
    layer6_outputs(5794) <= (layer5_outputs(471)) and (layer5_outputs(5868));
    layer6_outputs(5795) <= not(layer5_outputs(3725));
    layer6_outputs(5796) <= (layer5_outputs(6969)) and (layer5_outputs(771));
    layer6_outputs(5797) <= (layer5_outputs(6134)) and not (layer5_outputs(1127));
    layer6_outputs(5798) <= layer5_outputs(7211);
    layer6_outputs(5799) <= layer5_outputs(1739);
    layer6_outputs(5800) <= not(layer5_outputs(1223)) or (layer5_outputs(4311));
    layer6_outputs(5801) <= not(layer5_outputs(1594));
    layer6_outputs(5802) <= (layer5_outputs(1551)) or (layer5_outputs(6061));
    layer6_outputs(5803) <= layer5_outputs(1332);
    layer6_outputs(5804) <= not(layer5_outputs(5004)) or (layer5_outputs(6082));
    layer6_outputs(5805) <= not(layer5_outputs(223));
    layer6_outputs(5806) <= not((layer5_outputs(4013)) and (layer5_outputs(4738)));
    layer6_outputs(5807) <= (layer5_outputs(3443)) or (layer5_outputs(584));
    layer6_outputs(5808) <= (layer5_outputs(7031)) and not (layer5_outputs(854));
    layer6_outputs(5809) <= layer5_outputs(2245);
    layer6_outputs(5810) <= not(layer5_outputs(3062)) or (layer5_outputs(2219));
    layer6_outputs(5811) <= layer5_outputs(3973);
    layer6_outputs(5812) <= not((layer5_outputs(3817)) xor (layer5_outputs(4681)));
    layer6_outputs(5813) <= (layer5_outputs(689)) xor (layer5_outputs(6945));
    layer6_outputs(5814) <= not(layer5_outputs(146));
    layer6_outputs(5815) <= not(layer5_outputs(7397)) or (layer5_outputs(5933));
    layer6_outputs(5816) <= layer5_outputs(348);
    layer6_outputs(5817) <= (layer5_outputs(5494)) and not (layer5_outputs(6610));
    layer6_outputs(5818) <= not(layer5_outputs(4102));
    layer6_outputs(5819) <= not((layer5_outputs(4663)) xor (layer5_outputs(3636)));
    layer6_outputs(5820) <= not((layer5_outputs(3358)) or (layer5_outputs(6974)));
    layer6_outputs(5821) <= (layer5_outputs(1496)) and not (layer5_outputs(2451));
    layer6_outputs(5822) <= layer5_outputs(6346);
    layer6_outputs(5823) <= not(layer5_outputs(1930));
    layer6_outputs(5824) <= not(layer5_outputs(1998)) or (layer5_outputs(1867));
    layer6_outputs(5825) <= not((layer5_outputs(734)) and (layer5_outputs(243)));
    layer6_outputs(5826) <= (layer5_outputs(3582)) or (layer5_outputs(6630));
    layer6_outputs(5827) <= layer5_outputs(2561);
    layer6_outputs(5828) <= not(layer5_outputs(6355));
    layer6_outputs(5829) <= layer5_outputs(5785);
    layer6_outputs(5830) <= not((layer5_outputs(2748)) and (layer5_outputs(4233)));
    layer6_outputs(5831) <= not((layer5_outputs(855)) and (layer5_outputs(7645)));
    layer6_outputs(5832) <= layer5_outputs(3428);
    layer6_outputs(5833) <= layer5_outputs(7272);
    layer6_outputs(5834) <= layer5_outputs(1565);
    layer6_outputs(5835) <= (layer5_outputs(6293)) and not (layer5_outputs(6455));
    layer6_outputs(5836) <= not(layer5_outputs(954)) or (layer5_outputs(3960));
    layer6_outputs(5837) <= layer5_outputs(6158);
    layer6_outputs(5838) <= (layer5_outputs(7147)) and (layer5_outputs(6693));
    layer6_outputs(5839) <= layer5_outputs(4755);
    layer6_outputs(5840) <= not(layer5_outputs(1550)) or (layer5_outputs(6774));
    layer6_outputs(5841) <= not(layer5_outputs(2667));
    layer6_outputs(5842) <= not(layer5_outputs(4835));
    layer6_outputs(5843) <= not(layer5_outputs(4661));
    layer6_outputs(5844) <= not((layer5_outputs(2265)) xor (layer5_outputs(4308)));
    layer6_outputs(5845) <= not(layer5_outputs(1043));
    layer6_outputs(5846) <= layer5_outputs(2540);
    layer6_outputs(5847) <= (layer5_outputs(2227)) xor (layer5_outputs(3944));
    layer6_outputs(5848) <= (layer5_outputs(2993)) and not (layer5_outputs(3462));
    layer6_outputs(5849) <= not(layer5_outputs(1237)) or (layer5_outputs(4126));
    layer6_outputs(5850) <= not(layer5_outputs(87));
    layer6_outputs(5851) <= (layer5_outputs(4145)) and not (layer5_outputs(3308));
    layer6_outputs(5852) <= layer5_outputs(3654);
    layer6_outputs(5853) <= layer5_outputs(3541);
    layer6_outputs(5854) <= not(layer5_outputs(249));
    layer6_outputs(5855) <= layer5_outputs(6376);
    layer6_outputs(5856) <= layer5_outputs(3158);
    layer6_outputs(5857) <= not(layer5_outputs(125));
    layer6_outputs(5858) <= layer5_outputs(142);
    layer6_outputs(5859) <= layer5_outputs(2040);
    layer6_outputs(5860) <= layer5_outputs(6699);
    layer6_outputs(5861) <= not(layer5_outputs(98)) or (layer5_outputs(5586));
    layer6_outputs(5862) <= not(layer5_outputs(902));
    layer6_outputs(5863) <= not((layer5_outputs(6967)) or (layer5_outputs(7678)));
    layer6_outputs(5864) <= not(layer5_outputs(3183));
    layer6_outputs(5865) <= layer5_outputs(5059);
    layer6_outputs(5866) <= layer5_outputs(3897);
    layer6_outputs(5867) <= layer5_outputs(7490);
    layer6_outputs(5868) <= not((layer5_outputs(3929)) xor (layer5_outputs(3720)));
    layer6_outputs(5869) <= layer5_outputs(167);
    layer6_outputs(5870) <= not(layer5_outputs(1651)) or (layer5_outputs(1477));
    layer6_outputs(5871) <= not(layer5_outputs(2790)) or (layer5_outputs(3820));
    layer6_outputs(5872) <= not(layer5_outputs(7636));
    layer6_outputs(5873) <= (layer5_outputs(1522)) xor (layer5_outputs(303));
    layer6_outputs(5874) <= layer5_outputs(5503);
    layer6_outputs(5875) <= not(layer5_outputs(5856));
    layer6_outputs(5876) <= not(layer5_outputs(3943));
    layer6_outputs(5877) <= (layer5_outputs(6126)) xor (layer5_outputs(5431));
    layer6_outputs(5878) <= not(layer5_outputs(4716));
    layer6_outputs(5879) <= not(layer5_outputs(3169)) or (layer5_outputs(5263));
    layer6_outputs(5880) <= (layer5_outputs(1589)) and (layer5_outputs(5860));
    layer6_outputs(5881) <= not(layer5_outputs(5947));
    layer6_outputs(5882) <= layer5_outputs(2229);
    layer6_outputs(5883) <= layer5_outputs(620);
    layer6_outputs(5884) <= not((layer5_outputs(7048)) and (layer5_outputs(2435)));
    layer6_outputs(5885) <= not((layer5_outputs(635)) xor (layer5_outputs(7095)));
    layer6_outputs(5886) <= not(layer5_outputs(4344));
    layer6_outputs(5887) <= '1';
    layer6_outputs(5888) <= not(layer5_outputs(3361));
    layer6_outputs(5889) <= layer5_outputs(4723);
    layer6_outputs(5890) <= not((layer5_outputs(6935)) and (layer5_outputs(448)));
    layer6_outputs(5891) <= layer5_outputs(7268);
    layer6_outputs(5892) <= layer5_outputs(5368);
    layer6_outputs(5893) <= not(layer5_outputs(375));
    layer6_outputs(5894) <= not(layer5_outputs(3693));
    layer6_outputs(5895) <= (layer5_outputs(2586)) xor (layer5_outputs(2222));
    layer6_outputs(5896) <= layer5_outputs(6704);
    layer6_outputs(5897) <= not((layer5_outputs(5445)) xor (layer5_outputs(2843)));
    layer6_outputs(5898) <= layer5_outputs(2203);
    layer6_outputs(5899) <= not(layer5_outputs(4564)) or (layer5_outputs(4769));
    layer6_outputs(5900) <= (layer5_outputs(7517)) and not (layer5_outputs(5913));
    layer6_outputs(5901) <= layer5_outputs(3281);
    layer6_outputs(5902) <= not(layer5_outputs(912));
    layer6_outputs(5903) <= not(layer5_outputs(3655));
    layer6_outputs(5904) <= not(layer5_outputs(4621));
    layer6_outputs(5905) <= layer5_outputs(7474);
    layer6_outputs(5906) <= (layer5_outputs(1900)) xor (layer5_outputs(5911));
    layer6_outputs(5907) <= not(layer5_outputs(3043));
    layer6_outputs(5908) <= not(layer5_outputs(2547));
    layer6_outputs(5909) <= not((layer5_outputs(4287)) xor (layer5_outputs(1813)));
    layer6_outputs(5910) <= layer5_outputs(6558);
    layer6_outputs(5911) <= (layer5_outputs(4804)) or (layer5_outputs(2247));
    layer6_outputs(5912) <= (layer5_outputs(7232)) and (layer5_outputs(5061));
    layer6_outputs(5913) <= not(layer5_outputs(5193));
    layer6_outputs(5914) <= not(layer5_outputs(3934));
    layer6_outputs(5915) <= not(layer5_outputs(2918));
    layer6_outputs(5916) <= layer5_outputs(2688);
    layer6_outputs(5917) <= not(layer5_outputs(5611));
    layer6_outputs(5918) <= not(layer5_outputs(3465));
    layer6_outputs(5919) <= (layer5_outputs(7622)) and not (layer5_outputs(7321));
    layer6_outputs(5920) <= not(layer5_outputs(903));
    layer6_outputs(5921) <= layer5_outputs(1313);
    layer6_outputs(5922) <= not((layer5_outputs(6800)) and (layer5_outputs(6756)));
    layer6_outputs(5923) <= not(layer5_outputs(523));
    layer6_outputs(5924) <= layer5_outputs(4445);
    layer6_outputs(5925) <= layer5_outputs(2234);
    layer6_outputs(5926) <= not((layer5_outputs(4441)) xor (layer5_outputs(5930)));
    layer6_outputs(5927) <= layer5_outputs(6422);
    layer6_outputs(5928) <= not(layer5_outputs(6553)) or (layer5_outputs(4872));
    layer6_outputs(5929) <= layer5_outputs(1397);
    layer6_outputs(5930) <= layer5_outputs(6328);
    layer6_outputs(5931) <= not((layer5_outputs(469)) xor (layer5_outputs(6468)));
    layer6_outputs(5932) <= layer5_outputs(3905);
    layer6_outputs(5933) <= not(layer5_outputs(3232));
    layer6_outputs(5934) <= not(layer5_outputs(4183)) or (layer5_outputs(2421));
    layer6_outputs(5935) <= not((layer5_outputs(3402)) or (layer5_outputs(6056)));
    layer6_outputs(5936) <= not(layer5_outputs(3847));
    layer6_outputs(5937) <= not(layer5_outputs(6017)) or (layer5_outputs(1208));
    layer6_outputs(5938) <= not(layer5_outputs(1185));
    layer6_outputs(5939) <= not(layer5_outputs(3950));
    layer6_outputs(5940) <= layer5_outputs(5644);
    layer6_outputs(5941) <= (layer5_outputs(3767)) xor (layer5_outputs(7659));
    layer6_outputs(5942) <= not(layer5_outputs(528));
    layer6_outputs(5943) <= not((layer5_outputs(4558)) or (layer5_outputs(1873)));
    layer6_outputs(5944) <= not(layer5_outputs(4205));
    layer6_outputs(5945) <= layer5_outputs(1923);
    layer6_outputs(5946) <= not((layer5_outputs(908)) xor (layer5_outputs(496)));
    layer6_outputs(5947) <= (layer5_outputs(361)) xor (layer5_outputs(3013));
    layer6_outputs(5948) <= not(layer5_outputs(3669));
    layer6_outputs(5949) <= (layer5_outputs(2775)) xor (layer5_outputs(3398));
    layer6_outputs(5950) <= not(layer5_outputs(148));
    layer6_outputs(5951) <= (layer5_outputs(6694)) xor (layer5_outputs(3331));
    layer6_outputs(5952) <= not(layer5_outputs(3765));
    layer6_outputs(5953) <= (layer5_outputs(5640)) and not (layer5_outputs(3529));
    layer6_outputs(5954) <= layer5_outputs(2052);
    layer6_outputs(5955) <= layer5_outputs(4602);
    layer6_outputs(5956) <= layer5_outputs(5401);
    layer6_outputs(5957) <= not(layer5_outputs(3019));
    layer6_outputs(5958) <= not(layer5_outputs(4612));
    layer6_outputs(5959) <= not((layer5_outputs(5150)) or (layer5_outputs(5154)));
    layer6_outputs(5960) <= not((layer5_outputs(6729)) and (layer5_outputs(5815)));
    layer6_outputs(5961) <= layer5_outputs(291);
    layer6_outputs(5962) <= (layer5_outputs(7360)) xor (layer5_outputs(2313));
    layer6_outputs(5963) <= not((layer5_outputs(4782)) and (layer5_outputs(5649)));
    layer6_outputs(5964) <= (layer5_outputs(3093)) and not (layer5_outputs(4717));
    layer6_outputs(5965) <= not(layer5_outputs(3233));
    layer6_outputs(5966) <= layer5_outputs(3378);
    layer6_outputs(5967) <= not((layer5_outputs(4373)) xor (layer5_outputs(6616)));
    layer6_outputs(5968) <= not(layer5_outputs(6223));
    layer6_outputs(5969) <= not((layer5_outputs(1605)) xor (layer5_outputs(3129)));
    layer6_outputs(5970) <= not(layer5_outputs(4669));
    layer6_outputs(5971) <= not(layer5_outputs(2296));
    layer6_outputs(5972) <= not(layer5_outputs(4352));
    layer6_outputs(5973) <= layer5_outputs(7197);
    layer6_outputs(5974) <= (layer5_outputs(2785)) and not (layer5_outputs(919));
    layer6_outputs(5975) <= not(layer5_outputs(4392));
    layer6_outputs(5976) <= not(layer5_outputs(2583)) or (layer5_outputs(4840));
    layer6_outputs(5977) <= not((layer5_outputs(6962)) or (layer5_outputs(4461)));
    layer6_outputs(5978) <= layer5_outputs(3);
    layer6_outputs(5979) <= (layer5_outputs(2177)) and (layer5_outputs(4241));
    layer6_outputs(5980) <= '0';
    layer6_outputs(5981) <= layer5_outputs(5071);
    layer6_outputs(5982) <= '1';
    layer6_outputs(5983) <= not(layer5_outputs(7058));
    layer6_outputs(5984) <= (layer5_outputs(5978)) and (layer5_outputs(536));
    layer6_outputs(5985) <= (layer5_outputs(769)) and not (layer5_outputs(5683));
    layer6_outputs(5986) <= (layer5_outputs(5351)) xor (layer5_outputs(4853));
    layer6_outputs(5987) <= (layer5_outputs(5291)) or (layer5_outputs(2516));
    layer6_outputs(5988) <= layer5_outputs(1190);
    layer6_outputs(5989) <= not(layer5_outputs(1615));
    layer6_outputs(5990) <= not(layer5_outputs(4763));
    layer6_outputs(5991) <= not((layer5_outputs(6438)) xor (layer5_outputs(6215)));
    layer6_outputs(5992) <= (layer5_outputs(7309)) and (layer5_outputs(3334));
    layer6_outputs(5993) <= layer5_outputs(7679);
    layer6_outputs(5994) <= layer5_outputs(3467);
    layer6_outputs(5995) <= (layer5_outputs(5783)) or (layer5_outputs(5903));
    layer6_outputs(5996) <= not(layer5_outputs(2425));
    layer6_outputs(5997) <= layer5_outputs(4273);
    layer6_outputs(5998) <= (layer5_outputs(3251)) or (layer5_outputs(7585));
    layer6_outputs(5999) <= (layer5_outputs(1625)) and not (layer5_outputs(1645));
    layer6_outputs(6000) <= not(layer5_outputs(1993));
    layer6_outputs(6001) <= layer5_outputs(470);
    layer6_outputs(6002) <= not((layer5_outputs(7051)) xor (layer5_outputs(3876)));
    layer6_outputs(6003) <= layer5_outputs(1458);
    layer6_outputs(6004) <= not((layer5_outputs(972)) xor (layer5_outputs(6012)));
    layer6_outputs(6005) <= layer5_outputs(7044);
    layer6_outputs(6006) <= (layer5_outputs(7021)) xor (layer5_outputs(7351));
    layer6_outputs(6007) <= layer5_outputs(1263);
    layer6_outputs(6008) <= not(layer5_outputs(4065));
    layer6_outputs(6009) <= layer5_outputs(5411);
    layer6_outputs(6010) <= (layer5_outputs(4716)) and (layer5_outputs(6031));
    layer6_outputs(6011) <= (layer5_outputs(1973)) and not (layer5_outputs(6432));
    layer6_outputs(6012) <= not((layer5_outputs(544)) xor (layer5_outputs(2851)));
    layer6_outputs(6013) <= not(layer5_outputs(215)) or (layer5_outputs(3832));
    layer6_outputs(6014) <= layer5_outputs(4951);
    layer6_outputs(6015) <= layer5_outputs(7621);
    layer6_outputs(6016) <= (layer5_outputs(5040)) and (layer5_outputs(7326));
    layer6_outputs(6017) <= not(layer5_outputs(2029));
    layer6_outputs(6018) <= layer5_outputs(2092);
    layer6_outputs(6019) <= not((layer5_outputs(5725)) xor (layer5_outputs(547)));
    layer6_outputs(6020) <= layer5_outputs(6708);
    layer6_outputs(6021) <= not(layer5_outputs(3338)) or (layer5_outputs(436));
    layer6_outputs(6022) <= layer5_outputs(387);
    layer6_outputs(6023) <= not(layer5_outputs(3542));
    layer6_outputs(6024) <= not(layer5_outputs(4792));
    layer6_outputs(6025) <= not((layer5_outputs(6120)) or (layer5_outputs(2530)));
    layer6_outputs(6026) <= (layer5_outputs(1116)) or (layer5_outputs(6308));
    layer6_outputs(6027) <= layer5_outputs(21);
    layer6_outputs(6028) <= not(layer5_outputs(6705));
    layer6_outputs(6029) <= not(layer5_outputs(6933)) or (layer5_outputs(6519));
    layer6_outputs(6030) <= (layer5_outputs(1851)) xor (layer5_outputs(5309));
    layer6_outputs(6031) <= not(layer5_outputs(6927));
    layer6_outputs(6032) <= (layer5_outputs(5502)) xor (layer5_outputs(7417));
    layer6_outputs(6033) <= (layer5_outputs(1294)) and (layer5_outputs(3134));
    layer6_outputs(6034) <= not(layer5_outputs(7167));
    layer6_outputs(6035) <= not((layer5_outputs(3509)) or (layer5_outputs(6559)));
    layer6_outputs(6036) <= layer5_outputs(1866);
    layer6_outputs(6037) <= not(layer5_outputs(2715));
    layer6_outputs(6038) <= not((layer5_outputs(1622)) xor (layer5_outputs(4415)));
    layer6_outputs(6039) <= not(layer5_outputs(1724)) or (layer5_outputs(4686));
    layer6_outputs(6040) <= layer5_outputs(46);
    layer6_outputs(6041) <= layer5_outputs(3878);
    layer6_outputs(6042) <= not(layer5_outputs(1683)) or (layer5_outputs(7015));
    layer6_outputs(6043) <= not(layer5_outputs(4086));
    layer6_outputs(6044) <= not((layer5_outputs(4265)) and (layer5_outputs(2384)));
    layer6_outputs(6045) <= '0';
    layer6_outputs(6046) <= not(layer5_outputs(1240));
    layer6_outputs(6047) <= layer5_outputs(986);
    layer6_outputs(6048) <= (layer5_outputs(842)) and not (layer5_outputs(3592));
    layer6_outputs(6049) <= layer5_outputs(5343);
    layer6_outputs(6050) <= layer5_outputs(87);
    layer6_outputs(6051) <= not(layer5_outputs(2271));
    layer6_outputs(6052) <= not(layer5_outputs(5769));
    layer6_outputs(6053) <= not(layer5_outputs(7433));
    layer6_outputs(6054) <= not(layer5_outputs(2352));
    layer6_outputs(6055) <= layer5_outputs(2899);
    layer6_outputs(6056) <= (layer5_outputs(1717)) xor (layer5_outputs(3703));
    layer6_outputs(6057) <= (layer5_outputs(689)) and not (layer5_outputs(2678));
    layer6_outputs(6058) <= not((layer5_outputs(1638)) or (layer5_outputs(2093)));
    layer6_outputs(6059) <= layer5_outputs(6176);
    layer6_outputs(6060) <= not((layer5_outputs(4158)) xor (layer5_outputs(6607)));
    layer6_outputs(6061) <= layer5_outputs(818);
    layer6_outputs(6062) <= layer5_outputs(1780);
    layer6_outputs(6063) <= layer5_outputs(1427);
    layer6_outputs(6064) <= layer5_outputs(6566);
    layer6_outputs(6065) <= not(layer5_outputs(2128));
    layer6_outputs(6066) <= not((layer5_outputs(85)) xor (layer5_outputs(5527)));
    layer6_outputs(6067) <= layer5_outputs(7349);
    layer6_outputs(6068) <= not(layer5_outputs(1778)) or (layer5_outputs(5063));
    layer6_outputs(6069) <= (layer5_outputs(4951)) xor (layer5_outputs(4637));
    layer6_outputs(6070) <= not((layer5_outputs(5977)) and (layer5_outputs(6511)));
    layer6_outputs(6071) <= not(layer5_outputs(7489));
    layer6_outputs(6072) <= layer5_outputs(6904);
    layer6_outputs(6073) <= layer5_outputs(2358);
    layer6_outputs(6074) <= layer5_outputs(6847);
    layer6_outputs(6075) <= not(layer5_outputs(1831));
    layer6_outputs(6076) <= layer5_outputs(2438);
    layer6_outputs(6077) <= (layer5_outputs(2519)) xor (layer5_outputs(6724));
    layer6_outputs(6078) <= not(layer5_outputs(1347));
    layer6_outputs(6079) <= (layer5_outputs(4933)) and not (layer5_outputs(3910));
    layer6_outputs(6080) <= layer5_outputs(195);
    layer6_outputs(6081) <= not((layer5_outputs(7669)) and (layer5_outputs(7631)));
    layer6_outputs(6082) <= not((layer5_outputs(6451)) and (layer5_outputs(1879)));
    layer6_outputs(6083) <= (layer5_outputs(7388)) xor (layer5_outputs(4421));
    layer6_outputs(6084) <= not(layer5_outputs(411));
    layer6_outputs(6085) <= not((layer5_outputs(2088)) and (layer5_outputs(1850)));
    layer6_outputs(6086) <= layer5_outputs(7599);
    layer6_outputs(6087) <= layer5_outputs(7406);
    layer6_outputs(6088) <= not((layer5_outputs(939)) xor (layer5_outputs(4892)));
    layer6_outputs(6089) <= layer5_outputs(1219);
    layer6_outputs(6090) <= not(layer5_outputs(6754));
    layer6_outputs(6091) <= not(layer5_outputs(2700));
    layer6_outputs(6092) <= layer5_outputs(1389);
    layer6_outputs(6093) <= layer5_outputs(1653);
    layer6_outputs(6094) <= not((layer5_outputs(1747)) xor (layer5_outputs(4361)));
    layer6_outputs(6095) <= not(layer5_outputs(4223));
    layer6_outputs(6096) <= '1';
    layer6_outputs(6097) <= (layer5_outputs(2375)) xor (layer5_outputs(5920));
    layer6_outputs(6098) <= layer5_outputs(6008);
    layer6_outputs(6099) <= layer5_outputs(5512);
    layer6_outputs(6100) <= (layer5_outputs(4153)) or (layer5_outputs(2146));
    layer6_outputs(6101) <= not((layer5_outputs(5418)) xor (layer5_outputs(3771)));
    layer6_outputs(6102) <= (layer5_outputs(4225)) or (layer5_outputs(7301));
    layer6_outputs(6103) <= layer5_outputs(775);
    layer6_outputs(6104) <= layer5_outputs(5782);
    layer6_outputs(6105) <= layer5_outputs(7197);
    layer6_outputs(6106) <= (layer5_outputs(179)) and not (layer5_outputs(1532));
    layer6_outputs(6107) <= layer5_outputs(2176);
    layer6_outputs(6108) <= not(layer5_outputs(329));
    layer6_outputs(6109) <= not((layer5_outputs(2366)) or (layer5_outputs(3068)));
    layer6_outputs(6110) <= (layer5_outputs(6976)) and not (layer5_outputs(7281));
    layer6_outputs(6111) <= not(layer5_outputs(2991));
    layer6_outputs(6112) <= not(layer5_outputs(2254));
    layer6_outputs(6113) <= (layer5_outputs(4892)) xor (layer5_outputs(692));
    layer6_outputs(6114) <= layer5_outputs(3801);
    layer6_outputs(6115) <= not(layer5_outputs(556));
    layer6_outputs(6116) <= (layer5_outputs(4807)) or (layer5_outputs(2869));
    layer6_outputs(6117) <= layer5_outputs(4477);
    layer6_outputs(6118) <= not(layer5_outputs(451));
    layer6_outputs(6119) <= not(layer5_outputs(4828));
    layer6_outputs(6120) <= layer5_outputs(2483);
    layer6_outputs(6121) <= not(layer5_outputs(3010));
    layer6_outputs(6122) <= (layer5_outputs(2653)) and not (layer5_outputs(4698));
    layer6_outputs(6123) <= not((layer5_outputs(6899)) and (layer5_outputs(2262)));
    layer6_outputs(6124) <= (layer5_outputs(7602)) and (layer5_outputs(1741));
    layer6_outputs(6125) <= layer5_outputs(1100);
    layer6_outputs(6126) <= not(layer5_outputs(3390)) or (layer5_outputs(4691));
    layer6_outputs(6127) <= '0';
    layer6_outputs(6128) <= (layer5_outputs(4357)) and (layer5_outputs(6160));
    layer6_outputs(6129) <= not(layer5_outputs(2838));
    layer6_outputs(6130) <= not((layer5_outputs(3995)) or (layer5_outputs(1678)));
    layer6_outputs(6131) <= (layer5_outputs(4046)) and not (layer5_outputs(5839));
    layer6_outputs(6132) <= not((layer5_outputs(4764)) xor (layer5_outputs(1355)));
    layer6_outputs(6133) <= (layer5_outputs(929)) xor (layer5_outputs(4547));
    layer6_outputs(6134) <= layer5_outputs(4459);
    layer6_outputs(6135) <= (layer5_outputs(2318)) and (layer5_outputs(1029));
    layer6_outputs(6136) <= not(layer5_outputs(1307));
    layer6_outputs(6137) <= (layer5_outputs(7661)) and (layer5_outputs(3719));
    layer6_outputs(6138) <= layer5_outputs(2205);
    layer6_outputs(6139) <= not(layer5_outputs(54)) or (layer5_outputs(548));
    layer6_outputs(6140) <= not((layer5_outputs(4282)) xor (layer5_outputs(4984)));
    layer6_outputs(6141) <= layer5_outputs(5330);
    layer6_outputs(6142) <= layer5_outputs(327);
    layer6_outputs(6143) <= not(layer5_outputs(2277));
    layer6_outputs(6144) <= layer5_outputs(4255);
    layer6_outputs(6145) <= not((layer5_outputs(4829)) xor (layer5_outputs(373)));
    layer6_outputs(6146) <= (layer5_outputs(6545)) or (layer5_outputs(82));
    layer6_outputs(6147) <= not(layer5_outputs(526));
    layer6_outputs(6148) <= not(layer5_outputs(6446));
    layer6_outputs(6149) <= not(layer5_outputs(3378));
    layer6_outputs(6150) <= not(layer5_outputs(4582)) or (layer5_outputs(1929));
    layer6_outputs(6151) <= '1';
    layer6_outputs(6152) <= (layer5_outputs(3021)) xor (layer5_outputs(7655));
    layer6_outputs(6153) <= not(layer5_outputs(480));
    layer6_outputs(6154) <= not((layer5_outputs(7451)) and (layer5_outputs(6878)));
    layer6_outputs(6155) <= not(layer5_outputs(2348));
    layer6_outputs(6156) <= not((layer5_outputs(5865)) xor (layer5_outputs(3216)));
    layer6_outputs(6157) <= layer5_outputs(3055);
    layer6_outputs(6158) <= (layer5_outputs(243)) xor (layer5_outputs(2711));
    layer6_outputs(6159) <= layer5_outputs(7247);
    layer6_outputs(6160) <= not(layer5_outputs(3909));
    layer6_outputs(6161) <= layer5_outputs(6651);
    layer6_outputs(6162) <= layer5_outputs(5831);
    layer6_outputs(6163) <= not((layer5_outputs(1731)) xor (layer5_outputs(230)));
    layer6_outputs(6164) <= layer5_outputs(676);
    layer6_outputs(6165) <= not((layer5_outputs(3696)) and (layer5_outputs(4305)));
    layer6_outputs(6166) <= not(layer5_outputs(136));
    layer6_outputs(6167) <= layer5_outputs(2081);
    layer6_outputs(6168) <= (layer5_outputs(1987)) or (layer5_outputs(1012));
    layer6_outputs(6169) <= not(layer5_outputs(4685));
    layer6_outputs(6170) <= (layer5_outputs(2206)) and (layer5_outputs(2588));
    layer6_outputs(6171) <= not(layer5_outputs(4667)) or (layer5_outputs(6914));
    layer6_outputs(6172) <= not(layer5_outputs(1138));
    layer6_outputs(6173) <= not(layer5_outputs(1493));
    layer6_outputs(6174) <= (layer5_outputs(6186)) or (layer5_outputs(607));
    layer6_outputs(6175) <= not(layer5_outputs(5275)) or (layer5_outputs(1012));
    layer6_outputs(6176) <= not(layer5_outputs(6932));
    layer6_outputs(6177) <= (layer5_outputs(7391)) xor (layer5_outputs(1002));
    layer6_outputs(6178) <= (layer5_outputs(4122)) or (layer5_outputs(6568));
    layer6_outputs(6179) <= not(layer5_outputs(5786)) or (layer5_outputs(3598));
    layer6_outputs(6180) <= not(layer5_outputs(5932)) or (layer5_outputs(1141));
    layer6_outputs(6181) <= not((layer5_outputs(843)) or (layer5_outputs(480)));
    layer6_outputs(6182) <= not(layer5_outputs(4661));
    layer6_outputs(6183) <= not((layer5_outputs(7329)) xor (layer5_outputs(5447)));
    layer6_outputs(6184) <= not((layer5_outputs(5091)) xor (layer5_outputs(303)));
    layer6_outputs(6185) <= layer5_outputs(4266);
    layer6_outputs(6186) <= not(layer5_outputs(6475));
    layer6_outputs(6187) <= not(layer5_outputs(4674));
    layer6_outputs(6188) <= layer5_outputs(5788);
    layer6_outputs(6189) <= layer5_outputs(4053);
    layer6_outputs(6190) <= not(layer5_outputs(1509)) or (layer5_outputs(1462));
    layer6_outputs(6191) <= not(layer5_outputs(3469));
    layer6_outputs(6192) <= layer5_outputs(2459);
    layer6_outputs(6193) <= not(layer5_outputs(1235));
    layer6_outputs(6194) <= layer5_outputs(6233);
    layer6_outputs(6195) <= not(layer5_outputs(1533));
    layer6_outputs(6196) <= (layer5_outputs(1041)) and (layer5_outputs(673));
    layer6_outputs(6197) <= not((layer5_outputs(6218)) xor (layer5_outputs(824)));
    layer6_outputs(6198) <= not(layer5_outputs(5475)) or (layer5_outputs(5784));
    layer6_outputs(6199) <= not((layer5_outputs(2706)) and (layer5_outputs(5845)));
    layer6_outputs(6200) <= (layer5_outputs(7015)) and not (layer5_outputs(1953));
    layer6_outputs(6201) <= not(layer5_outputs(3333)) or (layer5_outputs(6618));
    layer6_outputs(6202) <= not(layer5_outputs(5446));
    layer6_outputs(6203) <= layer5_outputs(2252);
    layer6_outputs(6204) <= not(layer5_outputs(7353));
    layer6_outputs(6205) <= layer5_outputs(3081);
    layer6_outputs(6206) <= layer5_outputs(6236);
    layer6_outputs(6207) <= not((layer5_outputs(927)) xor (layer5_outputs(103)));
    layer6_outputs(6208) <= not((layer5_outputs(1216)) and (layer5_outputs(6124)));
    layer6_outputs(6209) <= (layer5_outputs(3629)) and not (layer5_outputs(5365));
    layer6_outputs(6210) <= layer5_outputs(6025);
    layer6_outputs(6211) <= not(layer5_outputs(3463));
    layer6_outputs(6212) <= (layer5_outputs(2602)) and not (layer5_outputs(6202));
    layer6_outputs(6213) <= (layer5_outputs(2375)) and (layer5_outputs(6475));
    layer6_outputs(6214) <= layer5_outputs(3831);
    layer6_outputs(6215) <= not(layer5_outputs(1973));
    layer6_outputs(6216) <= layer5_outputs(3453);
    layer6_outputs(6217) <= (layer5_outputs(5409)) or (layer5_outputs(2875));
    layer6_outputs(6218) <= not(layer5_outputs(2463));
    layer6_outputs(6219) <= layer5_outputs(4467);
    layer6_outputs(6220) <= layer5_outputs(1803);
    layer6_outputs(6221) <= layer5_outputs(1631);
    layer6_outputs(6222) <= not(layer5_outputs(6582)) or (layer5_outputs(7293));
    layer6_outputs(6223) <= (layer5_outputs(3397)) and not (layer5_outputs(2446));
    layer6_outputs(6224) <= layer5_outputs(2487);
    layer6_outputs(6225) <= not(layer5_outputs(2346)) or (layer5_outputs(2358));
    layer6_outputs(6226) <= not(layer5_outputs(371)) or (layer5_outputs(3363));
    layer6_outputs(6227) <= (layer5_outputs(650)) xor (layer5_outputs(4379));
    layer6_outputs(6228) <= (layer5_outputs(3967)) and not (layer5_outputs(3839));
    layer6_outputs(6229) <= not(layer5_outputs(2742)) or (layer5_outputs(2648));
    layer6_outputs(6230) <= layer5_outputs(7162);
    layer6_outputs(6231) <= (layer5_outputs(3267)) and not (layer5_outputs(447));
    layer6_outputs(6232) <= (layer5_outputs(6211)) or (layer5_outputs(1502));
    layer6_outputs(6233) <= (layer5_outputs(3698)) xor (layer5_outputs(3047));
    layer6_outputs(6234) <= not(layer5_outputs(568));
    layer6_outputs(6235) <= not(layer5_outputs(2650));
    layer6_outputs(6236) <= layer5_outputs(2231);
    layer6_outputs(6237) <= not(layer5_outputs(7578));
    layer6_outputs(6238) <= layer5_outputs(5247);
    layer6_outputs(6239) <= layer5_outputs(99);
    layer6_outputs(6240) <= layer5_outputs(5437);
    layer6_outputs(6241) <= not(layer5_outputs(105));
    layer6_outputs(6242) <= layer5_outputs(1560);
    layer6_outputs(6243) <= layer5_outputs(3609);
    layer6_outputs(6244) <= (layer5_outputs(5749)) or (layer5_outputs(1273));
    layer6_outputs(6245) <= (layer5_outputs(2385)) and not (layer5_outputs(2835));
    layer6_outputs(6246) <= not((layer5_outputs(4554)) xor (layer5_outputs(1144)));
    layer6_outputs(6247) <= (layer5_outputs(1146)) xor (layer5_outputs(5748));
    layer6_outputs(6248) <= not(layer5_outputs(3727)) or (layer5_outputs(6791));
    layer6_outputs(6249) <= (layer5_outputs(2986)) xor (layer5_outputs(7540));
    layer6_outputs(6250) <= layer5_outputs(1900);
    layer6_outputs(6251) <= (layer5_outputs(5201)) and not (layer5_outputs(2833));
    layer6_outputs(6252) <= not(layer5_outputs(4675));
    layer6_outputs(6253) <= layer5_outputs(1667);
    layer6_outputs(6254) <= not(layer5_outputs(5322));
    layer6_outputs(6255) <= (layer5_outputs(60)) and (layer5_outputs(3919));
    layer6_outputs(6256) <= not(layer5_outputs(949));
    layer6_outputs(6257) <= layer5_outputs(663);
    layer6_outputs(6258) <= (layer5_outputs(2124)) xor (layer5_outputs(6692));
    layer6_outputs(6259) <= layer5_outputs(3313);
    layer6_outputs(6260) <= layer5_outputs(1940);
    layer6_outputs(6261) <= not(layer5_outputs(4063));
    layer6_outputs(6262) <= (layer5_outputs(1401)) and not (layer5_outputs(312));
    layer6_outputs(6263) <= not((layer5_outputs(1573)) xor (layer5_outputs(2540)));
    layer6_outputs(6264) <= '1';
    layer6_outputs(6265) <= (layer5_outputs(1326)) and (layer5_outputs(5642));
    layer6_outputs(6266) <= not(layer5_outputs(2692)) or (layer5_outputs(3208));
    layer6_outputs(6267) <= layer5_outputs(4310);
    layer6_outputs(6268) <= (layer5_outputs(4511)) xor (layer5_outputs(2496));
    layer6_outputs(6269) <= not(layer5_outputs(2629)) or (layer5_outputs(2225));
    layer6_outputs(6270) <= not(layer5_outputs(3200));
    layer6_outputs(6271) <= not((layer5_outputs(675)) xor (layer5_outputs(1434)));
    layer6_outputs(6272) <= (layer5_outputs(1262)) and not (layer5_outputs(4418));
    layer6_outputs(6273) <= layer5_outputs(1159);
    layer6_outputs(6274) <= not(layer5_outputs(4894));
    layer6_outputs(6275) <= not(layer5_outputs(4941)) or (layer5_outputs(6175));
    layer6_outputs(6276) <= not(layer5_outputs(4900));
    layer6_outputs(6277) <= not(layer5_outputs(2452));
    layer6_outputs(6278) <= not(layer5_outputs(3241));
    layer6_outputs(6279) <= not(layer5_outputs(534)) or (layer5_outputs(7075));
    layer6_outputs(6280) <= not(layer5_outputs(7369)) or (layer5_outputs(5198));
    layer6_outputs(6281) <= not(layer5_outputs(6530)) or (layer5_outputs(1588));
    layer6_outputs(6282) <= (layer5_outputs(2856)) and not (layer5_outputs(6187));
    layer6_outputs(6283) <= not(layer5_outputs(350));
    layer6_outputs(6284) <= (layer5_outputs(7596)) and not (layer5_outputs(6722));
    layer6_outputs(6285) <= layer5_outputs(6068);
    layer6_outputs(6286) <= not(layer5_outputs(2059));
    layer6_outputs(6287) <= (layer5_outputs(7383)) and not (layer5_outputs(324));
    layer6_outputs(6288) <= (layer5_outputs(1452)) xor (layer5_outputs(4536));
    layer6_outputs(6289) <= not(layer5_outputs(3169)) or (layer5_outputs(4271));
    layer6_outputs(6290) <= not(layer5_outputs(6340));
    layer6_outputs(6291) <= (layer5_outputs(6156)) and not (layer5_outputs(1935));
    layer6_outputs(6292) <= (layer5_outputs(4244)) or (layer5_outputs(3608));
    layer6_outputs(6293) <= not(layer5_outputs(3325));
    layer6_outputs(6294) <= (layer5_outputs(2470)) or (layer5_outputs(6600));
    layer6_outputs(6295) <= layer5_outputs(3284);
    layer6_outputs(6296) <= layer5_outputs(326);
    layer6_outputs(6297) <= not(layer5_outputs(1931));
    layer6_outputs(6298) <= not(layer5_outputs(5406));
    layer6_outputs(6299) <= (layer5_outputs(3180)) and not (layer5_outputs(6259));
    layer6_outputs(6300) <= not(layer5_outputs(3953));
    layer6_outputs(6301) <= (layer5_outputs(1123)) xor (layer5_outputs(4985));
    layer6_outputs(6302) <= layer5_outputs(3447);
    layer6_outputs(6303) <= (layer5_outputs(4419)) xor (layer5_outputs(2043));
    layer6_outputs(6304) <= not(layer5_outputs(107));
    layer6_outputs(6305) <= (layer5_outputs(6424)) and not (layer5_outputs(2468));
    layer6_outputs(6306) <= not(layer5_outputs(6127)) or (layer5_outputs(454));
    layer6_outputs(6307) <= not(layer5_outputs(3873));
    layer6_outputs(6308) <= not((layer5_outputs(5442)) xor (layer5_outputs(353)));
    layer6_outputs(6309) <= not(layer5_outputs(6866));
    layer6_outputs(6310) <= not(layer5_outputs(2379));
    layer6_outputs(6311) <= layer5_outputs(6209);
    layer6_outputs(6312) <= layer5_outputs(5891);
    layer6_outputs(6313) <= not((layer5_outputs(5780)) and (layer5_outputs(4180)));
    layer6_outputs(6314) <= '0';
    layer6_outputs(6315) <= layer5_outputs(867);
    layer6_outputs(6316) <= not((layer5_outputs(2208)) xor (layer5_outputs(4119)));
    layer6_outputs(6317) <= layer5_outputs(7496);
    layer6_outputs(6318) <= (layer5_outputs(5973)) or (layer5_outputs(2087));
    layer6_outputs(6319) <= (layer5_outputs(2791)) and not (layer5_outputs(6732));
    layer6_outputs(6320) <= not(layer5_outputs(7566)) or (layer5_outputs(6389));
    layer6_outputs(6321) <= not((layer5_outputs(5994)) xor (layer5_outputs(917)));
    layer6_outputs(6322) <= not(layer5_outputs(3007));
    layer6_outputs(6323) <= (layer5_outputs(4884)) and not (layer5_outputs(5639));
    layer6_outputs(6324) <= layer5_outputs(6262);
    layer6_outputs(6325) <= not(layer5_outputs(3648));
    layer6_outputs(6326) <= not(layer5_outputs(1023));
    layer6_outputs(6327) <= (layer5_outputs(5449)) xor (layer5_outputs(4687));
    layer6_outputs(6328) <= not(layer5_outputs(4224));
    layer6_outputs(6329) <= layer5_outputs(2489);
    layer6_outputs(6330) <= not((layer5_outputs(719)) xor (layer5_outputs(2496)));
    layer6_outputs(6331) <= not(layer5_outputs(485));
    layer6_outputs(6332) <= not((layer5_outputs(3184)) xor (layer5_outputs(3938)));
    layer6_outputs(6333) <= not(layer5_outputs(3403)) or (layer5_outputs(7611));
    layer6_outputs(6334) <= (layer5_outputs(6526)) and not (layer5_outputs(6697));
    layer6_outputs(6335) <= not(layer5_outputs(2830)) or (layer5_outputs(5869));
    layer6_outputs(6336) <= not(layer5_outputs(2712));
    layer6_outputs(6337) <= layer5_outputs(3847);
    layer6_outputs(6338) <= layer5_outputs(7047);
    layer6_outputs(6339) <= not(layer5_outputs(3600));
    layer6_outputs(6340) <= layer5_outputs(3988);
    layer6_outputs(6341) <= not((layer5_outputs(7244)) and (layer5_outputs(6590)));
    layer6_outputs(6342) <= not(layer5_outputs(2008));
    layer6_outputs(6343) <= layer5_outputs(5297);
    layer6_outputs(6344) <= not((layer5_outputs(2657)) xor (layer5_outputs(7433)));
    layer6_outputs(6345) <= not(layer5_outputs(6615)) or (layer5_outputs(4725));
    layer6_outputs(6346) <= layer5_outputs(6286);
    layer6_outputs(6347) <= not((layer5_outputs(6317)) xor (layer5_outputs(6014)));
    layer6_outputs(6348) <= layer5_outputs(6053);
    layer6_outputs(6349) <= not(layer5_outputs(2479));
    layer6_outputs(6350) <= layer5_outputs(5569);
    layer6_outputs(6351) <= not(layer5_outputs(7241));
    layer6_outputs(6352) <= not(layer5_outputs(6595));
    layer6_outputs(6353) <= layer5_outputs(510);
    layer6_outputs(6354) <= not((layer5_outputs(4882)) xor (layer5_outputs(7546)));
    layer6_outputs(6355) <= (layer5_outputs(6080)) xor (layer5_outputs(7126));
    layer6_outputs(6356) <= not(layer5_outputs(4110));
    layer6_outputs(6357) <= (layer5_outputs(6525)) xor (layer5_outputs(5629));
    layer6_outputs(6358) <= not(layer5_outputs(4889));
    layer6_outputs(6359) <= layer5_outputs(4771);
    layer6_outputs(6360) <= layer5_outputs(1191);
    layer6_outputs(6361) <= not((layer5_outputs(1075)) xor (layer5_outputs(1463)));
    layer6_outputs(6362) <= (layer5_outputs(2648)) xor (layer5_outputs(2084));
    layer6_outputs(6363) <= (layer5_outputs(5372)) xor (layer5_outputs(3420));
    layer6_outputs(6364) <= not((layer5_outputs(1623)) and (layer5_outputs(724)));
    layer6_outputs(6365) <= not((layer5_outputs(843)) xor (layer5_outputs(735)));
    layer6_outputs(6366) <= layer5_outputs(5674);
    layer6_outputs(6367) <= not(layer5_outputs(7387));
    layer6_outputs(6368) <= not(layer5_outputs(3486));
    layer6_outputs(6369) <= layer5_outputs(6892);
    layer6_outputs(6370) <= not((layer5_outputs(6702)) or (layer5_outputs(3874)));
    layer6_outputs(6371) <= '0';
    layer6_outputs(6372) <= (layer5_outputs(232)) and not (layer5_outputs(4533));
    layer6_outputs(6373) <= layer5_outputs(4190);
    layer6_outputs(6374) <= layer5_outputs(262);
    layer6_outputs(6375) <= not(layer5_outputs(2623));
    layer6_outputs(6376) <= (layer5_outputs(5555)) xor (layer5_outputs(292));
    layer6_outputs(6377) <= '1';
    layer6_outputs(6378) <= not((layer5_outputs(3833)) xor (layer5_outputs(7041)));
    layer6_outputs(6379) <= not(layer5_outputs(1639));
    layer6_outputs(6380) <= not(layer5_outputs(1354)) or (layer5_outputs(2551));
    layer6_outputs(6381) <= not(layer5_outputs(1700));
    layer6_outputs(6382) <= not(layer5_outputs(4192));
    layer6_outputs(6383) <= not(layer5_outputs(429));
    layer6_outputs(6384) <= not(layer5_outputs(657));
    layer6_outputs(6385) <= not(layer5_outputs(838)) or (layer5_outputs(1584));
    layer6_outputs(6386) <= not(layer5_outputs(7676)) or (layer5_outputs(3430));
    layer6_outputs(6387) <= (layer5_outputs(3452)) xor (layer5_outputs(1569));
    layer6_outputs(6388) <= not(layer5_outputs(3029));
    layer6_outputs(6389) <= (layer5_outputs(4991)) or (layer5_outputs(3013));
    layer6_outputs(6390) <= layer5_outputs(4049);
    layer6_outputs(6391) <= not(layer5_outputs(2137));
    layer6_outputs(6392) <= not(layer5_outputs(1489));
    layer6_outputs(6393) <= layer5_outputs(412);
    layer6_outputs(6394) <= (layer5_outputs(6806)) and not (layer5_outputs(4281));
    layer6_outputs(6395) <= '0';
    layer6_outputs(6396) <= layer5_outputs(5792);
    layer6_outputs(6397) <= (layer5_outputs(2930)) and not (layer5_outputs(5114));
    layer6_outputs(6398) <= not((layer5_outputs(1472)) xor (layer5_outputs(6904)));
    layer6_outputs(6399) <= layer5_outputs(1686);
    layer6_outputs(6400) <= layer5_outputs(592);
    layer6_outputs(6401) <= (layer5_outputs(7496)) xor (layer5_outputs(1026));
    layer6_outputs(6402) <= layer5_outputs(5323);
    layer6_outputs(6403) <= layer5_outputs(6382);
    layer6_outputs(6404) <= not(layer5_outputs(5021));
    layer6_outputs(6405) <= layer5_outputs(3615);
    layer6_outputs(6406) <= (layer5_outputs(1266)) xor (layer5_outputs(3475));
    layer6_outputs(6407) <= not((layer5_outputs(209)) xor (layer5_outputs(320)));
    layer6_outputs(6408) <= not((layer5_outputs(4338)) xor (layer5_outputs(2824)));
    layer6_outputs(6409) <= not(layer5_outputs(4112));
    layer6_outputs(6410) <= not(layer5_outputs(778));
    layer6_outputs(6411) <= (layer5_outputs(7156)) xor (layer5_outputs(4631));
    layer6_outputs(6412) <= not(layer5_outputs(2482));
    layer6_outputs(6413) <= layer5_outputs(5816);
    layer6_outputs(6414) <= (layer5_outputs(4398)) and not (layer5_outputs(3098));
    layer6_outputs(6415) <= layer5_outputs(34);
    layer6_outputs(6416) <= not(layer5_outputs(3944));
    layer6_outputs(6417) <= not(layer5_outputs(3912));
    layer6_outputs(6418) <= '0';
    layer6_outputs(6419) <= not(layer5_outputs(58)) or (layer5_outputs(254));
    layer6_outputs(6420) <= not(layer5_outputs(4552));
    layer6_outputs(6421) <= not(layer5_outputs(7301));
    layer6_outputs(6422) <= (layer5_outputs(6679)) and not (layer5_outputs(4170));
    layer6_outputs(6423) <= not(layer5_outputs(6314));
    layer6_outputs(6424) <= not(layer5_outputs(6820));
    layer6_outputs(6425) <= not(layer5_outputs(6765));
    layer6_outputs(6426) <= not((layer5_outputs(5747)) xor (layer5_outputs(6230)));
    layer6_outputs(6427) <= not((layer5_outputs(6442)) or (layer5_outputs(6943)));
    layer6_outputs(6428) <= not((layer5_outputs(3858)) or (layer5_outputs(6171)));
    layer6_outputs(6429) <= not(layer5_outputs(5907)) or (layer5_outputs(1942));
    layer6_outputs(6430) <= not(layer5_outputs(4891));
    layer6_outputs(6431) <= not((layer5_outputs(2956)) and (layer5_outputs(7004)));
    layer6_outputs(6432) <= (layer5_outputs(4507)) xor (layer5_outputs(2907));
    layer6_outputs(6433) <= not(layer5_outputs(3805));
    layer6_outputs(6434) <= not((layer5_outputs(5289)) and (layer5_outputs(6060)));
    layer6_outputs(6435) <= not(layer5_outputs(5945));
    layer6_outputs(6436) <= not(layer5_outputs(3020));
    layer6_outputs(6437) <= not((layer5_outputs(4659)) xor (layer5_outputs(6013)));
    layer6_outputs(6438) <= not(layer5_outputs(1629));
    layer6_outputs(6439) <= not((layer5_outputs(403)) and (layer5_outputs(376)));
    layer6_outputs(6440) <= not(layer5_outputs(7641));
    layer6_outputs(6441) <= (layer5_outputs(4610)) or (layer5_outputs(4485));
    layer6_outputs(6442) <= layer5_outputs(6829);
    layer6_outputs(6443) <= not(layer5_outputs(382));
    layer6_outputs(6444) <= not(layer5_outputs(427));
    layer6_outputs(6445) <= not(layer5_outputs(7125));
    layer6_outputs(6446) <= layer5_outputs(7657);
    layer6_outputs(6447) <= not(layer5_outputs(3258)) or (layer5_outputs(5223));
    layer6_outputs(6448) <= layer5_outputs(4374);
    layer6_outputs(6449) <= not(layer5_outputs(1949));
    layer6_outputs(6450) <= layer5_outputs(5175);
    layer6_outputs(6451) <= (layer5_outputs(5144)) and not (layer5_outputs(815));
    layer6_outputs(6452) <= not((layer5_outputs(3367)) and (layer5_outputs(6648)));
    layer6_outputs(6453) <= layer5_outputs(3095);
    layer6_outputs(6454) <= not(layer5_outputs(595)) or (layer5_outputs(5331));
    layer6_outputs(6455) <= not(layer5_outputs(1436)) or (layer5_outputs(2513));
    layer6_outputs(6456) <= not(layer5_outputs(5512));
    layer6_outputs(6457) <= not(layer5_outputs(4476));
    layer6_outputs(6458) <= not((layer5_outputs(3392)) xor (layer5_outputs(5886)));
    layer6_outputs(6459) <= not(layer5_outputs(6242));
    layer6_outputs(6460) <= not(layer5_outputs(77));
    layer6_outputs(6461) <= (layer5_outputs(6091)) xor (layer5_outputs(379));
    layer6_outputs(6462) <= (layer5_outputs(2798)) xor (layer5_outputs(6240));
    layer6_outputs(6463) <= not((layer5_outputs(806)) or (layer5_outputs(254)));
    layer6_outputs(6464) <= layer5_outputs(2829);
    layer6_outputs(6465) <= not(layer5_outputs(1798));
    layer6_outputs(6466) <= (layer5_outputs(6110)) and not (layer5_outputs(6112));
    layer6_outputs(6467) <= '0';
    layer6_outputs(6468) <= layer5_outputs(1397);
    layer6_outputs(6469) <= (layer5_outputs(2912)) xor (layer5_outputs(1435));
    layer6_outputs(6470) <= (layer5_outputs(4413)) xor (layer5_outputs(2571));
    layer6_outputs(6471) <= not((layer5_outputs(4640)) xor (layer5_outputs(4212)));
    layer6_outputs(6472) <= layer5_outputs(5856);
    layer6_outputs(6473) <= (layer5_outputs(3337)) or (layer5_outputs(443));
    layer6_outputs(6474) <= (layer5_outputs(212)) or (layer5_outputs(860));
    layer6_outputs(6475) <= (layer5_outputs(841)) and not (layer5_outputs(7639));
    layer6_outputs(6476) <= layer5_outputs(4299);
    layer6_outputs(6477) <= not(layer5_outputs(3278)) or (layer5_outputs(5513));
    layer6_outputs(6478) <= (layer5_outputs(3035)) or (layer5_outputs(2174));
    layer6_outputs(6479) <= layer5_outputs(3784);
    layer6_outputs(6480) <= (layer5_outputs(7380)) and not (layer5_outputs(3166));
    layer6_outputs(6481) <= not((layer5_outputs(4184)) xor (layer5_outputs(4508)));
    layer6_outputs(6482) <= not(layer5_outputs(394));
    layer6_outputs(6483) <= not(layer5_outputs(2636)) or (layer5_outputs(3349));
    layer6_outputs(6484) <= not((layer5_outputs(4303)) xor (layer5_outputs(5464)));
    layer6_outputs(6485) <= not(layer5_outputs(5716));
    layer6_outputs(6486) <= layer5_outputs(642);
    layer6_outputs(6487) <= not(layer5_outputs(7362)) or (layer5_outputs(726));
    layer6_outputs(6488) <= (layer5_outputs(2273)) or (layer5_outputs(801));
    layer6_outputs(6489) <= layer5_outputs(357);
    layer6_outputs(6490) <= layer5_outputs(2838);
    layer6_outputs(6491) <= not(layer5_outputs(2819)) or (layer5_outputs(749));
    layer6_outputs(6492) <= not(layer5_outputs(5408));
    layer6_outputs(6493) <= not(layer5_outputs(3216));
    layer6_outputs(6494) <= layer5_outputs(2344);
    layer6_outputs(6495) <= (layer5_outputs(1654)) xor (layer5_outputs(4393));
    layer6_outputs(6496) <= not((layer5_outputs(1538)) and (layer5_outputs(7463)));
    layer6_outputs(6497) <= layer5_outputs(670);
    layer6_outputs(6498) <= not(layer5_outputs(7656));
    layer6_outputs(6499) <= not(layer5_outputs(4256)) or (layer5_outputs(7145));
    layer6_outputs(6500) <= not((layer5_outputs(3446)) or (layer5_outputs(844)));
    layer6_outputs(6501) <= not((layer5_outputs(237)) or (layer5_outputs(6660)));
    layer6_outputs(6502) <= layer5_outputs(3899);
    layer6_outputs(6503) <= layer5_outputs(5717);
    layer6_outputs(6504) <= not(layer5_outputs(1704));
    layer6_outputs(6505) <= (layer5_outputs(5572)) or (layer5_outputs(3412));
    layer6_outputs(6506) <= not(layer5_outputs(3593));
    layer6_outputs(6507) <= layer5_outputs(2608);
    layer6_outputs(6508) <= not(layer5_outputs(2031)) or (layer5_outputs(1117));
    layer6_outputs(6509) <= layer5_outputs(4524);
    layer6_outputs(6510) <= (layer5_outputs(7549)) and (layer5_outputs(6058));
    layer6_outputs(6511) <= (layer5_outputs(6380)) or (layer5_outputs(4125));
    layer6_outputs(6512) <= not(layer5_outputs(1510));
    layer6_outputs(6513) <= not((layer5_outputs(4569)) or (layer5_outputs(2270)));
    layer6_outputs(6514) <= not((layer5_outputs(6585)) and (layer5_outputs(6104)));
    layer6_outputs(6515) <= not(layer5_outputs(1351)) or (layer5_outputs(1268));
    layer6_outputs(6516) <= (layer5_outputs(1010)) and not (layer5_outputs(5035));
    layer6_outputs(6517) <= layer5_outputs(4252);
    layer6_outputs(6518) <= layer5_outputs(7084);
    layer6_outputs(6519) <= (layer5_outputs(1577)) and not (layer5_outputs(2401));
    layer6_outputs(6520) <= (layer5_outputs(4067)) xor (layer5_outputs(3876));
    layer6_outputs(6521) <= (layer5_outputs(3632)) xor (layer5_outputs(1374));
    layer6_outputs(6522) <= (layer5_outputs(5880)) and not (layer5_outputs(897));
    layer6_outputs(6523) <= layer5_outputs(4827);
    layer6_outputs(6524) <= layer5_outputs(1441);
    layer6_outputs(6525) <= not(layer5_outputs(5216));
    layer6_outputs(6526) <= not(layer5_outputs(3828));
    layer6_outputs(6527) <= (layer5_outputs(2593)) xor (layer5_outputs(6537));
    layer6_outputs(6528) <= (layer5_outputs(4875)) and not (layer5_outputs(2796));
    layer6_outputs(6529) <= not(layer5_outputs(1576)) or (layer5_outputs(4058));
    layer6_outputs(6530) <= (layer5_outputs(2864)) xor (layer5_outputs(1987));
    layer6_outputs(6531) <= (layer5_outputs(5202)) or (layer5_outputs(942));
    layer6_outputs(6532) <= not((layer5_outputs(1439)) or (layer5_outputs(6955)));
    layer6_outputs(6533) <= layer5_outputs(5347);
    layer6_outputs(6534) <= layer5_outputs(6219);
    layer6_outputs(6535) <= not((layer5_outputs(2057)) and (layer5_outputs(2715)));
    layer6_outputs(6536) <= not((layer5_outputs(672)) xor (layer5_outputs(500)));
    layer6_outputs(6537) <= (layer5_outputs(5065)) or (layer5_outputs(1760));
    layer6_outputs(6538) <= not((layer5_outputs(3518)) or (layer5_outputs(4438)));
    layer6_outputs(6539) <= not(layer5_outputs(5303));
    layer6_outputs(6540) <= not((layer5_outputs(6106)) or (layer5_outputs(4649)));
    layer6_outputs(6541) <= not((layer5_outputs(5003)) or (layer5_outputs(4121)));
    layer6_outputs(6542) <= layer5_outputs(7447);
    layer6_outputs(6543) <= layer5_outputs(4045);
    layer6_outputs(6544) <= not(layer5_outputs(5362));
    layer6_outputs(6545) <= not(layer5_outputs(7553));
    layer6_outputs(6546) <= (layer5_outputs(3850)) and not (layer5_outputs(2950));
    layer6_outputs(6547) <= not(layer5_outputs(2163));
    layer6_outputs(6548) <= layer5_outputs(7296);
    layer6_outputs(6549) <= layer5_outputs(5881);
    layer6_outputs(6550) <= (layer5_outputs(4646)) and not (layer5_outputs(3319));
    layer6_outputs(6551) <= layer5_outputs(4526);
    layer6_outputs(6552) <= layer5_outputs(5108);
    layer6_outputs(6553) <= not((layer5_outputs(6043)) or (layer5_outputs(4613)));
    layer6_outputs(6554) <= not(layer5_outputs(3524));
    layer6_outputs(6555) <= not(layer5_outputs(5080));
    layer6_outputs(6556) <= not(layer5_outputs(1086));
    layer6_outputs(6557) <= not(layer5_outputs(4221));
    layer6_outputs(6558) <= not(layer5_outputs(3551));
    layer6_outputs(6559) <= not(layer5_outputs(2192));
    layer6_outputs(6560) <= not(layer5_outputs(2749));
    layer6_outputs(6561) <= not((layer5_outputs(1922)) xor (layer5_outputs(2329)));
    layer6_outputs(6562) <= (layer5_outputs(5709)) xor (layer5_outputs(2574));
    layer6_outputs(6563) <= not(layer5_outputs(3285));
    layer6_outputs(6564) <= not(layer5_outputs(4174));
    layer6_outputs(6565) <= (layer5_outputs(745)) or (layer5_outputs(4340));
    layer6_outputs(6566) <= not(layer5_outputs(4890));
    layer6_outputs(6567) <= not((layer5_outputs(7262)) xor (layer5_outputs(561)));
    layer6_outputs(6568) <= not((layer5_outputs(1039)) xor (layer5_outputs(1941)));
    layer6_outputs(6569) <= not(layer5_outputs(6097));
    layer6_outputs(6570) <= (layer5_outputs(6041)) or (layer5_outputs(5448));
    layer6_outputs(6571) <= not(layer5_outputs(4881));
    layer6_outputs(6572) <= (layer5_outputs(7324)) and not (layer5_outputs(5766));
    layer6_outputs(6573) <= (layer5_outputs(2732)) xor (layer5_outputs(1926));
    layer6_outputs(6574) <= (layer5_outputs(6426)) xor (layer5_outputs(5305));
    layer6_outputs(6575) <= layer5_outputs(2524);
    layer6_outputs(6576) <= (layer5_outputs(5519)) and not (layer5_outputs(2141));
    layer6_outputs(6577) <= (layer5_outputs(5951)) or (layer5_outputs(6067));
    layer6_outputs(6578) <= (layer5_outputs(6699)) and not (layer5_outputs(1355));
    layer6_outputs(6579) <= (layer5_outputs(5771)) xor (layer5_outputs(4381));
    layer6_outputs(6580) <= not((layer5_outputs(968)) xor (layer5_outputs(1031)));
    layer6_outputs(6581) <= (layer5_outputs(5163)) or (layer5_outputs(805));
    layer6_outputs(6582) <= not(layer5_outputs(4721));
    layer6_outputs(6583) <= not(layer5_outputs(849)) or (layer5_outputs(960));
    layer6_outputs(6584) <= layer5_outputs(212);
    layer6_outputs(6585) <= not(layer5_outputs(4253));
    layer6_outputs(6586) <= not(layer5_outputs(7418));
    layer6_outputs(6587) <= (layer5_outputs(1953)) and (layer5_outputs(6329));
    layer6_outputs(6588) <= not((layer5_outputs(1167)) or (layer5_outputs(5571)));
    layer6_outputs(6589) <= layer5_outputs(5821);
    layer6_outputs(6590) <= not(layer5_outputs(6838));
    layer6_outputs(6591) <= not(layer5_outputs(260));
    layer6_outputs(6592) <= not((layer5_outputs(7467)) xor (layer5_outputs(7410)));
    layer6_outputs(6593) <= layer5_outputs(3380);
    layer6_outputs(6594) <= layer5_outputs(7311);
    layer6_outputs(6595) <= (layer5_outputs(807)) xor (layer5_outputs(5564));
    layer6_outputs(6596) <= not(layer5_outputs(367));
    layer6_outputs(6597) <= (layer5_outputs(538)) or (layer5_outputs(4338));
    layer6_outputs(6598) <= (layer5_outputs(3754)) and not (layer5_outputs(4572));
    layer6_outputs(6599) <= not(layer5_outputs(4586));
    layer6_outputs(6600) <= layer5_outputs(2124);
    layer6_outputs(6601) <= layer5_outputs(3183);
    layer6_outputs(6602) <= (layer5_outputs(6957)) or (layer5_outputs(1011));
    layer6_outputs(6603) <= not(layer5_outputs(4309));
    layer6_outputs(6604) <= not(layer5_outputs(936));
    layer6_outputs(6605) <= (layer5_outputs(145)) and not (layer5_outputs(5268));
    layer6_outputs(6606) <= (layer5_outputs(4828)) xor (layer5_outputs(3906));
    layer6_outputs(6607) <= layer5_outputs(1409);
    layer6_outputs(6608) <= layer5_outputs(5902);
    layer6_outputs(6609) <= (layer5_outputs(6803)) xor (layer5_outputs(1905));
    layer6_outputs(6610) <= not((layer5_outputs(837)) xor (layer5_outputs(5937)));
    layer6_outputs(6611) <= not(layer5_outputs(4674));
    layer6_outputs(6612) <= layer5_outputs(2195);
    layer6_outputs(6613) <= (layer5_outputs(1694)) and not (layer5_outputs(2709));
    layer6_outputs(6614) <= layer5_outputs(6661);
    layer6_outputs(6615) <= layer5_outputs(6916);
    layer6_outputs(6616) <= (layer5_outputs(2404)) xor (layer5_outputs(7023));
    layer6_outputs(6617) <= not(layer5_outputs(263));
    layer6_outputs(6618) <= not((layer5_outputs(4931)) xor (layer5_outputs(5832)));
    layer6_outputs(6619) <= layer5_outputs(6220);
    layer6_outputs(6620) <= (layer5_outputs(392)) and not (layer5_outputs(4573));
    layer6_outputs(6621) <= not((layer5_outputs(2190)) or (layer5_outputs(2089)));
    layer6_outputs(6622) <= not(layer5_outputs(4261));
    layer6_outputs(6623) <= not((layer5_outputs(356)) or (layer5_outputs(7359)));
    layer6_outputs(6624) <= layer5_outputs(2338);
    layer6_outputs(6625) <= layer5_outputs(2472);
    layer6_outputs(6626) <= layer5_outputs(5486);
    layer6_outputs(6627) <= not(layer5_outputs(3255)) or (layer5_outputs(7044));
    layer6_outputs(6628) <= (layer5_outputs(5506)) or (layer5_outputs(5194));
    layer6_outputs(6629) <= (layer5_outputs(6532)) and not (layer5_outputs(6272));
    layer6_outputs(6630) <= not(layer5_outputs(1903));
    layer6_outputs(6631) <= layer5_outputs(3170);
    layer6_outputs(6632) <= not((layer5_outputs(3716)) xor (layer5_outputs(1193)));
    layer6_outputs(6633) <= not(layer5_outputs(5227)) or (layer5_outputs(5156));
    layer6_outputs(6634) <= not(layer5_outputs(957));
    layer6_outputs(6635) <= not(layer5_outputs(1107));
    layer6_outputs(6636) <= not(layer5_outputs(64));
    layer6_outputs(6637) <= not(layer5_outputs(5055));
    layer6_outputs(6638) <= (layer5_outputs(6291)) and not (layer5_outputs(4401));
    layer6_outputs(6639) <= (layer5_outputs(5703)) and (layer5_outputs(130));
    layer6_outputs(6640) <= not(layer5_outputs(1531));
    layer6_outputs(6641) <= not(layer5_outputs(2248));
    layer6_outputs(6642) <= not(layer5_outputs(6578)) or (layer5_outputs(3440));
    layer6_outputs(6643) <= layer5_outputs(7557);
    layer6_outputs(6644) <= not(layer5_outputs(6826)) or (layer5_outputs(5246));
    layer6_outputs(6645) <= layer5_outputs(4284);
    layer6_outputs(6646) <= layer5_outputs(5275);
    layer6_outputs(6647) <= not(layer5_outputs(2208));
    layer6_outputs(6648) <= (layer5_outputs(7389)) xor (layer5_outputs(1198));
    layer6_outputs(6649) <= layer5_outputs(941);
    layer6_outputs(6650) <= not(layer5_outputs(4205));
    layer6_outputs(6651) <= '1';
    layer6_outputs(6652) <= not(layer5_outputs(956));
    layer6_outputs(6653) <= '1';
    layer6_outputs(6654) <= layer5_outputs(354);
    layer6_outputs(6655) <= not((layer5_outputs(1305)) xor (layer5_outputs(4667)));
    layer6_outputs(6656) <= not(layer5_outputs(1362));
    layer6_outputs(6657) <= (layer5_outputs(222)) xor (layer5_outputs(1796));
    layer6_outputs(6658) <= not(layer5_outputs(4525));
    layer6_outputs(6659) <= layer5_outputs(6329);
    layer6_outputs(6660) <= layer5_outputs(441);
    layer6_outputs(6661) <= (layer5_outputs(4793)) or (layer5_outputs(2937));
    layer6_outputs(6662) <= (layer5_outputs(5262)) xor (layer5_outputs(394));
    layer6_outputs(6663) <= (layer5_outputs(5039)) xor (layer5_outputs(4494));
    layer6_outputs(6664) <= not((layer5_outputs(337)) xor (layer5_outputs(5619)));
    layer6_outputs(6665) <= layer5_outputs(7591);
    layer6_outputs(6666) <= layer5_outputs(1975);
    layer6_outputs(6667) <= layer5_outputs(4221);
    layer6_outputs(6668) <= (layer5_outputs(5895)) and not (layer5_outputs(111));
    layer6_outputs(6669) <= (layer5_outputs(3888)) and not (layer5_outputs(5584));
    layer6_outputs(6670) <= not(layer5_outputs(981));
    layer6_outputs(6671) <= (layer5_outputs(6376)) or (layer5_outputs(759));
    layer6_outputs(6672) <= not(layer5_outputs(797));
    layer6_outputs(6673) <= layer5_outputs(4941);
    layer6_outputs(6674) <= not((layer5_outputs(343)) or (layer5_outputs(1982)));
    layer6_outputs(6675) <= not(layer5_outputs(7287));
    layer6_outputs(6676) <= layer5_outputs(625);
    layer6_outputs(6677) <= layer5_outputs(3619);
    layer6_outputs(6678) <= layer5_outputs(7461);
    layer6_outputs(6679) <= not(layer5_outputs(1633));
    layer6_outputs(6680) <= layer5_outputs(1122);
    layer6_outputs(6681) <= not(layer5_outputs(4806));
    layer6_outputs(6682) <= (layer5_outputs(1986)) or (layer5_outputs(1888));
    layer6_outputs(6683) <= layer5_outputs(3566);
    layer6_outputs(6684) <= not(layer5_outputs(6328));
    layer6_outputs(6685) <= layer5_outputs(629);
    layer6_outputs(6686) <= not(layer5_outputs(7451)) or (layer5_outputs(4918));
    layer6_outputs(6687) <= layer5_outputs(1562);
    layer6_outputs(6688) <= not(layer5_outputs(7246));
    layer6_outputs(6689) <= not((layer5_outputs(2396)) and (layer5_outputs(2249)));
    layer6_outputs(6690) <= layer5_outputs(6591);
    layer6_outputs(6691) <= not(layer5_outputs(5140));
    layer6_outputs(6692) <= layer5_outputs(5811);
    layer6_outputs(6693) <= '0';
    layer6_outputs(6694) <= layer5_outputs(5129);
    layer6_outputs(6695) <= not((layer5_outputs(2207)) xor (layer5_outputs(1197)));
    layer6_outputs(6696) <= not(layer5_outputs(2771));
    layer6_outputs(6697) <= (layer5_outputs(1745)) or (layer5_outputs(4714));
    layer6_outputs(6698) <= not(layer5_outputs(1613));
    layer6_outputs(6699) <= layer5_outputs(3300);
    layer6_outputs(6700) <= layer5_outputs(4773);
    layer6_outputs(6701) <= layer5_outputs(5456);
    layer6_outputs(6702) <= not((layer5_outputs(3870)) xor (layer5_outputs(794)));
    layer6_outputs(6703) <= layer5_outputs(2500);
    layer6_outputs(6704) <= not((layer5_outputs(5516)) xor (layer5_outputs(4705)));
    layer6_outputs(6705) <= not((layer5_outputs(7164)) xor (layer5_outputs(2952)));
    layer6_outputs(6706) <= not((layer5_outputs(4744)) xor (layer5_outputs(6510)));
    layer6_outputs(6707) <= layer5_outputs(6605);
    layer6_outputs(6708) <= not(layer5_outputs(1225));
    layer6_outputs(6709) <= (layer5_outputs(6751)) and (layer5_outputs(2047));
    layer6_outputs(6710) <= (layer5_outputs(3870)) xor (layer5_outputs(826));
    layer6_outputs(6711) <= not(layer5_outputs(3640)) or (layer5_outputs(5525));
    layer6_outputs(6712) <= (layer5_outputs(1555)) xor (layer5_outputs(7306));
    layer6_outputs(6713) <= not(layer5_outputs(7516)) or (layer5_outputs(2546));
    layer6_outputs(6714) <= not((layer5_outputs(5112)) and (layer5_outputs(7096)));
    layer6_outputs(6715) <= layer5_outputs(156);
    layer6_outputs(6716) <= not(layer5_outputs(7383));
    layer6_outputs(6717) <= not((layer5_outputs(5000)) xor (layer5_outputs(5423)));
    layer6_outputs(6718) <= (layer5_outputs(1311)) and not (layer5_outputs(6016));
    layer6_outputs(6719) <= not(layer5_outputs(5001));
    layer6_outputs(6720) <= (layer5_outputs(667)) xor (layer5_outputs(1655));
    layer6_outputs(6721) <= (layer5_outputs(3053)) and (layer5_outputs(3180));
    layer6_outputs(6722) <= not((layer5_outputs(2256)) and (layer5_outputs(4782)));
    layer6_outputs(6723) <= layer5_outputs(2810);
    layer6_outputs(6724) <= not(layer5_outputs(4531));
    layer6_outputs(6725) <= layer5_outputs(4495);
    layer6_outputs(6726) <= not(layer5_outputs(2578));
    layer6_outputs(6727) <= layer5_outputs(760);
    layer6_outputs(6728) <= (layer5_outputs(7560)) and not (layer5_outputs(383));
    layer6_outputs(6729) <= not(layer5_outputs(2259));
    layer6_outputs(6730) <= not(layer5_outputs(5651));
    layer6_outputs(6731) <= layer5_outputs(3159);
    layer6_outputs(6732) <= not(layer5_outputs(1260));
    layer6_outputs(6733) <= layer5_outputs(5703);
    layer6_outputs(6734) <= not((layer5_outputs(1396)) or (layer5_outputs(3695)));
    layer6_outputs(6735) <= not(layer5_outputs(5461));
    layer6_outputs(6736) <= '1';
    layer6_outputs(6737) <= not(layer5_outputs(6562)) or (layer5_outputs(4437));
    layer6_outputs(6738) <= (layer5_outputs(1315)) and not (layer5_outputs(5597));
    layer6_outputs(6739) <= (layer5_outputs(6128)) and not (layer5_outputs(5092));
    layer6_outputs(6740) <= not(layer5_outputs(7011));
    layer6_outputs(6741) <= not(layer5_outputs(7213));
    layer6_outputs(6742) <= layer5_outputs(6086);
    layer6_outputs(6743) <= layer5_outputs(472);
    layer6_outputs(6744) <= (layer5_outputs(7228)) xor (layer5_outputs(4858));
    layer6_outputs(6745) <= (layer5_outputs(4123)) or (layer5_outputs(3744));
    layer6_outputs(6746) <= not(layer5_outputs(5550));
    layer6_outputs(6747) <= not(layer5_outputs(3291));
    layer6_outputs(6748) <= (layer5_outputs(2574)) and (layer5_outputs(6265));
    layer6_outputs(6749) <= not(layer5_outputs(3575));
    layer6_outputs(6750) <= not((layer5_outputs(5823)) xor (layer5_outputs(5836)));
    layer6_outputs(6751) <= (layer5_outputs(1663)) and not (layer5_outputs(6740));
    layer6_outputs(6752) <= not((layer5_outputs(719)) or (layer5_outputs(5588)));
    layer6_outputs(6753) <= not(layer5_outputs(2826));
    layer6_outputs(6754) <= not(layer5_outputs(5746));
    layer6_outputs(6755) <= not(layer5_outputs(6392)) or (layer5_outputs(7049));
    layer6_outputs(6756) <= layer5_outputs(31);
    layer6_outputs(6757) <= not((layer5_outputs(5099)) xor (layer5_outputs(1410)));
    layer6_outputs(6758) <= layer5_outputs(7079);
    layer6_outputs(6759) <= not((layer5_outputs(3983)) xor (layer5_outputs(5829)));
    layer6_outputs(6760) <= not(layer5_outputs(1688)) or (layer5_outputs(1816));
    layer6_outputs(6761) <= not((layer5_outputs(5020)) xor (layer5_outputs(4500)));
    layer6_outputs(6762) <= (layer5_outputs(3690)) and not (layer5_outputs(6515));
    layer6_outputs(6763) <= not(layer5_outputs(2670));
    layer6_outputs(6764) <= not(layer5_outputs(6287));
    layer6_outputs(6765) <= not(layer5_outputs(7107));
    layer6_outputs(6766) <= layer5_outputs(4918);
    layer6_outputs(6767) <= (layer5_outputs(6601)) and not (layer5_outputs(4688));
    layer6_outputs(6768) <= layer5_outputs(3032);
    layer6_outputs(6769) <= not(layer5_outputs(5478));
    layer6_outputs(6770) <= not(layer5_outputs(6780));
    layer6_outputs(6771) <= not(layer5_outputs(7440)) or (layer5_outputs(2140));
    layer6_outputs(6772) <= layer5_outputs(4057);
    layer6_outputs(6773) <= layer5_outputs(2676);
    layer6_outputs(6774) <= (layer5_outputs(3200)) xor (layer5_outputs(3604));
    layer6_outputs(6775) <= layer5_outputs(1979);
    layer6_outputs(6776) <= not(layer5_outputs(5473)) or (layer5_outputs(4870));
    layer6_outputs(6777) <= (layer5_outputs(850)) xor (layer5_outputs(1549));
    layer6_outputs(6778) <= (layer5_outputs(1626)) or (layer5_outputs(902));
    layer6_outputs(6779) <= (layer5_outputs(5628)) and not (layer5_outputs(236));
    layer6_outputs(6780) <= (layer5_outputs(24)) and (layer5_outputs(2169));
    layer6_outputs(6781) <= (layer5_outputs(6406)) and (layer5_outputs(2806));
    layer6_outputs(6782) <= not((layer5_outputs(2781)) xor (layer5_outputs(983)));
    layer6_outputs(6783) <= not(layer5_outputs(3795));
    layer6_outputs(6784) <= not((layer5_outputs(6980)) and (layer5_outputs(7431)));
    layer6_outputs(6785) <= not(layer5_outputs(3246));
    layer6_outputs(6786) <= not((layer5_outputs(7038)) xor (layer5_outputs(6806)));
    layer6_outputs(6787) <= layer5_outputs(65);
    layer6_outputs(6788) <= (layer5_outputs(5892)) and not (layer5_outputs(2544));
    layer6_outputs(6789) <= layer5_outputs(6830);
    layer6_outputs(6790) <= layer5_outputs(1971);
    layer6_outputs(6791) <= not((layer5_outputs(1414)) and (layer5_outputs(3602)));
    layer6_outputs(6792) <= not((layer5_outputs(6487)) or (layer5_outputs(4050)));
    layer6_outputs(6793) <= not(layer5_outputs(6644));
    layer6_outputs(6794) <= not(layer5_outputs(5250));
    layer6_outputs(6795) <= (layer5_outputs(4753)) and not (layer5_outputs(4468));
    layer6_outputs(6796) <= layer5_outputs(5495);
    layer6_outputs(6797) <= not(layer5_outputs(5873)) or (layer5_outputs(1400));
    layer6_outputs(6798) <= not(layer5_outputs(5632));
    layer6_outputs(6799) <= not(layer5_outputs(3778));
    layer6_outputs(6800) <= layer5_outputs(5625);
    layer6_outputs(6801) <= not((layer5_outputs(409)) xor (layer5_outputs(1152)));
    layer6_outputs(6802) <= (layer5_outputs(2647)) and (layer5_outputs(1795));
    layer6_outputs(6803) <= not(layer5_outputs(7550));
    layer6_outputs(6804) <= (layer5_outputs(7537)) xor (layer5_outputs(6682));
    layer6_outputs(6805) <= not((layer5_outputs(3854)) or (layer5_outputs(135)));
    layer6_outputs(6806) <= (layer5_outputs(1908)) xor (layer5_outputs(4227));
    layer6_outputs(6807) <= layer5_outputs(5283);
    layer6_outputs(6808) <= (layer5_outputs(751)) and (layer5_outputs(7230));
    layer6_outputs(6809) <= layer5_outputs(2327);
    layer6_outputs(6810) <= layer5_outputs(7397);
    layer6_outputs(6811) <= layer5_outputs(1708);
    layer6_outputs(6812) <= layer5_outputs(2345);
    layer6_outputs(6813) <= not(layer5_outputs(4695));
    layer6_outputs(6814) <= (layer5_outputs(2567)) and not (layer5_outputs(6099));
    layer6_outputs(6815) <= (layer5_outputs(2859)) xor (layer5_outputs(2514));
    layer6_outputs(6816) <= layer5_outputs(5474);
    layer6_outputs(6817) <= not((layer5_outputs(1056)) or (layer5_outputs(642)));
    layer6_outputs(6818) <= not(layer5_outputs(753)) or (layer5_outputs(6261));
    layer6_outputs(6819) <= layer5_outputs(1021);
    layer6_outputs(6820) <= not(layer5_outputs(4761));
    layer6_outputs(6821) <= not(layer5_outputs(918));
    layer6_outputs(6822) <= not(layer5_outputs(5440)) or (layer5_outputs(654));
    layer6_outputs(6823) <= layer5_outputs(3631);
    layer6_outputs(6824) <= layer5_outputs(2278);
    layer6_outputs(6825) <= layer5_outputs(6134);
    layer6_outputs(6826) <= not(layer5_outputs(5184));
    layer6_outputs(6827) <= (layer5_outputs(4574)) and not (layer5_outputs(22));
    layer6_outputs(6828) <= not(layer5_outputs(3746));
    layer6_outputs(6829) <= layer5_outputs(3996);
    layer6_outputs(6830) <= (layer5_outputs(1820)) and not (layer5_outputs(442));
    layer6_outputs(6831) <= (layer5_outputs(1680)) and not (layer5_outputs(3125));
    layer6_outputs(6832) <= (layer5_outputs(6049)) xor (layer5_outputs(1176));
    layer6_outputs(6833) <= not(layer5_outputs(3116));
    layer6_outputs(6834) <= not((layer5_outputs(4295)) or (layer5_outputs(6199)));
    layer6_outputs(6835) <= not(layer5_outputs(2566));
    layer6_outputs(6836) <= (layer5_outputs(7128)) and not (layer5_outputs(5488));
    layer6_outputs(6837) <= not((layer5_outputs(2067)) xor (layer5_outputs(4399)));
    layer6_outputs(6838) <= not(layer5_outputs(420));
    layer6_outputs(6839) <= not(layer5_outputs(763));
    layer6_outputs(6840) <= not(layer5_outputs(2579));
    layer6_outputs(6841) <= layer5_outputs(7609);
    layer6_outputs(6842) <= not((layer5_outputs(386)) xor (layer5_outputs(5927)));
    layer6_outputs(6843) <= not(layer5_outputs(6950));
    layer6_outputs(6844) <= (layer5_outputs(2420)) or (layer5_outputs(6247));
    layer6_outputs(6845) <= not(layer5_outputs(880));
    layer6_outputs(6846) <= not(layer5_outputs(4456));
    layer6_outputs(6847) <= not(layer5_outputs(6977));
    layer6_outputs(6848) <= layer5_outputs(2233);
    layer6_outputs(6849) <= not((layer5_outputs(7319)) and (layer5_outputs(5581)));
    layer6_outputs(6850) <= layer5_outputs(7081);
    layer6_outputs(6851) <= (layer5_outputs(6705)) or (layer5_outputs(6449));
    layer6_outputs(6852) <= not(layer5_outputs(617));
    layer6_outputs(6853) <= layer5_outputs(3406);
    layer6_outputs(6854) <= not(layer5_outputs(6275));
    layer6_outputs(6855) <= layer5_outputs(1742);
    layer6_outputs(6856) <= not(layer5_outputs(6213));
    layer6_outputs(6857) <= layer5_outputs(5561);
    layer6_outputs(6858) <= layer5_outputs(3760);
    layer6_outputs(6859) <= not(layer5_outputs(2401));
    layer6_outputs(6860) <= (layer5_outputs(3740)) xor (layer5_outputs(1403));
    layer6_outputs(6861) <= not(layer5_outputs(7116)) or (layer5_outputs(5849));
    layer6_outputs(6862) <= layer5_outputs(166);
    layer6_outputs(6863) <= not(layer5_outputs(2753));
    layer6_outputs(6864) <= (layer5_outputs(489)) xor (layer5_outputs(2230));
    layer6_outputs(6865) <= (layer5_outputs(4291)) and (layer5_outputs(828));
    layer6_outputs(6866) <= (layer5_outputs(4006)) and (layer5_outputs(6775));
    layer6_outputs(6867) <= not(layer5_outputs(2588));
    layer6_outputs(6868) <= layer5_outputs(564);
    layer6_outputs(6869) <= not(layer5_outputs(7285));
    layer6_outputs(6870) <= not(layer5_outputs(1263));
    layer6_outputs(6871) <= layer5_outputs(423);
    layer6_outputs(6872) <= layer5_outputs(1079);
    layer6_outputs(6873) <= not(layer5_outputs(2880));
    layer6_outputs(6874) <= not(layer5_outputs(5971)) or (layer5_outputs(4885));
    layer6_outputs(6875) <= not((layer5_outputs(1659)) xor (layer5_outputs(4436)));
    layer6_outputs(6876) <= not(layer5_outputs(6583));
    layer6_outputs(6877) <= layer5_outputs(6416);
    layer6_outputs(6878) <= not((layer5_outputs(4601)) and (layer5_outputs(1161)));
    layer6_outputs(6879) <= layer5_outputs(2524);
    layer6_outputs(6880) <= layer5_outputs(3141);
    layer6_outputs(6881) <= (layer5_outputs(2180)) xor (layer5_outputs(3205));
    layer6_outputs(6882) <= (layer5_outputs(6415)) and not (layer5_outputs(6879));
    layer6_outputs(6883) <= not((layer5_outputs(7663)) xor (layer5_outputs(4999)));
    layer6_outputs(6884) <= layer5_outputs(2739);
    layer6_outputs(6885) <= not(layer5_outputs(3002));
    layer6_outputs(6886) <= layer5_outputs(952);
    layer6_outputs(6887) <= not(layer5_outputs(3314));
    layer6_outputs(6888) <= not(layer5_outputs(654));
    layer6_outputs(6889) <= (layer5_outputs(723)) and (layer5_outputs(4183));
    layer6_outputs(6890) <= not(layer5_outputs(7295));
    layer6_outputs(6891) <= layer5_outputs(3123);
    layer6_outputs(6892) <= not((layer5_outputs(5173)) or (layer5_outputs(2924)));
    layer6_outputs(6893) <= (layer5_outputs(2236)) and not (layer5_outputs(4045));
    layer6_outputs(6894) <= not((layer5_outputs(1652)) xor (layer5_outputs(5499)));
    layer6_outputs(6895) <= (layer5_outputs(3691)) xor (layer5_outputs(2261));
    layer6_outputs(6896) <= layer5_outputs(7084);
    layer6_outputs(6897) <= not(layer5_outputs(7395)) or (layer5_outputs(1476));
    layer6_outputs(6898) <= (layer5_outputs(4134)) xor (layer5_outputs(1705));
    layer6_outputs(6899) <= not(layer5_outputs(5898));
    layer6_outputs(6900) <= (layer5_outputs(5516)) xor (layer5_outputs(5684));
    layer6_outputs(6901) <= not(layer5_outputs(6518));
    layer6_outputs(6902) <= (layer5_outputs(7268)) and not (layer5_outputs(7637));
    layer6_outputs(6903) <= not(layer5_outputs(3796));
    layer6_outputs(6904) <= not(layer5_outputs(3174));
    layer6_outputs(6905) <= layer5_outputs(6193);
    layer6_outputs(6906) <= not(layer5_outputs(4214));
    layer6_outputs(6907) <= not(layer5_outputs(2670)) or (layer5_outputs(5292));
    layer6_outputs(6908) <= not(layer5_outputs(1146)) or (layer5_outputs(780));
    layer6_outputs(6909) <= not(layer5_outputs(191));
    layer6_outputs(6910) <= not(layer5_outputs(1363)) or (layer5_outputs(4475));
    layer6_outputs(6911) <= not(layer5_outputs(5306));
    layer6_outputs(6912) <= (layer5_outputs(359)) and not (layer5_outputs(3177));
    layer6_outputs(6913) <= not((layer5_outputs(4010)) or (layer5_outputs(1040)));
    layer6_outputs(6914) <= not(layer5_outputs(5010));
    layer6_outputs(6915) <= not((layer5_outputs(701)) and (layer5_outputs(5129)));
    layer6_outputs(6916) <= not(layer5_outputs(6045));
    layer6_outputs(6917) <= (layer5_outputs(6809)) and not (layer5_outputs(720));
    layer6_outputs(6918) <= not(layer5_outputs(4771));
    layer6_outputs(6919) <= not((layer5_outputs(6139)) xor (layer5_outputs(7267)));
    layer6_outputs(6920) <= layer5_outputs(2733);
    layer6_outputs(6921) <= not((layer5_outputs(3426)) xor (layer5_outputs(6214)));
    layer6_outputs(6922) <= not(layer5_outputs(6767));
    layer6_outputs(6923) <= layer5_outputs(2957);
    layer6_outputs(6924) <= not(layer5_outputs(738));
    layer6_outputs(6925) <= not((layer5_outputs(7454)) xor (layer5_outputs(7642)));
    layer6_outputs(6926) <= layer5_outputs(220);
    layer6_outputs(6927) <= layer5_outputs(2288);
    layer6_outputs(6928) <= not(layer5_outputs(7429));
    layer6_outputs(6929) <= not(layer5_outputs(2490));
    layer6_outputs(6930) <= not(layer5_outputs(6990));
    layer6_outputs(6931) <= layer5_outputs(5447);
    layer6_outputs(6932) <= not(layer5_outputs(2167));
    layer6_outputs(6933) <= not(layer5_outputs(2861));
    layer6_outputs(6934) <= not((layer5_outputs(246)) or (layer5_outputs(7505)));
    layer6_outputs(6935) <= not(layer5_outputs(5925));
    layer6_outputs(6936) <= layer5_outputs(6283);
    layer6_outputs(6937) <= layer5_outputs(6693);
    layer6_outputs(6938) <= not(layer5_outputs(6137));
    layer6_outputs(6939) <= layer5_outputs(4652);
    layer6_outputs(6940) <= not((layer5_outputs(5427)) or (layer5_outputs(5120)));
    layer6_outputs(6941) <= layer5_outputs(6479);
    layer6_outputs(6942) <= not((layer5_outputs(4937)) and (layer5_outputs(79)));
    layer6_outputs(6943) <= layer5_outputs(7400);
    layer6_outputs(6944) <= not(layer5_outputs(2878));
    layer6_outputs(6945) <= (layer5_outputs(3063)) xor (layer5_outputs(2726));
    layer6_outputs(6946) <= layer5_outputs(4984);
    layer6_outputs(6947) <= not(layer5_outputs(5682));
    layer6_outputs(6948) <= (layer5_outputs(4022)) and not (layer5_outputs(4292));
    layer6_outputs(6949) <= not((layer5_outputs(3980)) xor (layer5_outputs(6895)));
    layer6_outputs(6950) <= not((layer5_outputs(4363)) or (layer5_outputs(2664)));
    layer6_outputs(6951) <= layer5_outputs(5481);
    layer6_outputs(6952) <= not(layer5_outputs(468));
    layer6_outputs(6953) <= (layer5_outputs(6975)) and (layer5_outputs(786));
    layer6_outputs(6954) <= layer5_outputs(3244);
    layer6_outputs(6955) <= layer5_outputs(4373);
    layer6_outputs(6956) <= not((layer5_outputs(7471)) and (layer5_outputs(4098)));
    layer6_outputs(6957) <= layer5_outputs(7458);
    layer6_outputs(6958) <= not(layer5_outputs(5199));
    layer6_outputs(6959) <= (layer5_outputs(3346)) and not (layer5_outputs(4806));
    layer6_outputs(6960) <= not(layer5_outputs(4591));
    layer6_outputs(6961) <= not(layer5_outputs(6222));
    layer6_outputs(6962) <= layer5_outputs(6296);
    layer6_outputs(6963) <= layer5_outputs(1160);
    layer6_outputs(6964) <= not(layer5_outputs(7431));
    layer6_outputs(6965) <= layer5_outputs(6104);
    layer6_outputs(6966) <= layer5_outputs(1223);
    layer6_outputs(6967) <= layer5_outputs(161);
    layer6_outputs(6968) <= (layer5_outputs(6425)) and (layer5_outputs(4965));
    layer6_outputs(6969) <= layer5_outputs(6854);
    layer6_outputs(6970) <= layer5_outputs(2163);
    layer6_outputs(6971) <= not(layer5_outputs(7569)) or (layer5_outputs(4865));
    layer6_outputs(6972) <= layer5_outputs(3649);
    layer6_outputs(6973) <= not(layer5_outputs(4019)) or (layer5_outputs(2076));
    layer6_outputs(6974) <= not(layer5_outputs(1276));
    layer6_outputs(6975) <= not((layer5_outputs(5399)) xor (layer5_outputs(6214)));
    layer6_outputs(6976) <= layer5_outputs(7026);
    layer6_outputs(6977) <= not(layer5_outputs(1295));
    layer6_outputs(6978) <= not(layer5_outputs(1221));
    layer6_outputs(6979) <= not((layer5_outputs(6095)) xor (layer5_outputs(2622)));
    layer6_outputs(6980) <= (layer5_outputs(1009)) and not (layer5_outputs(4372));
    layer6_outputs(6981) <= not(layer5_outputs(6182));
    layer6_outputs(6982) <= (layer5_outputs(84)) and (layer5_outputs(6548));
    layer6_outputs(6983) <= not(layer5_outputs(4187));
    layer6_outputs(6984) <= not(layer5_outputs(6835));
    layer6_outputs(6985) <= layer5_outputs(5824);
    layer6_outputs(6986) <= not((layer5_outputs(2232)) xor (layer5_outputs(4416)));
    layer6_outputs(6987) <= not(layer5_outputs(2322));
    layer6_outputs(6988) <= (layer5_outputs(1819)) or (layer5_outputs(3620));
    layer6_outputs(6989) <= not(layer5_outputs(6975));
    layer6_outputs(6990) <= (layer5_outputs(3907)) and (layer5_outputs(6884));
    layer6_outputs(6991) <= layer5_outputs(3476);
    layer6_outputs(6992) <= layer5_outputs(2690);
    layer6_outputs(6993) <= not(layer5_outputs(5696));
    layer6_outputs(6994) <= layer5_outputs(2699);
    layer6_outputs(6995) <= not(layer5_outputs(192));
    layer6_outputs(6996) <= not((layer5_outputs(7165)) xor (layer5_outputs(2036)));
    layer6_outputs(6997) <= (layer5_outputs(7199)) or (layer5_outputs(5670));
    layer6_outputs(6998) <= layer5_outputs(1997);
    layer6_outputs(6999) <= not((layer5_outputs(5539)) xor (layer5_outputs(5545)));
    layer6_outputs(7000) <= not(layer5_outputs(166)) or (layer5_outputs(3905));
    layer6_outputs(7001) <= not(layer5_outputs(6935));
    layer6_outputs(7002) <= (layer5_outputs(3846)) and not (layer5_outputs(3580));
    layer6_outputs(7003) <= layer5_outputs(1377);
    layer6_outputs(7004) <= '0';
    layer6_outputs(7005) <= layer5_outputs(7054);
    layer6_outputs(7006) <= not(layer5_outputs(6258));
    layer6_outputs(7007) <= (layer5_outputs(5990)) and (layer5_outputs(6133));
    layer6_outputs(7008) <= layer5_outputs(3501);
    layer6_outputs(7009) <= layer5_outputs(904);
    layer6_outputs(7010) <= (layer5_outputs(593)) and (layer5_outputs(5190));
    layer6_outputs(7011) <= not(layer5_outputs(47)) or (layer5_outputs(6456));
    layer6_outputs(7012) <= not(layer5_outputs(5877));
    layer6_outputs(7013) <= not((layer5_outputs(4773)) xor (layer5_outputs(458)));
    layer6_outputs(7014) <= layer5_outputs(4068);
    layer6_outputs(7015) <= layer5_outputs(6298);
    layer6_outputs(7016) <= layer5_outputs(1440);
    layer6_outputs(7017) <= not(layer5_outputs(4441));
    layer6_outputs(7018) <= not(layer5_outputs(2935));
    layer6_outputs(7019) <= not(layer5_outputs(1785));
    layer6_outputs(7020) <= layer5_outputs(5064);
    layer6_outputs(7021) <= layer5_outputs(1178);
    layer6_outputs(7022) <= (layer5_outputs(3807)) and (layer5_outputs(5724));
    layer6_outputs(7023) <= layer5_outputs(1808);
    layer6_outputs(7024) <= not(layer5_outputs(7201));
    layer6_outputs(7025) <= not((layer5_outputs(376)) xor (layer5_outputs(4919)));
    layer6_outputs(7026) <= not(layer5_outputs(6358));
    layer6_outputs(7027) <= not((layer5_outputs(1624)) xor (layer5_outputs(5725)));
    layer6_outputs(7028) <= (layer5_outputs(4401)) or (layer5_outputs(6467));
    layer6_outputs(7029) <= layer5_outputs(803);
    layer6_outputs(7030) <= (layer5_outputs(5050)) xor (layer5_outputs(7412));
    layer6_outputs(7031) <= (layer5_outputs(2980)) xor (layer5_outputs(6010));
    layer6_outputs(7032) <= not((layer5_outputs(297)) and (layer5_outputs(945)));
    layer6_outputs(7033) <= not(layer5_outputs(3355));
    layer6_outputs(7034) <= not((layer5_outputs(3730)) xor (layer5_outputs(7518)));
    layer6_outputs(7035) <= not(layer5_outputs(7450));
    layer6_outputs(7036) <= layer5_outputs(7131);
    layer6_outputs(7037) <= layer5_outputs(3711);
    layer6_outputs(7038) <= not((layer5_outputs(5232)) and (layer5_outputs(1892)));
    layer6_outputs(7039) <= not((layer5_outputs(4997)) xor (layer5_outputs(984)));
    layer6_outputs(7040) <= not(layer5_outputs(3377));
    layer6_outputs(7041) <= not((layer5_outputs(1024)) xor (layer5_outputs(5212)));
    layer6_outputs(7042) <= not((layer5_outputs(3503)) or (layer5_outputs(5863)));
    layer6_outputs(7043) <= (layer5_outputs(6454)) and (layer5_outputs(1462));
    layer6_outputs(7044) <= not(layer5_outputs(1047));
    layer6_outputs(7045) <= not(layer5_outputs(6800)) or (layer5_outputs(2872));
    layer6_outputs(7046) <= not(layer5_outputs(1712));
    layer6_outputs(7047) <= not((layer5_outputs(211)) xor (layer5_outputs(1058)));
    layer6_outputs(7048) <= not(layer5_outputs(230));
    layer6_outputs(7049) <= not(layer5_outputs(2971));
    layer6_outputs(7050) <= layer5_outputs(4899);
    layer6_outputs(7051) <= not((layer5_outputs(6891)) or (layer5_outputs(2985)));
    layer6_outputs(7052) <= layer5_outputs(2429);
    layer6_outputs(7053) <= not(layer5_outputs(6105));
    layer6_outputs(7054) <= not(layer5_outputs(4073));
    layer6_outputs(7055) <= not((layer5_outputs(6157)) or (layer5_outputs(827)));
    layer6_outputs(7056) <= layer5_outputs(3844);
    layer6_outputs(7057) <= not(layer5_outputs(1671)) or (layer5_outputs(6901));
    layer6_outputs(7058) <= layer5_outputs(4299);
    layer6_outputs(7059) <= layer5_outputs(7236);
    layer6_outputs(7060) <= (layer5_outputs(2672)) or (layer5_outputs(4946));
    layer6_outputs(7061) <= layer5_outputs(6543);
    layer6_outputs(7062) <= (layer5_outputs(6327)) xor (layer5_outputs(3984));
    layer6_outputs(7063) <= not((layer5_outputs(6313)) xor (layer5_outputs(5230)));
    layer6_outputs(7064) <= (layer5_outputs(5295)) xor (layer5_outputs(4469));
    layer6_outputs(7065) <= (layer5_outputs(873)) or (layer5_outputs(7174));
    layer6_outputs(7066) <= not(layer5_outputs(5504));
    layer6_outputs(7067) <= layer5_outputs(5146);
    layer6_outputs(7068) <= not(layer5_outputs(2438));
    layer6_outputs(7069) <= not((layer5_outputs(2580)) and (layer5_outputs(3504)));
    layer6_outputs(7070) <= not(layer5_outputs(1414)) or (layer5_outputs(834));
    layer6_outputs(7071) <= layer5_outputs(3082);
    layer6_outputs(7072) <= not(layer5_outputs(4378));
    layer6_outputs(7073) <= layer5_outputs(2686);
    layer6_outputs(7074) <= not(layer5_outputs(7210)) or (layer5_outputs(7188));
    layer6_outputs(7075) <= (layer5_outputs(1485)) and not (layer5_outputs(918));
    layer6_outputs(7076) <= (layer5_outputs(6469)) and not (layer5_outputs(1662));
    layer6_outputs(7077) <= not(layer5_outputs(910)) or (layer5_outputs(1324));
    layer6_outputs(7078) <= (layer5_outputs(887)) and not (layer5_outputs(5668));
    layer6_outputs(7079) <= not((layer5_outputs(4530)) xor (layer5_outputs(3139)));
    layer6_outputs(7080) <= layer5_outputs(7545);
    layer6_outputs(7081) <= not((layer5_outputs(4603)) xor (layer5_outputs(497)));
    layer6_outputs(7082) <= (layer5_outputs(6359)) xor (layer5_outputs(1769));
    layer6_outputs(7083) <= (layer5_outputs(4260)) xor (layer5_outputs(748));
    layer6_outputs(7084) <= layer5_outputs(796);
    layer6_outputs(7085) <= layer5_outputs(7444);
    layer6_outputs(7086) <= layer5_outputs(2591);
    layer6_outputs(7087) <= layer5_outputs(7194);
    layer6_outputs(7088) <= not(layer5_outputs(6581)) or (layer5_outputs(5158));
    layer6_outputs(7089) <= layer5_outputs(4702);
    layer6_outputs(7090) <= layer5_outputs(284);
    layer6_outputs(7091) <= not(layer5_outputs(6378));
    layer6_outputs(7092) <= not(layer5_outputs(453));
    layer6_outputs(7093) <= (layer5_outputs(362)) or (layer5_outputs(4218));
    layer6_outputs(7094) <= not(layer5_outputs(5088));
    layer6_outputs(7095) <= layer5_outputs(916);
    layer6_outputs(7096) <= (layer5_outputs(1776)) and not (layer5_outputs(2789));
    layer6_outputs(7097) <= not(layer5_outputs(4478)) or (layer5_outputs(207));
    layer6_outputs(7098) <= not(layer5_outputs(1920));
    layer6_outputs(7099) <= (layer5_outputs(1346)) and not (layer5_outputs(2146));
    layer6_outputs(7100) <= (layer5_outputs(1000)) xor (layer5_outputs(123));
    layer6_outputs(7101) <= not(layer5_outputs(6038));
    layer6_outputs(7102) <= not((layer5_outputs(1068)) xor (layer5_outputs(6766)));
    layer6_outputs(7103) <= layer5_outputs(6602);
    layer6_outputs(7104) <= not(layer5_outputs(1570));
    layer6_outputs(7105) <= not((layer5_outputs(6683)) xor (layer5_outputs(1204)));
    layer6_outputs(7106) <= not(layer5_outputs(6031)) or (layer5_outputs(6542));
    layer6_outputs(7107) <= layer5_outputs(75);
    layer6_outputs(7108) <= layer5_outputs(3949);
    layer6_outputs(7109) <= not(layer5_outputs(3658));
    layer6_outputs(7110) <= not(layer5_outputs(1903));
    layer6_outputs(7111) <= layer5_outputs(2192);
    layer6_outputs(7112) <= not(layer5_outputs(5502));
    layer6_outputs(7113) <= not((layer5_outputs(374)) or (layer5_outputs(2234)));
    layer6_outputs(7114) <= not((layer5_outputs(4942)) and (layer5_outputs(5263)));
    layer6_outputs(7115) <= (layer5_outputs(6661)) or (layer5_outputs(2282));
    layer6_outputs(7116) <= (layer5_outputs(3682)) and (layer5_outputs(6248));
    layer6_outputs(7117) <= layer5_outputs(821);
    layer6_outputs(7118) <= not(layer5_outputs(5640));
    layer6_outputs(7119) <= (layer5_outputs(5604)) and (layer5_outputs(7454));
    layer6_outputs(7120) <= not(layer5_outputs(2972));
    layer6_outputs(7121) <= layer5_outputs(4274);
    layer6_outputs(7122) <= not(layer5_outputs(3019)) or (layer5_outputs(2662));
    layer6_outputs(7123) <= layer5_outputs(1661);
    layer6_outputs(7124) <= not(layer5_outputs(7524));
    layer6_outputs(7125) <= (layer5_outputs(3770)) xor (layer5_outputs(404));
    layer6_outputs(7126) <= not(layer5_outputs(452));
    layer6_outputs(7127) <= layer5_outputs(2745);
    layer6_outputs(7128) <= layer5_outputs(3538);
    layer6_outputs(7129) <= layer5_outputs(6657);
    layer6_outputs(7130) <= not(layer5_outputs(5834));
    layer6_outputs(7131) <= layer5_outputs(3172);
    layer6_outputs(7132) <= (layer5_outputs(2567)) or (layer5_outputs(4347));
    layer6_outputs(7133) <= not(layer5_outputs(1514));
    layer6_outputs(7134) <= not((layer5_outputs(2970)) xor (layer5_outputs(1330)));
    layer6_outputs(7135) <= not(layer5_outputs(6764));
    layer6_outputs(7136) <= layer5_outputs(6153);
    layer6_outputs(7137) <= layer5_outputs(4640);
    layer6_outputs(7138) <= not(layer5_outputs(4722));
    layer6_outputs(7139) <= (layer5_outputs(4449)) or (layer5_outputs(5086));
    layer6_outputs(7140) <= not((layer5_outputs(2229)) xor (layer5_outputs(6641)));
    layer6_outputs(7141) <= not(layer5_outputs(4309)) or (layer5_outputs(62));
    layer6_outputs(7142) <= not((layer5_outputs(1303)) xor (layer5_outputs(5900)));
    layer6_outputs(7143) <= not(layer5_outputs(3769));
    layer6_outputs(7144) <= layer5_outputs(6417);
    layer6_outputs(7145) <= layer5_outputs(1912);
    layer6_outputs(7146) <= layer5_outputs(7634);
    layer6_outputs(7147) <= '0';
    layer6_outputs(7148) <= not((layer5_outputs(1006)) xor (layer5_outputs(338)));
    layer6_outputs(7149) <= not(layer5_outputs(5537)) or (layer5_outputs(2698));
    layer6_outputs(7150) <= not(layer5_outputs(6759)) or (layer5_outputs(281));
    layer6_outputs(7151) <= not(layer5_outputs(1457));
    layer6_outputs(7152) <= not(layer5_outputs(7619));
    layer6_outputs(7153) <= layer5_outputs(3087);
    layer6_outputs(7154) <= layer5_outputs(6225);
    layer6_outputs(7155) <= not((layer5_outputs(6218)) xor (layer5_outputs(4038)));
    layer6_outputs(7156) <= (layer5_outputs(3079)) and (layer5_outputs(6850));
    layer6_outputs(7157) <= not(layer5_outputs(865));
    layer6_outputs(7158) <= not(layer5_outputs(1332));
    layer6_outputs(7159) <= not(layer5_outputs(608));
    layer6_outputs(7160) <= layer5_outputs(210);
    layer6_outputs(7161) <= layer5_outputs(2241);
    layer6_outputs(7162) <= not(layer5_outputs(1428));
    layer6_outputs(7163) <= not(layer5_outputs(6874));
    layer6_outputs(7164) <= (layer5_outputs(1614)) xor (layer5_outputs(641));
    layer6_outputs(7165) <= not(layer5_outputs(5355));
    layer6_outputs(7166) <= layer5_outputs(6706);
    layer6_outputs(7167) <= (layer5_outputs(2291)) and (layer5_outputs(4792));
    layer6_outputs(7168) <= (layer5_outputs(4978)) and not (layer5_outputs(4364));
    layer6_outputs(7169) <= not((layer5_outputs(6350)) and (layer5_outputs(2337)));
    layer6_outputs(7170) <= not((layer5_outputs(6284)) or (layer5_outputs(3353)));
    layer6_outputs(7171) <= not((layer5_outputs(4777)) or (layer5_outputs(5009)));
    layer6_outputs(7172) <= (layer5_outputs(3395)) and not (layer5_outputs(578));
    layer6_outputs(7173) <= not(layer5_outputs(6326));
    layer6_outputs(7174) <= layer5_outputs(3170);
    layer6_outputs(7175) <= not(layer5_outputs(7176));
    layer6_outputs(7176) <= not(layer5_outputs(1829));
    layer6_outputs(7177) <= not((layer5_outputs(6174)) xor (layer5_outputs(5484)));
    layer6_outputs(7178) <= not(layer5_outputs(7404));
    layer6_outputs(7179) <= not(layer5_outputs(3330));
    layer6_outputs(7180) <= (layer5_outputs(4427)) or (layer5_outputs(449));
    layer6_outputs(7181) <= layer5_outputs(970);
    layer6_outputs(7182) <= (layer5_outputs(5547)) xor (layer5_outputs(2960));
    layer6_outputs(7183) <= not(layer5_outputs(3199));
    layer6_outputs(7184) <= (layer5_outputs(1278)) xor (layer5_outputs(2117));
    layer6_outputs(7185) <= not(layer5_outputs(1937));
    layer6_outputs(7186) <= (layer5_outputs(6562)) xor (layer5_outputs(5272));
    layer6_outputs(7187) <= not((layer5_outputs(4760)) xor (layer5_outputs(2523)));
    layer6_outputs(7188) <= not(layer5_outputs(3878));
    layer6_outputs(7189) <= not(layer5_outputs(6902)) or (layer5_outputs(6735));
    layer6_outputs(7190) <= (layer5_outputs(17)) or (layer5_outputs(3692));
    layer6_outputs(7191) <= layer5_outputs(422);
    layer6_outputs(7192) <= layer5_outputs(1215);
    layer6_outputs(7193) <= not(layer5_outputs(1137));
    layer6_outputs(7194) <= not(layer5_outputs(4116)) or (layer5_outputs(165));
    layer6_outputs(7195) <= layer5_outputs(7083);
    layer6_outputs(7196) <= (layer5_outputs(1147)) and (layer5_outputs(5003));
    layer6_outputs(7197) <= not(layer5_outputs(5029));
    layer6_outputs(7198) <= not(layer5_outputs(81)) or (layer5_outputs(2852));
    layer6_outputs(7199) <= not(layer5_outputs(5667));
    layer6_outputs(7200) <= layer5_outputs(2816);
    layer6_outputs(7201) <= (layer5_outputs(5633)) and not (layer5_outputs(4599));
    layer6_outputs(7202) <= not(layer5_outputs(6720)) or (layer5_outputs(3966));
    layer6_outputs(7203) <= (layer5_outputs(1415)) and not (layer5_outputs(3810));
    layer6_outputs(7204) <= not(layer5_outputs(4020));
    layer6_outputs(7205) <= layer5_outputs(3620);
    layer6_outputs(7206) <= layer5_outputs(4140);
    layer6_outputs(7207) <= not(layer5_outputs(2899));
    layer6_outputs(7208) <= not(layer5_outputs(956));
    layer6_outputs(7209) <= not((layer5_outputs(5761)) xor (layer5_outputs(1575)));
    layer6_outputs(7210) <= not((layer5_outputs(6952)) and (layer5_outputs(7607)));
    layer6_outputs(7211) <= layer5_outputs(6638);
    layer6_outputs(7212) <= not(layer5_outputs(7350));
    layer6_outputs(7213) <= not(layer5_outputs(879));
    layer6_outputs(7214) <= layer5_outputs(7452);
    layer6_outputs(7215) <= layer5_outputs(3500);
    layer6_outputs(7216) <= layer5_outputs(7582);
    layer6_outputs(7217) <= layer5_outputs(6551);
    layer6_outputs(7218) <= layer5_outputs(3121);
    layer6_outputs(7219) <= not(layer5_outputs(7277)) or (layer5_outputs(5096));
    layer6_outputs(7220) <= not((layer5_outputs(4822)) xor (layer5_outputs(5056)));
    layer6_outputs(7221) <= layer5_outputs(5158);
    layer6_outputs(7222) <= (layer5_outputs(4397)) xor (layer5_outputs(2785));
    layer6_outputs(7223) <= (layer5_outputs(7)) and not (layer5_outputs(6772));
    layer6_outputs(7224) <= (layer5_outputs(3079)) xor (layer5_outputs(6131));
    layer6_outputs(7225) <= not(layer5_outputs(1787));
    layer6_outputs(7226) <= not(layer5_outputs(7638));
    layer6_outputs(7227) <= (layer5_outputs(2708)) and not (layer5_outputs(830));
    layer6_outputs(7228) <= (layer5_outputs(7172)) and (layer5_outputs(2260));
    layer6_outputs(7229) <= layer5_outputs(1375);
    layer6_outputs(7230) <= layer5_outputs(7240);
    layer6_outputs(7231) <= (layer5_outputs(6643)) and not (layer5_outputs(2445));
    layer6_outputs(7232) <= not(layer5_outputs(6047)) or (layer5_outputs(7090));
    layer6_outputs(7233) <= layer5_outputs(2812);
    layer6_outputs(7234) <= not(layer5_outputs(5790)) or (layer5_outputs(4949));
    layer6_outputs(7235) <= layer5_outputs(37);
    layer6_outputs(7236) <= (layer5_outputs(1488)) xor (layer5_outputs(1433));
    layer6_outputs(7237) <= (layer5_outputs(3182)) and (layer5_outputs(3571));
    layer6_outputs(7238) <= not((layer5_outputs(5394)) or (layer5_outputs(671)));
    layer6_outputs(7239) <= layer5_outputs(4619);
    layer6_outputs(7240) <= layer5_outputs(4371);
    layer6_outputs(7241) <= not((layer5_outputs(7478)) xor (layer5_outputs(65)));
    layer6_outputs(7242) <= (layer5_outputs(6234)) xor (layer5_outputs(3835));
    layer6_outputs(7243) <= not(layer5_outputs(5760));
    layer6_outputs(7244) <= not(layer5_outputs(4074));
    layer6_outputs(7245) <= not((layer5_outputs(5571)) and (layer5_outputs(2443)));
    layer6_outputs(7246) <= not((layer5_outputs(7626)) and (layer5_outputs(6435)));
    layer6_outputs(7247) <= not(layer5_outputs(2436));
    layer6_outputs(7248) <= (layer5_outputs(5236)) xor (layer5_outputs(1972));
    layer6_outputs(7249) <= (layer5_outputs(4397)) and not (layer5_outputs(3561));
    layer6_outputs(7250) <= layer5_outputs(4541);
    layer6_outputs(7251) <= not((layer5_outputs(5206)) or (layer5_outputs(5188)));
    layer6_outputs(7252) <= layer5_outputs(3283);
    layer6_outputs(7253) <= (layer5_outputs(5605)) xor (layer5_outputs(1477));
    layer6_outputs(7254) <= (layer5_outputs(3983)) and not (layer5_outputs(562));
    layer6_outputs(7255) <= not((layer5_outputs(4288)) xor (layer5_outputs(1647)));
    layer6_outputs(7256) <= not((layer5_outputs(644)) xor (layer5_outputs(1015)));
    layer6_outputs(7257) <= (layer5_outputs(1682)) and not (layer5_outputs(6506));
    layer6_outputs(7258) <= not(layer5_outputs(7139));
    layer6_outputs(7259) <= layer5_outputs(3848);
    layer6_outputs(7260) <= not(layer5_outputs(122));
    layer6_outputs(7261) <= not(layer5_outputs(6066));
    layer6_outputs(7262) <= not((layer5_outputs(7638)) or (layer5_outputs(7471)));
    layer6_outputs(7263) <= (layer5_outputs(7220)) and not (layer5_outputs(5768));
    layer6_outputs(7264) <= not(layer5_outputs(543));
    layer6_outputs(7265) <= not((layer5_outputs(4288)) or (layer5_outputs(7316)));
    layer6_outputs(7266) <= (layer5_outputs(5288)) xor (layer5_outputs(6688));
    layer6_outputs(7267) <= layer5_outputs(4915);
    layer6_outputs(7268) <= not(layer5_outputs(1165));
    layer6_outputs(7269) <= not(layer5_outputs(7138));
    layer6_outputs(7270) <= layer5_outputs(1619);
    layer6_outputs(7271) <= (layer5_outputs(1299)) or (layer5_outputs(7331));
    layer6_outputs(7272) <= (layer5_outputs(6318)) xor (layer5_outputs(1988));
    layer6_outputs(7273) <= '0';
    layer6_outputs(7274) <= (layer5_outputs(3815)) xor (layer5_outputs(6832));
    layer6_outputs(7275) <= layer5_outputs(5715);
    layer6_outputs(7276) <= not(layer5_outputs(4036));
    layer6_outputs(7277) <= layer5_outputs(711);
    layer6_outputs(7278) <= (layer5_outputs(5727)) xor (layer5_outputs(1632));
    layer6_outputs(7279) <= (layer5_outputs(1416)) or (layer5_outputs(118));
    layer6_outputs(7280) <= not(layer5_outputs(5971));
    layer6_outputs(7281) <= layer5_outputs(2650);
    layer6_outputs(7282) <= (layer5_outputs(6852)) and not (layer5_outputs(1672));
    layer6_outputs(7283) <= layer5_outputs(4433);
    layer6_outputs(7284) <= (layer5_outputs(410)) and not (layer5_outputs(4402));
    layer6_outputs(7285) <= not((layer5_outputs(766)) xor (layer5_outputs(4129)));
    layer6_outputs(7286) <= not(layer5_outputs(5179)) or (layer5_outputs(1343));
    layer6_outputs(7287) <= (layer5_outputs(4490)) or (layer5_outputs(2368));
    layer6_outputs(7288) <= (layer5_outputs(2689)) and not (layer5_outputs(5005));
    layer6_outputs(7289) <= not(layer5_outputs(227));
    layer6_outputs(7290) <= not(layer5_outputs(5147)) or (layer5_outputs(90));
    layer6_outputs(7291) <= not(layer5_outputs(7285));
    layer6_outputs(7292) <= (layer5_outputs(6877)) xor (layer5_outputs(6121));
    layer6_outputs(7293) <= layer5_outputs(4349);
    layer6_outputs(7294) <= (layer5_outputs(527)) and not (layer5_outputs(3471));
    layer6_outputs(7295) <= (layer5_outputs(6078)) and not (layer5_outputs(2840));
    layer6_outputs(7296) <= (layer5_outputs(4928)) or (layer5_outputs(6889));
    layer6_outputs(7297) <= (layer5_outputs(4505)) xor (layer5_outputs(7238));
    layer6_outputs(7298) <= layer5_outputs(6787);
    layer6_outputs(7299) <= not(layer5_outputs(6133)) or (layer5_outputs(6714));
    layer6_outputs(7300) <= layer5_outputs(4739);
    layer6_outputs(7301) <= layer5_outputs(3651);
    layer6_outputs(7302) <= (layer5_outputs(2534)) and not (layer5_outputs(5083));
    layer6_outputs(7303) <= (layer5_outputs(4098)) or (layer5_outputs(198));
    layer6_outputs(7304) <= not(layer5_outputs(6817));
    layer6_outputs(7305) <= not(layer5_outputs(4509));
    layer6_outputs(7306) <= not(layer5_outputs(2183));
    layer6_outputs(7307) <= not(layer5_outputs(5652));
    layer6_outputs(7308) <= layer5_outputs(4481);
    layer6_outputs(7309) <= not(layer5_outputs(154));
    layer6_outputs(7310) <= not(layer5_outputs(987));
    layer6_outputs(7311) <= not((layer5_outputs(3950)) and (layer5_outputs(5585)));
    layer6_outputs(7312) <= not((layer5_outputs(4583)) xor (layer5_outputs(7113)));
    layer6_outputs(7313) <= layer5_outputs(5530);
    layer6_outputs(7314) <= layer5_outputs(6321);
    layer6_outputs(7315) <= not(layer5_outputs(1110));
    layer6_outputs(7316) <= not(layer5_outputs(2150));
    layer6_outputs(7317) <= not(layer5_outputs(99)) or (layer5_outputs(3860));
    layer6_outputs(7318) <= not(layer5_outputs(4817));
    layer6_outputs(7319) <= (layer5_outputs(78)) and not (layer5_outputs(5663));
    layer6_outputs(7320) <= not(layer5_outputs(5746)) or (layer5_outputs(1183));
    layer6_outputs(7321) <= not(layer5_outputs(2104));
    layer6_outputs(7322) <= (layer5_outputs(4101)) and not (layer5_outputs(6986));
    layer6_outputs(7323) <= layer5_outputs(5329);
    layer6_outputs(7324) <= layer5_outputs(6411);
    layer6_outputs(7325) <= not(layer5_outputs(2642));
    layer6_outputs(7326) <= not(layer5_outputs(6049));
    layer6_outputs(7327) <= (layer5_outputs(1471)) or (layer5_outputs(5093));
    layer6_outputs(7328) <= (layer5_outputs(1964)) xor (layer5_outputs(6802));
    layer6_outputs(7329) <= not(layer5_outputs(542)) or (layer5_outputs(6525));
    layer6_outputs(7330) <= not((layer5_outputs(7253)) xor (layer5_outputs(1590)));
    layer6_outputs(7331) <= not(layer5_outputs(5805));
    layer6_outputs(7332) <= not(layer5_outputs(151));
    layer6_outputs(7333) <= layer5_outputs(6577);
    layer6_outputs(7334) <= layer5_outputs(2560);
    layer6_outputs(7335) <= not(layer5_outputs(5793));
    layer6_outputs(7336) <= not(layer5_outputs(2165));
    layer6_outputs(7337) <= (layer5_outputs(3142)) and not (layer5_outputs(2677));
    layer6_outputs(7338) <= layer5_outputs(53);
    layer6_outputs(7339) <= not((layer5_outputs(134)) or (layer5_outputs(691)));
    layer6_outputs(7340) <= layer5_outputs(3456);
    layer6_outputs(7341) <= not(layer5_outputs(1887));
    layer6_outputs(7342) <= layer5_outputs(4487);
    layer6_outputs(7343) <= (layer5_outputs(279)) or (layer5_outputs(6395));
    layer6_outputs(7344) <= (layer5_outputs(2486)) or (layer5_outputs(3399));
    layer6_outputs(7345) <= not(layer5_outputs(5164));
    layer6_outputs(7346) <= not((layer5_outputs(2620)) xor (layer5_outputs(5061)));
    layer6_outputs(7347) <= not(layer5_outputs(5636));
    layer6_outputs(7348) <= not((layer5_outputs(3247)) or (layer5_outputs(5837)));
    layer6_outputs(7349) <= (layer5_outputs(1519)) and not (layer5_outputs(1554));
    layer6_outputs(7350) <= layer5_outputs(4422);
    layer6_outputs(7351) <= not(layer5_outputs(1299));
    layer6_outputs(7352) <= not((layer5_outputs(4447)) xor (layer5_outputs(518)));
    layer6_outputs(7353) <= layer5_outputs(4988);
    layer6_outputs(7354) <= not(layer5_outputs(4365)) or (layer5_outputs(2025));
    layer6_outputs(7355) <= (layer5_outputs(4921)) and not (layer5_outputs(2109));
    layer6_outputs(7356) <= not(layer5_outputs(2835));
    layer6_outputs(7357) <= (layer5_outputs(6321)) and not (layer5_outputs(4811));
    layer6_outputs(7358) <= not((layer5_outputs(7575)) xor (layer5_outputs(4388)));
    layer6_outputs(7359) <= not(layer5_outputs(6569)) or (layer5_outputs(5751));
    layer6_outputs(7360) <= not((layer5_outputs(4945)) xor (layer5_outputs(1383)));
    layer6_outputs(7361) <= not(layer5_outputs(6142));
    layer6_outputs(7362) <= (layer5_outputs(666)) and not (layer5_outputs(239));
    layer6_outputs(7363) <= (layer5_outputs(5341)) xor (layer5_outputs(3224));
    layer6_outputs(7364) <= not((layer5_outputs(5514)) xor (layer5_outputs(307)));
    layer6_outputs(7365) <= not(layer5_outputs(3084));
    layer6_outputs(7366) <= not(layer5_outputs(999));
    layer6_outputs(7367) <= layer5_outputs(3486);
    layer6_outputs(7368) <= not(layer5_outputs(3489));
    layer6_outputs(7369) <= layer5_outputs(4616);
    layer6_outputs(7370) <= layer5_outputs(6527);
    layer6_outputs(7371) <= (layer5_outputs(611)) and (layer5_outputs(5433));
    layer6_outputs(7372) <= not(layer5_outputs(7235));
    layer6_outputs(7373) <= not(layer5_outputs(5019));
    layer6_outputs(7374) <= layer5_outputs(7587);
    layer6_outputs(7375) <= (layer5_outputs(1156)) xor (layer5_outputs(6164));
    layer6_outputs(7376) <= not((layer5_outputs(4917)) or (layer5_outputs(4826)));
    layer6_outputs(7377) <= not(layer5_outputs(2287)) or (layer5_outputs(5359));
    layer6_outputs(7378) <= not(layer5_outputs(4926));
    layer6_outputs(7379) <= not(layer5_outputs(6264));
    layer6_outputs(7380) <= layer5_outputs(3864);
    layer6_outputs(7381) <= (layer5_outputs(5864)) and not (layer5_outputs(5015));
    layer6_outputs(7382) <= (layer5_outputs(1461)) and not (layer5_outputs(5410));
    layer6_outputs(7383) <= layer5_outputs(1372);
    layer6_outputs(7384) <= not(layer5_outputs(3469));
    layer6_outputs(7385) <= not((layer5_outputs(1421)) xor (layer5_outputs(1087)));
    layer6_outputs(7386) <= not(layer5_outputs(6055));
    layer6_outputs(7387) <= (layer5_outputs(3563)) and not (layer5_outputs(7462));
    layer6_outputs(7388) <= not(layer5_outputs(858)) or (layer5_outputs(4121));
    layer6_outputs(7389) <= not(layer5_outputs(7422));
    layer6_outputs(7390) <= not(layer5_outputs(4103));
    layer6_outputs(7391) <= layer5_outputs(3);
    layer6_outputs(7392) <= not(layer5_outputs(7208));
    layer6_outputs(7393) <= (layer5_outputs(3492)) or (layer5_outputs(369));
    layer6_outputs(7394) <= layer5_outputs(1597);
    layer6_outputs(7395) <= layer5_outputs(3665);
    layer6_outputs(7396) <= not((layer5_outputs(4264)) xor (layer5_outputs(3513)));
    layer6_outputs(7397) <= layer5_outputs(6811);
    layer6_outputs(7398) <= not((layer5_outputs(1004)) xor (layer5_outputs(7364)));
    layer6_outputs(7399) <= not(layer5_outputs(7168));
    layer6_outputs(7400) <= (layer5_outputs(2389)) and not (layer5_outputs(5507));
    layer6_outputs(7401) <= not((layer5_outputs(5349)) or (layer5_outputs(302)));
    layer6_outputs(7402) <= not(layer5_outputs(3731)) or (layer5_outputs(7594));
    layer6_outputs(7403) <= not(layer5_outputs(5470));
    layer6_outputs(7404) <= (layer5_outputs(1969)) xor (layer5_outputs(718));
    layer6_outputs(7405) <= (layer5_outputs(14)) xor (layer5_outputs(6447));
    layer6_outputs(7406) <= layer5_outputs(3933);
    layer6_outputs(7407) <= (layer5_outputs(2627)) xor (layer5_outputs(3130));
    layer6_outputs(7408) <= (layer5_outputs(7385)) xor (layer5_outputs(3606));
    layer6_outputs(7409) <= (layer5_outputs(5006)) or (layer5_outputs(2110));
    layer6_outputs(7410) <= not((layer5_outputs(795)) or (layer5_outputs(6181)));
    layer6_outputs(7411) <= layer5_outputs(6524);
    layer6_outputs(7412) <= layer5_outputs(4303);
    layer6_outputs(7413) <= not((layer5_outputs(4497)) and (layer5_outputs(4966)));
    layer6_outputs(7414) <= (layer5_outputs(753)) and (layer5_outputs(6574));
    layer6_outputs(7415) <= (layer5_outputs(6231)) and not (layer5_outputs(1304));
    layer6_outputs(7416) <= (layer5_outputs(2191)) and (layer5_outputs(5079));
    layer6_outputs(7417) <= not(layer5_outputs(2040));
    layer6_outputs(7418) <= layer5_outputs(1239);
    layer6_outputs(7419) <= (layer5_outputs(5670)) and not (layer5_outputs(6909));
    layer6_outputs(7420) <= (layer5_outputs(4213)) and not (layer5_outputs(64));
    layer6_outputs(7421) <= not(layer5_outputs(6838));
    layer6_outputs(7422) <= not(layer5_outputs(1640));
    layer6_outputs(7423) <= layer5_outputs(5143);
    layer6_outputs(7424) <= layer5_outputs(7447);
    layer6_outputs(7425) <= layer5_outputs(6347);
    layer6_outputs(7426) <= not((layer5_outputs(2030)) xor (layer5_outputs(2683)));
    layer6_outputs(7427) <= (layer5_outputs(2742)) and (layer5_outputs(5665));
    layer6_outputs(7428) <= (layer5_outputs(4731)) or (layer5_outputs(4658));
    layer6_outputs(7429) <= not(layer5_outputs(2684));
    layer6_outputs(7430) <= not((layer5_outputs(3078)) or (layer5_outputs(3490)));
    layer6_outputs(7431) <= layer5_outputs(2950);
    layer6_outputs(7432) <= layer5_outputs(5073);
    layer6_outputs(7433) <= layer5_outputs(4742);
    layer6_outputs(7434) <= layer5_outputs(432);
    layer6_outputs(7435) <= not(layer5_outputs(1549)) or (layer5_outputs(5942));
    layer6_outputs(7436) <= layer5_outputs(2145);
    layer6_outputs(7437) <= not(layer5_outputs(5795));
    layer6_outputs(7438) <= layer5_outputs(6352);
    layer6_outputs(7439) <= not(layer5_outputs(6101));
    layer6_outputs(7440) <= not(layer5_outputs(6951));
    layer6_outputs(7441) <= (layer5_outputs(3466)) xor (layer5_outputs(3814));
    layer6_outputs(7442) <= layer5_outputs(2995);
    layer6_outputs(7443) <= not(layer5_outputs(1619));
    layer6_outputs(7444) <= (layer5_outputs(7436)) or (layer5_outputs(6731));
    layer6_outputs(7445) <= '1';
    layer6_outputs(7446) <= layer5_outputs(3674);
    layer6_outputs(7447) <= layer5_outputs(2847);
    layer6_outputs(7448) <= not((layer5_outputs(7021)) and (layer5_outputs(906)));
    layer6_outputs(7449) <= not(layer5_outputs(4115));
    layer6_outputs(7450) <= not(layer5_outputs(5616)) or (layer5_outputs(6749));
    layer6_outputs(7451) <= not(layer5_outputs(6813));
    layer6_outputs(7452) <= layer5_outputs(752);
    layer6_outputs(7453) <= not(layer5_outputs(7274));
    layer6_outputs(7454) <= not(layer5_outputs(3978));
    layer6_outputs(7455) <= (layer5_outputs(5531)) xor (layer5_outputs(4224));
    layer6_outputs(7456) <= not(layer5_outputs(606));
    layer6_outputs(7457) <= layer5_outputs(1437);
    layer6_outputs(7458) <= (layer5_outputs(6121)) or (layer5_outputs(3339));
    layer6_outputs(7459) <= not((layer5_outputs(7609)) or (layer5_outputs(1972)));
    layer6_outputs(7460) <= (layer5_outputs(1008)) and not (layer5_outputs(2104));
    layer6_outputs(7461) <= not(layer5_outputs(2906));
    layer6_outputs(7462) <= layer5_outputs(4474);
    layer6_outputs(7463) <= (layer5_outputs(2992)) xor (layer5_outputs(1761));
    layer6_outputs(7464) <= layer5_outputs(3306);
    layer6_outputs(7465) <= (layer5_outputs(5270)) and not (layer5_outputs(891));
    layer6_outputs(7466) <= (layer5_outputs(7476)) and (layer5_outputs(1096));
    layer6_outputs(7467) <= not(layer5_outputs(1830));
    layer6_outputs(7468) <= layer5_outputs(1735);
    layer6_outputs(7469) <= (layer5_outputs(3760)) xor (layer5_outputs(798));
    layer6_outputs(7470) <= not(layer5_outputs(2804));
    layer6_outputs(7471) <= (layer5_outputs(4241)) and not (layer5_outputs(2694));
    layer6_outputs(7472) <= not((layer5_outputs(7222)) or (layer5_outputs(925)));
    layer6_outputs(7473) <= not(layer5_outputs(581)) or (layer5_outputs(6734));
    layer6_outputs(7474) <= (layer5_outputs(6698)) xor (layer5_outputs(2841));
    layer6_outputs(7475) <= not(layer5_outputs(274));
    layer6_outputs(7476) <= layer5_outputs(1436);
    layer6_outputs(7477) <= not((layer5_outputs(391)) xor (layer5_outputs(5118)));
    layer6_outputs(7478) <= (layer5_outputs(2314)) xor (layer5_outputs(4611));
    layer6_outputs(7479) <= not(layer5_outputs(4066)) or (layer5_outputs(4977));
    layer6_outputs(7480) <= layer5_outputs(7331);
    layer6_outputs(7481) <= (layer5_outputs(2974)) xor (layer5_outputs(3935));
    layer6_outputs(7482) <= not(layer5_outputs(4555));
    layer6_outputs(7483) <= not(layer5_outputs(4432));
    layer6_outputs(7484) <= (layer5_outputs(4115)) and not (layer5_outputs(2012));
    layer6_outputs(7485) <= not(layer5_outputs(171));
    layer6_outputs(7486) <= not(layer5_outputs(191));
    layer6_outputs(7487) <= not(layer5_outputs(1882));
    layer6_outputs(7488) <= not(layer5_outputs(4896)) or (layer5_outputs(6977));
    layer6_outputs(7489) <= layer5_outputs(6260);
    layer6_outputs(7490) <= (layer5_outputs(5525)) xor (layer5_outputs(3429));
    layer6_outputs(7491) <= layer5_outputs(5259);
    layer6_outputs(7492) <= '1';
    layer6_outputs(7493) <= not((layer5_outputs(2469)) xor (layer5_outputs(2095)));
    layer6_outputs(7494) <= not(layer5_outputs(656));
    layer6_outputs(7495) <= not((layer5_outputs(1958)) or (layer5_outputs(3813)));
    layer6_outputs(7496) <= layer5_outputs(393);
    layer6_outputs(7497) <= layer5_outputs(1755);
    layer6_outputs(7498) <= (layer5_outputs(2231)) or (layer5_outputs(6795));
    layer6_outputs(7499) <= layer5_outputs(3778);
    layer6_outputs(7500) <= layer5_outputs(5326);
    layer6_outputs(7501) <= not(layer5_outputs(6741)) or (layer5_outputs(7647));
    layer6_outputs(7502) <= (layer5_outputs(3440)) xor (layer5_outputs(282));
    layer6_outputs(7503) <= layer5_outputs(1594);
    layer6_outputs(7504) <= not(layer5_outputs(1230));
    layer6_outputs(7505) <= not(layer5_outputs(6390));
    layer6_outputs(7506) <= layer5_outputs(1841);
    layer6_outputs(7507) <= not(layer5_outputs(1392));
    layer6_outputs(7508) <= not(layer5_outputs(2372));
    layer6_outputs(7509) <= not(layer5_outputs(3027));
    layer6_outputs(7510) <= not((layer5_outputs(825)) or (layer5_outputs(5980)));
    layer6_outputs(7511) <= not((layer5_outputs(5458)) or (layer5_outputs(3852)));
    layer6_outputs(7512) <= layer5_outputs(6887);
    layer6_outputs(7513) <= (layer5_outputs(6027)) xor (layer5_outputs(3056));
    layer6_outputs(7514) <= not(layer5_outputs(6403)) or (layer5_outputs(7215));
    layer6_outputs(7515) <= layer5_outputs(7390);
    layer6_outputs(7516) <= not((layer5_outputs(2691)) and (layer5_outputs(6960)));
    layer6_outputs(7517) <= not((layer5_outputs(6229)) and (layer5_outputs(1992)));
    layer6_outputs(7518) <= not(layer5_outputs(1574));
    layer6_outputs(7519) <= (layer5_outputs(1074)) and (layer5_outputs(1369));
    layer6_outputs(7520) <= not((layer5_outputs(3161)) xor (layer5_outputs(2659)));
    layer6_outputs(7521) <= not(layer5_outputs(2383));
    layer6_outputs(7522) <= (layer5_outputs(7025)) and (layer5_outputs(5858));
    layer6_outputs(7523) <= (layer5_outputs(4206)) or (layer5_outputs(5019));
    layer6_outputs(7524) <= not((layer5_outputs(7257)) xor (layer5_outputs(1438)));
    layer6_outputs(7525) <= not(layer5_outputs(1572)) or (layer5_outputs(5867));
    layer6_outputs(7526) <= layer5_outputs(7376);
    layer6_outputs(7527) <= layer5_outputs(1155);
    layer6_outputs(7528) <= layer5_outputs(2343);
    layer6_outputs(7529) <= not((layer5_outputs(4230)) xor (layer5_outputs(3528)));
    layer6_outputs(7530) <= not((layer5_outputs(4652)) xor (layer5_outputs(7351)));
    layer6_outputs(7531) <= not(layer5_outputs(4038));
    layer6_outputs(7532) <= not(layer5_outputs(5899));
    layer6_outputs(7533) <= layer5_outputs(4466);
    layer6_outputs(7534) <= not(layer5_outputs(6757));
    layer6_outputs(7535) <= not(layer5_outputs(2743));
    layer6_outputs(7536) <= layer5_outputs(6812);
    layer6_outputs(7537) <= layer5_outputs(1886);
    layer6_outputs(7538) <= (layer5_outputs(4282)) xor (layer5_outputs(3206));
    layer6_outputs(7539) <= not((layer5_outputs(199)) or (layer5_outputs(4625)));
    layer6_outputs(7540) <= not(layer5_outputs(1450));
    layer6_outputs(7541) <= layer5_outputs(2099);
    layer6_outputs(7542) <= layer5_outputs(4666);
    layer6_outputs(7543) <= layer5_outputs(5626);
    layer6_outputs(7544) <= not(layer5_outputs(5225));
    layer6_outputs(7545) <= not(layer5_outputs(5650));
    layer6_outputs(7546) <= (layer5_outputs(6605)) or (layer5_outputs(6612));
    layer6_outputs(7547) <= not(layer5_outputs(2327));
    layer6_outputs(7548) <= layer5_outputs(3025);
    layer6_outputs(7549) <= not(layer5_outputs(1929)) or (layer5_outputs(7151));
    layer6_outputs(7550) <= (layer5_outputs(2778)) or (layer5_outputs(3862));
    layer6_outputs(7551) <= (layer5_outputs(4724)) xor (layer5_outputs(3243));
    layer6_outputs(7552) <= not((layer5_outputs(4411)) and (layer5_outputs(179)));
    layer6_outputs(7553) <= (layer5_outputs(829)) and not (layer5_outputs(516));
    layer6_outputs(7554) <= not(layer5_outputs(6223));
    layer6_outputs(7555) <= (layer5_outputs(4915)) xor (layer5_outputs(278));
    layer6_outputs(7556) <= layer5_outputs(3298);
    layer6_outputs(7557) <= layer5_outputs(7379);
    layer6_outputs(7558) <= not(layer5_outputs(2017)) or (layer5_outputs(3229));
    layer6_outputs(7559) <= layer5_outputs(7179);
    layer6_outputs(7560) <= layer5_outputs(6622);
    layer6_outputs(7561) <= layer5_outputs(1999);
    layer6_outputs(7562) <= not(layer5_outputs(5098));
    layer6_outputs(7563) <= layer5_outputs(7357);
    layer6_outputs(7564) <= layer5_outputs(1212);
    layer6_outputs(7565) <= not(layer5_outputs(5177));
    layer6_outputs(7566) <= not(layer5_outputs(6063));
    layer6_outputs(7567) <= (layer5_outputs(2064)) xor (layer5_outputs(5597));
    layer6_outputs(7568) <= (layer5_outputs(995)) xor (layer5_outputs(846));
    layer6_outputs(7569) <= not((layer5_outputs(1561)) xor (layer5_outputs(7074)));
    layer6_outputs(7570) <= layer5_outputs(4095);
    layer6_outputs(7571) <= not(layer5_outputs(7231));
    layer6_outputs(7572) <= (layer5_outputs(6770)) or (layer5_outputs(7181));
    layer6_outputs(7573) <= not(layer5_outputs(1778));
    layer6_outputs(7574) <= (layer5_outputs(5935)) xor (layer5_outputs(3475));
    layer6_outputs(7575) <= not(layer5_outputs(1642));
    layer6_outputs(7576) <= (layer5_outputs(6799)) or (layer5_outputs(1229));
    layer6_outputs(7577) <= not(layer5_outputs(5063));
    layer6_outputs(7578) <= layer5_outputs(2654);
    layer6_outputs(7579) <= layer5_outputs(6007);
    layer6_outputs(7580) <= (layer5_outputs(7085)) and (layer5_outputs(4739));
    layer6_outputs(7581) <= (layer5_outputs(2136)) xor (layer5_outputs(3089));
    layer6_outputs(7582) <= (layer5_outputs(2960)) and not (layer5_outputs(6239));
    layer6_outputs(7583) <= (layer5_outputs(5040)) and not (layer5_outputs(770));
    layer6_outputs(7584) <= (layer5_outputs(570)) or (layer5_outputs(3120));
    layer6_outputs(7585) <= not(layer5_outputs(663));
    layer6_outputs(7586) <= (layer5_outputs(4735)) or (layer5_outputs(4609));
    layer6_outputs(7587) <= (layer5_outputs(1335)) and (layer5_outputs(6387));
    layer6_outputs(7588) <= (layer5_outputs(5984)) and not (layer5_outputs(7296));
    layer6_outputs(7589) <= not(layer5_outputs(3940));
    layer6_outputs(7590) <= not(layer5_outputs(7259));
    layer6_outputs(7591) <= layer5_outputs(4247);
    layer6_outputs(7592) <= layer5_outputs(4710);
    layer6_outputs(7593) <= (layer5_outputs(1553)) and not (layer5_outputs(4790));
    layer6_outputs(7594) <= layer5_outputs(6815);
    layer6_outputs(7595) <= not(layer5_outputs(5639));
    layer6_outputs(7596) <= not(layer5_outputs(2562)) or (layer5_outputs(705));
    layer6_outputs(7597) <= (layer5_outputs(1041)) xor (layer5_outputs(1218));
    layer6_outputs(7598) <= not((layer5_outputs(7128)) and (layer5_outputs(5658)));
    layer6_outputs(7599) <= not(layer5_outputs(4868));
    layer6_outputs(7600) <= layer5_outputs(128);
    layer6_outputs(7601) <= not(layer5_outputs(1184)) or (layer5_outputs(417));
    layer6_outputs(7602) <= (layer5_outputs(2212)) xor (layer5_outputs(1661));
    layer6_outputs(7603) <= not(layer5_outputs(5622));
    layer6_outputs(7604) <= '0';
    layer6_outputs(7605) <= (layer5_outputs(2201)) and not (layer5_outputs(3517));
    layer6_outputs(7606) <= (layer5_outputs(5690)) xor (layer5_outputs(3812));
    layer6_outputs(7607) <= layer5_outputs(6333);
    layer6_outputs(7608) <= layer5_outputs(6550);
    layer6_outputs(7609) <= not(layer5_outputs(3565));
    layer6_outputs(7610) <= not(layer5_outputs(3315));
    layer6_outputs(7611) <= (layer5_outputs(7445)) and not (layer5_outputs(6585));
    layer6_outputs(7612) <= layer5_outputs(5707);
    layer6_outputs(7613) <= not(layer5_outputs(481)) or (layer5_outputs(6112));
    layer6_outputs(7614) <= '1';
    layer6_outputs(7615) <= not(layer5_outputs(792));
    layer6_outputs(7616) <= not(layer5_outputs(2862));
    layer6_outputs(7617) <= layer5_outputs(7061);
    layer6_outputs(7618) <= not(layer5_outputs(3630));
    layer6_outputs(7619) <= (layer5_outputs(3117)) xor (layer5_outputs(2233));
    layer6_outputs(7620) <= not(layer5_outputs(2323));
    layer6_outputs(7621) <= not(layer5_outputs(5008)) or (layer5_outputs(1479));
    layer6_outputs(7622) <= not(layer5_outputs(6319));
    layer6_outputs(7623) <= (layer5_outputs(743)) and (layer5_outputs(4957));
    layer6_outputs(7624) <= layer5_outputs(6597);
    layer6_outputs(7625) <= not((layer5_outputs(7178)) and (layer5_outputs(3601)));
    layer6_outputs(7626) <= (layer5_outputs(492)) and (layer5_outputs(4513));
    layer6_outputs(7627) <= not((layer5_outputs(1693)) or (layer5_outputs(3471)));
    layer6_outputs(7628) <= not(layer5_outputs(6802));
    layer6_outputs(7629) <= (layer5_outputs(4522)) xor (layer5_outputs(5895));
    layer6_outputs(7630) <= not(layer5_outputs(5945));
    layer6_outputs(7631) <= layer5_outputs(2776);
    layer6_outputs(7632) <= (layer5_outputs(6305)) and (layer5_outputs(3017));
    layer6_outputs(7633) <= not(layer5_outputs(7161));
    layer6_outputs(7634) <= not(layer5_outputs(759));
    layer6_outputs(7635) <= not((layer5_outputs(7116)) and (layer5_outputs(6713)));
    layer6_outputs(7636) <= (layer5_outputs(6544)) xor (layer5_outputs(4193));
    layer6_outputs(7637) <= layer5_outputs(3798);
    layer6_outputs(7638) <= layer5_outputs(5463);
    layer6_outputs(7639) <= layer5_outputs(1417);
    layer6_outputs(7640) <= not((layer5_outputs(6025)) xor (layer5_outputs(4291)));
    layer6_outputs(7641) <= not((layer5_outputs(6)) xor (layer5_outputs(4146)));
    layer6_outputs(7642) <= '1';
    layer6_outputs(7643) <= (layer5_outputs(6810)) and not (layer5_outputs(992));
    layer6_outputs(7644) <= (layer5_outputs(2882)) and not (layer5_outputs(4922));
    layer6_outputs(7645) <= layer5_outputs(4389);
    layer6_outputs(7646) <= not(layer5_outputs(6465)) or (layer5_outputs(1689));
    layer6_outputs(7647) <= not(layer5_outputs(3586));
    layer6_outputs(7648) <= not(layer5_outputs(80));
    layer6_outputs(7649) <= layer5_outputs(3647);
    layer6_outputs(7650) <= not((layer5_outputs(3684)) or (layer5_outputs(502)));
    layer6_outputs(7651) <= (layer5_outputs(1844)) or (layer5_outputs(7261));
    layer6_outputs(7652) <= layer5_outputs(6531);
    layer6_outputs(7653) <= layer5_outputs(5991);
    layer6_outputs(7654) <= layer5_outputs(6497);
    layer6_outputs(7655) <= not(layer5_outputs(5773));
    layer6_outputs(7656) <= layer5_outputs(1049);
    layer6_outputs(7657) <= not((layer5_outputs(5110)) xor (layer5_outputs(682)));
    layer6_outputs(7658) <= layer5_outputs(5376);
    layer6_outputs(7659) <= layer5_outputs(3172);
    layer6_outputs(7660) <= not(layer5_outputs(2717));
    layer6_outputs(7661) <= not(layer5_outputs(6081));
    layer6_outputs(7662) <= not(layer5_outputs(6519));
    layer6_outputs(7663) <= not((layer5_outputs(186)) xor (layer5_outputs(6344)));
    layer6_outputs(7664) <= not((layer5_outputs(1281)) xor (layer5_outputs(5944)));
    layer6_outputs(7665) <= not((layer5_outputs(5294)) or (layer5_outputs(2464)));
    layer6_outputs(7666) <= layer5_outputs(4400);
    layer6_outputs(7667) <= layer5_outputs(6107);
    layer6_outputs(7668) <= not((layer5_outputs(1304)) xor (layer5_outputs(7590)));
    layer6_outputs(7669) <= layer5_outputs(4280);
    layer6_outputs(7670) <= layer5_outputs(3037);
    layer6_outputs(7671) <= (layer5_outputs(1032)) xor (layer5_outputs(2603));
    layer6_outputs(7672) <= not(layer5_outputs(3519)) or (layer5_outputs(2936));
    layer6_outputs(7673) <= not(layer5_outputs(4051)) or (layer5_outputs(1649));
    layer6_outputs(7674) <= layer5_outputs(499);
    layer6_outputs(7675) <= layer5_outputs(5162);
    layer6_outputs(7676) <= not(layer5_outputs(6778));
    layer6_outputs(7677) <= not(layer5_outputs(5118));
    layer6_outputs(7678) <= layer5_outputs(1746);
    layer6_outputs(7679) <= layer5_outputs(2382);
    outputs(0) <= (layer6_outputs(138)) xor (layer6_outputs(2667));
    outputs(1) <= (layer6_outputs(1796)) xor (layer6_outputs(6650));
    outputs(2) <= not(layer6_outputs(6058));
    outputs(3) <= (layer6_outputs(1604)) and not (layer6_outputs(5533));
    outputs(4) <= not((layer6_outputs(5165)) or (layer6_outputs(4935)));
    outputs(5) <= not(layer6_outputs(1543));
    outputs(6) <= not((layer6_outputs(3676)) xor (layer6_outputs(3250)));
    outputs(7) <= layer6_outputs(1454);
    outputs(8) <= layer6_outputs(309);
    outputs(9) <= layer6_outputs(684);
    outputs(10) <= (layer6_outputs(6978)) xor (layer6_outputs(1672));
    outputs(11) <= not(layer6_outputs(995));
    outputs(12) <= not(layer6_outputs(1222));
    outputs(13) <= layer6_outputs(1818);
    outputs(14) <= not(layer6_outputs(2685));
    outputs(15) <= (layer6_outputs(7388)) xor (layer6_outputs(1488));
    outputs(16) <= layer6_outputs(4171);
    outputs(17) <= layer6_outputs(1621);
    outputs(18) <= not(layer6_outputs(1950));
    outputs(19) <= layer6_outputs(7352);
    outputs(20) <= (layer6_outputs(6287)) xor (layer6_outputs(6143));
    outputs(21) <= not(layer6_outputs(4334));
    outputs(22) <= not((layer6_outputs(1918)) xor (layer6_outputs(4008)));
    outputs(23) <= not(layer6_outputs(7232)) or (layer6_outputs(2533));
    outputs(24) <= not(layer6_outputs(3321));
    outputs(25) <= layer6_outputs(5316);
    outputs(26) <= not((layer6_outputs(3691)) xor (layer6_outputs(1843)));
    outputs(27) <= not(layer6_outputs(7518));
    outputs(28) <= not((layer6_outputs(544)) xor (layer6_outputs(4087)));
    outputs(29) <= (layer6_outputs(1688)) and not (layer6_outputs(6620));
    outputs(30) <= (layer6_outputs(4311)) xor (layer6_outputs(22));
    outputs(31) <= (layer6_outputs(3422)) and (layer6_outputs(3406));
    outputs(32) <= layer6_outputs(445);
    outputs(33) <= layer6_outputs(375);
    outputs(34) <= layer6_outputs(6773);
    outputs(35) <= not(layer6_outputs(5815));
    outputs(36) <= not(layer6_outputs(4172)) or (layer6_outputs(7540));
    outputs(37) <= (layer6_outputs(3731)) and (layer6_outputs(4275));
    outputs(38) <= not(layer6_outputs(7291));
    outputs(39) <= not(layer6_outputs(26));
    outputs(40) <= layer6_outputs(6152);
    outputs(41) <= layer6_outputs(1276);
    outputs(42) <= not(layer6_outputs(2222));
    outputs(43) <= not((layer6_outputs(1947)) xor (layer6_outputs(6924)));
    outputs(44) <= not((layer6_outputs(6748)) xor (layer6_outputs(919)));
    outputs(45) <= not(layer6_outputs(441));
    outputs(46) <= (layer6_outputs(4247)) xor (layer6_outputs(601));
    outputs(47) <= not((layer6_outputs(2906)) xor (layer6_outputs(3847)));
    outputs(48) <= layer6_outputs(4286);
    outputs(49) <= layer6_outputs(2422);
    outputs(50) <= not(layer6_outputs(5998));
    outputs(51) <= layer6_outputs(5850);
    outputs(52) <= not(layer6_outputs(1094));
    outputs(53) <= not((layer6_outputs(6189)) xor (layer6_outputs(4897)));
    outputs(54) <= layer6_outputs(2104);
    outputs(55) <= layer6_outputs(1741);
    outputs(56) <= not(layer6_outputs(3592)) or (layer6_outputs(2189));
    outputs(57) <= not(layer6_outputs(702));
    outputs(58) <= layer6_outputs(35);
    outputs(59) <= layer6_outputs(1402);
    outputs(60) <= layer6_outputs(6388);
    outputs(61) <= not(layer6_outputs(5490));
    outputs(62) <= not(layer6_outputs(5841));
    outputs(63) <= not(layer6_outputs(7019));
    outputs(64) <= (layer6_outputs(5764)) and not (layer6_outputs(878));
    outputs(65) <= not(layer6_outputs(3805));
    outputs(66) <= layer6_outputs(4772);
    outputs(67) <= layer6_outputs(2058);
    outputs(68) <= not(layer6_outputs(1230));
    outputs(69) <= layer6_outputs(7378);
    outputs(70) <= not((layer6_outputs(5617)) xor (layer6_outputs(5156)));
    outputs(71) <= not(layer6_outputs(954));
    outputs(72) <= not(layer6_outputs(6629));
    outputs(73) <= (layer6_outputs(9)) or (layer6_outputs(1684));
    outputs(74) <= not(layer6_outputs(51));
    outputs(75) <= not((layer6_outputs(3336)) or (layer6_outputs(936)));
    outputs(76) <= not(layer6_outputs(6281));
    outputs(77) <= not(layer6_outputs(1350));
    outputs(78) <= not(layer6_outputs(4260));
    outputs(79) <= (layer6_outputs(6958)) xor (layer6_outputs(6506));
    outputs(80) <= layer6_outputs(5908);
    outputs(81) <= not((layer6_outputs(6995)) or (layer6_outputs(7564)));
    outputs(82) <= not(layer6_outputs(696));
    outputs(83) <= (layer6_outputs(2532)) xor (layer6_outputs(7185));
    outputs(84) <= layer6_outputs(3911);
    outputs(85) <= layer6_outputs(770);
    outputs(86) <= not(layer6_outputs(3108));
    outputs(87) <= not(layer6_outputs(6001));
    outputs(88) <= layer6_outputs(7073);
    outputs(89) <= not(layer6_outputs(686));
    outputs(90) <= layer6_outputs(3756);
    outputs(91) <= layer6_outputs(4552);
    outputs(92) <= (layer6_outputs(4362)) xor (layer6_outputs(3865));
    outputs(93) <= layer6_outputs(5113);
    outputs(94) <= not(layer6_outputs(75));
    outputs(95) <= not(layer6_outputs(480));
    outputs(96) <= not(layer6_outputs(3745));
    outputs(97) <= not((layer6_outputs(2268)) or (layer6_outputs(4464)));
    outputs(98) <= not(layer6_outputs(7472));
    outputs(99) <= not(layer6_outputs(6931));
    outputs(100) <= layer6_outputs(1140);
    outputs(101) <= not(layer6_outputs(2202));
    outputs(102) <= not(layer6_outputs(5384));
    outputs(103) <= (layer6_outputs(6508)) and not (layer6_outputs(1238));
    outputs(104) <= layer6_outputs(2214);
    outputs(105) <= (layer6_outputs(2627)) xor (layer6_outputs(2254));
    outputs(106) <= (layer6_outputs(2079)) or (layer6_outputs(7627));
    outputs(107) <= not(layer6_outputs(7272));
    outputs(108) <= layer6_outputs(5318);
    outputs(109) <= (layer6_outputs(1075)) xor (layer6_outputs(7109));
    outputs(110) <= not(layer6_outputs(7009));
    outputs(111) <= not((layer6_outputs(2232)) xor (layer6_outputs(1609)));
    outputs(112) <= not(layer6_outputs(1555));
    outputs(113) <= (layer6_outputs(6394)) xor (layer6_outputs(444));
    outputs(114) <= not((layer6_outputs(1540)) xor (layer6_outputs(5303)));
    outputs(115) <= not(layer6_outputs(67));
    outputs(116) <= layer6_outputs(5297);
    outputs(117) <= not((layer6_outputs(4744)) or (layer6_outputs(1128)));
    outputs(118) <= not((layer6_outputs(2640)) xor (layer6_outputs(3790)));
    outputs(119) <= layer6_outputs(1749);
    outputs(120) <= layer6_outputs(1248);
    outputs(121) <= not(layer6_outputs(6250));
    outputs(122) <= layer6_outputs(5854);
    outputs(123) <= (layer6_outputs(3446)) and not (layer6_outputs(4075));
    outputs(124) <= (layer6_outputs(6176)) xor (layer6_outputs(7526));
    outputs(125) <= not(layer6_outputs(4059));
    outputs(126) <= layer6_outputs(3944);
    outputs(127) <= (layer6_outputs(5536)) and not (layer6_outputs(3459));
    outputs(128) <= not((layer6_outputs(367)) and (layer6_outputs(1703)));
    outputs(129) <= not(layer6_outputs(1956));
    outputs(130) <= layer6_outputs(7458);
    outputs(131) <= (layer6_outputs(6891)) and not (layer6_outputs(5012));
    outputs(132) <= layer6_outputs(1890);
    outputs(133) <= layer6_outputs(1107);
    outputs(134) <= not((layer6_outputs(1197)) xor (layer6_outputs(4163)));
    outputs(135) <= (layer6_outputs(7121)) and (layer6_outputs(6041));
    outputs(136) <= not((layer6_outputs(65)) xor (layer6_outputs(7245)));
    outputs(137) <= layer6_outputs(2701);
    outputs(138) <= (layer6_outputs(2052)) xor (layer6_outputs(7565));
    outputs(139) <= (layer6_outputs(394)) xor (layer6_outputs(1216));
    outputs(140) <= layer6_outputs(432);
    outputs(141) <= not(layer6_outputs(5048));
    outputs(142) <= not(layer6_outputs(1968));
    outputs(143) <= not((layer6_outputs(1268)) xor (layer6_outputs(7308)));
    outputs(144) <= (layer6_outputs(1716)) xor (layer6_outputs(1071));
    outputs(145) <= not(layer6_outputs(1880));
    outputs(146) <= layer6_outputs(1759);
    outputs(147) <= layer6_outputs(2164);
    outputs(148) <= not((layer6_outputs(1364)) xor (layer6_outputs(3393)));
    outputs(149) <= not((layer6_outputs(3494)) xor (layer6_outputs(1574)));
    outputs(150) <= layer6_outputs(5199);
    outputs(151) <= (layer6_outputs(1591)) xor (layer6_outputs(4311));
    outputs(152) <= not(layer6_outputs(4205));
    outputs(153) <= layer6_outputs(945);
    outputs(154) <= not(layer6_outputs(2091));
    outputs(155) <= layer6_outputs(5892);
    outputs(156) <= (layer6_outputs(3518)) and (layer6_outputs(3348));
    outputs(157) <= layer6_outputs(7140);
    outputs(158) <= (layer6_outputs(6743)) and (layer6_outputs(648));
    outputs(159) <= layer6_outputs(7214);
    outputs(160) <= not(layer6_outputs(4283));
    outputs(161) <= not(layer6_outputs(5933));
    outputs(162) <= layer6_outputs(4655);
    outputs(163) <= not((layer6_outputs(3158)) xor (layer6_outputs(2542)));
    outputs(164) <= not((layer6_outputs(6669)) xor (layer6_outputs(7123)));
    outputs(165) <= layer6_outputs(4929);
    outputs(166) <= not(layer6_outputs(1120)) or (layer6_outputs(5748));
    outputs(167) <= not(layer6_outputs(482));
    outputs(168) <= (layer6_outputs(6630)) xor (layer6_outputs(7543));
    outputs(169) <= layer6_outputs(534);
    outputs(170) <= not(layer6_outputs(4130));
    outputs(171) <= not(layer6_outputs(4182));
    outputs(172) <= not(layer6_outputs(3775));
    outputs(173) <= (layer6_outputs(2043)) and not (layer6_outputs(4526));
    outputs(174) <= layer6_outputs(6337);
    outputs(175) <= (layer6_outputs(4553)) xor (layer6_outputs(1747));
    outputs(176) <= not(layer6_outputs(7592));
    outputs(177) <= not(layer6_outputs(6939));
    outputs(178) <= not(layer6_outputs(5052));
    outputs(179) <= not(layer6_outputs(710));
    outputs(180) <= layer6_outputs(1225);
    outputs(181) <= (layer6_outputs(2165)) and (layer6_outputs(6895));
    outputs(182) <= not((layer6_outputs(3605)) and (layer6_outputs(3553)));
    outputs(183) <= not((layer6_outputs(5010)) or (layer6_outputs(3768)));
    outputs(184) <= (layer6_outputs(5372)) and not (layer6_outputs(2094));
    outputs(185) <= not((layer6_outputs(1547)) xor (layer6_outputs(5929)));
    outputs(186) <= layer6_outputs(4956);
    outputs(187) <= (layer6_outputs(1353)) and (layer6_outputs(2136));
    outputs(188) <= not((layer6_outputs(1187)) xor (layer6_outputs(1715)));
    outputs(189) <= layer6_outputs(6374);
    outputs(190) <= not((layer6_outputs(5149)) or (layer6_outputs(3962)));
    outputs(191) <= layer6_outputs(223);
    outputs(192) <= (layer6_outputs(3460)) xor (layer6_outputs(2021));
    outputs(193) <= (layer6_outputs(866)) xor (layer6_outputs(1584));
    outputs(194) <= not((layer6_outputs(4752)) or (layer6_outputs(1210)));
    outputs(195) <= not((layer6_outputs(3630)) or (layer6_outputs(2140)));
    outputs(196) <= (layer6_outputs(6112)) and not (layer6_outputs(1921));
    outputs(197) <= (layer6_outputs(5762)) or (layer6_outputs(6785));
    outputs(198) <= layer6_outputs(7157);
    outputs(199) <= not(layer6_outputs(2907));
    outputs(200) <= not((layer6_outputs(6771)) xor (layer6_outputs(3207)));
    outputs(201) <= not(layer6_outputs(5905));
    outputs(202) <= not(layer6_outputs(7097));
    outputs(203) <= not(layer6_outputs(6086));
    outputs(204) <= layer6_outputs(3280);
    outputs(205) <= layer6_outputs(188);
    outputs(206) <= not(layer6_outputs(2512));
    outputs(207) <= (layer6_outputs(722)) xor (layer6_outputs(2997));
    outputs(208) <= not(layer6_outputs(1525));
    outputs(209) <= not(layer6_outputs(325));
    outputs(210) <= layer6_outputs(6642);
    outputs(211) <= layer6_outputs(5564);
    outputs(212) <= (layer6_outputs(5299)) xor (layer6_outputs(5308));
    outputs(213) <= not(layer6_outputs(1649));
    outputs(214) <= not(layer6_outputs(694));
    outputs(215) <= not((layer6_outputs(6660)) xor (layer6_outputs(5123)));
    outputs(216) <= (layer6_outputs(5562)) and (layer6_outputs(2781));
    outputs(217) <= layer6_outputs(913);
    outputs(218) <= layer6_outputs(198);
    outputs(219) <= layer6_outputs(3315);
    outputs(220) <= not(layer6_outputs(7279));
    outputs(221) <= not(layer6_outputs(5818));
    outputs(222) <= layer6_outputs(5147);
    outputs(223) <= not(layer6_outputs(6180));
    outputs(224) <= layer6_outputs(2394);
    outputs(225) <= not(layer6_outputs(6565));
    outputs(226) <= not(layer6_outputs(1407)) or (layer6_outputs(3916));
    outputs(227) <= not(layer6_outputs(7489));
    outputs(228) <= (layer6_outputs(2035)) xor (layer6_outputs(6869));
    outputs(229) <= not(layer6_outputs(4589));
    outputs(230) <= layer6_outputs(6324);
    outputs(231) <= not(layer6_outputs(4834));
    outputs(232) <= not((layer6_outputs(2788)) xor (layer6_outputs(1186)));
    outputs(233) <= (layer6_outputs(2451)) and not (layer6_outputs(5751));
    outputs(234) <= (layer6_outputs(7110)) xor (layer6_outputs(2228));
    outputs(235) <= (layer6_outputs(6185)) or (layer6_outputs(7192));
    outputs(236) <= not((layer6_outputs(5494)) or (layer6_outputs(5607)));
    outputs(237) <= not(layer6_outputs(7115));
    outputs(238) <= layer6_outputs(7475);
    outputs(239) <= layer6_outputs(2785);
    outputs(240) <= layer6_outputs(605);
    outputs(241) <= (layer6_outputs(1281)) xor (layer6_outputs(7130));
    outputs(242) <= not((layer6_outputs(7005)) or (layer6_outputs(788)));
    outputs(243) <= not(layer6_outputs(4542));
    outputs(244) <= layer6_outputs(770);
    outputs(245) <= not(layer6_outputs(2780));
    outputs(246) <= not(layer6_outputs(4775));
    outputs(247) <= layer6_outputs(3182);
    outputs(248) <= not(layer6_outputs(541));
    outputs(249) <= not(layer6_outputs(6406));
    outputs(250) <= not(layer6_outputs(655));
    outputs(251) <= (layer6_outputs(1599)) xor (layer6_outputs(4204));
    outputs(252) <= not(layer6_outputs(5665));
    outputs(253) <= (layer6_outputs(666)) xor (layer6_outputs(5187));
    outputs(254) <= not(layer6_outputs(3587));
    outputs(255) <= not(layer6_outputs(5015));
    outputs(256) <= (layer6_outputs(2341)) and not (layer6_outputs(1294));
    outputs(257) <= layer6_outputs(6061);
    outputs(258) <= (layer6_outputs(6135)) xor (layer6_outputs(1071));
    outputs(259) <= not(layer6_outputs(4682));
    outputs(260) <= layer6_outputs(5790);
    outputs(261) <= layer6_outputs(7392);
    outputs(262) <= not(layer6_outputs(1776));
    outputs(263) <= not(layer6_outputs(4140));
    outputs(264) <= not(layer6_outputs(783));
    outputs(265) <= not(layer6_outputs(2860));
    outputs(266) <= layer6_outputs(5526);
    outputs(267) <= not(layer6_outputs(7346));
    outputs(268) <= layer6_outputs(4447);
    outputs(269) <= (layer6_outputs(7340)) xor (layer6_outputs(2587));
    outputs(270) <= not(layer6_outputs(2145));
    outputs(271) <= not(layer6_outputs(3412)) or (layer6_outputs(6817));
    outputs(272) <= not(layer6_outputs(747));
    outputs(273) <= not((layer6_outputs(2253)) xor (layer6_outputs(6496)));
    outputs(274) <= not((layer6_outputs(5043)) xor (layer6_outputs(2256)));
    outputs(275) <= (layer6_outputs(1215)) xor (layer6_outputs(7601));
    outputs(276) <= layer6_outputs(2593);
    outputs(277) <= not(layer6_outputs(1025));
    outputs(278) <= not(layer6_outputs(4194));
    outputs(279) <= (layer6_outputs(2178)) xor (layer6_outputs(4290));
    outputs(280) <= not(layer6_outputs(827));
    outputs(281) <= not(layer6_outputs(411));
    outputs(282) <= not(layer6_outputs(2501));
    outputs(283) <= layer6_outputs(5638);
    outputs(284) <= (layer6_outputs(2609)) xor (layer6_outputs(6552));
    outputs(285) <= not((layer6_outputs(1133)) xor (layer6_outputs(844)));
    outputs(286) <= not((layer6_outputs(4659)) and (layer6_outputs(421)));
    outputs(287) <= not((layer6_outputs(6104)) xor (layer6_outputs(7353)));
    outputs(288) <= layer6_outputs(2205);
    outputs(289) <= layer6_outputs(321);
    outputs(290) <= not(layer6_outputs(5466));
    outputs(291) <= not((layer6_outputs(3099)) or (layer6_outputs(6789)));
    outputs(292) <= not(layer6_outputs(2715));
    outputs(293) <= not((layer6_outputs(5300)) or (layer6_outputs(4904)));
    outputs(294) <= layer6_outputs(490);
    outputs(295) <= not((layer6_outputs(5174)) xor (layer6_outputs(2422)));
    outputs(296) <= not((layer6_outputs(7105)) xor (layer6_outputs(5636)));
    outputs(297) <= not(layer6_outputs(7084));
    outputs(298) <= (layer6_outputs(7485)) and not (layer6_outputs(2117));
    outputs(299) <= not(layer6_outputs(2354));
    outputs(300) <= not(layer6_outputs(6662));
    outputs(301) <= layer6_outputs(1362);
    outputs(302) <= (layer6_outputs(4351)) xor (layer6_outputs(4199));
    outputs(303) <= not(layer6_outputs(3265));
    outputs(304) <= not(layer6_outputs(4608)) or (layer6_outputs(7339));
    outputs(305) <= layer6_outputs(3190);
    outputs(306) <= (layer6_outputs(2380)) and not (layer6_outputs(2286));
    outputs(307) <= not((layer6_outputs(5504)) and (layer6_outputs(1607)));
    outputs(308) <= not(layer6_outputs(7638));
    outputs(309) <= not((layer6_outputs(773)) xor (layer6_outputs(7438)));
    outputs(310) <= (layer6_outputs(6802)) xor (layer6_outputs(4936));
    outputs(311) <= layer6_outputs(349);
    outputs(312) <= (layer6_outputs(6377)) and not (layer6_outputs(4409));
    outputs(313) <= not(layer6_outputs(4791));
    outputs(314) <= not((layer6_outputs(1048)) xor (layer6_outputs(589)));
    outputs(315) <= layer6_outputs(1357);
    outputs(316) <= not((layer6_outputs(4421)) and (layer6_outputs(5246)));
    outputs(317) <= not(layer6_outputs(6310)) or (layer6_outputs(4757));
    outputs(318) <= not(layer6_outputs(2386));
    outputs(319) <= layer6_outputs(3740);
    outputs(320) <= (layer6_outputs(6477)) xor (layer6_outputs(7195));
    outputs(321) <= not(layer6_outputs(103));
    outputs(322) <= not(layer6_outputs(5615)) or (layer6_outputs(4949));
    outputs(323) <= not((layer6_outputs(7651)) xor (layer6_outputs(1568)));
    outputs(324) <= not(layer6_outputs(4093));
    outputs(325) <= not(layer6_outputs(190)) or (layer6_outputs(7602));
    outputs(326) <= (layer6_outputs(4971)) xor (layer6_outputs(1209));
    outputs(327) <= layer6_outputs(7331);
    outputs(328) <= not(layer6_outputs(4539));
    outputs(329) <= not(layer6_outputs(1636));
    outputs(330) <= layer6_outputs(817);
    outputs(331) <= not((layer6_outputs(5420)) xor (layer6_outputs(340)));
    outputs(332) <= layer6_outputs(365);
    outputs(333) <= not((layer6_outputs(4570)) xor (layer6_outputs(6763)));
    outputs(334) <= not((layer6_outputs(2920)) xor (layer6_outputs(4735)));
    outputs(335) <= layer6_outputs(5649);
    outputs(336) <= not(layer6_outputs(3991));
    outputs(337) <= not((layer6_outputs(5802)) xor (layer6_outputs(2999)));
    outputs(338) <= not((layer6_outputs(2146)) xor (layer6_outputs(1566)));
    outputs(339) <= layer6_outputs(1163);
    outputs(340) <= not((layer6_outputs(3803)) xor (layer6_outputs(1506)));
    outputs(341) <= (layer6_outputs(6168)) xor (layer6_outputs(2629));
    outputs(342) <= not(layer6_outputs(7280));
    outputs(343) <= layer6_outputs(6472);
    outputs(344) <= layer6_outputs(1677);
    outputs(345) <= layer6_outputs(7523);
    outputs(346) <= (layer6_outputs(43)) xor (layer6_outputs(3647));
    outputs(347) <= layer6_outputs(549);
    outputs(348) <= layer6_outputs(417);
    outputs(349) <= not(layer6_outputs(7267));
    outputs(350) <= not((layer6_outputs(4429)) xor (layer6_outputs(5997)));
    outputs(351) <= not(layer6_outputs(5446));
    outputs(352) <= (layer6_outputs(3897)) and (layer6_outputs(1466));
    outputs(353) <= (layer6_outputs(2580)) xor (layer6_outputs(3712));
    outputs(354) <= not(layer6_outputs(1224));
    outputs(355) <= not(layer6_outputs(1889)) or (layer6_outputs(474));
    outputs(356) <= (layer6_outputs(4747)) and not (layer6_outputs(6330));
    outputs(357) <= not((layer6_outputs(5013)) xor (layer6_outputs(427)));
    outputs(358) <= layer6_outputs(3363);
    outputs(359) <= not((layer6_outputs(4192)) xor (layer6_outputs(5519)));
    outputs(360) <= layer6_outputs(3307);
    outputs(361) <= not(layer6_outputs(998)) or (layer6_outputs(7416));
    outputs(362) <= not(layer6_outputs(6483));
    outputs(363) <= not(layer6_outputs(2129));
    outputs(364) <= not(layer6_outputs(4963));
    outputs(365) <= (layer6_outputs(7234)) xor (layer6_outputs(1013));
    outputs(366) <= layer6_outputs(5361);
    outputs(367) <= not(layer6_outputs(1758));
    outputs(368) <= not(layer6_outputs(2209));
    outputs(369) <= (layer6_outputs(4776)) xor (layer6_outputs(1608));
    outputs(370) <= not(layer6_outputs(6260)) or (layer6_outputs(1021));
    outputs(371) <= (layer6_outputs(1242)) and not (layer6_outputs(302));
    outputs(372) <= not((layer6_outputs(6263)) xor (layer6_outputs(2905)));
    outputs(373) <= layer6_outputs(4653);
    outputs(374) <= layer6_outputs(3152);
    outputs(375) <= layer6_outputs(1526);
    outputs(376) <= not(layer6_outputs(5106)) or (layer6_outputs(3274));
    outputs(377) <= not(layer6_outputs(3413));
    outputs(378) <= (layer6_outputs(2245)) xor (layer6_outputs(1396));
    outputs(379) <= not(layer6_outputs(6154));
    outputs(380) <= not(layer6_outputs(1801));
    outputs(381) <= (layer6_outputs(3444)) xor (layer6_outputs(2240));
    outputs(382) <= layer6_outputs(1872);
    outputs(383) <= not((layer6_outputs(946)) and (layer6_outputs(898)));
    outputs(384) <= layer6_outputs(3407);
    outputs(385) <= (layer6_outputs(4556)) xor (layer6_outputs(5054));
    outputs(386) <= not(layer6_outputs(5766));
    outputs(387) <= not(layer6_outputs(3535));
    outputs(388) <= layer6_outputs(3199);
    outputs(389) <= (layer6_outputs(4704)) and (layer6_outputs(885));
    outputs(390) <= (layer6_outputs(4686)) and not (layer6_outputs(6762));
    outputs(391) <= layer6_outputs(4854);
    outputs(392) <= not(layer6_outputs(2018));
    outputs(393) <= layer6_outputs(678);
    outputs(394) <= (layer6_outputs(4416)) xor (layer6_outputs(259));
    outputs(395) <= not((layer6_outputs(2245)) xor (layer6_outputs(694)));
    outputs(396) <= not((layer6_outputs(178)) xor (layer6_outputs(6836)));
    outputs(397) <= (layer6_outputs(6039)) and (layer6_outputs(6843));
    outputs(398) <= layer6_outputs(6890);
    outputs(399) <= layer6_outputs(3469);
    outputs(400) <= layer6_outputs(7138);
    outputs(401) <= not(layer6_outputs(5941));
    outputs(402) <= (layer6_outputs(627)) xor (layer6_outputs(7162));
    outputs(403) <= layer6_outputs(6277);
    outputs(404) <= (layer6_outputs(2221)) and not (layer6_outputs(3024));
    outputs(405) <= (layer6_outputs(5061)) xor (layer6_outputs(52));
    outputs(406) <= not((layer6_outputs(1708)) and (layer6_outputs(1665)));
    outputs(407) <= not((layer6_outputs(486)) or (layer6_outputs(5722)));
    outputs(408) <= not((layer6_outputs(6077)) xor (layer6_outputs(1800)));
    outputs(409) <= not(layer6_outputs(4605));
    outputs(410) <= not((layer6_outputs(1326)) xor (layer6_outputs(2712)));
    outputs(411) <= not(layer6_outputs(1520));
    outputs(412) <= (layer6_outputs(5849)) xor (layer6_outputs(2225));
    outputs(413) <= layer6_outputs(6850);
    outputs(414) <= not(layer6_outputs(1914));
    outputs(415) <= not((layer6_outputs(3537)) xor (layer6_outputs(6982)));
    outputs(416) <= not(layer6_outputs(4098));
    outputs(417) <= not((layer6_outputs(4010)) and (layer6_outputs(6341)));
    outputs(418) <= (layer6_outputs(6580)) xor (layer6_outputs(5806));
    outputs(419) <= not(layer6_outputs(2097));
    outputs(420) <= layer6_outputs(3429);
    outputs(421) <= not((layer6_outputs(6820)) xor (layer6_outputs(7348)));
    outputs(422) <= not(layer6_outputs(1082));
    outputs(423) <= not((layer6_outputs(4577)) xor (layer6_outputs(1926)));
    outputs(424) <= layer6_outputs(3771);
    outputs(425) <= not((layer6_outputs(2665)) or (layer6_outputs(6869)));
    outputs(426) <= not((layer6_outputs(1961)) xor (layer6_outputs(7678)));
    outputs(427) <= not(layer6_outputs(3752));
    outputs(428) <= not(layer6_outputs(1806));
    outputs(429) <= (layer6_outputs(1680)) and (layer6_outputs(5111));
    outputs(430) <= not(layer6_outputs(74));
    outputs(431) <= (layer6_outputs(1080)) xor (layer6_outputs(2436));
    outputs(432) <= not((layer6_outputs(6188)) or (layer6_outputs(5499)));
    outputs(433) <= (layer6_outputs(6861)) and (layer6_outputs(1038));
    outputs(434) <= not(layer6_outputs(98)) or (layer6_outputs(28));
    outputs(435) <= layer6_outputs(3128);
    outputs(436) <= not(layer6_outputs(5594));
    outputs(437) <= not((layer6_outputs(2375)) xor (layer6_outputs(3337)));
    outputs(438) <= layer6_outputs(1461);
    outputs(439) <= not(layer6_outputs(4098));
    outputs(440) <= not((layer6_outputs(5956)) xor (layer6_outputs(6705)));
    outputs(441) <= not(layer6_outputs(758));
    outputs(442) <= not(layer6_outputs(7063));
    outputs(443) <= layer6_outputs(3748);
    outputs(444) <= not(layer6_outputs(5417));
    outputs(445) <= layer6_outputs(5563);
    outputs(446) <= layer6_outputs(526);
    outputs(447) <= (layer6_outputs(4214)) xor (layer6_outputs(61));
    outputs(448) <= not(layer6_outputs(3624));
    outputs(449) <= layer6_outputs(3573);
    outputs(450) <= not(layer6_outputs(1837));
    outputs(451) <= not(layer6_outputs(6349));
    outputs(452) <= not(layer6_outputs(2351));
    outputs(453) <= (layer6_outputs(3020)) or (layer6_outputs(1549));
    outputs(454) <= (layer6_outputs(1353)) and (layer6_outputs(1809));
    outputs(455) <= layer6_outputs(2980);
    outputs(456) <= not((layer6_outputs(7347)) xor (layer6_outputs(6899)));
    outputs(457) <= (layer6_outputs(50)) xor (layer6_outputs(6396));
    outputs(458) <= (layer6_outputs(6092)) and not (layer6_outputs(5182));
    outputs(459) <= (layer6_outputs(3137)) xor (layer6_outputs(2452));
    outputs(460) <= not(layer6_outputs(4049));
    outputs(461) <= not(layer6_outputs(6448));
    outputs(462) <= not((layer6_outputs(7441)) xor (layer6_outputs(4350)));
    outputs(463) <= (layer6_outputs(1665)) xor (layer6_outputs(4797));
    outputs(464) <= layer6_outputs(3601);
    outputs(465) <= not(layer6_outputs(632));
    outputs(466) <= layer6_outputs(3058);
    outputs(467) <= layer6_outputs(808);
    outputs(468) <= not((layer6_outputs(3610)) xor (layer6_outputs(454)));
    outputs(469) <= not(layer6_outputs(2559)) or (layer6_outputs(3717));
    outputs(470) <= not(layer6_outputs(2802));
    outputs(471) <= (layer6_outputs(2322)) xor (layer6_outputs(6265));
    outputs(472) <= not(layer6_outputs(3762));
    outputs(473) <= layer6_outputs(6370);
    outputs(474) <= not(layer6_outputs(51));
    outputs(475) <= not((layer6_outputs(3514)) xor (layer6_outputs(2154)));
    outputs(476) <= not((layer6_outputs(7293)) xor (layer6_outputs(5474)));
    outputs(477) <= (layer6_outputs(203)) and not (layer6_outputs(6035));
    outputs(478) <= not((layer6_outputs(1083)) xor (layer6_outputs(6489)));
    outputs(479) <= '0';
    outputs(480) <= not(layer6_outputs(2478));
    outputs(481) <= not(layer6_outputs(4943));
    outputs(482) <= layer6_outputs(1446);
    outputs(483) <= not((layer6_outputs(1837)) xor (layer6_outputs(2806)));
    outputs(484) <= not(layer6_outputs(298));
    outputs(485) <= not(layer6_outputs(5052));
    outputs(486) <= (layer6_outputs(7226)) xor (layer6_outputs(2447));
    outputs(487) <= not(layer6_outputs(6084));
    outputs(488) <= not(layer6_outputs(7010));
    outputs(489) <= not(layer6_outputs(2923));
    outputs(490) <= (layer6_outputs(7402)) xor (layer6_outputs(1578));
    outputs(491) <= (layer6_outputs(2874)) xor (layer6_outputs(255));
    outputs(492) <= not(layer6_outputs(1223));
    outputs(493) <= layer6_outputs(287);
    outputs(494) <= not(layer6_outputs(201));
    outputs(495) <= layer6_outputs(6958);
    outputs(496) <= not(layer6_outputs(6966));
    outputs(497) <= (layer6_outputs(5451)) and not (layer6_outputs(5640));
    outputs(498) <= (layer6_outputs(489)) and not (layer6_outputs(314));
    outputs(499) <= not(layer6_outputs(1696));
    outputs(500) <= layer6_outputs(6703);
    outputs(501) <= layer6_outputs(6088);
    outputs(502) <= not(layer6_outputs(1814));
    outputs(503) <= layer6_outputs(4765);
    outputs(504) <= layer6_outputs(3430);
    outputs(505) <= (layer6_outputs(1572)) and (layer6_outputs(6544));
    outputs(506) <= (layer6_outputs(1902)) xor (layer6_outputs(6753));
    outputs(507) <= not(layer6_outputs(3326)) or (layer6_outputs(1));
    outputs(508) <= not(layer6_outputs(3292));
    outputs(509) <= (layer6_outputs(7480)) xor (layer6_outputs(2030));
    outputs(510) <= not(layer6_outputs(4911)) or (layer6_outputs(6989));
    outputs(511) <= not(layer6_outputs(5285));
    outputs(512) <= not(layer6_outputs(6249));
    outputs(513) <= not(layer6_outputs(5991));
    outputs(514) <= layer6_outputs(4615);
    outputs(515) <= (layer6_outputs(6661)) xor (layer6_outputs(2537));
    outputs(516) <= layer6_outputs(5385);
    outputs(517) <= not((layer6_outputs(5221)) xor (layer6_outputs(6171)));
    outputs(518) <= not(layer6_outputs(4000));
    outputs(519) <= not(layer6_outputs(4734));
    outputs(520) <= not(layer6_outputs(3535));
    outputs(521) <= (layer6_outputs(1887)) xor (layer6_outputs(3701));
    outputs(522) <= layer6_outputs(3903);
    outputs(523) <= not((layer6_outputs(1871)) xor (layer6_outputs(1285)));
    outputs(524) <= not((layer6_outputs(2978)) xor (layer6_outputs(6366)));
    outputs(525) <= not(layer6_outputs(120));
    outputs(526) <= layer6_outputs(5588);
    outputs(527) <= (layer6_outputs(6488)) xor (layer6_outputs(5657));
    outputs(528) <= not(layer6_outputs(5427));
    outputs(529) <= not(layer6_outputs(6042));
    outputs(530) <= not((layer6_outputs(6612)) xor (layer6_outputs(2743)));
    outputs(531) <= not(layer6_outputs(2159));
    outputs(532) <= (layer6_outputs(3502)) xor (layer6_outputs(4773));
    outputs(533) <= (layer6_outputs(6810)) xor (layer6_outputs(1085));
    outputs(534) <= layer6_outputs(672);
    outputs(535) <= layer6_outputs(3461);
    outputs(536) <= not(layer6_outputs(7085));
    outputs(537) <= not(layer6_outputs(3936));
    outputs(538) <= not(layer6_outputs(1656));
    outputs(539) <= not(layer6_outputs(7546));
    outputs(540) <= (layer6_outputs(5243)) and not (layer6_outputs(789));
    outputs(541) <= (layer6_outputs(765)) xor (layer6_outputs(2469));
    outputs(542) <= layer6_outputs(1771);
    outputs(543) <= not((layer6_outputs(6573)) xor (layer6_outputs(5458)));
    outputs(544) <= layer6_outputs(6631);
    outputs(545) <= not((layer6_outputs(2908)) xor (layer6_outputs(4593)));
    outputs(546) <= (layer6_outputs(905)) xor (layer6_outputs(6073));
    outputs(547) <= not((layer6_outputs(4544)) xor (layer6_outputs(965)));
    outputs(548) <= layer6_outputs(4272);
    outputs(549) <= (layer6_outputs(598)) xor (layer6_outputs(1412));
    outputs(550) <= layer6_outputs(3341);
    outputs(551) <= (layer6_outputs(282)) xor (layer6_outputs(2894));
    outputs(552) <= layer6_outputs(4976);
    outputs(553) <= not(layer6_outputs(4829));
    outputs(554) <= not((layer6_outputs(1732)) xor (layer6_outputs(7174)));
    outputs(555) <= not((layer6_outputs(7309)) xor (layer6_outputs(2978)));
    outputs(556) <= not((layer6_outputs(1064)) xor (layer6_outputs(3747)));
    outputs(557) <= not((layer6_outputs(6611)) or (layer6_outputs(2555)));
    outputs(558) <= not(layer6_outputs(7215));
    outputs(559) <= layer6_outputs(4181);
    outputs(560) <= not(layer6_outputs(6944));
    outputs(561) <= layer6_outputs(3585);
    outputs(562) <= not((layer6_outputs(5322)) xor (layer6_outputs(3538)));
    outputs(563) <= not(layer6_outputs(5060));
    outputs(564) <= layer6_outputs(7435);
    outputs(565) <= (layer6_outputs(7329)) xor (layer6_outputs(3321));
    outputs(566) <= not(layer6_outputs(2268));
    outputs(567) <= not(layer6_outputs(2783));
    outputs(568) <= (layer6_outputs(5394)) xor (layer6_outputs(7443));
    outputs(569) <= not((layer6_outputs(1842)) xor (layer6_outputs(1067)));
    outputs(570) <= (layer6_outputs(900)) xor (layer6_outputs(5180));
    outputs(571) <= (layer6_outputs(3033)) and not (layer6_outputs(1004));
    outputs(572) <= (layer6_outputs(1893)) xor (layer6_outputs(6257));
    outputs(573) <= not((layer6_outputs(593)) xor (layer6_outputs(4130)));
    outputs(574) <= not(layer6_outputs(2044));
    outputs(575) <= (layer6_outputs(4326)) xor (layer6_outputs(4414));
    outputs(576) <= not(layer6_outputs(7294)) or (layer6_outputs(662));
    outputs(577) <= (layer6_outputs(2331)) xor (layer6_outputs(6321));
    outputs(578) <= (layer6_outputs(683)) xor (layer6_outputs(6780));
    outputs(579) <= layer6_outputs(3039);
    outputs(580) <= (layer6_outputs(6607)) xor (layer6_outputs(3539));
    outputs(581) <= (layer6_outputs(2088)) xor (layer6_outputs(1136));
    outputs(582) <= layer6_outputs(2619);
    outputs(583) <= (layer6_outputs(439)) xor (layer6_outputs(6484));
    outputs(584) <= not((layer6_outputs(3974)) xor (layer6_outputs(1784)));
    outputs(585) <= layer6_outputs(6513);
    outputs(586) <= not((layer6_outputs(1299)) and (layer6_outputs(3203)));
    outputs(587) <= (layer6_outputs(5104)) and not (layer6_outputs(6564));
    outputs(588) <= layer6_outputs(6616);
    outputs(589) <= layer6_outputs(4313);
    outputs(590) <= layer6_outputs(1744);
    outputs(591) <= (layer6_outputs(7200)) xor (layer6_outputs(5047));
    outputs(592) <= (layer6_outputs(7480)) or (layer6_outputs(376));
    outputs(593) <= not((layer6_outputs(22)) and (layer6_outputs(7229)));
    outputs(594) <= not(layer6_outputs(3017));
    outputs(595) <= layer6_outputs(240);
    outputs(596) <= (layer6_outputs(7335)) xor (layer6_outputs(7661));
    outputs(597) <= not(layer6_outputs(428));
    outputs(598) <= not(layer6_outputs(4236));
    outputs(599) <= not((layer6_outputs(1252)) or (layer6_outputs(858)));
    outputs(600) <= not((layer6_outputs(4207)) xor (layer6_outputs(4022)));
    outputs(601) <= not(layer6_outputs(7323));
    outputs(602) <= (layer6_outputs(6893)) xor (layer6_outputs(2217));
    outputs(603) <= not((layer6_outputs(4518)) xor (layer6_outputs(384)));
    outputs(604) <= not(layer6_outputs(2500));
    outputs(605) <= layer6_outputs(5138);
    outputs(606) <= not(layer6_outputs(3864));
    outputs(607) <= not((layer6_outputs(7439)) xor (layer6_outputs(7462)));
    outputs(608) <= not(layer6_outputs(1220));
    outputs(609) <= not(layer6_outputs(5832)) or (layer6_outputs(4582));
    outputs(610) <= not((layer6_outputs(6678)) and (layer6_outputs(5174)));
    outputs(611) <= not(layer6_outputs(6711)) or (layer6_outputs(6251));
    outputs(612) <= (layer6_outputs(1684)) xor (layer6_outputs(2654));
    outputs(613) <= (layer6_outputs(6870)) and (layer6_outputs(1764));
    outputs(614) <= layer6_outputs(69);
    outputs(615) <= (layer6_outputs(5062)) xor (layer6_outputs(110));
    outputs(616) <= not((layer6_outputs(173)) xor (layer6_outputs(6003)));
    outputs(617) <= not(layer6_outputs(2631));
    outputs(618) <= not(layer6_outputs(2183));
    outputs(619) <= not(layer6_outputs(1752));
    outputs(620) <= layer6_outputs(6967);
    outputs(621) <= (layer6_outputs(5748)) or (layer6_outputs(3283));
    outputs(622) <= not((layer6_outputs(4905)) or (layer6_outputs(5121)));
    outputs(623) <= layer6_outputs(414);
    outputs(624) <= (layer6_outputs(161)) xor (layer6_outputs(674));
    outputs(625) <= not(layer6_outputs(2892));
    outputs(626) <= (layer6_outputs(6041)) xor (layer6_outputs(1173));
    outputs(627) <= (layer6_outputs(2267)) xor (layer6_outputs(1599));
    outputs(628) <= (layer6_outputs(4026)) or (layer6_outputs(2598));
    outputs(629) <= layer6_outputs(6610);
    outputs(630) <= layer6_outputs(5339);
    outputs(631) <= not(layer6_outputs(6020));
    outputs(632) <= layer6_outputs(1330);
    outputs(633) <= not((layer6_outputs(3497)) xor (layer6_outputs(1449)));
    outputs(634) <= not(layer6_outputs(2411));
    outputs(635) <= layer6_outputs(592);
    outputs(636) <= layer6_outputs(3868);
    outputs(637) <= layer6_outputs(4907);
    outputs(638) <= (layer6_outputs(1073)) and not (layer6_outputs(2636));
    outputs(639) <= (layer6_outputs(3213)) xor (layer6_outputs(7313));
    outputs(640) <= layer6_outputs(1870);
    outputs(641) <= (layer6_outputs(1239)) xor (layer6_outputs(3854));
    outputs(642) <= layer6_outputs(7474);
    outputs(643) <= not(layer6_outputs(3996));
    outputs(644) <= not((layer6_outputs(7523)) xor (layer6_outputs(6441)));
    outputs(645) <= layer6_outputs(990);
    outputs(646) <= layer6_outputs(2630);
    outputs(647) <= not((layer6_outputs(6186)) xor (layer6_outputs(7366)));
    outputs(648) <= not(layer6_outputs(2513));
    outputs(649) <= (layer6_outputs(4932)) and not (layer6_outputs(5095));
    outputs(650) <= not(layer6_outputs(5809));
    outputs(651) <= (layer6_outputs(5179)) xor (layer6_outputs(2787));
    outputs(652) <= layer6_outputs(5385);
    outputs(653) <= layer6_outputs(2526);
    outputs(654) <= not(layer6_outputs(10));
    outputs(655) <= not(layer6_outputs(5814)) or (layer6_outputs(3493));
    outputs(656) <= not(layer6_outputs(7127));
    outputs(657) <= not(layer6_outputs(2604));
    outputs(658) <= not(layer6_outputs(3952));
    outputs(659) <= (layer6_outputs(6175)) and not (layer6_outputs(3625));
    outputs(660) <= not(layer6_outputs(6944));
    outputs(661) <= layer6_outputs(6365);
    outputs(662) <= not((layer6_outputs(6003)) xor (layer6_outputs(147)));
    outputs(663) <= (layer6_outputs(6772)) xor (layer6_outputs(615));
    outputs(664) <= not((layer6_outputs(3185)) xor (layer6_outputs(1641)));
    outputs(665) <= layer6_outputs(3944);
    outputs(666) <= not(layer6_outputs(3773));
    outputs(667) <= (layer6_outputs(1807)) xor (layer6_outputs(898));
    outputs(668) <= layer6_outputs(6501);
    outputs(669) <= not(layer6_outputs(4396));
    outputs(670) <= not(layer6_outputs(5533));
    outputs(671) <= not(layer6_outputs(525));
    outputs(672) <= not(layer6_outputs(1157));
    outputs(673) <= not(layer6_outputs(7019));
    outputs(674) <= not(layer6_outputs(5976)) or (layer6_outputs(3157));
    outputs(675) <= (layer6_outputs(2264)) and not (layer6_outputs(3752));
    outputs(676) <= not((layer6_outputs(3000)) and (layer6_outputs(2366)));
    outputs(677) <= layer6_outputs(4322);
    outputs(678) <= layer6_outputs(7397);
    outputs(679) <= not((layer6_outputs(7006)) or (layer6_outputs(6808)));
    outputs(680) <= layer6_outputs(4717);
    outputs(681) <= layer6_outputs(7679);
    outputs(682) <= (layer6_outputs(433)) xor (layer6_outputs(5774));
    outputs(683) <= not(layer6_outputs(5447));
    outputs(684) <= not(layer6_outputs(3008));
    outputs(685) <= not(layer6_outputs(7016));
    outputs(686) <= (layer6_outputs(882)) xor (layer6_outputs(6241));
    outputs(687) <= (layer6_outputs(2731)) and (layer6_outputs(1069));
    outputs(688) <= layer6_outputs(5944);
    outputs(689) <= not(layer6_outputs(6384));
    outputs(690) <= not(layer6_outputs(6140));
    outputs(691) <= not(layer6_outputs(3912));
    outputs(692) <= not(layer6_outputs(4428));
    outputs(693) <= (layer6_outputs(156)) xor (layer6_outputs(3356));
    outputs(694) <= (layer6_outputs(4134)) and not (layer6_outputs(6040));
    outputs(695) <= (layer6_outputs(3456)) xor (layer6_outputs(2588));
    outputs(696) <= not(layer6_outputs(4479));
    outputs(697) <= not((layer6_outputs(3950)) or (layer6_outputs(4821)));
    outputs(698) <= not((layer6_outputs(3678)) xor (layer6_outputs(5870)));
    outputs(699) <= not((layer6_outputs(5814)) xor (layer6_outputs(734)));
    outputs(700) <= layer6_outputs(2426);
    outputs(701) <= (layer6_outputs(2046)) xor (layer6_outputs(3419));
    outputs(702) <= not((layer6_outputs(1630)) xor (layer6_outputs(7279)));
    outputs(703) <= (layer6_outputs(5900)) xor (layer6_outputs(5484));
    outputs(704) <= not(layer6_outputs(2336));
    outputs(705) <= not((layer6_outputs(6252)) xor (layer6_outputs(2176)));
    outputs(706) <= layer6_outputs(2940);
    outputs(707) <= layer6_outputs(1040);
    outputs(708) <= not(layer6_outputs(4622));
    outputs(709) <= (layer6_outputs(1542)) xor (layer6_outputs(3216));
    outputs(710) <= not(layer6_outputs(2277));
    outputs(711) <= not(layer6_outputs(2988));
    outputs(712) <= not(layer6_outputs(4994));
    outputs(713) <= not(layer6_outputs(3513));
    outputs(714) <= not((layer6_outputs(2769)) and (layer6_outputs(4524)));
    outputs(715) <= layer6_outputs(2810);
    outputs(716) <= not(layer6_outputs(2826));
    outputs(717) <= not((layer6_outputs(5922)) or (layer6_outputs(2142)));
    outputs(718) <= not(layer6_outputs(1710));
    outputs(719) <= not((layer6_outputs(6545)) xor (layer6_outputs(6547)));
    outputs(720) <= layer6_outputs(3177);
    outputs(721) <= not((layer6_outputs(263)) xor (layer6_outputs(6418)));
    outputs(722) <= not(layer6_outputs(4529));
    outputs(723) <= not(layer6_outputs(1510));
    outputs(724) <= layer6_outputs(6145);
    outputs(725) <= layer6_outputs(5682);
    outputs(726) <= layer6_outputs(1245);
    outputs(727) <= not((layer6_outputs(5885)) xor (layer6_outputs(7351)));
    outputs(728) <= not((layer6_outputs(240)) xor (layer6_outputs(2851)));
    outputs(729) <= layer6_outputs(5209);
    outputs(730) <= not(layer6_outputs(4334));
    outputs(731) <= layer6_outputs(5238);
    outputs(732) <= (layer6_outputs(4209)) xor (layer6_outputs(6888));
    outputs(733) <= layer6_outputs(5942);
    outputs(734) <= not(layer6_outputs(3130));
    outputs(735) <= layer6_outputs(5951);
    outputs(736) <= not(layer6_outputs(2435));
    outputs(737) <= layer6_outputs(924);
    outputs(738) <= not(layer6_outputs(5289));
    outputs(739) <= layer6_outputs(3565);
    outputs(740) <= (layer6_outputs(854)) xor (layer6_outputs(7196));
    outputs(741) <= layer6_outputs(6193);
    outputs(742) <= (layer6_outputs(1546)) xor (layer6_outputs(125));
    outputs(743) <= not(layer6_outputs(4455));
    outputs(744) <= not(layer6_outputs(1667));
    outputs(745) <= not((layer6_outputs(3244)) xor (layer6_outputs(5924)));
    outputs(746) <= (layer6_outputs(6651)) xor (layer6_outputs(6402));
    outputs(747) <= not((layer6_outputs(2113)) xor (layer6_outputs(6369)));
    outputs(748) <= layer6_outputs(5160);
    outputs(749) <= not(layer6_outputs(7042));
    outputs(750) <= not(layer6_outputs(7653));
    outputs(751) <= not((layer6_outputs(3282)) xor (layer6_outputs(6832)));
    outputs(752) <= layer6_outputs(1564);
    outputs(753) <= not(layer6_outputs(3150));
    outputs(754) <= not(layer6_outputs(330));
    outputs(755) <= not(layer6_outputs(2624));
    outputs(756) <= not((layer6_outputs(7078)) or (layer6_outputs(82)));
    outputs(757) <= not(layer6_outputs(6446));
    outputs(758) <= not(layer6_outputs(7267)) or (layer6_outputs(2451));
    outputs(759) <= not(layer6_outputs(1913));
    outputs(760) <= not(layer6_outputs(3644));
    outputs(761) <= not(layer6_outputs(4302));
    outputs(762) <= not(layer6_outputs(4120));
    outputs(763) <= layer6_outputs(2036);
    outputs(764) <= not((layer6_outputs(807)) xor (layer6_outputs(3052)));
    outputs(765) <= not(layer6_outputs(2757));
    outputs(766) <= (layer6_outputs(5307)) or (layer6_outputs(1997));
    outputs(767) <= (layer6_outputs(6235)) xor (layer6_outputs(4604));
    outputs(768) <= not(layer6_outputs(5378));
    outputs(769) <= not(layer6_outputs(7324));
    outputs(770) <= layer6_outputs(6692);
    outputs(771) <= not(layer6_outputs(6961));
    outputs(772) <= not((layer6_outputs(4175)) xor (layer6_outputs(5997)));
    outputs(773) <= layer6_outputs(6105);
    outputs(774) <= layer6_outputs(2898);
    outputs(775) <= layer6_outputs(6287);
    outputs(776) <= not((layer6_outputs(2762)) xor (layer6_outputs(3932)));
    outputs(777) <= not(layer6_outputs(7234));
    outputs(778) <= not((layer6_outputs(226)) xor (layer6_outputs(3837)));
    outputs(779) <= not((layer6_outputs(4041)) xor (layer6_outputs(5990)));
    outputs(780) <= not((layer6_outputs(3547)) xor (layer6_outputs(593)));
    outputs(781) <= not((layer6_outputs(5609)) xor (layer6_outputs(461)));
    outputs(782) <= layer6_outputs(4833);
    outputs(783) <= not(layer6_outputs(2182));
    outputs(784) <= not(layer6_outputs(3956));
    outputs(785) <= layer6_outputs(2987);
    outputs(786) <= not((layer6_outputs(7581)) xor (layer6_outputs(1960)));
    outputs(787) <= not(layer6_outputs(1387));
    outputs(788) <= layer6_outputs(5880);
    outputs(789) <= layer6_outputs(3074);
    outputs(790) <= (layer6_outputs(4333)) and not (layer6_outputs(100));
    outputs(791) <= layer6_outputs(3214);
    outputs(792) <= (layer6_outputs(7657)) xor (layer6_outputs(7568));
    outputs(793) <= not((layer6_outputs(2968)) xor (layer6_outputs(1377)));
    outputs(794) <= not(layer6_outputs(5426));
    outputs(795) <= not(layer6_outputs(3538));
    outputs(796) <= (layer6_outputs(7290)) and not (layer6_outputs(468));
    outputs(797) <= (layer6_outputs(2556)) and not (layer6_outputs(7593));
    outputs(798) <= not(layer6_outputs(1498));
    outputs(799) <= not(layer6_outputs(7227));
    outputs(800) <= layer6_outputs(5868);
    outputs(801) <= (layer6_outputs(328)) xor (layer6_outputs(1178));
    outputs(802) <= layer6_outputs(4059);
    outputs(803) <= (layer6_outputs(5928)) and not (layer6_outputs(7461));
    outputs(804) <= (layer6_outputs(7203)) xor (layer6_outputs(2292));
    outputs(805) <= not((layer6_outputs(3057)) xor (layer6_outputs(2843)));
    outputs(806) <= not((layer6_outputs(5144)) xor (layer6_outputs(5990)));
    outputs(807) <= not(layer6_outputs(835));
    outputs(808) <= (layer6_outputs(1978)) xor (layer6_outputs(4660));
    outputs(809) <= layer6_outputs(2546);
    outputs(810) <= not(layer6_outputs(6524));
    outputs(811) <= (layer6_outputs(4416)) and (layer6_outputs(437));
    outputs(812) <= not((layer6_outputs(6935)) or (layer6_outputs(2995)));
    outputs(813) <= not(layer6_outputs(4173));
    outputs(814) <= not(layer6_outputs(6348));
    outputs(815) <= (layer6_outputs(4893)) and (layer6_outputs(740));
    outputs(816) <= not(layer6_outputs(5663));
    outputs(817) <= not(layer6_outputs(2053)) or (layer6_outputs(4007));
    outputs(818) <= layer6_outputs(920);
    outputs(819) <= not(layer6_outputs(577));
    outputs(820) <= not((layer6_outputs(5683)) xor (layer6_outputs(5665)));
    outputs(821) <= not(layer6_outputs(4913));
    outputs(822) <= not(layer6_outputs(2153));
    outputs(823) <= not((layer6_outputs(3391)) xor (layer6_outputs(6630)));
    outputs(824) <= (layer6_outputs(5055)) xor (layer6_outputs(5129));
    outputs(825) <= not((layer6_outputs(4115)) xor (layer6_outputs(2206)));
    outputs(826) <= '0';
    outputs(827) <= (layer6_outputs(1158)) and (layer6_outputs(4103));
    outputs(828) <= layer6_outputs(7419);
    outputs(829) <= layer6_outputs(6020);
    outputs(830) <= (layer6_outputs(7574)) and not (layer6_outputs(1083));
    outputs(831) <= not(layer6_outputs(5107));
    outputs(832) <= not((layer6_outputs(4937)) xor (layer6_outputs(1917)));
    outputs(833) <= (layer6_outputs(1053)) xor (layer6_outputs(4297));
    outputs(834) <= not(layer6_outputs(6019));
    outputs(835) <= (layer6_outputs(3930)) and not (layer6_outputs(3033));
    outputs(836) <= layer6_outputs(1342);
    outputs(837) <= layer6_outputs(4509);
    outputs(838) <= not(layer6_outputs(6423));
    outputs(839) <= not((layer6_outputs(2224)) xor (layer6_outputs(976)));
    outputs(840) <= layer6_outputs(37);
    outputs(841) <= not((layer6_outputs(4781)) xor (layer6_outputs(612)));
    outputs(842) <= layer6_outputs(4174);
    outputs(843) <= not(layer6_outputs(7044));
    outputs(844) <= not(layer6_outputs(3869)) or (layer6_outputs(336));
    outputs(845) <= layer6_outputs(6904);
    outputs(846) <= not((layer6_outputs(768)) xor (layer6_outputs(7389)));
    outputs(847) <= not((layer6_outputs(5113)) xor (layer6_outputs(1507)));
    outputs(848) <= (layer6_outputs(3631)) and not (layer6_outputs(5910));
    outputs(849) <= not(layer6_outputs(4303));
    outputs(850) <= layer6_outputs(3379);
    outputs(851) <= not(layer6_outputs(4650));
    outputs(852) <= layer6_outputs(3112);
    outputs(853) <= (layer6_outputs(3309)) xor (layer6_outputs(5962));
    outputs(854) <= not(layer6_outputs(7621));
    outputs(855) <= layer6_outputs(1728);
    outputs(856) <= not((layer6_outputs(2359)) xor (layer6_outputs(3013)));
    outputs(857) <= not(layer6_outputs(23));
    outputs(858) <= not(layer6_outputs(5537)) or (layer6_outputs(5416));
    outputs(859) <= layer6_outputs(60);
    outputs(860) <= (layer6_outputs(2829)) xor (layer6_outputs(4125));
    outputs(861) <= not(layer6_outputs(2200));
    outputs(862) <= (layer6_outputs(1712)) and (layer6_outputs(1226));
    outputs(863) <= (layer6_outputs(604)) and not (layer6_outputs(7573));
    outputs(864) <= layer6_outputs(6783);
    outputs(865) <= layer6_outputs(11);
    outputs(866) <= (layer6_outputs(3685)) and not (layer6_outputs(6463));
    outputs(867) <= not(layer6_outputs(3440));
    outputs(868) <= not(layer6_outputs(7499));
    outputs(869) <= not(layer6_outputs(3677));
    outputs(870) <= not(layer6_outputs(155));
    outputs(871) <= layer6_outputs(2376);
    outputs(872) <= (layer6_outputs(2499)) xor (layer6_outputs(5946));
    outputs(873) <= not((layer6_outputs(4331)) xor (layer6_outputs(4598)));
    outputs(874) <= (layer6_outputs(4378)) and not (layer6_outputs(5407));
    outputs(875) <= not((layer6_outputs(7490)) xor (layer6_outputs(6510)));
    outputs(876) <= (layer6_outputs(1795)) or (layer6_outputs(2642));
    outputs(877) <= (layer6_outputs(372)) and not (layer6_outputs(4342));
    outputs(878) <= layer6_outputs(7357);
    outputs(879) <= not(layer6_outputs(6247));
    outputs(880) <= not(layer6_outputs(3804));
    outputs(881) <= not(layer6_outputs(343));
    outputs(882) <= layer6_outputs(6774);
    outputs(883) <= not(layer6_outputs(5330));
    outputs(884) <= (layer6_outputs(6677)) and not (layer6_outputs(1540));
    outputs(885) <= not(layer6_outputs(105));
    outputs(886) <= layer6_outputs(410);
    outputs(887) <= not(layer6_outputs(2684));
    outputs(888) <= not(layer6_outputs(6628));
    outputs(889) <= layer6_outputs(3127);
    outputs(890) <= not(layer6_outputs(6356));
    outputs(891) <= not((layer6_outputs(1486)) xor (layer6_outputs(6701)));
    outputs(892) <= not(layer6_outputs(3534));
    outputs(893) <= layer6_outputs(595);
    outputs(894) <= layer6_outputs(6684);
    outputs(895) <= not((layer6_outputs(597)) xor (layer6_outputs(2261)));
    outputs(896) <= layer6_outputs(3544);
    outputs(897) <= (layer6_outputs(1838)) and not (layer6_outputs(5563));
    outputs(898) <= not((layer6_outputs(6620)) xor (layer6_outputs(6478)));
    outputs(899) <= (layer6_outputs(6673)) xor (layer6_outputs(4302));
    outputs(900) <= (layer6_outputs(5387)) and not (layer6_outputs(210));
    outputs(901) <= (layer6_outputs(2554)) and (layer6_outputs(320));
    outputs(902) <= not(layer6_outputs(1296));
    outputs(903) <= not(layer6_outputs(2862));
    outputs(904) <= not((layer6_outputs(7566)) xor (layer6_outputs(5056)));
    outputs(905) <= layer6_outputs(1545);
    outputs(906) <= layer6_outputs(7176);
    outputs(907) <= (layer6_outputs(2468)) and not (layer6_outputs(3));
    outputs(908) <= (layer6_outputs(970)) or (layer6_outputs(3616));
    outputs(909) <= (layer6_outputs(4122)) and (layer6_outputs(7145));
    outputs(910) <= layer6_outputs(7630);
    outputs(911) <= (layer6_outputs(804)) xor (layer6_outputs(6784));
    outputs(912) <= not((layer6_outputs(1396)) and (layer6_outputs(6393)));
    outputs(913) <= not(layer6_outputs(6539));
    outputs(914) <= (layer6_outputs(4615)) xor (layer6_outputs(7361));
    outputs(915) <= layer6_outputs(3241);
    outputs(916) <= (layer6_outputs(1334)) xor (layer6_outputs(1507));
    outputs(917) <= not((layer6_outputs(4156)) xor (layer6_outputs(2923)));
    outputs(918) <= not(layer6_outputs(5331));
    outputs(919) <= not(layer6_outputs(4506));
    outputs(920) <= layer6_outputs(1062);
    outputs(921) <= (layer6_outputs(6056)) xor (layer6_outputs(6515));
    outputs(922) <= (layer6_outputs(1967)) and not (layer6_outputs(3654));
    outputs(923) <= not(layer6_outputs(5491));
    outputs(924) <= not(layer6_outputs(2625));
    outputs(925) <= layer6_outputs(6085);
    outputs(926) <= (layer6_outputs(1451)) and not (layer6_outputs(3925));
    outputs(927) <= layer6_outputs(6109);
    outputs(928) <= not(layer6_outputs(2943));
    outputs(929) <= not(layer6_outputs(1601));
    outputs(930) <= (layer6_outputs(4830)) and not (layer6_outputs(6043));
    outputs(931) <= layer6_outputs(5564);
    outputs(932) <= not(layer6_outputs(4956));
    outputs(933) <= not((layer6_outputs(5350)) xor (layer6_outputs(5444)));
    outputs(934) <= layer6_outputs(4808);
    outputs(935) <= layer6_outputs(792);
    outputs(936) <= (layer6_outputs(6099)) and (layer6_outputs(2844));
    outputs(937) <= layer6_outputs(4669);
    outputs(938) <= (layer6_outputs(2786)) and (layer6_outputs(3751));
    outputs(939) <= (layer6_outputs(7036)) and not (layer6_outputs(3238));
    outputs(940) <= (layer6_outputs(7145)) xor (layer6_outputs(7015));
    outputs(941) <= not((layer6_outputs(6256)) xor (layer6_outputs(4816)));
    outputs(942) <= not(layer6_outputs(2684));
    outputs(943) <= layer6_outputs(3892);
    outputs(944) <= not(layer6_outputs(7208));
    outputs(945) <= not((layer6_outputs(1240)) xor (layer6_outputs(5233)));
    outputs(946) <= not(layer6_outputs(4627));
    outputs(947) <= not(layer6_outputs(4300));
    outputs(948) <= not((layer6_outputs(3723)) xor (layer6_outputs(5366)));
    outputs(949) <= not(layer6_outputs(2884));
    outputs(950) <= not(layer6_outputs(342));
    outputs(951) <= layer6_outputs(6519);
    outputs(952) <= (layer6_outputs(4922)) xor (layer6_outputs(1127));
    outputs(953) <= (layer6_outputs(7033)) xor (layer6_outputs(4599));
    outputs(954) <= layer6_outputs(2927);
    outputs(955) <= layer6_outputs(1263);
    outputs(956) <= not(layer6_outputs(4135)) or (layer6_outputs(4086));
    outputs(957) <= layer6_outputs(4316);
    outputs(958) <= not(layer6_outputs(6820));
    outputs(959) <= (layer6_outputs(4700)) and not (layer6_outputs(1952));
    outputs(960) <= not((layer6_outputs(7248)) xor (layer6_outputs(4879)));
    outputs(961) <= (layer6_outputs(5523)) xor (layer6_outputs(7298));
    outputs(962) <= not(layer6_outputs(3426));
    outputs(963) <= not((layer6_outputs(6103)) xor (layer6_outputs(6878)));
    outputs(964) <= not(layer6_outputs(7062));
    outputs(965) <= not(layer6_outputs(2227));
    outputs(966) <= (layer6_outputs(3500)) xor (layer6_outputs(4202));
    outputs(967) <= not(layer6_outputs(5558));
    outputs(968) <= layer6_outputs(1164);
    outputs(969) <= not(layer6_outputs(876));
    outputs(970) <= not(layer6_outputs(335)) or (layer6_outputs(4505));
    outputs(971) <= layer6_outputs(5811);
    outputs(972) <= (layer6_outputs(4198)) xor (layer6_outputs(5152));
    outputs(973) <= not(layer6_outputs(3837));
    outputs(974) <= not(layer6_outputs(7493));
    outputs(975) <= (layer6_outputs(7525)) and (layer6_outputs(6164));
    outputs(976) <= (layer6_outputs(3849)) and not (layer6_outputs(6989));
    outputs(977) <= not((layer6_outputs(2964)) xor (layer6_outputs(4062)));
    outputs(978) <= layer6_outputs(3737);
    outputs(979) <= layer6_outputs(6794);
    outputs(980) <= (layer6_outputs(2590)) and not (layer6_outputs(6108));
    outputs(981) <= (layer6_outputs(5618)) xor (layer6_outputs(3646));
    outputs(982) <= (layer6_outputs(2707)) and not (layer6_outputs(3636));
    outputs(983) <= not((layer6_outputs(6900)) or (layer6_outputs(1403)));
    outputs(984) <= not(layer6_outputs(3866));
    outputs(985) <= (layer6_outputs(6522)) and not (layer6_outputs(1191));
    outputs(986) <= layer6_outputs(4449);
    outputs(987) <= layer6_outputs(7175);
    outputs(988) <= not(layer6_outputs(1830));
    outputs(989) <= not((layer6_outputs(3932)) or (layer6_outputs(7669)));
    outputs(990) <= not(layer6_outputs(2638));
    outputs(991) <= (layer6_outputs(5187)) and (layer6_outputs(4077));
    outputs(992) <= (layer6_outputs(1595)) and not (layer6_outputs(1307));
    outputs(993) <= not(layer6_outputs(6456));
    outputs(994) <= layer6_outputs(5499);
    outputs(995) <= (layer6_outputs(7228)) xor (layer6_outputs(3206));
    outputs(996) <= not(layer6_outputs(764));
    outputs(997) <= (layer6_outputs(2396)) xor (layer6_outputs(4945));
    outputs(998) <= not(layer6_outputs(7400)) or (layer6_outputs(7519));
    outputs(999) <= layer6_outputs(2348);
    outputs(1000) <= not(layer6_outputs(6422));
    outputs(1001) <= not(layer6_outputs(6578));
    outputs(1002) <= not(layer6_outputs(7520));
    outputs(1003) <= not((layer6_outputs(1430)) xor (layer6_outputs(4711)));
    outputs(1004) <= not(layer6_outputs(2768));
    outputs(1005) <= not(layer6_outputs(6626)) or (layer6_outputs(1280));
    outputs(1006) <= (layer6_outputs(3333)) xor (layer6_outputs(1582));
    outputs(1007) <= layer6_outputs(701);
    outputs(1008) <= (layer6_outputs(3234)) and not (layer6_outputs(5704));
    outputs(1009) <= not((layer6_outputs(5338)) xor (layer6_outputs(1098)));
    outputs(1010) <= not(layer6_outputs(2536));
    outputs(1011) <= (layer6_outputs(1032)) and (layer6_outputs(286));
    outputs(1012) <= not(layer6_outputs(5192));
    outputs(1013) <= (layer6_outputs(1896)) xor (layer6_outputs(713));
    outputs(1014) <= (layer6_outputs(3259)) xor (layer6_outputs(6475));
    outputs(1015) <= not((layer6_outputs(4812)) and (layer6_outputs(2782)));
    outputs(1016) <= not((layer6_outputs(2633)) or (layer6_outputs(3590)));
    outputs(1017) <= not(layer6_outputs(5203));
    outputs(1018) <= layer6_outputs(692);
    outputs(1019) <= layer6_outputs(3106);
    outputs(1020) <= not(layer6_outputs(2568));
    outputs(1021) <= layer6_outputs(6610);
    outputs(1022) <= layer6_outputs(5098);
    outputs(1023) <= layer6_outputs(7460);
    outputs(1024) <= (layer6_outputs(823)) and not (layer6_outputs(1790));
    outputs(1025) <= not(layer6_outputs(3909));
    outputs(1026) <= layer6_outputs(2981);
    outputs(1027) <= not(layer6_outputs(1606));
    outputs(1028) <= (layer6_outputs(4510)) xor (layer6_outputs(6975));
    outputs(1029) <= not(layer6_outputs(969));
    outputs(1030) <= not((layer6_outputs(3552)) xor (layer6_outputs(3657)));
    outputs(1031) <= not(layer6_outputs(5749));
    outputs(1032) <= (layer6_outputs(5791)) and (layer6_outputs(1936));
    outputs(1033) <= (layer6_outputs(940)) xor (layer6_outputs(1686));
    outputs(1034) <= layer6_outputs(262);
    outputs(1035) <= not(layer6_outputs(5332));
    outputs(1036) <= (layer6_outputs(1478)) xor (layer6_outputs(5293));
    outputs(1037) <= layer6_outputs(6923);
    outputs(1038) <= (layer6_outputs(6980)) xor (layer6_outputs(2037));
    outputs(1039) <= not(layer6_outputs(1642));
    outputs(1040) <= (layer6_outputs(4852)) and not (layer6_outputs(2799));
    outputs(1041) <= not((layer6_outputs(2850)) xor (layer6_outputs(663)));
    outputs(1042) <= (layer6_outputs(4447)) xor (layer6_outputs(3451));
    outputs(1043) <= not(layer6_outputs(4873));
    outputs(1044) <= not(layer6_outputs(3902)) or (layer6_outputs(6));
    outputs(1045) <= not((layer6_outputs(3967)) or (layer6_outputs(5022)));
    outputs(1046) <= not(layer6_outputs(5348));
    outputs(1047) <= not((layer6_outputs(3615)) xor (layer6_outputs(3078)));
    outputs(1048) <= not(layer6_outputs(2355));
    outputs(1049) <= layer6_outputs(5342);
    outputs(1050) <= not(layer6_outputs(4483));
    outputs(1051) <= not((layer6_outputs(4728)) xor (layer6_outputs(5537)));
    outputs(1052) <= not(layer6_outputs(279));
    outputs(1053) <= layer6_outputs(7243);
    outputs(1054) <= layer6_outputs(2737);
    outputs(1055) <= (layer6_outputs(1186)) and not (layer6_outputs(591));
    outputs(1056) <= not(layer6_outputs(5942));
    outputs(1057) <= layer6_outputs(1196);
    outputs(1058) <= not((layer6_outputs(5509)) xor (layer6_outputs(880)));
    outputs(1059) <= (layer6_outputs(7016)) and not (layer6_outputs(4163));
    outputs(1060) <= not(layer6_outputs(4127));
    outputs(1061) <= not(layer6_outputs(7194)) or (layer6_outputs(4662));
    outputs(1062) <= (layer6_outputs(1055)) and not (layer6_outputs(69));
    outputs(1063) <= not((layer6_outputs(7655)) xor (layer6_outputs(886)));
    outputs(1064) <= layer6_outputs(5154);
    outputs(1065) <= layer6_outputs(2622);
    outputs(1066) <= (layer6_outputs(2948)) or (layer6_outputs(7021));
    outputs(1067) <= not(layer6_outputs(2087));
    outputs(1068) <= (layer6_outputs(2561)) xor (layer6_outputs(950));
    outputs(1069) <= not(layer6_outputs(1998));
    outputs(1070) <= layer6_outputs(6681);
    outputs(1071) <= (layer6_outputs(3661)) and not (layer6_outputs(2188));
    outputs(1072) <= layer6_outputs(4806);
    outputs(1073) <= (layer6_outputs(5145)) xor (layer6_outputs(5991));
    outputs(1074) <= layer6_outputs(3102);
    outputs(1075) <= not(layer6_outputs(5660));
    outputs(1076) <= not(layer6_outputs(5620));
    outputs(1077) <= not((layer6_outputs(2401)) xor (layer6_outputs(1533)));
    outputs(1078) <= (layer6_outputs(1758)) and not (layer6_outputs(2172));
    outputs(1079) <= not(layer6_outputs(7627));
    outputs(1080) <= layer6_outputs(1160);
    outputs(1081) <= not(layer6_outputs(1989));
    outputs(1082) <= (layer6_outputs(2043)) xor (layer6_outputs(1195));
    outputs(1083) <= (layer6_outputs(6342)) and not (layer6_outputs(7221));
    outputs(1084) <= (layer6_outputs(3101)) and (layer6_outputs(7468));
    outputs(1085) <= layer6_outputs(3328);
    outputs(1086) <= (layer6_outputs(2605)) xor (layer6_outputs(7450));
    outputs(1087) <= (layer6_outputs(2120)) xor (layer6_outputs(2483));
    outputs(1088) <= not(layer6_outputs(5090));
    outputs(1089) <= not(layer6_outputs(6364));
    outputs(1090) <= layer6_outputs(6723);
    outputs(1091) <= layer6_outputs(2489);
    outputs(1092) <= layer6_outputs(3273);
    outputs(1093) <= layer6_outputs(1550);
    outputs(1094) <= layer6_outputs(339);
    outputs(1095) <= not(layer6_outputs(3286));
    outputs(1096) <= (layer6_outputs(1216)) xor (layer6_outputs(4501));
    outputs(1097) <= not(layer6_outputs(6007));
    outputs(1098) <= layer6_outputs(813);
    outputs(1099) <= not(layer6_outputs(3353));
    outputs(1100) <= layer6_outputs(6534);
    outputs(1101) <= not(layer6_outputs(1639));
    outputs(1102) <= layer6_outputs(4332);
    outputs(1103) <= not(layer6_outputs(7222));
    outputs(1104) <= layer6_outputs(6701);
    outputs(1105) <= (layer6_outputs(3962)) xor (layer6_outputs(5429));
    outputs(1106) <= layer6_outputs(409);
    outputs(1107) <= not(layer6_outputs(1530));
    outputs(1108) <= not((layer6_outputs(2212)) or (layer6_outputs(7478)));
    outputs(1109) <= (layer6_outputs(7169)) and not (layer6_outputs(7637));
    outputs(1110) <= not(layer6_outputs(3492));
    outputs(1111) <= not((layer6_outputs(5501)) or (layer6_outputs(2820)));
    outputs(1112) <= layer6_outputs(1394);
    outputs(1113) <= not((layer6_outputs(5186)) xor (layer6_outputs(4280)));
    outputs(1114) <= (layer6_outputs(6880)) or (layer6_outputs(1957));
    outputs(1115) <= not(layer6_outputs(2485));
    outputs(1116) <= layer6_outputs(3472);
    outputs(1117) <= not(layer6_outputs(2922));
    outputs(1118) <= layer6_outputs(6678);
    outputs(1119) <= not((layer6_outputs(3294)) xor (layer6_outputs(5350)));
    outputs(1120) <= not(layer6_outputs(4143));
    outputs(1121) <= layer6_outputs(6435);
    outputs(1122) <= (layer6_outputs(5450)) xor (layer6_outputs(4807));
    outputs(1123) <= layer6_outputs(6934);
    outputs(1124) <= (layer6_outputs(5431)) xor (layer6_outputs(2212));
    outputs(1125) <= (layer6_outputs(2498)) xor (layer6_outputs(5509));
    outputs(1126) <= (layer6_outputs(5288)) or (layer6_outputs(4857));
    outputs(1127) <= layer6_outputs(4469);
    outputs(1128) <= layer6_outputs(569);
    outputs(1129) <= layer6_outputs(1634);
    outputs(1130) <= not(layer6_outputs(2682)) or (layer6_outputs(2463));
    outputs(1131) <= layer6_outputs(6815);
    outputs(1132) <= not(layer6_outputs(6298)) or (layer6_outputs(2198));
    outputs(1133) <= not(layer6_outputs(6900)) or (layer6_outputs(7667));
    outputs(1134) <= (layer6_outputs(5515)) xor (layer6_outputs(4681));
    outputs(1135) <= not(layer6_outputs(5561));
    outputs(1136) <= not(layer6_outputs(6100));
    outputs(1137) <= (layer6_outputs(4946)) and not (layer6_outputs(3222));
    outputs(1138) <= layer6_outputs(2464);
    outputs(1139) <= layer6_outputs(3876);
    outputs(1140) <= not((layer6_outputs(2496)) xor (layer6_outputs(7597)));
    outputs(1141) <= (layer6_outputs(7672)) and (layer6_outputs(1623));
    outputs(1142) <= not((layer6_outputs(4119)) xor (layer6_outputs(4749)));
    outputs(1143) <= (layer6_outputs(5668)) and not (layer6_outputs(6856));
    outputs(1144) <= not((layer6_outputs(5878)) xor (layer6_outputs(7436)));
    outputs(1145) <= layer6_outputs(4790);
    outputs(1146) <= (layer6_outputs(5317)) and (layer6_outputs(520));
    outputs(1147) <= not((layer6_outputs(3961)) or (layer6_outputs(6469)));
    outputs(1148) <= (layer6_outputs(5951)) and not (layer6_outputs(3967));
    outputs(1149) <= (layer6_outputs(3323)) and (layer6_outputs(1572));
    outputs(1150) <= (layer6_outputs(4314)) and not (layer6_outputs(2294));
    outputs(1151) <= not(layer6_outputs(5400)) or (layer6_outputs(3548));
    outputs(1152) <= (layer6_outputs(1247)) xor (layer6_outputs(1290));
    outputs(1153) <= layer6_outputs(5697);
    outputs(1154) <= layer6_outputs(2947);
    outputs(1155) <= (layer6_outputs(177)) xor (layer6_outputs(4957));
    outputs(1156) <= not(layer6_outputs(6077));
    outputs(1157) <= (layer6_outputs(6618)) and not (layer6_outputs(3798));
    outputs(1158) <= not(layer6_outputs(6976));
    outputs(1159) <= (layer6_outputs(6647)) xor (layer6_outputs(124));
    outputs(1160) <= not((layer6_outputs(6740)) xor (layer6_outputs(4293)));
    outputs(1161) <= not(layer6_outputs(5670));
    outputs(1162) <= (layer6_outputs(3187)) xor (layer6_outputs(2223));
    outputs(1163) <= layer6_outputs(4958);
    outputs(1164) <= not(layer6_outputs(4323));
    outputs(1165) <= layer6_outputs(1925);
    outputs(1166) <= layer6_outputs(4522);
    outputs(1167) <= not(layer6_outputs(5484));
    outputs(1168) <= not((layer6_outputs(280)) xor (layer6_outputs(1972)));
    outputs(1169) <= not(layer6_outputs(6334));
    outputs(1170) <= layer6_outputs(7124);
    outputs(1171) <= not(layer6_outputs(2958));
    outputs(1172) <= not(layer6_outputs(2356));
    outputs(1173) <= not((layer6_outputs(4404)) xor (layer6_outputs(7086)));
    outputs(1174) <= (layer6_outputs(7341)) xor (layer6_outputs(2093));
    outputs(1175) <= (layer6_outputs(5597)) and (layer6_outputs(5183));
    outputs(1176) <= layer6_outputs(2316);
    outputs(1177) <= not((layer6_outputs(2108)) xor (layer6_outputs(3544)));
    outputs(1178) <= layer6_outputs(4289);
    outputs(1179) <= not(layer6_outputs(2334));
    outputs(1180) <= (layer6_outputs(235)) and not (layer6_outputs(2567));
    outputs(1181) <= not(layer6_outputs(2723));
    outputs(1182) <= layer6_outputs(4899);
    outputs(1183) <= (layer6_outputs(7659)) and not (layer6_outputs(572));
    outputs(1184) <= (layer6_outputs(5524)) and (layer6_outputs(369));
    outputs(1185) <= (layer6_outputs(4423)) and not (layer6_outputs(402));
    outputs(1186) <= (layer6_outputs(4915)) xor (layer6_outputs(5827));
    outputs(1187) <= not(layer6_outputs(3840));
    outputs(1188) <= not((layer6_outputs(5211)) or (layer6_outputs(6443)));
    outputs(1189) <= not(layer6_outputs(1755));
    outputs(1190) <= layer6_outputs(7099);
    outputs(1191) <= layer6_outputs(3117);
    outputs(1192) <= (layer6_outputs(6331)) and (layer6_outputs(4822));
    outputs(1193) <= (layer6_outputs(7360)) or (layer6_outputs(49));
    outputs(1194) <= not(layer6_outputs(7677));
    outputs(1195) <= (layer6_outputs(3060)) xor (layer6_outputs(7538));
    outputs(1196) <= not((layer6_outputs(6534)) xor (layer6_outputs(7479)));
    outputs(1197) <= layer6_outputs(7442);
    outputs(1198) <= layer6_outputs(7040);
    outputs(1199) <= not(layer6_outputs(3600));
    outputs(1200) <= layer6_outputs(6898);
    outputs(1201) <= layer6_outputs(1901);
    outputs(1202) <= not((layer6_outputs(5552)) xor (layer6_outputs(7133)));
    outputs(1203) <= layer6_outputs(925);
    outputs(1204) <= layer6_outputs(6934);
    outputs(1205) <= (layer6_outputs(230)) and not (layer6_outputs(6773));
    outputs(1206) <= not((layer6_outputs(2594)) or (layer6_outputs(6702)));
    outputs(1207) <= layer6_outputs(6226);
    outputs(1208) <= layer6_outputs(5015);
    outputs(1209) <= not(layer6_outputs(7296));
    outputs(1210) <= not(layer6_outputs(5270));
    outputs(1211) <= not((layer6_outputs(3115)) or (layer6_outputs(6204)));
    outputs(1212) <= not((layer6_outputs(4466)) xor (layer6_outputs(6409)));
    outputs(1213) <= not((layer6_outputs(1722)) xor (layer6_outputs(2720)));
    outputs(1214) <= not((layer6_outputs(6172)) xor (layer6_outputs(7142)));
    outputs(1215) <= (layer6_outputs(4392)) xor (layer6_outputs(2521));
    outputs(1216) <= layer6_outputs(2584);
    outputs(1217) <= not(layer6_outputs(6142));
    outputs(1218) <= not(layer6_outputs(6862));
    outputs(1219) <= not((layer6_outputs(5193)) xor (layer6_outputs(3393)));
    outputs(1220) <= layer6_outputs(7558);
    outputs(1221) <= (layer6_outputs(5824)) and (layer6_outputs(2977));
    outputs(1222) <= layer6_outputs(5739);
    outputs(1223) <= not(layer6_outputs(5878));
    outputs(1224) <= not(layer6_outputs(1182));
    outputs(1225) <= not((layer6_outputs(2012)) xor (layer6_outputs(2664)));
    outputs(1226) <= not(layer6_outputs(1685));
    outputs(1227) <= not(layer6_outputs(4743));
    outputs(1228) <= not(layer6_outputs(2092));
    outputs(1229) <= layer6_outputs(5957);
    outputs(1230) <= layer6_outputs(2385);
    outputs(1231) <= not(layer6_outputs(1939));
    outputs(1232) <= layer6_outputs(6272);
    outputs(1233) <= not(layer6_outputs(4814));
    outputs(1234) <= not(layer6_outputs(4200));
    outputs(1235) <= layer6_outputs(4547);
    outputs(1236) <= (layer6_outputs(2287)) and not (layer6_outputs(1704));
    outputs(1237) <= (layer6_outputs(1756)) and not (layer6_outputs(1005));
    outputs(1238) <= layer6_outputs(7594);
    outputs(1239) <= not(layer6_outputs(3656));
    outputs(1240) <= layer6_outputs(6828);
    outputs(1241) <= (layer6_outputs(5534)) xor (layer6_outputs(2005));
    outputs(1242) <= (layer6_outputs(4133)) and not (layer6_outputs(6664));
    outputs(1243) <= (layer6_outputs(6570)) and not (layer6_outputs(1583));
    outputs(1244) <= layer6_outputs(6449);
    outputs(1245) <= not((layer6_outputs(7235)) or (layer6_outputs(3984)));
    outputs(1246) <= layer6_outputs(3681);
    outputs(1247) <= (layer6_outputs(7530)) and (layer6_outputs(6457));
    outputs(1248) <= not(layer6_outputs(7456));
    outputs(1249) <= not((layer6_outputs(5281)) xor (layer6_outputs(2433)));
    outputs(1250) <= (layer6_outputs(4959)) xor (layer6_outputs(4053));
    outputs(1251) <= (layer6_outputs(906)) xor (layer6_outputs(5283));
    outputs(1252) <= layer6_outputs(4630);
    outputs(1253) <= not((layer6_outputs(4457)) xor (layer6_outputs(4366)));
    outputs(1254) <= not(layer6_outputs(3316));
    outputs(1255) <= layer6_outputs(6133);
    outputs(1256) <= (layer6_outputs(7612)) xor (layer6_outputs(5344));
    outputs(1257) <= layer6_outputs(1865);
    outputs(1258) <= not(layer6_outputs(4812)) or (layer6_outputs(7529));
    outputs(1259) <= not((layer6_outputs(5364)) xor (layer6_outputs(5119)));
    outputs(1260) <= not(layer6_outputs(5935));
    outputs(1261) <= layer6_outputs(2926);
    outputs(1262) <= layer6_outputs(4980);
    outputs(1263) <= not(layer6_outputs(6158));
    outputs(1264) <= layer6_outputs(7572);
    outputs(1265) <= layer6_outputs(2783);
    outputs(1266) <= (layer6_outputs(6597)) and not (layer6_outputs(211));
    outputs(1267) <= not(layer6_outputs(5418)) or (layer6_outputs(667));
    outputs(1268) <= (layer6_outputs(7390)) and (layer6_outputs(2148));
    outputs(1269) <= not((layer6_outputs(4409)) xor (layer6_outputs(2290)));
    outputs(1270) <= (layer6_outputs(7354)) and not (layer6_outputs(6382));
    outputs(1271) <= (layer6_outputs(6405)) and not (layer6_outputs(7417));
    outputs(1272) <= not(layer6_outputs(283));
    outputs(1273) <= layer6_outputs(5280);
    outputs(1274) <= layer6_outputs(366);
    outputs(1275) <= (layer6_outputs(3954)) xor (layer6_outputs(5979));
    outputs(1276) <= (layer6_outputs(4443)) and not (layer6_outputs(7611));
    outputs(1277) <= not((layer6_outputs(2755)) xor (layer6_outputs(2306)));
    outputs(1278) <= layer6_outputs(2976);
    outputs(1279) <= layer6_outputs(7591);
    outputs(1280) <= not(layer6_outputs(819));
    outputs(1281) <= (layer6_outputs(4955)) xor (layer6_outputs(1886));
    outputs(1282) <= not(layer6_outputs(209));
    outputs(1283) <= layer6_outputs(5122);
    outputs(1284) <= layer6_outputs(1305);
    outputs(1285) <= not(layer6_outputs(4206));
    outputs(1286) <= layer6_outputs(315);
    outputs(1287) <= not(layer6_outputs(5876));
    outputs(1288) <= not((layer6_outputs(4991)) xor (layer6_outputs(2064)));
    outputs(1289) <= (layer6_outputs(6837)) xor (layer6_outputs(5823));
    outputs(1290) <= layer6_outputs(6907);
    outputs(1291) <= layer6_outputs(7387);
    outputs(1292) <= not(layer6_outputs(5242));
    outputs(1293) <= layer6_outputs(5116);
    outputs(1294) <= not((layer6_outputs(5586)) xor (layer6_outputs(7139)));
    outputs(1295) <= not(layer6_outputs(7031));
    outputs(1296) <= not((layer6_outputs(1359)) xor (layer6_outputs(3479)));
    outputs(1297) <= layer6_outputs(4255);
    outputs(1298) <= (layer6_outputs(6714)) and not (layer6_outputs(5151));
    outputs(1299) <= (layer6_outputs(4182)) and not (layer6_outputs(557));
    outputs(1300) <= not(layer6_outputs(316));
    outputs(1301) <= (layer6_outputs(841)) xor (layer6_outputs(975));
    outputs(1302) <= layer6_outputs(596);
    outputs(1303) <= not(layer6_outputs(2315));
    outputs(1304) <= layer6_outputs(4536);
    outputs(1305) <= not(layer6_outputs(5705)) or (layer6_outputs(6953));
    outputs(1306) <= layer6_outputs(1573);
    outputs(1307) <= not(layer6_outputs(6443));
    outputs(1308) <= not((layer6_outputs(4042)) xor (layer6_outputs(7511)));
    outputs(1309) <= not((layer6_outputs(2704)) xor (layer6_outputs(2969)));
    outputs(1310) <= (layer6_outputs(1584)) xor (layer6_outputs(5925));
    outputs(1311) <= not(layer6_outputs(6445));
    outputs(1312) <= layer6_outputs(7477);
    outputs(1313) <= (layer6_outputs(4243)) and (layer6_outputs(2112));
    outputs(1314) <= not(layer6_outputs(932));
    outputs(1315) <= not(layer6_outputs(5527));
    outputs(1316) <= not((layer6_outputs(2055)) xor (layer6_outputs(5136)));
    outputs(1317) <= not(layer6_outputs(2842)) or (layer6_outputs(5494));
    outputs(1318) <= layer6_outputs(1259);
    outputs(1319) <= layer6_outputs(1419);
    outputs(1320) <= not(layer6_outputs(2257));
    outputs(1321) <= not(layer6_outputs(3559));
    outputs(1322) <= (layer6_outputs(6381)) and (layer6_outputs(4651));
    outputs(1323) <= (layer6_outputs(7413)) and not (layer6_outputs(3025));
    outputs(1324) <= layer6_outputs(6049);
    outputs(1325) <= layer6_outputs(1562);
    outputs(1326) <= (layer6_outputs(4552)) xor (layer6_outputs(940));
    outputs(1327) <= not((layer6_outputs(3668)) or (layer6_outputs(1792)));
    outputs(1328) <= not(layer6_outputs(6562));
    outputs(1329) <= not(layer6_outputs(6173));
    outputs(1330) <= (layer6_outputs(2580)) xor (layer6_outputs(4523));
    outputs(1331) <= layer6_outputs(3893);
    outputs(1332) <= layer6_outputs(4668);
    outputs(1333) <= (layer6_outputs(4624)) xor (layer6_outputs(1226));
    outputs(1334) <= layer6_outputs(3522);
    outputs(1335) <= not((layer6_outputs(1662)) xor (layer6_outputs(7491)));
    outputs(1336) <= not(layer6_outputs(4131));
    outputs(1337) <= not(layer6_outputs(3589));
    outputs(1338) <= (layer6_outputs(5469)) xor (layer6_outputs(2013));
    outputs(1339) <= layer6_outputs(2312);
    outputs(1340) <= (layer6_outputs(1274)) and not (layer6_outputs(2472));
    outputs(1341) <= layer6_outputs(1716);
    outputs(1342) <= layer6_outputs(5794);
    outputs(1343) <= not(layer6_outputs(6380));
    outputs(1344) <= layer6_outputs(4184);
    outputs(1345) <= (layer6_outputs(4711)) and not (layer6_outputs(358));
    outputs(1346) <= layer6_outputs(7667);
    outputs(1347) <= layer6_outputs(7675);
    outputs(1348) <= layer6_outputs(7154);
    outputs(1349) <= not(layer6_outputs(6317));
    outputs(1350) <= not((layer6_outputs(1466)) or (layer6_outputs(4486)));
    outputs(1351) <= not((layer6_outputs(1392)) xor (layer6_outputs(5839)));
    outputs(1352) <= not(layer6_outputs(1193));
    outputs(1353) <= not((layer6_outputs(3223)) xor (layer6_outputs(4841)));
    outputs(1354) <= not(layer6_outputs(2389));
    outputs(1355) <= layer6_outputs(7124);
    outputs(1356) <= layer6_outputs(2934);
    outputs(1357) <= not(layer6_outputs(6579));
    outputs(1358) <= layer6_outputs(5360);
    outputs(1359) <= not((layer6_outputs(3888)) or (layer6_outputs(2540)));
    outputs(1360) <= not(layer6_outputs(4665));
    outputs(1361) <= layer6_outputs(6655);
    outputs(1362) <= layer6_outputs(2080);
    outputs(1363) <= layer6_outputs(617);
    outputs(1364) <= layer6_outputs(752);
    outputs(1365) <= not((layer6_outputs(6560)) xor (layer6_outputs(4515)));
    outputs(1366) <= (layer6_outputs(5165)) xor (layer6_outputs(7051));
    outputs(1367) <= (layer6_outputs(4967)) and (layer6_outputs(6943));
    outputs(1368) <= layer6_outputs(2667);
    outputs(1369) <= (layer6_outputs(501)) and (layer6_outputs(6985));
    outputs(1370) <= (layer6_outputs(6208)) and not (layer6_outputs(5367));
    outputs(1371) <= not((layer6_outputs(7250)) xor (layer6_outputs(5496)));
    outputs(1372) <= layer6_outputs(215);
    outputs(1373) <= (layer6_outputs(571)) xor (layer6_outputs(7266));
    outputs(1374) <= (layer6_outputs(7459)) xor (layer6_outputs(423));
    outputs(1375) <= not((layer6_outputs(6415)) xor (layer6_outputs(5247)));
    outputs(1376) <= layer6_outputs(5369);
    outputs(1377) <= not((layer6_outputs(6068)) or (layer6_outputs(1876)));
    outputs(1378) <= (layer6_outputs(4114)) xor (layer6_outputs(6091));
    outputs(1379) <= (layer6_outputs(6858)) xor (layer6_outputs(6992));
    outputs(1380) <= layer6_outputs(7257);
    outputs(1381) <= not(layer6_outputs(7434));
    outputs(1382) <= (layer6_outputs(144)) and not (layer6_outputs(3109));
    outputs(1383) <= not(layer6_outputs(1729));
    outputs(1384) <= not((layer6_outputs(4744)) xor (layer6_outputs(2897)));
    outputs(1385) <= layer6_outputs(4179);
    outputs(1386) <= layer6_outputs(6692);
    outputs(1387) <= not((layer6_outputs(842)) xor (layer6_outputs(4018)));
    outputs(1388) <= not(layer6_outputs(5938));
    outputs(1389) <= not(layer6_outputs(2503));
    outputs(1390) <= (layer6_outputs(3625)) and (layer6_outputs(3198));
    outputs(1391) <= not(layer6_outputs(4686)) or (layer6_outputs(1181));
    outputs(1392) <= (layer6_outputs(3664)) and not (layer6_outputs(4842));
    outputs(1393) <= (layer6_outputs(436)) xor (layer6_outputs(6044));
    outputs(1394) <= layer6_outputs(1864);
    outputs(1395) <= not(layer6_outputs(6247));
    outputs(1396) <= not(layer6_outputs(7617));
    outputs(1397) <= not((layer6_outputs(994)) xor (layer6_outputs(3365)));
    outputs(1398) <= layer6_outputs(4222);
    outputs(1399) <= layer6_outputs(6663);
    outputs(1400) <= not((layer6_outputs(6428)) or (layer6_outputs(3516)));
    outputs(1401) <= (layer6_outputs(7500)) xor (layer6_outputs(5895));
    outputs(1402) <= (layer6_outputs(3834)) xor (layer6_outputs(1882));
    outputs(1403) <= (layer6_outputs(7512)) or (layer6_outputs(3187));
    outputs(1404) <= layer6_outputs(5552);
    outputs(1405) <= not(layer6_outputs(2330));
    outputs(1406) <= not(layer6_outputs(2059));
    outputs(1407) <= (layer6_outputs(47)) xor (layer6_outputs(3381));
    outputs(1408) <= not(layer6_outputs(1971));
    outputs(1409) <= (layer6_outputs(4763)) xor (layer6_outputs(173));
    outputs(1410) <= not(layer6_outputs(5844));
    outputs(1411) <= (layer6_outputs(2690)) and not (layer6_outputs(6579));
    outputs(1412) <= not(layer6_outputs(4125));
    outputs(1413) <= not(layer6_outputs(7095));
    outputs(1414) <= not(layer6_outputs(3726));
    outputs(1415) <= not(layer6_outputs(1265));
    outputs(1416) <= (layer6_outputs(5084)) xor (layer6_outputs(6721));
    outputs(1417) <= layer6_outputs(1918);
    outputs(1418) <= layer6_outputs(3090);
    outputs(1419) <= not(layer6_outputs(1987));
    outputs(1420) <= not(layer6_outputs(4131));
    outputs(1421) <= layer6_outputs(1663);
    outputs(1422) <= not((layer6_outputs(746)) xor (layer6_outputs(2420)));
    outputs(1423) <= not(layer6_outputs(6876)) or (layer6_outputs(6639));
    outputs(1424) <= not(layer6_outputs(3731));
    outputs(1425) <= layer6_outputs(3821);
    outputs(1426) <= not((layer6_outputs(7096)) xor (layer6_outputs(3047)));
    outputs(1427) <= (layer6_outputs(3011)) and not (layer6_outputs(762));
    outputs(1428) <= (layer6_outputs(2078)) xor (layer6_outputs(7368));
    outputs(1429) <= (layer6_outputs(3542)) and not (layer6_outputs(3899));
    outputs(1430) <= layer6_outputs(1190);
    outputs(1431) <= not(layer6_outputs(4983));
    outputs(1432) <= not(layer6_outputs(5974));
    outputs(1433) <= not(layer6_outputs(3547));
    outputs(1434) <= not(layer6_outputs(459));
    outputs(1435) <= layer6_outputs(2348);
    outputs(1436) <= not(layer6_outputs(389));
    outputs(1437) <= (layer6_outputs(406)) xor (layer6_outputs(6418));
    outputs(1438) <= not(layer6_outputs(1472));
    outputs(1439) <= layer6_outputs(6283);
    outputs(1440) <= layer6_outputs(6792);
    outputs(1441) <= layer6_outputs(2902);
    outputs(1442) <= (layer6_outputs(6714)) and not (layer6_outputs(1785));
    outputs(1443) <= layer6_outputs(2582);
    outputs(1444) <= (layer6_outputs(4573)) xor (layer6_outputs(7166));
    outputs(1445) <= not((layer6_outputs(5019)) xor (layer6_outputs(2638)));
    outputs(1446) <= layer6_outputs(3515);
    outputs(1447) <= (layer6_outputs(5064)) and not (layer6_outputs(5090));
    outputs(1448) <= not((layer6_outputs(1825)) or (layer6_outputs(3044)));
    outputs(1449) <= not(layer6_outputs(5389));
    outputs(1450) <= layer6_outputs(3947);
    outputs(1451) <= layer6_outputs(3363);
    outputs(1452) <= layer6_outputs(5383);
    outputs(1453) <= layer6_outputs(912);
    outputs(1454) <= not(layer6_outputs(157));
    outputs(1455) <= (layer6_outputs(2354)) xor (layer6_outputs(725));
    outputs(1456) <= layer6_outputs(5130);
    outputs(1457) <= (layer6_outputs(3369)) and not (layer6_outputs(4646));
    outputs(1458) <= (layer6_outputs(4222)) xor (layer6_outputs(3340));
    outputs(1459) <= not(layer6_outputs(3092));
    outputs(1460) <= not((layer6_outputs(3585)) xor (layer6_outputs(3452)));
    outputs(1461) <= layer6_outputs(4623);
    outputs(1462) <= not(layer6_outputs(4738));
    outputs(1463) <= (layer6_outputs(2429)) xor (layer6_outputs(1925));
    outputs(1464) <= (layer6_outputs(3409)) or (layer6_outputs(1519));
    outputs(1465) <= not((layer6_outputs(2833)) or (layer6_outputs(6464)));
    outputs(1466) <= layer6_outputs(6815);
    outputs(1467) <= (layer6_outputs(1617)) and not (layer6_outputs(4587));
    outputs(1468) <= layer6_outputs(6315);
    outputs(1469) <= layer6_outputs(2930);
    outputs(1470) <= not(layer6_outputs(1848));
    outputs(1471) <= not((layer6_outputs(1520)) xor (layer6_outputs(4901)));
    outputs(1472) <= not((layer6_outputs(4504)) xor (layer6_outputs(4360)));
    outputs(1473) <= not((layer6_outputs(4501)) xor (layer6_outputs(6322)));
    outputs(1474) <= layer6_outputs(1260);
    outputs(1475) <= not(layer6_outputs(1393));
    outputs(1476) <= not(layer6_outputs(2675));
    outputs(1477) <= (layer6_outputs(1154)) xor (layer6_outputs(2230));
    outputs(1478) <= not(layer6_outputs(7508));
    outputs(1479) <= not(layer6_outputs(6513)) or (layer6_outputs(5017));
    outputs(1480) <= layer6_outputs(1713);
    outputs(1481) <= layer6_outputs(5265);
    outputs(1482) <= (layer6_outputs(7209)) xor (layer6_outputs(7030));
    outputs(1483) <= not(layer6_outputs(4736));
    outputs(1484) <= (layer6_outputs(4674)) xor (layer6_outputs(5448));
    outputs(1485) <= layer6_outputs(1183);
    outputs(1486) <= not((layer6_outputs(5167)) xor (layer6_outputs(542)));
    outputs(1487) <= layer6_outputs(4185);
    outputs(1488) <= not((layer6_outputs(7211)) and (layer6_outputs(5462)));
    outputs(1489) <= layer6_outputs(6321);
    outputs(1490) <= (layer6_outputs(3819)) xor (layer6_outputs(3412));
    outputs(1491) <= layer6_outputs(3739);
    outputs(1492) <= layer6_outputs(215);
    outputs(1493) <= layer6_outputs(4336);
    outputs(1494) <= not((layer6_outputs(5400)) xor (layer6_outputs(1356)));
    outputs(1495) <= not(layer6_outputs(6177));
    outputs(1496) <= not(layer6_outputs(3579));
    outputs(1497) <= (layer6_outputs(6414)) xor (layer6_outputs(4412));
    outputs(1498) <= (layer6_outputs(3454)) xor (layer6_outputs(4704));
    outputs(1499) <= not((layer6_outputs(6779)) xor (layer6_outputs(535)));
    outputs(1500) <= not(layer6_outputs(3880));
    outputs(1501) <= (layer6_outputs(712)) and not (layer6_outputs(2077));
    outputs(1502) <= layer6_outputs(3633);
    outputs(1503) <= (layer6_outputs(7368)) xor (layer6_outputs(3044));
    outputs(1504) <= layer6_outputs(3403);
    outputs(1505) <= layer6_outputs(7408);
    outputs(1506) <= layer6_outputs(6770);
    outputs(1507) <= (layer6_outputs(916)) xor (layer6_outputs(6263));
    outputs(1508) <= not(layer6_outputs(5266)) or (layer6_outputs(7477));
    outputs(1509) <= layer6_outputs(5905);
    outputs(1510) <= (layer6_outputs(688)) and (layer6_outputs(1928));
    outputs(1511) <= layer6_outputs(989);
    outputs(1512) <= layer6_outputs(3872);
    outputs(1513) <= not((layer6_outputs(5216)) xor (layer6_outputs(4266)));
    outputs(1514) <= not(layer6_outputs(7150));
    outputs(1515) <= layer6_outputs(4668);
    outputs(1516) <= not((layer6_outputs(2111)) or (layer6_outputs(2744)));
    outputs(1517) <= layer6_outputs(7020);
    outputs(1518) <= not((layer6_outputs(1500)) or (layer6_outputs(7194)));
    outputs(1519) <= not(layer6_outputs(41));
    outputs(1520) <= layer6_outputs(5328);
    outputs(1521) <= not((layer6_outputs(1387)) xor (layer6_outputs(2162)));
    outputs(1522) <= not((layer6_outputs(1902)) xor (layer6_outputs(7549)));
    outputs(1523) <= '0';
    outputs(1524) <= not(layer6_outputs(610));
    outputs(1525) <= not(layer6_outputs(2024));
    outputs(1526) <= not((layer6_outputs(4088)) xor (layer6_outputs(4421)));
    outputs(1527) <= not(layer6_outputs(1091));
    outputs(1528) <= (layer6_outputs(3404)) xor (layer6_outputs(295));
    outputs(1529) <= not(layer6_outputs(1772));
    outputs(1530) <= (layer6_outputs(7518)) xor (layer6_outputs(6667));
    outputs(1531) <= not(layer6_outputs(2594));
    outputs(1532) <= layer6_outputs(2429);
    outputs(1533) <= layer6_outputs(322);
    outputs(1534) <= layer6_outputs(3783);
    outputs(1535) <= layer6_outputs(4602);
    outputs(1536) <= not((layer6_outputs(1903)) xor (layer6_outputs(3775)));
    outputs(1537) <= not(layer6_outputs(6190));
    outputs(1538) <= layer6_outputs(5661);
    outputs(1539) <= layer6_outputs(277);
    outputs(1540) <= layer6_outputs(711);
    outputs(1541) <= (layer6_outputs(2197)) or (layer6_outputs(5829));
    outputs(1542) <= not(layer6_outputs(1725));
    outputs(1543) <= layer6_outputs(5489);
    outputs(1544) <= (layer6_outputs(7190)) and not (layer6_outputs(1306));
    outputs(1545) <= not(layer6_outputs(3857));
    outputs(1546) <= not(layer6_outputs(2950));
    outputs(1547) <= layer6_outputs(4664);
    outputs(1548) <= not(layer6_outputs(5326)) or (layer6_outputs(2));
    outputs(1549) <= not(layer6_outputs(68));
    outputs(1550) <= not(layer6_outputs(2208)) or (layer6_outputs(4833));
    outputs(1551) <= not(layer6_outputs(6979));
    outputs(1552) <= not(layer6_outputs(5641));
    outputs(1553) <= not((layer6_outputs(3952)) and (layer6_outputs(312)));
    outputs(1554) <= layer6_outputs(7269);
    outputs(1555) <= layer6_outputs(354);
    outputs(1556) <= layer6_outputs(3884);
    outputs(1557) <= not(layer6_outputs(5839));
    outputs(1558) <= layer6_outputs(4318);
    outputs(1559) <= not(layer6_outputs(939));
    outputs(1560) <= not(layer6_outputs(2526));
    outputs(1561) <= not(layer6_outputs(1498));
    outputs(1562) <= layer6_outputs(6490);
    outputs(1563) <= not(layer6_outputs(4917));
    outputs(1564) <= not(layer6_outputs(2767));
    outputs(1565) <= not(layer6_outputs(4760));
    outputs(1566) <= not(layer6_outputs(4789));
    outputs(1567) <= not(layer6_outputs(5103));
    outputs(1568) <= not(layer6_outputs(6925)) or (layer6_outputs(3982));
    outputs(1569) <= not(layer6_outputs(1148));
    outputs(1570) <= (layer6_outputs(6770)) xor (layer6_outputs(198));
    outputs(1571) <= not(layer6_outputs(530));
    outputs(1572) <= (layer6_outputs(978)) xor (layer6_outputs(4787));
    outputs(1573) <= layer6_outputs(5475);
    outputs(1574) <= not(layer6_outputs(4913));
    outputs(1575) <= (layer6_outputs(6970)) xor (layer6_outputs(5708));
    outputs(1576) <= (layer6_outputs(2434)) xor (layer6_outputs(7052));
    outputs(1577) <= (layer6_outputs(395)) and not (layer6_outputs(6824));
    outputs(1578) <= not(layer6_outputs(619)) or (layer6_outputs(207));
    outputs(1579) <= (layer6_outputs(1757)) xor (layer6_outputs(4113));
    outputs(1580) <= not(layer6_outputs(6642)) or (layer6_outputs(7590));
    outputs(1581) <= (layer6_outputs(1272)) and not (layer6_outputs(1209));
    outputs(1582) <= (layer6_outputs(7555)) xor (layer6_outputs(4426));
    outputs(1583) <= (layer6_outputs(3253)) and (layer6_outputs(3866));
    outputs(1584) <= not(layer6_outputs(4378));
    outputs(1585) <= not(layer6_outputs(3903)) or (layer6_outputs(6959));
    outputs(1586) <= not((layer6_outputs(7613)) xor (layer6_outputs(5887)));
    outputs(1587) <= not(layer6_outputs(4935));
    outputs(1588) <= (layer6_outputs(7249)) or (layer6_outputs(4085));
    outputs(1589) <= not((layer6_outputs(270)) xor (layer6_outputs(5598)));
    outputs(1590) <= not(layer6_outputs(5048));
    outputs(1591) <= not((layer6_outputs(1284)) xor (layer6_outputs(7021)));
    outputs(1592) <= not(layer6_outputs(1731));
    outputs(1593) <= not((layer6_outputs(2105)) xor (layer6_outputs(2295)));
    outputs(1594) <= layer6_outputs(859);
    outputs(1595) <= layer6_outputs(3529);
    outputs(1596) <= (layer6_outputs(1438)) xor (layer6_outputs(6666));
    outputs(1597) <= not(layer6_outputs(4771));
    outputs(1598) <= not(layer6_outputs(412));
    outputs(1599) <= (layer6_outputs(1090)) or (layer6_outputs(7550));
    outputs(1600) <= not(layer6_outputs(1948));
    outputs(1601) <= layer6_outputs(128);
    outputs(1602) <= not(layer6_outputs(340));
    outputs(1603) <= (layer6_outputs(5960)) xor (layer6_outputs(7496));
    outputs(1604) <= layer6_outputs(2082);
    outputs(1605) <= layer6_outputs(1807);
    outputs(1606) <= not(layer6_outputs(5908));
    outputs(1607) <= not(layer6_outputs(405)) or (layer6_outputs(3628));
    outputs(1608) <= (layer6_outputs(11)) xor (layer6_outputs(5272));
    outputs(1609) <= (layer6_outputs(6389)) or (layer6_outputs(4341));
    outputs(1610) <= (layer6_outputs(5423)) xor (layer6_outputs(6048));
    outputs(1611) <= not(layer6_outputs(1120));
    outputs(1612) <= not(layer6_outputs(7152));
    outputs(1613) <= (layer6_outputs(5655)) xor (layer6_outputs(1558));
    outputs(1614) <= not(layer6_outputs(6429));
    outputs(1615) <= not((layer6_outputs(4055)) xor (layer6_outputs(2293)));
    outputs(1616) <= not(layer6_outputs(4585));
    outputs(1617) <= layer6_outputs(6854);
    outputs(1618) <= not(layer6_outputs(3614));
    outputs(1619) <= not((layer6_outputs(1852)) xor (layer6_outputs(4035)));
    outputs(1620) <= not(layer6_outputs(7168));
    outputs(1621) <= not(layer6_outputs(4912));
    outputs(1622) <= not((layer6_outputs(2093)) xor (layer6_outputs(1766)));
    outputs(1623) <= not(layer6_outputs(6777));
    outputs(1624) <= not(layer6_outputs(7291)) or (layer6_outputs(6541));
    outputs(1625) <= layer6_outputs(5954);
    outputs(1626) <= not((layer6_outputs(290)) xor (layer6_outputs(2651)));
    outputs(1627) <= not(layer6_outputs(6481));
    outputs(1628) <= not((layer6_outputs(6129)) or (layer6_outputs(2554)));
    outputs(1629) <= not((layer6_outputs(5593)) xor (layer6_outputs(7439)));
    outputs(1630) <= not(layer6_outputs(5666));
    outputs(1631) <= not(layer6_outputs(5885));
    outputs(1632) <= (layer6_outputs(5916)) xor (layer6_outputs(2633));
    outputs(1633) <= (layer6_outputs(6230)) and (layer6_outputs(3890));
    outputs(1634) <= not(layer6_outputs(6768));
    outputs(1635) <= layer6_outputs(3233);
    outputs(1636) <= (layer6_outputs(3350)) and not (layer6_outputs(7606));
    outputs(1637) <= layer6_outputs(7263);
    outputs(1638) <= not((layer6_outputs(3959)) xor (layer6_outputs(3299)));
    outputs(1639) <= (layer6_outputs(3570)) and not (layer6_outputs(3597));
    outputs(1640) <= layer6_outputs(2610);
    outputs(1641) <= not(layer6_outputs(5952));
    outputs(1642) <= (layer6_outputs(6552)) and not (layer6_outputs(832));
    outputs(1643) <= not(layer6_outputs(3794));
    outputs(1644) <= layer6_outputs(4967);
    outputs(1645) <= (layer6_outputs(1632)) xor (layer6_outputs(684));
    outputs(1646) <= not(layer6_outputs(2868));
    outputs(1647) <= (layer6_outputs(2981)) xor (layer6_outputs(4920));
    outputs(1648) <= (layer6_outputs(518)) and not (layer6_outputs(7043));
    outputs(1649) <= (layer6_outputs(5694)) xor (layer6_outputs(5334));
    outputs(1650) <= not((layer6_outputs(34)) xor (layer6_outputs(4599)));
    outputs(1651) <= layer6_outputs(2626);
    outputs(1652) <= not(layer6_outputs(4453));
    outputs(1653) <= (layer6_outputs(2458)) and (layer6_outputs(6920));
    outputs(1654) <= not(layer6_outputs(1914));
    outputs(1655) <= (layer6_outputs(6398)) xor (layer6_outputs(1459));
    outputs(1656) <= layer6_outputs(95);
    outputs(1657) <= not((layer6_outputs(1722)) xor (layer6_outputs(2270)));
    outputs(1658) <= layer6_outputs(4969);
    outputs(1659) <= not(layer6_outputs(2789));
    outputs(1660) <= not(layer6_outputs(874));
    outputs(1661) <= layer6_outputs(3763);
    outputs(1662) <= layer6_outputs(220);
    outputs(1663) <= layer6_outputs(3424);
    outputs(1664) <= not(layer6_outputs(4641));
    outputs(1665) <= layer6_outputs(524);
    outputs(1666) <= layer6_outputs(3365);
    outputs(1667) <= not((layer6_outputs(1622)) xor (layer6_outputs(7322)));
    outputs(1668) <= not(layer6_outputs(4712));
    outputs(1669) <= layer6_outputs(3895);
    outputs(1670) <= (layer6_outputs(1087)) xor (layer6_outputs(4840));
    outputs(1671) <= layer6_outputs(4853);
    outputs(1672) <= not(layer6_outputs(6469));
    outputs(1673) <= not(layer6_outputs(2519));
    outputs(1674) <= not((layer6_outputs(2511)) xor (layer6_outputs(766)));
    outputs(1675) <= not(layer6_outputs(6150));
    outputs(1676) <= not((layer6_outputs(5547)) and (layer6_outputs(6938)));
    outputs(1677) <= layer6_outputs(2608);
    outputs(1678) <= layer6_outputs(2857);
    outputs(1679) <= layer6_outputs(3225);
    outputs(1680) <= layer6_outputs(2023);
    outputs(1681) <= (layer6_outputs(3349)) and not (layer6_outputs(1010));
    outputs(1682) <= not((layer6_outputs(930)) or (layer6_outputs(2842)));
    outputs(1683) <= layer6_outputs(5526);
    outputs(1684) <= not(layer6_outputs(5613));
    outputs(1685) <= not(layer6_outputs(3891)) or (layer6_outputs(5848));
    outputs(1686) <= not((layer6_outputs(2971)) xor (layer6_outputs(3023)));
    outputs(1687) <= (layer6_outputs(3082)) xor (layer6_outputs(2029));
    outputs(1688) <= not(layer6_outputs(1351));
    outputs(1689) <= not(layer6_outputs(284));
    outputs(1690) <= not(layer6_outputs(2683));
    outputs(1691) <= (layer6_outputs(206)) xor (layer6_outputs(6804));
    outputs(1692) <= (layer6_outputs(5379)) or (layer6_outputs(151));
    outputs(1693) <= layer6_outputs(5251);
    outputs(1694) <= layer6_outputs(1980);
    outputs(1695) <= not(layer6_outputs(5361));
    outputs(1696) <= layer6_outputs(3616);
    outputs(1697) <= layer6_outputs(2308);
    outputs(1698) <= not(layer6_outputs(3437));
    outputs(1699) <= not(layer6_outputs(2222));
    outputs(1700) <= not((layer6_outputs(1142)) xor (layer6_outputs(645)));
    outputs(1701) <= layer6_outputs(5105);
    outputs(1702) <= (layer6_outputs(7594)) and (layer6_outputs(1259));
    outputs(1703) <= (layer6_outputs(3598)) xor (layer6_outputs(7410));
    outputs(1704) <= layer6_outputs(6441);
    outputs(1705) <= not((layer6_outputs(3773)) and (layer6_outputs(2705)));
    outputs(1706) <= not(layer6_outputs(6972));
    outputs(1707) <= not(layer6_outputs(249));
    outputs(1708) <= (layer6_outputs(6936)) and not (layer6_outputs(3848));
    outputs(1709) <= (layer6_outputs(6067)) or (layer6_outputs(4242));
    outputs(1710) <= layer6_outputs(6814);
    outputs(1711) <= not(layer6_outputs(1530));
    outputs(1712) <= layer6_outputs(7079);
    outputs(1713) <= not(layer6_outputs(1003));
    outputs(1714) <= (layer6_outputs(7444)) xor (layer6_outputs(6709));
    outputs(1715) <= not((layer6_outputs(455)) xor (layer6_outputs(5919)));
    outputs(1716) <= (layer6_outputs(3054)) or (layer6_outputs(6101));
    outputs(1717) <= not(layer6_outputs(5371));
    outputs(1718) <= (layer6_outputs(361)) and not (layer6_outputs(2272));
    outputs(1719) <= layer6_outputs(7494);
    outputs(1720) <= not(layer6_outputs(6525));
    outputs(1721) <= (layer6_outputs(6350)) and (layer6_outputs(4057));
    outputs(1722) <= layer6_outputs(7620);
    outputs(1723) <= not(layer6_outputs(3519));
    outputs(1724) <= layer6_outputs(2498);
    outputs(1725) <= layer6_outputs(752);
    outputs(1726) <= not(layer6_outputs(7343)) or (layer6_outputs(1529));
    outputs(1727) <= not(layer6_outputs(6425));
    outputs(1728) <= layer6_outputs(864);
    outputs(1729) <= layer6_outputs(4584);
    outputs(1730) <= not((layer6_outputs(1224)) and (layer6_outputs(7433)));
    outputs(1731) <= not(layer6_outputs(1845));
    outputs(1732) <= not(layer6_outputs(333));
    outputs(1733) <= not(layer6_outputs(7371));
    outputs(1734) <= layer6_outputs(4324);
    outputs(1735) <= layer6_outputs(7375);
    outputs(1736) <= not(layer6_outputs(5719));
    outputs(1737) <= (layer6_outputs(790)) xor (layer6_outputs(5162));
    outputs(1738) <= not(layer6_outputs(6169));
    outputs(1739) <= layer6_outputs(6654);
    outputs(1740) <= not(layer6_outputs(1705));
    outputs(1741) <= (layer6_outputs(7356)) xor (layer6_outputs(1469));
    outputs(1742) <= not(layer6_outputs(2340)) or (layer6_outputs(6160));
    outputs(1743) <= not(layer6_outputs(3487));
    outputs(1744) <= not(layer6_outputs(1148));
    outputs(1745) <= (layer6_outputs(4574)) and not (layer6_outputs(2675));
    outputs(1746) <= layer6_outputs(3392);
    outputs(1747) <= not(layer6_outputs(7425));
    outputs(1748) <= not(layer6_outputs(3329));
    outputs(1749) <= not(layer6_outputs(4389));
    outputs(1750) <= not((layer6_outputs(2383)) xor (layer6_outputs(4039)));
    outputs(1751) <= not(layer6_outputs(5239));
    outputs(1752) <= layer6_outputs(3395);
    outputs(1753) <= not(layer6_outputs(452));
    outputs(1754) <= layer6_outputs(2307);
    outputs(1755) <= not(layer6_outputs(4632));
    outputs(1756) <= not(layer6_outputs(4399));
    outputs(1757) <= not((layer6_outputs(3153)) xor (layer6_outputs(7117)));
    outputs(1758) <= (layer6_outputs(5217)) and not (layer6_outputs(4885));
    outputs(1759) <= not(layer6_outputs(6730));
    outputs(1760) <= not(layer6_outputs(463));
    outputs(1761) <= not((layer6_outputs(5492)) xor (layer6_outputs(370)));
    outputs(1762) <= layer6_outputs(2437);
    outputs(1763) <= not(layer6_outputs(2749));
    outputs(1764) <= not(layer6_outputs(861));
    outputs(1765) <= layer6_outputs(918);
    outputs(1766) <= not(layer6_outputs(3855));
    outputs(1767) <= layer6_outputs(519);
    outputs(1768) <= not(layer6_outputs(4973));
    outputs(1769) <= not((layer6_outputs(6853)) xor (layer6_outputs(5395)));
    outputs(1770) <= not(layer6_outputs(3686));
    outputs(1771) <= layer6_outputs(4424);
    outputs(1772) <= layer6_outputs(786);
    outputs(1773) <= not(layer6_outputs(5443));
    outputs(1774) <= (layer6_outputs(7093)) and not (layer6_outputs(4794));
    outputs(1775) <= layer6_outputs(2546);
    outputs(1776) <= layer6_outputs(1888);
    outputs(1777) <= not(layer6_outputs(6875));
    outputs(1778) <= not(layer6_outputs(5933));
    outputs(1779) <= not((layer6_outputs(5037)) xor (layer6_outputs(4258)));
    outputs(1780) <= (layer6_outputs(2889)) xor (layer6_outputs(2942));
    outputs(1781) <= layer6_outputs(7243);
    outputs(1782) <= not(layer6_outputs(5244));
    outputs(1783) <= layer6_outputs(7377);
    outputs(1784) <= not(layer6_outputs(6677)) or (layer6_outputs(2820));
    outputs(1785) <= not(layer6_outputs(7522));
    outputs(1786) <= (layer6_outputs(3120)) xor (layer6_outputs(589));
    outputs(1787) <= layer6_outputs(180);
    outputs(1788) <= (layer6_outputs(4075)) xor (layer6_outputs(6524));
    outputs(1789) <= layer6_outputs(3323);
    outputs(1790) <= not(layer6_outputs(5208));
    outputs(1791) <= layer6_outputs(5284);
    outputs(1792) <= not(layer6_outputs(6308));
    outputs(1793) <= layer6_outputs(4386);
    outputs(1794) <= not((layer6_outputs(6259)) xor (layer6_outputs(3925)));
    outputs(1795) <= not((layer6_outputs(182)) or (layer6_outputs(1526)));
    outputs(1796) <= layer6_outputs(5111);
    outputs(1797) <= not(layer6_outputs(1123));
    outputs(1798) <= layer6_outputs(7638);
    outputs(1799) <= not(layer6_outputs(234));
    outputs(1800) <= not(layer6_outputs(6140));
    outputs(1801) <= layer6_outputs(555);
    outputs(1802) <= layer6_outputs(7387);
    outputs(1803) <= layer6_outputs(5146);
    outputs(1804) <= layer6_outputs(4550);
    outputs(1805) <= layer6_outputs(1800);
    outputs(1806) <= not(layer6_outputs(7106));
    outputs(1807) <= not(layer6_outputs(5545));
    outputs(1808) <= (layer6_outputs(7223)) xor (layer6_outputs(4708));
    outputs(1809) <= not((layer6_outputs(5579)) xor (layer6_outputs(6511)));
    outputs(1810) <= (layer6_outputs(423)) and (layer6_outputs(786));
    outputs(1811) <= not(layer6_outputs(4155)) or (layer6_outputs(2049));
    outputs(1812) <= not(layer6_outputs(4372));
    outputs(1813) <= not(layer6_outputs(5397));
    outputs(1814) <= not(layer6_outputs(282));
    outputs(1815) <= (layer6_outputs(1958)) xor (layer6_outputs(6758));
    outputs(1816) <= not(layer6_outputs(2817));
    outputs(1817) <= layer6_outputs(7073);
    outputs(1818) <= (layer6_outputs(5927)) and not (layer6_outputs(2701));
    outputs(1819) <= not((layer6_outputs(1349)) xor (layer6_outputs(2774)));
    outputs(1820) <= (layer6_outputs(531)) xor (layer6_outputs(6130));
    outputs(1821) <= layer6_outputs(2974);
    outputs(1822) <= not(layer6_outputs(5967)) or (layer6_outputs(7379));
    outputs(1823) <= (layer6_outputs(5183)) xor (layer6_outputs(809));
    outputs(1824) <= layer6_outputs(6329);
    outputs(1825) <= not(layer6_outputs(7164));
    outputs(1826) <= not(layer6_outputs(3309));
    outputs(1827) <= (layer6_outputs(4500)) xor (layer6_outputs(4246));
    outputs(1828) <= layer6_outputs(649);
    outputs(1829) <= layer6_outputs(3144);
    outputs(1830) <= (layer6_outputs(7442)) and not (layer6_outputs(5721));
    outputs(1831) <= not(layer6_outputs(4652)) or (layer6_outputs(3976));
    outputs(1832) <= not((layer6_outputs(7157)) xor (layer6_outputs(1033)));
    outputs(1833) <= not(layer6_outputs(4565));
    outputs(1834) <= not(layer6_outputs(5664));
    outputs(1835) <= layer6_outputs(724);
    outputs(1836) <= (layer6_outputs(6514)) xor (layer6_outputs(897));
    outputs(1837) <= not((layer6_outputs(5723)) xor (layer6_outputs(6314)));
    outputs(1838) <= layer6_outputs(5707);
    outputs(1839) <= not(layer6_outputs(4396));
    outputs(1840) <= layer6_outputs(4164);
    outputs(1841) <= not((layer6_outputs(5551)) xor (layer6_outputs(4555)));
    outputs(1842) <= not(layer6_outputs(4029));
    outputs(1843) <= not(layer6_outputs(2787)) or (layer6_outputs(2125));
    outputs(1844) <= not((layer6_outputs(5457)) xor (layer6_outputs(3971)));
    outputs(1845) <= not(layer6_outputs(5724));
    outputs(1846) <= layer6_outputs(4321);
    outputs(1847) <= not(layer6_outputs(5194));
    outputs(1848) <= layer6_outputs(1422);
    outputs(1849) <= (layer6_outputs(1772)) and (layer6_outputs(4531));
    outputs(1850) <= layer6_outputs(2718);
    outputs(1851) <= layer6_outputs(1034);
    outputs(1852) <= not(layer6_outputs(2234));
    outputs(1853) <= layer6_outputs(3872);
    outputs(1854) <= not(layer6_outputs(4863));
    outputs(1855) <= layer6_outputs(2168);
    outputs(1856) <= (layer6_outputs(7065)) xor (layer6_outputs(5535));
    outputs(1857) <= layer6_outputs(7386);
    outputs(1858) <= layer6_outputs(5892);
    outputs(1859) <= not(layer6_outputs(5325));
    outputs(1860) <= layer6_outputs(982);
    outputs(1861) <= not(layer6_outputs(2161));
    outputs(1862) <= layer6_outputs(147);
    outputs(1863) <= not(layer6_outputs(3085));
    outputs(1864) <= not(layer6_outputs(5470));
    outputs(1865) <= (layer6_outputs(332)) xor (layer6_outputs(7589));
    outputs(1866) <= layer6_outputs(2481);
    outputs(1867) <= layer6_outputs(3506);
    outputs(1868) <= layer6_outputs(5632);
    outputs(1869) <= not(layer6_outputs(7087));
    outputs(1870) <= not((layer6_outputs(6829)) xor (layer6_outputs(2769)));
    outputs(1871) <= layer6_outputs(798);
    outputs(1872) <= (layer6_outputs(3399)) xor (layer6_outputs(5627));
    outputs(1873) <= (layer6_outputs(4)) xor (layer6_outputs(5170));
    outputs(1874) <= (layer6_outputs(5549)) and (layer6_outputs(3689));
    outputs(1875) <= layer6_outputs(4592);
    outputs(1876) <= layer6_outputs(1218);
    outputs(1877) <= layer6_outputs(3346);
    outputs(1878) <= (layer6_outputs(3970)) or (layer6_outputs(1080));
    outputs(1879) <= not(layer6_outputs(5100));
    outputs(1880) <= layer6_outputs(1219);
    outputs(1881) <= layer6_outputs(514);
    outputs(1882) <= not(layer6_outputs(48));
    outputs(1883) <= layer6_outputs(189);
    outputs(1884) <= layer6_outputs(7085);
    outputs(1885) <= not(layer6_outputs(4032));
    outputs(1886) <= layer6_outputs(7380);
    outputs(1887) <= (layer6_outputs(1869)) xor (layer6_outputs(1511));
    outputs(1888) <= not(layer6_outputs(5888));
    outputs(1889) <= layer6_outputs(6563);
    outputs(1890) <= not((layer6_outputs(5283)) xor (layer6_outputs(1600)));
    outputs(1891) <= not(layer6_outputs(4090));
    outputs(1892) <= (layer6_outputs(5894)) or (layer6_outputs(4340));
    outputs(1893) <= layer6_outputs(6698);
    outputs(1894) <= not(layer6_outputs(2873));
    outputs(1895) <= layer6_outputs(3993);
    outputs(1896) <= layer6_outputs(2083);
    outputs(1897) <= layer6_outputs(42);
    outputs(1898) <= layer6_outputs(3931);
    outputs(1899) <= layer6_outputs(1492);
    outputs(1900) <= not(layer6_outputs(4867));
    outputs(1901) <= not((layer6_outputs(1605)) xor (layer6_outputs(6565)));
    outputs(1902) <= not((layer6_outputs(7034)) xor (layer6_outputs(4753)));
    outputs(1903) <= layer6_outputs(7559);
    outputs(1904) <= layer6_outputs(5286);
    outputs(1905) <= not(layer6_outputs(1059));
    outputs(1906) <= not(layer6_outputs(1999));
    outputs(1907) <= not((layer6_outputs(1904)) and (layer6_outputs(2010)));
    outputs(1908) <= layer6_outputs(45);
    outputs(1909) <= not((layer6_outputs(2589)) xor (layer6_outputs(5391)));
    outputs(1910) <= (layer6_outputs(5988)) xor (layer6_outputs(80));
    outputs(1911) <= not((layer6_outputs(1258)) or (layer6_outputs(1302)));
    outputs(1912) <= layer6_outputs(5609);
    outputs(1913) <= layer6_outputs(3643);
    outputs(1914) <= layer6_outputs(927);
    outputs(1915) <= layer6_outputs(5243);
    outputs(1916) <= layer6_outputs(4805);
    outputs(1917) <= layer6_outputs(6118);
    outputs(1918) <= not(layer6_outputs(3354));
    outputs(1919) <= (layer6_outputs(588)) xor (layer6_outputs(1704));
    outputs(1920) <= not(layer6_outputs(5957));
    outputs(1921) <= (layer6_outputs(512)) and (layer6_outputs(4027));
    outputs(1922) <= not((layer6_outputs(4570)) xor (layer6_outputs(3667)));
    outputs(1923) <= layer6_outputs(1673);
    outputs(1924) <= layer6_outputs(6991);
    outputs(1925) <= not(layer6_outputs(5235)) or (layer6_outputs(289));
    outputs(1926) <= not(layer6_outputs(2411));
    outputs(1927) <= not(layer6_outputs(7509));
    outputs(1928) <= layer6_outputs(6564);
    outputs(1929) <= not(layer6_outputs(5169));
    outputs(1930) <= not(layer6_outputs(2792));
    outputs(1931) <= not((layer6_outputs(4269)) or (layer6_outputs(732)));
    outputs(1932) <= layer6_outputs(1903);
    outputs(1933) <= not(layer6_outputs(2063));
    outputs(1934) <= not(layer6_outputs(6841));
    outputs(1935) <= (layer6_outputs(2412)) xor (layer6_outputs(6136));
    outputs(1936) <= layer6_outputs(7159);
    outputs(1937) <= not(layer6_outputs(7413));
    outputs(1938) <= not(layer6_outputs(629));
    outputs(1939) <= not(layer6_outputs(3920));
    outputs(1940) <= layer6_outputs(6690);
    outputs(1941) <= layer6_outputs(202);
    outputs(1942) <= not((layer6_outputs(771)) xor (layer6_outputs(2487)));
    outputs(1943) <= not((layer6_outputs(7424)) and (layer6_outputs(4801)));
    outputs(1944) <= (layer6_outputs(2290)) and (layer6_outputs(4295));
    outputs(1945) <= not(layer6_outputs(6487));
    outputs(1946) <= not(layer6_outputs(7104));
    outputs(1947) <= layer6_outputs(1565);
    outputs(1948) <= (layer6_outputs(6754)) or (layer6_outputs(1048));
    outputs(1949) <= not(layer6_outputs(5724));
    outputs(1950) <= not(layer6_outputs(4695)) or (layer6_outputs(411));
    outputs(1951) <= not(layer6_outputs(2895));
    outputs(1952) <= not(layer6_outputs(5374));
    outputs(1953) <= layer6_outputs(5069);
    outputs(1954) <= layer6_outputs(4770);
    outputs(1955) <= not(layer6_outputs(1778));
    outputs(1956) <= not(layer6_outputs(6700));
    outputs(1957) <= (layer6_outputs(2364)) xor (layer6_outputs(1878));
    outputs(1958) <= (layer6_outputs(4810)) xor (layer6_outputs(4754));
    outputs(1959) <= layer6_outputs(2368);
    outputs(1960) <= (layer6_outputs(3991)) and not (layer6_outputs(5726));
    outputs(1961) <= (layer6_outputs(106)) and not (layer6_outputs(1630));
    outputs(1962) <= not(layer6_outputs(2003));
    outputs(1963) <= not(layer6_outputs(1611));
    outputs(1964) <= layer6_outputs(3253);
    outputs(1965) <= not((layer6_outputs(5020)) xor (layer6_outputs(4975)));
    outputs(1966) <= not(layer6_outputs(325));
    outputs(1967) <= layer6_outputs(5166);
    outputs(1968) <= not(layer6_outputs(7343));
    outputs(1969) <= not((layer6_outputs(4347)) xor (layer6_outputs(1314)));
    outputs(1970) <= (layer6_outputs(7090)) xor (layer6_outputs(2997));
    outputs(1971) <= not(layer6_outputs(2520));
    outputs(1972) <= not(layer6_outputs(975));
    outputs(1973) <= not((layer6_outputs(2810)) xor (layer6_outputs(2345)));
    outputs(1974) <= layer6_outputs(5680);
    outputs(1975) <= layer6_outputs(5973);
    outputs(1976) <= layer6_outputs(7596);
    outputs(1977) <= not(layer6_outputs(4123));
    outputs(1978) <= layer6_outputs(67);
    outputs(1979) <= not(layer6_outputs(5201));
    outputs(1980) <= not(layer6_outputs(324));
    outputs(1981) <= not(layer6_outputs(3600));
    outputs(1982) <= not(layer6_outputs(558));
    outputs(1983) <= not(layer6_outputs(4109));
    outputs(1984) <= (layer6_outputs(4608)) and not (layer6_outputs(2958));
    outputs(1985) <= not(layer6_outputs(1711));
    outputs(1986) <= not(layer6_outputs(2070));
    outputs(1987) <= not(layer6_outputs(3829));
    outputs(1988) <= not(layer6_outputs(536));
    outputs(1989) <= layer6_outputs(4455);
    outputs(1990) <= (layer6_outputs(5725)) and not (layer6_outputs(6471));
    outputs(1991) <= not(layer6_outputs(3507));
    outputs(1992) <= not(layer6_outputs(5953));
    outputs(1993) <= layer6_outputs(3108);
    outputs(1994) <= not(layer6_outputs(182));
    outputs(1995) <= not((layer6_outputs(5770)) or (layer6_outputs(169)));
    outputs(1996) <= not(layer6_outputs(6261));
    outputs(1997) <= (layer6_outputs(4355)) and not (layer6_outputs(6550));
    outputs(1998) <= layer6_outputs(4076);
    outputs(1999) <= (layer6_outputs(3939)) or (layer6_outputs(4888));
    outputs(2000) <= not((layer6_outputs(4809)) and (layer6_outputs(5457)));
    outputs(2001) <= (layer6_outputs(2277)) xor (layer6_outputs(6235));
    outputs(2002) <= not(layer6_outputs(7506));
    outputs(2003) <= not(layer6_outputs(2166));
    outputs(2004) <= layer6_outputs(4316);
    outputs(2005) <= not(layer6_outputs(5516));
    outputs(2006) <= layer6_outputs(476);
    outputs(2007) <= layer6_outputs(5534);
    outputs(2008) <= not(layer6_outputs(1811)) or (layer6_outputs(2462));
    outputs(2009) <= not((layer6_outputs(5771)) xor (layer6_outputs(4436)));
    outputs(2010) <= layer6_outputs(7143);
    outputs(2011) <= not((layer6_outputs(4878)) xor (layer6_outputs(4828)));
    outputs(2012) <= layer6_outputs(5591);
    outputs(2013) <= layer6_outputs(5687);
    outputs(2014) <= not(layer6_outputs(866));
    outputs(2015) <= not((layer6_outputs(4917)) xor (layer6_outputs(3980)));
    outputs(2016) <= layer6_outputs(2342);
    outputs(2017) <= (layer6_outputs(7114)) and (layer6_outputs(4487));
    outputs(2018) <= not((layer6_outputs(272)) or (layer6_outputs(3490)));
    outputs(2019) <= layer6_outputs(7559);
    outputs(2020) <= not(layer6_outputs(242));
    outputs(2021) <= not((layer6_outputs(6148)) xor (layer6_outputs(2446)));
    outputs(2022) <= not(layer6_outputs(5049));
    outputs(2023) <= not(layer6_outputs(4459));
    outputs(2024) <= not(layer6_outputs(5741)) or (layer6_outputs(7225));
    outputs(2025) <= not(layer6_outputs(5157));
    outputs(2026) <= layer6_outputs(2972);
    outputs(2027) <= layer6_outputs(1975);
    outputs(2028) <= layer6_outputs(3418);
    outputs(2029) <= not(layer6_outputs(7223));
    outputs(2030) <= layer6_outputs(6236);
    outputs(2031) <= not((layer6_outputs(5293)) or (layer6_outputs(6503)));
    outputs(2032) <= layer6_outputs(3067);
    outputs(2033) <= not(layer6_outputs(6334));
    outputs(2034) <= not(layer6_outputs(1110));
    outputs(2035) <= layer6_outputs(3123);
    outputs(2036) <= not(layer6_outputs(5727));
    outputs(2037) <= not((layer6_outputs(5575)) xor (layer6_outputs(5191)));
    outputs(2038) <= not(layer6_outputs(1553));
    outputs(2039) <= (layer6_outputs(2751)) xor (layer6_outputs(1688));
    outputs(2040) <= not((layer6_outputs(2365)) xor (layer6_outputs(5315)));
    outputs(2041) <= not((layer6_outputs(5656)) xor (layer6_outputs(4576)));
    outputs(2042) <= not(layer6_outputs(2174));
    outputs(2043) <= not(layer6_outputs(5673)) or (layer6_outputs(1039));
    outputs(2044) <= layer6_outputs(3394);
    outputs(2045) <= layer6_outputs(1104);
    outputs(2046) <= not(layer6_outputs(2440));
    outputs(2047) <= not(layer6_outputs(2996));
    outputs(2048) <= layer6_outputs(296);
    outputs(2049) <= (layer6_outputs(2550)) and not (layer6_outputs(3415));
    outputs(2050) <= not(layer6_outputs(6732));
    outputs(2051) <= not(layer6_outputs(7193));
    outputs(2052) <= not(layer6_outputs(3750));
    outputs(2053) <= (layer6_outputs(4071)) xor (layer6_outputs(6296));
    outputs(2054) <= not((layer6_outputs(4308)) xor (layer6_outputs(4796)));
    outputs(2055) <= layer6_outputs(5973);
    outputs(2056) <= not(layer6_outputs(7149));
    outputs(2057) <= layer6_outputs(2170);
    outputs(2058) <= not(layer6_outputs(4676));
    outputs(2059) <= not(layer6_outputs(3035));
    outputs(2060) <= layer6_outputs(4748);
    outputs(2061) <= not((layer6_outputs(6053)) xor (layer6_outputs(4592)));
    outputs(2062) <= not((layer6_outputs(5546)) xor (layer6_outputs(5681)));
    outputs(2063) <= not(layer6_outputs(5421));
    outputs(2064) <= layer6_outputs(1726);
    outputs(2065) <= (layer6_outputs(1763)) and not (layer6_outputs(39));
    outputs(2066) <= not(layer6_outputs(1046));
    outputs(2067) <= not(layer6_outputs(1367));
    outputs(2068) <= layer6_outputs(5305);
    outputs(2069) <= (layer6_outputs(782)) xor (layer6_outputs(2905));
    outputs(2070) <= not(layer6_outputs(2161));
    outputs(2071) <= (layer6_outputs(3743)) xor (layer6_outputs(6460));
    outputs(2072) <= not(layer6_outputs(7619));
    outputs(2073) <= not(layer6_outputs(4427));
    outputs(2074) <= not((layer6_outputs(1047)) xor (layer6_outputs(3933)));
    outputs(2075) <= not(layer6_outputs(7469));
    outputs(2076) <= not(layer6_outputs(7041));
    outputs(2077) <= layer6_outputs(6420);
    outputs(2078) <= (layer6_outputs(5267)) xor (layer6_outputs(3167));
    outputs(2079) <= not(layer6_outputs(761));
    outputs(2080) <= layer6_outputs(4747);
    outputs(2081) <= not(layer6_outputs(4044));
    outputs(2082) <= not(layer6_outputs(2558)) or (layer6_outputs(2155));
    outputs(2083) <= not((layer6_outputs(3482)) xor (layer6_outputs(1736)));
    outputs(2084) <= (layer6_outputs(5745)) and not (layer6_outputs(7070));
    outputs(2085) <= (layer6_outputs(6577)) and (layer6_outputs(6615));
    outputs(2086) <= (layer6_outputs(3687)) xor (layer6_outputs(4663));
    outputs(2087) <= (layer6_outputs(7447)) and (layer6_outputs(6807));
    outputs(2088) <= not(layer6_outputs(183));
    outputs(2089) <= layer6_outputs(5177);
    outputs(2090) <= not(layer6_outputs(7011));
    outputs(2091) <= not(layer6_outputs(2499));
    outputs(2092) <= not((layer6_outputs(4822)) xor (layer6_outputs(6318)));
    outputs(2093) <= not(layer6_outputs(1455));
    outputs(2094) <= (layer6_outputs(3760)) xor (layer6_outputs(4815));
    outputs(2095) <= layer6_outputs(902);
    outputs(2096) <= not(layer6_outputs(6170));
    outputs(2097) <= layer6_outputs(2331);
    outputs(2098) <= not((layer6_outputs(6914)) xor (layer6_outputs(2405)));
    outputs(2099) <= not(layer6_outputs(7126));
    outputs(2100) <= not(layer6_outputs(5993));
    outputs(2101) <= not(layer6_outputs(2669));
    outputs(2102) <= not((layer6_outputs(5711)) xor (layer6_outputs(6861)));
    outputs(2103) <= not(layer6_outputs(2861));
    outputs(2104) <= not(layer6_outputs(1092));
    outputs(2105) <= (layer6_outputs(2416)) and not (layer6_outputs(1423));
    outputs(2106) <= layer6_outputs(7000);
    outputs(2107) <= not(layer6_outputs(2478));
    outputs(2108) <= not(layer6_outputs(3751)) or (layer6_outputs(5764));
    outputs(2109) <= not((layer6_outputs(321)) xor (layer6_outputs(1122)));
    outputs(2110) <= layer6_outputs(2457);
    outputs(2111) <= not(layer6_outputs(199));
    outputs(2112) <= not(layer6_outputs(5167)) or (layer6_outputs(3510));
    outputs(2113) <= layer6_outputs(451);
    outputs(2114) <= not(layer6_outputs(5507));
    outputs(2115) <= not(layer6_outputs(857));
    outputs(2116) <= layer6_outputs(7301);
    outputs(2117) <= (layer6_outputs(4215)) and (layer6_outputs(290));
    outputs(2118) <= not(layer6_outputs(797));
    outputs(2119) <= not(layer6_outputs(1982));
    outputs(2120) <= not((layer6_outputs(2400)) xor (layer6_outputs(693)));
    outputs(2121) <= not((layer6_outputs(5879)) and (layer6_outputs(2629)));
    outputs(2122) <= not((layer6_outputs(4852)) xor (layer6_outputs(2575)));
    outputs(2123) <= layer6_outputs(7586);
    outputs(2124) <= layer6_outputs(3006);
    outputs(2125) <= layer6_outputs(1424);
    outputs(2126) <= not(layer6_outputs(4571));
    outputs(2127) <= layer6_outputs(2803);
    outputs(2128) <= not((layer6_outputs(105)) or (layer6_outputs(1612)));
    outputs(2129) <= layer6_outputs(6233);
    outputs(2130) <= not(layer6_outputs(3566));
    outputs(2131) <= not(layer6_outputs(408));
    outputs(2132) <= layer6_outputs(79);
    outputs(2133) <= not(layer6_outputs(1056)) or (layer6_outputs(2167));
    outputs(2134) <= not(layer6_outputs(3692));
    outputs(2135) <= not(layer6_outputs(2310));
    outputs(2136) <= not(layer6_outputs(281));
    outputs(2137) <= not(layer6_outputs(626));
    outputs(2138) <= not(layer6_outputs(5292)) or (layer6_outputs(2562));
    outputs(2139) <= not((layer6_outputs(5456)) xor (layer6_outputs(4875)));
    outputs(2140) <= not(layer6_outputs(5948));
    outputs(2141) <= layer6_outputs(6459);
    outputs(2142) <= (layer6_outputs(5261)) xor (layer6_outputs(1592));
    outputs(2143) <= not(layer6_outputs(2652));
    outputs(2144) <= layer6_outputs(6023);
    outputs(2145) <= not(layer6_outputs(1077));
    outputs(2146) <= not((layer6_outputs(7405)) xor (layer6_outputs(3390)));
    outputs(2147) <= not(layer6_outputs(193));
    outputs(2148) <= (layer6_outputs(5758)) and not (layer6_outputs(969));
    outputs(2149) <= not(layer6_outputs(1238));
    outputs(2150) <= not(layer6_outputs(6037));
    outputs(2151) <= not((layer6_outputs(1832)) and (layer6_outputs(6707)));
    outputs(2152) <= not(layer6_outputs(2398));
    outputs(2153) <= layer6_outputs(5716);
    outputs(2154) <= layer6_outputs(5363);
    outputs(2155) <= not(layer6_outputs(1385));
    outputs(2156) <= not(layer6_outputs(3330));
    outputs(2157) <= layer6_outputs(18);
    outputs(2158) <= (layer6_outputs(4930)) xor (layer6_outputs(4346));
    outputs(2159) <= not((layer6_outputs(4274)) xor (layer6_outputs(5867)));
    outputs(2160) <= not(layer6_outputs(224));
    outputs(2161) <= not(layer6_outputs(4607));
    outputs(2162) <= not(layer6_outputs(7102));
    outputs(2163) <= not((layer6_outputs(2571)) and (layer6_outputs(2627)));
    outputs(2164) <= not(layer6_outputs(7144));
    outputs(2165) <= not(layer6_outputs(2009));
    outputs(2166) <= layer6_outputs(6526);
    outputs(2167) <= '0';
    outputs(2168) <= not(layer6_outputs(2470));
    outputs(2169) <= layer6_outputs(6390);
    outputs(2170) <= (layer6_outputs(2553)) and (layer6_outputs(6437));
    outputs(2171) <= not(layer6_outputs(2192));
    outputs(2172) <= not(layer6_outputs(4208));
    outputs(2173) <= not((layer6_outputs(931)) xor (layer6_outputs(7028)));
    outputs(2174) <= not((layer6_outputs(3035)) xor (layer6_outputs(4465)));
    outputs(2175) <= layer6_outputs(1569);
    outputs(2176) <= (layer6_outputs(7026)) and (layer6_outputs(5754));
    outputs(2177) <= not(layer6_outputs(1615));
    outputs(2178) <= layer6_outputs(4124);
    outputs(2179) <= layer6_outputs(3425);
    outputs(2180) <= layer6_outputs(5342);
    outputs(2181) <= (layer6_outputs(2579)) and not (layer6_outputs(1102));
    outputs(2182) <= layer6_outputs(4836);
    outputs(2183) <= not(layer6_outputs(3620));
    outputs(2184) <= (layer6_outputs(6530)) xor (layer6_outputs(4094));
    outputs(2185) <= (layer6_outputs(1050)) xor (layer6_outputs(4566));
    outputs(2186) <= layer6_outputs(2953);
    outputs(2187) <= not(layer6_outputs(1302));
    outputs(2188) <= layer6_outputs(963);
    outputs(2189) <= layer6_outputs(4328);
    outputs(2190) <= layer6_outputs(5348);
    outputs(2191) <= not(layer6_outputs(2017));
    outputs(2192) <= not((layer6_outputs(4428)) xor (layer6_outputs(5092)));
    outputs(2193) <= layer6_outputs(2737);
    outputs(2194) <= not((layer6_outputs(4097)) xor (layer6_outputs(4177)));
    outputs(2195) <= (layer6_outputs(7554)) and not (layer6_outputs(2862));
    outputs(2196) <= not(layer6_outputs(6475));
    outputs(2197) <= not(layer6_outputs(6054)) or (layer6_outputs(1289));
    outputs(2198) <= not(layer6_outputs(7633));
    outputs(2199) <= layer6_outputs(5269);
    outputs(2200) <= not((layer6_outputs(6627)) xor (layer6_outputs(6971)));
    outputs(2201) <= not(layer6_outputs(4468));
    outputs(2202) <= not(layer6_outputs(5093));
    outputs(2203) <= not((layer6_outputs(462)) xor (layer6_outputs(2406)));
    outputs(2204) <= not(layer6_outputs(6902));
    outputs(2205) <= (layer6_outputs(7555)) and not (layer6_outputs(3581));
    outputs(2206) <= layer6_outputs(6490);
    outputs(2207) <= layer6_outputs(3466);
    outputs(2208) <= layer6_outputs(265);
    outputs(2209) <= layer6_outputs(3164);
    outputs(2210) <= (layer6_outputs(3730)) and not (layer6_outputs(3438));
    outputs(2211) <= layer6_outputs(6021);
    outputs(2212) <= not(layer6_outputs(2703));
    outputs(2213) <= (layer6_outputs(6583)) xor (layer6_outputs(3246));
    outputs(2214) <= layer6_outputs(4546);
    outputs(2215) <= layer6_outputs(4413);
    outputs(2216) <= not((layer6_outputs(7023)) xor (layer6_outputs(4556)));
    outputs(2217) <= not(layer6_outputs(6946));
    outputs(2218) <= layer6_outputs(476);
    outputs(2219) <= (layer6_outputs(6726)) and not (layer6_outputs(3660));
    outputs(2220) <= layer6_outputs(4341);
    outputs(2221) <= (layer6_outputs(3569)) xor (layer6_outputs(116));
    outputs(2222) <= layer6_outputs(735);
    outputs(2223) <= layer6_outputs(3312);
    outputs(2224) <= (layer6_outputs(5455)) xor (layer6_outputs(6750));
    outputs(2225) <= not((layer6_outputs(5314)) xor (layer6_outputs(6328)));
    outputs(2226) <= layer6_outputs(2356);
    outputs(2227) <= (layer6_outputs(6877)) and not (layer6_outputs(1086));
    outputs(2228) <= layer6_outputs(3195);
    outputs(2229) <= (layer6_outputs(4276)) xor (layer6_outputs(1709));
    outputs(2230) <= not(layer6_outputs(6613));
    outputs(2231) <= layer6_outputs(6191);
    outputs(2232) <= not((layer6_outputs(4225)) xor (layer6_outputs(3133)));
    outputs(2233) <= layer6_outputs(1927);
    outputs(2234) <= not(layer6_outputs(5744));
    outputs(2235) <= (layer6_outputs(6871)) xor (layer6_outputs(6806));
    outputs(2236) <= layer6_outputs(1739);
    outputs(2237) <= (layer6_outputs(3421)) and not (layer6_outputs(4412));
    outputs(2238) <= not(layer6_outputs(1659));
    outputs(2239) <= not(layer6_outputs(2414));
    outputs(2240) <= layer6_outputs(4041);
    outputs(2241) <= layer6_outputs(3634);
    outputs(2242) <= layer6_outputs(1762);
    outputs(2243) <= layer6_outputs(4963);
    outputs(2244) <= layer6_outputs(5508);
    outputs(2245) <= layer6_outputs(6491);
    outputs(2246) <= not(layer6_outputs(6402));
    outputs(2247) <= layer6_outputs(1036);
    outputs(2248) <= layer6_outputs(6274);
    outputs(2249) <= layer6_outputs(6021);
    outputs(2250) <= not(layer6_outputs(1323));
    outputs(2251) <= layer6_outputs(3846);
    outputs(2252) <= (layer6_outputs(5874)) xor (layer6_outputs(611));
    outputs(2253) <= layer6_outputs(3776);
    outputs(2254) <= not(layer6_outputs(7046));
    outputs(2255) <= layer6_outputs(720);
    outputs(2256) <= not(layer6_outputs(2367));
    outputs(2257) <= not((layer6_outputs(3403)) xor (layer6_outputs(6177)));
    outputs(2258) <= layer6_outputs(4549);
    outputs(2259) <= layer6_outputs(5339);
    outputs(2260) <= not((layer6_outputs(6704)) xor (layer6_outputs(3696)));
    outputs(2261) <= layer6_outputs(1378);
    outputs(2262) <= not(layer6_outputs(3327));
    outputs(2263) <= layer6_outputs(6137);
    outputs(2264) <= not(layer6_outputs(2235));
    outputs(2265) <= not(layer6_outputs(504));
    outputs(2266) <= layer6_outputs(3784);
    outputs(2267) <= not(layer6_outputs(3147));
    outputs(2268) <= not((layer6_outputs(3254)) xor (layer6_outputs(1706)));
    outputs(2269) <= layer6_outputs(1146);
    outputs(2270) <= not((layer6_outputs(1987)) and (layer6_outputs(4203)));
    outputs(2271) <= not(layer6_outputs(527));
    outputs(2272) <= not(layer6_outputs(1670));
    outputs(2273) <= not(layer6_outputs(2813));
    outputs(2274) <= not(layer6_outputs(253));
    outputs(2275) <= layer6_outputs(1598);
    outputs(2276) <= not(layer6_outputs(2836));
    outputs(2277) <= (layer6_outputs(7304)) xor (layer6_outputs(7038));
    outputs(2278) <= not(layer6_outputs(2585));
    outputs(2279) <= not(layer6_outputs(3739));
    outputs(2280) <= layer6_outputs(6442);
    outputs(2281) <= not(layer6_outputs(6380));
    outputs(2282) <= layer6_outputs(2758);
    outputs(2283) <= not(layer6_outputs(7211));
    outputs(2284) <= not(layer6_outputs(214));
    outputs(2285) <= layer6_outputs(6807);
    outputs(2286) <= not(layer6_outputs(4558));
    outputs(2287) <= not((layer6_outputs(1873)) xor (layer6_outputs(2486)));
    outputs(2288) <= not(layer6_outputs(604));
    outputs(2289) <= layer6_outputs(2257);
    outputs(2290) <= (layer6_outputs(6893)) xor (layer6_outputs(1964));
    outputs(2291) <= not(layer6_outputs(2763));
    outputs(2292) <= layer6_outputs(2347);
    outputs(2293) <= layer6_outputs(2968);
    outputs(2294) <= not(layer6_outputs(1389));
    outputs(2295) <= (layer6_outputs(6737)) and not (layer6_outputs(959));
    outputs(2296) <= not((layer6_outputs(4829)) xor (layer6_outputs(342)));
    outputs(2297) <= not(layer6_outputs(4764));
    outputs(2298) <= layer6_outputs(1657);
    outputs(2299) <= layer6_outputs(4670);
    outputs(2300) <= not((layer6_outputs(2463)) or (layer6_outputs(3335)));
    outputs(2301) <= not(layer6_outputs(1819));
    outputs(2302) <= layer6_outputs(2110);
    outputs(2303) <= layer6_outputs(6984);
    outputs(2304) <= layer6_outputs(2854);
    outputs(2305) <= not((layer6_outputs(6716)) xor (layer6_outputs(4786)));
    outputs(2306) <= not(layer6_outputs(1161));
    outputs(2307) <= layer6_outputs(3649);
    outputs(2308) <= (layer6_outputs(243)) and (layer6_outputs(987));
    outputs(2309) <= layer6_outputs(1177);
    outputs(2310) <= not((layer6_outputs(5643)) xor (layer6_outputs(1436)));
    outputs(2311) <= (layer6_outputs(2021)) and not (layer6_outputs(4387));
    outputs(2312) <= (layer6_outputs(1754)) xor (layer6_outputs(134));
    outputs(2313) <= layer6_outputs(5329);
    outputs(2314) <= layer6_outputs(5502);
    outputs(2315) <= layer6_outputs(7171);
    outputs(2316) <= not((layer6_outputs(5096)) xor (layer6_outputs(690)));
    outputs(2317) <= not(layer6_outputs(5137));
    outputs(2318) <= (layer6_outputs(6640)) and not (layer6_outputs(4569));
    outputs(2319) <= (layer6_outputs(1151)) xor (layer6_outputs(7351));
    outputs(2320) <= layer6_outputs(1341);
    outputs(2321) <= layer6_outputs(4397);
    outputs(2322) <= not((layer6_outputs(1368)) xor (layer6_outputs(1184)));
    outputs(2323) <= (layer6_outputs(4369)) or (layer6_outputs(6045));
    outputs(2324) <= not((layer6_outputs(3742)) xor (layer6_outputs(6295)));
    outputs(2325) <= not(layer6_outputs(4590));
    outputs(2326) <= layer6_outputs(253);
    outputs(2327) <= layer6_outputs(1888);
    outputs(2328) <= not(layer6_outputs(4001));
    outputs(2329) <= not(layer6_outputs(5488)) or (layer6_outputs(5023));
    outputs(2330) <= not((layer6_outputs(5505)) xor (layer6_outputs(3132)));
    outputs(2331) <= layer6_outputs(2628);
    outputs(2332) <= layer6_outputs(3007);
    outputs(2333) <= not(layer6_outputs(7434));
    outputs(2334) <= layer6_outputs(4305);
    outputs(2335) <= (layer6_outputs(2337)) and not (layer6_outputs(5437));
    outputs(2336) <= not(layer6_outputs(6826));
    outputs(2337) <= not((layer6_outputs(6574)) and (layer6_outputs(5995)));
    outputs(2338) <= not(layer6_outputs(354));
    outputs(2339) <= not(layer6_outputs(6771));
    outputs(2340) <= (layer6_outputs(5373)) xor (layer6_outputs(7025));
    outputs(2341) <= layer6_outputs(1600);
    outputs(2342) <= not(layer6_outputs(361));
    outputs(2343) <= layer6_outputs(3071);
    outputs(2344) <= not(layer6_outputs(3829));
    outputs(2345) <= layer6_outputs(5397);
    outputs(2346) <= not(layer6_outputs(2116));
    outputs(2347) <= not(layer6_outputs(7180));
    outputs(2348) <= (layer6_outputs(4718)) and (layer6_outputs(7034));
    outputs(2349) <= layer6_outputs(3489);
    outputs(2350) <= layer6_outputs(3123);
    outputs(2351) <= layer6_outputs(88);
    outputs(2352) <= (layer6_outputs(6447)) and not (layer6_outputs(5739));
    outputs(2353) <= not((layer6_outputs(5620)) or (layer6_outputs(459)));
    outputs(2354) <= not(layer6_outputs(2229)) or (layer6_outputs(7113));
    outputs(2355) <= not(layer6_outputs(485));
    outputs(2356) <= not(layer6_outputs(6204));
    outputs(2357) <= (layer6_outputs(4973)) xor (layer6_outputs(1989));
    outputs(2358) <= not(layer6_outputs(3457));
    outputs(2359) <= not(layer6_outputs(4713));
    outputs(2360) <= not((layer6_outputs(7318)) xor (layer6_outputs(237)));
    outputs(2361) <= (layer6_outputs(6592)) and not (layer6_outputs(6410));
    outputs(2362) <= not((layer6_outputs(62)) or (layer6_outputs(4756)));
    outputs(2363) <= (layer6_outputs(3630)) xor (layer6_outputs(4751));
    outputs(2364) <= layer6_outputs(4401);
    outputs(2365) <= not((layer6_outputs(1435)) or (layer6_outputs(360)));
    outputs(2366) <= not((layer6_outputs(4666)) and (layer6_outputs(1778)));
    outputs(2367) <= (layer6_outputs(19)) xor (layer6_outputs(2119));
    outputs(2368) <= layer6_outputs(3533);
    outputs(2369) <= (layer6_outputs(6431)) and not (layer6_outputs(6948));
    outputs(2370) <= layer6_outputs(1773);
    outputs(2371) <= not(layer6_outputs(7548));
    outputs(2372) <= not(layer6_outputs(5598));
    outputs(2373) <= not(layer6_outputs(324));
    outputs(2374) <= not(layer6_outputs(441));
    outputs(2375) <= layer6_outputs(7079);
    outputs(2376) <= layer6_outputs(4871);
    outputs(2377) <= not(layer6_outputs(3639));
    outputs(2378) <= layer6_outputs(7237);
    outputs(2379) <= (layer6_outputs(4167)) and (layer6_outputs(2909));
    outputs(2380) <= layer6_outputs(232);
    outputs(2381) <= not(layer6_outputs(2190));
    outputs(2382) <= not(layer6_outputs(3389));
    outputs(2383) <= layer6_outputs(2710);
    outputs(2384) <= (layer6_outputs(6599)) or (layer6_outputs(5722));
    outputs(2385) <= (layer6_outputs(4925)) xor (layer6_outputs(3275));
    outputs(2386) <= layer6_outputs(2261);
    outputs(2387) <= not((layer6_outputs(2490)) xor (layer6_outputs(4278)));
    outputs(2388) <= (layer6_outputs(4232)) xor (layer6_outputs(7642));
    outputs(2389) <= (layer6_outputs(676)) and not (layer6_outputs(2134));
    outputs(2390) <= layer6_outputs(4076);
    outputs(2391) <= layer6_outputs(4731);
    outputs(2392) <= layer6_outputs(1813);
    outputs(2393) <= (layer6_outputs(6191)) and not (layer6_outputs(5343));
    outputs(2394) <= not(layer6_outputs(3442));
    outputs(2395) <= not(layer6_outputs(7567));
    outputs(2396) <= not(layer6_outputs(2374));
    outputs(2397) <= (layer6_outputs(2563)) and (layer6_outputs(1885));
    outputs(2398) <= not(layer6_outputs(5194));
    outputs(2399) <= not((layer6_outputs(7423)) or (layer6_outputs(864)));
    outputs(2400) <= not(layer6_outputs(7629));
    outputs(2401) <= not((layer6_outputs(6637)) xor (layer6_outputs(1628)));
    outputs(2402) <= (layer6_outputs(1343)) xor (layer6_outputs(1389));
    outputs(2403) <= (layer6_outputs(424)) and not (layer6_outputs(3503));
    outputs(2404) <= (layer6_outputs(7254)) and (layer6_outputs(6775));
    outputs(2405) <= (layer6_outputs(5001)) and not (layer6_outputs(5812));
    outputs(2406) <= not(layer6_outputs(5352));
    outputs(2407) <= (layer6_outputs(2831)) xor (layer6_outputs(6746));
    outputs(2408) <= not(layer6_outputs(1664));
    outputs(2409) <= not(layer6_outputs(1876));
    outputs(2410) <= layer6_outputs(6201);
    outputs(2411) <= not((layer6_outputs(2034)) xor (layer6_outputs(6451)));
    outputs(2412) <= layer6_outputs(5881);
    outputs(2413) <= (layer6_outputs(5662)) and not (layer6_outputs(5675));
    outputs(2414) <= not(layer6_outputs(2129));
    outputs(2415) <= layer6_outputs(1382);
    outputs(2416) <= (layer6_outputs(5418)) and not (layer6_outputs(6472));
    outputs(2417) <= not((layer6_outputs(383)) xor (layer6_outputs(3500)));
    outputs(2418) <= not(layer6_outputs(170));
    outputs(2419) <= layer6_outputs(2370);
    outputs(2420) <= (layer6_outputs(6952)) xor (layer6_outputs(5219));
    outputs(2421) <= not(layer6_outputs(7184));
    outputs(2422) <= not((layer6_outputs(7453)) xor (layer6_outputs(2618)));
    outputs(2423) <= (layer6_outputs(7562)) and not (layer6_outputs(6684));
    outputs(2424) <= not(layer6_outputs(2952));
    outputs(2425) <= layer6_outputs(2972);
    outputs(2426) <= not((layer6_outputs(2653)) xor (layer6_outputs(1208)));
    outputs(2427) <= layer6_outputs(1052);
    outputs(2428) <= not((layer6_outputs(4680)) or (layer6_outputs(3202)));
    outputs(2429) <= layer6_outputs(1465);
    outputs(2430) <= layer6_outputs(3453);
    outputs(2431) <= layer6_outputs(2928);
    outputs(2432) <= (layer6_outputs(6547)) and (layer6_outputs(4149));
    outputs(2433) <= (layer6_outputs(6670)) and not (layer6_outputs(6647));
    outputs(2434) <= (layer6_outputs(1072)) xor (layer6_outputs(4986));
    outputs(2435) <= layer6_outputs(4349);
    outputs(2436) <= layer6_outputs(2249);
    outputs(2437) <= (layer6_outputs(3667)) xor (layer6_outputs(2664));
    outputs(2438) <= (layer6_outputs(2652)) xor (layer6_outputs(2612));
    outputs(2439) <= (layer6_outputs(2845)) and not (layer6_outputs(4021));
    outputs(2440) <= not(layer6_outputs(4157));
    outputs(2441) <= layer6_outputs(4066);
    outputs(2442) <= not(layer6_outputs(4847));
    outputs(2443) <= layer6_outputs(1049);
    outputs(2444) <= not(layer6_outputs(358));
    outputs(2445) <= layer6_outputs(4079);
    outputs(2446) <= (layer6_outputs(3579)) and (layer6_outputs(5680));
    outputs(2447) <= not(layer6_outputs(1065));
    outputs(2448) <= not((layer6_outputs(1246)) xor (layer6_outputs(1515)));
    outputs(2449) <= not(layer6_outputs(3984));
    outputs(2450) <= not(layer6_outputs(2474)) or (layer6_outputs(5703));
    outputs(2451) <= not(layer6_outputs(1501));
    outputs(2452) <= not(layer6_outputs(4788));
    outputs(2453) <= layer6_outputs(6080);
    outputs(2454) <= layer6_outputs(3853);
    outputs(2455) <= not(layer6_outputs(2127)) or (layer6_outputs(7137));
    outputs(2456) <= not((layer6_outputs(2207)) xor (layer6_outputs(6480)));
    outputs(2457) <= layer6_outputs(2109);
    outputs(2458) <= not((layer6_outputs(6111)) and (layer6_outputs(2167)));
    outputs(2459) <= not(layer6_outputs(5901));
    outputs(2460) <= not(layer6_outputs(6482));
    outputs(2461) <= (layer6_outputs(532)) xor (layer6_outputs(638));
    outputs(2462) <= not(layer6_outputs(5612));
    outputs(2463) <= not(layer6_outputs(6093));
    outputs(2464) <= not(layer6_outputs(3144));
    outputs(2465) <= (layer6_outputs(812)) and (layer6_outputs(3662));
    outputs(2466) <= not(layer6_outputs(2130));
    outputs(2467) <= not(layer6_outputs(1459));
    outputs(2468) <= not(layer6_outputs(451)) or (layer6_outputs(7422));
    outputs(2469) <= layer6_outputs(5238);
    outputs(2470) <= layer6_outputs(5553);
    outputs(2471) <= layer6_outputs(762);
    outputs(2472) <= not(layer6_outputs(2461));
    outputs(2473) <= layer6_outputs(4699);
    outputs(2474) <= not((layer6_outputs(3793)) or (layer6_outputs(1280)));
    outputs(2475) <= not((layer6_outputs(227)) and (layer6_outputs(3610)));
    outputs(2476) <= not(layer6_outputs(421));
    outputs(2477) <= layer6_outputs(2548);
    outputs(2478) <= (layer6_outputs(7290)) and (layer6_outputs(4707));
    outputs(2479) <= not(layer6_outputs(654));
    outputs(2480) <= not(layer6_outputs(2615));
    outputs(2481) <= layer6_outputs(7615);
    outputs(2482) <= not(layer6_outputs(5791));
    outputs(2483) <= layer6_outputs(3395);
    outputs(2484) <= not(layer6_outputs(1235));
    outputs(2485) <= not(layer6_outputs(1857));
    outputs(2486) <= not((layer6_outputs(62)) or (layer6_outputs(6834)));
    outputs(2487) <= not((layer6_outputs(5746)) xor (layer6_outputs(5656)));
    outputs(2488) <= layer6_outputs(733);
    outputs(2489) <= (layer6_outputs(4047)) and not (layer6_outputs(624));
    outputs(2490) <= layer6_outputs(4073);
    outputs(2491) <= not(layer6_outputs(142));
    outputs(2492) <= not(layer6_outputs(2380));
    outputs(2493) <= not(layer6_outputs(6474)) or (layer6_outputs(6428));
    outputs(2494) <= not((layer6_outputs(2378)) xor (layer6_outputs(5463)));
    outputs(2495) <= layer6_outputs(4533);
    outputs(2496) <= not((layer6_outputs(5713)) or (layer6_outputs(4141)));
    outputs(2497) <= not((layer6_outputs(649)) or (layer6_outputs(2574)));
    outputs(2498) <= not(layer6_outputs(3919));
    outputs(2499) <= (layer6_outputs(6529)) xor (layer6_outputs(725));
    outputs(2500) <= layer6_outputs(7319);
    outputs(2501) <= layer6_outputs(4434);
    outputs(2502) <= not((layer6_outputs(1361)) or (layer6_outputs(6055)));
    outputs(2503) <= not(layer6_outputs(1927));
    outputs(2504) <= not(layer6_outputs(5072));
    outputs(2505) <= layer6_outputs(3415);
    outputs(2506) <= (layer6_outputs(879)) and not (layer6_outputs(6585));
    outputs(2507) <= (layer6_outputs(759)) and not (layer6_outputs(6757));
    outputs(2508) <= not(layer6_outputs(1225)) or (layer6_outputs(3352));
    outputs(2509) <= not(layer6_outputs(3442));
    outputs(2510) <= layer6_outputs(2877);
    outputs(2511) <= layer6_outputs(1023);
    outputs(2512) <= not(layer6_outputs(4727));
    outputs(2513) <= not(layer6_outputs(6835));
    outputs(2514) <= (layer6_outputs(6676)) and (layer6_outputs(2613));
    outputs(2515) <= not(layer6_outputs(1089));
    outputs(2516) <= layer6_outputs(4456);
    outputs(2517) <= not((layer6_outputs(1384)) xor (layer6_outputs(3261)));
    outputs(2518) <= not(layer6_outputs(1179));
    outputs(2519) <= not((layer6_outputs(7236)) or (layer6_outputs(518)));
    outputs(2520) <= layer6_outputs(4997);
    outputs(2521) <= layer6_outputs(1061);
    outputs(2522) <= layer6_outputs(3084);
    outputs(2523) <= layer6_outputs(3023);
    outputs(2524) <= not(layer6_outputs(5877));
    outputs(2525) <= not(layer6_outputs(4777)) or (layer6_outputs(1931));
    outputs(2526) <= layer6_outputs(1193);
    outputs(2527) <= not(layer6_outputs(5148));
    outputs(2528) <= (layer6_outputs(7081)) xor (layer6_outputs(3214));
    outputs(2529) <= (layer6_outputs(1638)) and not (layer6_outputs(7365));
    outputs(2530) <= layer6_outputs(6872);
    outputs(2531) <= not(layer6_outputs(7287));
    outputs(2532) <= not(layer6_outputs(6444));
    outputs(2533) <= not(layer6_outputs(3255));
    outputs(2534) <= not(layer6_outputs(1628));
    outputs(2535) <= not(layer6_outputs(3235));
    outputs(2536) <= layer6_outputs(7346);
    outputs(2537) <= not(layer6_outputs(6520));
    outputs(2538) <= (layer6_outputs(1173)) and (layer6_outputs(3635));
    outputs(2539) <= layer6_outputs(6128);
    outputs(2540) <= not(layer6_outputs(6411));
    outputs(2541) <= not(layer6_outputs(1827));
    outputs(2542) <= (layer6_outputs(880)) xor (layer6_outputs(78));
    outputs(2543) <= '0';
    outputs(2544) <= (layer6_outputs(2448)) and not (layer6_outputs(7056));
    outputs(2545) <= not(layer6_outputs(3553)) or (layer6_outputs(3818));
    outputs(2546) <= (layer6_outputs(5465)) and (layer6_outputs(1998));
    outputs(2547) <= not((layer6_outputs(4398)) xor (layer6_outputs(1279)));
    outputs(2548) <= not((layer6_outputs(392)) xor (layer6_outputs(4635)));
    outputs(2549) <= layer6_outputs(3143);
    outputs(2550) <= not(layer6_outputs(4620));
    outputs(2551) <= (layer6_outputs(6779)) or (layer6_outputs(1691));
    outputs(2552) <= (layer6_outputs(4870)) and not (layer6_outputs(5611));
    outputs(2553) <= layer6_outputs(1432);
    outputs(2554) <= layer6_outputs(278);
    outputs(2555) <= layer6_outputs(7649);
    outputs(2556) <= not(layer6_outputs(6760));
    outputs(2557) <= layer6_outputs(4236);
    outputs(2558) <= layer6_outputs(6497);
    outputs(2559) <= (layer6_outputs(84)) and (layer6_outputs(5040));
    outputs(2560) <= layer6_outputs(6566);
    outputs(2561) <= layer6_outputs(1613);
    outputs(2562) <= not(layer6_outputs(3470));
    outputs(2563) <= layer6_outputs(6052);
    outputs(2564) <= not(layer6_outputs(6102));
    outputs(2565) <= not((layer6_outputs(632)) xor (layer6_outputs(6450)));
    outputs(2566) <= not(layer6_outputs(2333));
    outputs(2567) <= layer6_outputs(6369);
    outputs(2568) <= (layer6_outputs(5359)) or (layer6_outputs(1237));
    outputs(2569) <= not(layer6_outputs(7580));
    outputs(2570) <= not((layer6_outputs(515)) xor (layer6_outputs(2121)));
    outputs(2571) <= (layer6_outputs(5332)) and (layer6_outputs(5922));
    outputs(2572) <= not((layer6_outputs(6515)) or (layer6_outputs(6093)));
    outputs(2573) <= not(layer6_outputs(1441));
    outputs(2574) <= (layer6_outputs(7561)) xor (layer6_outputs(3753));
    outputs(2575) <= (layer6_outputs(7677)) and not (layer6_outputs(5036));
    outputs(2576) <= not(layer6_outputs(6631));
    outputs(2577) <= layer6_outputs(3951);
    outputs(2578) <= not(layer6_outputs(7490));
    outputs(2579) <= (layer6_outputs(5962)) and (layer6_outputs(3672));
    outputs(2580) <= not(layer6_outputs(5463));
    outputs(2581) <= not(layer6_outputs(2901));
    outputs(2582) <= layer6_outputs(821);
    outputs(2583) <= not((layer6_outputs(5632)) and (layer6_outputs(6601)));
    outputs(2584) <= layer6_outputs(158);
    outputs(2585) <= not(layer6_outputs(2216));
    outputs(2586) <= not(layer6_outputs(1139)) or (layer6_outputs(4078));
    outputs(2587) <= (layer6_outputs(6153)) xor (layer6_outputs(6674));
    outputs(2588) <= (layer6_outputs(5890)) xor (layer6_outputs(7577));
    outputs(2589) <= not(layer6_outputs(2544));
    outputs(2590) <= (layer6_outputs(2186)) or (layer6_outputs(6665));
    outputs(2591) <= not(layer6_outputs(4958));
    outputs(2592) <= (layer6_outputs(413)) and (layer6_outputs(4932));
    outputs(2593) <= not(layer6_outputs(3172)) or (layer6_outputs(4237));
    outputs(2594) <= not((layer6_outputs(2387)) xor (layer6_outputs(6649)));
    outputs(2595) <= layer6_outputs(362);
    outputs(2596) <= not(layer6_outputs(6956));
    outputs(2597) <= not((layer6_outputs(7361)) xor (layer6_outputs(2444)));
    outputs(2598) <= not(layer6_outputs(3994));
    outputs(2599) <= (layer6_outputs(602)) or (layer6_outputs(6872));
    outputs(2600) <= layer6_outputs(1738);
    outputs(2601) <= not(layer6_outputs(113));
    outputs(2602) <= (layer6_outputs(705)) xor (layer6_outputs(2646));
    outputs(2603) <= not(layer6_outputs(207)) or (layer6_outputs(6286));
    outputs(2604) <= not(layer6_outputs(5896));
    outputs(2605) <= not(layer6_outputs(7411)) or (layer6_outputs(1686));
    outputs(2606) <= layer6_outputs(4290);
    outputs(2607) <= layer6_outputs(3269);
    outputs(2608) <= layer6_outputs(4927);
    outputs(2609) <= (layer6_outputs(5911)) and not (layer6_outputs(5893));
    outputs(2610) <= not((layer6_outputs(716)) or (layer6_outputs(1390)));
    outputs(2611) <= not((layer6_outputs(3465)) xor (layer6_outputs(2661)));
    outputs(2612) <= not((layer6_outputs(1521)) or (layer6_outputs(2475)));
    outputs(2613) <= not(layer6_outputs(904));
    outputs(2614) <= layer6_outputs(5132);
    outputs(2615) <= not((layer6_outputs(7589)) xor (layer6_outputs(3582)));
    outputs(2616) <= layer6_outputs(4889);
    outputs(2617) <= layer6_outputs(3325);
    outputs(2618) <= (layer6_outputs(1152)) xor (layer6_outputs(3149));
    outputs(2619) <= not(layer6_outputs(6383));
    outputs(2620) <= not((layer6_outputs(1137)) xor (layer6_outputs(3878)));
    outputs(2621) <= (layer6_outputs(3641)) or (layer6_outputs(3959));
    outputs(2622) <= not((layer6_outputs(4023)) xor (layer6_outputs(3521)));
    outputs(2623) <= layer6_outputs(5333);
    outputs(2624) <= layer6_outputs(6941);
    outputs(2625) <= not(layer6_outputs(200));
    outputs(2626) <= not(layer6_outputs(17));
    outputs(2627) <= layer6_outputs(5250);
    outputs(2628) <= layer6_outputs(6424);
    outputs(2629) <= layer6_outputs(7556);
    outputs(2630) <= layer6_outputs(6162);
    outputs(2631) <= layer6_outputs(6827);
    outputs(2632) <= (layer6_outputs(2720)) xor (layer6_outputs(6646));
    outputs(2633) <= (layer6_outputs(2886)) and not (layer6_outputs(7173));
    outputs(2634) <= not(layer6_outputs(5265));
    outputs(2635) <= not((layer6_outputs(1252)) xor (layer6_outputs(4209)));
    outputs(2636) <= not((layer6_outputs(4343)) xor (layer6_outputs(6450)));
    outputs(2637) <= layer6_outputs(7370);
    outputs(2638) <= not((layer6_outputs(4865)) xor (layer6_outputs(2079)));
    outputs(2639) <= not(layer6_outputs(3942));
    outputs(2640) <= not(layer6_outputs(4690));
    outputs(2641) <= layer6_outputs(938);
    outputs(2642) <= (layer6_outputs(4083)) xor (layer6_outputs(6509));
    outputs(2643) <= (layer6_outputs(1895)) xor (layer6_outputs(1733));
    outputs(2644) <= (layer6_outputs(5974)) xor (layer6_outputs(3207));
    outputs(2645) <= not(layer6_outputs(4040));
    outputs(2646) <= layer6_outputs(3377);
    outputs(2647) <= not(layer6_outputs(2796)) or (layer6_outputs(3320));
    outputs(2648) <= not((layer6_outputs(4064)) xor (layer6_outputs(6914)));
    outputs(2649) <= (layer6_outputs(6427)) xor (layer6_outputs(5044));
    outputs(2650) <= not((layer6_outputs(1624)) xor (layer6_outputs(4795)));
    outputs(2651) <= not((layer6_outputs(2460)) xor (layer6_outputs(6060)));
    outputs(2652) <= (layer6_outputs(6500)) xor (layer6_outputs(5031));
    outputs(2653) <= layer6_outputs(7240);
    outputs(2654) <= not((layer6_outputs(4513)) or (layer6_outputs(6957)));
    outputs(2655) <= layer6_outputs(3608);
    outputs(2656) <= layer6_outputs(4990);
    outputs(2657) <= (layer6_outputs(415)) and (layer6_outputs(1941));
    outputs(2658) <= not(layer6_outputs(7186));
    outputs(2659) <= (layer6_outputs(7265)) and not (layer6_outputs(1288));
    outputs(2660) <= not(layer6_outputs(547));
    outputs(2661) <= layer6_outputs(4142);
    outputs(2662) <= (layer6_outputs(192)) or (layer6_outputs(1395));
    outputs(2663) <= layer6_outputs(2547);
    outputs(2664) <= not(layer6_outputs(2572));
    outputs(2665) <= layer6_outputs(4664);
    outputs(2666) <= (layer6_outputs(5958)) or (layer6_outputs(7129));
    outputs(2667) <= layer6_outputs(5558);
    outputs(2668) <= not((layer6_outputs(6144)) xor (layer6_outputs(2619)));
    outputs(2669) <= not((layer6_outputs(5359)) xor (layer6_outputs(5118)));
    outputs(2670) <= not(layer6_outputs(1288));
    outputs(2671) <= layer6_outputs(3066);
    outputs(2672) <= not(layer6_outputs(2998));
    outputs(2673) <= not((layer6_outputs(5105)) xor (layer6_outputs(4817)));
    outputs(2674) <= (layer6_outputs(1810)) or (layer6_outputs(3286));
    outputs(2675) <= layer6_outputs(6854);
    outputs(2676) <= layer6_outputs(7134);
    outputs(2677) <= (layer6_outputs(4850)) xor (layer6_outputs(7353));
    outputs(2678) <= (layer6_outputs(5999)) xor (layer6_outputs(3520));
    outputs(2679) <= layer6_outputs(879);
    outputs(2680) <= (layer6_outputs(4750)) and not (layer6_outputs(695));
    outputs(2681) <= not((layer6_outputs(2965)) xor (layer6_outputs(1131)));
    outputs(2682) <= not(layer6_outputs(2586)) or (layer6_outputs(5363));
    outputs(2683) <= (layer6_outputs(7502)) xor (layer6_outputs(3433));
    outputs(2684) <= layer6_outputs(4710);
    outputs(2685) <= layer6_outputs(7461);
    outputs(2686) <= layer6_outputs(4434);
    outputs(2687) <= not(layer6_outputs(7248));
    outputs(2688) <= layer6_outputs(4315);
    outputs(2689) <= not((layer6_outputs(5815)) xor (layer6_outputs(3810)));
    outputs(2690) <= not((layer6_outputs(2151)) xor (layer6_outputs(2408)));
    outputs(2691) <= layer6_outputs(3770);
    outputs(2692) <= not(layer6_outputs(2000));
    outputs(2693) <= (layer6_outputs(3859)) xor (layer6_outputs(1342));
    outputs(2694) <= layer6_outputs(6963);
    outputs(2695) <= layer6_outputs(6855);
    outputs(2696) <= layer6_outputs(6906);
    outputs(2697) <= not(layer6_outputs(3276));
    outputs(2698) <= not(layer6_outputs(4071));
    outputs(2699) <= not(layer6_outputs(6155)) or (layer6_outputs(6670));
    outputs(2700) <= not(layer6_outputs(3068));
    outputs(2701) <= layer6_outputs(7371);
    outputs(2702) <= not((layer6_outputs(3463)) xor (layer6_outputs(634)));
    outputs(2703) <= layer6_outputs(3278);
    outputs(2704) <= layer6_outputs(3565);
    outputs(2705) <= not(layer6_outputs(5219));
    outputs(2706) <= not(layer6_outputs(1254));
    outputs(2707) <= not((layer6_outputs(4896)) xor (layer6_outputs(6148)));
    outputs(2708) <= not(layer6_outputs(1501));
    outputs(2709) <= not((layer6_outputs(7504)) xor (layer6_outputs(716)));
    outputs(2710) <= not(layer6_outputs(3276));
    outputs(2711) <= layer6_outputs(4299);
    outputs(2712) <= not(layer6_outputs(6212));
    outputs(2713) <= not(layer6_outputs(486));
    outputs(2714) <= not(layer6_outputs(356));
    outputs(2715) <= (layer6_outputs(5362)) and not (layer6_outputs(7295));
    outputs(2716) <= layer6_outputs(154);
    outputs(2717) <= not((layer6_outputs(3360)) and (layer6_outputs(4752)));
    outputs(2718) <= not(layer6_outputs(7389));
    outputs(2719) <= not((layer6_outputs(3588)) xor (layer6_outputs(7449)));
    outputs(2720) <= not(layer6_outputs(3100)) or (layer6_outputs(4002));
    outputs(2721) <= not((layer6_outputs(3764)) xor (layer6_outputs(5806)));
    outputs(2722) <= (layer6_outputs(446)) xor (layer6_outputs(514));
    outputs(2723) <= (layer6_outputs(4715)) xor (layer6_outputs(7599));
    outputs(2724) <= not((layer6_outputs(2663)) xor (layer6_outputs(1988)));
    outputs(2725) <= not(layer6_outputs(1150));
    outputs(2726) <= not((layer6_outputs(3191)) and (layer6_outputs(4631)));
    outputs(2727) <= (layer6_outputs(7063)) xor (layer6_outputs(4837));
    outputs(2728) <= layer6_outputs(2822);
    outputs(2729) <= layer6_outputs(4551);
    outputs(2730) <= not((layer6_outputs(2326)) xor (layer6_outputs(2672)));
    outputs(2731) <= layer6_outputs(3199);
    outputs(2732) <= not(layer6_outputs(3960)) or (layer6_outputs(382));
    outputs(2733) <= layer6_outputs(5268);
    outputs(2734) <= (layer6_outputs(5409)) xor (layer6_outputs(4235));
    outputs(2735) <= layer6_outputs(2492);
    outputs(2736) <= not(layer6_outputs(1263)) or (layer6_outputs(6553));
    outputs(2737) <= not(layer6_outputs(690));
    outputs(2738) <= not((layer6_outputs(1326)) or (layer6_outputs(3632)));
    outputs(2739) <= layer6_outputs(3435);
    outputs(2740) <= not(layer6_outputs(271));
    outputs(2741) <= (layer6_outputs(7126)) xor (layer6_outputs(7043));
    outputs(2742) <= (layer6_outputs(6277)) and (layer6_outputs(6207));
    outputs(2743) <= layer6_outputs(7037);
    outputs(2744) <= not((layer6_outputs(5134)) xor (layer6_outputs(3390)));
    outputs(2745) <= layer6_outputs(4055);
    outputs(2746) <= layer6_outputs(6421);
    outputs(2747) <= layer6_outputs(3559);
    outputs(2748) <= (layer6_outputs(3961)) or (layer6_outputs(7519));
    outputs(2749) <= not(layer6_outputs(1278)) or (layer6_outputs(2203));
    outputs(2750) <= layer6_outputs(2169);
    outputs(2751) <= not(layer6_outputs(6504)) or (layer6_outputs(1051));
    outputs(2752) <= not((layer6_outputs(6104)) and (layer6_outputs(5376)));
    outputs(2753) <= not((layer6_outputs(2471)) xor (layer6_outputs(3358)));
    outputs(2754) <= not(layer6_outputs(6452));
    outputs(2755) <= not(layer6_outputs(6926));
    outputs(2756) <= not(layer6_outputs(3086));
    outputs(2757) <= not(layer6_outputs(5655));
    outputs(2758) <= not(layer6_outputs(4046));
    outputs(2759) <= not(layer6_outputs(6002));
    outputs(2760) <= not((layer6_outputs(3191)) xor (layer6_outputs(2821)));
    outputs(2761) <= not((layer6_outputs(4974)) or (layer6_outputs(1529)));
    outputs(2762) <= layer6_outputs(5807);
    outputs(2763) <= layer6_outputs(2472);
    outputs(2764) <= layer6_outputs(223);
    outputs(2765) <= (layer6_outputs(1539)) and not (layer6_outputs(4993));
    outputs(2766) <= not(layer6_outputs(1481));
    outputs(2767) <= not(layer6_outputs(6603));
    outputs(2768) <= (layer6_outputs(1281)) and (layer6_outputs(4991));
    outputs(2769) <= (layer6_outputs(7298)) xor (layer6_outputs(2734));
    outputs(2770) <= layer6_outputs(4614);
    outputs(2771) <= layer6_outputs(5669);
    outputs(2772) <= (layer6_outputs(6855)) xor (layer6_outputs(450));
    outputs(2773) <= not(layer6_outputs(768));
    outputs(2774) <= not(layer6_outputs(1890));
    outputs(2775) <= (layer6_outputs(7059)) and not (layer6_outputs(3449));
    outputs(2776) <= layer6_outputs(1480);
    outputs(2777) <= layer6_outputs(3);
    outputs(2778) <= not((layer6_outputs(597)) and (layer6_outputs(300)));
    outputs(2779) <= not((layer6_outputs(333)) or (layer6_outputs(832)));
    outputs(2780) <= layer6_outputs(3430);
    outputs(2781) <= layer6_outputs(4210);
    outputs(2782) <= not((layer6_outputs(4337)) xor (layer6_outputs(983)));
    outputs(2783) <= (layer6_outputs(6439)) xor (layer6_outputs(245));
    outputs(2784) <= layer6_outputs(6632);
    outputs(2785) <= layer6_outputs(149);
    outputs(2786) <= not(layer6_outputs(3551));
    outputs(2787) <= layer6_outputs(1956);
    outputs(2788) <= (layer6_outputs(7134)) and not (layer6_outputs(1251));
    outputs(2789) <= not(layer6_outputs(557)) or (layer6_outputs(6373));
    outputs(2790) <= layer6_outputs(230);
    outputs(2791) <= not(layer6_outputs(7276));
    outputs(2792) <= not(layer6_outputs(3306));
    outputs(2793) <= not(layer6_outputs(3831));
    outputs(2794) <= not((layer6_outputs(2985)) xor (layer6_outputs(5604)));
    outputs(2795) <= (layer6_outputs(1613)) and not (layer6_outputs(191));
    outputs(2796) <= not(layer6_outputs(7557));
    outputs(2797) <= (layer6_outputs(4315)) and (layer6_outputs(3042));
    outputs(2798) <= layer6_outputs(5967);
    outputs(2799) <= layer6_outputs(7441);
    outputs(2800) <= layer6_outputs(6927);
    outputs(2801) <= not(layer6_outputs(4909));
    outputs(2802) <= not(layer6_outputs(2597));
    outputs(2803) <= not(layer6_outputs(5351));
    outputs(2804) <= not(layer6_outputs(3525));
    outputs(2805) <= not((layer6_outputs(6724)) xor (layer6_outputs(4259)));
    outputs(2806) <= not(layer6_outputs(4090));
    outputs(2807) <= not((layer6_outputs(4737)) xor (layer6_outputs(183)));
    outputs(2808) <= not(layer6_outputs(674));
    outputs(2809) <= layer6_outputs(2753);
    outputs(2810) <= layer6_outputs(3626);
    outputs(2811) <= layer6_outputs(5481);
    outputs(2812) <= layer6_outputs(3232);
    outputs(2813) <= (layer6_outputs(5886)) or (layer6_outputs(143));
    outputs(2814) <= not(layer6_outputs(5542)) or (layer6_outputs(1279));
    outputs(2815) <= not((layer6_outputs(3316)) xor (layer6_outputs(4543)));
    outputs(2816) <= not((layer6_outputs(2880)) xor (layer6_outputs(3194)));
    outputs(2817) <= not(layer6_outputs(3038)) or (layer6_outputs(2203));
    outputs(2818) <= not((layer6_outputs(7165)) xor (layer6_outputs(810)));
    outputs(2819) <= not((layer6_outputs(6033)) xor (layer6_outputs(5710)));
    outputs(2820) <= not((layer6_outputs(2493)) xor (layer6_outputs(2059)));
    outputs(2821) <= layer6_outputs(4093);
    outputs(2822) <= not(layer6_outputs(3337));
    outputs(2823) <= layer6_outputs(4977);
    outputs(2824) <= not((layer6_outputs(4474)) xor (layer6_outputs(2353)));
    outputs(2825) <= (layer6_outputs(1171)) xor (layer6_outputs(2148));
    outputs(2826) <= not((layer6_outputs(7404)) xor (layer6_outputs(3602)));
    outputs(2827) <= not(layer6_outputs(1826));
    outputs(2828) <= (layer6_outputs(5582)) xor (layer6_outputs(6276));
    outputs(2829) <= not(layer6_outputs(517));
    outputs(2830) <= not((layer6_outputs(3849)) or (layer6_outputs(4618)));
    outputs(2831) <= layer6_outputs(7210);
    outputs(2832) <= not((layer6_outputs(5480)) xor (layer6_outputs(4232)));
    outputs(2833) <= layer6_outputs(3543);
    outputs(2834) <= not(layer6_outputs(2181)) or (layer6_outputs(5835));
    outputs(2835) <= (layer6_outputs(5208)) xor (layer6_outputs(4694));
    outputs(2836) <= layer6_outputs(894);
    outputs(2837) <= layer6_outputs(2062);
    outputs(2838) <= not((layer6_outputs(4637)) xor (layer6_outputs(7652)));
    outputs(2839) <= not(layer6_outputs(4807));
    outputs(2840) <= not(layer6_outputs(2155)) or (layer6_outputs(2346));
    outputs(2841) <= not(layer6_outputs(2464));
    outputs(2842) <= not((layer6_outputs(1640)) xor (layer6_outputs(4376)));
    outputs(2843) <= not((layer6_outputs(7001)) or (layer6_outputs(6956)));
    outputs(2844) <= layer6_outputs(2311);
    outputs(2845) <= (layer6_outputs(369)) xor (layer6_outputs(6928));
    outputs(2846) <= (layer6_outputs(2253)) xor (layer6_outputs(6643));
    outputs(2847) <= (layer6_outputs(5024)) xor (layer6_outputs(5047));
    outputs(2848) <= not(layer6_outputs(4391));
    outputs(2849) <= not(layer6_outputs(5948));
    outputs(2850) <= not((layer6_outputs(191)) xor (layer6_outputs(6131)));
    outputs(2851) <= not(layer6_outputs(5120));
    outputs(2852) <= not(layer6_outputs(5513));
    outputs(2853) <= (layer6_outputs(38)) xor (layer6_outputs(2078));
    outputs(2854) <= (layer6_outputs(7268)) and (layer6_outputs(5875));
    outputs(2855) <= not((layer6_outputs(509)) xor (layer6_outputs(6483)));
    outputs(2856) <= layer6_outputs(466);
    outputs(2857) <= (layer6_outputs(52)) and not (layer6_outputs(3946));
    outputs(2858) <= not((layer6_outputs(7380)) and (layer6_outputs(1555)));
    outputs(2859) <= not(layer6_outputs(3943));
    outputs(2860) <= not(layer6_outputs(5370));
    outputs(2861) <= not((layer6_outputs(4259)) xor (layer6_outputs(4200)));
    outputs(2862) <= not(layer6_outputs(4466));
    outputs(2863) <= not(layer6_outputs(6756));
    outputs(2864) <= (layer6_outputs(2045)) or (layer6_outputs(1309));
    outputs(2865) <= layer6_outputs(2492);
    outputs(2866) <= (layer6_outputs(1784)) xor (layer6_outputs(4010));
    outputs(2867) <= not(layer6_outputs(6269));
    outputs(2868) <= (layer6_outputs(5026)) and not (layer6_outputs(1196));
    outputs(2869) <= (layer6_outputs(4288)) and not (layer6_outputs(635));
    outputs(2870) <= layer6_outputs(1258);
    outputs(2871) <= not(layer6_outputs(5955));
    outputs(2872) <= (layer6_outputs(5319)) and not (layer6_outputs(6269));
    outputs(2873) <= layer6_outputs(4453);
    outputs(2874) <= not(layer6_outputs(973));
    outputs(2875) <= layer6_outputs(2053);
    outputs(2876) <= layer6_outputs(5742);
    outputs(2877) <= (layer6_outputs(7250)) and not (layer6_outputs(347));
    outputs(2878) <= not(layer6_outputs(4415));
    outputs(2879) <= layer6_outputs(717);
    outputs(2880) <= (layer6_outputs(127)) or (layer6_outputs(7664));
    outputs(2881) <= not((layer6_outputs(6873)) xor (layer6_outputs(5096)));
    outputs(2882) <= not(layer6_outputs(464));
    outputs(2883) <= layer6_outputs(2027);
    outputs(2884) <= layer6_outputs(7482);
    outputs(2885) <= not(layer6_outputs(5830)) or (layer6_outputs(4253));
    outputs(2886) <= layer6_outputs(5616);
    outputs(2887) <= (layer6_outputs(5601)) and not (layer6_outputs(6196));
    outputs(2888) <= layer6_outputs(5433);
    outputs(2889) <= layer6_outputs(3411);
    outputs(2890) <= (layer6_outputs(6563)) and (layer6_outputs(6976));
    outputs(2891) <= layer6_outputs(2423);
    outputs(2892) <= not((layer6_outputs(168)) xor (layer6_outputs(2879)));
    outputs(2893) <= not(layer6_outputs(1817));
    outputs(2894) <= not((layer6_outputs(3521)) xor (layer6_outputs(2886)));
    outputs(2895) <= not((layer6_outputs(3446)) xor (layer6_outputs(7655)));
    outputs(2896) <= not((layer6_outputs(5473)) or (layer6_outputs(966)));
    outputs(2897) <= not(layer6_outputs(4746)) or (layer6_outputs(5556));
    outputs(2898) <= not(layer6_outputs(3389));
    outputs(2899) <= not(layer6_outputs(3576)) or (layer6_outputs(5835));
    outputs(2900) <= not(layer6_outputs(3118));
    outputs(2901) <= not(layer6_outputs(66)) or (layer6_outputs(96));
    outputs(2902) <= not(layer6_outputs(5759));
    outputs(2903) <= layer6_outputs(5605);
    outputs(2904) <= not(layer6_outputs(679));
    outputs(2905) <= not(layer6_outputs(1461));
    outputs(2906) <= not(layer6_outputs(3501));
    outputs(2907) <= (layer6_outputs(3339)) xor (layer6_outputs(2056));
    outputs(2908) <= not(layer6_outputs(5490));
    outputs(2909) <= not(layer6_outputs(5828));
    outputs(2910) <= (layer6_outputs(3703)) xor (layer6_outputs(6627));
    outputs(2911) <= not((layer6_outputs(4612)) xor (layer6_outputs(5185)));
    outputs(2912) <= not(layer6_outputs(4773));
    outputs(2913) <= not(layer6_outputs(5038));
    outputs(2914) <= layer6_outputs(6237);
    outputs(2915) <= not(layer6_outputs(3055));
    outputs(2916) <= not(layer6_outputs(6047));
    outputs(2917) <= (layer6_outputs(1426)) xor (layer6_outputs(6889));
    outputs(2918) <= (layer6_outputs(39)) xor (layer6_outputs(7138));
    outputs(2919) <= (layer6_outputs(2358)) and not (layer6_outputs(7066));
    outputs(2920) <= layer6_outputs(4903);
    outputs(2921) <= not(layer6_outputs(1631));
    outputs(2922) <= not(layer6_outputs(6942));
    outputs(2923) <= not(layer6_outputs(2302));
    outputs(2924) <= layer6_outputs(5866);
    outputs(2925) <= layer6_outputs(5723);
    outputs(2926) <= not(layer6_outputs(5736));
    outputs(2927) <= not(layer6_outputs(4765));
    outputs(2928) <= layer6_outputs(757);
    outputs(2929) <= not(layer6_outputs(1178));
    outputs(2930) <= not(layer6_outputs(2144));
    outputs(2931) <= not(layer6_outputs(2177));
    outputs(2932) <= not((layer6_outputs(5309)) or (layer6_outputs(6681)));
    outputs(2933) <= not(layer6_outputs(1018));
    outputs(2934) <= not(layer6_outputs(5530));
    outputs(2935) <= layer6_outputs(4089);
    outputs(2936) <= not(layer6_outputs(6926));
    outputs(2937) <= (layer6_outputs(5037)) xor (layer6_outputs(1815));
    outputs(2938) <= (layer6_outputs(5085)) and not (layer6_outputs(6250));
    outputs(2939) <= not(layer6_outputs(2437));
    outputs(2940) <= layer6_outputs(3195);
    outputs(2941) <= layer6_outputs(3530);
    outputs(2942) <= layer6_outputs(7096);
    outputs(2943) <= not(layer6_outputs(5586));
    outputs(2944) <= (layer6_outputs(642)) and (layer6_outputs(6470));
    outputs(2945) <= layer6_outputs(488);
    outputs(2946) <= layer6_outputs(4830);
    outputs(2947) <= (layer6_outputs(2960)) or (layer6_outputs(6464));
    outputs(2948) <= (layer6_outputs(3518)) xor (layer6_outputs(1971));
    outputs(2949) <= (layer6_outputs(1364)) xor (layer6_outputs(5786));
    outputs(2950) <= not(layer6_outputs(1544));
    outputs(2951) <= not(layer6_outputs(3768));
    outputs(2952) <= not(layer6_outputs(3766));
    outputs(2953) <= layer6_outputs(7245);
    outputs(2954) <= layer6_outputs(5372);
    outputs(2955) <= (layer6_outputs(7146)) and not (layer6_outputs(505));
    outputs(2956) <= not((layer6_outputs(5595)) xor (layer6_outputs(1003)));
    outputs(2957) <= (layer6_outputs(3333)) xor (layer6_outputs(2801));
    outputs(2958) <= (layer6_outputs(2584)) and (layer6_outputs(6658));
    outputs(2959) <= not(layer6_outputs(4968));
    outputs(2960) <= layer6_outputs(1421);
    outputs(2961) <= not(layer6_outputs(57));
    outputs(2962) <= not((layer6_outputs(5626)) xor (layer6_outputs(5410)));
    outputs(2963) <= not(layer6_outputs(1664));
    outputs(2964) <= layer6_outputs(6821);
    outputs(2965) <= (layer6_outputs(1355)) xor (layer6_outputs(563));
    outputs(2966) <= not(layer6_outputs(40));
    outputs(2967) <= (layer6_outputs(4891)) xor (layer6_outputs(6005));
    outputs(2968) <= (layer6_outputs(7337)) xor (layer6_outputs(7521));
    outputs(2969) <= layer6_outputs(7471);
    outputs(2970) <= layer6_outputs(5337);
    outputs(2971) <= (layer6_outputs(2419)) xor (layer6_outputs(3112));
    outputs(2972) <= not(layer6_outputs(811));
    outputs(2973) <= not(layer6_outputs(3840));
    outputs(2974) <= (layer6_outputs(4952)) xor (layer6_outputs(7197));
    outputs(2975) <= not((layer6_outputs(3483)) xor (layer6_outputs(2772)));
    outputs(2976) <= not(layer6_outputs(3505));
    outputs(2977) <= layer6_outputs(6489);
    outputs(2978) <= not((layer6_outputs(7342)) xor (layer6_outputs(5761)));
    outputs(2979) <= not(layer6_outputs(228));
    outputs(2980) <= not((layer6_outputs(1024)) xor (layer6_outputs(2184)));
    outputs(2981) <= layer6_outputs(6187);
    outputs(2982) <= (layer6_outputs(1782)) and not (layer6_outputs(2455));
    outputs(2983) <= (layer6_outputs(3349)) xor (layer6_outputs(3618));
    outputs(2984) <= layer6_outputs(4393);
    outputs(2985) <= not(layer6_outputs(3351));
    outputs(2986) <= (layer6_outputs(1745)) xor (layer6_outputs(618));
    outputs(2987) <= not(layer6_outputs(2765));
    outputs(2988) <= not(layer6_outputs(7464));
    outputs(2989) <= not(layer6_outputs(4804));
    outputs(2990) <= layer6_outputs(928);
    outputs(2991) <= not(layer6_outputs(5257));
    outputs(2992) <= not((layer6_outputs(6752)) xor (layer6_outputs(7580)));
    outputs(2993) <= not(layer6_outputs(2538));
    outputs(2994) <= not(layer6_outputs(5273));
    outputs(2995) <= (layer6_outputs(3558)) and not (layer6_outputs(2009));
    outputs(2996) <= layer6_outputs(7146);
    outputs(2997) <= (layer6_outputs(2888)) xor (layer6_outputs(6720));
    outputs(2998) <= not(layer6_outputs(579)) or (layer6_outputs(3320));
    outputs(2999) <= not((layer6_outputs(2834)) xor (layer6_outputs(4573)));
    outputs(3000) <= not(layer6_outputs(7446));
    outputs(3001) <= not(layer6_outputs(1875));
    outputs(3002) <= (layer6_outputs(4825)) or (layer6_outputs(1292));
    outputs(3003) <= not(layer6_outputs(2785)) or (layer6_outputs(6165));
    outputs(3004) <= not((layer6_outputs(7060)) xor (layer6_outputs(197)));
    outputs(3005) <= not((layer6_outputs(2004)) or (layer6_outputs(1503)));
    outputs(3006) <= not(layer6_outputs(2487));
    outputs(3007) <= not(layer6_outputs(5500));
    outputs(3008) <= (layer6_outputs(3825)) and not (layer6_outputs(5890));
    outputs(3009) <= not((layer6_outputs(7573)) and (layer6_outputs(132)));
    outputs(3010) <= (layer6_outputs(1322)) xor (layer6_outputs(5975));
    outputs(3011) <= layer6_outputs(1880);
    outputs(3012) <= (layer6_outputs(3828)) xor (layer6_outputs(2899));
    outputs(3013) <= layer6_outputs(4079);
    outputs(3014) <= (layer6_outputs(821)) and not (layer6_outputs(4866));
    outputs(3015) <= layer6_outputs(1579);
    outputs(3016) <= not((layer6_outputs(5518)) xor (layer6_outputs(1447)));
    outputs(3017) <= not(layer6_outputs(2581));
    outputs(3018) <= layer6_outputs(5108);
    outputs(3019) <= not((layer6_outputs(6586)) xor (layer6_outputs(4339)));
    outputs(3020) <= layer6_outputs(7119);
    outputs(3021) <= not((layer6_outputs(5478)) xor (layer6_outputs(3757)));
    outputs(3022) <= layer6_outputs(1292);
    outputs(3023) <= not((layer6_outputs(923)) or (layer6_outputs(6860)));
    outputs(3024) <= (layer6_outputs(5521)) and not (layer6_outputs(6729));
    outputs(3025) <= layer6_outputs(6968);
    outputs(3026) <= layer6_outputs(6960);
    outputs(3027) <= layer6_outputs(6766);
    outputs(3028) <= not(layer6_outputs(5773)) or (layer6_outputs(7007));
    outputs(3029) <= (layer6_outputs(6817)) xor (layer6_outputs(7));
    outputs(3030) <= layer6_outputs(6829);
    outputs(3031) <= not(layer6_outputs(2302));
    outputs(3032) <= not((layer6_outputs(4199)) or (layer6_outputs(1892)));
    outputs(3033) <= (layer6_outputs(394)) xor (layer6_outputs(3427));
    outputs(3034) <= not((layer6_outputs(2893)) xor (layer6_outputs(4080)));
    outputs(3035) <= (layer6_outputs(3018)) xor (layer6_outputs(6028));
    outputs(3036) <= not(layer6_outputs(936));
    outputs(3037) <= layer6_outputs(6358);
    outputs(3038) <= layer6_outputs(2481);
    outputs(3039) <= (layer6_outputs(7396)) xor (layer6_outputs(7321));
    outputs(3040) <= not(layer6_outputs(562));
    outputs(3041) <= not((layer6_outputs(3564)) or (layer6_outputs(65)));
    outputs(3042) <= layer6_outputs(4667);
    outputs(3043) <= not((layer6_outputs(3721)) xor (layer6_outputs(7544)));
    outputs(3044) <= layer6_outputs(4312);
    outputs(3045) <= (layer6_outputs(5716)) and not (layer6_outputs(1000));
    outputs(3046) <= (layer6_outputs(6625)) and not (layer6_outputs(3688));
    outputs(3047) <= not(layer6_outputs(4313));
    outputs(3048) <= layer6_outputs(7324);
    outputs(3049) <= not(layer6_outputs(1907));
    outputs(3050) <= not(layer6_outputs(598));
    outputs(3051) <= (layer6_outputs(6264)) xor (layer6_outputs(5229));
    outputs(3052) <= (layer6_outputs(1313)) and not (layer6_outputs(6055));
    outputs(3053) <= layer6_outputs(5011);
    outputs(3054) <= layer6_outputs(625);
    outputs(3055) <= not(layer6_outputs(7659));
    outputs(3056) <= (layer6_outputs(5109)) or (layer6_outputs(1596));
    outputs(3057) <= (layer6_outputs(1524)) xor (layer6_outputs(5408));
    outputs(3058) <= not((layer6_outputs(4197)) or (layer6_outputs(3790)));
    outputs(3059) <= (layer6_outputs(3924)) and not (layer6_outputs(180));
    outputs(3060) <= layer6_outputs(1125);
    outputs(3061) <= (layer6_outputs(2994)) xor (layer6_outputs(7521));
    outputs(3062) <= layer6_outputs(5644);
    outputs(3063) <= not(layer6_outputs(2246)) or (layer6_outputs(344));
    outputs(3064) <= layer6_outputs(322);
    outputs(3065) <= layer6_outputs(5920);
    outputs(3066) <= not(layer6_outputs(1505));
    outputs(3067) <= not(layer6_outputs(921)) or (layer6_outputs(1237));
    outputs(3068) <= (layer6_outputs(7325)) xor (layer6_outputs(5511));
    outputs(3069) <= (layer6_outputs(4941)) xor (layer6_outputs(5406));
    outputs(3070) <= layer6_outputs(359);
    outputs(3071) <= not(layer6_outputs(6685));
    outputs(3072) <= not((layer6_outputs(794)) xor (layer6_outputs(1753)));
    outputs(3073) <= not(layer6_outputs(1789));
    outputs(3074) <= not(layer6_outputs(4408));
    outputs(3075) <= layer6_outputs(3138);
    outputs(3076) <= not(layer6_outputs(6456));
    outputs(3077) <= (layer6_outputs(6909)) and not (layer6_outputs(962));
    outputs(3078) <= (layer6_outputs(4347)) xor (layer6_outputs(3941));
    outputs(3079) <= not((layer6_outputs(1541)) xor (layer6_outputs(5864)));
    outputs(3080) <= not(layer6_outputs(3531));
    outputs(3081) <= layer6_outputs(5721);
    outputs(3082) <= layer6_outputs(5810);
    outputs(3083) <= not(layer6_outputs(148));
    outputs(3084) <= not(layer6_outputs(3863));
    outputs(3085) <= (layer6_outputs(3850)) and (layer6_outputs(400));
    outputs(3086) <= not((layer6_outputs(2683)) and (layer6_outputs(1980)));
    outputs(3087) <= layer6_outputs(135);
    outputs(3088) <= not((layer6_outputs(4541)) xor (layer6_outputs(6650)));
    outputs(3089) <= not(layer6_outputs(2952));
    outputs(3090) <= not(layer6_outputs(6906));
    outputs(3091) <= layer6_outputs(3417);
    outputs(3092) <= not((layer6_outputs(6812)) xor (layer6_outputs(5407)));
    outputs(3093) <= not(layer6_outputs(5917));
    outputs(3094) <= (layer6_outputs(4122)) and not (layer6_outputs(6751));
    outputs(3095) <= not(layer6_outputs(3949));
    outputs(3096) <= layer6_outputs(1253);
    outputs(3097) <= not(layer6_outputs(1094));
    outputs(3098) <= not((layer6_outputs(2776)) or (layer6_outputs(668)));
    outputs(3099) <= not(layer6_outputs(5192));
    outputs(3100) <= (layer6_outputs(2248)) xor (layer6_outputs(903));
    outputs(3101) <= layer6_outputs(4938);
    outputs(3102) <= not(layer6_outputs(2350));
    outputs(3103) <= not((layer6_outputs(7083)) xor (layer6_outputs(7653)));
    outputs(3104) <= (layer6_outputs(6384)) and (layer6_outputs(4361));
    outputs(3105) <= (layer6_outputs(3392)) xor (layer6_outputs(767));
    outputs(3106) <= (layer6_outputs(2443)) xor (layer6_outputs(2962));
    outputs(3107) <= layer6_outputs(4419);
    outputs(3108) <= layer6_outputs(141);
    outputs(3109) <= not(layer6_outputs(4616)) or (layer6_outputs(313));
    outputs(3110) <= layer6_outputs(5294);
    outputs(3111) <= (layer6_outputs(6604)) xor (layer6_outputs(4443));
    outputs(3112) <= not(layer6_outputs(3972));
    outputs(3113) <= (layer6_outputs(3170)) xor (layer6_outputs(3229));
    outputs(3114) <= (layer6_outputs(7135)) xor (layer6_outputs(5040));
    outputs(3115) <= layer6_outputs(3719);
    outputs(3116) <= layer6_outputs(5833);
    outputs(3117) <= layer6_outputs(303);
    outputs(3118) <= layer6_outputs(3182);
    outputs(3119) <= layer6_outputs(3650);
    outputs(3120) <= not(layer6_outputs(3143));
    outputs(3121) <= not((layer6_outputs(3468)) and (layer6_outputs(2708)));
    outputs(3122) <= not(layer6_outputs(3715));
    outputs(3123) <= layer6_outputs(6567);
    outputs(3124) <= (layer6_outputs(85)) xor (layer6_outputs(7013));
    outputs(3125) <= (layer6_outputs(319)) xor (layer6_outputs(7643));
    outputs(3126) <= not(layer6_outputs(5963));
    outputs(3127) <= (layer6_outputs(1460)) and not (layer6_outputs(430));
    outputs(3128) <= layer6_outputs(5734);
    outputs(3129) <= (layer6_outputs(3666)) xor (layer6_outputs(7224));
    outputs(3130) <= not(layer6_outputs(6695));
    outputs(3131) <= (layer6_outputs(6116)) xor (layer6_outputs(4965));
    outputs(3132) <= not(layer6_outputs(3003));
    outputs(3133) <= not(layer6_outputs(5800));
    outputs(3134) <= (layer6_outputs(7114)) xor (layer6_outputs(1137));
    outputs(3135) <= not(layer6_outputs(1480));
    outputs(3136) <= not(layer6_outputs(1069)) or (layer6_outputs(2962));
    outputs(3137) <= not(layer6_outputs(3718)) or (layer6_outputs(7564));
    outputs(3138) <= layer6_outputs(6946);
    outputs(3139) <= not(layer6_outputs(6608));
    outputs(3140) <= (layer6_outputs(1220)) xor (layer6_outputs(4138));
    outputs(3141) <= layer6_outputs(1060);
    outputs(3142) <= layer6_outputs(4855);
    outputs(3143) <= (layer6_outputs(2413)) and not (layer6_outputs(429));
    outputs(3144) <= layer6_outputs(1242);
    outputs(3145) <= (layer6_outputs(2625)) xor (layer6_outputs(600));
    outputs(3146) <= layer6_outputs(1597);
    outputs(3147) <= not(layer6_outputs(3196));
    outputs(3148) <= (layer6_outputs(6466)) xor (layer6_outputs(2681));
    outputs(3149) <= layer6_outputs(2957);
    outputs(3150) <= layer6_outputs(3245);
    outputs(3151) <= (layer6_outputs(1783)) xor (layer6_outputs(427));
    outputs(3152) <= layer6_outputs(5952);
    outputs(3153) <= layer6_outputs(6344);
    outputs(3154) <= not(layer6_outputs(4033));
    outputs(3155) <= not((layer6_outputs(6973)) xor (layer6_outputs(3970)));
    outputs(3156) <= layer6_outputs(1571);
    outputs(3157) <= not(layer6_outputs(1293));
    outputs(3158) <= not(layer6_outputs(3169)) or (layer6_outputs(4268));
    outputs(3159) <= layer6_outputs(855);
    outputs(3160) <= (layer6_outputs(2543)) xor (layer6_outputs(2967));
    outputs(3161) <= not(layer6_outputs(3359));
    outputs(3162) <= layer6_outputs(6392);
    outputs(3163) <= layer6_outputs(6591);
    outputs(3164) <= (layer6_outputs(312)) xor (layer6_outputs(612));
    outputs(3165) <= layer6_outputs(3113);
    outputs(3166) <= (layer6_outputs(3564)) and not (layer6_outputs(1166));
    outputs(3167) <= layer6_outputs(4909);
    outputs(3168) <= not(layer6_outputs(5652));
    outputs(3169) <= layer6_outputs(2654);
    outputs(3170) <= not(layer6_outputs(1969));
    outputs(3171) <= not(layer6_outputs(5917));
    outputs(3172) <= layer6_outputs(3609);
    outputs(3173) <= layer6_outputs(1743);
    outputs(3174) <= not((layer6_outputs(3270)) xor (layer6_outputs(5912)));
    outputs(3175) <= layer6_outputs(6091);
    outputs(3176) <= not(layer6_outputs(3251));
    outputs(3177) <= layer6_outputs(4147);
    outputs(3178) <= (layer6_outputs(6718)) xor (layer6_outputs(1721));
    outputs(3179) <= not(layer6_outputs(6307));
    outputs(3180) <= not(layer6_outputs(1130));
    outputs(3181) <= not(layer6_outputs(1318));
    outputs(3182) <= layer6_outputs(6309);
    outputs(3183) <= not(layer6_outputs(5489));
    outputs(3184) <= not((layer6_outputs(3039)) or (layer6_outputs(3232)));
    outputs(3185) <= layer6_outputs(3416);
    outputs(3186) <= layer6_outputs(2031);
    outputs(3187) <= not(layer6_outputs(5000));
    outputs(3188) <= (layer6_outputs(7133)) xor (layer6_outputs(5146));
    outputs(3189) <= not(layer6_outputs(5130));
    outputs(3190) <= not(layer6_outputs(1832));
    outputs(3191) <= layer6_outputs(4669);
    outputs(3192) <= not(layer6_outputs(112));
    outputs(3193) <= (layer6_outputs(3178)) and not (layer6_outputs(5771));
    outputs(3194) <= not((layer6_outputs(2527)) xor (layer6_outputs(5230)));
    outputs(3195) <= (layer6_outputs(5345)) and not (layer6_outputs(1753));
    outputs(3196) <= layer6_outputs(1650);
    outputs(3197) <= not((layer6_outputs(2112)) xor (layer6_outputs(7224)));
    outputs(3198) <= not(layer6_outputs(1591));
    outputs(3199) <= not(layer6_outputs(7503));
    outputs(3200) <= layer6_outputs(916);
    outputs(3201) <= layer6_outputs(3609);
    outputs(3202) <= (layer6_outputs(1067)) xor (layer6_outputs(396));
    outputs(3203) <= (layer6_outputs(3102)) xor (layer6_outputs(1666));
    outputs(3204) <= (layer6_outputs(5493)) xor (layer6_outputs(1212));
    outputs(3205) <= layer6_outputs(4645);
    outputs(3206) <= not(layer6_outputs(7414));
    outputs(3207) <= not(layer6_outputs(179));
    outputs(3208) <= not(layer6_outputs(7233));
    outputs(3209) <= (layer6_outputs(2838)) and (layer6_outputs(4516));
    outputs(3210) <= not(layer6_outputs(3955));
    outputs(3211) <= not((layer6_outputs(4500)) xor (layer6_outputs(6276)));
    outputs(3212) <= not(layer6_outputs(3051));
    outputs(3213) <= layer6_outputs(3476);
    outputs(3214) <= layer6_outputs(5600);
    outputs(3215) <= not(layer6_outputs(7658));
    outputs(3216) <= (layer6_outputs(4774)) and (layer6_outputs(3660));
    outputs(3217) <= layer6_outputs(6224);
    outputs(3218) <= layer6_outputs(3203);
    outputs(3219) <= not((layer6_outputs(3303)) xor (layer6_outputs(401)));
    outputs(3220) <= not((layer6_outputs(2755)) xor (layer6_outputs(1206)));
    outputs(3221) <= not(layer6_outputs(5237));
    outputs(3222) <= not(layer6_outputs(563)) or (layer6_outputs(6555));
    outputs(3223) <= not((layer6_outputs(2681)) or (layer6_outputs(6568)));
    outputs(3224) <= not(layer6_outputs(5963));
    outputs(3225) <= (layer6_outputs(6004)) and not (layer6_outputs(5788));
    outputs(3226) <= (layer6_outputs(561)) xor (layer6_outputs(6791));
    outputs(3227) <= layer6_outputs(2944);
    outputs(3228) <= not(layer6_outputs(3526));
    outputs(3229) <= (layer6_outputs(3823)) xor (layer6_outputs(2041));
    outputs(3230) <= not((layer6_outputs(2846)) and (layer6_outputs(877)));
    outputs(3231) <= layer6_outputs(6323);
    outputs(3232) <= not((layer6_outputs(5660)) or (layer6_outputs(412)));
    outputs(3233) <= layer6_outputs(2104);
    outputs(3234) <= (layer6_outputs(4656)) and not (layer6_outputs(6033));
    outputs(3235) <= not(layer6_outputs(350));
    outputs(3236) <= not(layer6_outputs(661));
    outputs(3237) <= layer6_outputs(1503);
    outputs(3238) <= not((layer6_outputs(4309)) or (layer6_outputs(3611)));
    outputs(3239) <= (layer6_outputs(7147)) xor (layer6_outputs(2164));
    outputs(3240) <= not((layer6_outputs(5765)) xor (layer6_outputs(3376)));
    outputs(3241) <= not(layer6_outputs(6986));
    outputs(3242) <= not((layer6_outputs(3318)) xor (layer6_outputs(1314)));
    outputs(3243) <= layer6_outputs(1332);
    outputs(3244) <= not((layer6_outputs(4831)) xor (layer6_outputs(1011)));
    outputs(3245) <= not(layer6_outputs(241)) or (layer6_outputs(7459));
    outputs(3246) <= not((layer6_outputs(7632)) or (layer6_outputs(64)));
    outputs(3247) <= layer6_outputs(2947);
    outputs(3248) <= layer6_outputs(3766);
    outputs(3249) <= not(layer6_outputs(4407));
    outputs(3250) <= (layer6_outputs(2798)) xor (layer6_outputs(6037));
    outputs(3251) <= layer6_outputs(2033);
    outputs(3252) <= not((layer6_outputs(4438)) xor (layer6_outputs(958)));
    outputs(3253) <= layer6_outputs(785);
    outputs(3254) <= layer6_outputs(3138);
    outputs(3255) <= (layer6_outputs(5072)) and (layer6_outputs(3093));
    outputs(3256) <= not(layer6_outputs(7103));
    outputs(3257) <= not(layer6_outputs(895)) or (layer6_outputs(55));
    outputs(3258) <= (layer6_outputs(1920)) and not (layer6_outputs(3210));
    outputs(3259) <= (layer6_outputs(2508)) and (layer6_outputs(3652));
    outputs(3260) <= not(layer6_outputs(4584));
    outputs(3261) <= layer6_outputs(1386);
    outputs(3262) <= not(layer6_outputs(4872));
    outputs(3263) <= layer6_outputs(761);
    outputs(3264) <= layer6_outputs(6050);
    outputs(3265) <= (layer6_outputs(2195)) xor (layer6_outputs(6583));
    outputs(3266) <= (layer6_outputs(6672)) xor (layer6_outputs(4230));
    outputs(3267) <= layer6_outputs(546);
    outputs(3268) <= not(layer6_outputs(1816));
    outputs(3269) <= not(layer6_outputs(4472));
    outputs(3270) <= not(layer6_outputs(1337));
    outputs(3271) <= not(layer6_outputs(3458));
    outputs(3272) <= not(layer6_outputs(2733));
    outputs(3273) <= not(layer6_outputs(6290));
    outputs(3274) <= not(layer6_outputs(229));
    outputs(3275) <= not(layer6_outputs(6118));
    outputs(3276) <= layer6_outputs(2793);
    outputs(3277) <= not(layer6_outputs(1109));
    outputs(3278) <= not(layer6_outputs(1440));
    outputs(3279) <= (layer6_outputs(3351)) and (layer6_outputs(7276));
    outputs(3280) <= layer6_outputs(4213);
    outputs(3281) <= not(layer6_outputs(932));
    outputs(3282) <= (layer6_outputs(4998)) or (layer6_outputs(2233));
    outputs(3283) <= not((layer6_outputs(4176)) or (layer6_outputs(6007)));
    outputs(3284) <= (layer6_outputs(4806)) xor (layer6_outputs(3202));
    outputs(3285) <= not(layer6_outputs(6134));
    outputs(3286) <= (layer6_outputs(554)) xor (layer6_outputs(2106));
    outputs(3287) <= not((layer6_outputs(6816)) xor (layer6_outputs(2937)));
    outputs(3288) <= not((layer6_outputs(503)) xor (layer6_outputs(1912)));
    outputs(3289) <= not(layer6_outputs(7487));
    outputs(3290) <= layer6_outputs(5549);
    outputs(3291) <= (layer6_outputs(3489)) and not (layer6_outputs(1359));
    outputs(3292) <= layer6_outputs(1512);
    outputs(3293) <= (layer6_outputs(4158)) xor (layer6_outputs(7673));
    outputs(3294) <= (layer6_outputs(5877)) xor (layer6_outputs(3561));
    outputs(3295) <= layer6_outputs(4441);
    outputs(3296) <= not(layer6_outputs(7218));
    outputs(3297) <= not(layer6_outputs(7421));
    outputs(3298) <= not(layer6_outputs(3209));
    outputs(3299) <= layer6_outputs(1911);
    outputs(3300) <= (layer6_outputs(3161)) xor (layer6_outputs(417));
    outputs(3301) <= not(layer6_outputs(4350));
    outputs(3302) <= layer6_outputs(4179);
    outputs(3303) <= not((layer6_outputs(6058)) xor (layer6_outputs(6609)));
    outputs(3304) <= layer6_outputs(6225);
    outputs(3305) <= layer6_outputs(3904);
    outputs(3306) <= not(layer6_outputs(3435)) or (layer6_outputs(2890));
    outputs(3307) <= not(layer6_outputs(5969));
    outputs(3308) <= (layer6_outputs(6830)) xor (layer6_outputs(323));
    outputs(3309) <= layer6_outputs(1452);
    outputs(3310) <= not(layer6_outputs(1021));
    outputs(3311) <= (layer6_outputs(4994)) and not (layer6_outputs(4097));
    outputs(3312) <= (layer6_outputs(4597)) and (layer6_outputs(477));
    outputs(3313) <= not(layer6_outputs(2715));
    outputs(3314) <= (layer6_outputs(7541)) xor (layer6_outputs(3720));
    outputs(3315) <= layer6_outputs(7072);
    outputs(3316) <= (layer6_outputs(1251)) or (layer6_outputs(7410));
    outputs(3317) <= not(layer6_outputs(5386)) or (layer6_outputs(1620));
    outputs(3318) <= not(layer6_outputs(892));
    outputs(3319) <= not((layer6_outputs(6184)) xor (layer6_outputs(5862)));
    outputs(3320) <= layer6_outputs(4750);
    outputs(3321) <= (layer6_outputs(4135)) xor (layer6_outputs(6558));
    outputs(3322) <= (layer6_outputs(2011)) and (layer6_outputs(1027));
    outputs(3323) <= (layer6_outputs(7022)) or (layer6_outputs(4050));
    outputs(3324) <= layer6_outputs(4743);
    outputs(3325) <= not(layer6_outputs(3226));
    outputs(3326) <= (layer6_outputs(3329)) xor (layer6_outputs(79));
    outputs(3327) <= not(layer6_outputs(741));
    outputs(3328) <= layer6_outputs(7087);
    outputs(3329) <= not((layer6_outputs(5823)) xor (layer6_outputs(332)));
    outputs(3330) <= (layer6_outputs(2068)) and (layer6_outputs(5767));
    outputs(3331) <= (layer6_outputs(2814)) xor (layer6_outputs(3808));
    outputs(3332) <= not(layer6_outputs(7347));
    outputs(3333) <= not(layer6_outputs(7630));
    outputs(3334) <= layer6_outputs(360);
    outputs(3335) <= (layer6_outputs(5625)) and not (layer6_outputs(1365));
    outputs(3336) <= not((layer6_outputs(2915)) xor (layer6_outputs(5226)));
    outputs(3337) <= layer6_outputs(7312);
    outputs(3338) <= layer6_outputs(5136);
    outputs(3339) <= layer6_outputs(1619);
    outputs(3340) <= layer6_outputs(4067);
    outputs(3341) <= not(layer6_outputs(6072));
    outputs(3342) <= layer6_outputs(2937);
    outputs(3343) <= not(layer6_outputs(741)) or (layer6_outputs(3874));
    outputs(3344) <= (layer6_outputs(5585)) xor (layer6_outputs(6598));
    outputs(3345) <= (layer6_outputs(833)) and (layer6_outputs(5482));
    outputs(3346) <= (layer6_outputs(4165)) xor (layer6_outputs(6666));
    outputs(3347) <= layer6_outputs(2408);
    outputs(3348) <= layer6_outputs(493);
    outputs(3349) <= not(layer6_outputs(7331));
    outputs(3350) <= not(layer6_outputs(3882)) or (layer6_outputs(4495));
    outputs(3351) <= not((layer6_outputs(4364)) xor (layer6_outputs(7464)));
    outputs(3352) <= layer6_outputs(1062);
    outputs(3353) <= (layer6_outputs(2668)) xor (layer6_outputs(4782));
    outputs(3354) <= layer6_outputs(6016);
    outputs(3355) <= not(layer6_outputs(1938));
    outputs(3356) <= not(layer6_outputs(2866));
    outputs(3357) <= not(layer6_outputs(3606));
    outputs(3358) <= (layer6_outputs(5304)) xor (layer6_outputs(5506));
    outputs(3359) <= (layer6_outputs(381)) xor (layer6_outputs(4460));
    outputs(3360) <= not(layer6_outputs(6796));
    outputs(3361) <= not((layer6_outputs(2743)) xor (layer6_outputs(3012)));
    outputs(3362) <= layer6_outputs(6953);
    outputs(3363) <= not((layer6_outputs(671)) xor (layer6_outputs(2916)));
    outputs(3364) <= layer6_outputs(6485);
    outputs(3365) <= layer6_outputs(6521);
    outputs(3366) <= not((layer6_outputs(555)) or (layer6_outputs(1874)));
    outputs(3367) <= not(layer6_outputs(687));
    outputs(3368) <= layer6_outputs(1429);
    outputs(3369) <= not(layer6_outputs(1274));
    outputs(3370) <= not((layer6_outputs(7051)) xor (layer6_outputs(3797)));
    outputs(3371) <= not(layer6_outputs(2595));
    outputs(3372) <= not(layer6_outputs(300)) or (layer6_outputs(2051));
    outputs(3373) <= layer6_outputs(913);
    outputs(3374) <= layer6_outputs(5539);
    outputs(3375) <= not(layer6_outputs(3935));
    outputs(3376) <= not(layer6_outputs(2267));
    outputs(3377) <= not(layer6_outputs(4282)) or (layer6_outputs(4721));
    outputs(3378) <= not(layer6_outputs(1149));
    outputs(3379) <= layer6_outputs(161);
    outputs(3380) <= layer6_outputs(2944);
    outputs(3381) <= not(layer6_outputs(5206));
    outputs(3382) <= not(layer6_outputs(2640));
    outputs(3383) <= not(layer6_outputs(1354));
    outputs(3384) <= not(layer6_outputs(860));
    outputs(3385) <= layer6_outputs(5274);
    outputs(3386) <= not(layer6_outputs(5532)) or (layer6_outputs(247));
    outputs(3387) <= layer6_outputs(6205);
    outputs(3388) <= layer6_outputs(928);
    outputs(3389) <= (layer6_outputs(6786)) and (layer6_outputs(2165));
    outputs(3390) <= (layer6_outputs(5394)) xor (layer6_outputs(1323));
    outputs(3391) <= layer6_outputs(7591);
    outputs(3392) <= not(layer6_outputs(351));
    outputs(3393) <= layer6_outputs(6266);
    outputs(3394) <= layer6_outputs(1470);
    outputs(3395) <= (layer6_outputs(7283)) and (layer6_outputs(7449));
    outputs(3396) <= (layer6_outputs(1725)) and (layer6_outputs(6782));
    outputs(3397) <= not(layer6_outputs(5452));
    outputs(3398) <= not((layer6_outputs(6800)) and (layer6_outputs(4448)));
    outputs(3399) <= (layer6_outputs(3383)) xor (layer6_outputs(3258));
    outputs(3400) <= (layer6_outputs(2610)) xor (layer6_outputs(2604));
    outputs(3401) <= layer6_outputs(345);
    outputs(3402) <= not(layer6_outputs(5622));
    outputs(3403) <= not(layer6_outputs(3419));
    outputs(3404) <= not(layer6_outputs(6986));
    outputs(3405) <= not(layer6_outputs(7160));
    outputs(3406) <= not(layer6_outputs(6797));
    outputs(3407) <= not(layer6_outputs(5353));
    outputs(3408) <= layer6_outputs(5638);
    outputs(3409) <= (layer6_outputs(4899)) xor (layer6_outputs(1627));
    outputs(3410) <= not((layer6_outputs(4625)) xor (layer6_outputs(1766)));
    outputs(3411) <= (layer6_outputs(2522)) and not (layer6_outputs(2387));
    outputs(3412) <= not((layer6_outputs(3824)) xor (layer6_outputs(2151)));
    outputs(3413) <= not(layer6_outputs(2368));
    outputs(3414) <= not(layer6_outputs(625));
    outputs(3415) <= (layer6_outputs(7258)) and not (layer6_outputs(5924));
    outputs(3416) <= not(layer6_outputs(6206));
    outputs(3417) <= layer6_outputs(2840);
    outputs(3418) <= layer6_outputs(4992);
    outputs(3419) <= layer6_outputs(87);
    outputs(3420) <= layer6_outputs(5324);
    outputs(3421) <= not(layer6_outputs(2229));
    outputs(3422) <= layer6_outputs(6062);
    outputs(3423) <= layer6_outputs(3537);
    outputs(3424) <= not(layer6_outputs(2641));
    outputs(3425) <= layer6_outputs(5569);
    outputs(3426) <= layer6_outputs(6991);
    outputs(3427) <= not((layer6_outputs(6196)) xor (layer6_outputs(1230)));
    outputs(3428) <= not((layer6_outputs(5337)) xor (layer6_outputs(3160)));
    outputs(3429) <= not((layer6_outputs(2002)) or (layer6_outputs(1702)));
    outputs(3430) <= not(layer6_outputs(2319));
    outputs(3431) <= layer6_outputs(1727);
    outputs(3432) <= not((layer6_outputs(4508)) xor (layer6_outputs(1504)));
    outputs(3433) <= (layer6_outputs(2013)) xor (layer6_outputs(3814));
    outputs(3434) <= (layer6_outputs(4137)) and not (layer6_outputs(4411));
    outputs(3435) <= not(layer6_outputs(3735));
    outputs(3436) <= not((layer6_outputs(1863)) or (layer6_outputs(6391)));
    outputs(3437) <= not((layer6_outputs(6209)) xor (layer6_outputs(3694)));
    outputs(3438) <= not(layer6_outputs(7054));
    outputs(3439) <= layer6_outputs(5239);
    outputs(3440) <= (layer6_outputs(122)) xor (layer6_outputs(5152));
    outputs(3441) <= layer6_outputs(3567);
    outputs(3442) <= layer6_outputs(7176);
    outputs(3443) <= layer6_outputs(6166);
    outputs(3444) <= layer6_outputs(658);
    outputs(3445) <= not(layer6_outputs(3931));
    outputs(3446) <= not(layer6_outputs(6897)) or (layer6_outputs(3084));
    outputs(3447) <= (layer6_outputs(6826)) and not (layer6_outputs(5790));
    outputs(3448) <= not(layer6_outputs(6699));
    outputs(3449) <= not((layer6_outputs(3186)) xor (layer6_outputs(3682)));
    outputs(3450) <= not((layer6_outputs(2114)) xor (layer6_outputs(3867)));
    outputs(3451) <= not(layer6_outputs(3370));
    outputs(3452) <= not(layer6_outputs(7622));
    outputs(3453) <= layer6_outputs(6203);
    outputs(3454) <= layer6_outputs(4352);
    outputs(3455) <= layer6_outputs(546);
    outputs(3456) <= not(layer6_outputs(5706));
    outputs(3457) <= not(layer6_outputs(3063));
    outputs(3458) <= layer6_outputs(2103);
    outputs(3459) <= (layer6_outputs(7528)) or (layer6_outputs(5602));
    outputs(3460) <= not(layer6_outputs(6665));
    outputs(3461) <= (layer6_outputs(4755)) and (layer6_outputs(1211));
    outputs(3462) <= layer6_outputs(4928);
    outputs(3463) <= not(layer6_outputs(4403));
    outputs(3464) <= not((layer6_outputs(6749)) xor (layer6_outputs(2296)));
    outputs(3465) <= not(layer6_outputs(2007));
    outputs(3466) <= (layer6_outputs(1363)) and not (layer6_outputs(5702));
    outputs(3467) <= (layer6_outputs(7052)) or (layer6_outputs(3572));
    outputs(3468) <= layer6_outputs(3434);
    outputs(3469) <= not(layer6_outputs(6098));
    outputs(3470) <= (layer6_outputs(6149)) xor (layer6_outputs(5228));
    outputs(3471) <= not(layer6_outputs(6715));
    outputs(3472) <= not(layer6_outputs(25));
    outputs(3473) <= not((layer6_outputs(7118)) or (layer6_outputs(4497)));
    outputs(3474) <= not(layer6_outputs(4004));
    outputs(3475) <= layer6_outputs(2172);
    outputs(3476) <= layer6_outputs(3148);
    outputs(3477) <= layer6_outputs(5161);
    outputs(3478) <= not(layer6_outputs(1040));
    outputs(3479) <= not(layer6_outputs(4161));
    outputs(3480) <= layer6_outputs(511);
    outputs(3481) <= not(layer6_outputs(2276));
    outputs(3482) <= not(layer6_outputs(7483));
    outputs(3483) <= (layer6_outputs(1587)) and not (layer6_outputs(1412));
    outputs(3484) <= layer6_outputs(3675);
    outputs(3485) <= not((layer6_outputs(256)) xor (layer6_outputs(6499)));
    outputs(3486) <= (layer6_outputs(30)) or (layer6_outputs(5947));
    outputs(3487) <= not((layer6_outputs(7563)) xor (layer6_outputs(6734)));
    outputs(3488) <= layer6_outputs(4371);
    outputs(3489) <= not(layer6_outputs(5180)) or (layer6_outputs(169));
    outputs(3490) <= (layer6_outputs(1100)) and not (layer6_outputs(1489));
    outputs(3491) <= not(layer6_outputs(4889));
    outputs(3492) <= layer6_outputs(3297);
    outputs(3493) <= (layer6_outputs(7363)) xor (layer6_outputs(1551));
    outputs(3494) <= layer6_outputs(4533);
    outputs(3495) <= (layer6_outputs(3432)) xor (layer6_outputs(238));
    outputs(3496) <= layer6_outputs(1707);
    outputs(3497) <= (layer6_outputs(2608)) xor (layer6_outputs(1457));
    outputs(3498) <= not((layer6_outputs(3091)) xor (layer6_outputs(5346)));
    outputs(3499) <= not((layer6_outputs(6360)) or (layer6_outputs(1473)));
    outputs(3500) <= not(layer6_outputs(6899));
    outputs(3501) <= not(layer6_outputs(650));
    outputs(3502) <= not((layer6_outputs(4798)) xor (layer6_outputs(7195)));
    outputs(3503) <= not((layer6_outputs(6218)) xor (layer6_outputs(7577)));
    outputs(3504) <= not((layer6_outputs(4205)) and (layer6_outputs(5780)));
    outputs(3505) <= not(layer6_outputs(3347));
    outputs(3506) <= (layer6_outputs(3836)) or (layer6_outputs(5404));
    outputs(3507) <= layer6_outputs(4869);
    outputs(3508) <= not((layer6_outputs(7050)) xor (layer6_outputs(4933)));
    outputs(3509) <= layer6_outputs(7012);
    outputs(3510) <= not(layer6_outputs(5702));
    outputs(3511) <= not(layer6_outputs(6320));
    outputs(3512) <= layer6_outputs(4080);
    outputs(3513) <= (layer6_outputs(1950)) xor (layer6_outputs(789));
    outputs(3514) <= not((layer6_outputs(4086)) or (layer6_outputs(3042)));
    outputs(3515) <= layer6_outputs(4211);
    outputs(3516) <= not(layer6_outputs(6840));
    outputs(3517) <= (layer6_outputs(2982)) xor (layer6_outputs(3555));
    outputs(3518) <= layer6_outputs(7426);
    outputs(3519) <= layer6_outputs(1922);
    outputs(3520) <= (layer6_outputs(2280)) xor (layer6_outputs(3671));
    outputs(3521) <= layer6_outputs(1913);
    outputs(3522) <= not(layer6_outputs(1130));
    outputs(3523) <= layer6_outputs(3491);
    outputs(3524) <= layer6_outputs(3372);
    outputs(3525) <= layer6_outputs(3896);
    outputs(3526) <= not((layer6_outputs(4924)) xor (layer6_outputs(3705)));
    outputs(3527) <= (layer6_outputs(1967)) or (layer6_outputs(3706));
    outputs(3528) <= not(layer6_outputs(1));
    outputs(3529) <= not(layer6_outputs(1844));
    outputs(3530) <= layer6_outputs(6106);
    outputs(3531) <= not((layer6_outputs(7156)) xor (layer6_outputs(3139)));
    outputs(3532) <= not(layer6_outputs(1030));
    outputs(3533) <= layer6_outputs(4639);
    outputs(3534) <= layer6_outputs(234);
    outputs(3535) <= layer6_outputs(2088);
    outputs(3536) <= layer6_outputs(1721);
    outputs(3537) <= not((layer6_outputs(5327)) xor (layer6_outputs(111)));
    outputs(3538) <= not(layer6_outputs(1401));
    outputs(3539) <= not((layer6_outputs(288)) and (layer6_outputs(3193)));
    outputs(3540) <= layer6_outputs(1096);
    outputs(3541) <= (layer6_outputs(2271)) xor (layer6_outputs(3029));
    outputs(3542) <= not(layer6_outputs(2179));
    outputs(3543) <= (layer6_outputs(5889)) or (layer6_outputs(7400));
    outputs(3544) <= layer6_outputs(6977);
    outputs(3545) <= not(layer6_outputs(5276));
    outputs(3546) <= layer6_outputs(4666);
    outputs(3547) <= not(layer6_outputs(4762));
    outputs(3548) <= not(layer6_outputs(4823));
    outputs(3549) <= layer6_outputs(3779);
    outputs(3550) <= layer6_outputs(4594);
    outputs(3551) <= not((layer6_outputs(5291)) xor (layer6_outputs(5713)));
    outputs(3552) <= not(layer6_outputs(730));
    outputs(3553) <= not(layer6_outputs(6649));
    outputs(3554) <= (layer6_outputs(5647)) xor (layer6_outputs(1930));
    outputs(3555) <= not(layer6_outputs(5176));
    outputs(3556) <= not((layer6_outputs(7415)) xor (layer6_outputs(3174)));
    outputs(3557) <= not(layer6_outputs(5055));
    outputs(3558) <= layer6_outputs(4531);
    outputs(3559) <= (layer6_outputs(6451)) xor (layer6_outputs(6798));
    outputs(3560) <= (layer6_outputs(1295)) and not (layer6_outputs(6169));
    outputs(3561) <= (layer6_outputs(3620)) and not (layer6_outputs(4395));
    outputs(3562) <= (layer6_outputs(5618)) xor (layer6_outputs(1340));
    outputs(3563) <= not((layer6_outputs(3641)) xor (layer6_outputs(6460)));
    outputs(3564) <= not(layer6_outputs(6346));
    outputs(3565) <= not(layer6_outputs(2086));
    outputs(3566) <= not(layer6_outputs(3589));
    outputs(3567) <= (layer6_outputs(4601)) xor (layer6_outputs(4355));
    outputs(3568) <= layer6_outputs(5343);
    outputs(3569) <= layer6_outputs(2564);
    outputs(3570) <= layer6_outputs(4457);
    outputs(3571) <= layer6_outputs(281);
    outputs(3572) <= (layer6_outputs(947)) xor (layer6_outputs(7241));
    outputs(3573) <= layer6_outputs(2044);
    outputs(3574) <= layer6_outputs(3966);
    outputs(3575) <= layer6_outputs(7671);
    outputs(3576) <= (layer6_outputs(137)) and (layer6_outputs(1559));
    outputs(3577) <= not(layer6_outputs(4520));
    outputs(3578) <= layer6_outputs(2443);
    outputs(3579) <= not((layer6_outputs(3690)) xor (layer6_outputs(4697)));
    outputs(3580) <= not((layer6_outputs(5234)) xor (layer6_outputs(3481)));
    outputs(3581) <= layer6_outputs(3031);
    outputs(3582) <= layer6_outputs(2695);
    outputs(3583) <= not(layer6_outputs(4587));
    outputs(3584) <= not(layer6_outputs(6430));
    outputs(3585) <= not((layer6_outputs(3570)) xor (layer6_outputs(1812)));
    outputs(3586) <= layer6_outputs(7274);
    outputs(3587) <= (layer6_outputs(2051)) or (layer6_outputs(5619));
    outputs(3588) <= layer6_outputs(5689);
    outputs(3589) <= (layer6_outputs(1448)) xor (layer6_outputs(7407));
    outputs(3590) <= layer6_outputs(2519);
    outputs(3591) <= layer6_outputs(743);
    outputs(3592) <= (layer6_outputs(3771)) xor (layer6_outputs(5217));
    outputs(3593) <= layer6_outputs(3402);
    outputs(3594) <= not(layer6_outputs(6928));
    outputs(3595) <= not(layer6_outputs(4129));
    outputs(3596) <= not(layer6_outputs(2547));
    outputs(3597) <= (layer6_outputs(1862)) and not (layer6_outputs(6350));
    outputs(3598) <= layer6_outputs(1959);
    outputs(3599) <= layer6_outputs(3501);
    outputs(3600) <= layer6_outputs(1602);
    outputs(3601) <= layer6_outputs(4191);
    outputs(3602) <= layer6_outputs(2064);
    outputs(3603) <= layer6_outputs(3745);
    outputs(3604) <= not(layer6_outputs(393));
    outputs(3605) <= layer6_outputs(5110);
    outputs(3606) <= layer6_outputs(6907);
    outputs(3607) <= not(layer6_outputs(5417));
    outputs(3608) <= not(layer6_outputs(158));
    outputs(3609) <= layer6_outputs(7251);
    outputs(3610) <= layer6_outputs(3627);
    outputs(3611) <= (layer6_outputs(737)) xor (layer6_outputs(122));
    outputs(3612) <= layer6_outputs(3581);
    outputs(3613) <= layer6_outputs(5732);
    outputs(3614) <= layer6_outputs(7148);
    outputs(3615) <= layer6_outputs(4603);
    outputs(3616) <= layer6_outputs(2749);
    outputs(3617) <= not(layer6_outputs(1421));
    outputs(3618) <= not(layer6_outputs(3410));
    outputs(3619) <= layer6_outputs(3498);
    outputs(3620) <= layer6_outputs(5645);
    outputs(3621) <= not(layer6_outputs(25));
    outputs(3622) <= not(layer6_outputs(263));
    outputs(3623) <= not((layer6_outputs(5438)) and (layer6_outputs(2965)));
    outputs(3624) <= not(layer6_outputs(5181));
    outputs(3625) <= not(layer6_outputs(4887));
    outputs(3626) <= (layer6_outputs(5031)) and not (layer6_outputs(1872));
    outputs(3627) <= not(layer6_outputs(436));
    outputs(3628) <= not(layer6_outputs(7654)) or (layer6_outputs(1472));
    outputs(3629) <= not(layer6_outputs(2687));
    outputs(3630) <= layer6_outputs(6326);
    outputs(3631) <= layer6_outputs(7540);
    outputs(3632) <= layer6_outputs(4869);
    outputs(3633) <= not(layer6_outputs(949));
    outputs(3634) <= (layer6_outputs(4658)) xor (layer6_outputs(3181));
    outputs(3635) <= not(layer6_outputs(4277));
    outputs(3636) <= (layer6_outputs(715)) xor (layer6_outputs(448));
    outputs(3637) <= not((layer6_outputs(5259)) xor (layer6_outputs(7236)));
    outputs(3638) <= not(layer6_outputs(5477));
    outputs(3639) <= layer6_outputs(2901);
    outputs(3640) <= not(layer6_outputs(1261));
    outputs(3641) <= not((layer6_outputs(1801)) xor (layer6_outputs(4577)));
    outputs(3642) <= not(layer6_outputs(1891));
    outputs(3643) <= layer6_outputs(83);
    outputs(3644) <= layer6_outputs(2955);
    outputs(3645) <= layer6_outputs(3242);
    outputs(3646) <= not(layer6_outputs(2054));
    outputs(3647) <= not((layer6_outputs(1310)) xor (layer6_outputs(1879)));
    outputs(3648) <= (layer6_outputs(3850)) xor (layer6_outputs(4841));
    outputs(3649) <= not(layer6_outputs(6615));
    outputs(3650) <= not((layer6_outputs(3918)) xor (layer6_outputs(6851)));
    outputs(3651) <= (layer6_outputs(5462)) xor (layer6_outputs(2005));
    outputs(3652) <= not((layer6_outputs(965)) xor (layer6_outputs(3951)));
    outputs(3653) <= layer6_outputs(6910);
    outputs(3654) <= layer6_outputs(2460);
    outputs(3655) <= not((layer6_outputs(4157)) or (layer6_outputs(2073)));
    outputs(3656) <= not(layer6_outputs(5028));
    outputs(3657) <= not(layer6_outputs(953));
    outputs(3658) <= not(layer6_outputs(1150));
    outputs(3659) <= not(layer6_outputs(6852));
    outputs(3660) <= layer6_outputs(5569);
    outputs(3661) <= not((layer6_outputs(5592)) xor (layer6_outputs(185)));
    outputs(3662) <= not(layer6_outputs(4250));
    outputs(3663) <= not((layer6_outputs(533)) xor (layer6_outputs(5547)));
    outputs(3664) <= layer6_outputs(677);
    outputs(3665) <= not((layer6_outputs(6094)) xor (layer6_outputs(1580)));
    outputs(3666) <= not((layer6_outputs(5177)) or (layer6_outputs(3475)));
    outputs(3667) <= not((layer6_outputs(7089)) xor (layer6_outputs(5579)));
    outputs(3668) <= (layer6_outputs(750)) xor (layer6_outputs(7330));
    outputs(3669) <= not(layer6_outputs(3129));
    outputs(3670) <= (layer6_outputs(5046)) xor (layer6_outputs(7297));
    outputs(3671) <= (layer6_outputs(3477)) xor (layer6_outputs(2975));
    outputs(3672) <= not(layer6_outputs(7679));
    outputs(3673) <= not(layer6_outputs(6603));
    outputs(3674) <= (layer6_outputs(5341)) and not (layer6_outputs(2291));
    outputs(3675) <= not(layer6_outputs(5139)) or (layer6_outputs(7108));
    outputs(3676) <= not((layer6_outputs(6253)) xor (layer6_outputs(5204)));
    outputs(3677) <= not(layer6_outputs(1141));
    outputs(3678) <= layer6_outputs(3663);
    outputs(3679) <= layer6_outputs(1286);
    outputs(3680) <= not(layer6_outputs(5799));
    outputs(3681) <= (layer6_outputs(3734)) xor (layer6_outputs(6911));
    outputs(3682) <= not(layer6_outputs(5870));
    outputs(3683) <= not((layer6_outputs(2427)) and (layer6_outputs(7431)));
    outputs(3684) <= (layer6_outputs(4062)) xor (layer6_outputs(5275));
    outputs(3685) <= layer6_outputs(2599);
    outputs(3686) <= not((layer6_outputs(5469)) xor (layer6_outputs(2128)));
    outputs(3687) <= not(layer6_outputs(6226));
    outputs(3688) <= (layer6_outputs(4970)) xor (layer6_outputs(6977));
    outputs(3689) <= layer6_outputs(3693);
    outputs(3690) <= not(layer6_outputs(5438));
    outputs(3691) <= layer6_outputs(2920);
    outputs(3692) <= (layer6_outputs(1532)) and not (layer6_outputs(930));
    outputs(3693) <= (layer6_outputs(4061)) xor (layer6_outputs(6572));
    outputs(3694) <= not(layer6_outputs(3634));
    outputs(3695) <= layer6_outputs(7633);
    outputs(3696) <= not(layer6_outputs(4201));
    outputs(3697) <= (layer6_outputs(7018)) and not (layer6_outputs(6523));
    outputs(3698) <= not(layer6_outputs(2352)) or (layer6_outputs(480));
    outputs(3699) <= (layer6_outputs(2190)) and (layer6_outputs(6262));
    outputs(3700) <= (layer6_outputs(233)) xor (layer6_outputs(1213));
    outputs(3701) <= not(layer6_outputs(985));
    outputs(3702) <= (layer6_outputs(3156)) and not (layer6_outputs(5762));
    outputs(3703) <= not((layer6_outputs(3710)) xor (layer6_outputs(573)));
    outputs(3704) <= not(layer6_outputs(1447));
    outputs(3705) <= not(layer6_outputs(5252));
    outputs(3706) <= (layer6_outputs(7241)) xor (layer6_outputs(4111));
    outputs(3707) <= layer6_outputs(3490);
    outputs(3708) <= not(layer6_outputs(2863));
    outputs(3709) <= not(layer6_outputs(2152));
    outputs(3710) <= layer6_outputs(3948);
    outputs(3711) <= (layer6_outputs(1730)) xor (layer6_outputs(6359));
    outputs(3712) <= (layer6_outputs(7582)) or (layer6_outputs(740));
    outputs(3713) <= layer6_outputs(4728);
    outputs(3714) <= (layer6_outputs(6795)) xor (layer6_outputs(7379));
    outputs(3715) <= layer6_outputs(7158);
    outputs(3716) <= layer6_outputs(1707);
    outputs(3717) <= layer6_outputs(5578);
    outputs(3718) <= not((layer6_outputs(2693)) xor (layer6_outputs(4718)));
    outputs(3719) <= not(layer6_outputs(3428));
    outputs(3720) <= layer6_outputs(691);
    outputs(3721) <= (layer6_outputs(4454)) xor (layer6_outputs(541));
    outputs(3722) <= not(layer6_outputs(6248));
    outputs(3723) <= not(layer6_outputs(6454));
    outputs(3724) <= (layer6_outputs(4469)) or (layer6_outputs(1812));
    outputs(3725) <= not(layer6_outputs(6268));
    outputs(3726) <= (layer6_outputs(2695)) and not (layer6_outputs(519));
    outputs(3727) <= not(layer6_outputs(4698));
    outputs(3728) <= not(layer6_outputs(5930));
    outputs(3729) <= not((layer6_outputs(382)) or (layer6_outputs(6834)));
    outputs(3730) <= not(layer6_outputs(5147)) or (layer6_outputs(6337));
    outputs(3731) <= not((layer6_outputs(2285)) xor (layer6_outputs(6805)));
    outputs(3732) <= (layer6_outputs(2439)) xor (layer6_outputs(3863));
    outputs(3733) <= not(layer6_outputs(1720));
    outputs(3734) <= not(layer6_outputs(7620));
    outputs(3735) <= not((layer6_outputs(3824)) xor (layer6_outputs(4820)));
    outputs(3736) <= not(layer6_outputs(6010));
    outputs(3737) <= layer6_outputs(7354);
    outputs(3738) <= not(layer6_outputs(5850));
    outputs(3739) <= (layer6_outputs(7456)) xor (layer6_outputs(3714));
    outputs(3740) <= layer6_outputs(3811);
    outputs(3741) <= not(layer6_outputs(5230));
    outputs(3742) <= not(layer6_outputs(4714)) or (layer6_outputs(749));
    outputs(3743) <= not((layer6_outputs(1462)) xor (layer6_outputs(993)));
    outputs(3744) <= layer6_outputs(3527);
    outputs(3745) <= (layer6_outputs(7584)) and not (layer6_outputs(4000));
    outputs(3746) <= layer6_outputs(3663);
    outputs(3747) <= not((layer6_outputs(3898)) xor (layer6_outputs(884)));
    outputs(3748) <= layer6_outputs(1057);
    outputs(3749) <= not((layer6_outputs(1055)) xor (layer6_outputs(2441)));
    outputs(3750) <= (layer6_outputs(6054)) xor (layer6_outputs(1275));
    outputs(3751) <= (layer6_outputs(1489)) xor (layer6_outputs(6671));
    outputs(3752) <= layer6_outputs(7676);
    outputs(3753) <= (layer6_outputs(7119)) xor (layer6_outputs(2929));
    outputs(3754) <= not(layer6_outputs(6847));
    outputs(3755) <= (layer6_outputs(3336)) and not (layer6_outputs(6368));
    outputs(3756) <= not(layer6_outputs(4929));
    outputs(3757) <= layer6_outputs(4720);
    outputs(3758) <= layer6_outputs(5287);
    outputs(3759) <= not(layer6_outputs(6348));
    outputs(3760) <= not(layer6_outputs(6405));
    outputs(3761) <= not(layer6_outputs(7054));
    outputs(3762) <= not(layer6_outputs(7316));
    outputs(3763) <= not((layer6_outputs(5903)) xor (layer6_outputs(4048)));
    outputs(3764) <= layer6_outputs(4380);
    outputs(3765) <= not((layer6_outputs(3072)) xor (layer6_outputs(3014)));
    outputs(3766) <= layer6_outputs(1483);
    outputs(3767) <= layer6_outputs(587);
    outputs(3768) <= not(layer6_outputs(2276));
    outputs(3769) <= not(layer6_outputs(4218));
    outputs(3770) <= not(layer6_outputs(5855));
    outputs(3771) <= not((layer6_outputs(5220)) xor (layer6_outputs(6653)));
    outputs(3772) <= (layer6_outputs(1231)) and not (layer6_outputs(6025));
    outputs(3773) <= (layer6_outputs(3957)) xor (layer6_outputs(2963));
    outputs(3774) <= not(layer6_outputs(5050));
    outputs(3775) <= (layer6_outputs(2795)) xor (layer6_outputs(805));
    outputs(3776) <= layer6_outputs(4160);
    outputs(3777) <= not((layer6_outputs(5752)) xor (layer6_outputs(5496)));
    outputs(3778) <= layer6_outputs(1344);
    outputs(3779) <= layer6_outputs(131);
    outputs(3780) <= (layer6_outputs(874)) and (layer6_outputs(7385));
    outputs(3781) <= not(layer6_outputs(4813));
    outputs(3782) <= not(layer6_outputs(2991));
    outputs(3783) <= not(layer6_outputs(1624));
    outputs(3784) <= layer6_outputs(4228);
    outputs(3785) <= not(layer6_outputs(4941));
    outputs(3786) <= (layer6_outputs(57)) and not (layer6_outputs(1894));
    outputs(3787) <= layer6_outputs(252);
    outputs(3788) <= not((layer6_outputs(6258)) xor (layer6_outputs(6444)));
    outputs(3789) <= layer6_outputs(697);
    outputs(3790) <= not(layer6_outputs(6840));
    outputs(3791) <= (layer6_outputs(4661)) and not (layer6_outputs(5657));
    outputs(3792) <= layer6_outputs(5241);
    outputs(3793) <= layer6_outputs(6948);
    outputs(3794) <= layer6_outputs(6029);
    outputs(3795) <= layer6_outputs(2934);
    outputs(3796) <= (layer6_outputs(2889)) xor (layer6_outputs(2891));
    outputs(3797) <= layer6_outputs(1429);
    outputs(3798) <= layer6_outputs(1575);
    outputs(3799) <= not(layer6_outputs(4151));
    outputs(3800) <= not(layer6_outputs(1609));
    outputs(3801) <= (layer6_outputs(5190)) and not (layer6_outputs(7314));
    outputs(3802) <= not(layer6_outputs(2314));
    outputs(3803) <= not(layer6_outputs(320));
    outputs(3804) <= not(layer6_outputs(3384));
    outputs(3805) <= not((layer6_outputs(738)) xor (layer6_outputs(877)));
    outputs(3806) <= not((layer6_outputs(4012)) xor (layer6_outputs(7258)));
    outputs(3807) <= layer6_outputs(6047);
    outputs(3808) <= not((layer6_outputs(3886)) xor (layer6_outputs(1917)));
    outputs(3809) <= (layer6_outputs(572)) xor (layer6_outputs(3825));
    outputs(3810) <= not(layer6_outputs(7370));
    outputs(3811) <= layer6_outputs(1430);
    outputs(3812) <= (layer6_outputs(4267)) xor (layer6_outputs(118));
    outputs(3813) <= layer6_outputs(7000);
    outputs(3814) <= layer6_outputs(6655);
    outputs(3815) <= not(layer6_outputs(2014)) or (layer6_outputs(2835));
    outputs(3816) <= (layer6_outputs(3361)) and not (layer6_outputs(5284));
    outputs(3817) <= layer6_outputs(3058);
    outputs(3818) <= layer6_outputs(2194);
    outputs(3819) <= not(layer6_outputs(2288));
    outputs(3820) <= layer6_outputs(3496);
    outputs(3821) <= not(layer6_outputs(6366));
    outputs(3822) <= not(layer6_outputs(6199));
    outputs(3823) <= (layer6_outputs(6694)) and (layer6_outputs(5531));
    outputs(3824) <= not(layer6_outputs(4890));
    outputs(3825) <= not(layer6_outputs(5277));
    outputs(3826) <= layer6_outputs(4983);
    outputs(3827) <= (layer6_outputs(2135)) xor (layer6_outputs(7238));
    outputs(3828) <= not(layer6_outputs(664));
    outputs(3829) <= (layer6_outputs(66)) and not (layer6_outputs(3920));
    outputs(3830) <= not(layer6_outputs(990));
    outputs(3831) <= (layer6_outputs(5430)) xor (layer6_outputs(5779));
    outputs(3832) <= not(layer6_outputs(112));
    outputs(3833) <= layer6_outputs(950);
    outputs(3834) <= (layer6_outputs(432)) xor (layer6_outputs(1983));
    outputs(3835) <= layer6_outputs(1349);
    outputs(3836) <= not(layer6_outputs(3971));
    outputs(3837) <= not((layer6_outputs(2846)) and (layer6_outputs(306)));
    outputs(3838) <= layer6_outputs(4526);
    outputs(3839) <= not(layer6_outputs(2259));
    outputs(3840) <= layer6_outputs(7210);
    outputs(3841) <= not(layer6_outputs(6758));
    outputs(3842) <= layer6_outputs(1799);
    outputs(3843) <= (layer6_outputs(3285)) xor (layer6_outputs(3780));
    outputs(3844) <= not(layer6_outputs(4293));
    outputs(3845) <= (layer6_outputs(6883)) xor (layer6_outputs(4139));
    outputs(3846) <= not(layer6_outputs(7666));
    outputs(3847) <= not(layer6_outputs(3396));
    outputs(3848) <= layer6_outputs(726);
    outputs(3849) <= (layer6_outputs(6316)) xor (layer6_outputs(249));
    outputs(3850) <= layer6_outputs(6739);
    outputs(3851) <= not(layer6_outputs(7314));
    outputs(3852) <= not(layer6_outputs(4679));
    outputs(3853) <= layer6_outputs(7113);
    outputs(3854) <= (layer6_outputs(6997)) and not (layer6_outputs(374));
    outputs(3855) <= (layer6_outputs(2119)) xor (layer6_outputs(4074));
    outputs(3856) <= not(layer6_outputs(3296));
    outputs(3857) <= not((layer6_outputs(7498)) xor (layer6_outputs(6980)));
    outputs(3858) <= layer6_outputs(4939);
    outputs(3859) <= not(layer6_outputs(2938));
    outputs(3860) <= layer6_outputs(3607);
    outputs(3861) <= layer6_outputs(2673);
    outputs(3862) <= not((layer6_outputs(4835)) xor (layer6_outputs(6440)));
    outputs(3863) <= (layer6_outputs(1715)) and not (layer6_outputs(1986));
    outputs(3864) <= not(layer6_outputs(837)) or (layer6_outputs(4406));
    outputs(3865) <= (layer6_outputs(498)) or (layer6_outputs(681));
    outputs(3866) <= not(layer6_outputs(993));
    outputs(3867) <= layer6_outputs(6311);
    outputs(3868) <= layer6_outputs(4277);
    outputs(3869) <= layer6_outputs(792);
    outputs(3870) <= not((layer6_outputs(3985)) xor (layer6_outputs(3420)));
    outputs(3871) <= not(layer6_outputs(6823));
    outputs(3872) <= layer6_outputs(849);
    outputs(3873) <= (layer6_outputs(6216)) and not (layer6_outputs(438));
    outputs(3874) <= (layer6_outputs(6295)) or (layer6_outputs(7554));
    outputs(3875) <= (layer6_outputs(7432)) xor (layer6_outputs(4015));
    outputs(3876) <= (layer6_outputs(3912)) or (layer6_outputs(7201));
    outputs(3877) <= not(layer6_outputs(4795));
    outputs(3878) <= not(layer6_outputs(7623));
    outputs(3879) <= layer6_outputs(4940);
    outputs(3880) <= not(layer6_outputs(4332)) or (layer6_outputs(3062));
    outputs(3881) <= layer6_outputs(889);
    outputs(3882) <= (layer6_outputs(3302)) xor (layer6_outputs(5681));
    outputs(3883) <= (layer6_outputs(4002)) xor (layer6_outputs(5209));
    outputs(3884) <= not(layer6_outputs(3142));
    outputs(3885) <= not(layer6_outputs(2355));
    outputs(3886) <= (layer6_outputs(1154)) xor (layer6_outputs(6643));
    outputs(3887) <= layer6_outputs(3361);
    outputs(3888) <= not(layer6_outputs(283)) or (layer6_outputs(2588));
    outputs(3889) <= not(layer6_outputs(3001));
    outputs(3890) <= not((layer6_outputs(6549)) xor (layer6_outputs(2798)));
    outputs(3891) <= not(layer6_outputs(1061));
    outputs(3892) <= not((layer6_outputs(1556)) xor (layer6_outputs(2067)));
    outputs(3893) <= not((layer6_outputs(5102)) xor (layer6_outputs(6793)));
    outputs(3894) <= (layer6_outputs(831)) xor (layer6_outputs(6291));
    outputs(3895) <= not(layer6_outputs(5134));
    outputs(3896) <= (layer6_outputs(568)) xor (layer6_outputs(3072));
    outputs(3897) <= (layer6_outputs(1802)) xor (layer6_outputs(7286));
    outputs(3898) <= layer6_outputs(6576);
    outputs(3899) <= not(layer6_outputs(3719));
    outputs(3900) <= not((layer6_outputs(6717)) xor (layer6_outputs(5784)));
    outputs(3901) <= not(layer6_outputs(5387));
    outputs(3902) <= (layer6_outputs(4719)) xor (layer6_outputs(3769));
    outputs(3903) <= not(layer6_outputs(1710));
    outputs(3904) <= (layer6_outputs(3077)) xor (layer6_outputs(6157));
    outputs(3905) <= layer6_outputs(2753);
    outputs(3906) <= not(layer6_outputs(801));
    outputs(3907) <= (layer6_outputs(7333)) xor (layer6_outputs(6230));
    outputs(3908) <= (layer6_outputs(1919)) xor (layer6_outputs(3479));
    outputs(3909) <= layer6_outputs(703);
    outputs(3910) <= layer6_outputs(405);
    outputs(3911) <= not(layer6_outputs(845));
    outputs(3912) <= not(layer6_outputs(1164));
    outputs(3913) <= not((layer6_outputs(1653)) xor (layer6_outputs(6895)));
    outputs(3914) <= not((layer6_outputs(6533)) xor (layer6_outputs(7646)));
    outputs(3915) <= not(layer6_outputs(3503));
    outputs(3916) <= not(layer6_outputs(1233));
    outputs(3917) <= not(layer6_outputs(5225));
    outputs(3918) <= (layer6_outputs(7282)) xor (layer6_outputs(1026));
    outputs(3919) <= (layer6_outputs(4818)) or (layer6_outputs(5057));
    outputs(3920) <= not(layer6_outputs(5690));
    outputs(3921) <= (layer6_outputs(5572)) xor (layer6_outputs(6887));
    outputs(3922) <= not(layer6_outputs(5701));
    outputs(3923) <= not(layer6_outputs(4904));
    outputs(3924) <= not(layer6_outputs(6913));
    outputs(3925) <= (layer6_outputs(4143)) xor (layer6_outputs(1443));
    outputs(3926) <= not(layer6_outputs(6781));
    outputs(3927) <= layer6_outputs(3741);
    outputs(3928) <= not(layer6_outputs(7111));
    outputs(3929) <= layer6_outputs(7443);
    outputs(3930) <= (layer6_outputs(893)) and not (layer6_outputs(6667));
    outputs(3931) <= not(layer6_outputs(2316));
    outputs(3932) <= not(layer6_outputs(1594)) or (layer6_outputs(4641));
    outputs(3933) <= not(layer6_outputs(5148));
    outputs(3934) <= not(layer6_outputs(3162));
    outputs(3935) <= (layer6_outputs(3171)) and not (layer6_outputs(4942));
    outputs(3936) <= not(layer6_outputs(4677));
    outputs(3937) <= not(layer6_outputs(7621)) or (layer6_outputs(7086));
    outputs(3938) <= not(layer6_outputs(2805));
    outputs(3939) <= (layer6_outputs(3643)) xor (layer6_outputs(232));
    outputs(3940) <= (layer6_outputs(3666)) xor (layer6_outputs(284));
    outputs(3941) <= not((layer6_outputs(6842)) xor (layer6_outputs(3713)));
    outputs(3942) <= not((layer6_outputs(4824)) xor (layer6_outputs(3958)));
    outputs(3943) <= (layer6_outputs(5931)) xor (layer6_outputs(4300));
    outputs(3944) <= (layer6_outputs(4081)) xor (layer6_outputs(4908));
    outputs(3945) <= not((layer6_outputs(1409)) xor (layer6_outputs(3575)));
    outputs(3946) <= not((layer6_outputs(4809)) and (layer6_outputs(1916)));
    outputs(3947) <= (layer6_outputs(4636)) xor (layer6_outputs(348));
    outputs(3948) <= not((layer6_outputs(1864)) or (layer6_outputs(5290)));
    outputs(3949) <= (layer6_outputs(5476)) and not (layer6_outputs(3869));
    outputs(3950) <= (layer6_outputs(4365)) xor (layer6_outputs(428));
    outputs(3951) <= (layer6_outputs(4031)) and not (layer6_outputs(5258));
    outputs(3952) <= not((layer6_outputs(899)) xor (layer6_outputs(4861)));
    outputs(3953) <= layer6_outputs(7571);
    outputs(3954) <= (layer6_outputs(5825)) and (layer6_outputs(710));
    outputs(3955) <= (layer6_outputs(7607)) xor (layer6_outputs(471));
    outputs(3956) <= not((layer6_outputs(2403)) xor (layer6_outputs(6161)));
    outputs(3957) <= not(layer6_outputs(5297));
    outputs(3958) <= layer6_outputs(6929);
    outputs(3959) <= (layer6_outputs(3081)) xor (layer6_outputs(6521));
    outputs(3960) <= (layer6_outputs(6957)) xor (layer6_outputs(5384));
    outputs(3961) <= (layer6_outputs(6516)) xor (layer6_outputs(3076));
    outputs(3962) <= not((layer6_outputs(4517)) xor (layer6_outputs(6641)));
    outputs(3963) <= not((layer6_outputs(6192)) xor (layer6_outputs(4292)));
    outputs(3964) <= (layer6_outputs(4025)) and not (layer6_outputs(1976));
    outputs(3965) <= not(layer6_outputs(2988));
    outputs(3966) <= not(layer6_outputs(115));
    outputs(3967) <= not((layer6_outputs(5554)) xor (layer6_outputs(5667)));
    outputs(3968) <= layer6_outputs(7550);
    outputs(3969) <= layer6_outputs(3756);
    outputs(3970) <= not(layer6_outputs(1833));
    outputs(3971) <= layer6_outputs(3759);
    outputs(3972) <= not((layer6_outputs(908)) xor (layer6_outputs(1651)));
    outputs(3973) <= not(layer6_outputs(6679));
    outputs(3974) <= layer6_outputs(6324);
    outputs(3975) <= not(layer6_outputs(6764)) or (layer6_outputs(5743));
    outputs(3976) <= not(layer6_outputs(1476));
    outputs(3977) <= layer6_outputs(1149);
    outputs(3978) <= not((layer6_outputs(3319)) and (layer6_outputs(496)));
    outputs(3979) <= not((layer6_outputs(2686)) xor (layer6_outputs(472)));
    outputs(3980) <= (layer6_outputs(7055)) xor (layer6_outputs(6937));
    outputs(3981) <= not((layer6_outputs(7514)) xor (layer6_outputs(1042)));
    outputs(3982) <= not((layer6_outputs(6499)) xor (layer6_outputs(7153)));
    outputs(3983) <= not((layer6_outputs(2882)) and (layer6_outputs(5653)));
    outputs(3984) <= layer6_outputs(7372);
    outputs(3985) <= not(layer6_outputs(2645));
    outputs(3986) <= layer6_outputs(7552);
    outputs(3987) <= not((layer6_outputs(3017)) xor (layer6_outputs(641)));
    outputs(3988) <= layer6_outputs(5986);
    outputs(3989) <= layer6_outputs(5777);
    outputs(3990) <= not((layer6_outputs(2680)) xor (layer6_outputs(2778)));
    outputs(3991) <= layer6_outputs(6368);
    outputs(3992) <= not(layer6_outputs(3230));
    outputs(3993) <= layer6_outputs(3680);
    outputs(3994) <= not(layer6_outputs(3894)) or (layer6_outputs(7524));
    outputs(3995) <= not((layer6_outputs(4548)) xor (layer6_outputs(7438)));
    outputs(3996) <= (layer6_outputs(2689)) xor (layer6_outputs(1680));
    outputs(3997) <= not((layer6_outputs(1668)) xor (layer6_outputs(3016)));
    outputs(3998) <= layer6_outputs(4382);
    outputs(3999) <= not(layer6_outputs(4296));
    outputs(4000) <= not(layer6_outputs(4417));
    outputs(4001) <= not(layer6_outputs(4578));
    outputs(4002) <= layer6_outputs(4992);
    outputs(4003) <= not(layer6_outputs(3218));
    outputs(4004) <= layer6_outputs(4418);
    outputs(4005) <= layer6_outputs(6545);
    outputs(4006) <= not((layer6_outputs(164)) xor (layer6_outputs(2226)));
    outputs(4007) <= (layer6_outputs(1441)) xor (layer6_outputs(5590));
    outputs(4008) <= (layer6_outputs(2871)) xor (layer6_outputs(571));
    outputs(4009) <= not(layer6_outputs(2382));
    outputs(4010) <= not((layer6_outputs(498)) xor (layer6_outputs(5801)));
    outputs(4011) <= not((layer6_outputs(6385)) xor (layer6_outputs(4230)));
    outputs(4012) <= not(layer6_outputs(2431));
    outputs(4013) <= (layer6_outputs(4390)) xor (layer6_outputs(2233));
    outputs(4014) <= not(layer6_outputs(6641));
    outputs(4015) <= not((layer6_outputs(4789)) xor (layer6_outputs(5705)));
    outputs(4016) <= (layer6_outputs(365)) or (layer6_outputs(453));
    outputs(4017) <= not((layer6_outputs(3914)) xor (layer6_outputs(1576)));
    outputs(4018) <= layer6_outputs(244);
    outputs(4019) <= (layer6_outputs(636)) and not (layer6_outputs(1453));
    outputs(4020) <= layer6_outputs(876);
    outputs(4021) <= not(layer6_outputs(7072));
    outputs(4022) <= not(layer6_outputs(4520));
    outputs(4023) <= layer6_outputs(3087);
    outputs(4024) <= (layer6_outputs(1283)) xor (layer6_outputs(7120));
    outputs(4025) <= not(layer6_outputs(4532));
    outputs(4026) <= (layer6_outputs(3724)) xor (layer6_outputs(999));
    outputs(4027) <= layer6_outputs(4794);
    outputs(4028) <= layer6_outputs(2971);
    outputs(4029) <= not(layer6_outputs(2686));
    outputs(4030) <= layer6_outputs(5517);
    outputs(4031) <= (layer6_outputs(800)) xor (layer6_outputs(4418));
    outputs(4032) <= (layer6_outputs(2949)) and not (layer6_outputs(6360));
    outputs(4033) <= not((layer6_outputs(239)) xor (layer6_outputs(1934)));
    outputs(4034) <= layer6_outputs(2551);
    outputs(4035) <= not(layer6_outputs(4051));
    outputs(4036) <= not(layer6_outputs(1039));
    outputs(4037) <= (layer6_outputs(5902)) xor (layer6_outputs(5302));
    outputs(4038) <= not(layer6_outputs(3025));
    outputs(4039) <= layer6_outputs(6381);
    outputs(4040) <= (layer6_outputs(5497)) xor (layer6_outputs(2717));
    outputs(4041) <= layer6_outputs(6536);
    outputs(4042) <= not((layer6_outputs(2286)) xor (layer6_outputs(1400)));
    outputs(4043) <= not(layer6_outputs(7512));
    outputs(4044) <= (layer6_outputs(4921)) xor (layer6_outputs(5020));
    outputs(4045) <= layer6_outputs(3428);
    outputs(4046) <= (layer6_outputs(3708)) xor (layer6_outputs(4516));
    outputs(4047) <= not((layer6_outputs(847)) xor (layer6_outputs(1547)));
    outputs(4048) <= not(layer6_outputs(4663));
    outputs(4049) <= layer6_outputs(4285);
    outputs(4050) <= layer6_outputs(7608);
    outputs(4051) <= not((layer6_outputs(3596)) xor (layer6_outputs(6733)));
    outputs(4052) <= layer6_outputs(296);
    outputs(4053) <= not(layer6_outputs(6548));
    outputs(4054) <= not((layer6_outputs(2714)) xor (layer6_outputs(1657)));
    outputs(4055) <= layer6_outputs(3638);
    outputs(4056) <= layer6_outputs(6609);
    outputs(4057) <= not(layer6_outputs(1761));
    outputs(4058) <= layer6_outputs(5318);
    outputs(4059) <= not((layer6_outputs(1297)) xor (layer6_outputs(1308)));
    outputs(4060) <= not((layer6_outputs(2467)) xor (layer6_outputs(3184)));
    outputs(4061) <= not(layer6_outputs(267));
    outputs(4062) <= not((layer6_outputs(3090)) xor (layer6_outputs(688)));
    outputs(4063) <= not((layer6_outputs(1228)) xor (layer6_outputs(5028)));
    outputs(4064) <= layer6_outputs(5978);
    outputs(4065) <= layer6_outputs(5844);
    outputs(4066) <= (layer6_outputs(788)) xor (layer6_outputs(4168));
    outputs(4067) <= layer6_outputs(992);
    outputs(4068) <= not((layer6_outputs(506)) xor (layer6_outputs(181)));
    outputs(4069) <= not(layer6_outputs(1994));
    outputs(4070) <= (layer6_outputs(7252)) xor (layer6_outputs(7417));
    outputs(4071) <= layer6_outputs(1265);
    outputs(4072) <= (layer6_outputs(994)) xor (layer6_outputs(2150));
    outputs(4073) <= not((layer6_outputs(2728)) xor (layer6_outputs(825)));
    outputs(4074) <= not((layer6_outputs(3707)) xor (layer6_outputs(5452)));
    outputs(4075) <= (layer6_outputs(4648)) xor (layer6_outputs(2095));
    outputs(4076) <= layer6_outputs(4031);
    outputs(4077) <= not(layer6_outputs(5936));
    outputs(4078) <= not((layer6_outputs(5432)) xor (layer6_outputs(5472)));
    outputs(4079) <= (layer6_outputs(1370)) xor (layer6_outputs(1910));
    outputs(4080) <= (layer6_outputs(6194)) and not (layer6_outputs(4771));
    outputs(4081) <= (layer6_outputs(6710)) xor (layer6_outputs(3753));
    outputs(4082) <= not((layer6_outputs(670)) xor (layer6_outputs(1964)));
    outputs(4083) <= '1';
    outputs(4084) <= layer6_outputs(2505);
    outputs(4085) <= (layer6_outputs(4109)) xor (layer6_outputs(2709));
    outputs(4086) <= not(layer6_outputs(4439));
    outputs(4087) <= layer6_outputs(1352);
    outputs(4088) <= (layer6_outputs(6316)) xor (layer6_outputs(5587));
    outputs(4089) <= not(layer6_outputs(5915));
    outputs(4090) <= (layer6_outputs(2038)) and not (layer6_outputs(2637));
    outputs(4091) <= not(layer6_outputs(2466)) or (layer6_outputs(1943));
    outputs(4092) <= layer6_outputs(5646);
    outputs(4093) <= layer6_outputs(636);
    outputs(4094) <= not(layer6_outputs(3910));
    outputs(4095) <= not(layer6_outputs(3458)) or (layer6_outputs(2230));
    outputs(4096) <= layer6_outputs(3927);
    outputs(4097) <= not(layer6_outputs(5286));
    outputs(4098) <= not(layer6_outputs(5467));
    outputs(4099) <= (layer6_outputs(6951)) xor (layer6_outputs(4270));
    outputs(4100) <= not((layer6_outputs(7111)) or (layer6_outputs(5943)));
    outputs(4101) <= (layer6_outputs(2509)) xor (layer6_outputs(3687));
    outputs(4102) <= not(layer6_outputs(2060));
    outputs(4103) <= not(layer6_outputs(3549));
    outputs(4104) <= layer6_outputs(5847);
    outputs(4105) <= not(layer6_outputs(3599));
    outputs(4106) <= layer6_outputs(2814);
    outputs(4107) <= not(layer6_outputs(7451));
    outputs(4108) <= layer6_outputs(7192);
    outputs(4109) <= (layer6_outputs(3189)) xor (layer6_outputs(3983));
    outputs(4110) <= not(layer6_outputs(524)) or (layer6_outputs(3190));
    outputs(4111) <= layer6_outputs(6198);
    outputs(4112) <= not((layer6_outputs(2095)) and (layer6_outputs(6153)));
    outputs(4113) <= not(layer6_outputs(4261));
    outputs(4114) <= layer6_outputs(6279);
    outputs(4115) <= (layer6_outputs(5474)) or (layer6_outputs(444));
    outputs(4116) <= layer6_outputs(2282);
    outputs(4117) <= not((layer6_outputs(5335)) and (layer6_outputs(3830)));
    outputs(4118) <= (layer6_outputs(7239)) and not (layer6_outputs(87));
    outputs(4119) <= layer6_outputs(3101);
    outputs(4120) <= not(layer6_outputs(5610));
    outputs(4121) <= (layer6_outputs(2592)) xor (layer6_outputs(2369));
    outputs(4122) <= layer6_outputs(184);
    outputs(4123) <= (layer6_outputs(4224)) xor (layer6_outputs(2006));
    outputs(4124) <= not(layer6_outputs(7486));
    outputs(4125) <= not((layer6_outputs(3009)) xor (layer6_outputs(5961)));
    outputs(4126) <= layer6_outputs(6354);
    outputs(4127) <= layer6_outputs(7302);
    outputs(4128) <= not(layer6_outputs(929));
    outputs(4129) <= not(layer6_outputs(3124));
    outputs(4130) <= layer6_outputs(1146);
    outputs(4131) <= layer6_outputs(739);
    outputs(4132) <= (layer6_outputs(1129)) and not (layer6_outputs(1027));
    outputs(4133) <= layer6_outputs(1970);
    outputs(4134) <= not((layer6_outputs(3655)) xor (layer6_outputs(5125)));
    outputs(4135) <= (layer6_outputs(1794)) xor (layer6_outputs(4156));
    outputs(4136) <= layer6_outputs(1734);
    outputs(4137) <= layer6_outputs(2703);
    outputs(4138) <= not((layer6_outputs(5009)) and (layer6_outputs(4383)));
    outputs(4139) <= layer6_outputs(3445);
    outputs(4140) <= not((layer6_outputs(2500)) xor (layer6_outputs(7515)));
    outputs(4141) <= layer6_outputs(3803);
    outputs(4142) <= (layer6_outputs(3271)) and not (layer6_outputs(6242));
    outputs(4143) <= (layer6_outputs(6081)) xor (layer6_outputs(4105));
    outputs(4144) <= not(layer6_outputs(4260));
    outputs(4145) <= layer6_outputs(162);
    outputs(4146) <= (layer6_outputs(3188)) xor (layer6_outputs(5779));
    outputs(4147) <= not(layer6_outputs(1127));
    outputs(4148) <= (layer6_outputs(2062)) xor (layer6_outputs(4931));
    outputs(4149) <= not(layer6_outputs(6200));
    outputs(4150) <= layer6_outputs(456);
    outputs(4151) <= (layer6_outputs(50)) xor (layer6_outputs(6645));
    outputs(4152) <= layer6_outputs(1402);
    outputs(4153) <= (layer6_outputs(3197)) xor (layer6_outputs(5264));
    outputs(4154) <= (layer6_outputs(1050)) and not (layer6_outputs(4190));
    outputs(4155) <= (layer6_outputs(3509)) and (layer6_outputs(6674));
    outputs(4156) <= not(layer6_outputs(3817)) or (layer6_outputs(3082));
    outputs(4157) <= not(layer6_outputs(6925));
    outputs(4158) <= not(layer6_outputs(3716));
    outputs(4159) <= layer6_outputs(6922);
    outputs(4160) <= layer6_outputs(4445);
    outputs(4161) <= layer6_outputs(261);
    outputs(4162) <= not(layer6_outputs(714));
    outputs(4163) <= layer6_outputs(6052);
    outputs(4164) <= not((layer6_outputs(2522)) xor (layer6_outputs(5641)));
    outputs(4165) <= (layer6_outputs(5642)) or (layer6_outputs(4560));
    outputs(4166) <= not((layer6_outputs(4764)) xor (layer6_outputs(811)));
    outputs(4167) <= (layer6_outputs(2673)) and not (layer6_outputs(749));
    outputs(4168) <= not((layer6_outputs(2269)) xor (layer6_outputs(4269)));
    outputs(4169) <= (layer6_outputs(7437)) xor (layer6_outputs(2376));
    outputs(4170) <= layer6_outputs(7098);
    outputs(4171) <= layer6_outputs(6747);
    outputs(4172) <= layer6_outputs(7433);
    outputs(4173) <= not(layer6_outputs(3852));
    outputs(4174) <= not(layer6_outputs(1835));
    outputs(4175) <= layer6_outputs(1297);
    outputs(4176) <= not(layer6_outputs(345));
    outputs(4177) <= not(layer6_outputs(5296));
    outputs(4178) <= not((layer6_outputs(7535)) or (layer6_outputs(3918)));
    outputs(4179) <= not(layer6_outputs(7662));
    outputs(4180) <= not(layer6_outputs(5202));
    outputs(4181) <= layer6_outputs(4344);
    outputs(4182) <= not(layer6_outputs(3852));
    outputs(4183) <= not(layer6_outputs(1511));
    outputs(4184) <= not((layer6_outputs(1162)) xor (layer6_outputs(5725)));
    outputs(4185) <= (layer6_outputs(6954)) xor (layer6_outputs(3111));
    outputs(4186) <= not((layer6_outputs(1868)) xor (layer6_outputs(4885)));
    outputs(4187) <= not((layer6_outputs(3689)) xor (layer6_outputs(5327)));
    outputs(4188) <= not((layer6_outputs(5900)) and (layer6_outputs(3146)));
    outputs(4189) <= not((layer6_outputs(6913)) or (layer6_outputs(6828)));
    outputs(4190) <= (layer6_outputs(6008)) xor (layer6_outputs(3955));
    outputs(4191) <= layer6_outputs(5205);
    outputs(4192) <= not((layer6_outputs(1065)) xor (layer6_outputs(5695)));
    outputs(4193) <= not((layer6_outputs(287)) and (layer6_outputs(4287)));
    outputs(4194) <= (layer6_outputs(4413)) xor (layer6_outputs(623));
    outputs(4195) <= (layer6_outputs(2830)) or (layer6_outputs(6016));
    outputs(4196) <= (layer6_outputs(3340)) xor (layer6_outputs(6685));
    outputs(4197) <= not((layer6_outputs(5398)) xor (layer6_outputs(323)));
    outputs(4198) <= (layer6_outputs(5008)) and not (layer6_outputs(7586));
    outputs(4199) <= layer6_outputs(2669);
    outputs(4200) <= layer6_outputs(6430);
    outputs(4201) <= not(layer6_outputs(6824));
    outputs(4202) <= not(layer6_outputs(6404));
    outputs(4203) <= (layer6_outputs(6996)) xor (layer6_outputs(5161));
    outputs(4204) <= layer6_outputs(6306);
    outputs(4205) <= not((layer6_outputs(4715)) xor (layer6_outputs(6570)));
    outputs(4206) <= not((layer6_outputs(5975)) xor (layer6_outputs(3557)));
    outputs(4207) <= not(layer6_outputs(7303));
    outputs(4208) <= not(layer6_outputs(5759));
    outputs(4209) <= layer6_outputs(1470);
    outputs(4210) <= (layer6_outputs(635)) xor (layer6_outputs(2343));
    outputs(4211) <= not(layer6_outputs(6910));
    outputs(4212) <= not(layer6_outputs(6090));
    outputs(4213) <= not(layer6_outputs(3801));
    outputs(4214) <= not(layer6_outputs(4381)) or (layer6_outputs(7640));
    outputs(4215) <= layer6_outputs(1223);
    outputs(4216) <= layer6_outputs(4877);
    outputs(4217) <= not(layer6_outputs(97));
    outputs(4218) <= (layer6_outputs(7578)) and not (layer6_outputs(2716));
    outputs(4219) <= layer6_outputs(5380);
    outputs(4220) <= not((layer6_outputs(6862)) xor (layer6_outputs(1718)));
    outputs(4221) <= not(layer6_outputs(6462));
    outputs(4222) <= layer6_outputs(5837);
    outputs(4223) <= not(layer6_outputs(6050));
    outputs(4224) <= not((layer6_outputs(3894)) xor (layer6_outputs(479)));
    outputs(4225) <= (layer6_outputs(3355)) xor (layer6_outputs(7155));
    outputs(4226) <= not(layer6_outputs(6301));
    outputs(4227) <= (layer6_outputs(1544)) or (layer6_outputs(1358));
    outputs(4228) <= not(layer6_outputs(1774));
    outputs(4229) <= (layer6_outputs(6006)) or (layer6_outputs(1905));
    outputs(4230) <= layer6_outputs(6921);
    outputs(4231) <= not((layer6_outputs(2757)) xor (layer6_outputs(3670)));
    outputs(4232) <= not((layer6_outputs(1442)) xor (layer6_outputs(1625)));
    outputs(4233) <= not(layer6_outputs(4519));
    outputs(4234) <= not(layer6_outputs(6742));
    outputs(4235) <= (layer6_outputs(3998)) xor (layer6_outputs(1037));
    outputs(4236) <= layer6_outputs(2822);
    outputs(4237) <= not(layer6_outputs(6764));
    outputs(4238) <= layer6_outputs(6787);
    outputs(4239) <= layer6_outputs(5860);
    outputs(4240) <= (layer6_outputs(4946)) xor (layer6_outputs(1986));
    outputs(4241) <= not((layer6_outputs(5449)) xor (layer6_outputs(1654)));
    outputs(4242) <= layer6_outputs(1431);
    outputs(4243) <= not((layer6_outputs(6075)) xor (layer6_outputs(500)));
    outputs(4244) <= not((layer6_outputs(304)) xor (layer6_outputs(934)));
    outputs(4245) <= layer6_outputs(3262);
    outputs(4246) <= not(layer6_outputs(4839));
    outputs(4247) <= (layer6_outputs(3901)) xor (layer6_outputs(7614));
    outputs(4248) <= (layer6_outputs(5292)) and (layer6_outputs(2748));
    outputs(4249) <= layer6_outputs(5141);
    outputs(4250) <= layer6_outputs(6353);
    outputs(4251) <= not(layer6_outputs(1169));
    outputs(4252) <= (layer6_outputs(5505)) xor (layer6_outputs(5290));
    outputs(4253) <= not(layer6_outputs(134));
    outputs(4254) <= (layer6_outputs(4851)) xor (layer6_outputs(3308));
    outputs(4255) <= not((layer6_outputs(3068)) xor (layer6_outputs(5911)));
    outputs(4256) <= not(layer6_outputs(594));
    outputs(4257) <= (layer6_outputs(1471)) xor (layer6_outputs(1496));
    outputs(4258) <= not(layer6_outputs(754));
    outputs(4259) <= not(layer6_outputs(5482));
    outputs(4260) <= not((layer6_outputs(4210)) xor (layer6_outputs(3906)));
    outputs(4261) <= not(layer6_outputs(1192));
    outputs(4262) <= (layer6_outputs(13)) and (layer6_outputs(3669));
    outputs(4263) <= not(layer6_outputs(2069));
    outputs(4264) <= layer6_outputs(6098);
    outputs(4265) <= layer6_outputs(4855);
    outputs(4266) <= layer6_outputs(5016);
    outputs(4267) <= layer6_outputs(5248);
    outputs(4268) <= not(layer6_outputs(4786));
    outputs(4269) <= layer6_outputs(1795);
    outputs(4270) <= layer6_outputs(1776);
    outputs(4271) <= not((layer6_outputs(1514)) or (layer6_outputs(3313)));
    outputs(4272) <= not(layer6_outputs(4057));
    outputs(4273) <= not(layer6_outputs(840));
    outputs(4274) <= not(layer6_outputs(4702));
    outputs(4275) <= not(layer6_outputs(6532));
    outputs(4276) <= layer6_outputs(4848);
    outputs(4277) <= not(layer6_outputs(6210));
    outputs(4278) <= layer6_outputs(5664);
    outputs(4279) <= not(layer6_outputs(2479));
    outputs(4280) <= layer6_outputs(5125);
    outputs(4281) <= (layer6_outputs(7468)) xor (layer6_outputs(6170));
    outputs(4282) <= layer6_outputs(5099);
    outputs(4283) <= layer6_outputs(5658);
    outputs(4284) <= layer6_outputs(119);
    outputs(4285) <= layer6_outputs(7216);
    outputs(4286) <= layer6_outputs(5728);
    outputs(4287) <= not(layer6_outputs(306));
    outputs(4288) <= not(layer6_outputs(5530)) or (layer6_outputs(4020));
    outputs(4289) <= layer6_outputs(2288);
    outputs(4290) <= layer6_outputs(3269);
    outputs(4291) <= not(layer6_outputs(7020));
    outputs(4292) <= not((layer6_outputs(875)) or (layer6_outputs(495)));
    outputs(4293) <= not((layer6_outputs(3688)) xor (layer6_outputs(6017)));
    outputs(4294) <= not(layer6_outputs(5599));
    outputs(4295) <= not(layer6_outputs(5059));
    outputs(4296) <= not((layer6_outputs(984)) and (layer6_outputs(1107)));
    outputs(4297) <= not(layer6_outputs(7498));
    outputs(4298) <= layer6_outputs(1581);
    outputs(4299) <= (layer6_outputs(3141)) xor (layer6_outputs(4649));
    outputs(4300) <= not(layer6_outputs(1032));
    outputs(4301) <= not(layer6_outputs(907));
    outputs(4302) <= (layer6_outputs(2279)) xor (layer6_outputs(2626));
    outputs(4303) <= layer6_outputs(5926);
    outputs(4304) <= (layer6_outputs(3000)) and not (layer6_outputs(5178));
    outputs(4305) <= layer6_outputs(7332);
    outputs(4306) <= not(layer6_outputs(2117));
    outputs(4307) <= (layer6_outputs(5772)) xor (layer6_outputs(7150));
    outputs(4308) <= not(layer6_outputs(2795));
    outputs(4309) <= not(layer6_outputs(5670)) or (layer6_outputs(6440));
    outputs(4310) <= (layer6_outputs(5164)) xor (layer6_outputs(6036));
    outputs(4311) <= layer6_outputs(4279);
    outputs(4312) <= layer6_outputs(1210);
    outputs(4313) <= not((layer6_outputs(4648)) xor (layer6_outputs(7285)));
    outputs(4314) <= (layer6_outputs(3678)) and (layer6_outputs(5555));
    outputs(4315) <= (layer6_outputs(7289)) xor (layer6_outputs(3900));
    outputs(4316) <= not((layer6_outputs(1090)) and (layer6_outputs(2082)));
    outputs(4317) <= layer6_outputs(1621);
    outputs(4318) <= layer6_outputs(2824);
    outputs(4319) <= not(layer6_outputs(6585));
    outputs(4320) <= layer6_outputs(2514);
    outputs(4321) <= layer6_outputs(1751);
    outputs(4322) <= not(layer6_outputs(523));
    outputs(4323) <= (layer6_outputs(2722)) xor (layer6_outputs(5160));
    outputs(4324) <= layer6_outputs(2247);
    outputs(4325) <= not(layer6_outputs(5355));
    outputs(4326) <= not(layer6_outputs(8));
    outputs(4327) <= (layer6_outputs(7162)) or (layer6_outputs(4900));
    outputs(4328) <= not(layer6_outputs(3901));
    outputs(4329) <= layer6_outputs(7082);
    outputs(4330) <= (layer6_outputs(301)) and (layer6_outputs(6852));
    outputs(4331) <= layer6_outputs(5453);
    outputs(4332) <= layer6_outputs(1394);
    outputs(4333) <= (layer6_outputs(2265)) and not (layer6_outputs(4970));
    outputs(4334) <= not(layer6_outputs(5852)) or (layer6_outputs(6063));
    outputs(4335) <= (layer6_outputs(63)) xor (layer6_outputs(440));
    outputs(4336) <= not(layer6_outputs(2449));
    outputs(4337) <= not((layer6_outputs(5064)) xor (layer6_outputs(4860)));
    outputs(4338) <= (layer6_outputs(3422)) and not (layer6_outputs(85));
    outputs(4339) <= layer6_outputs(222);
    outputs(4340) <= layer6_outputs(431);
    outputs(4341) <= layer6_outputs(6278);
    outputs(4342) <= not(layer6_outputs(586)) or (layer6_outputs(7545));
    outputs(4343) <= not((layer6_outputs(5875)) xor (layer6_outputs(2657)));
    outputs(4344) <= not(layer6_outputs(2764));
    outputs(4345) <= layer6_outputs(5584);
    outputs(4346) <= not((layer6_outputs(4064)) and (layer6_outputs(7161)));
    outputs(4347) <= not(layer6_outputs(2281));
    outputs(4348) <= not(layer6_outputs(5915));
    outputs(4349) <= not(layer6_outputs(1782)) or (layer6_outputs(590));
    outputs(4350) <= (layer6_outputs(7513)) xor (layer6_outputs(4782));
    outputs(4351) <= layer6_outputs(7366);
    outputs(4352) <= (layer6_outputs(4880)) or (layer6_outputs(4043));
    outputs(4353) <= layer6_outputs(813);
    outputs(4354) <= (layer6_outputs(5869)) and not (layer6_outputs(606));
    outputs(4355) <= not((layer6_outputs(1681)) xor (layer6_outputs(140)));
    outputs(4356) <= not(layer6_outputs(275));
    outputs(4357) <= not((layer6_outputs(47)) xor (layer6_outputs(82)));
    outputs(4358) <= not(layer6_outputs(4327));
    outputs(4359) <= not(layer6_outputs(5089));
    outputs(4360) <= not(layer6_outputs(578)) or (layer6_outputs(3761));
    outputs(4361) <= layer6_outputs(4285);
    outputs(4362) <= (layer6_outputs(5486)) and not (layer6_outputs(2827));
    outputs(4363) <= layer6_outputs(6061);
    outputs(4364) <= layer6_outputs(4554);
    outputs(4365) <= not(layer6_outputs(3192));
    outputs(4366) <= not((layer6_outputs(6896)) xor (layer6_outputs(7006)));
    outputs(4367) <= (layer6_outputs(2793)) xor (layer6_outputs(5061));
    outputs(4368) <= layer6_outputs(2149);
    outputs(4369) <= not((layer6_outputs(1978)) xor (layer6_outputs(4740)));
    outputs(4370) <= not(layer6_outputs(1603));
    outputs(4371) <= (layer6_outputs(7664)) and (layer6_outputs(7319));
    outputs(4372) <= not(layer6_outputs(3252));
    outputs(4373) <= not((layer6_outputs(6187)) xor (layer6_outputs(1206)));
    outputs(4374) <= layer6_outputs(7528);
    outputs(4375) <= not((layer6_outputs(1413)) or (layer6_outputs(6463)));
    outputs(4376) <= not((layer6_outputs(2036)) and (layer6_outputs(395)));
    outputs(4377) <= not(layer6_outputs(3700));
    outputs(4378) <= not(layer6_outputs(2366));
    outputs(4379) <= not((layer6_outputs(5025)) or (layer6_outputs(2847)));
    outputs(4380) <= not((layer6_outputs(4151)) xor (layer6_outputs(2488)));
    outputs(4381) <= not(layer6_outputs(4359));
    outputs(4382) <= (layer6_outputs(6336)) xor (layer6_outputs(3239));
    outputs(4383) <= layer6_outputs(4685);
    outputs(4384) <= (layer6_outputs(2946)) xor (layer6_outputs(353));
    outputs(4385) <= not(layer6_outputs(4003));
    outputs(4386) <= layer6_outputs(2196);
    outputs(4387) <= layer6_outputs(4180);
    outputs(4388) <= layer6_outputs(5340);
    outputs(4389) <= layer6_outputs(6389);
    outputs(4390) <= layer6_outputs(5787);
    outputs(4391) <= not(layer6_outputs(5789));
    outputs(4392) <= layer6_outputs(2816);
    outputs(4393) <= (layer6_outputs(4551)) xor (layer6_outputs(4108));
    outputs(4394) <= not((layer6_outputs(1900)) and (layer6_outputs(294)));
    outputs(4395) <= (layer6_outputs(7622)) xor (layer6_outputs(6937));
    outputs(4396) <= layer6_outputs(587);
    outputs(4397) <= not(layer6_outputs(3584));
    outputs(4398) <= not(layer6_outputs(3936));
    outputs(4399) <= layer6_outputs(1006);
    outputs(4400) <= not(layer6_outputs(5630));
    outputs(4401) <= layer6_outputs(5008);
    outputs(4402) <= (layer6_outputs(1513)) xor (layer6_outputs(6974));
    outputs(4403) <= (layer6_outputs(660)) xor (layer6_outputs(4502));
    outputs(4404) <= not(layer6_outputs(7186));
    outputs(4405) <= (layer6_outputs(892)) xor (layer6_outputs(5659));
    outputs(4406) <= not(layer6_outputs(4015));
    outputs(4407) <= not(layer6_outputs(3624));
    outputs(4408) <= (layer6_outputs(1587)) xor (layer6_outputs(3990));
    outputs(4409) <= layer6_outputs(2797);
    outputs(4410) <= (layer6_outputs(3204)) xor (layer6_outputs(7474));
    outputs(4411) <= not(layer6_outputs(3809));
    outputs(4412) <= layer6_outputs(5070);
    outputs(4413) <= layer6_outputs(2816);
    outputs(4414) <= not((layer6_outputs(1820)) or (layer6_outputs(3241)));
    outputs(4415) <= not(layer6_outputs(6849));
    outputs(4416) <= not(layer6_outputs(4286));
    outputs(4417) <= not((layer6_outputs(5021)) xor (layer6_outputs(783)));
    outputs(4418) <= (layer6_outputs(5768)) xor (layer6_outputs(4494));
    outputs(4419) <= (layer6_outputs(5758)) xor (layer6_outputs(1553));
    outputs(4420) <= not((layer6_outputs(7247)) xor (layer6_outputs(4021)));
    outputs(4421) <= not((layer6_outputs(6387)) xor (layer6_outputs(4291)));
    outputs(4422) <= not((layer6_outputs(785)) or (layer6_outputs(3325)));
    outputs(4423) <= layer6_outputs(2630);
    outputs(4424) <= (layer6_outputs(3441)) or (layer6_outputs(882));
    outputs(4425) <= layer6_outputs(986);
    outputs(4426) <= not(layer6_outputs(5320));
    outputs(4427) <= (layer6_outputs(1542)) xor (layer6_outputs(3917));
    outputs(4428) <= not(layer6_outputs(4231));
    outputs(4429) <= not(layer6_outputs(2048));
    outputs(4430) <= not((layer6_outputs(1299)) and (layer6_outputs(7069)));
    outputs(4431) <= not((layer6_outputs(203)) and (layer6_outputs(3669)));
    outputs(4432) <= (layer6_outputs(5832)) xor (layer6_outputs(2586));
    outputs(4433) <= (layer6_outputs(5826)) xor (layer6_outputs(2980));
    outputs(4434) <= not(layer6_outputs(4564));
    outputs(4435) <= not((layer6_outputs(3629)) xor (layer6_outputs(5016)));
    outputs(4436) <= not(layer6_outputs(7660)) or (layer6_outputs(711));
    outputs(4437) <= (layer6_outputs(5778)) xor (layer6_outputs(2534));
    outputs(4438) <= not(layer6_outputs(2494));
    outputs(4439) <= (layer6_outputs(814)) and not (layer6_outputs(359));
    outputs(4440) <= not((layer6_outputs(7167)) xor (layer6_outputs(6783)));
    outputs(4441) <= not(layer6_outputs(2067));
    outputs(4442) <= (layer6_outputs(871)) xor (layer6_outputs(2076));
    outputs(4443) <= (layer6_outputs(1187)) and not (layer6_outputs(1862));
    outputs(4444) <= not(layer6_outputs(7652));
    outputs(4445) <= layer6_outputs(7458);
    outputs(4446) <= not(layer6_outputs(6697));
    outputs(4447) <= layer6_outputs(6561);
    outputs(4448) <= not(layer6_outputs(6242));
    outputs(4449) <= (layer6_outputs(1058)) xor (layer6_outputs(5220));
    outputs(4450) <= not(layer6_outputs(2320));
    outputs(4451) <= layer6_outputs(6919);
    outputs(4452) <= not(layer6_outputs(5816)) or (layer6_outputs(1348));
    outputs(4453) <= not(layer6_outputs(56));
    outputs(4454) <= (layer6_outputs(2154)) xor (layer6_outputs(3065));
    outputs(4455) <= layer6_outputs(6238);
    outputs(4456) <= not(layer6_outputs(1156));
    outputs(4457) <= not(layer6_outputs(2370)) or (layer6_outputs(530));
    outputs(4458) <= not((layer6_outputs(4088)) xor (layer6_outputs(4009)));
    outputs(4459) <= (layer6_outputs(544)) and not (layer6_outputs(7273));
    outputs(4460) <= layer6_outputs(3347);
    outputs(4461) <= not((layer6_outputs(4020)) xor (layer6_outputs(12)));
    outputs(4462) <= layer6_outputs(1227);
    outputs(4463) <= not(layer6_outputs(5053));
    outputs(4464) <= layer6_outputs(1028);
    outputs(4465) <= (layer6_outputs(560)) xor (layer6_outputs(926));
    outputs(4466) <= layer6_outputs(904);
    outputs(4467) <= not((layer6_outputs(2573)) xor (layer6_outputs(2406)));
    outputs(4468) <= layer6_outputs(434);
    outputs(4469) <= not((layer6_outputs(5969)) xor (layer6_outputs(961)));
    outputs(4470) <= (layer6_outputs(1201)) and (layer6_outputs(4037));
    outputs(4471) <= not(layer6_outputs(2255));
    outputs(4472) <= not(layer6_outputs(6952));
    outputs(4473) <= not(layer6_outputs(4280));
    outputs(4474) <= layer6_outputs(6596);
    outputs(4475) <= not(layer6_outputs(7367)) or (layer6_outputs(1638));
    outputs(4476) <= not(layer6_outputs(7488));
    outputs(4477) <= not(layer6_outputs(7067));
    outputs(4478) <= not(layer6_outputs(2747));
    outputs(4479) <= not(layer6_outputs(1607)) or (layer6_outputs(7008));
    outputs(4480) <= (layer6_outputs(1623)) xor (layer6_outputs(760));
    outputs(4481) <= layer6_outputs(3978);
    outputs(4482) <= not(layer6_outputs(7611));
    outputs(4483) <= layer6_outputs(7253);
    outputs(4484) <= not(layer6_outputs(3284));
    outputs(4485) <= (layer6_outputs(5567)) and (layer6_outputs(317));
    outputs(4486) <= (layer6_outputs(2990)) xor (layer6_outputs(3488));
    outputs(4487) <= not(layer6_outputs(1698));
    outputs(4488) <= layer6_outputs(6311);
    outputs(4489) <= not(layer6_outputs(3871));
    outputs(4490) <= not(layer6_outputs(4527));
    outputs(4491) <= (layer6_outputs(6156)) xor (layer6_outputs(747));
    outputs(4492) <= (layer6_outputs(2567)) xor (layer6_outputs(2143));
    outputs(4493) <= not((layer6_outputs(4901)) xor (layer6_outputs(6608)));
    outputs(4494) <= layer6_outputs(869);
    outputs(4495) <= not(layer6_outputs(3560));
    outputs(4496) <= not(layer6_outputs(274));
    outputs(4497) <= (layer6_outputs(6831)) xor (layer6_outputs(1829));
    outputs(4498) <= layer6_outputs(3027);
    outputs(4499) <= layer6_outputs(4372);
    outputs(4500) <= not(layer6_outputs(5114)) or (layer6_outputs(3698));
    outputs(4501) <= layer6_outputs(2819);
    outputs(4502) <= (layer6_outputs(3273)) and not (layer6_outputs(5218));
    outputs(4503) <= not(layer6_outputs(7143));
    outputs(4504) <= not((layer6_outputs(4819)) or (layer6_outputs(4245)));
    outputs(4505) <= not(layer6_outputs(445));
    outputs(4506) <= not(layer6_outputs(4954));
    outputs(4507) <= not(layer6_outputs(6947));
    outputs(4508) <= not((layer6_outputs(6519)) xor (layer6_outputs(7030)));
    outputs(4509) <= layer6_outputs(3520);
    outputs(4510) <= not((layer6_outputs(961)) xor (layer6_outputs(4481)));
    outputs(4511) <= layer6_outputs(618);
    outputs(4512) <= layer6_outputs(3095);
    outputs(4513) <= layer6_outputs(1732);
    outputs(4514) <= not(layer6_outputs(2047));
    outputs(4515) <= (layer6_outputs(1115)) xor (layer6_outputs(6213));
    outputs(4516) <= (layer6_outputs(3522)) and not (layer6_outputs(5124));
    outputs(4517) <= layer6_outputs(613);
    outputs(4518) <= not((layer6_outputs(5245)) xor (layer6_outputs(3827)));
    outputs(4519) <= (layer6_outputs(2727)) and not (layer6_outputs(6429));
    outputs(4520) <= (layer6_outputs(6154)) xor (layer6_outputs(6863));
    outputs(4521) <= not(layer6_outputs(2642));
    outputs(4522) <= not(layer6_outputs(219)) or (layer6_outputs(2634));
    outputs(4523) <= not(layer6_outputs(4245));
    outputs(4524) <= layer6_outputs(1588);
    outputs(4525) <= not((layer6_outputs(6560)) xor (layer6_outputs(5943)));
    outputs(4526) <= not(layer6_outputs(5853));
    outputs(4527) <= not((layer6_outputs(6813)) xor (layer6_outputs(6275)));
    outputs(4528) <= not(layer6_outputs(20));
    outputs(4529) <= (layer6_outputs(4123)) xor (layer6_outputs(6309));
    outputs(4530) <= layer6_outputs(5471);
    outputs(4531) <= layer6_outputs(1153);
    outputs(4532) <= (layer6_outputs(3754)) xor (layer6_outputs(927));
    outputs(4533) <= layer6_outputs(2913);
    outputs(4534) <= layer6_outputs(2909);
    outputs(4535) <= not(layer6_outputs(1502));
    outputs(4536) <= not(layer6_outputs(1915)) or (layer6_outputs(3774));
    outputs(4537) <= layer6_outputs(1118);
    outputs(4538) <= layer6_outputs(1375);
    outputs(4539) <= layer6_outputs(6682);
    outputs(4540) <= layer6_outputs(7026);
    outputs(4541) <= (layer6_outputs(4044)) xor (layer6_outputs(5982));
    outputs(4542) <= layer6_outputs(5403);
    outputs(4543) <= not(layer6_outputs(5089));
    outputs(4544) <= not(layer6_outputs(305));
    outputs(4545) <= not(layer6_outputs(4303));
    outputs(4546) <= layer6_outputs(6868);
    outputs(4547) <= layer6_outputs(5950);
    outputs(4548) <= not(layer6_outputs(455));
    outputs(4549) <= not(layer6_outputs(1453));
    outputs(4550) <= layer6_outputs(5658);
    outputs(4551) <= (layer6_outputs(7254)) xor (layer6_outputs(5866));
    outputs(4552) <= (layer6_outputs(5041)) xor (layer6_outputs(1899));
    outputs(4553) <= not(layer6_outputs(7108)) or (layer6_outputs(3486));
    outputs(4554) <= not((layer6_outputs(3332)) xor (layer6_outputs(1212)));
    outputs(4555) <= not((layer6_outputs(5367)) xor (layer6_outputs(2490)));
    outputs(4556) <= (layer6_outputs(6150)) and not (layer6_outputs(7205));
    outputs(4557) <= layer6_outputs(487);
    outputs(4558) <= not(layer6_outputs(7396));
    outputs(4559) <= not(layer6_outputs(899));
    outputs(4560) <= layer6_outputs(4233);
    outputs(4561) <= not((layer6_outputs(4184)) xor (layer6_outputs(1923)));
    outputs(4562) <= not((layer6_outputs(7311)) xor (layer6_outputs(822)));
    outputs(4563) <= layer6_outputs(4058);
    outputs(4564) <= not(layer6_outputs(3651));
    outputs(4565) <= layer6_outputs(6331);
    outputs(4566) <= not((layer6_outputs(3314)) xor (layer6_outputs(4197)));
    outputs(4567) <= not(layer6_outputs(6433));
    outputs(4568) <= layer6_outputs(2410);
    outputs(4569) <= layer6_outputs(3519);
    outputs(4570) <= (layer6_outputs(7590)) xor (layer6_outputs(1475));
    outputs(4571) <= (layer6_outputs(1081)) xor (layer6_outputs(3949));
    outputs(4572) <= not(layer6_outputs(3510));
    outputs(4573) <= (layer6_outputs(4141)) or (layer6_outputs(6414));
    outputs(4574) <= not((layer6_outputs(4990)) xor (layer6_outputs(1687)));
    outputs(4575) <= (layer6_outputs(3733)) xor (layer6_outputs(2692));
    outputs(4576) <= not(layer6_outputs(1484));
    outputs(4577) <= (layer6_outputs(7239)) or (layer6_outputs(6083));
    outputs(4578) <= not(layer6_outputs(988));
    outputs(4579) <= not((layer6_outputs(1634)) xor (layer6_outputs(4709)));
    outputs(4580) <= not((layer6_outputs(818)) xor (layer6_outputs(4257)));
    outputs(4581) <= not(layer6_outputs(1096));
    outputs(4582) <= (layer6_outputs(53)) xor (layer6_outputs(7532));
    outputs(4583) <= (layer6_outputs(6635)) xor (layer6_outputs(439));
    outputs(4584) <= not(layer6_outputs(2358));
    outputs(4585) <= not(layer6_outputs(4928));
    outputs(4586) <= layer6_outputs(6505);
    outputs(4587) <= (layer6_outputs(1345)) and not (layer6_outputs(2213));
    outputs(4588) <= (layer6_outputs(6424)) and (layer6_outputs(3029));
    outputs(4589) <= layer6_outputs(7349);
    outputs(4590) <= not(layer6_outputs(3517));
    outputs(4591) <= (layer6_outputs(4918)) and (layer6_outputs(1088));
    outputs(4592) <= not((layer6_outputs(2445)) xor (layer6_outputs(2773)));
    outputs(4593) <= not(layer6_outputs(3627));
    outputs(4594) <= layer6_outputs(3881);
    outputs(4595) <= not(layer6_outputs(2736));
    outputs(4596) <= layer6_outputs(5);
    outputs(4597) <= layer6_outputs(697);
    outputs(4598) <= not((layer6_outputs(4658)) xor (layer6_outputs(2529)));
    outputs(4599) <= not(layer6_outputs(5143));
    outputs(4600) <= layer6_outputs(6998);
    outputs(4601) <= layer6_outputs(2386);
    outputs(4602) <= (layer6_outputs(619)) xor (layer6_outputs(6769));
    outputs(4603) <= (layer6_outputs(2560)) and not (layer6_outputs(5857));
    outputs(4604) <= not((layer6_outputs(305)) xor (layer6_outputs(5801)));
    outputs(4605) <= layer6_outputs(2132);
    outputs(4606) <= not(layer6_outputs(1843));
    outputs(4607) <= not(layer6_outputs(3287));
    outputs(4608) <= not((layer6_outputs(3212)) and (layer6_outputs(278)));
    outputs(4609) <= not(layer6_outputs(6601));
    outputs(4610) <= (layer6_outputs(4579)) xor (layer6_outputs(3675));
    outputs(4611) <= not(layer6_outputs(175));
    outputs(4612) <= (layer6_outputs(1648)) and not (layer6_outputs(1847));
    outputs(4613) <= layer6_outputs(7548);
    outputs(4614) <= not(layer6_outputs(1194));
    outputs(4615) <= not(layer6_outputs(6702));
    outputs(4616) <= layer6_outputs(973);
    outputs(4617) <= not(layer6_outputs(5464));
    outputs(4618) <= not(layer6_outputs(6166));
    outputs(4619) <= (layer6_outputs(1391)) xor (layer6_outputs(7055));
    outputs(4620) <= not(layer6_outputs(2943));
    outputs(4621) <= (layer6_outputs(2055)) xor (layer6_outputs(2635));
    outputs(4622) <= (layer6_outputs(7326)) xor (layer6_outputs(4651));
    outputs(4623) <= not(layer6_outputs(1731));
    outputs(4624) <= not((layer6_outputs(772)) or (layer6_outputs(404)));
    outputs(4625) <= layer6_outputs(4367);
    outputs(4626) <= layer6_outputs(4945);
    outputs(4627) <= layer6_outputs(6753);
    outputs(4628) <= (layer6_outputs(5792)) or (layer6_outputs(5783));
    outputs(4629) <= (layer6_outputs(7130)) and (layer6_outputs(1535));
    outputs(4630) <= layer6_outputs(72);
    outputs(4631) <= not((layer6_outputs(2037)) and (layer6_outputs(1134)));
    outputs(4632) <= not(layer6_outputs(2739));
    outputs(4633) <= not(layer6_outputs(2595));
    outputs(4634) <= layer6_outputs(0);
    outputs(4635) <= not(layer6_outputs(3209));
    outputs(4636) <= (layer6_outputs(1427)) xor (layer6_outputs(3921));
    outputs(4637) <= layer6_outputs(4117);
    outputs(4638) <= not(layer6_outputs(2072));
    outputs(4639) <= not(layer6_outputs(2694));
    outputs(4640) <= (layer6_outputs(1376)) and not (layer6_outputs(2719));
    outputs(4641) <= not(layer6_outputs(4851)) or (layer6_outputs(4708));
    outputs(4642) <= layer6_outputs(3312);
    outputs(4643) <= (layer6_outputs(1897)) and (layer6_outputs(4462));
    outputs(4644) <= layer6_outputs(605);
    outputs(4645) <= (layer6_outputs(4767)) xor (layer6_outputs(7587));
    outputs(4646) <= layer6_outputs(3013);
    outputs(4647) <= not(layer6_outputs(1380));
    outputs(4648) <= not(layer6_outputs(2940));
    outputs(4649) <= not(layer6_outputs(5841));
    outputs(4650) <= not((layer6_outputs(5612)) xor (layer6_outputs(2579)));
    outputs(4651) <= not((layer6_outputs(5880)) and (layer6_outputs(7602)));
    outputs(4652) <= not(layer6_outputs(2545));
    outputs(4653) <= (layer6_outputs(1622)) xor (layer6_outputs(2388));
    outputs(4654) <= layer6_outputs(915);
    outputs(4655) <= (layer6_outputs(1631)) and (layer6_outputs(3213));
    outputs(4656) <= not(layer6_outputs(2423));
    outputs(4657) <= (layer6_outputs(2827)) and (layer6_outputs(7216));
    outputs(4658) <= layer6_outputs(640);
    outputs(4659) <= (layer6_outputs(1147)) and not (layer6_outputs(6120));
    outputs(4660) <= (layer6_outputs(4680)) and (layer6_outputs(3701));
    outputs(4661) <= not(layer6_outputs(7246));
    outputs(4662) <= not(layer6_outputs(6234));
    outputs(4663) <= layer6_outputs(5478);
    outputs(4664) <= layer6_outputs(2742);
    outputs(4665) <= layer6_outputs(5591);
    outputs(4666) <= not(layer6_outputs(4473));
    outputs(4667) <= not(layer6_outputs(5693));
    outputs(4668) <= layer6_outputs(2542);
    outputs(4669) <= not(layer6_outputs(4720));
    outputs(4670) <= layer6_outputs(3777);
    outputs(4671) <= (layer6_outputs(6326)) xor (layer6_outputs(5045));
    outputs(4672) <= not(layer6_outputs(999));
    outputs(4673) <= layer6_outputs(1767);
    outputs(4674) <= not(layer6_outputs(5319));
    outputs(4675) <= (layer6_outputs(1775)) or (layer6_outputs(1440));
    outputs(4676) <= layer6_outputs(200);
    outputs(4677) <= layer6_outputs(7605);
    outputs(4678) <= layer6_outputs(24);
    outputs(4679) <= not(layer6_outputs(5914));
    outputs(4680) <= (layer6_outputs(2182)) xor (layer6_outputs(2688));
    outputs(4681) <= (layer6_outputs(7177)) xor (layer6_outputs(4406));
    outputs(4682) <= (layer6_outputs(7294)) and not (layer6_outputs(6312));
    outputs(4683) <= layer6_outputs(2269);
    outputs(4684) <= not(layer6_outputs(4611));
    outputs(4685) <= (layer6_outputs(3083)) xor (layer6_outputs(4104));
    outputs(4686) <= layer6_outputs(1172);
    outputs(4687) <= not(layer6_outputs(1551));
    outputs(4688) <= (layer6_outputs(1643)) xor (layer6_outputs(4638));
    outputs(4689) <= not((layer6_outputs(6403)) xor (layer6_outputs(704)));
    outputs(4690) <= not(layer6_outputs(4647));
    outputs(4691) <= (layer6_outputs(7225)) and not (layer6_outputs(7188));
    outputs(4692) <= not(layer6_outputs(4180));
    outputs(4693) <= not(layer6_outputs(7472));
    outputs(4694) <= layer6_outputs(3423);
    outputs(4695) <= not(layer6_outputs(3517));
    outputs(4696) <= not((layer6_outputs(5128)) xor (layer6_outputs(3387)));
    outputs(4697) <= layer6_outputs(4729);
    outputs(4698) <= not(layer6_outputs(5026));
    outputs(4699) <= layer6_outputs(7307);
    outputs(4700) <= not((layer6_outputs(5311)) xor (layer6_outputs(7492)));
    outputs(4701) <= not(layer6_outputs(5709));
    outputs(4702) <= layer6_outputs(671);
    outputs(4703) <= not((layer6_outputs(809)) xor (layer6_outputs(5637)));
    outputs(4704) <= (layer6_outputs(4569)) and not (layer6_outputs(6553));
    outputs(4705) <= not(layer6_outputs(3577));
    outputs(4706) <= layer6_outputs(5575);
    outputs(4707) <= not(layer6_outputs(3580));
    outputs(4708) <= layer6_outputs(4850);
    outputs(4709) <= not((layer6_outputs(1165)) xor (layer6_outputs(3262)));
    outputs(4710) <= layer6_outputs(887);
    outputs(4711) <= layer6_outputs(3945);
    outputs(4712) <= layer6_outputs(6274);
    outputs(4713) <= not((layer6_outputs(1990)) xor (layer6_outputs(4534)));
    outputs(4714) <= not(layer6_outputs(3602));
    outputs(4715) <= not(layer6_outputs(4978));
    outputs(4716) <= (layer6_outputs(7560)) xor (layer6_outputs(7009));
    outputs(4717) <= not(layer6_outputs(2221));
    outputs(4718) <= layer6_outputs(5798);
    outputs(4719) <= layer6_outputs(3786);
    outputs(4720) <= layer6_outputs(6987);
    outputs(4721) <= not(layer6_outputs(7344));
    outputs(4722) <= (layer6_outputs(2461)) xor (layer6_outputs(2702));
    outputs(4723) <= not(layer6_outputs(2869));
    outputs(4724) <= not(layer6_outputs(4585));
    outputs(4725) <= not(layer6_outputs(1320));
    outputs(4726) <= not((layer6_outputs(6988)) and (layer6_outputs(2724)));
    outputs(4727) <= not((layer6_outputs(2313)) xor (layer6_outputs(1834)));
    outputs(4728) <= not(layer6_outputs(5550));
    outputs(4729) <= not(layer6_outputs(3192));
    outputs(4730) <= layer6_outputs(2047);
    outputs(4731) <= layer6_outputs(1113);
    outputs(4732) <= not((layer6_outputs(6299)) xor (layer6_outputs(1808)));
    outputs(4733) <= not(layer6_outputs(5694));
    outputs(4734) <= layer6_outputs(1962);
    outputs(4735) <= (layer6_outputs(6303)) and not (layer6_outputs(5140));
    outputs(4736) <= (layer6_outputs(3052)) xor (layer6_outputs(4023));
    outputs(4737) <= layer6_outputs(3036);
    outputs(4738) <= not(layer6_outputs(4162));
    outputs(4739) <= layer6_outputs(3784);
    outputs(4740) <= not(layer6_outputs(4984));
    outputs(4741) <= (layer6_outputs(5483)) xor (layer6_outputs(204));
    outputs(4742) <= layer6_outputs(3639);
    outputs(4743) <= not(layer6_outputs(2574));
    outputs(4744) <= not(layer6_outputs(2019));
    outputs(4745) <= not((layer6_outputs(4463)) or (layer6_outputs(4995)));
    outputs(4746) <= not(layer6_outputs(2616));
    outputs(4747) <= layer6_outputs(2379);
    outputs(4748) <= not(layer6_outputs(6259));
    outputs(4749) <= (layer6_outputs(218)) xor (layer6_outputs(3434));
    outputs(4750) <= layer6_outputs(7293);
    outputs(4751) <= (layer6_outputs(6089)) xor (layer6_outputs(4395));
    outputs(4752) <= (layer6_outputs(1360)) xor (layer6_outputs(1380));
    outputs(4753) <= not((layer6_outputs(7215)) xor (layer6_outputs(6494)));
    outputs(4754) <= layer6_outputs(4100);
    outputs(4755) <= layer6_outputs(5063);
    outputs(4756) <= layer6_outputs(4320);
    outputs(4757) <= not(layer6_outputs(4678));
    outputs(4758) <= layer6_outputs(4454);
    outputs(4759) <= layer6_outputs(4169);
    outputs(4760) <= (layer6_outputs(6777)) and (layer6_outputs(2685));
    outputs(4761) <= (layer6_outputs(6178)) and (layer6_outputs(3730));
    outputs(4762) <= not(layer6_outputs(4248));
    outputs(4763) <= not((layer6_outputs(4950)) and (layer6_outputs(20)));
    outputs(4764) <= layer6_outputs(4729);
    outputs(4765) <= layer6_outputs(2651);
    outputs(4766) <= not(layer6_outputs(3908));
    outputs(4767) <= (layer6_outputs(6536)) and not (layer6_outputs(7607));
    outputs(4768) <= not(layer6_outputs(4325));
    outputs(4769) <= not(layer6_outputs(6983));
    outputs(4770) <= layer6_outputs(6589);
    outputs(4771) <= not(layer6_outputs(6835));
    outputs(4772) <= not(layer6_outputs(6789));
    outputs(4773) <= not(layer6_outputs(824));
    outputs(4774) <= (layer6_outputs(3623)) and not (layer6_outputs(1979));
    outputs(4775) <= not(layer6_outputs(7634));
    outputs(4776) <= layer6_outputs(5101);
    outputs(4777) <= (layer6_outputs(4866)) xor (layer6_outputs(4139));
    outputs(4778) <= not(layer6_outputs(7081));
    outputs(4779) <= not(layer6_outputs(603));
    outputs(4780) <= (layer6_outputs(2436)) xor (layer6_outputs(3491));
    outputs(4781) <= not(layer6_outputs(6740));
    outputs(4782) <= not(layer6_outputs(1311));
    outputs(4783) <= layer6_outputs(4442);
    outputs(4784) <= not((layer6_outputs(91)) xor (layer6_outputs(4490)));
    outputs(4785) <= layer6_outputs(5189);
    outputs(4786) <= layer6_outputs(7038);
    outputs(4787) <= layer6_outputs(1814);
    outputs(4788) <= not(layer6_outputs(424));
    outputs(4789) <= not(layer6_outputs(6147)) or (layer6_outputs(5912));
    outputs(4790) <= not(layer6_outputs(5859));
    outputs(4791) <= not((layer6_outputs(7301)) or (layer6_outputs(5310)));
    outputs(4792) <= (layer6_outputs(2020)) xor (layer6_outputs(6333));
    outputs(4793) <= (layer6_outputs(1756)) xor (layer6_outputs(7240));
    outputs(4794) <= layer6_outputs(1689);
    outputs(4795) <= (layer6_outputs(774)) xor (layer6_outputs(1897));
    outputs(4796) <= not(layer6_outputs(6979));
    outputs(4797) <= not((layer6_outputs(2848)) xor (layer6_outputs(6251)));
    outputs(4798) <= layer6_outputs(718);
    outputs(4799) <= not((layer6_outputs(5876)) xor (layer6_outputs(6419)));
    outputs(4800) <= not(layer6_outputs(5433));
    outputs(4801) <= not((layer6_outputs(4475)) xor (layer6_outputs(647)));
    outputs(4802) <= not(layer6_outputs(2371));
    outputs(4803) <= not((layer6_outputs(777)) xor (layer6_outputs(7598)));
    outputs(4804) <= not(layer6_outputs(5634));
    outputs(4805) <= layer6_outputs(2056);
    outputs(4806) <= (layer6_outputs(567)) xor (layer6_outputs(1018));
    outputs(4807) <= (layer6_outputs(124)) and not (layer6_outputs(6415));
    outputs(4808) <= (layer6_outputs(5240)) and not (layer6_outputs(3098));
    outputs(4809) <= not(layer6_outputs(3277));
    outputs(4810) <= not(layer6_outputs(5178));
    outputs(4811) <= layer6_outputs(2926);
    outputs(4812) <= not(layer6_outputs(60));
    outputs(4813) <= not(layer6_outputs(7207)) or (layer6_outputs(3913));
    outputs(4814) <= (layer6_outputs(5520)) and not (layer6_outputs(5207));
    outputs(4815) <= (layer6_outputs(7151)) and not (layer6_outputs(6724));
    outputs(4816) <= not(layer6_outputs(3964));
    outputs(4817) <= not(layer6_outputs(1478));
    outputs(4818) <= not(layer6_outputs(4908)) or (layer6_outputs(6272));
    outputs(4819) <= (layer6_outputs(2632)) and not (layer6_outputs(7542));
    outputs(4820) <= layer6_outputs(5441);
    outputs(4821) <= (layer6_outputs(2517)) and not (layer6_outputs(7335));
    outputs(4822) <= layer6_outputs(2933);
    outputs(4823) <= (layer6_outputs(1886)) xor (layer6_outputs(5195));
    outputs(4824) <= not((layer6_outputs(373)) xor (layer6_outputs(6876)));
    outputs(4825) <= layer6_outputs(1219);
    outputs(4826) <= not((layer6_outputs(7491)) xor (layer6_outputs(1675)));
    outputs(4827) <= layer6_outputs(926);
    outputs(4828) <= (layer6_outputs(6139)) and (layer6_outputs(1157));
    outputs(4829) <= not(layer6_outputs(7529));
    outputs(4830) <= not((layer6_outputs(872)) xor (layer6_outputs(3801)));
    outputs(4831) <= not(layer6_outputs(5139));
    outputs(4832) <= not((layer6_outputs(4099)) or (layer6_outputs(1468)));
    outputs(4833) <= not(layer6_outputs(1909));
    outputs(4834) <= (layer6_outputs(404)) xor (layer6_outputs(3043));
    outputs(4835) <= (layer6_outputs(2799)) xor (layer6_outputs(6833));
    outputs(4836) <= (layer6_outputs(960)) xor (layer6_outputs(1689));
    outputs(4837) <= not((layer6_outputs(1213)) xor (layer6_outputs(5129)));
    outputs(4838) <= not(layer6_outputs(7315));
    outputs(4839) <= layer6_outputs(2353);
    outputs(4840) <= (layer6_outputs(997)) xor (layer6_outputs(212));
    outputs(4841) <= not(layer6_outputs(4884));
    outputs(4842) <= not(layer6_outputs(6215));
    outputs(4843) <= not(layer6_outputs(4263));
    outputs(4844) <= (layer6_outputs(4873)) and not (layer6_outputs(2639));
    outputs(4845) <= (layer6_outputs(2409)) and not (layer6_outputs(2441));
    outputs(4846) <= layer6_outputs(3083);
    outputs(4847) <= not(layer6_outputs(495));
    outputs(4848) <= not((layer6_outputs(675)) xor (layer6_outputs(1590)));
    outputs(4849) <= not(layer6_outputs(6043));
    outputs(4850) <= layer6_outputs(7131);
    outputs(4851) <= (layer6_outputs(3612)) xor (layer6_outputs(2791));
    outputs(4852) <= (layer6_outputs(6399)) and (layer6_outputs(804));
    outputs(4853) <= layer6_outputs(151);
    outputs(4854) <= (layer6_outputs(4482)) xor (layer6_outputs(5043));
    outputs(4855) <= (layer6_outputs(7074)) xor (layer6_outputs(5886));
    outputs(4856) <= layer6_outputs(4872);
    outputs(4857) <= not(layer6_outputs(6632));
    outputs(4858) <= not(layer6_outputs(101));
    outputs(4859) <= layer6_outputs(1172);
    outputs(4860) <= (layer6_outputs(1797)) and not (layer6_outputs(5368));
    outputs(4861) <= not(layer6_outputs(6927));
    outputs(4862) <= layer6_outputs(7530);
    outputs(4863) <= layer6_outputs(4719);
    outputs(4864) <= not((layer6_outputs(2693)) or (layer6_outputs(7218)));
    outputs(4865) <= not(layer6_outputs(946));
    outputs(4866) <= not((layer6_outputs(3583)) xor (layer6_outputs(7676)));
    outputs(4867) <= not(layer6_outputs(3587));
    outputs(4868) <= (layer6_outputs(2434)) and (layer6_outputs(4014));
    outputs(4869) <= layer6_outputs(5812);
    outputs(4870) <= layer6_outputs(4944);
    outputs(4871) <= not(layer6_outputs(4261));
    outputs(4872) <= not(layer6_outputs(5565));
    outputs(4873) <= not(layer6_outputs(5965));
    outputs(4874) <= layer6_outputs(5559);
    outputs(4875) <= not(layer6_outputs(1458));
    outputs(4876) <= not(layer6_outputs(5215));
    outputs(4877) <= not(layer6_outputs(224));
    outputs(4878) <= layer6_outputs(1798);
    outputs(4879) <= (layer6_outputs(5068)) and not (layer6_outputs(1477));
    outputs(4880) <= layer6_outputs(2529);
    outputs(4881) <= layer6_outputs(5034);
    outputs(4882) <= (layer6_outputs(2788)) and not (layer6_outputs(3533));
    outputs(4883) <= (layer6_outputs(1629)) and not (layer6_outputs(2916));
    outputs(4884) <= not(layer6_outputs(5424));
    outputs(4885) <= not(layer6_outputs(7344));
    outputs(4886) <= not((layer6_outputs(7533)) xor (layer6_outputs(5603)));
    outputs(4887) <= layer6_outputs(652);
    outputs(4888) <= (layer6_outputs(1068)) and not (layer6_outputs(1403));
    outputs(4889) <= not(layer6_outputs(5901));
    outputs(4890) <= layer6_outputs(5522);
    outputs(4891) <= layer6_outputs(3155);
    outputs(4892) <= (layer6_outputs(3799)) xor (layer6_outputs(2791));
    outputs(4893) <= not(layer6_outputs(3110));
    outputs(4894) <= layer6_outputs(1995);
    outputs(4895) <= layer6_outputs(1007);
    outputs(4896) <= not(layer6_outputs(4672));
    outputs(4897) <= (layer6_outputs(2931)) and not (layer6_outputs(1011));
    outputs(4898) <= layer6_outputs(1166);
    outputs(4899) <= layer6_outputs(46);
    outputs(4900) <= layer6_outputs(977);
    outputs(4901) <= not(layer6_outputs(4432));
    outputs(4902) <= not((layer6_outputs(7570)) and (layer6_outputs(1654)));
    outputs(4903) <= (layer6_outputs(746)) xor (layer6_outputs(7588));
    outputs(4904) <= not(layer6_outputs(1350));
    outputs(4905) <= (layer6_outputs(4379)) and (layer6_outputs(7517));
    outputs(4906) <= layer6_outputs(5205);
    outputs(4907) <= not(layer6_outputs(4927));
    outputs(4908) <= layer6_outputs(5328);
    outputs(4909) <= (layer6_outputs(4244)) xor (layer6_outputs(734));
    outputs(4910) <= not((layer6_outputs(897)) or (layer6_outputs(4385)));
    outputs(4911) <= not(layer6_outputs(3927));
    outputs(4912) <= not(layer6_outputs(1450));
    outputs(4913) <= not(layer6_outputs(7014));
    outputs(4914) <= layer6_outputs(2917);
    outputs(4915) <= (layer6_outputs(113)) or (layer6_outputs(652));
    outputs(4916) <= not(layer6_outputs(2624));
    outputs(4917) <= not(layer6_outputs(1539));
    outputs(4918) <= not(layer6_outputs(2845));
    outputs(4919) <= layer6_outputs(5067);
    outputs(4920) <= (layer6_outputs(1757)) xor (layer6_outputs(7141));
    outputs(4921) <= layer6_outputs(4891);
    outputs(4922) <= (layer6_outputs(2936)) or (layer6_outputs(293));
    outputs(4923) <= not((layer6_outputs(363)) and (layer6_outputs(4026)));
    outputs(4924) <= not(layer6_outputs(3367));
    outputs(4925) <= not((layer6_outputs(1576)) and (layer6_outputs(4388)));
    outputs(4926) <= not((layer6_outputs(4557)) xor (layer6_outputs(3867)));
    outputs(4927) <= layer6_outputs(6629);
    outputs(4928) <= not(layer6_outputs(127));
    outputs(4929) <= (layer6_outputs(2605)) xor (layer6_outputs(5542));
    outputs(4930) <= layer6_outputs(1324);
    outputs(4931) <= not((layer6_outputs(7598)) and (layer6_outputs(129)));
    outputs(4932) <= (layer6_outputs(6039)) xor (layer6_outputs(2297));
    outputs(4933) <= layer6_outputs(2100);
    outputs(4934) <= not(layer6_outputs(63));
    outputs(4935) <= not((layer6_outputs(6122)) xor (layer6_outputs(2759)));
    outputs(4936) <= not(layer6_outputs(3603));
    outputs(4937) <= layer6_outputs(303);
    outputs(4938) <= (layer6_outputs(4544)) xor (layer6_outputs(6371));
    outputs(4939) <= layer6_outputs(1158);
    outputs(4940) <= not((layer6_outputs(3121)) or (layer6_outputs(4757)));
    outputs(4941) <= (layer6_outputs(1381)) or (layer6_outputs(5792));
    outputs(4942) <= layer6_outputs(7032);
    outputs(4943) <= layer6_outputs(7507);
    outputs(4944) <= layer6_outputs(3205);
    outputs(4945) <= not(layer6_outputs(3819));
    outputs(4946) <= layer6_outputs(2191);
    outputs(4947) <= not(layer6_outputs(2283));
    outputs(4948) <= not(layer6_outputs(5329));
    outputs(4949) <= not((layer6_outputs(1205)) or (layer6_outputs(6730)));
    outputs(4950) <= not(layer6_outputs(4955));
    outputs(4951) <= layer6_outputs(2623);
    outputs(4952) <= not(layer6_outputs(3159)) or (layer6_outputs(7084));
    outputs(4953) <= not(layer6_outputs(1804));
    outputs(4954) <= layer6_outputs(2514);
    outputs(4955) <= layer6_outputs(7610);
    outputs(4956) <= layer6_outputs(4619);
    outputs(4957) <= layer6_outputs(7494);
    outputs(4958) <= not(layer6_outputs(1175));
    outputs(4959) <= layer6_outputs(3665);
    outputs(4960) <= layer6_outputs(7537);
    outputs(4961) <= not((layer6_outputs(779)) and (layer6_outputs(5252)));
    outputs(4962) <= not(layer6_outputs(41));
    outputs(4963) <= not((layer6_outputs(5750)) xor (layer6_outputs(2921)));
    outputs(4964) <= not(layer6_outputs(71));
    outputs(4965) <= (layer6_outputs(5615)) and not (layer6_outputs(3729));
    outputs(4966) <= not((layer6_outputs(3019)) xor (layer6_outputs(2539)));
    outputs(4967) <= not((layer6_outputs(2456)) xor (layer6_outputs(6359)));
    outputs(4968) <= not(layer6_outputs(1121));
    outputs(4969) <= (layer6_outputs(7148)) xor (layer6_outputs(3711));
    outputs(4970) <= layer6_outputs(6491);
    outputs(4971) <= not(layer6_outputs(5149));
    outputs(4972) <= not(layer6_outputs(3727));
    outputs(4973) <= layer6_outputs(7666);
    outputs(4974) <= not(layer6_outputs(5902));
    outputs(4975) <= layer6_outputs(6512);
    outputs(4976) <= not((layer6_outputs(1791)) xor (layer6_outputs(6141)));
    outputs(4977) <= not((layer6_outputs(4530)) xor (layer6_outputs(997)));
    outputs(4978) <= layer6_outputs(6210);
    outputs(4979) <= layer6_outputs(4411);
    outputs(4980) <= layer6_outputs(2687);
    outputs(4981) <= layer6_outputs(2925);
    outputs(4982) <= not(layer6_outputs(3595));
    outputs(4983) <= not(layer6_outputs(1972));
    outputs(4984) <= not(layer6_outputs(6159));
    outputs(4985) <= not(layer6_outputs(3122));
    outputs(4986) <= (layer6_outputs(3742)) xor (layer6_outputs(1481));
    outputs(4987) <= layer6_outputs(7593);
    outputs(4988) <= layer6_outputs(643);
    outputs(4989) <= (layer6_outputs(5487)) xor (layer6_outputs(2853));
    outputs(4990) <= not(layer6_outputs(4957));
    outputs(4991) <= layer6_outputs(5944);
    outputs(4992) <= not(layer6_outputs(1450));
    outputs(4993) <= layer6_outputs(6506);
    outputs(4994) <= (layer6_outputs(968)) xor (layer6_outputs(4066));
    outputs(4995) <= layer6_outputs(6504);
    outputs(4996) <= not(layer6_outputs(7308));
    outputs(4997) <= not(layer6_outputs(2397));
    outputs(4998) <= layer6_outputs(6074);
    outputs(4999) <= (layer6_outputs(5358)) xor (layer6_outputs(4192));
    outputs(5000) <= not((layer6_outputs(2237)) xor (layer6_outputs(5964)));
    outputs(5001) <= not(layer6_outputs(6215));
    outputs(5002) <= not((layer6_outputs(895)) and (layer6_outputs(1476)));
    outputs(5003) <= not(layer6_outputs(2309));
    outputs(5004) <= not(layer6_outputs(3180));
    outputs(5005) <= (layer6_outputs(341)) xor (layer6_outputs(1639));
    outputs(5006) <= not(layer6_outputs(5511));
    outputs(5007) <= layer6_outputs(6246);
    outputs(5008) <= not(layer6_outputs(7628));
    outputs(5009) <= layer6_outputs(3464);
    outputs(5010) <= layer6_outputs(1954);
    outputs(5011) <= (layer6_outputs(160)) xor (layer6_outputs(3571));
    outputs(5012) <= (layer6_outputs(6179)) and not (layer6_outputs(4484));
    outputs(5013) <= not(layer6_outputs(812));
    outputs(5014) <= not(layer6_outputs(7662));
    outputs(5015) <= layer6_outputs(166);
    outputs(5016) <= not((layer6_outputs(3405)) and (layer6_outputs(6660)));
    outputs(5017) <= not(layer6_outputs(4095));
    outputs(5018) <= (layer6_outputs(914)) and not (layer6_outputs(6765));
    outputs(5019) <= not(layer6_outputs(5428));
    outputs(5020) <= layer6_outputs(6182);
    outputs(5021) <= (layer6_outputs(7501)) and not (layer6_outputs(4092));
    outputs(5022) <= not(layer6_outputs(3964));
    outputs(5023) <= (layer6_outputs(4792)) and not (layer6_outputs(5155));
    outputs(5024) <= not(layer6_outputs(6106));
    outputs(5025) <= layer6_outputs(7483);
    outputs(5026) <= (layer6_outputs(5411)) and not (layer6_outputs(5154));
    outputs(5027) <= layer6_outputs(4365);
    outputs(5028) <= layer6_outputs(3973);
    outputs(5029) <= (layer6_outputs(6879)) xor (layer6_outputs(1521));
    outputs(5030) <= layer6_outputs(1376);
    outputs(5031) <= (layer6_outputs(3092)) and not (layer6_outputs(1932));
    outputs(5032) <= not((layer6_outputs(5550)) xor (layer6_outputs(2762)));
    outputs(5033) <= (layer6_outputs(7077)) and not (layer6_outputs(4263));
    outputs(5034) <= not(layer6_outputs(6908));
    outputs(5035) <= not(layer6_outputs(2863));
    outputs(5036) <= not(layer6_outputs(430));
    outputs(5037) <= layer6_outputs(4459);
    outputs(5038) <= (layer6_outputs(1408)) xor (layer6_outputs(425));
    outputs(5039) <= not(layer6_outputs(6793));
    outputs(5040) <= (layer6_outputs(1879)) xor (layer6_outputs(6516));
    outputs(5041) <= not((layer6_outputs(294)) xor (layer6_outputs(2834)));
    outputs(5042) <= not(layer6_outputs(7572));
    outputs(5043) <= not(layer6_outputs(1132));
    outputs(5044) <= not(layer6_outputs(1519));
    outputs(5045) <= (layer6_outputs(7270)) and not (layer6_outputs(1316));
    outputs(5046) <= layer6_outputs(1842);
    outputs(5047) <= layer6_outputs(1355);
    outputs(5048) <= not((layer6_outputs(7260)) xor (layer6_outputs(54)));
    outputs(5049) <= layer6_outputs(3527);
    outputs(5050) <= not(layer6_outputs(5035));
    outputs(5051) <= layer6_outputs(6844);
    outputs(5052) <= layer6_outputs(389);
    outputs(5053) <= not(layer6_outputs(93));
    outputs(5054) <= layer6_outputs(2644);
    outputs(5055) <= not(layer6_outputs(941));
    outputs(5056) <= not(layer6_outputs(4784));
    outputs(5057) <= (layer6_outputs(5039)) and not (layer6_outputs(963));
    outputs(5058) <= layer6_outputs(5777);
    outputs(5059) <= not(layer6_outputs(7488));
    outputs(5060) <= (layer6_outputs(665)) xor (layer6_outputs(2405));
    outputs(5061) <= not((layer6_outputs(1486)) or (layer6_outputs(5254)));
    outputs(5062) <= layer6_outputs(1768);
    outputs(5063) <= layer6_outputs(860);
    outputs(5064) <= layer6_outputs(4121);
    outputs(5065) <= not((layer6_outputs(7516)) xor (layer6_outputs(1951)));
    outputs(5066) <= layer6_outputs(3968);
    outputs(5067) <= layer6_outputs(5135);
    outputs(5068) <= not(layer6_outputs(2543));
    outputs(5069) <= layer6_outputs(443);
    outputs(5070) <= layer6_outputs(7562);
    outputs(5071) <= (layer6_outputs(3317)) xor (layer6_outputs(6668));
    outputs(5072) <= not((layer6_outputs(374)) or (layer6_outputs(2825)));
    outputs(5073) <= not((layer6_outputs(3807)) xor (layer6_outputs(3820)));
    outputs(5074) <= not(layer6_outputs(5861));
    outputs(5075) <= (layer6_outputs(2976)) xor (layer6_outputs(3281));
    outputs(5076) <= not(layer6_outputs(4681));
    outputs(5077) <= layer6_outputs(1406);
    outputs(5078) <= layer6_outputs(2141);
    outputs(5079) <= not((layer6_outputs(5276)) xor (layer6_outputs(5171)));
    outputs(5080) <= not(layer6_outputs(7071));
    outputs(5081) <= (layer6_outputs(4304)) xor (layer6_outputs(585));
    outputs(5082) <= (layer6_outputs(4330)) xor (layer6_outputs(2895));
    outputs(5083) <= (layer6_outputs(3567)) and (layer6_outputs(1234));
    outputs(5084) <= layer6_outputs(6257);
    outputs(5085) <= layer6_outputs(4690);
    outputs(5086) <= (layer6_outputs(4730)) xor (layer6_outputs(539));
    outputs(5087) <= not(layer6_outputs(4423));
    outputs(5088) <= not(layer6_outputs(1205));
    outputs(5089) <= layer6_outputs(1074);
    outputs(5090) <= (layer6_outputs(1097)) xor (layer6_outputs(5572));
    outputs(5091) <= not(layer6_outputs(2175));
    outputs(5092) <= not((layer6_outputs(1462)) xor (layer6_outputs(6355)));
    outputs(5093) <= (layer6_outputs(1298)) xor (layer6_outputs(4820));
    outputs(5094) <= not(layer6_outputs(1774));
    outputs(5095) <= not(layer6_outputs(2242));
    outputs(5096) <= not(layer6_outputs(4966));
    outputs(5097) <= layer6_outputs(4767);
    outputs(5098) <= not((layer6_outputs(4422)) and (layer6_outputs(676)));
    outputs(5099) <= (layer6_outputs(4975)) xor (layer6_outputs(6069));
    outputs(5100) <= not((layer6_outputs(337)) xor (layer6_outputs(4400)));
    outputs(5101) <= not(layer6_outputs(6750)) or (layer6_outputs(6427));
    outputs(5102) <= not((layer6_outputs(489)) xor (layer6_outputs(6581)));
    outputs(5103) <= layer6_outputs(6246);
    outputs(5104) <= not(layer6_outputs(5476)) or (layer6_outputs(769));
    outputs(5105) <= not(layer6_outputs(1485)) or (layer6_outputs(3356));
    outputs(5106) <= layer6_outputs(3506);
    outputs(5107) <= not(layer6_outputs(7526));
    outputs(5108) <= (layer6_outputs(3418)) or (layer6_outputs(7618));
    outputs(5109) <= (layer6_outputs(1676)) and (layer6_outputs(748));
    outputs(5110) <= layer6_outputs(5222);
    outputs(5111) <= layer6_outputs(1231);
    outputs(5112) <= layer6_outputs(1645);
    outputs(5113) <= not(layer6_outputs(1175));
    outputs(5114) <= not((layer6_outputs(2156)) or (layer6_outputs(5965)));
    outputs(5115) <= not(layer6_outputs(6434));
    outputs(5116) <= layer6_outputs(2040);
    outputs(5117) <= not(layer6_outputs(984));
    outputs(5118) <= not(layer6_outputs(4294));
    outputs(5119) <= (layer6_outputs(7394)) xor (layer6_outputs(5080));
    outputs(5120) <= (layer6_outputs(167)) and not (layer6_outputs(1013));
    outputs(5121) <= not(layer6_outputs(1729)) or (layer6_outputs(3496));
    outputs(5122) <= (layer6_outputs(4461)) xor (layer6_outputs(2033));
    outputs(5123) <= (layer6_outputs(5577)) and not (layer6_outputs(7094));
    outputs(5124) <= not(layer6_outputs(301));
    outputs(5125) <= not((layer6_outputs(392)) and (layer6_outputs(5336)));
    outputs(5126) <= not(layer6_outputs(5800));
    outputs(5127) <= not(layer6_outputs(4104));
    outputs(5128) <= not(layer6_outputs(2482));
    outputs(5129) <= not(layer6_outputs(5749));
    outputs(5130) <= not(layer6_outputs(3728));
    outputs(5131) <= (layer6_outputs(4430)) xor (layer6_outputs(1029));
    outputs(5132) <= layer6_outputs(1905);
    outputs(5133) <= layer6_outputs(2094);
    outputs(5134) <= not(layer6_outputs(2193));
    outputs(5135) <= not(layer6_outputs(7205));
    outputs(5136) <= layer6_outputs(4240);
    outputs(5137) <= not(layer6_outputs(6375));
    outputs(5138) <= layer6_outputs(2409);
    outputs(5139) <= not(layer6_outputs(4058));
    outputs(5140) <= not(layer6_outputs(2752));
    outputs(5141) <= (layer6_outputs(6283)) or (layer6_outputs(1093));
    outputs(5142) <= (layer6_outputs(1082)) and (layer6_outputs(3120));
    outputs(5143) <= layer6_outputs(6107);
    outputs(5144) <= not(layer6_outputs(4035));
    outputs(5145) <= layer6_outputs(4923);
    outputs(5146) <= (layer6_outputs(4683)) or (layer6_outputs(2723));
    outputs(5147) <= layer6_outputs(2733);
    outputs(5148) <= not((layer6_outputs(2828)) or (layer6_outputs(3614)));
    outputs(5149) <= layer6_outputs(4583);
    outputs(5150) <= layer6_outputs(1188);
    outputs(5151) <= layer6_outputs(2631);
    outputs(5152) <= not(layer6_outputs(842));
    outputs(5153) <= (layer6_outputs(3702)) xor (layer6_outputs(953));
    outputs(5154) <= (layer6_outputs(7044)) and not (layer6_outputs(4859));
    outputs(5155) <= layer6_outputs(2504);
    outputs(5156) <= layer6_outputs(264);
    outputs(5157) <= (layer6_outputs(2397)) xor (layer6_outputs(111));
    outputs(5158) <= (layer6_outputs(6689)) and (layer6_outputs(6577));
    outputs(5159) <= not(layer6_outputs(5200));
    outputs(5160) <= (layer6_outputs(885)) and not (layer6_outputs(5022));
    outputs(5161) <= layer6_outputs(4320);
    outputs(5162) <= not((layer6_outputs(5715)) xor (layer6_outputs(2763)));
    outputs(5163) <= layer6_outputs(4753);
    outputs(5164) <= layer6_outputs(1191);
    outputs(5165) <= not((layer6_outputs(3541)) or (layer6_outputs(6768)));
    outputs(5166) <= (layer6_outputs(2141)) and (layer6_outputs(5557));
    outputs(5167) <= (layer6_outputs(6652)) xor (layer6_outputs(657));
    outputs(5168) <= not((layer6_outputs(372)) and (layer6_outputs(6896)));
    outputs(5169) <= not(layer6_outputs(4894));
    outputs(5170) <= layer6_outputs(4493);
    outputs(5171) <= not((layer6_outputs(6905)) xor (layer6_outputs(3495)));
    outputs(5172) <= not(layer6_outputs(1793));
    outputs(5173) <= (layer6_outputs(6220)) and not (layer6_outputs(6465));
    outputs(5174) <= not(layer6_outputs(5855));
    outputs(5175) <= not(layer6_outputs(6969)) or (layer6_outputs(1532));
    outputs(5176) <= not(layer6_outputs(3934));
    outputs(5177) <= (layer6_outputs(5625)) and (layer6_outputs(7584));
    outputs(5178) <= (layer6_outputs(3882)) and not (layer6_outputs(7328));
    outputs(5179) <= layer6_outputs(3059);
    outputs(5180) <= not((layer6_outputs(6473)) xor (layer6_outputs(4537)));
    outputs(5181) <= (layer6_outputs(4948)) and not (layer6_outputs(5436));
    outputs(5182) <= (layer6_outputs(7604)) xor (layer6_outputs(6867));
    outputs(5183) <= layer6_outputs(4030);
    outputs(5184) <= layer6_outputs(3910);
    outputs(5185) <= layer6_outputs(2841);
    outputs(5186) <= layer6_outputs(5232);
    outputs(5187) <= layer6_outputs(6800);
    outputs(5188) <= layer6_outputs(894);
    outputs(5189) <= not((layer6_outputs(2706)) xor (layer6_outputs(7045)));
    outputs(5190) <= layer6_outputs(720);
    outputs(5191) <= (layer6_outputs(4656)) and not (layer6_outputs(2216));
    outputs(5192) <= not(layer6_outputs(3887));
    outputs(5193) <= not(layer6_outputs(4449));
    outputs(5194) <= layer6_outputs(4596);
    outputs(5195) <= layer6_outputs(5906);
    outputs(5196) <= not((layer6_outputs(2955)) or (layer6_outputs(853)));
    outputs(5197) <= layer6_outputs(977);
    outputs(5198) <= layer6_outputs(6576);
    outputs(5199) <= layer6_outputs(2649);
    outputs(5200) <= (layer6_outputs(4646)) xor (layer6_outputs(7125));
    outputs(5201) <= (layer6_outputs(510)) xor (layer6_outputs(2219));
    outputs(5202) <= not(layer6_outputs(7505));
    outputs(5203) <= (layer6_outputs(7365)) or (layer6_outputs(5078));
    outputs(5204) <= not(layer6_outputs(7585));
    outputs(5205) <= layer6_outputs(3324);
    outputs(5206) <= layer6_outputs(3130);
    outputs(5207) <= layer6_outputs(3946);
    outputs(5208) <= not((layer6_outputs(3380)) xor (layer6_outputs(2495)));
    outputs(5209) <= layer6_outputs(7556);
    outputs(5210) <= layer6_outputs(4014);
    outputs(5211) <= not(layer6_outputs(7175));
    outputs(5212) <= not(layer6_outputs(6625));
    outputs(5213) <= layer6_outputs(929);
    outputs(5214) <= layer6_outputs(4645);
    outputs(5215) <= (layer6_outputs(5751)) xor (layer6_outputs(89));
    outputs(5216) <= not((layer6_outputs(4433)) xor (layer6_outputs(7463)));
    outputs(5217) <= not(layer6_outputs(3280));
    outputs(5218) <= not(layer6_outputs(6386));
    outputs(5219) <= (layer6_outputs(5988)) and not (layer6_outputs(1192));
    outputs(5220) <= layer6_outputs(1702);
    outputs(5221) <= not((layer6_outputs(917)) or (layer6_outputs(4012)));
    outputs(5222) <= not((layer6_outputs(4383)) xor (layer6_outputs(5691)));
    outputs(5223) <= (layer6_outputs(3915)) xor (layer6_outputs(5002));
    outputs(5224) <= layer6_outputs(5602);
    outputs(5225) <= not(layer6_outputs(2118));
    outputs(5226) <= not(layer6_outputs(7209));
    outputs(5227) <= (layer6_outputs(5114)) and (layer6_outputs(1740));
    outputs(5228) <= (layer6_outputs(5622)) xor (layer6_outputs(3233));
    outputs(5229) <= (layer6_outputs(5142)) xor (layer6_outputs(1337));
    outputs(5230) <= not((layer6_outputs(7144)) or (layer6_outputs(6133)));
    outputs(5231) <= layer6_outputs(2644);
    outputs(5232) <= layer6_outputs(4960);
    outputs(5233) <= layer6_outputs(6731);
    outputs(5234) <= layer6_outputs(5019);
    outputs(5235) <= layer6_outputs(2260);
    outputs(5236) <= not(layer6_outputs(3750)) or (layer6_outputs(1333));
    outputs(5237) <= layer6_outputs(937);
    outputs(5238) <= layer6_outputs(943);
    outputs(5239) <= not(layer6_outputs(1593));
    outputs(5240) <= not((layer6_outputs(2705)) xor (layer6_outputs(221)));
    outputs(5241) <= (layer6_outputs(3048)) and not (layer6_outputs(7295));
    outputs(5242) <= not(layer6_outputs(1966));
    outputs(5243) <= not(layer6_outputs(6134));
    outputs(5244) <= (layer6_outputs(3299)) xor (layer6_outputs(6544));
    outputs(5245) <= layer6_outputs(3398);
    outputs(5246) <= layer6_outputs(5838);
    outputs(5247) <= layer6_outputs(4227);
    outputs(5248) <= (layer6_outputs(3802)) xor (layer6_outputs(3095));
    outputs(5249) <= not(layer6_outputs(5744));
    outputs(5250) <= layer6_outputs(3292);
    outputs(5251) <= not(layer6_outputs(1373));
    outputs(5252) <= not((layer6_outputs(5080)) xor (layer6_outputs(2818)));
    outputs(5253) <= layer6_outputs(6500);
    outputs(5254) <= layer6_outputs(5927);
    outputs(5255) <= not(layer6_outputs(7374));
    outputs(5256) <= not((layer6_outputs(4643)) xor (layer6_outputs(6794)));
    outputs(5257) <= (layer6_outputs(7117)) and not (layer6_outputs(5131));
    outputs(5258) <= not(layer6_outputs(1086));
    outputs(5259) <= layer6_outputs(6860);
    outputs(5260) <= layer6_outputs(2970);
    outputs(5261) <= layer6_outputs(2832);
    outputs(5262) <= (layer6_outputs(4972)) and not (layer6_outputs(2873));
    outputs(5263) <= not(layer6_outputs(2032));
    outputs(5264) <= (layer6_outputs(6523)) and not (layer6_outputs(5633));
    outputs(5265) <= (layer6_outputs(1089)) and (layer6_outputs(4673));
    outputs(5266) <= layer6_outputs(678);
    outputs(5267) <= not(layer6_outputs(4299));
    outputs(5268) <= layer6_outputs(1960);
    outputs(5269) <= (layer6_outputs(2395)) and not (layer6_outputs(3248));
    outputs(5270) <= not(layer6_outputs(3737));
    outputs(5271) <= layer6_outputs(7487);
    outputs(5272) <= not(layer6_outputs(2003));
    outputs(5273) <= (layer6_outputs(3586)) and not (layer6_outputs(6727));
    outputs(5274) <= not(layer6_outputs(7670));
    outputs(5275) <= layer6_outputs(399);
    outputs(5276) <= not(layer6_outputs(7208));
    outputs(5277) <= not(layer6_outputs(2074));
    outputs(5278) <= not((layer6_outputs(7631)) xor (layer6_outputs(1904)));
    outputs(5279) <= not((layer6_outputs(7345)) xor (layer6_outputs(7395)));
    outputs(5280) <= layer6_outputs(3371);
    outputs(5281) <= layer6_outputs(777);
    outputs(5282) <= not(layer6_outputs(7142));
    outputs(5283) <= not((layer6_outputs(3376)) or (layer6_outputs(3245)));
    outputs(5284) <= layer6_outputs(3282);
    outputs(5285) <= not(layer6_outputs(7628));
    outputs(5286) <= not((layer6_outputs(5312)) or (layer6_outputs(6298)));
    outputs(5287) <= not(layer6_outputs(4349));
    outputs(5288) <= layer6_outputs(4493);
    outputs(5289) <= (layer6_outputs(473)) xor (layer6_outputs(1340));
    outputs(5290) <= not(layer6_outputs(580));
    outputs(5291) <= (layer6_outputs(700)) and not (layer6_outputs(4828));
    outputs(5292) <= not(layer6_outputs(6386));
    outputs(5293) <= (layer6_outputs(2770)) and (layer6_outputs(1099));
    outputs(5294) <= not((layer6_outputs(3047)) and (layer6_outputs(2184)));
    outputs(5295) <= layer6_outputs(3096);
    outputs(5296) <= layer6_outputs(2100);
    outputs(5297) <= not(layer6_outputs(4949));
    outputs(5298) <= not(layer6_outputs(535));
    outputs(5299) <= not(layer6_outputs(5164));
    outputs(5300) <= (layer6_outputs(3658)) and not (layer6_outputs(529));
    outputs(5301) <= (layer6_outputs(4317)) xor (layer6_outputs(5249));
    outputs(5302) <= (layer6_outputs(3735)) and not (layer6_outputs(6823));
    outputs(5303) <= not(layer6_outputs(450));
    outputs(5304) <= not(layer6_outputs(6004));
    outputs(5305) <= (layer6_outputs(5629)) and not (layer6_outputs(3791));
    outputs(5306) <= (layer6_outputs(5525)) xor (layer6_outputs(1485));
    outputs(5307) <= (layer6_outputs(7541)) or (layer6_outputs(6376));
    outputs(5308) <= not(layer6_outputs(921)) or (layer6_outputs(2634));
    outputs(5309) <= (layer6_outputs(2989)) xor (layer6_outputs(3374));
    outputs(5310) <= layer6_outputs(5269);
    outputs(5311) <= not((layer6_outputs(5435)) or (layer6_outputs(6988)));
    outputs(5312) <= layer6_outputs(2110);
    outputs(5313) <= layer6_outputs(4874);
    outputs(5314) <= (layer6_outputs(6776)) xor (layer6_outputs(5634));
    outputs(5315) <= not(layer6_outputs(1199));
    outputs(5316) <= layer6_outputs(3049);
    outputs(5317) <= (layer6_outputs(7350)) xor (layer6_outputs(1852));
    outputs(5318) <= not((layer6_outputs(3917)) xor (layer6_outputs(6939)));
    outputs(5319) <= not(layer6_outputs(2287));
    outputs(5320) <= layer6_outputs(739);
    outputs(5321) <= layer6_outputs(1762);
    outputs(5322) <= not(layer6_outputs(6904));
    outputs(5323) <= layer6_outputs(4644);
    outputs(5324) <= not(layer6_outputs(5390));
    outputs(5325) <= layer6_outputs(6379);
    outputs(5326) <= not((layer6_outputs(1881)) xor (layer6_outputs(549)));
    outputs(5327) <= layer6_outputs(3673);
    outputs(5328) <= not((layer6_outputs(1595)) xor (layer6_outputs(2560)));
    outputs(5329) <= not((layer6_outputs(2525)) xor (layer6_outputs(49)));
    outputs(5330) <= (layer6_outputs(6626)) and not (layer6_outputs(7424));
    outputs(5331) <= not(layer6_outputs(3504));
    outputs(5332) <= layer6_outputs(846);
    outputs(5333) <= layer6_outputs(6343);
    outputs(5334) <= not(layer6_outputs(7264));
    outputs(5335) <= not(layer6_outputs(4863));
    outputs(5336) <= not(layer6_outputs(2690));
    outputs(5337) <= layer6_outputs(3201);
    outputs(5338) <= (layer6_outputs(3978)) xor (layer6_outputs(4221));
    outputs(5339) <= layer6_outputs(4775);
    outputs(5340) <= layer6_outputs(2209);
    outputs(5341) <= not(layer6_outputs(5153));
    outputs(5342) <= layer6_outputs(4916);
    outputs(5343) <= not(layer6_outputs(5466));
    outputs(5344) <= layer6_outputs(7193);
    outputs(5345) <= (layer6_outputs(4696)) xor (layer6_outputs(5299));
    outputs(5346) <= not(layer6_outputs(4884));
    outputs(5347) <= (layer6_outputs(582)) and (layer6_outputs(1076));
    outputs(5348) <= layer6_outputs(5197);
    outputs(5349) <= layer6_outputs(3400);
    outputs(5350) <= layer6_outputs(7484);
    outputs(5351) <= (layer6_outputs(3528)) and not (layer6_outputs(2038));
    outputs(5352) <= (layer6_outputs(3685)) xor (layer6_outputs(3075));
    outputs(5353) <= layer6_outputs(362);
    outputs(5354) <= layer6_outputs(1500);
    outputs(5355) <= not(layer6_outputs(3455)) or (layer6_outputs(4225));
    outputs(5356) <= not((layer6_outputs(1955)) xor (layer6_outputs(6636)));
    outputs(5357) <= (layer6_outputs(164)) and (layer6_outputs(6990));
    outputs(5358) <= layer6_outputs(4618);
    outputs(5359) <= not(layer6_outputs(1266));
    outputs(5360) <= not(layer6_outputs(2493)) or (layer6_outputs(7648));
    outputs(5361) <= not(layer6_outputs(831));
    outputs(5362) <= not(layer6_outputs(344));
    outputs(5363) <= not(layer6_outputs(2485));
    outputs(5364) <= (layer6_outputs(3817)) xor (layer6_outputs(2071));
    outputs(5365) <= not(layer6_outputs(2903));
    outputs(5366) <= not(layer6_outputs(458));
    outputs(5367) <= not(layer6_outputs(2085));
    outputs(5368) <= not(layer6_outputs(186));
    outputs(5369) <= not(layer6_outputs(6208));
    outputs(5370) <= not(layer6_outputs(2977));
    outputs(5371) <= not((layer6_outputs(5212)) xor (layer6_outputs(2179)));
    outputs(5372) <= (layer6_outputs(6778)) xor (layer6_outputs(2213));
    outputs(5373) <= layer6_outputs(4462);
    outputs(5374) <= layer6_outputs(7275);
    outputs(5375) <= layer6_outputs(2187);
    outputs(5376) <= layer6_outputs(1906);
    outputs(5377) <= layer6_outputs(2682);
    outputs(5378) <= not(layer6_outputs(1474));
    outputs(5379) <= layer6_outputs(2144);
    outputs(5380) <= not(layer6_outputs(376));
    outputs(5381) <= not(layer6_outputs(4011));
    outputs(5382) <= not(layer6_outputs(6214));
    outputs(5383) <= not(layer6_outputs(7297));
    outputs(5384) <= layer6_outputs(2896);
    outputs(5385) <= not(layer6_outputs(3695));
    outputs(5386) <= not((layer6_outputs(3278)) xor (layer6_outputs(3926)));
    outputs(5387) <= layer6_outputs(1582);
    outputs(5388) <= layer6_outputs(2913);
    outputs(5389) <= layer6_outputs(501);
    outputs(5390) <= not(layer6_outputs(7268));
    outputs(5391) <= not(layer6_outputs(1853));
    outputs(5392) <= not((layer6_outputs(1641)) or (layer6_outputs(7605)));
    outputs(5393) <= not(layer6_outputs(1585));
    outputs(5394) <= layer6_outputs(5370);
    outputs(5395) <= layer6_outputs(37);
    outputs(5396) <= (layer6_outputs(3097)) and not (layer6_outputs(704));
    outputs(5397) <= (layer6_outputs(6841)) and (layer6_outputs(1830));
    outputs(5398) <= not(layer6_outputs(2817));
    outputs(5399) <= not(layer6_outputs(3919));
    outputs(5400) <= not(layer6_outputs(956));
    outputs(5401) <= (layer6_outputs(2525)) and (layer6_outputs(1227));
    outputs(5402) <= not(layer6_outputs(4613));
    outputs(5403) <= not(layer6_outputs(6688));
    outputs(5404) <= (layer6_outputs(3218)) xor (layer6_outputs(852));
    outputs(5405) <= (layer6_outputs(179)) and not (layer6_outputs(7639));
    outputs(5406) <= layer6_outputs(2371);
    outputs(5407) <= not(layer6_outputs(3369));
    outputs(5408) <= layer6_outputs(6186);
    outputs(5409) <= not(layer6_outputs(5169));
    outputs(5410) <= not((layer6_outputs(490)) xor (layer6_outputs(3604)));
    outputs(5411) <= (layer6_outputs(2201)) and (layer6_outputs(5320));
    outputs(5412) <= not((layer6_outputs(6659)) or (layer6_outputs(5843)));
    outputs(5413) <= not(layer6_outputs(7359));
    outputs(5414) <= not((layer6_outputs(5242)) or (layer6_outputs(945)));
    outputs(5415) <= layer6_outputs(4414);
    outputs(5416) <= not(layer6_outputs(731));
    outputs(5417) <= not(layer6_outputs(1257));
    outputs(5418) <= not(layer6_outputs(442));
    outputs(5419) <= not(layer6_outputs(796));
    outputs(5420) <= layer6_outputs(269);
    outputs(5421) <= not(layer6_outputs(6811)) or (layer6_outputs(1053));
    outputs(5422) <= not(layer6_outputs(4538));
    outputs(5423) <= not((layer6_outputs(839)) xor (layer6_outputs(1051)));
    outputs(5424) <= not(layer6_outputs(1685)) or (layer6_outputs(790));
    outputs(5425) <= layer6_outputs(5633);
    outputs(5426) <= not(layer6_outputs(4389));
    outputs(5427) <= not((layer6_outputs(5071)) xor (layer6_outputs(2540)));
    outputs(5428) <= not(layer6_outputs(2760)) or (layer6_outputs(1506));
    outputs(5429) <= not((layer6_outputs(3330)) or (layer6_outputs(380)));
    outputs(5430) <= layer6_outputs(6833);
    outputs(5431) <= (layer6_outputs(6936)) and not (layer6_outputs(2192));
    outputs(5432) <= (layer6_outputs(1889)) xor (layer6_outputs(2400));
    outputs(5433) <= layer6_outputs(2603);
    outputs(5434) <= not((layer6_outputs(1992)) xor (layer6_outputs(5984)));
    outputs(5435) <= not(layer6_outputs(7256));
    outputs(5436) <= (layer6_outputs(2325)) xor (layer6_outputs(3302));
    outputs(5437) <= not(layer6_outputs(1924)) or (layer6_outputs(6774));
    outputs(5438) <= not((layer6_outputs(2122)) xor (layer6_outputs(5898)));
    outputs(5439) <= not(layer6_outputs(3374));
    outputs(5440) <= not(layer6_outputs(3028));
    outputs(5441) <= (layer6_outputs(3136)) and (layer6_outputs(6940));
    outputs(5442) <= layer6_outputs(2357);
    outputs(5443) <= layer6_outputs(3113);
    outputs(5444) <= not(layer6_outputs(1099)) or (layer6_outputs(1635));
    outputs(5445) <= layer6_outputs(4819);
    outputs(5446) <= layer6_outputs(4856);
    outputs(5447) <= (layer6_outputs(4905)) xor (layer6_outputs(4999));
    outputs(5448) <= (layer6_outputs(1818)) or (layer6_outputs(176));
    outputs(5449) <= layer6_outputs(6633);
    outputs(5450) <= layer6_outputs(7524);
    outputs(5451) <= layer6_outputs(6886);
    outputs(5452) <= layer6_outputs(5358);
    outputs(5453) <= (layer6_outputs(1009)) xor (layer6_outputs(5861));
    outputs(5454) <= not((layer6_outputs(4054)) or (layer6_outputs(6401)));
    outputs(5455) <= (layer6_outputs(2539)) xor (layer6_outputs(6001));
    outputs(5456) <= layer6_outputs(5223);
    outputs(5457) <= not((layer6_outputs(6698)) xor (layer6_outputs(4643)));
    outputs(5458) <= not((layer6_outputs(3622)) xor (layer6_outputs(327)));
    outputs(5459) <= (layer6_outputs(2877)) and not (layer6_outputs(2102));
    outputs(5460) <= not(layer6_outputs(6918));
    outputs(5461) <= not(layer6_outputs(2756));
    outputs(5462) <= not(layer6_outputs(2103));
    outputs(5463) <= not(layer6_outputs(4553));
    outputs(5464) <= layer6_outputs(4706);
    outputs(5465) <= not(layer6_outputs(4838));
    outputs(5466) <= (layer6_outputs(1111)) and not (layer6_outputs(2745));
    outputs(5467) <= (layer6_outputs(1824)) xor (layer6_outputs(3473));
    outputs(5468) <= layer6_outputs(3815);
    outputs(5469) <= (layer6_outputs(2896)) xor (layer6_outputs(4579));
    outputs(5470) <= not(layer6_outputs(2146));
    outputs(5471) <= not((layer6_outputs(4662)) xor (layer6_outputs(5150)));
    outputs(5472) <= not(layer6_outputs(3650));
    outputs(5473) <= layer6_outputs(7097);
    outputs(5474) <= not(layer6_outputs(6566));
    outputs(5475) <= not((layer6_outputs(3573)) xor (layer6_outputs(5094)));
    outputs(5476) <= not((layer6_outputs(1979)) xor (layer6_outputs(2200)));
    outputs(5477) <= not(layer6_outputs(986));
    outputs(5478) <= not(layer6_outputs(7384));
    outputs(5479) <= layer6_outputs(5842);
    outputs(5480) <= not(layer6_outputs(5032));
    outputs(5481) <= layer6_outputs(5305);
    outputs(5482) <= layer6_outputs(6315);
    outputs(5483) <= not((layer6_outputs(2907)) or (layer6_outputs(7339)));
    outputs(5484) <= layer6_outputs(5075);
    outputs(5485) <= layer6_outputs(4238);
    outputs(5486) <= layer6_outputs(461);
    outputs(5487) <= not(layer6_outputs(2520));
    outputs(5488) <= layer6_outputs(6699);
    outputs(5489) <= not(layer6_outputs(3424));
    outputs(5490) <= not(layer6_outputs(756));
    outputs(5491) <= layer6_outputs(5847);
    outputs(5492) <= not((layer6_outputs(6741)) xor (layer6_outputs(2655)));
    outputs(5493) <= layer6_outputs(5707);
    outputs(5494) <= not(layer6_outputs(3360));
    outputs(5495) <= layer6_outputs(128);
    outputs(5496) <= layer6_outputs(7401);
    outputs(5497) <= layer6_outputs(1327);
    outputs(5498) <= not(layer6_outputs(5996));
    outputs(5499) <= layer6_outputs(1777);
    outputs(5500) <= not(layer6_outputs(4547));
    outputs(5501) <= not(layer6_outputs(5860));
    outputs(5502) <= not(layer6_outputs(6998));
    outputs(5503) <= not(layer6_outputs(4042));
    outputs(5504) <= layer6_outputs(3133);
    outputs(5505) <= not(layer6_outputs(159));
    outputs(5506) <= not((layer6_outputs(4360)) xor (layer6_outputs(621)));
    outputs(5507) <= not(layer6_outputs(2284));
    outputs(5508) <= layer6_outputs(4403);
    outputs(5509) <= not(layer6_outputs(1841));
    outputs(5510) <= (layer6_outputs(3436)) xor (layer6_outputs(2744));
    outputs(5511) <= not(layer6_outputs(5768)) or (layer6_outputs(454));
    outputs(5512) <= not((layer6_outputs(7041)) and (layer6_outputs(5939)));
    outputs(5513) <= not(layer6_outputs(4572));
    outputs(5514) <= not(layer6_outputs(1548));
    outputs(5515) <= not(layer6_outputs(1129)) or (layer6_outputs(5701));
    outputs(5516) <= not(layer6_outputs(270));
    outputs(5517) <= not((layer6_outputs(3698)) or (layer6_outputs(3300)));
    outputs(5518) <= (layer6_outputs(1853)) xor (layer6_outputs(1054));
    outputs(5519) <= (layer6_outputs(4687)) xor (layer6_outputs(2041));
    outputs(5520) <= layer6_outputs(2993);
    outputs(5521) <= not(layer6_outputs(1618));
    outputs(5522) <= not(layer6_outputs(4297));
    outputs(5523) <= (layer6_outputs(3871)) and (layer6_outputs(1752));
    outputs(5524) <= not((layer6_outputs(5836)) and (layer6_outputs(4056)));
    outputs(5525) <= layer6_outputs(1804);
    outputs(5526) <= layer6_outputs(7122);
    outputs(5527) <= not((layer6_outputs(941)) and (layer6_outputs(2162)));
    outputs(5528) <= layer6_outputs(6438);
    outputs(5529) <= layer6_outputs(3062);
    outputs(5530) <= layer6_outputs(3211);
    outputs(5531) <= not(layer6_outputs(3343));
    outputs(5532) <= not(layer6_outputs(2149));
    outputs(5533) <= (layer6_outputs(6535)) and not (layer6_outputs(5103));
    outputs(5534) <= not(layer6_outputs(217));
    outputs(5535) <= (layer6_outputs(3114)) xor (layer6_outputs(6711));
    outputs(5536) <= not(layer6_outputs(507));
    outputs(5537) <= not(layer6_outputs(4011));
    outputs(5538) <= not((layer6_outputs(210)) xor (layer6_outputs(2876)));
    outputs(5539) <= (layer6_outputs(5545)) and not (layer6_outputs(2326));
    outputs(5540) <= not((layer6_outputs(3408)) xor (layer6_outputs(6943)));
    outputs(5541) <= not(layer6_outputs(5352));
    outputs(5542) <= (layer6_outputs(7566)) xor (layer6_outputs(385));
    outputs(5543) <= not((layer6_outputs(4660)) xor (layer6_outputs(3350)));
    outputs(5544) <= not(layer6_outputs(6161));
    outputs(5545) <= layer6_outputs(2800);
    outputs(5546) <= layer6_outputs(1159);
    outputs(5547) <= not(layer6_outputs(5065)) or (layer6_outputs(3578));
    outputs(5548) <= not(layer6_outputs(6302));
    outputs(5549) <= layer6_outputs(123);
    outputs(5550) <= not(layer6_outputs(4961));
    outputs(5551) <= not(layer6_outputs(1077));
    outputs(5552) <= layer6_outputs(2906);
    outputs(5553) <= layer6_outputs(1637);
    outputs(5554) <= layer6_outputs(479);
    outputs(5555) <= layer6_outputs(379);
    outputs(5556) <= (layer6_outputs(2678)) and (layer6_outputs(4943));
    outputs(5557) <= not(layer6_outputs(7383));
    outputs(5558) <= not((layer6_outputs(4016)) xor (layer6_outputs(1709)));
    outputs(5559) <= not((layer6_outputs(5126)) xor (layer6_outputs(90)));
    outputs(5560) <= not(layer6_outputs(5859));
    outputs(5561) <= layer6_outputs(3795);
    outputs(5562) <= not((layer6_outputs(4346)) or (layer6_outputs(2274)));
    outputs(5563) <= layer6_outputs(6413);
    outputs(5564) <= not(layer6_outputs(2918));
    outputs(5565) <= layer6_outputs(1348);
    outputs(5566) <= layer6_outputs(4511);
    outputs(5567) <= (layer6_outputs(7017)) and (layer6_outputs(3568));
    outputs(5568) <= (layer6_outputs(2369)) and (layer6_outputs(257));
    outputs(5569) <= layer6_outputs(3550);
    outputs(5570) <= not((layer6_outputs(2416)) or (layer6_outputs(5222)));
    outputs(5571) <= not(layer6_outputs(5737));
    outputs(5572) <= layer6_outputs(4758);
    outputs(5573) <= not((layer6_outputs(4600)) or (layer6_outputs(5784)));
    outputs(5574) <= layer6_outputs(2775);
    outputs(5575) <= layer6_outputs(642);
    outputs(5576) <= not((layer6_outputs(7132)) xor (layer6_outputs(3366)));
    outputs(5577) <= not(layer6_outputs(214));
    outputs(5578) <= (layer6_outputs(5934)) and not (layer6_outputs(4684));
    outputs(5579) <= not(layer6_outputs(3317));
    outputs(5580) <= (layer6_outputs(3009)) or (layer6_outputs(673));
    outputs(5581) <= not((layer6_outputs(2852)) or (layer6_outputs(4352)));
    outputs(5582) <= not(layer6_outputs(3989)) or (layer6_outputs(503));
    outputs(5583) <= layer6_outputs(6595);
    outputs(5584) <= not(layer6_outputs(5581));
    outputs(5585) <= not(layer6_outputs(4185));
    outputs(5586) <= (layer6_outputs(1528)) or (layer6_outputs(1102));
    outputs(5587) <= layer6_outputs(3426);
    outputs(5588) <= not(layer6_outputs(1797));
    outputs(5589) <= not(layer6_outputs(6370));
    outputs(5590) <= not(layer6_outputs(1070));
    outputs(5591) <= layer6_outputs(2349);
    outputs(5592) <= layer6_outputs(5443);
    outputs(5593) <= (layer6_outputs(7132)) and (layer6_outputs(2097));
    outputs(5594) <= not((layer6_outputs(2766)) and (layer6_outputs(1577)));
    outputs(5595) <= layer6_outputs(5913);
    outputs(5596) <= not((layer6_outputs(2399)) or (layer6_outputs(6189)));
    outputs(5597) <= not(layer6_outputs(3134));
    outputs(5598) <= not((layer6_outputs(2223)) xor (layer6_outputs(2098)));
    outputs(5599) <= layer6_outputs(4401);
    outputs(5600) <= layer6_outputs(6634);
    outputs(5601) <= not(layer6_outputs(1677));
    outputs(5602) <= (layer6_outputs(2281)) xor (layer6_outputs(10));
    outputs(5603) <= layer6_outputs(5382);
    outputs(5604) <= not(layer6_outputs(4101));
    outputs(5605) <= (layer6_outputs(691)) xor (layer6_outputs(5788));
    outputs(5606) <= (layer6_outputs(2002)) or (layer6_outputs(4742));
    outputs(5607) <= layer6_outputs(5498);
    outputs(5608) <= not(layer6_outputs(3493));
    outputs(5609) <= not(layer6_outputs(2410));
    outputs(5610) <= not(layer6_outputs(1992));
    outputs(5611) <= (layer6_outputs(3999)) and not (layer6_outputs(5405));
    outputs(5612) <= not(layer6_outputs(2513)) or (layer6_outputs(4478));
    outputs(5613) <= layer6_outputs(4126);
    outputs(5614) <= (layer6_outputs(6032)) or (layer6_outputs(3478));
    outputs(5615) <= not((layer6_outputs(6198)) and (layer6_outputs(6313)));
    outputs(5616) <= layer6_outputs(3640);
    outputs(5617) <= layer6_outputs(1052);
    outputs(5618) <= layer6_outputs(4375);
    outputs(5619) <= not(layer6_outputs(58));
    outputs(5620) <= (layer6_outputs(2994)) and (layer6_outputs(5447));
    outputs(5621) <= (layer6_outputs(1755)) and not (layer6_outputs(7014));
    outputs(5622) <= not(layer6_outputs(3793));
    outputs(5623) <= not(layer6_outputs(5259));
    outputs(5624) <= (layer6_outputs(4781)) and (layer6_outputs(6232));
    outputs(5625) <= layer6_outputs(4824);
    outputs(5626) <= layer6_outputs(2665);
    outputs(5627) <= not((layer6_outputs(6234)) xor (layer6_outputs(2573)));
    outputs(5628) <= not(layer6_outputs(3285));
    outputs(5629) <= layer6_outputs(7531);
    outputs(5630) <= layer6_outputs(2740);
    outputs(5631) <= not(layer6_outputs(2932));
    outputs(5632) <= (layer6_outputs(2648)) xor (layer6_outputs(3939));
    outputs(5633) <= layer6_outputs(3504);
    outputs(5634) <= layer6_outputs(791);
    outputs(5635) <= (layer6_outputs(2885)) xor (layer6_outputs(2407));
    outputs(5636) <= not((layer6_outputs(6203)) xor (layer6_outputs(5360)));
    outputs(5637) <= not(layer6_outputs(6092));
    outputs(5638) <= layer6_outputs(4769);
    outputs(5639) <= (layer6_outputs(6008)) and (layer6_outputs(1908));
    outputs(5640) <= not(layer6_outputs(5747));
    outputs(5641) <= not(layer6_outputs(3956));
    outputs(5642) <= layer6_outputs(2134);
    outputs(5643) <= layer6_outputs(6465);
    outputs(5644) <= (layer6_outputs(7418)) and not (layer6_outputs(1610));
    outputs(5645) <= (layer6_outputs(2177)) and not (layer6_outputs(6847));
    outputs(5646) <= not((layer6_outputs(2535)) or (layer6_outputs(846)));
    outputs(5647) <= not((layer6_outputs(719)) xor (layer6_outputs(5017)));
    outputs(5648) <= (layer6_outputs(3450)) xor (layer6_outputs(2240));
    outputs(5649) <= not(layer6_outputs(2671));
    outputs(5650) <= not(layer6_outputs(562));
    outputs(5651) <= not(layer6_outputs(6288));
    outputs(5652) <= (layer6_outputs(2116)) or (layer6_outputs(7362));
    outputs(5653) <= layer6_outputs(1808);
    outputs(5654) <= layer6_outputs(591);
    outputs(5655) <= layer6_outputs(5688);
    outputs(5656) <= layer6_outputs(3996);
    outputs(5657) <= (layer6_outputs(133)) xor (layer6_outputs(4513));
    outputs(5658) <= not(layer6_outputs(5029));
    outputs(5659) <= layer6_outputs(3034);
    outputs(5660) <= not(layer6_outputs(7470));
    outputs(5661) <= layer6_outputs(2278);
    outputs(5662) <= layer6_outputs(17);
    outputs(5663) <= not((layer6_outputs(6819)) xor (layer6_outputs(3826)));
    outputs(5664) <= not(layer6_outputs(1577));
    outputs(5665) <= not(layer6_outputs(4034));
    outputs(5666) <= not((layer6_outputs(1819)) xor (layer6_outputs(6884)));
    outputs(5667) <= not((layer6_outputs(3802)) xor (layer6_outputs(2677)));
    outputs(5668) <= layer6_outputs(4783);
    outputs(5669) <= not(layer6_outputs(3252));
    outputs(5670) <= layer6_outputs(4450);
    outputs(5671) <= (layer6_outputs(7035)) and not (layer6_outputs(4559));
    outputs(5672) <= (layer6_outputs(7603)) or (layer6_outputs(1874));
    outputs(5673) <= not(layer6_outputs(2660));
    outputs(5674) <= not((layer6_outputs(4262)) xor (layer6_outputs(7661)));
    outputs(5675) <= layer6_outputs(3560);
    outputs(5676) <= (layer6_outputs(5121)) or (layer6_outputs(136));
    outputs(5677) <= layer6_outputs(850);
    outputs(5678) <= (layer6_outputs(5601)) xor (layer6_outputs(4623));
    outputs(5679) <= not(layer6_outputs(4849));
    outputs(5680) <= not(layer6_outputs(4947));
    outputs(5681) <= not(layer6_outputs(2674));
    outputs(5682) <= layer6_outputs(1347);
    outputs(5683) <= layer6_outputs(4882);
    outputs(5684) <= not(layer6_outputs(6479)) or (layer6_outputs(6763));
    outputs(5685) <= not(layer6_outputs(27));
    outputs(5686) <= not(layer6_outputs(46));
    outputs(5687) <= not((layer6_outputs(1282)) xor (layer6_outputs(3166)));
    outputs(5688) <= not(layer6_outputs(2694));
    outputs(5689) <= not(layer6_outputs(7348));
    outputs(5690) <= (layer6_outputs(7141)) xor (layer6_outputs(5246));
    outputs(5691) <= (layer6_outputs(6982)) xor (layer6_outputs(5065));
    outputs(5692) <= not(layer6_outputs(5728));
    outputs(5693) <= not(layer6_outputs(3026));
    outputs(5694) <= not(layer6_outputs(2881)) or (layer6_outputs(1327));
    outputs(5695) <= (layer6_outputs(4445)) and not (layer6_outputs(4467));
    outputs(5696) <= not(layer6_outputs(5144));
    outputs(5697) <= (layer6_outputs(3257)) and (layer6_outputs(622));
    outputs(5698) <= not(layer6_outputs(4431));
    outputs(5699) <= (layer6_outputs(5949)) and not (layer6_outputs(4780));
    outputs(5700) <= layer6_outputs(1147);
    outputs(5701) <= (layer6_outputs(2747)) xor (layer6_outputs(5983));
    outputs(5702) <= layer6_outputs(709);
    outputs(5703) <= not(layer6_outputs(3003)) or (layer6_outputs(6445));
    outputs(5704) <= (layer6_outputs(1661)) xor (layer6_outputs(6600));
    outputs(5705) <= layer6_outputs(5087);
    outputs(5706) <= not(layer6_outputs(1614));
    outputs(5707) <= (layer6_outputs(4149)) xor (layer6_outputs(1301));
    outputs(5708) <= layer6_outputs(4087);
    outputs(5709) <= not((layer6_outputs(2811)) xor (layer6_outputs(208)));
    outputs(5710) <= layer6_outputs(1596);
    outputs(5711) <= (layer6_outputs(7646)) xor (layer6_outputs(4147));
    outputs(5712) <= (layer6_outputs(4512)) and (layer6_outputs(3098));
    outputs(5713) <= not(layer6_outputs(1409));
    outputs(5714) <= (layer6_outputs(5570)) and (layer6_outputs(6728));
    outputs(5715) <= layer6_outputs(3451);
    outputs(5716) <= (layer6_outputs(3835)) and not (layer6_outputs(4562));
    outputs(5717) <= layer6_outputs(3672);
    outputs(5718) <= not(layer6_outputs(6903));
    outputs(5719) <= layer6_outputs(6256);
    outputs(5720) <= not((layer6_outputs(5699)) xor (layer6_outputs(4282)));
    outputs(5721) <= layer6_outputs(5766);
    outputs(5722) <= not((layer6_outputs(5007)) xor (layer6_outputs(6965)));
    outputs(5723) <= not(layer6_outputs(5935));
    outputs(5724) <= not(layer6_outputs(6258));
    outputs(5725) <= not(layer6_outputs(3937));
    outputs(5726) <= not(layer6_outputs(2291));
    outputs(5727) <= not(layer6_outputs(3440));
    outputs(5728) <= not(layer6_outputs(7481));
    outputs(5729) <= (layer6_outputs(7229)) and not (layer6_outputs(181));
    outputs(5730) <= (layer6_outputs(6164)) and not (layer6_outputs(5186));
    outputs(5731) <= not((layer6_outputs(262)) xor (layer6_outputs(1810)));
    outputs(5732) <= (layer6_outputs(4013)) xor (layer6_outputs(7647));
    outputs(5733) <= not(layer6_outputs(914));
    outputs(5734) <= not(layer6_outputs(4022));
    outputs(5735) <= layer6_outputs(1637);
    outputs(5736) <= not((layer6_outputs(1878)) xor (layer6_outputs(5883)));
    outputs(5737) <= not(layer6_outputs(1618));
    outputs(5738) <= not(layer6_outputs(3807));
    outputs(5739) <= (layer6_outputs(3543)) and not (layer6_outputs(1484));
    outputs(5740) <= not(layer6_outputs(1727));
    outputs(5741) <= layer6_outputs(1700);
    outputs(5742) <= not(layer6_outputs(873));
    outputs(5743) <= not(layer6_outputs(6178));
    outputs(5744) <= layer6_outputs(2868);
    outputs(5745) <= layer6_outputs(3883);
    outputs(5746) <= not((layer6_outputs(6518)) xor (layer6_outputs(728)));
    outputs(5747) <= not(layer6_outputs(3930));
    outputs(5748) <= (layer6_outputs(6838)) xor (layer6_outputs(4494));
    outputs(5749) <= layer6_outputs(4805);
    outputs(5750) <= not(layer6_outputs(370));
    outputs(5751) <= layer6_outputs(1411);
    outputs(5752) <= not(layer6_outputs(2556));
    outputs(5753) <= not(layer6_outputs(7600)) or (layer6_outputs(6845));
    outputs(5754) <= (layer6_outputs(1508)) and not (layer6_outputs(7103));
    outputs(5755) <= not(layer6_outputs(1267));
    outputs(5756) <= (layer6_outputs(3975)) and (layer6_outputs(6129));
    outputs(5757) <= (layer6_outputs(3997)) and (layer6_outputs(4068));
    outputs(5758) <= not(layer6_outputs(3487));
    outputs(5759) <= not((layer6_outputs(2870)) xor (layer6_outputs(2157)));
    outputs(5760) <= not((layer6_outputs(1942)) xor (layer6_outputs(2025)));
    outputs(5761) <= (layer6_outputs(6237)) and not (layer6_outputs(5481));
    outputs(5762) <= (layer6_outputs(6358)) or (layer6_outputs(5603));
    outputs(5763) <= layer6_outputs(4089);
    outputs(5764) <= not(layer6_outputs(2986));
    outputs(5765) <= layer6_outputs(577);
    outputs(5766) <= layer6_outputs(3858);
    outputs(5767) <= not(layer6_outputs(1963));
    outputs(5768) <= not(layer6_outputs(1517));
    outputs(5769) <= layer6_outputs(1031);
    outputs(5770) <= not(layer6_outputs(4188));
    outputs(5771) <= (layer6_outputs(5778)) xor (layer6_outputs(884));
    outputs(5772) <= layer6_outputs(2183);
    outputs(5773) <= not((layer6_outputs(456)) or (layer6_outputs(6593)));
    outputs(5774) <= not(layer6_outputs(4431));
    outputs(5775) <= layer6_outputs(5295);
    outputs(5776) <= layer6_outputs(2581);
    outputs(5777) <= not((layer6_outputs(388)) xor (layer6_outputs(4617)));
    outputs(5778) <= layer6_outputs(5087);
    outputs(5779) <= layer6_outputs(1769);
    outputs(5780) <= (layer6_outputs(1815)) xor (layer6_outputs(992));
    outputs(5781) <= not(layer6_outputs(7131));
    outputs(5782) <= not((layer6_outputs(4759)) xor (layer6_outputs(4353)));
    outputs(5783) <= (layer6_outputs(3782)) and not (layer6_outputs(1135));
    outputs(5784) <= (layer6_outputs(1494)) or (layer6_outputs(2418));
    outputs(5785) <= layer6_outputs(5796);
    outputs(5786) <= not(layer6_outputs(375));
    outputs(5787) <= not((layer6_outputs(702)) xor (layer6_outputs(3761)));
    outputs(5788) <= not(layer6_outputs(185));
    outputs(5789) <= (layer6_outputs(917)) xor (layer6_outputs(192));
    outputs(5790) <= (layer6_outputs(699)) xor (layer6_outputs(3089));
    outputs(5791) <= layer6_outputs(5700);
    outputs(5792) <= (layer6_outputs(2852)) xor (layer6_outputs(907));
    outputs(5793) <= not(layer6_outputs(6176));
    outputs(5794) <= not(layer6_outputs(7199));
    outputs(5795) <= layer6_outputs(890);
    outputs(5796) <= not((layer6_outputs(6557)) and (layer6_outputs(6791)));
    outputs(5797) <= layer6_outputs(7623);
    outputs(5798) <= not(layer6_outputs(117));
    outputs(5799) <= not(layer6_outputs(393));
    outputs(5800) <= (layer6_outputs(5142)) xor (layer6_outputs(4470));
    outputs(5801) <= layer6_outputs(5916);
    outputs(5802) <= not((layer6_outputs(104)) xor (layer6_outputs(6284)));
    outputs(5803) <= layer6_outputs(7029);
    outputs(5804) <= not((layer6_outputs(5854)) or (layer6_outputs(1177)));
    outputs(5805) <= layer6_outputs(3574);
    outputs(5806) <= layer6_outputs(4189);
    outputs(5807) <= layer6_outputs(3174);
    outputs(5808) <= layer6_outputs(2299);
    outputs(5809) <= not(layer6_outputs(5232));
    outputs(5810) <= layer6_outputs(396);
    outputs(5811) <= (layer6_outputs(3953)) xor (layer6_outputs(2123));
    outputs(5812) <= not(layer6_outputs(3690));
    outputs(5813) <= not((layer6_outputs(4294)) xor (layer6_outputs(5786)));
    outputs(5814) <= layer6_outputs(6069);
    outputs(5815) <= not(layer6_outputs(2936));
    outputs(5816) <= layer6_outputs(6062);
    outputs(5817) <= not(layer6_outputs(5532));
    outputs(5818) <= not((layer6_outputs(6335)) and (layer6_outputs(3242)));
    outputs(5819) <= not(layer6_outputs(2034));
    outputs(5820) <= not(layer6_outputs(1824)) or (layer6_outputs(2898));
    outputs(5821) <= not((layer6_outputs(5580)) xor (layer6_outputs(1691)));
    outputs(5822) <= not(layer6_outputs(3115));
    outputs(5823) <= layer6_outputs(3848);
    outputs(5824) <= layer6_outputs(7446);
    outputs(5825) <= not(layer6_outputs(3821));
    outputs(5826) <= not(layer6_outputs(2964));
    outputs(5827) <= (layer6_outputs(5936)) and not (layer6_outputs(2378));
    outputs(5828) <= not((layer6_outputs(6555)) xor (layer6_outputs(2738)));
    outputs(5829) <= not((layer6_outputs(4561)) xor (layer6_outputs(2392)));
    outputs(5830) <= not((layer6_outputs(4246)) xor (layer6_outputs(7502)));
    outputs(5831) <= not(layer6_outputs(2541));
    outputs(5832) <= (layer6_outputs(6915)) and (layer6_outputs(157));
    outputs(5833) <= not((layer6_outputs(5651)) xor (layer6_outputs(6135)));
    outputs(5834) <= (layer6_outputs(3129)) and not (layer6_outputs(135));
    outputs(5835) <= not(layer6_outputs(3397));
    outputs(5836) <= layer6_outputs(7028);
    outputs(5837) <= (layer6_outputs(258)) and not (layer6_outputs(5454));
    outputs(5838) <= layer6_outputs(1475);
    outputs(5839) <= layer6_outputs(4065);
    outputs(5840) <= (layer6_outputs(1514)) xor (layer6_outputs(229));
    outputs(5841) <= not((layer6_outputs(4798)) xor (layer6_outputs(4440)));
    outputs(5842) <= layer6_outputs(1397);
    outputs(5843) <= not(layer6_outputs(7338));
    outputs(5844) <= not(layer6_outputs(4040));
    outputs(5845) <= layer6_outputs(2805);
    outputs(5846) <= layer6_outputs(4610);
    outputs(5847) <= (layer6_outputs(3969)) xor (layer6_outputs(3220));
    outputs(5848) <= layer6_outputs(6543);
    outputs(5849) <= layer6_outputs(4248);
    outputs(5850) <= not((layer6_outputs(496)) xor (layer6_outputs(1746)));
    outputs(5851) <= (layer6_outputs(4760)) and not (layer6_outputs(4136));
    outputs(5852) <= not(layer6_outputs(6141));
    outputs(5853) <= (layer6_outputs(3221)) xor (layer6_outputs(2390));
    outputs(5854) <= (layer6_outputs(4438)) or (layer6_outputs(7036));
    outputs(5855) <= not(layer6_outputs(2147));
    outputs(5856) <= (layer6_outputs(5377)) and not (layer6_outputs(902));
    outputs(5857) <= not(layer6_outputs(3011));
    outputs(5858) <= not(layer6_outputs(1410));
    outputs(5859) <= not(layer6_outputs(1833)) or (layer6_outputs(6613));
    outputs(5860) <= (layer6_outputs(6267)) and (layer6_outputs(5555));
    outputs(5861) <= not((layer6_outputs(6901)) or (layer6_outputs(6830)));
    outputs(5862) <= layer6_outputs(1670);
    outputs(5863) <= layer6_outputs(5464);
    outputs(5864) <= (layer6_outputs(1779)) xor (layer6_outputs(3606));
    outputs(5865) <= layer6_outputs(3189);
    outputs(5866) <= not(layer6_outputs(5431));
    outputs(5867) <= not(layer6_outputs(193));
    outputs(5868) <= not(layer6_outputs(2140));
    outputs(5869) <= not((layer6_outputs(6310)) or (layer6_outputs(2250)));
    outputs(5870) <= not(layer6_outputs(3995));
    outputs(5871) <= layer6_outputs(7173);
    outputs(5872) <= not((layer6_outputs(202)) xor (layer6_outputs(3457)));
    outputs(5873) <= layer6_outputs(3155);
    outputs(5874) <= not((layer6_outputs(1781)) xor (layer6_outputs(7027)));
    outputs(5875) <= layer6_outputs(5109);
    outputs(5876) <= layer6_outputs(5693);
    outputs(5877) <= layer6_outputs(7076);
    outputs(5878) <= not(layer6_outputs(6624));
    outputs(5879) <= layer6_outputs(7369);
    outputs(5880) <= not(layer6_outputs(487)) or (layer6_outputs(1929));
    outputs(5881) <= not(layer6_outputs(1215));
    outputs(5882) <= not(layer6_outputs(672));
    outputs(5883) <= not((layer6_outputs(4613)) xor (layer6_outputs(3711)));
    outputs(5884) <= layer6_outputs(3976);
    outputs(5885) <= not(layer6_outputs(2158));
    outputs(5886) <= layer6_outputs(1681);
    outputs(5887) <= not((layer6_outputs(4883)) xor (layer6_outputs(6219)));
    outputs(5888) <= layer6_outputs(74);
    outputs(5889) <= layer6_outputs(2616);
    outputs(5890) <= not((layer6_outputs(3888)) xor (layer6_outputs(4566)));
    outputs(5891) <= (layer6_outputs(3294)) xor (layer6_outputs(1054));
    outputs(5892) <= (layer6_outputs(4804)) and (layer6_outputs(4166));
    outputs(5893) <= (layer6_outputs(4966)) and not (layer6_outputs(5115));
    outputs(5894) <= layer6_outputs(4594);
    outputs(5895) <= not((layer6_outputs(435)) xor (layer6_outputs(1256)));
    outputs(5896) <= layer6_outputs(1002);
    outputs(5897) <= (layer6_outputs(1181)) xor (layer6_outputs(3474));
    outputs(5898) <= (layer6_outputs(3160)) xor (layer6_outputs(5661));
    outputs(5899) <= (layer6_outputs(4691)) and not (layer6_outputs(6866));
    outputs(5900) <= not(layer6_outputs(5347));
    outputs(5901) <= layer6_outputs(6799);
    outputs(5902) <= not(layer6_outputs(7270));
    outputs(5903) <= not(layer6_outputs(5340));
    outputs(5904) <= not(layer6_outputs(2298));
    outputs(5905) <= (layer6_outputs(2363)) and (layer6_outputs(35));
    outputs(5906) <= not((layer6_outputs(2639)) xor (layer6_outputs(3394)));
    outputs(5907) <= not(layer6_outputs(2998));
    outputs(5908) <= layer6_outputs(1811);
    outputs(5909) <= (layer6_outputs(6452)) and not (layer6_outputs(251));
    outputs(5910) <= not(layer6_outputs(6590));
    outputs(5911) <= (layer6_outputs(4252)) xor (layer6_outputs(4742));
    outputs(5912) <= layer6_outputs(7040);
    outputs(5913) <= not(layer6_outputs(474));
    outputs(5914) <= (layer6_outputs(3070)) and (layer6_outputs(118));
    outputs(5915) <= (layer6_outputs(5650)) xor (layer6_outputs(6243));
    outputs(5916) <= (layer6_outputs(5260)) and not (layer6_outputs(3885));
    outputs(5917) <= layer6_outputs(4095);
    outputs(5918) <= layer6_outputs(3679);
    outputs(5919) <= layer6_outputs(5958);
    outputs(5920) <= (layer6_outputs(121)) and (layer6_outputs(4586));
    outputs(5921) <= not(layer6_outputs(4620));
    outputs(5922) <= layer6_outputs(1043);
    outputs(5923) <= layer6_outputs(7083);
    outputs(5924) <= not(layer6_outputs(3551));
    outputs(5925) <= not(layer6_outputs(3135));
    outputs(5926) <= (layer6_outputs(7255)) xor (layer6_outputs(793));
    outputs(5927) <= not(layer6_outputs(2941));
    outputs(5928) <= layer6_outputs(3853);
    outputs(5929) <= not(layer6_outputs(4329));
    outputs(5930) <= not(layer6_outputs(5819));
    outputs(5931) <= (layer6_outputs(7032)) xor (layer6_outputs(1141));
    outputs(5932) <= not(layer6_outputs(4127));
    outputs(5933) <= not(layer6_outputs(1416));
    outputs(5934) <= layer6_outputs(2339);
    outputs(5935) <= not((layer6_outputs(5029)) or (layer6_outputs(5793)));
    outputs(5936) <= (layer6_outputs(4732)) and (layer6_outputs(2847));
    outputs(5937) <= not(layer6_outputs(1951));
    outputs(5938) <= not((layer6_outputs(6498)) xor (layer6_outputs(1457)));
    outputs(5939) <= not((layer6_outputs(1742)) xor (layer6_outputs(2180)));
    outputs(5940) <= layer6_outputs(1840);
    outputs(5941) <= not(layer6_outputs(1060));
    outputs(5942) <= not((layer6_outputs(3201)) xor (layer6_outputs(3342)));
    outputs(5943) <= not(layer6_outputs(630));
    outputs(5944) <= not(layer6_outputs(6505));
    outputs(5945) <= (layer6_outputs(2228)) xor (layer6_outputs(7579));
    outputs(5946) <= layer6_outputs(458);
    outputs(5947) <= not(layer6_outputs(1268)) or (layer6_outputs(309));
    outputs(5948) <= (layer6_outputs(2662)) xor (layer6_outputs(2016));
    outputs(5949) <= (layer6_outputs(3179)) and not (layer6_outputs(1211));
    outputs(5950) <= not(layer6_outputs(2680));
    outputs(5951) <= not(layer6_outputs(5539));
    outputs(5952) <= not(layer6_outputs(347));
    outputs(5953) <= not(layer6_outputs(3454));
    outputs(5954) <= not((layer6_outputs(3344)) xor (layer6_outputs(5673)));
    outputs(5955) <= not(layer6_outputs(756));
    outputs(5956) <= layer6_outputs(2453);
    outputs(5957) <= layer6_outputs(2341);
    outputs(5958) <= layer6_outputs(2809);
    outputs(5959) <= layer6_outputs(3963);
    outputs(5960) <= (layer6_outputs(1156)) xor (layer6_outputs(5920));
    outputs(5961) <= (layer6_outputs(1678)) xor (layer6_outputs(6993));
    outputs(5962) <= not(layer6_outputs(2660));
    outputs(5963) <= (layer6_outputs(5141)) xor (layer6_outputs(346));
    outputs(5964) <= layer6_outputs(5492);
    outputs(5965) <= not(layer6_outputs(5945));
    outputs(5966) <= layer6_outputs(6181);
    outputs(5967) <= not(layer6_outputs(4834));
    outputs(5968) <= not(layer6_outputs(2450));
    outputs(5969) <= not(layer6_outputs(1783));
    outputs(5970) <= layer6_outputs(4898);
    outputs(5971) <= layer6_outputs(5268);
    outputs(5972) <= not(layer6_outputs(2391));
    outputs(5973) <= not((layer6_outputs(3414)) xor (layer6_outputs(4017)));
    outputs(5974) <= not(layer6_outputs(4548)) or (layer6_outputs(3584));
    outputs(5975) <= not((layer6_outputs(1159)) xor (layer6_outputs(7492)));
    outputs(5976) <= layer6_outputs(7168);
    outputs(5977) <= (layer6_outputs(4791)) and not (layer6_outputs(109));
    outputs(5978) <= (layer6_outputs(2774)) xor (layer6_outputs(1045));
    outputs(5979) <= (layer6_outputs(2357)) and not (layer6_outputs(109));
    outputs(5980) <= not((layer6_outputs(7256)) xor (layer6_outputs(3845)));
    outputs(5981) <= layer6_outputs(4511);
    outputs(5982) <= layer6_outputs(837);
    outputs(5983) <= not((layer6_outputs(7219)) xor (layer6_outputs(4924)));
    outputs(5984) <= not(layer6_outputs(1659));
    outputs(5985) <= (layer6_outputs(3107)) xor (layer6_outputs(6511));
    outputs(5986) <= not(layer6_outputs(4509));
    outputs(5987) <= not(layer6_outputs(6868));
    outputs(5988) <= (layer6_outputs(31)) xor (layer6_outputs(386));
    outputs(5989) <= layer6_outputs(2930);
    outputs(5990) <= not((layer6_outputs(5837)) xor (layer6_outputs(2839)));
    outputs(5991) <= layer6_outputs(3846);
    outputs(5992) <= not(layer6_outputs(5003));
    outputs(5993) <= layer6_outputs(2621);
    outputs(5994) <= layer6_outputs(3982);
    outputs(5995) <= layer6_outputs(6723);
    outputs(5996) <= (layer6_outputs(5091)) xor (layer6_outputs(6712));
    outputs(5997) <= (layer6_outputs(5840)) and (layer6_outputs(7059));
    outputs(5998) <= not((layer6_outputs(6801)) or (layer6_outputs(6252)));
    outputs(5999) <= layer6_outputs(3603);
    outputs(6000) <= (layer6_outputs(4467)) xor (layer6_outputs(664));
    outputs(6001) <= (layer6_outputs(1592)) or (layer6_outputs(56));
    outputs(6002) <= not((layer6_outputs(2147)) or (layer6_outputs(4113)));
    outputs(6003) <= not(layer6_outputs(6602));
    outputs(6004) <= layer6_outputs(2068);
    outputs(6005) <= not((layer6_outputs(2091)) xor (layer6_outputs(3792)));
    outputs(6006) <= not(layer6_outputs(7003));
    outputs(6007) <= (layer6_outputs(6595)) and not (layer6_outputs(3665));
    outputs(6008) <= layer6_outputs(2524);
    outputs(6009) <= not(layer6_outputs(5596));
    outputs(6010) <= not(layer6_outputs(1188));
    outputs(6011) <= (layer6_outputs(1000)) and not (layer6_outputs(3916));
    outputs(6012) <= layer6_outputs(7080);
    outputs(6013) <= not((layer6_outputs(4272)) xor (layer6_outputs(4598)));
    outputs(6014) <= (layer6_outputs(5399)) xor (layer6_outputs(5176));
    outputs(6015) <= layer6_outputs(422);
    outputs(6016) <= (layer6_outputs(1943)) and (layer6_outputs(6356));
    outputs(6017) <= layer6_outputs(5274);
    outputs(6018) <= layer6_outputs(1981);
    outputs(6019) <= not(layer6_outputs(4174)) or (layer6_outputs(3611));
    outputs(6020) <= not((layer6_outputs(680)) xor (layer6_outputs(6225)));
    outputs(6021) <= layer6_outputs(1492);
    outputs(6022) <= (layer6_outputs(16)) xor (layer6_outputs(6801));
    outputs(6023) <= not(layer6_outputs(2950)) or (layer6_outputs(7510));
    outputs(6024) <= not((layer6_outputs(3281)) xor (layer6_outputs(4839)));
    outputs(6025) <= not(layer6_outputs(3512)) or (layer6_outputs(4868));
    outputs(6026) <= layer6_outputs(5395);
    outputs(6027) <= (layer6_outputs(5627)) xor (layer6_outputs(654));
    outputs(6028) <= (layer6_outputs(7466)) xor (layer6_outputs(3833));
    outputs(6029) <= (layer6_outputs(7635)) and not (layer6_outputs(3197));
    outputs(6030) <= not(layer6_outputs(1125));
    outputs(6031) <= not(layer6_outputs(6722));
    outputs(6032) <= (layer6_outputs(7005)) xor (layer6_outputs(5808));
    outputs(6033) <= (layer6_outputs(5767)) and (layer6_outputs(7473));
    outputs(6034) <= (layer6_outputs(4084)) xor (layer6_outputs(7316));
    outputs(6035) <= not(layer6_outputs(1934));
    outputs(6036) <= not((layer6_outputs(4508)) xor (layer6_outputs(830)));
    outputs(6037) <= layer6_outputs(538);
    outputs(6038) <= (layer6_outputs(4032)) xor (layer6_outputs(5266));
    outputs(6039) <= (layer6_outputs(7430)) and (layer6_outputs(4008));
    outputs(6040) <= (layer6_outputs(3007)) and (layer6_outputs(2335));
    outputs(6041) <= not(layer6_outputs(2052));
    outputs(6042) <= not((layer6_outputs(1597)) and (layer6_outputs(5231)));
    outputs(6043) <= (layer6_outputs(745)) and not (layer6_outputs(1446));
    outputs(6044) <= layer6_outputs(1325);
    outputs(6045) <= (layer6_outputs(905)) and not (layer6_outputs(5950));
    outputs(6046) <= layer6_outputs(4189);
    outputs(6047) <= layer6_outputs(1849);
    outputs(6048) <= not(layer6_outputs(4707));
    outputs(6049) <= layer6_outputs(527);
    outputs(6050) <= layer6_outputs(6408);
    outputs(6051) <= layer6_outputs(121);
    outputs(6052) <= not((layer6_outputs(3334)) xor (layer6_outputs(1779)));
    outputs(6053) <= not(layer6_outputs(1406));
    outputs(6054) <= (layer6_outputs(3396)) xor (layer6_outputs(1723));
    outputs(6055) <= not((layer6_outputs(1970)) xor (layer6_outputs(3215)));
    outputs(6056) <= (layer6_outputs(3277)) xor (layer6_outputs(4937));
    outputs(6057) <= (layer6_outputs(2332)) xor (layer6_outputs(6617));
    outputs(6058) <= layer6_outputs(833);
    outputs(6059) <= not(layer6_outputs(2447));
    outputs(6060) <= layer6_outputs(7183);
    outputs(6061) <= (layer6_outputs(1898)) xor (layer6_outputs(371));
    outputs(6062) <= not((layer6_outputs(4410)) xor (layer6_outputs(3746)));
    outputs(6063) <= (layer6_outputs(3623)) xor (layer6_outputs(433));
    outputs(6064) <= not(layer6_outputs(1153));
    outputs(6065) <= not(layer6_outputs(6923));
    outputs(6066) <= not(layer6_outputs(2426));
    outputs(6067) <= layer6_outputs(3217);
    outputs(6068) <= (layer6_outputs(3758)) xor (layer6_outputs(5831));
    outputs(6069) <= not(layer6_outputs(6067));
    outputs(6070) <= (layer6_outputs(6026)) and (layer6_outputs(422));
    outputs(6071) <= layer6_outputs(4783);
    outputs(6072) <= layer6_outputs(2911);
    outputs(6073) <= layer6_outputs(3580);
    outputs(6074) <= not(layer6_outputs(7202));
    outputs(6075) <= not((layer6_outputs(2530)) or (layer6_outputs(4155)));
    outputs(6076) <= not(layer6_outputs(89));
    outputs(6077) <= (layer6_outputs(6471)) and not (layer6_outputs(4961));
    outputs(6078) <= not(layer6_outputs(1735));
    outputs(6079) <= not(layer6_outputs(13));
    outputs(6080) <= layer6_outputs(2698);
    outputs(6081) <= not((layer6_outputs(6787)) or (layer6_outputs(4312)));
    outputs(6082) <= not(layer6_outputs(5874));
    outputs(6083) <= (layer6_outputs(1655)) and not (layer6_outputs(2307));
    outputs(6084) <= not(layer6_outputs(1788));
    outputs(6085) <= layer6_outputs(5717);
    outputs(6086) <= not(layer6_outputs(6880));
    outputs(6087) <= layer6_outputs(3986);
    outputs(6088) <= layer6_outputs(407);
    outputs(6089) <= not(layer6_outputs(2274));
    outputs(6090) <= (layer6_outputs(7069)) and not (layer6_outputs(3443));
    outputs(6091) <= layer6_outputs(7109);
    outputs(6092) <= layer6_outputs(3599);
    outputs(6093) <= not(layer6_outputs(2764));
    outputs(6094) <= (layer6_outputs(3550)) and not (layer6_outputs(1615));
    outputs(6095) <= not((layer6_outputs(2676)) or (layer6_outputs(665)));
    outputs(6096) <= not(layer6_outputs(4124));
    outputs(6097) <= layer6_outputs(390);
    outputs(6098) <= not(layer6_outputs(4345));
    outputs(6099) <= layer6_outputs(96);
    outputs(6100) <= not(layer6_outputs(4456));
    outputs(6101) <= layer6_outputs(7017);
    outputs(6102) <= layer6_outputs(3782);
    outputs(6103) <= not((layer6_outputs(6662)) xor (layer6_outputs(5937)));
    outputs(6104) <= not(layer6_outputs(6308));
    outputs(6105) <= layer6_outputs(5821);
    outputs(6106) <= (layer6_outputs(6125)) and not (layer6_outputs(4107));
    outputs(6107) <= layer6_outputs(6223);
    outputs(6108) <= (layer6_outputs(1892)) xor (layer6_outputs(1601));
    outputs(6109) <= not(layer6_outputs(5366));
    outputs(6110) <= (layer6_outputs(3832)) and not (layer6_outputs(274));
    outputs(6111) <= not(layer6_outputs(5004));
    outputs(6112) <= not((layer6_outputs(352)) xor (layer6_outputs(1661)));
    outputs(6113) <= layer6_outputs(7122);
    outputs(6114) <= not(layer6_outputs(3370));
    outputs(6115) <= layer6_outputs(3693);
    outputs(6116) <= not(layer6_outputs(1286));
    outputs(6117) <= not(layer6_outputs(2770));
    outputs(6118) <= not((layer6_outputs(5909)) xor (layer6_outputs(5294)));
    outputs(6119) <= not(layer6_outputs(609));
    outputs(6120) <= (layer6_outputs(621)) xor (layer6_outputs(2668));
    outputs(6121) <= not(layer6_outputs(6607));
    outputs(6122) <= not((layer6_outputs(6332)) xor (layer6_outputs(7606)));
    outputs(6123) <= layer6_outputs(2334);
    outputs(6124) <= not(layer6_outputs(6139));
    outputs(6125) <= (layer6_outputs(6540)) xor (layer6_outputs(1315));
    outputs(6126) <= not(layer6_outputs(967));
    outputs(6127) <= not(layer6_outputs(891));
    outputs(6128) <= not((layer6_outputs(3977)) and (layer6_outputs(5525)));
    outputs(6129) <= layer6_outputs(4997);
    outputs(6130) <= (layer6_outputs(4947)) xor (layer6_outputs(7334));
    outputs(6131) <= (layer6_outputs(1361)) xor (layer6_outputs(4309));
    outputs(6132) <= not(layer6_outputs(4521));
    outputs(6133) <= not(layer6_outputs(543));
    outputs(6134) <= layer6_outputs(6120);
    outputs(6135) <= not(layer6_outputs(5972));
    outputs(6136) <= (layer6_outputs(1649)) xor (layer6_outputs(3485));
    outputs(6137) <= layer6_outputs(1330);
    outputs(6138) <= not(layer6_outputs(3484));
    outputs(6139) <= (layer6_outputs(4254)) xor (layer6_outputs(378));
    outputs(6140) <= layer6_outputs(4331);
    outputs(6141) <= not((layer6_outputs(4490)) or (layer6_outputs(3746)));
    outputs(6142) <= not(layer6_outputs(76));
    outputs(6143) <= not((layer6_outputs(657)) xor (layer6_outputs(5821)));
    outputs(6144) <= (layer6_outputs(974)) xor (layer6_outputs(7170));
    outputs(6145) <= not((layer6_outputs(3119)) and (layer6_outputs(1198)));
    outputs(6146) <= layer6_outputs(3400);
    outputs(6147) <= (layer6_outputs(4802)) xor (layer6_outputs(493));
    outputs(6148) <= (layer6_outputs(4208)) xor (layer6_outputs(4497));
    outputs(6149) <= not((layer6_outputs(3447)) xor (layer6_outputs(5365)));
    outputs(6150) <= (layer6_outputs(6507)) and not (layer6_outputs(836));
    outputs(6151) <= not(layer6_outputs(377));
    outputs(6152) <= not((layer6_outputs(4242)) xor (layer6_outputs(6846)));
    outputs(6153) <= (layer6_outputs(2430)) xor (layer6_outputs(2231));
    outputs(6154) <= not(layer6_outputs(4769)) or (layer6_outputs(1167));
    outputs(6155) <= layer6_outputs(2016);
    outputs(6156) <= (layer6_outputs(1916)) and (layer6_outputs(4562));
    outputs(6157) <= not(layer6_outputs(4790));
    outputs(6158) <= not(layer6_outputs(4452));
    outputs(6159) <= layer6_outputs(3224);
    outputs(6160) <= not(layer6_outputs(4840)) or (layer6_outputs(2024));
    outputs(6161) <= (layer6_outputs(3838)) xor (layer6_outputs(1255));
    outputs(6162) <= not((layer6_outputs(1439)) xor (layer6_outputs(3397)));
    outputs(6163) <= not(layer6_outputs(7151)) or (layer6_outputs(1723));
    outputs(6164) <= not(layer6_outputs(329));
    outputs(6165) <= not(layer6_outputs(1603));
    outputs(6166) <= layer6_outputs(2474);
    outputs(6167) <= (layer6_outputs(580)) xor (layer6_outputs(981));
    outputs(6168) <= (layer6_outputs(7068)) and not (layer6_outputs(6379));
    outputs(6169) <= (layer6_outputs(4709)) xor (layer6_outputs(2073));
    outputs(6170) <= layer6_outputs(6207);
    outputs(6171) <= not((layer6_outputs(7644)) xor (layer6_outputs(1236)));
    outputs(6172) <= (layer6_outputs(6599)) xor (layer6_outputs(911));
    outputs(6173) <= not((layer6_outputs(5306)) xor (layer6_outputs(3438)));
    outputs(6174) <= not(layer6_outputs(4996));
    outputs(6175) <= (layer6_outputs(2864)) xor (layer6_outputs(5050));
    outputs(6176) <= layer6_outputs(6095);
    outputs(6177) <= not((layer6_outputs(1930)) xor (layer6_outputs(2741)));
    outputs(6178) <= not((layer6_outputs(4900)) xor (layer6_outputs(1132)));
    outputs(6179) <= layer6_outputs(2904);
    outputs(6180) <= not(layer6_outputs(1893));
    outputs(6181) <= layer6_outputs(5930);
    outputs(6182) <= (layer6_outputs(2782)) xor (layer6_outputs(7214));
    outputs(6183) <= not(layer6_outputs(4787));
    outputs(6184) <= layer6_outputs(4538);
    outputs(6185) <= not(layer6_outputs(3134));
    outputs(6186) <= not((layer6_outputs(144)) xor (layer6_outputs(1944)));
    outputs(6187) <= not(layer6_outputs(1885)) or (layer6_outputs(7397));
    outputs(6188) <= (layer6_outputs(700)) xor (layer6_outputs(4048));
    outputs(6189) <= not(layer6_outputs(4674));
    outputs(6190) <= not((layer6_outputs(5516)) xor (layer6_outputs(2524)));
    outputs(6191) <= not((layer6_outputs(1883)) or (layer6_outputs(1953)));
    outputs(6192) <= (layer6_outputs(5102)) and (layer6_outputs(483));
    outputs(6193) <= not((layer6_outputs(2825)) or (layer6_outputs(1780)));
    outputs(6194) <= not(layer6_outputs(909));
    outputs(6195) <= not(layer6_outputs(292));
    outputs(6196) <= (layer6_outputs(7272)) xor (layer6_outputs(92));
    outputs(6197) <= layer6_outputs(5434);
    outputs(6198) <= not(layer6_outputs(1247)) or (layer6_outputs(2696));
    outputs(6199) <= layer6_outputs(5098);
    outputs(6200) <= not(layer6_outputs(1214));
    outputs(6201) <= layer6_outputs(6743);
    outputs(6202) <= (layer6_outputs(4045)) xor (layer6_outputs(5971));
    outputs(6203) <= not(layer6_outputs(1919));
    outputs(6204) <= not(layer6_outputs(1769)) or (layer6_outputs(447));
    outputs(6205) <= (layer6_outputs(2902)) and (layer6_outputs(6132));
    outputs(6206) <= layer6_outputs(5279);
    outputs(6207) <= layer6_outputs(840);
    outputs(6208) <= layer6_outputs(7010);
    outputs(6209) <= '1';
    outputs(6210) <= layer6_outputs(5247);
    outputs(6211) <= not((layer6_outputs(1559)) xor (layer6_outputs(138)));
    outputs(6212) <= not(layer6_outputs(5852)) or (layer6_outputs(1900));
    outputs(6213) <= layer6_outputs(4241);
    outputs(6214) <= (layer6_outputs(4611)) xor (layer6_outputs(6162));
    outputs(6215) <= layer6_outputs(956);
    outputs(6216) <= not(layer6_outputs(3823));
    outputs(6217) <= not(layer6_outputs(7650));
    outputs(6218) <= layer6_outputs(5813);
    outputs(6219) <= not((layer6_outputs(6657)) xor (layer6_outputs(3612)));
    outputs(6220) <= not((layer6_outputs(1786)) xor (layer6_outputs(1505)));
    outputs(6221) <= layer6_outputs(33);
    outputs(6222) <= not(layer6_outputs(668));
    outputs(6223) <= layer6_outputs(4004);
    outputs(6224) <= not((layer6_outputs(3385)) xor (layer6_outputs(7668)));
    outputs(6225) <= not(layer6_outputs(5882)) or (layer6_outputs(1399));
    outputs(6226) <= layer6_outputs(5083);
    outputs(6227) <= (layer6_outputs(7078)) xor (layer6_outputs(3744));
    outputs(6228) <= not((layer6_outputs(449)) and (layer6_outputs(5414)));
    outputs(6229) <= not((layer6_outputs(165)) xor (layer6_outputs(2430)));
    outputs(6230) <= (layer6_outputs(3231)) xor (layer6_outputs(3413));
    outputs(6231) <= not((layer6_outputs(633)) xor (layer6_outputs(5864)));
    outputs(6232) <= (layer6_outputs(7665)) or (layer6_outputs(5684));
    outputs(6233) <= (layer6_outputs(4480)) xor (layer6_outputs(4024));
    outputs(6234) <= not(layer6_outputs(4468));
    outputs(6235) <= not((layer6_outputs(250)) xor (layer6_outputs(2741)));
    outputs(6236) <= layer6_outputs(4278);
    outputs(6237) <= not(layer6_outputs(1075));
    outputs(6238) <= layer6_outputs(2545);
    outputs(6239) <= not((layer6_outputs(556)) xor (layer6_outputs(5133)));
    outputs(6240) <= not(layer6_outputs(5624));
    outputs(6241) <= layer6_outputs(5582);
    outputs(6242) <= not(layer6_outputs(2266));
    outputs(6243) <= layer6_outputs(3362);
    outputs(6244) <= not(layer6_outputs(2107));
    outputs(6245) <= not(layer6_outputs(1863));
    outputs(6246) <= layer6_outputs(6214);
    outputs(6247) <= not(layer6_outputs(7182));
    outputs(6248) <= not(layer6_outputs(7045));
    outputs(6249) <= not(layer6_outputs(5166));
    outputs(6250) <= not(layer6_outputs(2361));
    outputs(6251) <= layer6_outputs(6303);
    outputs(6252) <= layer6_outputs(3346);
    outputs(6253) <= layer6_outputs(1816);
    outputs(6254) <= not(layer6_outputs(1871)) or (layer6_outputs(5932));
    outputs(6255) <= not(layer6_outputs(4898)) or (layer6_outputs(1952));
    outputs(6256) <= not((layer6_outputs(7180)) and (layer6_outputs(6038)));
    outputs(6257) <= (layer6_outputs(6903)) xor (layer6_outputs(4203));
    outputs(6258) <= layer6_outputs(32);
    outputs(6259) <= not(layer6_outputs(1932));
    outputs(6260) <= layer6_outputs(7001);
    outputs(6261) <= not(layer6_outputs(1922)) or (layer6_outputs(3900));
    outputs(6262) <= layer6_outputs(4971);
    outputs(6263) <= not(layer6_outputs(246));
    outputs(6264) <= not(layer6_outputs(4861));
    outputs(6265) <= (layer6_outputs(1217)) or (layer6_outputs(5314));
    outputs(6266) <= not((layer6_outputs(3514)) xor (layer6_outputs(4918)));
    outputs(6267) <= (layer6_outputs(1740)) xor (layer6_outputs(6484));
    outputs(6268) <= (layer6_outputs(1728)) or (layer6_outputs(1103));
    outputs(6269) <= not(layer6_outputs(385));
    outputs(6270) <= (layer6_outputs(4451)) xor (layer6_outputs(4793));
    outputs(6271) <= layer6_outputs(5223);
    outputs(6272) <= layer6_outputs(6752);
    outputs(6273) <= not(layer6_outputs(6497));
    outputs(6274) <= (layer6_outputs(7177)) and (layer6_outputs(1310));
    outputs(6275) <= not(layer6_outputs(3128)) or (layer6_outputs(3681));
    outputs(6276) <= (layer6_outputs(6741)) xor (layer6_outputs(3061));
    outputs(6277) <= not(layer6_outputs(156)) or (layer6_outputs(356));
    outputs(6278) <= not(layer6_outputs(3806));
    outputs(6279) <= not(layer6_outputs(4356));
    outputs(6280) <= layer6_outputs(3799);
    outputs(6281) <= layer6_outputs(3056);
    outputs(6282) <= not(layer6_outputs(6474)) or (layer6_outputs(6168));
    outputs(6283) <= layer6_outputs(4629);
    outputs(6284) <= not((layer6_outputs(388)) xor (layer6_outputs(2535)));
    outputs(6285) <= not(layer6_outputs(1322)) or (layer6_outputs(6550));
    outputs(6286) <= (layer6_outputs(1095)) xor (layer6_outputs(6962));
    outputs(6287) <= layer6_outputs(5619);
    outputs(6288) <= not((layer6_outputs(3732)) xor (layer6_outputs(4051)));
    outputs(6289) <= not(layer6_outputs(5529));
    outputs(6290) <= not((layer6_outputs(6180)) xor (layer6_outputs(2251)));
    outputs(6291) <= (layer6_outputs(5822)) xor (layer6_outputs(5225));
    outputs(6292) <= (layer6_outputs(3338)) xor (layer6_outputs(32));
    outputs(6293) <= layer6_outputs(5421);
    outputs(6294) <= not(layer6_outputs(426));
    outputs(6295) <= layer6_outputs(703);
    outputs(6296) <= layer6_outputs(938);
    outputs(6297) <= not(layer6_outputs(6782)) or (layer6_outputs(3588));
    outputs(6298) <= not((layer6_outputs(800)) xor (layer6_outputs(4698)));
    outputs(6299) <= layer6_outputs(3272);
    outputs(6300) <= not(layer6_outputs(2188));
    outputs(6301) <= not((layer6_outputs(5730)) and (layer6_outputs(4481)));
    outputs(6302) <= not((layer6_outputs(712)) and (layer6_outputs(7039)));
    outputs(6303) <= not((layer6_outputs(5596)) xor (layer6_outputs(2418)));
    outputs(6304) <= (layer6_outputs(6097)) xor (layer6_outputs(3462));
    outputs(6305) <= not((layer6_outputs(567)) xor (layer6_outputs(7378)));
    outputs(6306) <= layer6_outputs(2505);
    outputs(6307) <= not(layer6_outputs(6227));
    outputs(6308) <= not(layer6_outputs(933));
    outputs(6309) <= not(layer6_outputs(1100));
    outputs(6310) <= not((layer6_outputs(1204)) xor (layer6_outputs(4440)));
    outputs(6311) <= layer6_outputs(5184);
    outputs(6312) <= not(layer6_outputs(6353));
    outputs(6313) <= not(layer6_outputs(1277));
    outputs(6314) <= not(layer6_outputs(5214));
    outputs(6315) <= (layer6_outputs(7088)) and not (layer6_outputs(5413));
    outputs(6316) <= not(layer6_outputs(5470));
    outputs(6317) <= layer6_outputs(2404);
    outputs(6318) <= not(layer6_outputs(7634));
    outputs(6319) <= not(layer6_outputs(1015)) or (layer6_outputs(6149));
    outputs(6320) <= layer6_outputs(4962);
    outputs(6321) <= layer6_outputs(3172);
    outputs(6322) <= (layer6_outputs(1363)) xor (layer6_outputs(3067));
    outputs(6323) <= layer6_outputs(2217);
    outputs(6324) <= not(layer6_outputs(6922));
    outputs(6325) <= layer6_outputs(2019);
    outputs(6326) <= layer6_outputs(1456);
    outputs(6327) <= layer6_outputs(3595);
    outputs(6328) <= not(layer6_outputs(211));
    outputs(6329) <= layer6_outputs(3091);
    outputs(6330) <= not(layer6_outputs(4882));
    outputs(6331) <= not(layer6_outputs(7408));
    outputs(6332) <= not(layer6_outputs(1240));
    outputs(6333) <= not(layer6_outputs(2125));
    outputs(6334) <= layer6_outputs(5132);
    outputs(6335) <= not(layer6_outputs(607)) or (layer6_outputs(5062));
    outputs(6336) <= layer6_outputs(2549);
    outputs(6337) <= not(layer6_outputs(6442));
    outputs(6338) <= (layer6_outputs(5709)) and (layer6_outputs(6419));
    outputs(6339) <= (layer6_outputs(5440)) xor (layer6_outputs(4121));
    outputs(6340) <= layer6_outputs(4077);
    outputs(6341) <= not((layer6_outputs(6654)) xor (layer6_outputs(6772)));
    outputs(6342) <= not((layer6_outputs(3808)) xor (layer6_outputs(1126)));
    outputs(6343) <= layer6_outputs(3864);
    outputs(6344) <= not((layer6_outputs(1255)) xor (layer6_outputs(4479)));
    outputs(6345) <= layer6_outputs(9);
    outputs(6346) <= layer6_outputs(1966);
    outputs(6347) <= (layer6_outputs(1300)) xor (layer6_outputs(2611));
    outputs(6348) <= not(layer6_outputs(6011));
    outputs(6349) <= (layer6_outputs(478)) xor (layer6_outputs(3744));
    outputs(6350) <= not((layer6_outputs(4914)) xor (layer6_outputs(1270)));
    outputs(6351) <= not((layer6_outputs(3834)) xor (layer6_outputs(2528)));
    outputs(6352) <= not(layer6_outputs(4238));
    outputs(6353) <= not(layer6_outputs(6804));
    outputs(6354) <= (layer6_outputs(3406)) xor (layer6_outputs(2646));
    outputs(6355) <= not(layer6_outputs(6867));
    outputs(6356) <= not((layer6_outputs(403)) xor (layer6_outputs(5227)));
    outputs(6357) <= not(layer6_outputs(1846));
    outputs(6358) <= not((layer6_outputs(867)) xor (layer6_outputs(6708)));
    outputs(6359) <= not((layer6_outputs(4564)) and (layer6_outputs(1969)));
    outputs(6360) <= (layer6_outputs(6675)) xor (layer6_outputs(7369));
    outputs(6361) <= layer6_outputs(6508);
    outputs(6362) <= layer6_outputs(3715);
    outputs(6363) <= not(layer6_outputs(6810));
    outputs(6364) <= not(layer6_outputs(5440));
    outputs(6365) <= layer6_outputs(2726);
    outputs(6366) <= (layer6_outputs(1339)) xor (layer6_outputs(257));
    outputs(6367) <= not(layer6_outputs(3769));
    outputs(6368) <= layer6_outputs(6345);
    outputs(6369) <= not((layer6_outputs(5865)) xor (layer6_outputs(3994)));
    outputs(6370) <= (layer6_outputs(4255)) or (layer6_outputs(6790));
    outputs(6371) <= not(layer6_outputs(145));
    outputs(6372) <= not(layer6_outputs(682));
    outputs(6373) <= layer6_outputs(3923);
    outputs(6374) <= not((layer6_outputs(3488)) xor (layer6_outputs(4144)));
    outputs(6375) <= not(layer6_outputs(4766));
    outputs(6376) <= not(layer6_outputs(4693));
    outputs(6377) <= layer6_outputs(3523);
    outputs(6378) <= not(layer6_outputs(4654)) or (layer6_outputs(1882));
    outputs(6379) <= (layer6_outputs(5756)) xor (layer6_outputs(5014));
    outputs(6380) <= not(layer6_outputs(7137)) or (layer6_outputs(6461));
    outputs(6381) <= (layer6_outputs(3056)) and (layer6_outputs(7046));
    outputs(6382) <= (layer6_outputs(742)) xor (layer6_outputs(6680));
    outputs(6383) <= not(layer6_outputs(5513));
    outputs(6384) <= not(layer6_outputs(5278));
    outputs(6385) <= (layer6_outputs(6482)) xor (layer6_outputs(195));
    outputs(6386) <= (layer6_outputs(3145)) xor (layer6_outputs(7110));
    outputs(6387) <= not(layer6_outputs(2160));
    outputs(6388) <= (layer6_outputs(5714)) xor (layer6_outputs(4802));
    outputs(6389) <= layer6_outputs(3523);
    outputs(6390) <= not(layer6_outputs(2054)) or (layer6_outputs(1518));
    outputs(6391) <= layer6_outputs(2536);
    outputs(6392) <= (layer6_outputs(5851)) xor (layer6_outputs(6811));
    outputs(6393) <= (layer6_outputs(1552)) xor (layer6_outputs(629));
    outputs(6394) <= not(layer6_outputs(5108));
    outputs(6395) <= (layer6_outputs(1262)) xor (layer6_outputs(4348));
    outputs(6396) <= not(layer6_outputs(317));
    outputs(6397) <= not((layer6_outputs(2114)) xor (layer6_outputs(3064)));
    outputs(6398) <= not(layer6_outputs(7011));
    outputs(6399) <= (layer6_outputs(5163)) xor (layer6_outputs(3822));
    outputs(6400) <= layer6_outputs(443);
    outputs(6401) <= (layer6_outputs(4976)) or (layer6_outputs(5696));
    outputs(6402) <= not(layer6_outputs(613));
    outputs(6403) <= (layer6_outputs(5822)) xor (layer6_outputs(1926));
    outputs(6404) <= not(layer6_outputs(7265));
    outputs(6405) <= not(layer6_outputs(2636)) or (layer6_outputs(3826));
    outputs(6406) <= not(layer6_outputs(3993));
    outputs(6407) <= layer6_outputs(251);
    outputs(6408) <= not(layer6_outputs(3593));
    outputs(6409) <= not(layer6_outputs(3378));
    outputs(6410) <= not(layer6_outputs(3240));
    outputs(6411) <= (layer6_outputs(569)) xor (layer6_outputs(367));
    outputs(6412) <= not(layer6_outputs(6584)) or (layer6_outputs(550));
    outputs(6413) <= layer6_outputs(2263);
    outputs(6414) <= not(layer6_outputs(2992));
    outputs(6415) <= not((layer6_outputs(6963)) xor (layer6_outputs(7388)));
    outputs(6416) <= layer6_outputs(5996);
    outputs(6417) <= not((layer6_outputs(6165)) xor (layer6_outputs(4424)));
    outputs(6418) <= layer6_outputs(4865);
    outputs(6419) <= (layer6_outputs(6213)) xor (layer6_outputs(3456));
    outputs(6420) <= not(layer6_outputs(5926));
    outputs(6421) <= not((layer6_outputs(1445)) xor (layer6_outputs(6559)));
    outputs(6422) <= layer6_outputs(4198);
    outputs(6423) <= layer6_outputs(4433);
    outputs(6424) <= layer6_outputs(3592);
    outputs(6425) <= layer6_outputs(7070);
    outputs(6426) <= layer6_outputs(7204);
    outputs(6427) <= (layer6_outputs(7470)) xor (layer6_outputs(4527));
    outputs(6428) <= not(layer6_outputs(4903));
    outputs(6429) <= (layer6_outputs(7345)) xor (layer6_outputs(1985));
    outputs(6430) <= layer6_outputs(5005);
    outputs(6431) <= (layer6_outputs(481)) or (layer6_outputs(5347));
    outputs(6432) <= layer6_outputs(3699);
    outputs(6433) <= not(layer6_outputs(98));
    outputs(6434) <= not((layer6_outputs(4426)) xor (layer6_outputs(7385)));
    outputs(6435) <= not(layer6_outputs(6735));
    outputs(6436) <= layer6_outputs(6090);
    outputs(6437) <= layer6_outputs(3471);
    outputs(6438) <= not(layer6_outputs(256));
    outputs(6439) <= layer6_outputs(120);
    outputs(6440) <= (layer6_outputs(3385)) xor (layer6_outputs(4402));
    outputs(6441) <= layer6_outputs(7191);
    outputs(6442) <= not(layer6_outputs(1170));
    outputs(6443) <= (layer6_outputs(1516)) xor (layer6_outputs(845));
    outputs(6444) <= (layer6_outputs(7576)) xor (layer6_outputs(4504));
    outputs(6445) <= (layer6_outputs(1745)) xor (layer6_outputs(5451));
    outputs(6446) <= not(layer6_outputs(6347));
    outputs(6447) <= layer6_outputs(7517);
    outputs(6448) <= (layer6_outputs(5437)) xor (layer6_outputs(304));
    outputs(6449) <= not((layer6_outputs(1593)) xor (layer6_outputs(2137)));
    outputs(6450) <= not((layer6_outputs(7182)) and (layer6_outputs(4772)));
    outputs(6451) <= (layer6_outputs(3099)) xor (layer6_outputs(4405));
    outputs(6452) <= (layer6_outputs(2578)) xor (layer6_outputs(2118));
    outputs(6453) <= not((layer6_outputs(3552)) xor (layer6_outputs(7053)));
    outputs(6454) <= not((layer6_outputs(937)) xor (layer6_outputs(550)));
    outputs(6455) <= not(layer6_outputs(4906));
    outputs(6456) <= not((layer6_outputs(925)) xor (layer6_outputs(4920)));
    outputs(6457) <= layer6_outputs(4256);
    outputs(6458) <= layer6_outputs(1386);
    outputs(6459) <= not(layer6_outputs(1668));
    outputs(6460) <= (layer6_outputs(6623)) xor (layer6_outputs(3654));
    outputs(6461) <= not((layer6_outputs(6961)) xor (layer6_outputs(1674)));
    outputs(6462) <= not(layer6_outputs(1946)) or (layer6_outputs(2516));
    outputs(6463) <= (layer6_outputs(5803)) xor (layer6_outputs(3844));
    outputs(6464) <= layer6_outputs(6856);
    outputs(6465) <= not((layer6_outputs(1289)) and (layer6_outputs(2786)));
    outputs(6466) <= (layer6_outputs(7273)) xor (layer6_outputs(2583));
    outputs(6467) <= (layer6_outputs(626)) xor (layer6_outputs(1331));
    outputs(6468) <= (layer6_outputs(3892)) xor (layer6_outputs(5907));
    outputs(6469) <= (layer6_outputs(2773)) xor (layer6_outputs(2815));
    outputs(6470) <= not(layer6_outputs(7395));
    outputs(6471) <= (layer6_outputs(1881)) or (layer6_outputs(3377));
    outputs(6472) <= layer6_outputs(6056);
    outputs(6473) <= not(layer6_outputs(308));
    outputs(6474) <= layer6_outputs(3300);
    outputs(6475) <= layer6_outputs(2497);
    outputs(6476) <= (layer6_outputs(7431)) xor (layer6_outputs(1644));
    outputs(6477) <= not(layer6_outputs(6857));
    outputs(6478) <= layer6_outputs(5280);
    outputs(6479) <= layer6_outputs(6412);
    outputs(6480) <= layer6_outputs(594);
    outputs(6481) <= not(layer6_outputs(7159));
    outputs(6482) <= (layer6_outputs(1737)) xor (layer6_outputs(4622));
    outputs(6483) <= not(layer6_outputs(4117));
    outputs(6484) <= layer6_outputs(4563);
    outputs(6485) <= (layer6_outputs(3407)) xor (layer6_outputs(6270));
    outputs(6486) <= layer6_outputs(7338);
    outputs(6487) <= not(layer6_outputs(2111));
    outputs(6488) <= not((layer6_outputs(7088)) xor (layer6_outputs(5960)));
    outputs(6489) <= (layer6_outputs(4726)) xor (layer6_outputs(648));
    outputs(6490) <= not(layer6_outputs(2023)) or (layer6_outputs(6255));
    outputs(6491) <= not((layer6_outputs(3022)) xor (layer6_outputs(4600)));
    outputs(6492) <= layer6_outputs(2728);
    outputs(6493) <= not(layer6_outputs(2262));
    outputs(6494) <= layer6_outputs(781);
    outputs(6495) <= not(layer6_outputs(1014));
    outputs(6496) <= (layer6_outputs(3314)) or (layer6_outputs(6727));
    outputs(6497) <= layer6_outputs(4858);
    outputs(6498) <= layer6_outputs(129);
    outputs(6499) <= not(layer6_outputs(5893));
    outputs(6500) <= (layer6_outputs(7538)) and not (layer6_outputs(1748));
    outputs(6501) <= layer6_outputs(3789);
    outputs(6502) <= not((layer6_outputs(5069)) xor (layer6_outputs(543)));
    outputs(6503) <= (layer6_outputs(7199)) xor (layer6_outputs(512));
    outputs(6504) <= (layer6_outputs(130)) and not (layer6_outputs(576));
    outputs(6505) <= layer6_outputs(6477);
    outputs(6506) <= (layer6_outputs(1136)) xor (layer6_outputs(2042));
    outputs(6507) <= not(layer6_outputs(1410)) or (layer6_outputs(1793));
    outputs(6508) <= layer6_outputs(1110);
    outputs(6509) <= not(layer6_outputs(2729));
    outputs(6510) <= (layer6_outputs(5663)) and not (layer6_outputs(2377));
    outputs(6511) <= not(layer6_outputs(6488));
    outputs(6512) <= not(layer6_outputs(2340));
    outputs(6513) <= not((layer6_outputs(4848)) xor (layer6_outputs(101)));
    outputs(6514) <= not(layer6_outputs(1374));
    outputs(6515) <= (layer6_outputs(5626)) xor (layer6_outputs(482));
    outputs(6516) <= layer6_outputs(7024);
    outputs(6517) <= (layer6_outputs(2790)) and not (layer6_outputs(1434));
    outputs(6518) <= layer6_outputs(6113);
    outputs(6519) <= not((layer6_outputs(6232)) xor (layer6_outputs(4682)));
    outputs(6520) <= not((layer6_outputs(6738)) or (layer6_outputs(377)));
    outputs(6521) <= not(layer6_outputs(5357)) or (layer6_outputs(6282));
    outputs(6522) <= layer6_outputs(2933);
    outputs(6523) <= not((layer6_outputs(1384)) xor (layer6_outputs(7255)));
    outputs(6524) <= not(layer6_outputs(3468)) or (layer6_outputs(2477));
    outputs(6525) <= layer6_outputs(6992);
    outputs(6526) <= not((layer6_outputs(460)) xor (layer6_outputs(6319)));
    outputs(6527) <= not(layer6_outputs(4417));
    outputs(6528) <= layer6_outputs(5497);
    outputs(6529) <= not((layer6_outputs(7190)) xor (layer6_outputs(268)));
    outputs(6530) <= not(layer6_outputs(2092));
    outputs(6531) <= (layer6_outputs(4169)) xor (layer6_outputs(7612));
    outputs(6532) <= (layer6_outputs(6507)) and not (layer6_outputs(3388));
    outputs(6533) <= not(layer6_outputs(5084));
    outputs(6534) <= (layer6_outputs(3012)) and not (layer6_outputs(3557));
    outputs(6535) <= not(layer6_outputs(6304));
    outputs(6536) <= layer6_outputs(4231);
    outputs(6537) <= not(layer6_outputs(1134));
    outputs(6538) <= not(layer6_outputs(886));
    outputs(6539) <= layer6_outputs(3166);
    outputs(6540) <= layer6_outputs(3915);
    outputs(6541) <= layer6_outputs(4826);
    outputs(6542) <= (layer6_outputs(728)) xor (layer6_outputs(5685));
    outputs(6543) <= not(layer6_outputs(1750));
    outputs(6544) <= not(layer6_outputs(6211));
    outputs(6545) <= not((layer6_outputs(556)) xor (layer6_outputs(5495)));
    outputs(6546) <= layer6_outputs(2557);
    outputs(6547) <= layer6_outputs(4060);
    outputs(6548) <= layer6_outputs(3662);
    outputs(6549) <= layer6_outputs(3652);
    outputs(6550) <= layer6_outputs(3880);
    outputs(6551) <= layer6_outputs(7233);
    outputs(6552) <= not(layer6_outputs(3776));
    outputs(6553) <= layer6_outputs(4811);
    outputs(6554) <= not((layer6_outputs(3162)) xor (layer6_outputs(5033)));
    outputs(6555) <= layer6_outputs(3860);
    outputs(6556) <= layer6_outputs(5679);
    outputs(6557) <= not((layer6_outputs(3427)) xor (layer6_outputs(1182)));
    outputs(6558) <= not(layer6_outputs(4843)) or (layer6_outputs(620));
    outputs(6559) <= (layer6_outputs(1287)) and not (layer6_outputs(4338));
    outputs(6560) <= not((layer6_outputs(1669)) xor (layer6_outputs(236)));
    outputs(6561) <= (layer6_outputs(464)) xor (layer6_outputs(6119));
    outputs(6562) <= (layer6_outputs(2365)) or (layer6_outputs(2127));
    outputs(6563) <= layer6_outputs(7323);
    outputs(6564) <= not(layer6_outputs(466));
    outputs(6565) <= layer6_outputs(651);
    outputs(6566) <= not(layer6_outputs(1579));
    outputs(6567) <= not(layer6_outputs(4948));
    outputs(6568) <= not(layer6_outputs(6012));
    outputs(6569) <= not(layer6_outputs(5295));
    outputs(6570) <= (layer6_outputs(631)) xor (layer6_outputs(3911));
    outputs(6571) <= not((layer6_outputs(4224)) xor (layer6_outputs(3030)));
    outputs(6572) <= layer6_outputs(5263);
    outputs(6573) <= not((layer6_outputs(6290)) xor (layer6_outputs(2778)));
    outputs(6574) <= not((layer6_outputs(715)) xor (layer6_outputs(3094)));
    outputs(6575) <= layer6_outputs(6881);
    outputs(6576) <= not((layer6_outputs(3227)) xor (layer6_outputs(4099)));
    outputs(6577) <= (layer6_outputs(6527)) or (layer6_outputs(2932));
    outputs(6578) <= (layer6_outputs(6611)) xor (layer6_outputs(1038));
    outputs(6579) <= not(layer6_outputs(2750));
    outputs(6580) <= layer6_outputs(3691);
    outputs(6581) <= (layer6_outputs(6338)) xor (layer6_outputs(2578));
    outputs(6582) <= not(layer6_outputs(329));
    outputs(6583) <= not(layer6_outputs(6076));
    outputs(6584) <= not(layer6_outputs(4140));
    outputs(6585) <= not((layer6_outputs(1667)) xor (layer6_outputs(6728)));
    outputs(6586) <= not((layer6_outputs(7476)) xor (layer6_outputs(7094)));
    outputs(6587) <= layer6_outputs(2844);
    outputs(6588) <= (layer6_outputs(7102)) xor (layer6_outputs(3684));
    outputs(6589) <= not((layer6_outputs(5522)) xor (layer6_outputs(6188)));
    outputs(6590) <= (layer6_outputs(4567)) and not (layer6_outputs(815));
    outputs(6591) <= not((layer6_outputs(1393)) xor (layer6_outputs(7465)));
    outputs(6592) <= (layer6_outputs(4217)) xor (layer6_outputs(1543));
    outputs(6593) <= (layer6_outputs(5248)) and not (layer6_outputs(1452));
    outputs(6594) <= layer6_outputs(3153);
    outputs(6595) <= layer6_outputs(6569);
    outputs(6596) <= not(layer6_outputs(5375)) or (layer6_outputs(6040));
    outputs(6597) <= not((layer6_outputs(3169)) xor (layer6_outputs(3885)));
    outputs(6598) <= not(layer6_outputs(7139));
    outputs(6599) <= not(layer6_outputs(3556));
    outputs(6600) <= (layer6_outputs(6624)) xor (layer6_outputs(3582));
    outputs(6601) <= not((layer6_outputs(2495)) xor (layer6_outputs(4614)));
    outputs(6602) <= layer6_outputs(3679);
    outputs(6603) <= not((layer6_outputs(729)) xor (layer6_outputs(2175)));
    outputs(6604) <= (layer6_outputs(4972)) and (layer6_outputs(2659));
    outputs(6605) <= not(layer6_outputs(3021)) or (layer6_outputs(3591));
    outputs(6606) <= layer6_outputs(3455);
    outputs(6607) <= (layer6_outputs(171)) or (layer6_outputs(1993));
    outputs(6608) <= layer6_outputs(3953);
    outputs(6609) <= not((layer6_outputs(3032)) xor (layer6_outputs(6938)));
    outputs(6610) <= layer6_outputs(1117);
    outputs(6611) <= not(layer6_outputs(4628));
    outputs(6612) <= (layer6_outputs(4067)) xor (layer6_outputs(1675));
    outputs(6613) <= not(layer6_outputs(4628));
    outputs(6614) <= not((layer6_outputs(3839)) xor (layer6_outputs(4394)));
    outputs(6615) <= not(layer6_outputs(6076));
    outputs(6616) <= (layer6_outputs(5414)) xor (layer6_outputs(2484));
    outputs(6617) <= not(layer6_outputs(7336));
    outputs(6618) <= (layer6_outputs(2264)) xor (layer6_outputs(3922));
    outputs(6619) <= (layer6_outputs(5235)) and not (layer6_outputs(7647));
    outputs(6620) <= layer6_outputs(3788);
    outputs(6621) <= not(layer6_outputs(4337));
    outputs(6622) <= not(layer6_outputs(419));
    outputs(6623) <= not(layer6_outputs(4984));
    outputs(6624) <= not(layer6_outputs(1424));
    outputs(6625) <= (layer6_outputs(6756)) xor (layer6_outputs(6892));
    outputs(6626) <= not(layer6_outputs(4329));
    outputs(6627) <= layer6_outputs(1787);
    outputs(6628) <= layer6_outputs(4465);
    outputs(6629) <= (layer6_outputs(2838)) and not (layer6_outputs(4603));
    outputs(6630) <= layer6_outputs(5523);
    outputs(6631) <= layer6_outputs(5998);
    outputs(6632) <= (layer6_outputs(4110)) xor (layer6_outputs(6686));
    outputs(6633) <= (layer6_outputs(4780)) xor (layer6_outputs(5465));
    outputs(6634) <= not((layer6_outputs(4244)) xor (layer6_outputs(6696)));
    outputs(6635) <= (layer6_outputs(4404)) or (layer6_outputs(7167));
    outputs(6636) <= (layer6_outputs(2568)) xor (layer6_outputs(3344));
    outputs(6637) <= not(layer6_outputs(6673));
    outputs(6638) <= (layer6_outputs(6871)) xor (layer6_outputs(2352));
    outputs(6639) <= not(layer6_outputs(5833));
    outputs(6640) <= layer6_outputs(2533);
    outputs(6641) <= (layer6_outputs(7415)) xor (layer6_outputs(4358));
    outputs(6642) <= not(layer6_outputs(5979));
    outputs(6643) <= not(layer6_outputs(1463));
    outputs(6644) <= (layer6_outputs(2775)) and not (layer6_outputs(1121));
    outputs(6645) <= layer6_outputs(93);
    outputs(6646) <= (layer6_outputs(6776)) and (layer6_outputs(416));
    outputs(6647) <= (layer6_outputs(5450)) xor (layer6_outputs(3512));
    outputs(6648) <= (layer6_outputs(6183)) xor (layer6_outputs(6108));
    outputs(6649) <= (layer6_outputs(152)) and (layer6_outputs(1185));
    outputs(6650) <= layer6_outputs(3332);
    outputs(6651) <= layer6_outputs(1482);
    outputs(6652) <= not((layer6_outputs(1034)) xor (layer6_outputs(5486)));
    outputs(6653) <= not((layer6_outputs(6080)) xor (layer6_outputs(3295)));
    outputs(6654) <= layer6_outputs(2399);
    outputs(6655) <= (layer6_outputs(4165)) xor (layer6_outputs(3842));
    outputs(6656) <= not(layer6_outputs(2462));
    outputs(6657) <= not(layer6_outputs(6431)) or (layer6_outputs(1360));
    outputs(6658) <= not((layer6_outputs(6387)) xor (layer6_outputs(2373)));
    outputs(6659) <= (layer6_outputs(5070)) xor (layer6_outputs(4746));
    outputs(6660) <= layer6_outputs(1241);
    outputs(6661) <= not((layer6_outputs(2583)) xor (layer6_outputs(548)));
    outputs(6662) <= not(layer6_outputs(6582));
    outputs(6663) <= not(layer6_outputs(330));
    outputs(6664) <= layer6_outputs(3619);
    outputs(6665) <= not(layer6_outputs(7418));
    outputs(6666) <= (layer6_outputs(2015)) xor (layer6_outputs(2698));
    outputs(6667) <= layer6_outputs(2882);
    outputs(6668) <= (layer6_outputs(4601)) xor (layer6_outputs(2606));
    outputs(6669) <= (layer6_outputs(3063)) or (layer6_outputs(776));
    outputs(6670) <= layer6_outputs(1276);
    outputs(6671) <= not(layer6_outputs(6822));
    outputs(6672) <= layer6_outputs(6688);
    outputs(6673) <= layer6_outputs(6022);
    outputs(6674) <= (layer6_outputs(5541)) xor (layer6_outputs(3545));
    outputs(6675) <= layer6_outputs(3703);
    outputs(6676) <= (layer6_outputs(72)) xor (layer6_outputs(1895));
    outputs(6677) <= not(layer6_outputs(1365));
    outputs(6678) <= not(layer6_outputs(3470));
    outputs(6679) <= layer6_outputs(1301);
    outputs(6680) <= layer6_outputs(3800);
    outputs(6681) <= layer6_outputs(5879);
    outputs(6682) <= (layer6_outputs(5057)) xor (layer6_outputs(4724));
    outputs(6683) <= layer6_outputs(5386);
    outputs(6684) <= layer6_outputs(1531);
    outputs(6685) <= layer6_outputs(4590);
    outputs(6686) <= (layer6_outputs(6693)) or (layer6_outputs(7392));
    outputs(6687) <= not(layer6_outputs(5224)) or (layer6_outputs(7583));
    outputs(6688) <= not((layer6_outputs(2028)) xor (layer6_outputs(574)));
    outputs(6689) <= not((layer6_outputs(2609)) xor (layer6_outputs(2444)));
    outputs(6690) <= layer6_outputs(2509);
    outputs(6691) <= layer6_outputs(4202);
    outputs(6692) <= (layer6_outputs(6744)) or (layer6_outputs(4888));
    outputs(6693) <= (layer6_outputs(175)) xor (layer6_outputs(6510));
    outputs(6694) <= not(layer6_outputs(4886));
    outputs(6695) <= not(layer6_outputs(867));
    outputs(6696) <= (layer6_outputs(7284)) or (layer6_outputs(7665));
    outputs(6697) <= layer6_outputs(7629);
    outputs(6698) <= not(layer6_outputs(3161));
    outputs(6699) <= layer6_outputs(891);
    outputs(6700) <= not(layer6_outputs(3549));
    outputs(6701) <= not(layer6_outputs(5955));
    outputs(6702) <= not(layer6_outputs(2314));
    outputs(6703) <= (layer6_outputs(6843)) and not (layer6_outputs(2241));
    outputs(6704) <= not(layer6_outputs(1418));
    outputs(6705) <= layer6_outputs(1373);
    outputs(6706) <= not((layer6_outputs(1647)) xor (layer6_outputs(4219)));
    outputs(6707) <= not((layer6_outputs(2425)) xor (layer6_outputs(826)));
    outputs(6708) <= not((layer6_outputs(2346)) xor (layer6_outputs(1965)));
    outputs(6709) <= layer6_outputs(4558);
    outputs(6710) <= not(layer6_outputs(6509));
    outputs(6711) <= layer6_outputs(7292);
    outputs(6712) <= not((layer6_outputs(4270)) xor (layer6_outputs(187)));
    outputs(6713) <= layer6_outputs(1244);
    outputs(6714) <= not((layer6_outputs(639)) xor (layer6_outputs(1947)));
    outputs(6715) <= not(layer6_outputs(4359));
    outputs(6716) <= not((layer6_outputs(1249)) or (layer6_outputs(6745)));
    outputs(6717) <= layer6_outputs(5416);
    outputs(6718) <= not(layer6_outputs(5651));
    outputs(6719) <= (layer6_outputs(5546)) xor (layer6_outputs(1698));
    outputs(6720) <= (layer6_outputs(177)) xor (layer6_outputs(420));
    outputs(6721) <= not(layer6_outputs(6070)) or (layer6_outputs(3475));
    outputs(6722) <= (layer6_outputs(5763)) xor (layer6_outputs(1112));
    outputs(6723) <= not((layer6_outputs(1195)) xor (layer6_outputs(4731)));
    outputs(6724) <= not(layer6_outputs(827));
    outputs(6725) <= (layer6_outputs(2672)) xor (layer6_outputs(7062));
    outputs(6726) <= not(layer6_outputs(787));
    outputs(6727) <= (layer6_outputs(4425)) xor (layer6_outputs(5928));
    outputs(6728) <= layer6_outputs(4239);
    outputs(6729) <= (layer6_outputs(4567)) and not (layer6_outputs(6236));
    outputs(6730) <= not(layer6_outputs(5000));
    outputs(6731) <= not((layer6_outputs(3905)) xor (layer6_outputs(3572)));
    outputs(6732) <= layer6_outputs(5270);
    outputs(6733) <= layer6_outputs(4145);
    outputs(6734) <= layer6_outputs(5356);
    outputs(6735) <= (layer6_outputs(4201)) and not (layer6_outputs(4919));
    outputs(6736) <= (layer6_outputs(3653)) or (layer6_outputs(3183));
    outputs(6737) <= not(layer6_outputs(6722));
    outputs(6738) <= layer6_outputs(2645);
    outputs(6739) <= not((layer6_outputs(5461)) xor (layer6_outputs(6993)));
    outputs(6740) <= layer6_outputs(540);
    outputs(6741) <= not(layer6_outputs(308));
    outputs(6742) <= not(layer6_outputs(7656));
    outputs(6743) <= layer6_outputs(5679);
    outputs(6744) <= not(layer6_outputs(3367));
    outputs(6745) <= not(layer6_outputs(4193));
    outputs(6746) <= layer6_outputs(5120);
    outputs(6747) <= not((layer6_outputs(6734)) xor (layer6_outputs(7499)));
    outputs(6748) <= not((layer6_outputs(1143)) xor (layer6_outputs(219)));
    outputs(6749) <= not((layer6_outputs(7553)) xor (layer6_outputs(4142)));
    outputs(6750) <= not((layer6_outputs(721)) xor (layer6_outputs(5781)));
    outputs(6751) <= not(layer6_outputs(6143));
    outputs(6752) <= layer6_outputs(856);
    outputs(6753) <= not(layer6_outputs(6554));
    outputs(6754) <= not(layer6_outputs(4922));
    outputs(6755) <= not(layer6_outputs(3755));
    outputs(6756) <= layer6_outputs(1163);
    outputs(6757) <= not((layer6_outputs(5112)) xor (layer6_outputs(6306)));
    outputs(6758) <= layer6_outputs(521);
    outputs(6759) <= not(layer6_outputs(2992));
    outputs(6760) <= not((layer6_outputs(5355)) xor (layer6_outputs(4094)));
    outputs(6761) <= layer6_outputs(1076);
    outputs(6762) <= not((layer6_outputs(5733)) xor (layer6_outputs(59)));
    outputs(6763) <= not((layer6_outputs(5809)) xor (layer6_outputs(5313)));
    outputs(6764) <= not(layer6_outputs(7166));
    outputs(6765) <= layer6_outputs(4178);
    outputs(6766) <= layer6_outputs(6117);
    outputs(6767) <= layer6_outputs(3379);
    outputs(6768) <= not(layer6_outputs(523));
    outputs(6769) <= not(layer6_outputs(5301)) or (layer6_outputs(781));
    outputs(6770) <= not(layer6_outputs(4693)) or (layer6_outputs(5699));
    outputs(6771) <= layer6_outputs(1845);
    outputs(6772) <= not((layer6_outputs(3648)) and (layer6_outputs(1291)));
    outputs(6773) <= layer6_outputs(4878);
    outputs(6774) <= not(layer6_outputs(4478));
    outputs(6775) <= not(layer6_outputs(4951));
    outputs(6776) <= layer6_outputs(4450);
    outputs(6777) <= layer6_outputs(1417);
    outputs(6778) <= layer6_outputs(5382);
    outputs(6779) <= not(layer6_outputs(5254));
    outputs(6780) <= layer6_outputs(4557);
    outputs(6781) <= (layer6_outputs(7120)) and not (layer6_outputs(4422));
    outputs(6782) <= layer6_outputs(2797);
    outputs(6783) <= layer6_outputs(1933);
    outputs(6784) <= not(layer6_outputs(7042));
    outputs(6785) <= not(layer6_outputs(2917)) or (layer6_outputs(2275));
    outputs(6786) <= not((layer6_outputs(502)) xor (layer6_outputs(6006)));
    outputs(6787) <= (layer6_outputs(4181)) or (layer6_outputs(2351));
    outputs(6788) <= layer6_outputs(2028);
    outputs(6789) <= not(layer6_outputs(2061));
    outputs(6790) <= not(layer6_outputs(1203));
    outputs(6791) <= not(layer6_outputs(2768));
    outputs(6792) <= layer6_outputs(5374);
    outputs(6793) <= not(layer6_outputs(4249));
    outputs(6794) <= (layer6_outputs(2204)) xor (layer6_outputs(5704));
    outputs(6795) <= not(layer6_outputs(6446));
    outputs(6796) <= not(layer6_outputs(1269));
    outputs(6797) <= (layer6_outputs(820)) or (layer6_outputs(5846));
    outputs(6798) <= layer6_outputs(1260);
    outputs(6799) <= not(layer6_outputs(1935));
    outputs(6800) <= (layer6_outputs(5190)) xor (layer6_outputs(982));
    outputs(6801) <= layer6_outputs(4499);
    outputs(6802) <= not((layer6_outputs(2564)) xor (layer6_outputs(868)));
    outputs(6803) <= not((layer6_outputs(3983)) xor (layer6_outputs(7501)));
    outputs(6804) <= (layer6_outputs(2362)) xor (layer6_outputs(6818));
    outputs(6805) <= layer6_outputs(1785);
    outputs(6806) <= layer6_outputs(2000);
    outputs(6807) <= (layer6_outputs(3874)) xor (layer6_outputs(2849));
    outputs(6808) <= layer6_outputs(5904);
    outputs(6809) <= layer6_outputs(5211);
    outputs(6810) <= not((layer6_outputs(6842)) xor (layer6_outputs(5448)));
    outputs(6811) <= layer6_outputs(6894);
    outputs(6812) <= not(layer6_outputs(3291));
    outputs(6813) <= (layer6_outputs(1296)) xor (layer6_outputs(6912));
    outputs(6814) <= (layer6_outputs(3508)) xor (layer6_outputs(4233));
    outputs(6815) <= not(layer6_outputs(588)) or (layer6_outputs(947));
    outputs(6816) <= not(layer6_outputs(6866));
    outputs(6817) <= not(layer6_outputs(806));
    outputs(6818) <= not(layer6_outputs(4691));
    outputs(6819) <= (layer6_outputs(918)) xor (layer6_outputs(6950));
    outputs(6820) <= layer6_outputs(1417);
    outputs(6821) <= layer6_outputs(3256);
    outputs(6822) <= not(layer6_outputs(7558));
    outputs(6823) <= layer6_outputs(1432);
    outputs(6824) <= (layer6_outputs(7451)) xor (layer6_outputs(2255));
    outputs(6825) <= not(layer6_outputs(4779));
    outputs(6826) <= layer6_outputs(3217);
    outputs(6827) <= not(layer6_outputs(1495));
    outputs(6828) <= layer6_outputs(3935);
    outputs(6829) <= not(layer6_outputs(5769));
    outputs(6830) <= (layer6_outputs(2954)) xor (layer6_outputs(4137));
    outputs(6831) <= not(layer6_outputs(2872));
    outputs(6832) <= not(layer6_outputs(6909));
    outputs(6833) <= (layer6_outputs(3755)) xor (layer6_outputs(4858));
    outputs(6834) <= (layer6_outputs(6679)) and (layer6_outputs(410));
    outputs(6835) <= not(layer6_outputs(4432));
    outputs(6836) <= not((layer6_outputs(6304)) xor (layer6_outputs(553)));
    outputs(6837) <= not(layer6_outputs(3069)) or (layer6_outputs(6286));
    outputs(6838) <= not(layer6_outputs(2840));
    outputs(6839) <= layer6_outputs(4190);
    outputs(6840) <= (layer6_outputs(1516)) xor (layer6_outputs(2570));
    outputs(6841) <= (layer6_outputs(4050)) or (layer6_outputs(7213));
    outputs(6842) <= not((layer6_outputs(3257)) and (layer6_outputs(4803)));
    outputs(6843) <= layer6_outputs(4545);
    outputs(6844) <= (layer6_outputs(4214)) xor (layer6_outputs(1101));
    outputs(6845) <= not(layer6_outputs(3368));
    outputs(6846) <= not((layer6_outputs(5257)) xor (layer6_outputs(6435)));
    outputs(6847) <= (layer6_outputs(2143)) xor (layer6_outputs(948));
    outputs(6848) <= not((layer6_outputs(4677)) or (layer6_outputs(5527)));
    outputs(6849) <= not((layer6_outputs(4223)) xor (layer6_outputs(817)));
    outputs(6850) <= not((layer6_outputs(3208)) and (layer6_outputs(1269)));
    outputs(6851) <= (layer6_outputs(3002)) xor (layer6_outputs(1298));
    outputs(6852) <= (layer6_outputs(582)) and not (layer6_outputs(4030));
    outputs(6853) <= not(layer6_outputs(6111)) or (layer6_outputs(5471));
    outputs(6854) <= not(layer6_outputs(18));
    outputs(6855) <= layer6_outputs(3224);
    outputs(6856) <= (layer6_outputs(102)) and not (layer6_outputs(247));
    outputs(6857) <= (layer6_outputs(7349)) xor (layer6_outputs(6103));
    outputs(6858) <= not(layer6_outputs(2393));
    outputs(6859) <= (layer6_outputs(4559)) and (layer6_outputs(7674));
    outputs(6860) <= not((layer6_outputs(1548)) xor (layer6_outputs(5018)));
    outputs(6861) <= not((layer6_outputs(4212)) xor (layer6_outputs(923)));
    outputs(6862) <= (layer6_outputs(2538)) xor (layer6_outputs(4491));
    outputs(6863) <= not((layer6_outputs(2792)) xor (layer6_outputs(6713)));
    outputs(6864) <= not((layer6_outputs(5442)) xor (layer6_outputs(7454)));
    outputs(6865) <= not((layer6_outputs(3154)) xor (layer6_outputs(1128)));
    outputs(6866) <= not((layer6_outputs(1085)) xor (layer6_outputs(196)));
    outputs(6867) <= not(layer6_outputs(1328));
    outputs(6868) <= (layer6_outputs(5514)) xor (layer6_outputs(2289));
    outputs(6869) <= not((layer6_outputs(5124)) xor (layer6_outputs(5818)));
    outputs(6870) <= not((layer6_outputs(4514)) xor (layer6_outputs(2027)));
    outputs(6871) <= layer6_outputs(1854);
    outputs(6872) <= layer6_outputs(387);
    outputs(6873) <= not(layer6_outputs(2199)) or (layer6_outputs(910));
    outputs(6874) <= layer6_outputs(5856);
    outputs(6875) <= layer6_outputs(6917);
    outputs(6876) <= not((layer6_outputs(4154)) and (layer6_outputs(6347)));
    outputs(6877) <= (layer6_outputs(1834)) and not (layer6_outputs(2706));
    outputs(6878) <= not((layer6_outputs(6458)) xor (layer6_outputs(3481)));
    outputs(6879) <= not(layer6_outputs(4496));
    outputs(6880) <= (layer6_outputs(751)) xor (layer6_outputs(4586));
    outputs(6881) <= not(layer6_outputs(5324)) or (layer6_outputs(6327));
    outputs(6882) <= not(layer6_outputs(1617)) or (layer6_outputs(5956));
    outputs(6883) <= not(layer6_outputs(2959));
    outputs(6884) <= not((layer6_outputs(6413)) xor (layer6_outputs(331)));
    outputs(6885) <= (layer6_outputs(6142)) xor (layer6_outputs(5117));
    outputs(6886) <= (layer6_outputs(7557)) xor (layer6_outputs(3310));
    outputs(6887) <= layer6_outputs(402);
    outputs(6888) <= layer6_outputs(2659);
    outputs(6889) <= not(layer6_outputs(7091));
    outputs(6890) <= layer6_outputs(4732);
    outputs(6891) <= layer6_outputs(1614);
    outputs(6892) <= not((layer6_outputs(415)) and (layer6_outputs(2721)));
    outputs(6893) <= not((layer6_outputs(107)) and (layer6_outputs(828)));
    outputs(6894) <= layer6_outputs(2494);
    outputs(6895) <= not(layer6_outputs(3338)) or (layer6_outputs(782));
    outputs(6896) <= layer6_outputs(4926);
    outputs(6897) <= layer6_outputs(6848);
    outputs(6898) <= layer6_outputs(3100);
    outputs(6899) <= not((layer6_outputs(3267)) xor (layer6_outputs(1563)));
    outputs(6900) <= layer6_outputs(3322);
    outputs(6901) <= not(layer6_outputs(763));
    outputs(6902) <= not(layer6_outputs(6644));
    outputs(6903) <= layer6_outputs(6731);
    outputs(6904) <= layer6_outputs(3371);
    outputs(6905) <= not(layer6_outputs(5399));
    outputs(6906) <= not((layer6_outputs(3037)) xor (layer6_outputs(6849)));
    outputs(6907) <= layer6_outputs(5557);
    outputs(6908) <= (layer6_outputs(4879)) xor (layer6_outputs(753));
    outputs(6909) <= not((layer6_outputs(1724)) xor (layer6_outputs(2227)));
    outputs(6910) <= not(layer6_outputs(6809));
    outputs(6911) <= (layer6_outputs(3717)) or (layer6_outputs(1008));
    outputs(6912) <= not(layer6_outputs(1527));
    outputs(6913) <= layer6_outputs(677);
    outputs(6914) <= layer6_outputs(2855);
    outputs(6915) <= (layer6_outputs(1813)) and (layer6_outputs(5760));
    outputs(6916) <= (layer6_outputs(5820)) xor (layer6_outputs(3873));
    outputs(6917) <= not(layer6_outputs(4351));
    outputs(6918) <= not(layer6_outputs(5987));
    outputs(6919) <= not(layer6_outputs(148));
    outputs(6920) <= not(layer6_outputs(2360));
    outputs(6921) <= not(layer6_outputs(1938));
    outputs(6922) <= not(layer6_outputs(2910));
    outputs(6923) <= (layer6_outputs(3387)) and not (layer6_outputs(1405));
    outputs(6924) <= (layer6_outputs(4738)) xor (layer6_outputs(5066));
    outputs(6925) <= layer6_outputs(5287);
    outputs(6926) <= layer6_outputs(6697);
    outputs(6927) <= layer6_outputs(2020);
    outputs(6928) <= not((layer6_outputs(2700)) xor (layer6_outputs(15)));
    outputs(6929) <= not(layer6_outputs(2771));
    outputs(6930) <= (layer6_outputs(7278)) and not (layer6_outputs(2697));
    outputs(6931) <= not((layer6_outputs(3721)) and (layer6_outputs(1965)));
    outputs(6932) <= layer6_outputs(5086);
    outputs(6933) <= not((layer6_outputs(2870)) xor (layer6_outputs(5810)));
    outputs(6934) <= layer6_outputs(6949);
    outputs(6935) <= layer6_outputs(4938);
    outputs(6936) <= not((layer6_outputs(7320)) xor (layer6_outputs(3375)));
    outputs(6937) <= not(layer6_outputs(4310));
    outputs(6938) <= (layer6_outputs(1580)) and not (layer6_outputs(2837));
    outputs(6939) <= layer6_outputs(2393);
    outputs(6940) <= (layer6_outputs(819)) and not (layer6_outputs(5097));
    outputs(6941) <= not(layer6_outputs(2121));
    outputs(6942) <= not(layer6_outputs(2384));
    outputs(6943) <= not(layer6_outputs(19));
    outputs(6944) <= (layer6_outputs(784)) xor (layer6_outputs(4755));
    outputs(6945) <= not(layer6_outputs(3879));
    outputs(6946) <= layer6_outputs(6260);
    outputs(6947) <= layer6_outputs(4871);
    outputs(6948) <= not(layer6_outputs(5213));
    outputs(6949) <= layer6_outputs(4512);
    outputs(6950) <= layer6_outputs(615);
    outputs(6951) <= not(layer6_outputs(3335));
    outputs(6952) <= not((layer6_outputs(1278)) and (layer6_outputs(45)));
    outputs(6953) <= layer6_outputs(6066);
    outputs(6954) <= not(layer6_outputs(601));
    outputs(6955) <= layer6_outputs(5888);
    outputs(6956) <= (layer6_outputs(7412)) xor (layer6_outputs(3764));
    outputs(6957) <= layer6_outputs(1290);
    outputs(6958) <= layer6_outputs(3868);
    outputs(6959) <= layer6_outputs(7364);
    outputs(6960) <= not(layer6_outputs(3495)) or (layer6_outputs(7340));
    outputs(6961) <= (layer6_outputs(5727)) xor (layer6_outputs(4688));
    outputs(6962) <= not((layer6_outputs(870)) or (layer6_outputs(1973)));
    outputs(6963) <= layer6_outputs(5613);
    outputs(6964) <= (layer6_outputs(5296)) and (layer6_outputs(5510));
    outputs(6965) <= (layer6_outputs(6466)) xor (layer6_outputs(3077));
    outputs(6966) <= not(layer6_outputs(2137));
    outputs(6967) <= (layer6_outputs(1859)) xor (layer6_outputs(2197));
    outputs(6968) <= not(layer6_outputs(42));
    outputs(6969) <= not(layer6_outputs(4193));
    outputs(6970) <= not(layer6_outputs(4129)) or (layer6_outputs(7189));
    outputs(6971) <= layer6_outputs(3116);
    outputs(6972) <= not(layer6_outputs(5082));
    outputs(6973) <= layer6_outputs(6075);
    outputs(6974) <= layer6_outputs(2323);
    outputs(6975) <= not(layer6_outputs(3283));
    outputs(6976) <= (layer6_outputs(4649)) xor (layer6_outputs(4864));
    outputs(6977) <= (layer6_outputs(2666)) xor (layer6_outputs(2615));
    outputs(6978) <= layer6_outputs(7247);
    outputs(6979) <= not((layer6_outputs(7066)) or (layer6_outputs(5783)));
    outputs(6980) <= not(layer6_outputs(1860));
    outputs(6981) <= not(layer6_outputs(1140));
    outputs(6982) <= not(layer6_outputs(4902));
    outputs(6983) <= (layer6_outputs(3482)) and (layer6_outputs(6707));
    outputs(6984) <= not(layer6_outputs(1464));
    outputs(6985) <= not((layer6_outputs(4480)) xor (layer6_outputs(2807)));
    outputs(6986) <= (layer6_outputs(6116)) and not (layer6_outputs(644));
    outputs(6987) <= layer6_outputs(48);
    outputs(6988) <= layer6_outputs(4388);
    outputs(6989) <= not((layer6_outputs(499)) or (layer6_outputs(3210)));
    outputs(6990) <= layer6_outputs(6218);
    outputs(6991) <= not(layer6_outputs(2196));
    outputs(6992) <= not(layer6_outputs(1415)) or (layer6_outputs(2374));
    outputs(6993) <= layer6_outputs(416);
    outputs(6994) <= (layer6_outputs(4153)) and not (layer6_outputs(6916));
    outputs(6995) <= (layer6_outputs(3763)) xor (layer6_outputs(5567));
    outputs(6996) <= (layer6_outputs(4275)) and (layer6_outputs(3645));
    outputs(6997) <= not(layer6_outputs(4295));
    outputs(6998) <= not((layer6_outputs(4876)) xor (layer6_outputs(2866)));
    outputs(6999) <= (layer6_outputs(2796)) xor (layer6_outputs(1309));
    outputs(7000) <= (layer6_outputs(7227)) or (layer6_outputs(355));
    outputs(7001) <= layer6_outputs(2138);
    outputs(7002) <= not(layer6_outputs(828)) or (layer6_outputs(5585));
    outputs(7003) <= layer6_outputs(5742);
    outputs(7004) <= not(layer6_outputs(6181));
    outputs(7005) <= (layer6_outputs(2319)) and not (layer6_outputs(4213));
    outputs(7006) <= not(layer6_outputs(6345)) or (layer6_outputs(4384));
    outputs(7007) <= layer6_outputs(6549);
    outputs(7008) <= layer6_outputs(5341);
    outputs(7009) <= (layer6_outputs(6495)) xor (layer6_outputs(6930));
    outputs(7010) <= not(layer6_outputs(7625));
    outputs(7011) <= not(layer6_outputs(3152));
    outputs(7012) <= layer6_outputs(2553);
    outputs(7013) <= not(layer6_outputs(146));
    outputs(7014) <= not(layer6_outputs(1726));
    outputs(7015) <= not(layer6_outputs(1126));
    outputs(7016) <= (layer6_outputs(1256)) or (layer6_outputs(1370));
    outputs(7017) <= layer6_outputs(2794);
    outputs(7018) <= layer6_outputs(847);
    outputs(7019) <= not(layer6_outputs(7393)) or (layer6_outputs(1235));
    outputs(7020) <= (layer6_outputs(3507)) and (layer6_outputs(909));
    outputs(7021) <= not((layer6_outputs(5642)) and (layer6_outputs(3414)));
    outputs(7022) <= (layer6_outputs(6908)) and (layer6_outputs(6762));
    outputs(7023) <= layer6_outputs(5773);
    outputs(7024) <= not(layer6_outputs(713)) or (layer6_outputs(4684));
    outputs(7025) <= layer6_outputs(1717);
    outputs(7026) <= (layer6_outputs(5719)) and (layer6_outputs(3811));
    outputs(7027) <= layer6_outputs(7399);
    outputs(7028) <= layer6_outputs(4761);
    outputs(7029) <= not((layer6_outputs(3556)) and (layer6_outputs(5662)));
    outputs(7030) <= not(layer6_outputs(5961));
    outputs(7031) <= not(layer6_outputs(1963));
    outputs(7032) <= layer6_outputs(5371);
    outputs(7033) <= layer6_outputs(2946);
    outputs(7034) <= (layer6_outputs(4832)) and (layer6_outputs(4588));
    outputs(7035) <= layer6_outputs(2414);
    outputs(7036) <= not((layer6_outputs(3637)) xor (layer6_outputs(5435)));
    outputs(7037) <= (layer6_outputs(4399)) and not (layer6_outputs(4472));
    outputs(7038) <= not(layer6_outputs(7237));
    outputs(7039) <= not(layer6_outputs(7537));
    outputs(7040) <= not(layer6_outputs(3450));
    outputs(7041) <= layer6_outputs(3040);
    outputs(7042) <= not(layer6_outputs(216));
    outputs(7043) <= not(layer6_outputs(5682));
    outputs(7044) <= (layer6_outputs(7457)) xor (layer6_outputs(5671));
    outputs(7045) <= not(layer6_outputs(4626));
    outputs(7046) <= layer6_outputs(3832);
    outputs(7047) <= layer6_outputs(4306);
    outputs(7048) <= not(layer6_outputs(5045));
    outputs(7049) <= not((layer6_outputs(7082)) xor (layer6_outputs(4007)));
    outputs(7050) <= not(layer6_outputs(2308)) or (layer6_outputs(94));
    outputs(7051) <= layer6_outputs(6894);
    outputs(7052) <= (layer6_outputs(4854)) and not (layer6_outputs(2927));
    outputs(7053) <= layer6_outputs(408);
    outputs(7054) <= not(layer6_outputs(5981));
    outputs(7055) <= (layer6_outputs(5763)) and not (layer6_outputs(4685));
    outputs(7056) <= layer6_outputs(7412);
    outputs(7057) <= layer6_outputs(6300);
    outputs(7058) <= not(layer6_outputs(1975));
    outputs(7059) <= not(layer6_outputs(4053));
    outputs(7060) <= not(layer6_outputs(6514)) or (layer6_outputs(291));
    outputs(7061) <= layer6_outputs(599);
    outputs(7062) <= not(layer6_outputs(6285));
    outputs(7063) <= not(layer6_outputs(1541));
    outputs(7064) <= (layer6_outputs(6622)) and not (layer6_outputs(3525));
    outputs(7065) <= not(layer6_outputs(4549));
    outputs(7066) <= not(layer6_outputs(1313)) or (layer6_outputs(3896));
    outputs(7067) <= layer6_outputs(4006);
    outputs(7068) <= layer6_outputs(565);
    outputs(7069) <= (layer6_outputs(4768)) and (layer6_outputs(3447));
    outputs(7070) <= layer6_outputs(6318);
    outputs(7071) <= not(layer6_outputs(326));
    outputs(7072) <= not(layer6_outputs(7341));
    outputs(7073) <= (layer6_outputs(2063)) and not (layer6_outputs(5869));
    outputs(7074) <= not((layer6_outputs(2928)) xor (layer6_outputs(4725)));
    outputs(7075) <= layer6_outputs(5666);
    outputs(7076) <= (layer6_outputs(6294)) xor (layer6_outputs(5599));
    outputs(7077) <= layer6_outputs(4758);
    outputs(7078) <= not((layer6_outputs(2489)) xor (layer6_outputs(7125)));
    outputs(7079) <= (layer6_outputs(4034)) xor (layer6_outputs(1200));
    outputs(7080) <= not((layer6_outputs(561)) xor (layer6_outputs(2491)));
    outputs(7081) <= not(layer6_outputs(4818));
    outputs(7082) <= layer6_outputs(6932);
    outputs(7083) <= (layer6_outputs(7286)) xor (layer6_outputs(6775));
    outputs(7084) <= not((layer6_outputs(3988)) xor (layer6_outputs(5041)));
    outputs(7085) <= not(layer6_outputs(6590));
    outputs(7086) <= layer6_outputs(5202);
    outputs(7087) <= not(layer6_outputs(7567));
    outputs(7088) <= (layer6_outputs(1695)) and not (layer6_outputs(3352));
    outputs(7089) <= layer6_outputs(3040);
    outputs(7090) <= not((layer6_outputs(1700)) xor (layer6_outputs(6107)));
    outputs(7091) <= not(layer6_outputs(6612));
    outputs(7092) <= layer6_outputs(4921);
    outputs(7093) <= layer6_outputs(3541);
    outputs(7094) <= layer6_outputs(1552);
    outputs(7095) <= layer6_outputs(5140);
    outputs(7096) <= layer6_outputs(7364);
    outputs(7097) <= layer6_outputs(7522);
    outputs(7098) <= layer6_outputs(1955);
    outputs(7099) <= not((layer6_outputs(1946)) xor (layer6_outputs(1737)));
    outputs(7100) <= layer6_outputs(5215);
    outputs(7101) <= not(layer6_outputs(2202));
    outputs(7102) <= not(layer6_outputs(7545));
    outputs(7103) <= layer6_outputs(6887);
    outputs(7104) <= layer6_outputs(55);
    outputs(7105) <= layer6_outputs(6572);
    outputs(7106) <= layer6_outputs(4368);
    outputs(7107) <= not(layer6_outputs(3382));
    outputs(7108) <= (layer6_outputs(6265)) xor (layer6_outputs(1694));
    outputs(7109) <= not(layer6_outputs(7154));
    outputs(7110) <= (layer6_outputs(2207)) xor (layer6_outputs(7658));
    outputs(7111) <= layer6_outputs(4471);
    outputs(7112) <= not((layer6_outputs(68)) xor (layer6_outputs(3291)));
    outputs(7113) <= not((layer6_outputs(1066)) xor (layer6_outputs(1546)));
    outputs(7114) <= layer6_outputs(3194);
    outputs(7115) <= (layer6_outputs(4319)) and (layer6_outputs(5700));
    outputs(7116) <= not(layer6_outputs(3165));
    outputs(7117) <= not((layer6_outputs(6036)) xor (layer6_outputs(7288)));
    outputs(7118) <= not(layer6_outputs(6220));
    outputs(7119) <= (layer6_outputs(3653)) and (layer6_outputs(4532));
    outputs(7120) <= not((layer6_outputs(4844)) xor (layer6_outputs(4016)));
    outputs(7121) <= not(layer6_outputs(3157));
    outputs(7122) <= not(layer6_outputs(6086));
    outputs(7123) <= not((layer6_outputs(6767)) xor (layer6_outputs(5279)));
    outputs(7124) <= layer6_outputs(5288);
    outputs(7125) <= not(layer6_outputs(5811));
    outputs(7126) <= layer6_outputs(3883);
    outputs(7127) <= layer6_outputs(3529);
    outputs(7128) <= not((layer6_outputs(3032)) or (layer6_outputs(6206)));
    outputs(7129) <= not(layer6_outputs(787));
    outputs(7130) <= not(layer6_outputs(5175));
    outputs(7131) <= not((layer6_outputs(3695)) xor (layer6_outputs(4657)));
    outputs(7132) <= not(layer6_outputs(5158));
    outputs(7133) <= not(layer6_outputs(4138));
    outputs(7134) <= not((layer6_outputs(5669)) xor (layer6_outputs(3569)));
    outputs(7135) <= layer6_outputs(2911);
    outputs(7136) <= layer6_outputs(3366);
    outputs(7137) <= not(layer6_outputs(2303));
    outputs(7138) <= (layer6_outputs(3692)) and not (layer6_outputs(3484));
    outputs(7139) <= not(layer6_outputs(4314));
    outputs(7140) <= (layer6_outputs(4716)) xor (layer6_outputs(6074));
    outputs(7141) <= not(layer6_outputs(260));
    outputs(7142) <= not(layer6_outputs(5843));
    outputs(7143) <= not(layer6_outputs(6288));
    outputs(7144) <= layer6_outputs(599);
    outputs(7145) <= layer6_outputs(2199);
    outputs(7146) <= (layer6_outputs(7428)) xor (layer6_outputs(5093));
    outputs(7147) <= not((layer6_outputs(3516)) xor (layer6_outputs(5068)));
    outputs(7148) <= not((layer6_outputs(6011)) xor (layer6_outputs(468)));
    outputs(7149) <= not((layer6_outputs(6000)) xor (layer6_outputs(5336)));
    outputs(7150) <= layer6_outputs(1046);
    outputs(7151) <= not((layer6_outputs(502)) xor (layer6_outputs(3644)));
    outputs(7152) <= layer6_outputs(6542);
    outputs(7153) <= layer6_outputs(5059);
    outputs(7154) <= not((layer6_outputs(5831)) xor (layer6_outputs(5212)));
    outputs(7155) <= (layer6_outputs(508)) xor (layer6_outputs(2008));
    outputs(7156) <= not(layer6_outputs(7650));
    outputs(7157) <= layer6_outputs(1840);
    outputs(7158) <= layer6_outputs(4826);
    outputs(7159) <= layer6_outputs(7012);
    outputs(7160) <= (layer6_outputs(123)) and not (layer6_outputs(4070));
    outputs(7161) <= layer6_outputs(7430);
    outputs(7162) <= layer6_outputs(4188);
    outputs(7163) <= not(layer6_outputs(5780));
    outputs(7164) <= layer6_outputs(2022);
    outputs(7165) <= layer6_outputs(2502);
    outputs(7166) <= not((layer6_outputs(1115)) or (layer6_outputs(757)));
    outputs(7167) <= not(layer6_outputs(188));
    outputs(7168) <= (layer6_outputs(1250)) and not (layer6_outputs(3249));
    outputs(7169) <= (layer6_outputs(2421)) xor (layer6_outputs(4273));
    outputs(7170) <= not(layer6_outputs(7101));
    outputs(7171) <= (layer6_outputs(742)) xor (layer6_outputs(7510));
    outputs(7172) <= not(layer6_outputs(3699));
    outputs(7173) <= not(layer6_outputs(540));
    outputs(7174) <= layer6_outputs(3554);
    outputs(7175) <= not(layer6_outputs(5629)) or (layer6_outputs(1633));
    outputs(7176) <= layer6_outputs(5390);
    outputs(7177) <= not(layer6_outputs(398));
    outputs(7178) <= (layer6_outputs(221)) or (layer6_outputs(4523));
    outputs(7179) <= not(layer6_outputs(1354)) or (layer6_outputs(6364));
    outputs(7180) <= not(layer6_outputs(1418)) or (layer6_outputs(1221));
    outputs(7181) <= layer6_outputs(7075);
    outputs(7182) <= layer6_outputs(2159);
    outputs(7183) <= layer6_outputs(6373);
    outputs(7184) <= layer6_outputs(7035);
    outputs(7185) <= layer6_outputs(3554);
    outputs(7186) <= not(layer6_outputs(92));
    outputs(7187) <= not((layer6_outputs(3279)) xor (layer6_outputs(7560)));
    outputs(7188) <= (layer6_outputs(4028)) and not (layer6_outputs(3502));
    outputs(7189) <= (layer6_outputs(2712)) or (layer6_outputs(581));
    outputs(7190) <= not(layer6_outputs(1798));
    outputs(7191) <= not((layer6_outputs(2854)) xor (layer6_outputs(6706)));
    outputs(7192) <= not((layer6_outputs(6987)) xor (layer6_outputs(6031)));
    outputs(7193) <= layer6_outputs(75);
    outputs(7194) <= not((layer6_outputs(3979)) xor (layer6_outputs(7118)));
    outputs(7195) <= not(layer6_outputs(6094)) or (layer6_outputs(4881));
    outputs(7196) <= not(layer6_outputs(5453));
    outputs(7197) <= (layer6_outputs(343)) and not (layer6_outputs(5714));
    outputs(7198) <= layer6_outputs(4697);
    outputs(7199) <= not((layer6_outputs(1167)) xor (layer6_outputs(5913)));
    outputs(7200) <= layer6_outputs(7570);
    outputs(7201) <= layer6_outputs(6656);
    outputs(7202) <= layer6_outputs(162);
    outputs(7203) <= not(layer6_outputs(5652));
    outputs(7204) <= (layer6_outputs(2301)) or (layer6_outputs(2157));
    outputs(7205) <= not(layer6_outputs(1378));
    outputs(7206) <= layer6_outputs(2099);
    outputs(7207) <= not((layer6_outputs(3237)) xor (layer6_outputs(765)));
    outputs(7208) <= (layer6_outputs(4575)) xor (layer6_outputs(4054));
    outputs(7209) <= (layer6_outputs(2075)) xor (layer6_outputs(2424));
    outputs(7210) <= not(layer6_outputs(6742));
    outputs(7211) <= layer6_outputs(7440);
    outputs(7212) <= (layer6_outputs(6765)) or (layer6_outputs(2848));
    outputs(7213) <= not((layer6_outputs(2746)) xor (layer6_outputs(5614)));
    outputs(7214) <= layer6_outputs(3181);
    outputs(7215) <= layer6_outputs(3841);
    outputs(7216) <= not(layer6_outputs(4923));
    outputs(7217) <= not((layer6_outputs(620)) xor (layer6_outputs(5298)));
    outputs(7218) <= (layer6_outputs(2808)) or (layer6_outputs(3429));
    outputs(7219) <= (layer6_outputs(7263)) xor (layer6_outputs(6874));
    outputs(7220) <= layer6_outputs(4575);
    outputs(7221) <= layer6_outputs(3734);
    outputs(7222) <= layer6_outputs(3640);
    outputs(7223) <= layer6_outputs(6159);
    outputs(7224) <= (layer6_outputs(2679)) xor (layer6_outputs(2232));
    outputs(7225) <= layer6_outputs(102);
    outputs(7226) <= layer6_outputs(7399);
    outputs(7227) <= not(layer6_outputs(1962));
    outputs(7228) <= layer6_outputs(4237);
    outputs(7229) <= layer6_outputs(2996);
    outputs(7230) <= not(layer6_outputs(4120));
    outputs(7231) <= not(layer6_outputs(5373));
    outputs(7232) <= (layer6_outputs(1531)) and (layer6_outputs(989));
    outputs(7233) <= not(layer6_outputs(6338));
    outputs(7234) <= not((layer6_outputs(3508)) and (layer6_outputs(4265)));
    outputs(7235) <= layer6_outputs(5891);
    outputs(7236) <= (layer6_outputs(2039)) xor (layer6_outputs(2641));
    outputs(7237) <= not((layer6_outputs(1428)) xor (layer6_outputs(1477)));
    outputs(7238) <= not(layer6_outputs(3724)) or (layer6_outputs(1019));
    outputs(7239) <= not(layer6_outputs(972));
    outputs(7240) <= (layer6_outputs(7095)) and not (layer6_outputs(1844));
    outputs(7241) <= not(layer6_outputs(6737)) or (layer6_outputs(1865));
    outputs(7242) <= not((layer6_outputs(3178)) or (layer6_outputs(4701)));
    outputs(7243) <= not((layer6_outputs(6323)) xor (layer6_outputs(5236)));
    outputs(7244) <= not((layer6_outputs(5005)) xor (layer6_outputs(4392)));
    outputs(7245) <= not(layer6_outputs(3326));
    outputs(7246) <= not((layer6_outputs(979)) xor (layer6_outputs(6719)));
    outputs(7247) <= layer6_outputs(209);
    outputs(7248) <= (layer6_outputs(1116)) xor (layer6_outputs(1435));
    outputs(7249) <= layer6_outputs(4650);
    outputs(7250) <= not(layer6_outputs(7482));
    outputs(7251) <= (layer6_outputs(7334)) xor (layer6_outputs(6850));
    outputs(7252) <= not((layer6_outputs(5018)) xor (layer6_outputs(4510)));
    outputs(7253) <= (layer6_outputs(4845)) xor (layer6_outputs(3200));
    outputs(7254) <= layer6_outputs(6805);
    outputs(7255) <= layer6_outputs(5865);
    outputs(7256) <= not(layer6_outputs(2158));
    outputs(7257) <= layer6_outputs(4571);
    outputs(7258) <= not((layer6_outputs(537)) xor (layer6_outputs(1312)));
    outputs(7259) <= (layer6_outputs(484)) xor (layer6_outputs(3893));
    outputs(7260) <= (layer6_outputs(7374)) and (layer6_outputs(6212));
    outputs(7261) <= not(layer6_outputs(465)) or (layer6_outputs(5303));
    outputs(7262) <= layer6_outputs(7136);
    outputs(7263) <= not(layer6_outputs(2395)) or (layer6_outputs(5277));
    outputs(7264) <= not(layer6_outputs(297)) or (layer6_outputs(888));
    outputs(7265) <= not((layer6_outputs(6147)) xor (layer6_outputs(3726)));
    outputs(7266) <= not(layer6_outputs(2812));
    outputs(7267) <= not(layer6_outputs(2225));
    outputs(7268) <= (layer6_outputs(7089)) and not (layer6_outputs(5858));
    outputs(7269) <= layer6_outputs(4604);
    outputs(7270) <= not(layer6_outputs(4763));
    outputs(7271) <= (layer6_outputs(4634)) xor (layer6_outputs(3004));
    outputs(7272) <= not(layer6_outputs(1714));
    outputs(7273) <= (layer6_outputs(3539)) xor (layer6_outputs(2491));
    outputs(7274) <= not(layer6_outputs(5159));
    outputs(7275) <= not(layer6_outputs(531));
    outputs(7276) <= not(layer6_outputs(859));
    outputs(7277) <= not(layer6_outputs(7165));
    outputs(7278) <= not(layer6_outputs(310));
    outputs(7279) <= layer6_outputs(5608);
    outputs(7280) <= not(layer6_outputs(2304));
    outputs(7281) <= (layer6_outputs(7327)) xor (layer6_outputs(1777));
    outputs(7282) <= layer6_outputs(875);
    outputs(7283) <= layer6_outputs(3812);
    outputs(7284) <= layer6_outputs(5953);
    outputs(7285) <= (layer6_outputs(1095)) xor (layer6_outputs(6367));
    outputs(7286) <= not(layer6_outputs(6812));
    outputs(7287) <= not((layer6_outputs(3345)) xor (layer6_outputs(1200)));
    outputs(7288) <= layer6_outputs(3841);
    outputs(7289) <= not(layer6_outputs(1870));
    outputs(7290) <= not(layer6_outputs(2991));
    outputs(7291) <= layer6_outputs(3513);
    outputs(7292) <= (layer6_outputs(4944)) and not (layer6_outputs(5507));
    outputs(7293) <= not(layer6_outputs(3404));
    outputs(7294) <= (layer6_outputs(143)) xor (layer6_outputs(5628));
    outputs(7295) <= layer6_outputs(1123);
    outputs(7296) <= layer6_outputs(4568);
    outputs(7297) <= not(layer6_outputs(1416));
    outputs(7298) <= (layer6_outputs(3810)) xor (layer6_outputs(176));
    outputs(7299) <= not((layer6_outputs(1648)) xor (layer6_outputs(637)));
    outputs(7300) <= layer6_outputs(6468);
    outputs(7301) <= (layer6_outputs(7355)) xor (layer6_outputs(2761));
    outputs(7302) <= not((layer6_outputs(3940)) or (layer6_outputs(1171)));
    outputs(7303) <= not(layer6_outputs(2593));
    outputs(7304) <= not(layer6_outputs(2771));
    outputs(7305) <= layer6_outputs(955);
    outputs(7306) <= not(layer6_outputs(2317)) or (layer6_outputs(851));
    outputs(7307) <= not((layer6_outputs(964)) xor (layer6_outputs(2507)));
    outputs(7308) <= (layer6_outputs(7508)) and not (layer6_outputs(1640));
    outputs(7309) <= (layer6_outputs(5794)) xor (layer6_outputs(2057));
    outputs(7310) <= not(layer6_outputs(1490));
    outputs(7311) <= layer6_outputs(1358);
    outputs(7312) <= layer6_outputs(793);
    outputs(7313) <= layer6_outputs(1608);
    outputs(7314) <= not(layer6_outputs(7056));
    outputs(7315) <= not(layer6_outputs(5597));
    outputs(7316) <= layer6_outputs(2908);
    outputs(7317) <= layer6_outputs(6057);
    outputs(7318) <= not(layer6_outputs(3373));
    outputs(7319) <= not(layer6_outputs(5392));
    outputs(7320) <= (layer6_outputs(5271)) and (layer6_outputs(3816));
    outputs(7321) <= layer6_outputs(5155);
    outputs(7322) <= (layer6_outputs(4634)) and not (layer6_outputs(6034));
    outputs(7323) <= not(layer6_outputs(6278));
    outputs(7324) <= layer6_outputs(311);
    outputs(7325) <= not(layer6_outputs(1750));
    outputs(7326) <= layer6_outputs(6935);
    outputs(7327) <= (layer6_outputs(7563)) and not (layer6_outputs(686));
    outputs(7328) <= (layer6_outputs(6473)) and not (layer6_outputs(2607));
    outputs(7329) <= layer6_outputs(14);
    outputs(7330) <= layer6_outputs(3886);
    outputs(7331) <= (layer6_outputs(7152)) and not (layer6_outputs(4289));
    outputs(7332) <= not((layer6_outputs(1190)) xor (layer6_outputs(6238)));
    outputs(7333) <= (layer6_outputs(2587)) and (layer6_outputs(1111));
    outputs(7334) <= not(layer6_outputs(4583));
    outputs(7335) <= (layer6_outputs(7200)) xor (layer6_outputs(3381));
    outputs(7336) <= (layer6_outputs(1249)) xor (layer6_outputs(3022));
    outputs(7337) <= layer6_outputs(1763);
    outputs(7338) <= not(layer6_outputs(2126));
    outputs(7339) <= (layer6_outputs(5406)) or (layer6_outputs(5740));
    outputs(7340) <= not(layer6_outputs(2238));
    outputs(7341) <= not((layer6_outputs(3264)) or (layer6_outputs(3884)));
    outputs(7342) <= (layer6_outputs(3364)) and not (layer6_outputs(5799));
    outputs(7343) <= not(layer6_outputs(4503));
    outputs(7344) <= not((layer6_outputs(823)) or (layer6_outputs(6802)));
    outputs(7345) <= layer6_outputs(6378);
    outputs(7346) <= layer6_outputs(4919);
    outputs(7347) <= not((layer6_outputs(1165)) xor (layer6_outputs(7429)));
    outputs(7348) <= not((layer6_outputs(3968)) or (layer6_outputs(1381)));
    outputs(7349) <= layer6_outputs(3605);
    outputs(7350) <= not(layer6_outputs(6924));
    outputs(7351) <= layer6_outputs(3686);
    outputs(7352) <= (layer6_outputs(7156)) xor (layer6_outputs(778));
    outputs(7353) <= (layer6_outputs(5755)) or (layer6_outputs(4369));
    outputs(7354) <= (layer6_outputs(3524)) and not (layer6_outputs(5188));
    outputs(7355) <= layer6_outputs(1491);
    outputs(7356) <= (layer6_outputs(7184)) xor (layer6_outputs(948));
    outputs(7357) <= not(layer6_outputs(3304));
    outputs(7358) <= not(layer6_outputs(1016));
    outputs(7359) <= layer6_outputs(2558);
    outputs(7360) <= not((layer6_outputs(194)) xor (layer6_outputs(33)));
    outputs(7361) <= (layer6_outputs(5676)) xor (layer6_outputs(1616));
    outputs(7362) <= (layer6_outputs(6019)) and not (layer6_outputs(3941));
    outputs(7363) <= not(layer6_outputs(5697));
    outputs(7364) <= (layer6_outputs(2328)) xor (layer6_outputs(6951));
    outputs(7365) <= (layer6_outputs(4056)) xor (layer6_outputs(4740));
    outputs(7366) <= (layer6_outputs(6447)) and (layer6_outputs(1108));
    outputs(7367) <= layer6_outputs(1139);
    outputs(7368) <= layer6_outputs(5151);
    outputs(7369) <= layer6_outputs(2662);
    outputs(7370) <= not(layer6_outputs(2885));
    outputs(7371) <= layer6_outputs(1510);
    outputs(7372) <= not(layer6_outputs(6710)) or (layer6_outputs(7147));
    outputs(7373) <= (layer6_outputs(1043)) and not (layer6_outputs(7534));
    outputs(7374) <= not(layer6_outputs(3247));
    outputs(7375) <= (layer6_outputs(2263)) and not (layer6_outputs(814));
    outputs(7376) <= not((layer6_outputs(3696)) xor (layer6_outputs(6597)));
    outputs(7377) <= not((layer6_outputs(4254)) xor (layer6_outputs(153)));
    outputs(7378) <= not(layer6_outputs(6877));
    outputs(7379) <= layer6_outputs(6273);
    outputs(7380) <= not(layer6_outputs(7613));
    outputs(7381) <= layer6_outputs(3010);
    outputs(7382) <= not((layer6_outputs(5803)) xor (layer6_outputs(4799)));
    outputs(7383) <= not(layer6_outputs(7485));
    outputs(7384) <= layer6_outputs(5013);
    outputs(7385) <= not(layer6_outputs(3131));
    outputs(7386) <= not((layer6_outputs(7251)) xor (layer6_outputs(7320)));
    outputs(7387) <= (layer6_outputs(3264)) xor (layer6_outputs(1161));
    outputs(7388) <= layer6_outputs(1306);
    outputs(7389) <= (layer6_outputs(7497)) xor (layer6_outputs(4191));
    outputs(7390) <= (layer6_outputs(4108)) and (layer6_outputs(4370));
    outputs(7391) <= (layer6_outputs(4978)) xor (layer6_outputs(780));
    outputs(7392) <= not(layer6_outputs(6971));
    outputs(7393) <= layer6_outputs(2696);
    outputs(7394) <= not((layer6_outputs(5540)) or (layer6_outputs(896)));
    outputs(7395) <= layer6_outputs(6716);
    outputs(7396) <= not((layer6_outputs(3563)) or (layer6_outputs(1736)));
    outputs(7397) <= not(layer6_outputs(4748)) or (layer6_outputs(5460));
    outputs(7398) <= not(layer6_outputs(4745));
    outputs(7399) <= not((layer6_outputs(3831)) xor (layer6_outputs(2456)));
    outputs(7400) <= layer6_outputs(420);
    outputs(7401) <= not(layer6_outputs(1248));
    outputs(7402) <= not(layer6_outputs(5434));
    outputs(7403) <= not((layer6_outputs(7416)) xor (layer6_outputs(3445)));
    outputs(7404) <= layer6_outputs(2465);
    outputs(7405) <= not(layer6_outputs(5589));
    outputs(7406) <= not(layer6_outputs(2804));
    outputs(7407) <= not(layer6_outputs(1857)) or (layer6_outputs(1442));
    outputs(7408) <= layer6_outputs(5503);
    outputs(7409) <= not((layer6_outputs(3055)) or (layer6_outputs(1113)));
    outputs(7410) <= layer6_outputs(5621);
    outputs(7411) <= not((layer6_outputs(5092)) xor (layer6_outputs(6024)));
    outputs(7412) <= not(layer6_outputs(1990));
    outputs(7413) <= layer6_outputs(7511);
    outputs(7414) <= not(layer6_outputs(6367));
    outputs(7415) <= not(layer6_outputs(1257));
    outputs(7416) <= layer6_outputs(1004);
    outputs(7417) <= (layer6_outputs(2050)) or (layer6_outputs(4886));
    outputs(7418) <= layer6_outputs(100);
    outputs(7419) <= not(layer6_outputs(3173));
    outputs(7420) <= (layer6_outputs(500)) and (layer6_outputs(3184));
    outputs(7421) <= not(layer6_outputs(3530));
    outputs(7422) <= not((layer6_outputs(2236)) xor (layer6_outputs(2327)));
    outputs(7423) <= not(layer6_outputs(7325));
    outputs(7424) <= not((layer6_outputs(1928)) or (layer6_outputs(644)));
    outputs(7425) <= layer6_outputs(3298);
    outputs(7426) <= layer6_outputs(1122);
    outputs(7427) <= not((layer6_outputs(554)) and (layer6_outputs(5493)));
    outputs(7428) <= (layer6_outputs(2956)) xor (layer6_outputs(3375));
    outputs(7429) <= layer6_outputs(4249);
    outputs(7430) <= not((layer6_outputs(3274)) xor (layer6_outputs(4065)));
    outputs(7431) <= (layer6_outputs(3972)) and (layer6_outputs(3878));
    outputs(7432) <= layer6_outputs(2085);
    outputs(7433) <= (layer6_outputs(4288)) xor (layer6_outputs(53));
    outputs(7434) <= not(layer6_outputs(1625));
    outputs(7435) <= (layer6_outputs(881)) and (layer6_outputs(5030));
    outputs(7436) <= (layer6_outputs(2541)) xor (layer6_outputs(4046));
    outputs(7437) <= layer6_outputs(4862);
    outputs(7438) <= layer6_outputs(4119);
    outputs(7439) <= not(layer6_outputs(4194));
    outputs(7440) <= not(layer6_outputs(3778));
    outputs(7441) <= not(layer6_outputs(6648)) or (layer6_outputs(5740));
    outputs(7442) <= layer6_outputs(1949);
    outputs(7443) <= layer6_outputs(2235);
    outputs(7444) <= not(layer6_outputs(609));
    outputs(7445) <= layer6_outputs(6340);
    outputs(7446) <= layer6_outputs(7553);
    outputs(7447) <= (layer6_outputs(2577)) and (layer6_outputs(1589));
    outputs(7448) <= (layer6_outputs(5335)) and not (layer6_outputs(6382));
    outputs(7449) <= (layer6_outputs(6253)) xor (layer6_outputs(3670));
    outputs(7450) <= not((layer6_outputs(5774)) or (layer6_outputs(7217)));
    outputs(7451) <= not(layer6_outputs(3206));
    outputs(7452) <= layer6_outputs(3906);
    outputs(7453) <= layer6_outputs(7531);
    outputs(7454) <= layer6_outputs(5842);
    outputs(7455) <= layer6_outputs(6372);
    outputs(7456) <= layer6_outputs(3760);
    outputs(7457) <= not(layer6_outputs(943));
    outputs(7458) <= not(layer6_outputs(2718));
    outputs(7459) <= not((layer6_outputs(3219)) or (layer6_outputs(2555)));
    outputs(7460) <= layer6_outputs(6);
    outputs(7461) <= (layer6_outputs(1791)) xor (layer6_outputs(1585));
    outputs(7462) <= layer6_outputs(5570);
    outputs(7463) <= layer6_outputs(2166);
    outputs(7464) <= (layer6_outputs(6691)) and not (layer6_outputs(5726));
    outputs(7465) <= (layer6_outputs(2731)) and not (layer6_outputs(6929));
    outputs(7466) <= not(layer6_outputs(4735));
    outputs(7467) <= (layer6_outputs(5830)) and not (layer6_outputs(1703));
    outputs(7468) <= layer6_outputs(357);
    outputs(7469) <= layer6_outputs(4811);
    outputs(7470) <= (layer6_outputs(2295)) or (layer6_outputs(3024));
    outputs(7471) <= not(layer6_outputs(5306));
    outputs(7472) <= layer6_outputs(4287);
    outputs(7473) <= layer6_outputs(849);
    outputs(7474) <= (layer6_outputs(5863)) xor (layer6_outputs(4572));
    outputs(7475) <= (layer6_outputs(721)) and not (layer6_outputs(4228));
    outputs(7476) <= layer6_outputs(4152);
    outputs(7477) <= not(layer6_outputs(6857)) or (layer6_outputs(6748));
    outputs(7478) <= not(layer6_outputs(4609));
    outputs(7479) <= (layer6_outputs(4785)) or (layer6_outputs(1846));
    outputs(7480) <= layer6_outputs(3497);
    outputs(7481) <= not(layer6_outputs(848)) or (layer6_outputs(3114));
    outputs(7482) <= not((layer6_outputs(1300)) or (layer6_outputs(4070)));
    outputs(7483) <= not(layer6_outputs(4581)) or (layer6_outputs(4845));
    outputs(7484) <= (layer6_outputs(2884)) and (layer6_outputs(6197));
    outputs(7485) <= not((layer6_outputs(4488)) xor (layer6_outputs(2084)));
    outputs(7486) <= not(layer6_outputs(3131));
    outputs(7487) <= not((layer6_outputs(3416)) xor (layer6_outputs(7222)));
    outputs(7488) <= layer6_outputs(6160);
    outputs(7489) <= not((layer6_outputs(2133)) and (layer6_outputs(4393)));
    outputs(7490) <= not((layer6_outputs(3088)) and (layer6_outputs(6600)));
    outputs(7491) <= not(layer6_outputs(7394));
    outputs(7492) <= not(layer6_outputs(1285));
    outputs(7493) <= not(layer6_outputs(3806));
    outputs(7494) <= (layer6_outputs(526)) or (layer6_outputs(4216));
    outputs(7495) <= layer6_outputs(5753);
    outputs(7496) <= not(layer6_outputs(448));
    outputs(7497) <= (layer6_outputs(3311)) and not (layer6_outputs(2575));
    outputs(7498) <= not((layer6_outputs(1861)) xor (layer6_outputs(1025)));
    outputs(7499) <= (layer6_outputs(1026)) xor (layer6_outputs(748));
    outputs(7500) <= not(layer6_outputs(429));
    outputs(7501) <= (layer6_outputs(6538)) or (layer6_outputs(2099));
    outputs(7502) <= not((layer6_outputs(4766)) xor (layer6_outputs(348)));
    outputs(7503) <= not(layer6_outputs(6571));
    outputs(7504) <= layer6_outputs(6669);
    outputs(7505) <= not(layer6_outputs(5528));
    outputs(7506) <= not(layer6_outputs(5104)) or (layer6_outputs(7440));
    outputs(7507) <= not(layer6_outputs(3862));
    outputs(7508) <= not(layer6_outputs(5088)) or (layer6_outputs(2017));
    outputs(7509) <= not(layer6_outputs(6596));
    outputs(7510) <= layer6_outputs(2826);
    outputs(7511) <= layer6_outputs(1207);
    outputs(7512) <= not((layer6_outputs(1775)) xor (layer6_outputs(3897)));
    outputs(7513) <= layer6_outputs(4632);
    outputs(7514) <= (layer6_outputs(3716)) and not (layer6_outputs(3444));
    outputs(7515) <= not((layer6_outputs(328)) xor (layer6_outputs(5250)));
    outputs(7516) <= layer6_outputs(2389);
    outputs(7517) <= not(layer6_outputs(1241));
    outputs(7518) <= not(layer6_outputs(7552));
    outputs(7519) <= not(layer6_outputs(7536));
    outputs(7520) <= not(layer6_outputs(7381));
    outputs(7521) <= not(layer6_outputs(5528));
    outputs(7522) <= not((layer6_outputs(3842)) or (layer6_outputs(5587)));
    outputs(7523) <= layer6_outputs(6557);
    outputs(7524) <= not(layer6_outputs(4602));
    outputs(7525) <= layer6_outputs(106);
    outputs(7526) <= not(layer6_outputs(1036));
    outputs(7527) <= layer6_outputs(4800);
    outputs(7528) <= layer6_outputs(3231);
    outputs(7529) <= layer6_outputs(6588);
    outputs(7530) <= not(layer6_outputs(1217));
    outputs(7531) <= (layer6_outputs(7047)) xor (layer6_outputs(5675));
    outputs(7532) <= layer6_outputs(269);
    outputs(7533) <= (layer6_outputs(4241)) xor (layer6_outputs(5592));
    outputs(7534) <= layer6_outputs(6245);
    outputs(7535) <= layer6_outputs(7674);
    outputs(7536) <= not(layer6_outputs(2342));
    outputs(7537) <= (layer6_outputs(4333)) and not (layer6_outputs(5735));
    outputs(7538) <= layer6_outputs(4536);
    outputs(7539) <= not(layer6_outputs(4911));
    outputs(7540) <= layer6_outputs(4887);
    outputs(7541) <= not(layer6_outputs(5099));
    outputs(7542) <= layer6_outputs(2800);
    outputs(7543) <= layer6_outputs(2301);
    outputs(7544) <= not(layer6_outputs(2823)) or (layer6_outputs(150));
    outputs(7545) <= not(layer6_outputs(1826));
    outputs(7546) <= layer6_outputs(6411);
    outputs(7547) <= not((layer6_outputs(608)) xor (layer6_outputs(335)));
    outputs(7548) <= (layer6_outputs(6809)) and not (layer6_outputs(3657));
    outputs(7549) <= (layer6_outputs(6123)) xor (layer6_outputs(2904));
    outputs(7550) <= not(layer6_outputs(2572));
    outputs(7551) <= not(layer6_outputs(6302));
    outputs(7552) <= not(layer6_outputs(7057));
    outputs(7553) <= layer6_outputs(6121);
    outputs(7554) <= (layer6_outputs(16)) and not (layer6_outputs(3749));
    outputs(7555) <= (layer6_outputs(5630)) or (layer6_outputs(7585));
    outputs(7556) <= not(layer6_outputs(1275));
    outputs(7557) <= not(layer6_outputs(6457));
    outputs(7558) <= not(layer6_outputs(6459));
    outputs(7559) <= (layer6_outputs(2699)) and (layer6_outputs(6449));
    outputs(7560) <= layer6_outputs(4427);
    outputs(7561) <= not(layer6_outputs(4554));
    outputs(7562) <= layer6_outputs(4473);
    outputs(7563) <= (layer6_outputs(5498)) and (layer6_outputs(6083));
    outputs(7564) <= not((layer6_outputs(5934)) xor (layer6_outputs(6174)));
    outputs(7565) <= not(layer6_outputs(558));
    outputs(7566) <= not((layer6_outputs(3240)) xor (layer6_outputs(2321)));
    outputs(7567) <= layer6_outputs(5873);
    outputs(7568) <= not((layer6_outputs(2090)) xor (layer6_outputs(1414)));
    outputs(7569) <= not((layer6_outputs(4136)) xor (layer6_outputs(5117)));
    outputs(7570) <= not(layer6_outputs(7507));
    outputs(7571) <= layer6_outputs(5312);
    outputs(7572) <= not(layer6_outputs(3053));
    outputs(7573) <= not(layer6_outputs(3633));
    outputs(7574) <= not(layer6_outputs(2880));
    outputs(7575) <= not((layer6_outputs(7478)) xor (layer6_outputs(7163)));
    outputs(7576) <= not((layer6_outputs(3088)) xor (layer6_outputs(5221)));
    outputs(7577) <= not(layer6_outputs(145));
    outputs(7578) <= layer6_outputs(1647);
    outputs(7579) <= layer6_outputs(2722);
    outputs(7580) <= not(layer6_outputs(6919));
    outputs(7581) <= not(layer6_outputs(1545));
    outputs(7582) <= not(layer6_outputs(7171));
    outputs(7583) <= layer6_outputs(6696);
    outputs(7584) <= (layer6_outputs(1583)) xor (layer6_outputs(1131));
    outputs(7585) <= not((layer6_outputs(1329)) and (layer6_outputs(7384)));
    outputs(7586) <= not(layer6_outputs(919));
    outputs(7587) <= not((layer6_outputs(6394)) xor (layer6_outputs(7444)));
    outputs(7588) <= (layer6_outputs(1114)) and not (layer6_outputs(1994));
    outputs(7589) <= (layer6_outputs(1538)) xor (layer6_outputs(7025));
    outputs(7590) <= layer6_outputs(853);
    outputs(7591) <= not(layer6_outputs(3135));
    outputs(7592) <= not(layer6_outputs(4148));
    outputs(7593) <= layer6_outputs(481);
    outputs(7594) <= not(layer6_outputs(7625));
    outputs(7595) <= not(layer6_outputs(3511));
    outputs(7596) <= layer6_outputs(364);
    outputs(7597) <= (layer6_outputs(7277)) xor (layer6_outputs(6589));
    outputs(7598) <= (layer6_outputs(4940)) xor (layer6_outputs(5436));
    outputs(7599) <= (layer6_outputs(3907)) xor (layer6_outputs(4675));
    outputs(7600) <= layer6_outputs(2875);
    outputs(7601) <= layer6_outputs(3401);
    outputs(7602) <= (layer6_outputs(3436)) xor (layer6_outputs(1933));
    outputs(7603) <= not(layer6_outputs(510));
    outputs(7604) <= not((layer6_outputs(255)) xor (layer6_outputs(1806)));
    outputs(7605) <= not(layer6_outputs(1868));
    outputs(7606) <= (layer6_outputs(2361)) or (layer6_outputs(4633));
    outputs(7607) <= not(layer6_outputs(1829));
    outputs(7608) <= (layer6_outputs(6068)) xor (layer6_outputs(3757));
    outputs(7609) <= not(layer6_outputs(2611));
    outputs(7610) <= not((layer6_outputs(2250)) xor (layer6_outputs(3423)));
    outputs(7611) <= (layer6_outputs(2781)) xor (layer6_outputs(3709));
    outputs(7612) <= (layer6_outputs(7264)) and not (layer6_outputs(3697));
    outputs(7613) <= layer6_outputs(3110);
    outputs(7614) <= not(layer6_outputs(1734));
    outputs(7615) <= layer6_outputs(6675);
    outputs(7616) <= not(layer6_outputs(7454));
    outputs(7617) <= (layer6_outputs(3536)) xor (layer6_outputs(6241));
    outputs(7618) <= not(layer6_outputs(807));
    outputs(7619) <= layer6_outputs(14);
    outputs(7620) <= layer6_outputs(5775);
    outputs(7621) <= not(layer6_outputs(1035));
    outputs(7622) <= (layer6_outputs(3636)) xor (layer6_outputs(4778));
    outputs(7623) <= layer6_outputs(1019);
    outputs(7624) <= (layer6_outputs(5488)) xor (layer6_outputs(802));
    outputs(7625) <= not((layer6_outputs(6432)) xor (layer6_outputs(457)));
    outputs(7626) <= not(layer6_outputs(2293));
    outputs(7627) <= not(layer6_outputs(6365));
    outputs(7628) <= (layer6_outputs(7471)) and (layer6_outputs(3170));
    outputs(7629) <= not((layer6_outputs(4229)) xor (layer6_outputs(6881)));
    outputs(7630) <= not(layer6_outputs(6997));
    outputs(7631) <= layer6_outputs(3740);
    outputs(7632) <= not(layer6_outputs(730));
    outputs(7633) <= layer6_outputs(6018);
    outputs(7634) <= (layer6_outputs(2132)) and (layer6_outputs(81));
    outputs(7635) <= not(layer6_outputs(4836));
    outputs(7636) <= layer6_outputs(3086);
    outputs(7637) <= layer6_outputs(4345);
    outputs(7638) <= not(layer6_outputs(3914));
    outputs(7639) <= layer6_outputs(2931);
    outputs(7640) <= layer6_outputs(6293);
    outputs(7641) <= not(layer6_outputs(1017));
    outputs(7642) <= not((layer6_outputs(3388)) xor (layer6_outputs(2819)));
    outputs(7643) <= (layer6_outputs(2677)) and not (layer6_outputs(7336));
    outputs(7644) <= (layer6_outputs(7569)) xor (layer6_outputs(2708));
    outputs(7645) <= not((layer6_outputs(3704)) xor (layer6_outputs(5696)));
    outputs(7646) <= not((layer6_outputs(2336)) or (layer6_outputs(73)));
    outputs(7647) <= not(layer6_outputs(1676));
    outputs(7648) <= not((layer6_outputs(3709)) xor (layer6_outputs(6397)));
    outputs(7649) <= not(layer6_outputs(1425));
    outputs(7650) <= not(layer6_outputs(1423));
    outputs(7651) <= not(layer6_outputs(769));
    outputs(7652) <= layer6_outputs(1817);
    outputs(7653) <= layer6_outputs(6071);
    outputs(7654) <= (layer6_outputs(6343)) or (layer6_outputs(1371));
    outputs(7655) <= (layer6_outputs(5282)) xor (layer6_outputs(1556));
    outputs(7656) <= layer6_outputs(2855);
    outputs(7657) <= layer6_outputs(511);
    outputs(7658) <= not(layer6_outputs(5747));
    outputs(7659) <= layer6_outputs(568);
    outputs(7660) <= (layer6_outputs(6231)) or (layer6_outputs(4954));
    outputs(7661) <= not(layer6_outputs(4102));
    outputs(7662) <= layer6_outputs(4271);
    outputs(7663) <= layer6_outputs(1590);
    outputs(7664) <= (layer6_outputs(6376)) xor (layer6_outputs(2973));
    outputs(7665) <= (layer6_outputs(2323)) xor (layer6_outputs(3722));
    outputs(7666) <= layer6_outputs(5173);
    outputs(7667) <= not((layer6_outputs(958)) xor (layer6_outputs(3453)));
    outputs(7668) <= not(layer6_outputs(4110));
    outputs(7669) <= not((layer6_outputs(2910)) xor (layer6_outputs(3958)));
    outputs(7670) <= (layer6_outputs(5058)) xor (layer6_outputs(6015));
    outputs(7671) <= (layer6_outputs(3656)) xor (layer6_outputs(7561));
    outputs(7672) <= layer6_outputs(1344);
    outputs(7673) <= not((layer6_outputs(2087)) or (layer6_outputs(6593)));
    outputs(7674) <= not((layer6_outputs(1388)) xor (layer6_outputs(4377)));
    outputs(7675) <= not(layer6_outputs(3205));
    outputs(7676) <= not(layer6_outputs(1317));
    outputs(7677) <= not(layer6_outputs(5729));
    outputs(7678) <= layer6_outputs(6254);
    outputs(7679) <= layer6_outputs(497);

end Behavioral;
