library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs: in std_logic_vector(1023 downto 0);
        outputs: out std_logic_vector(9 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs: std_logic_vector(2559 downto 0);

begin
    layer0_outputs(0) <= a;
    layer0_outputs(1) <= b and not a;
    layer0_outputs(2) <= not (a xor b);
    layer0_outputs(3) <= a and not b;
    layer0_outputs(4) <= a xor b;
    layer0_outputs(5) <= not b;
    layer0_outputs(6) <= a or b;
    layer0_outputs(7) <= a or b;
    layer0_outputs(8) <= a;
    layer0_outputs(9) <= not a;
    layer0_outputs(10) <= b and not a;
    layer0_outputs(11) <= not (a or b);
    layer0_outputs(12) <= not a or b;
    layer0_outputs(13) <= a xor b;
    layer0_outputs(14) <= a xor b;
    layer0_outputs(15) <= a or b;
    layer0_outputs(16) <= not (a and b);
    layer0_outputs(17) <= b;
    layer0_outputs(18) <= a or b;
    layer0_outputs(19) <= b and not a;
    layer0_outputs(20) <= not (a xor b);
    layer0_outputs(21) <= b and not a;
    layer0_outputs(22) <= not a;
    layer0_outputs(23) <= a xor b;
    layer0_outputs(24) <= a and not b;
    layer0_outputs(25) <= not b or a;
    layer0_outputs(26) <= not b;
    layer0_outputs(27) <= not a or b;
    layer0_outputs(28) <= not b;
    layer0_outputs(29) <= a;
    layer0_outputs(30) <= not (a xor b);
    layer0_outputs(31) <= a or b;
    layer0_outputs(32) <= not b;
    layer0_outputs(33) <= not (a or b);
    layer0_outputs(34) <= b;
    layer0_outputs(35) <= 1'b1;
    layer0_outputs(36) <= a;
    layer0_outputs(37) <= a or b;
    layer0_outputs(38) <= not a or b;
    layer0_outputs(39) <= not b or a;
    layer0_outputs(40) <= not b;
    layer0_outputs(41) <= a and b;
    layer0_outputs(42) <= 1'b0;
    layer0_outputs(43) <= b and not a;
    layer0_outputs(44) <= not (a or b);
    layer0_outputs(45) <= not (a or b);
    layer0_outputs(46) <= not b or a;
    layer0_outputs(47) <= not (a or b);
    layer0_outputs(48) <= b;
    layer0_outputs(49) <= not b;
    layer0_outputs(50) <= a or b;
    layer0_outputs(51) <= not (a or b);
    layer0_outputs(52) <= a and b;
    layer0_outputs(53) <= not a;
    layer0_outputs(54) <= a;
    layer0_outputs(55) <= not a or b;
    layer0_outputs(56) <= a;
    layer0_outputs(57) <= not (a xor b);
    layer0_outputs(58) <= a or b;
    layer0_outputs(59) <= not (a and b);
    layer0_outputs(60) <= a or b;
    layer0_outputs(61) <= a and b;
    layer0_outputs(62) <= not (a or b);
    layer0_outputs(63) <= not (a or b);
    layer0_outputs(64) <= a or b;
    layer0_outputs(65) <= not a or b;
    layer0_outputs(66) <= a and not b;
    layer0_outputs(67) <= not a or b;
    layer0_outputs(68) <= not a;
    layer0_outputs(69) <= not b;
    layer0_outputs(70) <= a or b;
    layer0_outputs(71) <= not (a or b);
    layer0_outputs(72) <= not a or b;
    layer0_outputs(73) <= b and not a;
    layer0_outputs(74) <= a or b;
    layer0_outputs(75) <= not (a or b);
    layer0_outputs(76) <= a or b;
    layer0_outputs(77) <= not b or a;
    layer0_outputs(78) <= not (a or b);
    layer0_outputs(79) <= a or b;
    layer0_outputs(80) <= b and not a;
    layer0_outputs(81) <= not (a or b);
    layer0_outputs(82) <= not (a or b);
    layer0_outputs(83) <= not a or b;
    layer0_outputs(84) <= not (a xor b);
    layer0_outputs(85) <= not (a or b);
    layer0_outputs(86) <= a and not b;
    layer0_outputs(87) <= b;
    layer0_outputs(88) <= a xor b;
    layer0_outputs(89) <= not a;
    layer0_outputs(90) <= not (a or b);
    layer0_outputs(91) <= a or b;
    layer0_outputs(92) <= not (a xor b);
    layer0_outputs(93) <= a xor b;
    layer0_outputs(94) <= not (a xor b);
    layer0_outputs(95) <= not b;
    layer0_outputs(96) <= not (a xor b);
    layer0_outputs(97) <= 1'b0;
    layer0_outputs(98) <= a or b;
    layer0_outputs(99) <= not b or a;
    layer0_outputs(100) <= not (a or b);
    layer0_outputs(101) <= a and not b;
    layer0_outputs(102) <= not (a or b);
    layer0_outputs(103) <= b and not a;
    layer0_outputs(104) <= a and not b;
    layer0_outputs(105) <= not (a or b);
    layer0_outputs(106) <= not (a xor b);
    layer0_outputs(107) <= a and not b;
    layer0_outputs(108) <= not (a or b);
    layer0_outputs(109) <= not (a or b);
    layer0_outputs(110) <= a;
    layer0_outputs(111) <= not (a or b);
    layer0_outputs(112) <= 1'b1;
    layer0_outputs(113) <= not (a xor b);
    layer0_outputs(114) <= not (a xor b);
    layer0_outputs(115) <= not (a or b);
    layer0_outputs(116) <= b and not a;
    layer0_outputs(117) <= not b;
    layer0_outputs(118) <= a or b;
    layer0_outputs(119) <= b;
    layer0_outputs(120) <= not (a or b);
    layer0_outputs(121) <= b;
    layer0_outputs(122) <= a or b;
    layer0_outputs(123) <= not a or b;
    layer0_outputs(124) <= a or b;
    layer0_outputs(125) <= not a or b;
    layer0_outputs(126) <= not (a xor b);
    layer0_outputs(127) <= b and not a;
    layer0_outputs(128) <= a or b;
    layer0_outputs(129) <= not (a or b);
    layer0_outputs(130) <= not a;
    layer0_outputs(131) <= 1'b1;
    layer0_outputs(132) <= not b or a;
    layer0_outputs(133) <= not b;
    layer0_outputs(134) <= a;
    layer0_outputs(135) <= not (a or b);
    layer0_outputs(136) <= not b or a;
    layer0_outputs(137) <= not b;
    layer0_outputs(138) <= b and not a;
    layer0_outputs(139) <= not b or a;
    layer0_outputs(140) <= not (a xor b);
    layer0_outputs(141) <= not b or a;
    layer0_outputs(142) <= a or b;
    layer0_outputs(143) <= not (a or b);
    layer0_outputs(144) <= 1'b1;
    layer0_outputs(145) <= not b;
    layer0_outputs(146) <= a or b;
    layer0_outputs(147) <= a or b;
    layer0_outputs(148) <= a or b;
    layer0_outputs(149) <= a xor b;
    layer0_outputs(150) <= a xor b;
    layer0_outputs(151) <= not (a and b);
    layer0_outputs(152) <= a or b;
    layer0_outputs(153) <= b and not a;
    layer0_outputs(154) <= not a;
    layer0_outputs(155) <= b and not a;
    layer0_outputs(156) <= b;
    layer0_outputs(157) <= not a;
    layer0_outputs(158) <= not b or a;
    layer0_outputs(159) <= a xor b;
    layer0_outputs(160) <= not (a xor b);
    layer0_outputs(161) <= not b or a;
    layer0_outputs(162) <= not b;
    layer0_outputs(163) <= not b;
    layer0_outputs(164) <= not (a xor b);
    layer0_outputs(165) <= a xor b;
    layer0_outputs(166) <= a or b;
    layer0_outputs(167) <= b and not a;
    layer0_outputs(168) <= b;
    layer0_outputs(169) <= b;
    layer0_outputs(170) <= not (a or b);
    layer0_outputs(171) <= not a or b;
    layer0_outputs(172) <= not b;
    layer0_outputs(173) <= not a;
    layer0_outputs(174) <= a xor b;
    layer0_outputs(175) <= b;
    layer0_outputs(176) <= not (a xor b);
    layer0_outputs(177) <= a and not b;
    layer0_outputs(178) <= a;
    layer0_outputs(179) <= not (a or b);
    layer0_outputs(180) <= not (a or b);
    layer0_outputs(181) <= a or b;
    layer0_outputs(182) <= a or b;
    layer0_outputs(183) <= not (a or b);
    layer0_outputs(184) <= not (a or b);
    layer0_outputs(185) <= not a or b;
    layer0_outputs(186) <= a xor b;
    layer0_outputs(187) <= a or b;
    layer0_outputs(188) <= a and not b;
    layer0_outputs(189) <= not b or a;
    layer0_outputs(190) <= not a;
    layer0_outputs(191) <= not b or a;
    layer0_outputs(192) <= a or b;
    layer0_outputs(193) <= not a;
    layer0_outputs(194) <= b and not a;
    layer0_outputs(195) <= a;
    layer0_outputs(196) <= a or b;
    layer0_outputs(197) <= not b or a;
    layer0_outputs(198) <= not (a or b);
    layer0_outputs(199) <= not (a or b);
    layer0_outputs(200) <= not (a or b);
    layer0_outputs(201) <= a or b;
    layer0_outputs(202) <= not (a or b);
    layer0_outputs(203) <= a and not b;
    layer0_outputs(204) <= not b;
    layer0_outputs(205) <= a or b;
    layer0_outputs(206) <= not (a or b);
    layer0_outputs(207) <= a and not b;
    layer0_outputs(208) <= not (a or b);
    layer0_outputs(209) <= a or b;
    layer0_outputs(210) <= a or b;
    layer0_outputs(211) <= a or b;
    layer0_outputs(212) <= not b;
    layer0_outputs(213) <= not (a xor b);
    layer0_outputs(214) <= not b or a;
    layer0_outputs(215) <= a;
    layer0_outputs(216) <= a;
    layer0_outputs(217) <= not a or b;
    layer0_outputs(218) <= a or b;
    layer0_outputs(219) <= not a;
    layer0_outputs(220) <= not b;
    layer0_outputs(221) <= not a;
    layer0_outputs(222) <= a or b;
    layer0_outputs(223) <= a or b;
    layer0_outputs(224) <= not a or b;
    layer0_outputs(225) <= not b or a;
    layer0_outputs(226) <= not (a and b);
    layer0_outputs(227) <= a xor b;
    layer0_outputs(228) <= not (a xor b);
    layer0_outputs(229) <= not (a xor b);
    layer0_outputs(230) <= a or b;
    layer0_outputs(231) <= 1'b0;
    layer0_outputs(232) <= 1'b1;
    layer0_outputs(233) <= a;
    layer0_outputs(234) <= not (a or b);
    layer0_outputs(235) <= not (a or b);
    layer0_outputs(236) <= a or b;
    layer0_outputs(237) <= a and not b;
    layer0_outputs(238) <= b;
    layer0_outputs(239) <= not b or a;
    layer0_outputs(240) <= a or b;
    layer0_outputs(241) <= a or b;
    layer0_outputs(242) <= not (a or b);
    layer0_outputs(243) <= a or b;
    layer0_outputs(244) <= b and not a;
    layer0_outputs(245) <= a xor b;
    layer0_outputs(246) <= not a;
    layer0_outputs(247) <= not a;
    layer0_outputs(248) <= b;
    layer0_outputs(249) <= not b;
    layer0_outputs(250) <= not b;
    layer0_outputs(251) <= not b or a;
    layer0_outputs(252) <= a and b;
    layer0_outputs(253) <= not (a xor b);
    layer0_outputs(254) <= not (a or b);
    layer0_outputs(255) <= a or b;
    layer0_outputs(256) <= not (a or b);
    layer0_outputs(257) <= a xor b;
    layer0_outputs(258) <= a and b;
    layer0_outputs(259) <= not (a or b);
    layer0_outputs(260) <= b and not a;
    layer0_outputs(261) <= b and not a;
    layer0_outputs(262) <= a or b;
    layer0_outputs(263) <= a;
    layer0_outputs(264) <= not (a or b);
    layer0_outputs(265) <= not (a and b);
    layer0_outputs(266) <= not a or b;
    layer0_outputs(267) <= a xor b;
    layer0_outputs(268) <= a xor b;
    layer0_outputs(269) <= a or b;
    layer0_outputs(270) <= not a;
    layer0_outputs(271) <= a and b;
    layer0_outputs(272) <= not (a or b);
    layer0_outputs(273) <= b;
    layer0_outputs(274) <= a and not b;
    layer0_outputs(275) <= not (a xor b);
    layer0_outputs(276) <= b and not a;
    layer0_outputs(277) <= not (a or b);
    layer0_outputs(278) <= a and not b;
    layer0_outputs(279) <= not a;
    layer0_outputs(280) <= not a or b;
    layer0_outputs(281) <= not b;
    layer0_outputs(282) <= a or b;
    layer0_outputs(283) <= not (a or b);
    layer0_outputs(284) <= b and not a;
    layer0_outputs(285) <= a or b;
    layer0_outputs(286) <= a and not b;
    layer0_outputs(287) <= a and not b;
    layer0_outputs(288) <= a or b;
    layer0_outputs(289) <= b and not a;
    layer0_outputs(290) <= not b or a;
    layer0_outputs(291) <= not (a or b);
    layer0_outputs(292) <= not b or a;
    layer0_outputs(293) <= b and not a;
    layer0_outputs(294) <= a xor b;
    layer0_outputs(295) <= a;
    layer0_outputs(296) <= a xor b;
    layer0_outputs(297) <= not (a or b);
    layer0_outputs(298) <= b and not a;
    layer0_outputs(299) <= not b;
    layer0_outputs(300) <= b;
    layer0_outputs(301) <= not (a xor b);
    layer0_outputs(302) <= not a;
    layer0_outputs(303) <= not a or b;
    layer0_outputs(304) <= b and not a;
    layer0_outputs(305) <= 1'b0;
    layer0_outputs(306) <= a and b;
    layer0_outputs(307) <= 1'b0;
    layer0_outputs(308) <= not a or b;
    layer0_outputs(309) <= a or b;
    layer0_outputs(310) <= not a;
    layer0_outputs(311) <= not a;
    layer0_outputs(312) <= a or b;
    layer0_outputs(313) <= a or b;
    layer0_outputs(314) <= a xor b;
    layer0_outputs(315) <= b;
    layer0_outputs(316) <= a or b;
    layer0_outputs(317) <= not b or a;
    layer0_outputs(318) <= b;
    layer0_outputs(319) <= a xor b;
    layer0_outputs(320) <= b and not a;
    layer0_outputs(321) <= a or b;
    layer0_outputs(322) <= a and b;
    layer0_outputs(323) <= a and not b;
    layer0_outputs(324) <= not (a or b);
    layer0_outputs(325) <= not (a or b);
    layer0_outputs(326) <= not b or a;
    layer0_outputs(327) <= b;
    layer0_outputs(328) <= a or b;
    layer0_outputs(329) <= b and not a;
    layer0_outputs(330) <= b and not a;
    layer0_outputs(331) <= a or b;
    layer0_outputs(332) <= not b;
    layer0_outputs(333) <= not (a or b);
    layer0_outputs(334) <= not (a or b);
    layer0_outputs(335) <= a or b;
    layer0_outputs(336) <= not b or a;
    layer0_outputs(337) <= not (a xor b);
    layer0_outputs(338) <= not b;
    layer0_outputs(339) <= a;
    layer0_outputs(340) <= b;
    layer0_outputs(341) <= not a or b;
    layer0_outputs(342) <= not (a or b);
    layer0_outputs(343) <= not b or a;
    layer0_outputs(344) <= not a or b;
    layer0_outputs(345) <= not a;
    layer0_outputs(346) <= not (a xor b);
    layer0_outputs(347) <= not a or b;
    layer0_outputs(348) <= a or b;
    layer0_outputs(349) <= b and not a;
    layer0_outputs(350) <= a and b;
    layer0_outputs(351) <= not (a or b);
    layer0_outputs(352) <= not a;
    layer0_outputs(353) <= a or b;
    layer0_outputs(354) <= not a;
    layer0_outputs(355) <= not b;
    layer0_outputs(356) <= not b;
    layer0_outputs(357) <= a or b;
    layer0_outputs(358) <= a or b;
    layer0_outputs(359) <= a or b;
    layer0_outputs(360) <= not b;
    layer0_outputs(361) <= not a;
    layer0_outputs(362) <= not (a or b);
    layer0_outputs(363) <= 1'b0;
    layer0_outputs(364) <= not (a xor b);
    layer0_outputs(365) <= 1'b1;
    layer0_outputs(366) <= a and not b;
    layer0_outputs(367) <= not b;
    layer0_outputs(368) <= not a;
    layer0_outputs(369) <= b;
    layer0_outputs(370) <= not a;
    layer0_outputs(371) <= not (a and b);
    layer0_outputs(372) <= not a or b;
    layer0_outputs(373) <= a or b;
    layer0_outputs(374) <= a xor b;
    layer0_outputs(375) <= b and not a;
    layer0_outputs(376) <= a;
    layer0_outputs(377) <= not b;
    layer0_outputs(378) <= not (a or b);
    layer0_outputs(379) <= b;
    layer0_outputs(380) <= a and not b;
    layer0_outputs(381) <= a and not b;
    layer0_outputs(382) <= a or b;
    layer0_outputs(383) <= a or b;
    layer0_outputs(384) <= not a or b;
    layer0_outputs(385) <= not (a xor b);
    layer0_outputs(386) <= a or b;
    layer0_outputs(387) <= a or b;
    layer0_outputs(388) <= a and not b;
    layer0_outputs(389) <= a or b;
    layer0_outputs(390) <= a and b;
    layer0_outputs(391) <= not (a or b);
    layer0_outputs(392) <= not b;
    layer0_outputs(393) <= not (a or b);
    layer0_outputs(394) <= a;
    layer0_outputs(395) <= not a;
    layer0_outputs(396) <= not a;
    layer0_outputs(397) <= not b or a;
    layer0_outputs(398) <= not b;
    layer0_outputs(399) <= a or b;
    layer0_outputs(400) <= a;
    layer0_outputs(401) <= not (a or b);
    layer0_outputs(402) <= b and not a;
    layer0_outputs(403) <= not b;
    layer0_outputs(404) <= not (a or b);
    layer0_outputs(405) <= a or b;
    layer0_outputs(406) <= a or b;
    layer0_outputs(407) <= a xor b;
    layer0_outputs(408) <= a or b;
    layer0_outputs(409) <= a or b;
    layer0_outputs(410) <= a and not b;
    layer0_outputs(411) <= a or b;
    layer0_outputs(412) <= a and not b;
    layer0_outputs(413) <= not (a or b);
    layer0_outputs(414) <= not (a or b);
    layer0_outputs(415) <= a and not b;
    layer0_outputs(416) <= not (a or b);
    layer0_outputs(417) <= not (a or b);
    layer0_outputs(418) <= not (a xor b);
    layer0_outputs(419) <= not a or b;
    layer0_outputs(420) <= not (a or b);
    layer0_outputs(421) <= not a or b;
    layer0_outputs(422) <= a and not b;
    layer0_outputs(423) <= a or b;
    layer0_outputs(424) <= a and b;
    layer0_outputs(425) <= not a or b;
    layer0_outputs(426) <= not a;
    layer0_outputs(427) <= not a or b;
    layer0_outputs(428) <= not (a or b);
    layer0_outputs(429) <= not (a and b);
    layer0_outputs(430) <= a and not b;
    layer0_outputs(431) <= not b;
    layer0_outputs(432) <= not a;
    layer0_outputs(433) <= a or b;
    layer0_outputs(434) <= not (a or b);
    layer0_outputs(435) <= b;
    layer0_outputs(436) <= a and not b;
    layer0_outputs(437) <= not (a or b);
    layer0_outputs(438) <= not (a or b);
    layer0_outputs(439) <= not b or a;
    layer0_outputs(440) <= a or b;
    layer0_outputs(441) <= a and not b;
    layer0_outputs(442) <= not (a xor b);
    layer0_outputs(443) <= a xor b;
    layer0_outputs(444) <= not a;
    layer0_outputs(445) <= a or b;
    layer0_outputs(446) <= a and not b;
    layer0_outputs(447) <= not (a or b);
    layer0_outputs(448) <= a or b;
    layer0_outputs(449) <= not (a or b);
    layer0_outputs(450) <= 1'b1;
    layer0_outputs(451) <= not (a or b);
    layer0_outputs(452) <= b;
    layer0_outputs(453) <= not b or a;
    layer0_outputs(454) <= a or b;
    layer0_outputs(455) <= a or b;
    layer0_outputs(456) <= 1'b1;
    layer0_outputs(457) <= a or b;
    layer0_outputs(458) <= a or b;
    layer0_outputs(459) <= not b;
    layer0_outputs(460) <= not a or b;
    layer0_outputs(461) <= not a;
    layer0_outputs(462) <= not b or a;
    layer0_outputs(463) <= not b;
    layer0_outputs(464) <= not a;
    layer0_outputs(465) <= b;
    layer0_outputs(466) <= not a;
    layer0_outputs(467) <= not (a or b);
    layer0_outputs(468) <= b;
    layer0_outputs(469) <= not (a xor b);
    layer0_outputs(470) <= a;
    layer0_outputs(471) <= b and not a;
    layer0_outputs(472) <= b;
    layer0_outputs(473) <= not b or a;
    layer0_outputs(474) <= not (a or b);
    layer0_outputs(475) <= a or b;
    layer0_outputs(476) <= not b or a;
    layer0_outputs(477) <= not b;
    layer0_outputs(478) <= not (a or b);
    layer0_outputs(479) <= not b or a;
    layer0_outputs(480) <= b;
    layer0_outputs(481) <= 1'b1;
    layer0_outputs(482) <= not (a or b);
    layer0_outputs(483) <= not a;
    layer0_outputs(484) <= a and not b;
    layer0_outputs(485) <= not (a xor b);
    layer0_outputs(486) <= 1'b0;
    layer0_outputs(487) <= a or b;
    layer0_outputs(488) <= a and not b;
    layer0_outputs(489) <= b;
    layer0_outputs(490) <= a or b;
    layer0_outputs(491) <= not a;
    layer0_outputs(492) <= not (a xor b);
    layer0_outputs(493) <= not (a or b);
    layer0_outputs(494) <= not (a or b);
    layer0_outputs(495) <= not (a or b);
    layer0_outputs(496) <= b;
    layer0_outputs(497) <= not b;
    layer0_outputs(498) <= not (a xor b);
    layer0_outputs(499) <= not (a or b);
    layer0_outputs(500) <= not a;
    layer0_outputs(501) <= b;
    layer0_outputs(502) <= a;
    layer0_outputs(503) <= not (a xor b);
    layer0_outputs(504) <= a and not b;
    layer0_outputs(505) <= not b;
    layer0_outputs(506) <= not (a or b);
    layer0_outputs(507) <= 1'b1;
    layer0_outputs(508) <= 1'b0;
    layer0_outputs(509) <= a and not b;
    layer0_outputs(510) <= a or b;
    layer0_outputs(511) <= not b;
    layer0_outputs(512) <= not b;
    layer0_outputs(513) <= not a;
    layer0_outputs(514) <= b and not a;
    layer0_outputs(515) <= not (a or b);
    layer0_outputs(516) <= not a;
    layer0_outputs(517) <= not (a and b);
    layer0_outputs(518) <= not a or b;
    layer0_outputs(519) <= b and not a;
    layer0_outputs(520) <= a xor b;
    layer0_outputs(521) <= not b or a;
    layer0_outputs(522) <= a or b;
    layer0_outputs(523) <= not a or b;
    layer0_outputs(524) <= not a;
    layer0_outputs(525) <= a or b;
    layer0_outputs(526) <= not b;
    layer0_outputs(527) <= not (a or b);
    layer0_outputs(528) <= not (a or b);
    layer0_outputs(529) <= not (a or b);
    layer0_outputs(530) <= not (a xor b);
    layer0_outputs(531) <= a;
    layer0_outputs(532) <= a;
    layer0_outputs(533) <= not (a or b);
    layer0_outputs(534) <= b;
    layer0_outputs(535) <= a;
    layer0_outputs(536) <= a xor b;
    layer0_outputs(537) <= not b;
    layer0_outputs(538) <= a xor b;
    layer0_outputs(539) <= 1'b1;
    layer0_outputs(540) <= 1'b1;
    layer0_outputs(541) <= not (a or b);
    layer0_outputs(542) <= a or b;
    layer0_outputs(543) <= a or b;
    layer0_outputs(544) <= not b or a;
    layer0_outputs(545) <= not (a or b);
    layer0_outputs(546) <= b and not a;
    layer0_outputs(547) <= not a;
    layer0_outputs(548) <= not a;
    layer0_outputs(549) <= not b;
    layer0_outputs(550) <= not b or a;
    layer0_outputs(551) <= a;
    layer0_outputs(552) <= a or b;
    layer0_outputs(553) <= a xor b;
    layer0_outputs(554) <= a or b;
    layer0_outputs(555) <= not (a xor b);
    layer0_outputs(556) <= not b or a;
    layer0_outputs(557) <= b;
    layer0_outputs(558) <= not (a and b);
    layer0_outputs(559) <= not (a or b);
    layer0_outputs(560) <= not b or a;
    layer0_outputs(561) <= not a or b;
    layer0_outputs(562) <= not b;
    layer0_outputs(563) <= b and not a;
    layer0_outputs(564) <= not b;
    layer0_outputs(565) <= b;
    layer0_outputs(566) <= a or b;
    layer0_outputs(567) <= b;
    layer0_outputs(568) <= a or b;
    layer0_outputs(569) <= a;
    layer0_outputs(570) <= not (a or b);
    layer0_outputs(571) <= not (a or b);
    layer0_outputs(572) <= a;
    layer0_outputs(573) <= not (a or b);
    layer0_outputs(574) <= b;
    layer0_outputs(575) <= not (a xor b);
    layer0_outputs(576) <= not a;
    layer0_outputs(577) <= a or b;
    layer0_outputs(578) <= not a;
    layer0_outputs(579) <= a and not b;
    layer0_outputs(580) <= not (a or b);
    layer0_outputs(581) <= b and not a;
    layer0_outputs(582) <= a and b;
    layer0_outputs(583) <= a xor b;
    layer0_outputs(584) <= b and not a;
    layer0_outputs(585) <= 1'b1;
    layer0_outputs(586) <= a or b;
    layer0_outputs(587) <= a xor b;
    layer0_outputs(588) <= not (a or b);
    layer0_outputs(589) <= a xor b;
    layer0_outputs(590) <= a or b;
    layer0_outputs(591) <= not a;
    layer0_outputs(592) <= a or b;
    layer0_outputs(593) <= b and not a;
    layer0_outputs(594) <= a xor b;
    layer0_outputs(595) <= not b;
    layer0_outputs(596) <= a or b;
    layer0_outputs(597) <= a or b;
    layer0_outputs(598) <= not b or a;
    layer0_outputs(599) <= a or b;
    layer0_outputs(600) <= not (a and b);
    layer0_outputs(601) <= not b;
    layer0_outputs(602) <= not b or a;
    layer0_outputs(603) <= not (a xor b);
    layer0_outputs(604) <= not (a xor b);
    layer0_outputs(605) <= not a or b;
    layer0_outputs(606) <= 1'b0;
    layer0_outputs(607) <= not b;
    layer0_outputs(608) <= b and not a;
    layer0_outputs(609) <= not (a xor b);
    layer0_outputs(610) <= not (a or b);
    layer0_outputs(611) <= a;
    layer0_outputs(612) <= a;
    layer0_outputs(613) <= b and not a;
    layer0_outputs(614) <= not (a xor b);
    layer0_outputs(615) <= not a;
    layer0_outputs(616) <= not a;
    layer0_outputs(617) <= not (a or b);
    layer0_outputs(618) <= not (a or b);
    layer0_outputs(619) <= 1'b1;
    layer0_outputs(620) <= a;
    layer0_outputs(621) <= a xor b;
    layer0_outputs(622) <= a or b;
    layer0_outputs(623) <= not (a or b);
    layer0_outputs(624) <= not b or a;
    layer0_outputs(625) <= a xor b;
    layer0_outputs(626) <= a or b;
    layer0_outputs(627) <= b and not a;
    layer0_outputs(628) <= not (a or b);
    layer0_outputs(629) <= b and not a;
    layer0_outputs(630) <= not (a or b);
    layer0_outputs(631) <= not b or a;
    layer0_outputs(632) <= not (a xor b);
    layer0_outputs(633) <= not a;
    layer0_outputs(634) <= not b or a;
    layer0_outputs(635) <= not b or a;
    layer0_outputs(636) <= a;
    layer0_outputs(637) <= b and not a;
    layer0_outputs(638) <= not (a or b);
    layer0_outputs(639) <= not a;
    layer0_outputs(640) <= not (a or b);
    layer0_outputs(641) <= b;
    layer0_outputs(642) <= a and not b;
    layer0_outputs(643) <= not b;
    layer0_outputs(644) <= not (a or b);
    layer0_outputs(645) <= not b or a;
    layer0_outputs(646) <= not (a or b);
    layer0_outputs(647) <= a and b;
    layer0_outputs(648) <= a xor b;
    layer0_outputs(649) <= not a or b;
    layer0_outputs(650) <= a xor b;
    layer0_outputs(651) <= not a;
    layer0_outputs(652) <= not a or b;
    layer0_outputs(653) <= b;
    layer0_outputs(654) <= a or b;
    layer0_outputs(655) <= not (a xor b);
    layer0_outputs(656) <= b;
    layer0_outputs(657) <= b and not a;
    layer0_outputs(658) <= a or b;
    layer0_outputs(659) <= not b;
    layer0_outputs(660) <= 1'b1;
    layer0_outputs(661) <= a;
    layer0_outputs(662) <= a;
    layer0_outputs(663) <= not b;
    layer0_outputs(664) <= a or b;
    layer0_outputs(665) <= not (a or b);
    layer0_outputs(666) <= b;
    layer0_outputs(667) <= a;
    layer0_outputs(668) <= not b or a;
    layer0_outputs(669) <= b and not a;
    layer0_outputs(670) <= not (a and b);
    layer0_outputs(671) <= not (a or b);
    layer0_outputs(672) <= a;
    layer0_outputs(673) <= not b;
    layer0_outputs(674) <= not b or a;
    layer0_outputs(675) <= a or b;
    layer0_outputs(676) <= 1'b1;
    layer0_outputs(677) <= 1'b0;
    layer0_outputs(678) <= not (a or b);
    layer0_outputs(679) <= a xor b;
    layer0_outputs(680) <= a;
    layer0_outputs(681) <= not a or b;
    layer0_outputs(682) <= a or b;
    layer0_outputs(683) <= a and not b;
    layer0_outputs(684) <= not b or a;
    layer0_outputs(685) <= not b or a;
    layer0_outputs(686) <= not a or b;
    layer0_outputs(687) <= not a;
    layer0_outputs(688) <= not a or b;
    layer0_outputs(689) <= b and not a;
    layer0_outputs(690) <= not (a xor b);
    layer0_outputs(691) <= not a or b;
    layer0_outputs(692) <= not (a or b);
    layer0_outputs(693) <= not (a xor b);
    layer0_outputs(694) <= not a;
    layer0_outputs(695) <= b;
    layer0_outputs(696) <= a and not b;
    layer0_outputs(697) <= a or b;
    layer0_outputs(698) <= not a or b;
    layer0_outputs(699) <= a and not b;
    layer0_outputs(700) <= not (a and b);
    layer0_outputs(701) <= not (a xor b);
    layer0_outputs(702) <= a or b;
    layer0_outputs(703) <= not a or b;
    layer0_outputs(704) <= a and not b;
    layer0_outputs(705) <= a or b;
    layer0_outputs(706) <= b;
    layer0_outputs(707) <= a or b;
    layer0_outputs(708) <= not (a and b);
    layer0_outputs(709) <= not a or b;
    layer0_outputs(710) <= not b;
    layer0_outputs(711) <= 1'b0;
    layer0_outputs(712) <= not b;
    layer0_outputs(713) <= b;
    layer0_outputs(714) <= not b or a;
    layer0_outputs(715) <= not (a or b);
    layer0_outputs(716) <= not a or b;
    layer0_outputs(717) <= b;
    layer0_outputs(718) <= b;
    layer0_outputs(719) <= not b;
    layer0_outputs(720) <= not a or b;
    layer0_outputs(721) <= not (a xor b);
    layer0_outputs(722) <= a and not b;
    layer0_outputs(723) <= b and not a;
    layer0_outputs(724) <= not a;
    layer0_outputs(725) <= not b;
    layer0_outputs(726) <= not (a or b);
    layer0_outputs(727) <= not (a or b);
    layer0_outputs(728) <= a xor b;
    layer0_outputs(729) <= not (a or b);
    layer0_outputs(730) <= b;
    layer0_outputs(731) <= a and not b;
    layer0_outputs(732) <= a;
    layer0_outputs(733) <= not (a xor b);
    layer0_outputs(734) <= not (a xor b);
    layer0_outputs(735) <= not a or b;
    layer0_outputs(736) <= a or b;
    layer0_outputs(737) <= not b or a;
    layer0_outputs(738) <= not b;
    layer0_outputs(739) <= not b;
    layer0_outputs(740) <= not (a xor b);
    layer0_outputs(741) <= a or b;
    layer0_outputs(742) <= a xor b;
    layer0_outputs(743) <= b;
    layer0_outputs(744) <= not b;
    layer0_outputs(745) <= a and not b;
    layer0_outputs(746) <= not (a xor b);
    layer0_outputs(747) <= not b;
    layer0_outputs(748) <= not (a or b);
    layer0_outputs(749) <= not a or b;
    layer0_outputs(750) <= not (a or b);
    layer0_outputs(751) <= not (a and b);
    layer0_outputs(752) <= not a;
    layer0_outputs(753) <= not a;
    layer0_outputs(754) <= not a or b;
    layer0_outputs(755) <= not b;
    layer0_outputs(756) <= not (a or b);
    layer0_outputs(757) <= not b or a;
    layer0_outputs(758) <= a xor b;
    layer0_outputs(759) <= not (a and b);
    layer0_outputs(760) <= a or b;
    layer0_outputs(761) <= a or b;
    layer0_outputs(762) <= b;
    layer0_outputs(763) <= not b;
    layer0_outputs(764) <= a;
    layer0_outputs(765) <= a xor b;
    layer0_outputs(766) <= not (a or b);
    layer0_outputs(767) <= not (a xor b);
    layer0_outputs(768) <= not (a or b);
    layer0_outputs(769) <= not b;
    layer0_outputs(770) <= not (a or b);
    layer0_outputs(771) <= not b;
    layer0_outputs(772) <= not (a xor b);
    layer0_outputs(773) <= b and not a;
    layer0_outputs(774) <= not (a xor b);
    layer0_outputs(775) <= not b;
    layer0_outputs(776) <= not a;
    layer0_outputs(777) <= a or b;
    layer0_outputs(778) <= not (a or b);
    layer0_outputs(779) <= b;
    layer0_outputs(780) <= a or b;
    layer0_outputs(781) <= 1'b0;
    layer0_outputs(782) <= b;
    layer0_outputs(783) <= b and not a;
    layer0_outputs(784) <= a;
    layer0_outputs(785) <= a or b;
    layer0_outputs(786) <= not b or a;
    layer0_outputs(787) <= a and not b;
    layer0_outputs(788) <= not (a or b);
    layer0_outputs(789) <= not (a xor b);
    layer0_outputs(790) <= not (a or b);
    layer0_outputs(791) <= not b or a;
    layer0_outputs(792) <= b;
    layer0_outputs(793) <= a or b;
    layer0_outputs(794) <= a xor b;
    layer0_outputs(795) <= not (a or b);
    layer0_outputs(796) <= not (a xor b);
    layer0_outputs(797) <= not b;
    layer0_outputs(798) <= not (a xor b);
    layer0_outputs(799) <= a or b;
    layer0_outputs(800) <= not (a or b);
    layer0_outputs(801) <= a;
    layer0_outputs(802) <= a and not b;
    layer0_outputs(803) <= 1'b0;
    layer0_outputs(804) <= a xor b;
    layer0_outputs(805) <= not (a or b);
    layer0_outputs(806) <= not b;
    layer0_outputs(807) <= not (a xor b);
    layer0_outputs(808) <= not (a or b);
    layer0_outputs(809) <= a or b;
    layer0_outputs(810) <= 1'b0;
    layer0_outputs(811) <= not b;
    layer0_outputs(812) <= b and not a;
    layer0_outputs(813) <= not a;
    layer0_outputs(814) <= b;
    layer0_outputs(815) <= not (a xor b);
    layer0_outputs(816) <= not a;
    layer0_outputs(817) <= b;
    layer0_outputs(818) <= not (a xor b);
    layer0_outputs(819) <= not (a or b);
    layer0_outputs(820) <= not a or b;
    layer0_outputs(821) <= not (a xor b);
    layer0_outputs(822) <= not a or b;
    layer0_outputs(823) <= a;
    layer0_outputs(824) <= not a or b;
    layer0_outputs(825) <= a xor b;
    layer0_outputs(826) <= not (a or b);
    layer0_outputs(827) <= a or b;
    layer0_outputs(828) <= not a;
    layer0_outputs(829) <= a and b;
    layer0_outputs(830) <= not a;
    layer0_outputs(831) <= not (a or b);
    layer0_outputs(832) <= not (a or b);
    layer0_outputs(833) <= not (a or b);
    layer0_outputs(834) <= b;
    layer0_outputs(835) <= a xor b;
    layer0_outputs(836) <= b and not a;
    layer0_outputs(837) <= not (a or b);
    layer0_outputs(838) <= a xor b;
    layer0_outputs(839) <= not (a xor b);
    layer0_outputs(840) <= not (a or b);
    layer0_outputs(841) <= b;
    layer0_outputs(842) <= a or b;
    layer0_outputs(843) <= not (a or b);
    layer0_outputs(844) <= a and not b;
    layer0_outputs(845) <= not a;
    layer0_outputs(846) <= a and not b;
    layer0_outputs(847) <= a;
    layer0_outputs(848) <= b;
    layer0_outputs(849) <= a xor b;
    layer0_outputs(850) <= not (a or b);
    layer0_outputs(851) <= a and not b;
    layer0_outputs(852) <= not (a xor b);
    layer0_outputs(853) <= not a or b;
    layer0_outputs(854) <= a xor b;
    layer0_outputs(855) <= not a or b;
    layer0_outputs(856) <= not (a or b);
    layer0_outputs(857) <= not (a or b);
    layer0_outputs(858) <= b and not a;
    layer0_outputs(859) <= a or b;
    layer0_outputs(860) <= not a;
    layer0_outputs(861) <= not a;
    layer0_outputs(862) <= not b;
    layer0_outputs(863) <= a or b;
    layer0_outputs(864) <= a or b;
    layer0_outputs(865) <= a xor b;
    layer0_outputs(866) <= a xor b;
    layer0_outputs(867) <= a xor b;
    layer0_outputs(868) <= not (a or b);
    layer0_outputs(869) <= b and not a;
    layer0_outputs(870) <= a;
    layer0_outputs(871) <= not b;
    layer0_outputs(872) <= a or b;
    layer0_outputs(873) <= not (a or b);
    layer0_outputs(874) <= not b;
    layer0_outputs(875) <= a and b;
    layer0_outputs(876) <= a;
    layer0_outputs(877) <= a or b;
    layer0_outputs(878) <= a or b;
    layer0_outputs(879) <= not (a xor b);
    layer0_outputs(880) <= not (a or b);
    layer0_outputs(881) <= not b;
    layer0_outputs(882) <= a or b;
    layer0_outputs(883) <= not (a or b);
    layer0_outputs(884) <= not (a or b);
    layer0_outputs(885) <= not a or b;
    layer0_outputs(886) <= not a or b;
    layer0_outputs(887) <= a or b;
    layer0_outputs(888) <= b and not a;
    layer0_outputs(889) <= 1'b1;
    layer0_outputs(890) <= not (a or b);
    layer0_outputs(891) <= not a or b;
    layer0_outputs(892) <= a xor b;
    layer0_outputs(893) <= not b;
    layer0_outputs(894) <= not (a xor b);
    layer0_outputs(895) <= b;
    layer0_outputs(896) <= not (a or b);
    layer0_outputs(897) <= a xor b;
    layer0_outputs(898) <= not a;
    layer0_outputs(899) <= a;
    layer0_outputs(900) <= 1'b0;
    layer0_outputs(901) <= not (a and b);
    layer0_outputs(902) <= a;
    layer0_outputs(903) <= a or b;
    layer0_outputs(904) <= 1'b1;
    layer0_outputs(905) <= a or b;
    layer0_outputs(906) <= a or b;
    layer0_outputs(907) <= not (a or b);
    layer0_outputs(908) <= a and not b;
    layer0_outputs(909) <= a or b;
    layer0_outputs(910) <= a or b;
    layer0_outputs(911) <= a or b;
    layer0_outputs(912) <= a and not b;
    layer0_outputs(913) <= a or b;
    layer0_outputs(914) <= a or b;
    layer0_outputs(915) <= a or b;
    layer0_outputs(916) <= not a;
    layer0_outputs(917) <= not a or b;
    layer0_outputs(918) <= not a;
    layer0_outputs(919) <= a;
    layer0_outputs(920) <= a xor b;
    layer0_outputs(921) <= not a or b;
    layer0_outputs(922) <= a or b;
    layer0_outputs(923) <= not b;
    layer0_outputs(924) <= not (a or b);
    layer0_outputs(925) <= a xor b;
    layer0_outputs(926) <= a or b;
    layer0_outputs(927) <= b;
    layer0_outputs(928) <= b and not a;
    layer0_outputs(929) <= not (a or b);
    layer0_outputs(930) <= a or b;
    layer0_outputs(931) <= not b or a;
    layer0_outputs(932) <= not a or b;
    layer0_outputs(933) <= a or b;
    layer0_outputs(934) <= not b;
    layer0_outputs(935) <= not (a xor b);
    layer0_outputs(936) <= not b;
    layer0_outputs(937) <= a and not b;
    layer0_outputs(938) <= a or b;
    layer0_outputs(939) <= a and b;
    layer0_outputs(940) <= not a;
    layer0_outputs(941) <= a and not b;
    layer0_outputs(942) <= not a or b;
    layer0_outputs(943) <= a and not b;
    layer0_outputs(944) <= 1'b1;
    layer0_outputs(945) <= a and not b;
    layer0_outputs(946) <= b;
    layer0_outputs(947) <= not (a xor b);
    layer0_outputs(948) <= 1'b0;
    layer0_outputs(949) <= a xor b;
    layer0_outputs(950) <= b;
    layer0_outputs(951) <= not (a xor b);
    layer0_outputs(952) <= a and b;
    layer0_outputs(953) <= not b;
    layer0_outputs(954) <= b;
    layer0_outputs(955) <= not b;
    layer0_outputs(956) <= a or b;
    layer0_outputs(957) <= a and not b;
    layer0_outputs(958) <= not b or a;
    layer0_outputs(959) <= a or b;
    layer0_outputs(960) <= not b or a;
    layer0_outputs(961) <= 1'b1;
    layer0_outputs(962) <= not (a or b);
    layer0_outputs(963) <= not a or b;
    layer0_outputs(964) <= 1'b0;
    layer0_outputs(965) <= not a or b;
    layer0_outputs(966) <= not (a or b);
    layer0_outputs(967) <= a;
    layer0_outputs(968) <= not (a or b);
    layer0_outputs(969) <= a and not b;
    layer0_outputs(970) <= not (a or b);
    layer0_outputs(971) <= not (a or b);
    layer0_outputs(972) <= a and not b;
    layer0_outputs(973) <= a or b;
    layer0_outputs(974) <= not (a or b);
    layer0_outputs(975) <= not b or a;
    layer0_outputs(976) <= not (a or b);
    layer0_outputs(977) <= not (a xor b);
    layer0_outputs(978) <= b and not a;
    layer0_outputs(979) <= b;
    layer0_outputs(980) <= a;
    layer0_outputs(981) <= not b;
    layer0_outputs(982) <= not (a or b);
    layer0_outputs(983) <= not a;
    layer0_outputs(984) <= not (a or b);
    layer0_outputs(985) <= b;
    layer0_outputs(986) <= a or b;
    layer0_outputs(987) <= not b;
    layer0_outputs(988) <= a;
    layer0_outputs(989) <= not (a or b);
    layer0_outputs(990) <= a or b;
    layer0_outputs(991) <= not (a or b);
    layer0_outputs(992) <= b and not a;
    layer0_outputs(993) <= b;
    layer0_outputs(994) <= not b;
    layer0_outputs(995) <= not (a xor b);
    layer0_outputs(996) <= not (a xor b);
    layer0_outputs(997) <= not (a xor b);
    layer0_outputs(998) <= a;
    layer0_outputs(999) <= b;
    layer0_outputs(1000) <= not (a xor b);
    layer0_outputs(1001) <= a and not b;
    layer0_outputs(1002) <= not a;
    layer0_outputs(1003) <= not (a or b);
    layer0_outputs(1004) <= 1'b0;
    layer0_outputs(1005) <= b;
    layer0_outputs(1006) <= not (a xor b);
    layer0_outputs(1007) <= a and not b;
    layer0_outputs(1008) <= not (a or b);
    layer0_outputs(1009) <= not b;
    layer0_outputs(1010) <= b and not a;
    layer0_outputs(1011) <= a or b;
    layer0_outputs(1012) <= b;
    layer0_outputs(1013) <= not (a or b);
    layer0_outputs(1014) <= b and not a;
    layer0_outputs(1015) <= a and not b;
    layer0_outputs(1016) <= not b or a;
    layer0_outputs(1017) <= not (a xor b);
    layer0_outputs(1018) <= not b or a;
    layer0_outputs(1019) <= not a;
    layer0_outputs(1020) <= a and not b;
    layer0_outputs(1021) <= a or b;
    layer0_outputs(1022) <= a or b;
    layer0_outputs(1023) <= not b or a;
    layer0_outputs(1024) <= a;
    layer0_outputs(1025) <= a xor b;
    layer0_outputs(1026) <= not (a or b);
    layer0_outputs(1027) <= not (a or b);
    layer0_outputs(1028) <= not (a or b);
    layer0_outputs(1029) <= a and not b;
    layer0_outputs(1030) <= not b;
    layer0_outputs(1031) <= 1'b1;
    layer0_outputs(1032) <= not b or a;
    layer0_outputs(1033) <= not b;
    layer0_outputs(1034) <= not (a or b);
    layer0_outputs(1035) <= a or b;
    layer0_outputs(1036) <= a xor b;
    layer0_outputs(1037) <= not b;
    layer0_outputs(1038) <= not b or a;
    layer0_outputs(1039) <= a or b;
    layer0_outputs(1040) <= not b;
    layer0_outputs(1041) <= b;
    layer0_outputs(1042) <= not a or b;
    layer0_outputs(1043) <= b and not a;
    layer0_outputs(1044) <= not a or b;
    layer0_outputs(1045) <= not a;
    layer0_outputs(1046) <= a and not b;
    layer0_outputs(1047) <= not b;
    layer0_outputs(1048) <= not (a or b);
    layer0_outputs(1049) <= a or b;
    layer0_outputs(1050) <= a or b;
    layer0_outputs(1051) <= 1'b0;
    layer0_outputs(1052) <= a;
    layer0_outputs(1053) <= b and not a;
    layer0_outputs(1054) <= a or b;
    layer0_outputs(1055) <= a;
    layer0_outputs(1056) <= a;
    layer0_outputs(1057) <= a and not b;
    layer0_outputs(1058) <= a or b;
    layer0_outputs(1059) <= not (a or b);
    layer0_outputs(1060) <= not (a or b);
    layer0_outputs(1061) <= not (a xor b);
    layer0_outputs(1062) <= a and not b;
    layer0_outputs(1063) <= not a;
    layer0_outputs(1064) <= a xor b;
    layer0_outputs(1065) <= a;
    layer0_outputs(1066) <= 1'b1;
    layer0_outputs(1067) <= not b or a;
    layer0_outputs(1068) <= not (a or b);
    layer0_outputs(1069) <= a and not b;
    layer0_outputs(1070) <= not (a or b);
    layer0_outputs(1071) <= a and b;
    layer0_outputs(1072) <= not a or b;
    layer0_outputs(1073) <= b and not a;
    layer0_outputs(1074) <= a;
    layer0_outputs(1075) <= a xor b;
    layer0_outputs(1076) <= b and not a;
    layer0_outputs(1077) <= b and not a;
    layer0_outputs(1078) <= not b or a;
    layer0_outputs(1079) <= a and b;
    layer0_outputs(1080) <= a or b;
    layer0_outputs(1081) <= 1'b1;
    layer0_outputs(1082) <= b;
    layer0_outputs(1083) <= not a;
    layer0_outputs(1084) <= not a;
    layer0_outputs(1085) <= not (a or b);
    layer0_outputs(1086) <= b and not a;
    layer0_outputs(1087) <= not b or a;
    layer0_outputs(1088) <= not (a xor b);
    layer0_outputs(1089) <= a or b;
    layer0_outputs(1090) <= 1'b0;
    layer0_outputs(1091) <= not (a or b);
    layer0_outputs(1092) <= a xor b;
    layer0_outputs(1093) <= b and not a;
    layer0_outputs(1094) <= not a or b;
    layer0_outputs(1095) <= b and not a;
    layer0_outputs(1096) <= not (a or b);
    layer0_outputs(1097) <= b;
    layer0_outputs(1098) <= not b;
    layer0_outputs(1099) <= not (a xor b);
    layer0_outputs(1100) <= a and b;
    layer0_outputs(1101) <= not (a xor b);
    layer0_outputs(1102) <= a or b;
    layer0_outputs(1103) <= not (a or b);
    layer0_outputs(1104) <= not (a or b);
    layer0_outputs(1105) <= not (a or b);
    layer0_outputs(1106) <= not (a or b);
    layer0_outputs(1107) <= a and not b;
    layer0_outputs(1108) <= not b or a;
    layer0_outputs(1109) <= a;
    layer0_outputs(1110) <= not (a or b);
    layer0_outputs(1111) <= not a or b;
    layer0_outputs(1112) <= b;
    layer0_outputs(1113) <= not b;
    layer0_outputs(1114) <= not b;
    layer0_outputs(1115) <= 1'b1;
    layer0_outputs(1116) <= a and not b;
    layer0_outputs(1117) <= a and b;
    layer0_outputs(1118) <= b and not a;
    layer0_outputs(1119) <= a or b;
    layer0_outputs(1120) <= a or b;
    layer0_outputs(1121) <= b;
    layer0_outputs(1122) <= not b or a;
    layer0_outputs(1123) <= a or b;
    layer0_outputs(1124) <= not a;
    layer0_outputs(1125) <= not a or b;
    layer0_outputs(1126) <= not (a or b);
    layer0_outputs(1127) <= not a;
    layer0_outputs(1128) <= 1'b1;
    layer0_outputs(1129) <= not (a xor b);
    layer0_outputs(1130) <= a xor b;
    layer0_outputs(1131) <= a and b;
    layer0_outputs(1132) <= a or b;
    layer0_outputs(1133) <= 1'b1;
    layer0_outputs(1134) <= a and b;
    layer0_outputs(1135) <= not a;
    layer0_outputs(1136) <= 1'b0;
    layer0_outputs(1137) <= not (a or b);
    layer0_outputs(1138) <= a;
    layer0_outputs(1139) <= not a or b;
    layer0_outputs(1140) <= not b;
    layer0_outputs(1141) <= a;
    layer0_outputs(1142) <= b and not a;
    layer0_outputs(1143) <= not a or b;
    layer0_outputs(1144) <= a and not b;
    layer0_outputs(1145) <= a and not b;
    layer0_outputs(1146) <= not a;
    layer0_outputs(1147) <= b;
    layer0_outputs(1148) <= b and not a;
    layer0_outputs(1149) <= not (a or b);
    layer0_outputs(1150) <= b and not a;
    layer0_outputs(1151) <= not (a xor b);
    layer0_outputs(1152) <= a or b;
    layer0_outputs(1153) <= not (a or b);
    layer0_outputs(1154) <= not (a xor b);
    layer0_outputs(1155) <= a or b;
    layer0_outputs(1156) <= 1'b0;
    layer0_outputs(1157) <= not a;
    layer0_outputs(1158) <= not b;
    layer0_outputs(1159) <= a and not b;
    layer0_outputs(1160) <= a;
    layer0_outputs(1161) <= not (a or b);
    layer0_outputs(1162) <= a xor b;
    layer0_outputs(1163) <= not a or b;
    layer0_outputs(1164) <= not b;
    layer0_outputs(1165) <= a or b;
    layer0_outputs(1166) <= not a or b;
    layer0_outputs(1167) <= a;
    layer0_outputs(1168) <= 1'b0;
    layer0_outputs(1169) <= not (a or b);
    layer0_outputs(1170) <= a xor b;
    layer0_outputs(1171) <= not (a or b);
    layer0_outputs(1172) <= not b;
    layer0_outputs(1173) <= a and b;
    layer0_outputs(1174) <= a or b;
    layer0_outputs(1175) <= not (a xor b);
    layer0_outputs(1176) <= not b;
    layer0_outputs(1177) <= a or b;
    layer0_outputs(1178) <= not a or b;
    layer0_outputs(1179) <= a;
    layer0_outputs(1180) <= not b;
    layer0_outputs(1181) <= not (a or b);
    layer0_outputs(1182) <= b;
    layer0_outputs(1183) <= a;
    layer0_outputs(1184) <= b and not a;
    layer0_outputs(1185) <= a;
    layer0_outputs(1186) <= a xor b;
    layer0_outputs(1187) <= b;
    layer0_outputs(1188) <= a or b;
    layer0_outputs(1189) <= not (a or b);
    layer0_outputs(1190) <= a and not b;
    layer0_outputs(1191) <= not a or b;
    layer0_outputs(1192) <= not a;
    layer0_outputs(1193) <= a or b;
    layer0_outputs(1194) <= a or b;
    layer0_outputs(1195) <= a xor b;
    layer0_outputs(1196) <= not (a or b);
    layer0_outputs(1197) <= not (a or b);
    layer0_outputs(1198) <= b;
    layer0_outputs(1199) <= a or b;
    layer0_outputs(1200) <= a or b;
    layer0_outputs(1201) <= a;
    layer0_outputs(1202) <= not (a xor b);
    layer0_outputs(1203) <= not a or b;
    layer0_outputs(1204) <= a and not b;
    layer0_outputs(1205) <= a or b;
    layer0_outputs(1206) <= not (a or b);
    layer0_outputs(1207) <= not b or a;
    layer0_outputs(1208) <= a or b;
    layer0_outputs(1209) <= b;
    layer0_outputs(1210) <= 1'b1;
    layer0_outputs(1211) <= not b;
    layer0_outputs(1212) <= a or b;
    layer0_outputs(1213) <= a and not b;
    layer0_outputs(1214) <= not b or a;
    layer0_outputs(1215) <= a and not b;
    layer0_outputs(1216) <= a xor b;
    layer0_outputs(1217) <= a;
    layer0_outputs(1218) <= not (a or b);
    layer0_outputs(1219) <= a xor b;
    layer0_outputs(1220) <= a and not b;
    layer0_outputs(1221) <= a or b;
    layer0_outputs(1222) <= b;
    layer0_outputs(1223) <= not (a or b);
    layer0_outputs(1224) <= not a;
    layer0_outputs(1225) <= not a;
    layer0_outputs(1226) <= not b;
    layer0_outputs(1227) <= not (a or b);
    layer0_outputs(1228) <= a or b;
    layer0_outputs(1229) <= not (a xor b);
    layer0_outputs(1230) <= b;
    layer0_outputs(1231) <= not b;
    layer0_outputs(1232) <= not (a and b);
    layer0_outputs(1233) <= a;
    layer0_outputs(1234) <= not (a or b);
    layer0_outputs(1235) <= a or b;
    layer0_outputs(1236) <= not b or a;
    layer0_outputs(1237) <= a;
    layer0_outputs(1238) <= not a;
    layer0_outputs(1239) <= a;
    layer0_outputs(1240) <= not a;
    layer0_outputs(1241) <= a or b;
    layer0_outputs(1242) <= 1'b1;
    layer0_outputs(1243) <= a;
    layer0_outputs(1244) <= b;
    layer0_outputs(1245) <= a or b;
    layer0_outputs(1246) <= not (a or b);
    layer0_outputs(1247) <= a or b;
    layer0_outputs(1248) <= not a;
    layer0_outputs(1249) <= not (a or b);
    layer0_outputs(1250) <= not (a or b);
    layer0_outputs(1251) <= not b or a;
    layer0_outputs(1252) <= b;
    layer0_outputs(1253) <= b;
    layer0_outputs(1254) <= not (a xor b);
    layer0_outputs(1255) <= not (a or b);
    layer0_outputs(1256) <= a xor b;
    layer0_outputs(1257) <= not (a xor b);
    layer0_outputs(1258) <= b;
    layer0_outputs(1259) <= not b;
    layer0_outputs(1260) <= b;
    layer0_outputs(1261) <= not b;
    layer0_outputs(1262) <= not b or a;
    layer0_outputs(1263) <= not (a or b);
    layer0_outputs(1264) <= a or b;
    layer0_outputs(1265) <= a or b;
    layer0_outputs(1266) <= a and not b;
    layer0_outputs(1267) <= not (a xor b);
    layer0_outputs(1268) <= not (a or b);
    layer0_outputs(1269) <= not (a or b);
    layer0_outputs(1270) <= a or b;
    layer0_outputs(1271) <= not b or a;
    layer0_outputs(1272) <= not (a xor b);
    layer0_outputs(1273) <= not a;
    layer0_outputs(1274) <= not b or a;
    layer0_outputs(1275) <= not a;
    layer0_outputs(1276) <= not (a or b);
    layer0_outputs(1277) <= not (a and b);
    layer0_outputs(1278) <= 1'b1;
    layer0_outputs(1279) <= not (a xor b);
    layer0_outputs(1280) <= not (a or b);
    layer0_outputs(1281) <= not (a or b);
    layer0_outputs(1282) <= a or b;
    layer0_outputs(1283) <= a xor b;
    layer0_outputs(1284) <= 1'b0;
    layer0_outputs(1285) <= not (a or b);
    layer0_outputs(1286) <= a and b;
    layer0_outputs(1287) <= not a;
    layer0_outputs(1288) <= not (a xor b);
    layer0_outputs(1289) <= a;
    layer0_outputs(1290) <= not b or a;
    layer0_outputs(1291) <= not a or b;
    layer0_outputs(1292) <= b and not a;
    layer0_outputs(1293) <= a or b;
    layer0_outputs(1294) <= not (a or b);
    layer0_outputs(1295) <= not a;
    layer0_outputs(1296) <= b;
    layer0_outputs(1297) <= not b;
    layer0_outputs(1298) <= not (a xor b);
    layer0_outputs(1299) <= a xor b;
    layer0_outputs(1300) <= not (a xor b);
    layer0_outputs(1301) <= not a or b;
    layer0_outputs(1302) <= a or b;
    layer0_outputs(1303) <= not (a or b);
    layer0_outputs(1304) <= a and not b;
    layer0_outputs(1305) <= not (a and b);
    layer0_outputs(1306) <= a and not b;
    layer0_outputs(1307) <= a and not b;
    layer0_outputs(1308) <= not (a and b);
    layer0_outputs(1309) <= a;
    layer0_outputs(1310) <= not (a and b);
    layer0_outputs(1311) <= not (a xor b);
    layer0_outputs(1312) <= a or b;
    layer0_outputs(1313) <= a or b;
    layer0_outputs(1314) <= not b or a;
    layer0_outputs(1315) <= a or b;
    layer0_outputs(1316) <= not a;
    layer0_outputs(1317) <= a or b;
    layer0_outputs(1318) <= not b;
    layer0_outputs(1319) <= not (a or b);
    layer0_outputs(1320) <= a or b;
    layer0_outputs(1321) <= not a;
    layer0_outputs(1322) <= b and not a;
    layer0_outputs(1323) <= a or b;
    layer0_outputs(1324) <= a xor b;
    layer0_outputs(1325) <= b;
    layer0_outputs(1326) <= not (a or b);
    layer0_outputs(1327) <= not (a or b);
    layer0_outputs(1328) <= not a;
    layer0_outputs(1329) <= a and not b;
    layer0_outputs(1330) <= a or b;
    layer0_outputs(1331) <= b;
    layer0_outputs(1332) <= not a;
    layer0_outputs(1333) <= not (a or b);
    layer0_outputs(1334) <= a xor b;
    layer0_outputs(1335) <= not (a or b);
    layer0_outputs(1336) <= a or b;
    layer0_outputs(1337) <= a xor b;
    layer0_outputs(1338) <= not b or a;
    layer0_outputs(1339) <= not (a xor b);
    layer0_outputs(1340) <= a;
    layer0_outputs(1341) <= not a or b;
    layer0_outputs(1342) <= a or b;
    layer0_outputs(1343) <= not b;
    layer0_outputs(1344) <= not (a or b);
    layer0_outputs(1345) <= a or b;
    layer0_outputs(1346) <= not b;
    layer0_outputs(1347) <= not (a or b);
    layer0_outputs(1348) <= not b;
    layer0_outputs(1349) <= a and not b;
    layer0_outputs(1350) <= not (a or b);
    layer0_outputs(1351) <= not b or a;
    layer0_outputs(1352) <= a or b;
    layer0_outputs(1353) <= a;
    layer0_outputs(1354) <= not (a xor b);
    layer0_outputs(1355) <= not b or a;
    layer0_outputs(1356) <= not b or a;
    layer0_outputs(1357) <= a and not b;
    layer0_outputs(1358) <= not a or b;
    layer0_outputs(1359) <= not a;
    layer0_outputs(1360) <= a or b;
    layer0_outputs(1361) <= 1'b1;
    layer0_outputs(1362) <= a or b;
    layer0_outputs(1363) <= not b or a;
    layer0_outputs(1364) <= b;
    layer0_outputs(1365) <= a or b;
    layer0_outputs(1366) <= a xor b;
    layer0_outputs(1367) <= not b or a;
    layer0_outputs(1368) <= not a;
    layer0_outputs(1369) <= not b or a;
    layer0_outputs(1370) <= b and not a;
    layer0_outputs(1371) <= not b;
    layer0_outputs(1372) <= 1'b0;
    layer0_outputs(1373) <= not (a or b);
    layer0_outputs(1374) <= a or b;
    layer0_outputs(1375) <= a;
    layer0_outputs(1376) <= b and not a;
    layer0_outputs(1377) <= b;
    layer0_outputs(1378) <= not a;
    layer0_outputs(1379) <= 1'b1;
    layer0_outputs(1380) <= not (a and b);
    layer0_outputs(1381) <= b and not a;
    layer0_outputs(1382) <= a;
    layer0_outputs(1383) <= not (a xor b);
    layer0_outputs(1384) <= a;
    layer0_outputs(1385) <= a xor b;
    layer0_outputs(1386) <= not a or b;
    layer0_outputs(1387) <= not (a xor b);
    layer0_outputs(1388) <= a;
    layer0_outputs(1389) <= not b;
    layer0_outputs(1390) <= 1'b0;
    layer0_outputs(1391) <= not (a or b);
    layer0_outputs(1392) <= a and not b;
    layer0_outputs(1393) <= a or b;
    layer0_outputs(1394) <= not b or a;
    layer0_outputs(1395) <= a or b;
    layer0_outputs(1396) <= a or b;
    layer0_outputs(1397) <= a;
    layer0_outputs(1398) <= not b;
    layer0_outputs(1399) <= b;
    layer0_outputs(1400) <= not b or a;
    layer0_outputs(1401) <= not (a or b);
    layer0_outputs(1402) <= b and not a;
    layer0_outputs(1403) <= a xor b;
    layer0_outputs(1404) <= a xor b;
    layer0_outputs(1405) <= not (a or b);
    layer0_outputs(1406) <= not a;
    layer0_outputs(1407) <= not b or a;
    layer0_outputs(1408) <= a or b;
    layer0_outputs(1409) <= a or b;
    layer0_outputs(1410) <= a and not b;
    layer0_outputs(1411) <= not (a or b);
    layer0_outputs(1412) <= a and b;
    layer0_outputs(1413) <= not a or b;
    layer0_outputs(1414) <= not (a xor b);
    layer0_outputs(1415) <= a xor b;
    layer0_outputs(1416) <= not b;
    layer0_outputs(1417) <= a;
    layer0_outputs(1418) <= not b or a;
    layer0_outputs(1419) <= b;
    layer0_outputs(1420) <= not a or b;
    layer0_outputs(1421) <= not a;
    layer0_outputs(1422) <= not (a and b);
    layer0_outputs(1423) <= not (a xor b);
    layer0_outputs(1424) <= a or b;
    layer0_outputs(1425) <= not b or a;
    layer0_outputs(1426) <= a or b;
    layer0_outputs(1427) <= a or b;
    layer0_outputs(1428) <= a and not b;
    layer0_outputs(1429) <= a or b;
    layer0_outputs(1430) <= not (a or b);
    layer0_outputs(1431) <= not a;
    layer0_outputs(1432) <= b;
    layer0_outputs(1433) <= not a or b;
    layer0_outputs(1434) <= a;
    layer0_outputs(1435) <= not b;
    layer0_outputs(1436) <= b;
    layer0_outputs(1437) <= not b;
    layer0_outputs(1438) <= not (a or b);
    layer0_outputs(1439) <= b;
    layer0_outputs(1440) <= not a;
    layer0_outputs(1441) <= not (a or b);
    layer0_outputs(1442) <= a;
    layer0_outputs(1443) <= b;
    layer0_outputs(1444) <= not b;
    layer0_outputs(1445) <= 1'b1;
    layer0_outputs(1446) <= a;
    layer0_outputs(1447) <= not b or a;
    layer0_outputs(1448) <= b;
    layer0_outputs(1449) <= a or b;
    layer0_outputs(1450) <= not a;
    layer0_outputs(1451) <= 1'b1;
    layer0_outputs(1452) <= b and not a;
    layer0_outputs(1453) <= a xor b;
    layer0_outputs(1454) <= not (a or b);
    layer0_outputs(1455) <= b;
    layer0_outputs(1456) <= b;
    layer0_outputs(1457) <= b and not a;
    layer0_outputs(1458) <= not (a or b);
    layer0_outputs(1459) <= not a or b;
    layer0_outputs(1460) <= a;
    layer0_outputs(1461) <= not b;
    layer0_outputs(1462) <= a and not b;
    layer0_outputs(1463) <= not (a xor b);
    layer0_outputs(1464) <= not a or b;
    layer0_outputs(1465) <= a xor b;
    layer0_outputs(1466) <= a and not b;
    layer0_outputs(1467) <= a xor b;
    layer0_outputs(1468) <= b;
    layer0_outputs(1469) <= a and not b;
    layer0_outputs(1470) <= not (a and b);
    layer0_outputs(1471) <= not a or b;
    layer0_outputs(1472) <= a or b;
    layer0_outputs(1473) <= not (a xor b);
    layer0_outputs(1474) <= not b;
    layer0_outputs(1475) <= a xor b;
    layer0_outputs(1476) <= not (a or b);
    layer0_outputs(1477) <= a and not b;
    layer0_outputs(1478) <= b;
    layer0_outputs(1479) <= a and b;
    layer0_outputs(1480) <= b and not a;
    layer0_outputs(1481) <= b and not a;
    layer0_outputs(1482) <= a or b;
    layer0_outputs(1483) <= a;
    layer0_outputs(1484) <= not (a xor b);
    layer0_outputs(1485) <= not (a or b);
    layer0_outputs(1486) <= a xor b;
    layer0_outputs(1487) <= not (a xor b);
    layer0_outputs(1488) <= a;
    layer0_outputs(1489) <= not (a or b);
    layer0_outputs(1490) <= a;
    layer0_outputs(1491) <= a and b;
    layer0_outputs(1492) <= a or b;
    layer0_outputs(1493) <= b;
    layer0_outputs(1494) <= not (a or b);
    layer0_outputs(1495) <= a or b;
    layer0_outputs(1496) <= 1'b1;
    layer0_outputs(1497) <= not (a or b);
    layer0_outputs(1498) <= a or b;
    layer0_outputs(1499) <= a and not b;
    layer0_outputs(1500) <= not (a or b);
    layer0_outputs(1501) <= not (a xor b);
    layer0_outputs(1502) <= a and not b;
    layer0_outputs(1503) <= a and not b;
    layer0_outputs(1504) <= not (a or b);
    layer0_outputs(1505) <= not (a or b);
    layer0_outputs(1506) <= not a;
    layer0_outputs(1507) <= a and b;
    layer0_outputs(1508) <= a;
    layer0_outputs(1509) <= not a;
    layer0_outputs(1510) <= not a or b;
    layer0_outputs(1511) <= a;
    layer0_outputs(1512) <= b and not a;
    layer0_outputs(1513) <= b;
    layer0_outputs(1514) <= not a or b;
    layer0_outputs(1515) <= not a or b;
    layer0_outputs(1516) <= a or b;
    layer0_outputs(1517) <= not a;
    layer0_outputs(1518) <= not (a xor b);
    layer0_outputs(1519) <= a or b;
    layer0_outputs(1520) <= a or b;
    layer0_outputs(1521) <= not (a and b);
    layer0_outputs(1522) <= not a;
    layer0_outputs(1523) <= not (a or b);
    layer0_outputs(1524) <= not (a xor b);
    layer0_outputs(1525) <= not (a or b);
    layer0_outputs(1526) <= not b or a;
    layer0_outputs(1527) <= a or b;
    layer0_outputs(1528) <= b;
    layer0_outputs(1529) <= not a;
    layer0_outputs(1530) <= not (a or b);
    layer0_outputs(1531) <= not a or b;
    layer0_outputs(1532) <= not a;
    layer0_outputs(1533) <= not (a or b);
    layer0_outputs(1534) <= a and not b;
    layer0_outputs(1535) <= not (a and b);
    layer0_outputs(1536) <= not b or a;
    layer0_outputs(1537) <= a or b;
    layer0_outputs(1538) <= a or b;
    layer0_outputs(1539) <= not b or a;
    layer0_outputs(1540) <= a or b;
    layer0_outputs(1541) <= a or b;
    layer0_outputs(1542) <= b;
    layer0_outputs(1543) <= not (a and b);
    layer0_outputs(1544) <= a xor b;
    layer0_outputs(1545) <= a or b;
    layer0_outputs(1546) <= a and not b;
    layer0_outputs(1547) <= not b or a;
    layer0_outputs(1548) <= not b;
    layer0_outputs(1549) <= not (a or b);
    layer0_outputs(1550) <= a;
    layer0_outputs(1551) <= b;
    layer0_outputs(1552) <= a xor b;
    layer0_outputs(1553) <= a xor b;
    layer0_outputs(1554) <= not a;
    layer0_outputs(1555) <= a or b;
    layer0_outputs(1556) <= b;
    layer0_outputs(1557) <= not (a and b);
    layer0_outputs(1558) <= a and b;
    layer0_outputs(1559) <= not b or a;
    layer0_outputs(1560) <= not (a xor b);
    layer0_outputs(1561) <= not (a xor b);
    layer0_outputs(1562) <= not (a xor b);
    layer0_outputs(1563) <= 1'b1;
    layer0_outputs(1564) <= not (a or b);
    layer0_outputs(1565) <= not a;
    layer0_outputs(1566) <= not (a or b);
    layer0_outputs(1567) <= a or b;
    layer0_outputs(1568) <= not (a or b);
    layer0_outputs(1569) <= not a;
    layer0_outputs(1570) <= b;
    layer0_outputs(1571) <= a;
    layer0_outputs(1572) <= a xor b;
    layer0_outputs(1573) <= b and not a;
    layer0_outputs(1574) <= a or b;
    layer0_outputs(1575) <= a and not b;
    layer0_outputs(1576) <= a;
    layer0_outputs(1577) <= b;
    layer0_outputs(1578) <= not (a or b);
    layer0_outputs(1579) <= a xor b;
    layer0_outputs(1580) <= not b or a;
    layer0_outputs(1581) <= not (a or b);
    layer0_outputs(1582) <= not b;
    layer0_outputs(1583) <= a or b;
    layer0_outputs(1584) <= not b or a;
    layer0_outputs(1585) <= b and not a;
    layer0_outputs(1586) <= not a;
    layer0_outputs(1587) <= not a;
    layer0_outputs(1588) <= not (a or b);
    layer0_outputs(1589) <= a or b;
    layer0_outputs(1590) <= not (a or b);
    layer0_outputs(1591) <= a or b;
    layer0_outputs(1592) <= b and not a;
    layer0_outputs(1593) <= b;
    layer0_outputs(1594) <= a or b;
    layer0_outputs(1595) <= not a or b;
    layer0_outputs(1596) <= b;
    layer0_outputs(1597) <= a or b;
    layer0_outputs(1598) <= not (a or b);
    layer0_outputs(1599) <= not b or a;
    layer0_outputs(1600) <= not a or b;
    layer0_outputs(1601) <= a or b;
    layer0_outputs(1602) <= not a;
    layer0_outputs(1603) <= a xor b;
    layer0_outputs(1604) <= b and not a;
    layer0_outputs(1605) <= a and not b;
    layer0_outputs(1606) <= a or b;
    layer0_outputs(1607) <= a xor b;
    layer0_outputs(1608) <= not (a or b);
    layer0_outputs(1609) <= not (a or b);
    layer0_outputs(1610) <= not (a or b);
    layer0_outputs(1611) <= a or b;
    layer0_outputs(1612) <= b;
    layer0_outputs(1613) <= b and not a;
    layer0_outputs(1614) <= 1'b1;
    layer0_outputs(1615) <= b and not a;
    layer0_outputs(1616) <= not (a xor b);
    layer0_outputs(1617) <= a;
    layer0_outputs(1618) <= not b or a;
    layer0_outputs(1619) <= a or b;
    layer0_outputs(1620) <= a or b;
    layer0_outputs(1621) <= not (a or b);
    layer0_outputs(1622) <= not (a or b);
    layer0_outputs(1623) <= not a or b;
    layer0_outputs(1624) <= not a or b;
    layer0_outputs(1625) <= a xor b;
    layer0_outputs(1626) <= not (a xor b);
    layer0_outputs(1627) <= not (a or b);
    layer0_outputs(1628) <= a or b;
    layer0_outputs(1629) <= not (a or b);
    layer0_outputs(1630) <= b and not a;
    layer0_outputs(1631) <= a;
    layer0_outputs(1632) <= a and not b;
    layer0_outputs(1633) <= not (a xor b);
    layer0_outputs(1634) <= a and not b;
    layer0_outputs(1635) <= a and not b;
    layer0_outputs(1636) <= a and not b;
    layer0_outputs(1637) <= not a or b;
    layer0_outputs(1638) <= not (a or b);
    layer0_outputs(1639) <= a or b;
    layer0_outputs(1640) <= a xor b;
    layer0_outputs(1641) <= not (a or b);
    layer0_outputs(1642) <= not a or b;
    layer0_outputs(1643) <= a and not b;
    layer0_outputs(1644) <= a xor b;
    layer0_outputs(1645) <= a;
    layer0_outputs(1646) <= not (a xor b);
    layer0_outputs(1647) <= not a;
    layer0_outputs(1648) <= not a or b;
    layer0_outputs(1649) <= not b;
    layer0_outputs(1650) <= not (a and b);
    layer0_outputs(1651) <= a or b;
    layer0_outputs(1652) <= not (a xor b);
    layer0_outputs(1653) <= a or b;
    layer0_outputs(1654) <= 1'b0;
    layer0_outputs(1655) <= a;
    layer0_outputs(1656) <= not b or a;
    layer0_outputs(1657) <= not b;
    layer0_outputs(1658) <= b;
    layer0_outputs(1659) <= b;
    layer0_outputs(1660) <= not a;
    layer0_outputs(1661) <= a or b;
    layer0_outputs(1662) <= not (a xor b);
    layer0_outputs(1663) <= b and not a;
    layer0_outputs(1664) <= a;
    layer0_outputs(1665) <= a and not b;
    layer0_outputs(1666) <= not (a or b);
    layer0_outputs(1667) <= a xor b;
    layer0_outputs(1668) <= b and not a;
    layer0_outputs(1669) <= a;
    layer0_outputs(1670) <= a and not b;
    layer0_outputs(1671) <= a or b;
    layer0_outputs(1672) <= a or b;
    layer0_outputs(1673) <= not b;
    layer0_outputs(1674) <= b and not a;
    layer0_outputs(1675) <= not (a or b);
    layer0_outputs(1676) <= not b;
    layer0_outputs(1677) <= a and b;
    layer0_outputs(1678) <= a and not b;
    layer0_outputs(1679) <= a xor b;
    layer0_outputs(1680) <= not b;
    layer0_outputs(1681) <= not a or b;
    layer0_outputs(1682) <= not a;
    layer0_outputs(1683) <= not b;
    layer0_outputs(1684) <= not a;
    layer0_outputs(1685) <= a or b;
    layer0_outputs(1686) <= b and not a;
    layer0_outputs(1687) <= not (a xor b);
    layer0_outputs(1688) <= a;
    layer0_outputs(1689) <= not (a xor b);
    layer0_outputs(1690) <= a or b;
    layer0_outputs(1691) <= not (a xor b);
    layer0_outputs(1692) <= a and b;
    layer0_outputs(1693) <= b;
    layer0_outputs(1694) <= a or b;
    layer0_outputs(1695) <= not a;
    layer0_outputs(1696) <= b;
    layer0_outputs(1697) <= b;
    layer0_outputs(1698) <= not b;
    layer0_outputs(1699) <= not (a or b);
    layer0_outputs(1700) <= not b;
    layer0_outputs(1701) <= a xor b;
    layer0_outputs(1702) <= not (a xor b);
    layer0_outputs(1703) <= b;
    layer0_outputs(1704) <= a and not b;
    layer0_outputs(1705) <= a and b;
    layer0_outputs(1706) <= a xor b;
    layer0_outputs(1707) <= a and not b;
    layer0_outputs(1708) <= not b;
    layer0_outputs(1709) <= not (a or b);
    layer0_outputs(1710) <= 1'b0;
    layer0_outputs(1711) <= not a or b;
    layer0_outputs(1712) <= not a;
    layer0_outputs(1713) <= b and not a;
    layer0_outputs(1714) <= 1'b0;
    layer0_outputs(1715) <= a or b;
    layer0_outputs(1716) <= not (a or b);
    layer0_outputs(1717) <= a and not b;
    layer0_outputs(1718) <= not b;
    layer0_outputs(1719) <= not a;
    layer0_outputs(1720) <= a or b;
    layer0_outputs(1721) <= not (a or b);
    layer0_outputs(1722) <= not a or b;
    layer0_outputs(1723) <= a and b;
    layer0_outputs(1724) <= not (a or b);
    layer0_outputs(1725) <= not (a xor b);
    layer0_outputs(1726) <= b and not a;
    layer0_outputs(1727) <= a xor b;
    layer0_outputs(1728) <= b and not a;
    layer0_outputs(1729) <= a or b;
    layer0_outputs(1730) <= 1'b0;
    layer0_outputs(1731) <= not (a or b);
    layer0_outputs(1732) <= not b;
    layer0_outputs(1733) <= a and not b;
    layer0_outputs(1734) <= not (a or b);
    layer0_outputs(1735) <= not a or b;
    layer0_outputs(1736) <= not a;
    layer0_outputs(1737) <= not (a xor b);
    layer0_outputs(1738) <= not a or b;
    layer0_outputs(1739) <= not (a or b);
    layer0_outputs(1740) <= not (a xor b);
    layer0_outputs(1741) <= not a;
    layer0_outputs(1742) <= b;
    layer0_outputs(1743) <= not a or b;
    layer0_outputs(1744) <= b;
    layer0_outputs(1745) <= a;
    layer0_outputs(1746) <= a and not b;
    layer0_outputs(1747) <= not (a or b);
    layer0_outputs(1748) <= a or b;
    layer0_outputs(1749) <= b;
    layer0_outputs(1750) <= not a;
    layer0_outputs(1751) <= b and not a;
    layer0_outputs(1752) <= a or b;
    layer0_outputs(1753) <= not a or b;
    layer0_outputs(1754) <= a;
    layer0_outputs(1755) <= b and not a;
    layer0_outputs(1756) <= not b;
    layer0_outputs(1757) <= a and not b;
    layer0_outputs(1758) <= a xor b;
    layer0_outputs(1759) <= not a;
    layer0_outputs(1760) <= a or b;
    layer0_outputs(1761) <= b;
    layer0_outputs(1762) <= not (a or b);
    layer0_outputs(1763) <= a or b;
    layer0_outputs(1764) <= not (a and b);
    layer0_outputs(1765) <= a;
    layer0_outputs(1766) <= not b;
    layer0_outputs(1767) <= b;
    layer0_outputs(1768) <= b and not a;
    layer0_outputs(1769) <= not a;
    layer0_outputs(1770) <= b;
    layer0_outputs(1771) <= a xor b;
    layer0_outputs(1772) <= a or b;
    layer0_outputs(1773) <= not (a xor b);
    layer0_outputs(1774) <= b and not a;
    layer0_outputs(1775) <= a or b;
    layer0_outputs(1776) <= not b or a;
    layer0_outputs(1777) <= not (a or b);
    layer0_outputs(1778) <= a and not b;
    layer0_outputs(1779) <= b;
    layer0_outputs(1780) <= not b or a;
    layer0_outputs(1781) <= not a or b;
    layer0_outputs(1782) <= b and not a;
    layer0_outputs(1783) <= not (a or b);
    layer0_outputs(1784) <= not a;
    layer0_outputs(1785) <= not b or a;
    layer0_outputs(1786) <= not (a xor b);
    layer0_outputs(1787) <= a and not b;
    layer0_outputs(1788) <= not (a or b);
    layer0_outputs(1789) <= a and not b;
    layer0_outputs(1790) <= not b or a;
    layer0_outputs(1791) <= not a or b;
    layer0_outputs(1792) <= not (a or b);
    layer0_outputs(1793) <= not a or b;
    layer0_outputs(1794) <= b and not a;
    layer0_outputs(1795) <= not (a or b);
    layer0_outputs(1796) <= not (a xor b);
    layer0_outputs(1797) <= a and not b;
    layer0_outputs(1798) <= not (a or b);
    layer0_outputs(1799) <= not a or b;
    layer0_outputs(1800) <= a;
    layer0_outputs(1801) <= not b or a;
    layer0_outputs(1802) <= a and not b;
    layer0_outputs(1803) <= not a or b;
    layer0_outputs(1804) <= not b;
    layer0_outputs(1805) <= not (a xor b);
    layer0_outputs(1806) <= not (a xor b);
    layer0_outputs(1807) <= not b;
    layer0_outputs(1808) <= a xor b;
    layer0_outputs(1809) <= not a;
    layer0_outputs(1810) <= not (a and b);
    layer0_outputs(1811) <= not b or a;
    layer0_outputs(1812) <= not a;
    layer0_outputs(1813) <= not b;
    layer0_outputs(1814) <= not a or b;
    layer0_outputs(1815) <= not (a xor b);
    layer0_outputs(1816) <= not a;
    layer0_outputs(1817) <= b;
    layer0_outputs(1818) <= not (a or b);
    layer0_outputs(1819) <= not (a or b);
    layer0_outputs(1820) <= not (a or b);
    layer0_outputs(1821) <= not b or a;
    layer0_outputs(1822) <= a xor b;
    layer0_outputs(1823) <= not (a or b);
    layer0_outputs(1824) <= a or b;
    layer0_outputs(1825) <= not (a xor b);
    layer0_outputs(1826) <= not b or a;
    layer0_outputs(1827) <= not b or a;
    layer0_outputs(1828) <= not (a and b);
    layer0_outputs(1829) <= not b or a;
    layer0_outputs(1830) <= a and not b;
    layer0_outputs(1831) <= a or b;
    layer0_outputs(1832) <= a or b;
    layer0_outputs(1833) <= not a;
    layer0_outputs(1834) <= a xor b;
    layer0_outputs(1835) <= not (a or b);
    layer0_outputs(1836) <= not a;
    layer0_outputs(1837) <= not b or a;
    layer0_outputs(1838) <= not b;
    layer0_outputs(1839) <= not (a and b);
    layer0_outputs(1840) <= b and not a;
    layer0_outputs(1841) <= not a;
    layer0_outputs(1842) <= a or b;
    layer0_outputs(1843) <= not (a or b);
    layer0_outputs(1844) <= b;
    layer0_outputs(1845) <= not (a or b);
    layer0_outputs(1846) <= a and not b;
    layer0_outputs(1847) <= not b;
    layer0_outputs(1848) <= a and not b;
    layer0_outputs(1849) <= not (a xor b);
    layer0_outputs(1850) <= not (a xor b);
    layer0_outputs(1851) <= a or b;
    layer0_outputs(1852) <= not (a or b);
    layer0_outputs(1853) <= not a or b;
    layer0_outputs(1854) <= not (a and b);
    layer0_outputs(1855) <= b and not a;
    layer0_outputs(1856) <= a or b;
    layer0_outputs(1857) <= b and not a;
    layer0_outputs(1858) <= b;
    layer0_outputs(1859) <= a;
    layer0_outputs(1860) <= a;
    layer0_outputs(1861) <= not b or a;
    layer0_outputs(1862) <= a;
    layer0_outputs(1863) <= not (a or b);
    layer0_outputs(1864) <= a and not b;
    layer0_outputs(1865) <= a or b;
    layer0_outputs(1866) <= not (a or b);
    layer0_outputs(1867) <= a xor b;
    layer0_outputs(1868) <= not b;
    layer0_outputs(1869) <= not (a or b);
    layer0_outputs(1870) <= b and not a;
    layer0_outputs(1871) <= a or b;
    layer0_outputs(1872) <= not a;
    layer0_outputs(1873) <= a or b;
    layer0_outputs(1874) <= a or b;
    layer0_outputs(1875) <= not (a or b);
    layer0_outputs(1876) <= a or b;
    layer0_outputs(1877) <= a or b;
    layer0_outputs(1878) <= b;
    layer0_outputs(1879) <= a xor b;
    layer0_outputs(1880) <= not b or a;
    layer0_outputs(1881) <= a or b;
    layer0_outputs(1882) <= b and not a;
    layer0_outputs(1883) <= b;
    layer0_outputs(1884) <= not (a xor b);
    layer0_outputs(1885) <= a or b;
    layer0_outputs(1886) <= not (a and b);
    layer0_outputs(1887) <= not (a or b);
    layer0_outputs(1888) <= a or b;
    layer0_outputs(1889) <= a;
    layer0_outputs(1890) <= b and not a;
    layer0_outputs(1891) <= not a or b;
    layer0_outputs(1892) <= not (a or b);
    layer0_outputs(1893) <= not a;
    layer0_outputs(1894) <= a and not b;
    layer0_outputs(1895) <= not a or b;
    layer0_outputs(1896) <= not (a xor b);
    layer0_outputs(1897) <= not (a or b);
    layer0_outputs(1898) <= not (a or b);
    layer0_outputs(1899) <= not a or b;
    layer0_outputs(1900) <= a xor b;
    layer0_outputs(1901) <= not b or a;
    layer0_outputs(1902) <= not (a or b);
    layer0_outputs(1903) <= a and b;
    layer0_outputs(1904) <= not (a xor b);
    layer0_outputs(1905) <= not (a or b);
    layer0_outputs(1906) <= a and b;
    layer0_outputs(1907) <= not (a xor b);
    layer0_outputs(1908) <= a and not b;
    layer0_outputs(1909) <= b and not a;
    layer0_outputs(1910) <= not (a or b);
    layer0_outputs(1911) <= a;
    layer0_outputs(1912) <= a or b;
    layer0_outputs(1913) <= b;
    layer0_outputs(1914) <= not (a xor b);
    layer0_outputs(1915) <= a and not b;
    layer0_outputs(1916) <= not b or a;
    layer0_outputs(1917) <= b;
    layer0_outputs(1918) <= not a or b;
    layer0_outputs(1919) <= not (a or b);
    layer0_outputs(1920) <= a;
    layer0_outputs(1921) <= b;
    layer0_outputs(1922) <= b and not a;
    layer0_outputs(1923) <= a or b;
    layer0_outputs(1924) <= not (a or b);
    layer0_outputs(1925) <= a or b;
    layer0_outputs(1926) <= not (a or b);
    layer0_outputs(1927) <= not (a xor b);
    layer0_outputs(1928) <= not (a or b);
    layer0_outputs(1929) <= 1'b1;
    layer0_outputs(1930) <= a or b;
    layer0_outputs(1931) <= b;
    layer0_outputs(1932) <= not (a xor b);
    layer0_outputs(1933) <= a or b;
    layer0_outputs(1934) <= not b or a;
    layer0_outputs(1935) <= not (a xor b);
    layer0_outputs(1936) <= a or b;
    layer0_outputs(1937) <= a or b;
    layer0_outputs(1938) <= a or b;
    layer0_outputs(1939) <= not b or a;
    layer0_outputs(1940) <= a or b;
    layer0_outputs(1941) <= b and not a;
    layer0_outputs(1942) <= a xor b;
    layer0_outputs(1943) <= b and not a;
    layer0_outputs(1944) <= a and not b;
    layer0_outputs(1945) <= not a or b;
    layer0_outputs(1946) <= a and not b;
    layer0_outputs(1947) <= not b;
    layer0_outputs(1948) <= not a or b;
    layer0_outputs(1949) <= a or b;
    layer0_outputs(1950) <= a and not b;
    layer0_outputs(1951) <= not b or a;
    layer0_outputs(1952) <= a xor b;
    layer0_outputs(1953) <= not (a and b);
    layer0_outputs(1954) <= a and not b;
    layer0_outputs(1955) <= b;
    layer0_outputs(1956) <= not b or a;
    layer0_outputs(1957) <= not a or b;
    layer0_outputs(1958) <= not (a xor b);
    layer0_outputs(1959) <= not a or b;
    layer0_outputs(1960) <= a xor b;
    layer0_outputs(1961) <= not (a xor b);
    layer0_outputs(1962) <= a;
    layer0_outputs(1963) <= not (a xor b);
    layer0_outputs(1964) <= not (a or b);
    layer0_outputs(1965) <= not a or b;
    layer0_outputs(1966) <= b;
    layer0_outputs(1967) <= not b;
    layer0_outputs(1968) <= not (a xor b);
    layer0_outputs(1969) <= b;
    layer0_outputs(1970) <= not (a or b);
    layer0_outputs(1971) <= a and b;
    layer0_outputs(1972) <= a or b;
    layer0_outputs(1973) <= not (a or b);
    layer0_outputs(1974) <= not a or b;
    layer0_outputs(1975) <= not a;
    layer0_outputs(1976) <= b;
    layer0_outputs(1977) <= a or b;
    layer0_outputs(1978) <= not (a or b);
    layer0_outputs(1979) <= not (a or b);
    layer0_outputs(1980) <= a or b;
    layer0_outputs(1981) <= not b or a;
    layer0_outputs(1982) <= a and not b;
    layer0_outputs(1983) <= not a;
    layer0_outputs(1984) <= not (a or b);
    layer0_outputs(1985) <= a and not b;
    layer0_outputs(1986) <= a or b;
    layer0_outputs(1987) <= not a;
    layer0_outputs(1988) <= not a;
    layer0_outputs(1989) <= not (a or b);
    layer0_outputs(1990) <= not (a xor b);
    layer0_outputs(1991) <= not (a or b);
    layer0_outputs(1992) <= a and not b;
    layer0_outputs(1993) <= not a or b;
    layer0_outputs(1994) <= a;
    layer0_outputs(1995) <= a and b;
    layer0_outputs(1996) <= a or b;
    layer0_outputs(1997) <= a and not b;
    layer0_outputs(1998) <= not (a xor b);
    layer0_outputs(1999) <= a or b;
    layer0_outputs(2000) <= not (a or b);
    layer0_outputs(2001) <= a and b;
    layer0_outputs(2002) <= not a;
    layer0_outputs(2003) <= b;
    layer0_outputs(2004) <= a or b;
    layer0_outputs(2005) <= a or b;
    layer0_outputs(2006) <= a or b;
    layer0_outputs(2007) <= not (a or b);
    layer0_outputs(2008) <= b and not a;
    layer0_outputs(2009) <= not a;
    layer0_outputs(2010) <= not (a or b);
    layer0_outputs(2011) <= a and b;
    layer0_outputs(2012) <= a;
    layer0_outputs(2013) <= not a;
    layer0_outputs(2014) <= b and not a;
    layer0_outputs(2015) <= not a or b;
    layer0_outputs(2016) <= not (a xor b);
    layer0_outputs(2017) <= not (a xor b);
    layer0_outputs(2018) <= not (a or b);
    layer0_outputs(2019) <= not (a xor b);
    layer0_outputs(2020) <= not a;
    layer0_outputs(2021) <= not a;
    layer0_outputs(2022) <= a or b;
    layer0_outputs(2023) <= not (a xor b);
    layer0_outputs(2024) <= not (a or b);
    layer0_outputs(2025) <= a or b;
    layer0_outputs(2026) <= not b;
    layer0_outputs(2027) <= a or b;
    layer0_outputs(2028) <= not a or b;
    layer0_outputs(2029) <= 1'b0;
    layer0_outputs(2030) <= not (a or b);
    layer0_outputs(2031) <= a and not b;
    layer0_outputs(2032) <= not b or a;
    layer0_outputs(2033) <= not a;
    layer0_outputs(2034) <= not b;
    layer0_outputs(2035) <= not a or b;
    layer0_outputs(2036) <= a or b;
    layer0_outputs(2037) <= not (a xor b);
    layer0_outputs(2038) <= a or b;
    layer0_outputs(2039) <= b;
    layer0_outputs(2040) <= a xor b;
    layer0_outputs(2041) <= not (a or b);
    layer0_outputs(2042) <= a or b;
    layer0_outputs(2043) <= not a or b;
    layer0_outputs(2044) <= a xor b;
    layer0_outputs(2045) <= not (a xor b);
    layer0_outputs(2046) <= a or b;
    layer0_outputs(2047) <= not a or b;
    layer0_outputs(2048) <= not a;
    layer0_outputs(2049) <= b and not a;
    layer0_outputs(2050) <= b;
    layer0_outputs(2051) <= b and not a;
    layer0_outputs(2052) <= a xor b;
    layer0_outputs(2053) <= not (a or b);
    layer0_outputs(2054) <= a and not b;
    layer0_outputs(2055) <= a;
    layer0_outputs(2056) <= not (a or b);
    layer0_outputs(2057) <= not (a xor b);
    layer0_outputs(2058) <= not a;
    layer0_outputs(2059) <= not a or b;
    layer0_outputs(2060) <= b and not a;
    layer0_outputs(2061) <= not (a xor b);
    layer0_outputs(2062) <= not a or b;
    layer0_outputs(2063) <= not (a xor b);
    layer0_outputs(2064) <= not b;
    layer0_outputs(2065) <= not (a or b);
    layer0_outputs(2066) <= not (a or b);
    layer0_outputs(2067) <= b;
    layer0_outputs(2068) <= b and not a;
    layer0_outputs(2069) <= a;
    layer0_outputs(2070) <= a;
    layer0_outputs(2071) <= not a or b;
    layer0_outputs(2072) <= b and not a;
    layer0_outputs(2073) <= not b;
    layer0_outputs(2074) <= not (a xor b);
    layer0_outputs(2075) <= a xor b;
    layer0_outputs(2076) <= 1'b1;
    layer0_outputs(2077) <= a and not b;
    layer0_outputs(2078) <= a or b;
    layer0_outputs(2079) <= not a or b;
    layer0_outputs(2080) <= a;
    layer0_outputs(2081) <= not (a xor b);
    layer0_outputs(2082) <= a or b;
    layer0_outputs(2083) <= a xor b;
    layer0_outputs(2084) <= a or b;
    layer0_outputs(2085) <= b and not a;
    layer0_outputs(2086) <= not (a or b);
    layer0_outputs(2087) <= not a;
    layer0_outputs(2088) <= a xor b;
    layer0_outputs(2089) <= not a or b;
    layer0_outputs(2090) <= a;
    layer0_outputs(2091) <= b;
    layer0_outputs(2092) <= b and not a;
    layer0_outputs(2093) <= a or b;
    layer0_outputs(2094) <= not a or b;
    layer0_outputs(2095) <= not a;
    layer0_outputs(2096) <= not (a or b);
    layer0_outputs(2097) <= a and not b;
    layer0_outputs(2098) <= not a;
    layer0_outputs(2099) <= a or b;
    layer0_outputs(2100) <= not (a or b);
    layer0_outputs(2101) <= not (a or b);
    layer0_outputs(2102) <= 1'b0;
    layer0_outputs(2103) <= b and not a;
    layer0_outputs(2104) <= b and not a;
    layer0_outputs(2105) <= a;
    layer0_outputs(2106) <= a or b;
    layer0_outputs(2107) <= 1'b1;
    layer0_outputs(2108) <= 1'b0;
    layer0_outputs(2109) <= a and not b;
    layer0_outputs(2110) <= a or b;
    layer0_outputs(2111) <= not (a or b);
    layer0_outputs(2112) <= not a or b;
    layer0_outputs(2113) <= not (a or b);
    layer0_outputs(2114) <= not a;
    layer0_outputs(2115) <= a and not b;
    layer0_outputs(2116) <= not (a and b);
    layer0_outputs(2117) <= a or b;
    layer0_outputs(2118) <= not b;
    layer0_outputs(2119) <= a and not b;
    layer0_outputs(2120) <= not b;
    layer0_outputs(2121) <= not b;
    layer0_outputs(2122) <= a xor b;
    layer0_outputs(2123) <= a xor b;
    layer0_outputs(2124) <= a;
    layer0_outputs(2125) <= a and not b;
    layer0_outputs(2126) <= not a;
    layer0_outputs(2127) <= not (a or b);
    layer0_outputs(2128) <= a and not b;
    layer0_outputs(2129) <= not b;
    layer0_outputs(2130) <= not a;
    layer0_outputs(2131) <= not b or a;
    layer0_outputs(2132) <= not (a xor b);
    layer0_outputs(2133) <= a or b;
    layer0_outputs(2134) <= a;
    layer0_outputs(2135) <= not b;
    layer0_outputs(2136) <= a;
    layer0_outputs(2137) <= a xor b;
    layer0_outputs(2138) <= a or b;
    layer0_outputs(2139) <= not (a or b);
    layer0_outputs(2140) <= b and not a;
    layer0_outputs(2141) <= not a;
    layer0_outputs(2142) <= not (a xor b);
    layer0_outputs(2143) <= a and b;
    layer0_outputs(2144) <= 1'b1;
    layer0_outputs(2145) <= a xor b;
    layer0_outputs(2146) <= not a or b;
    layer0_outputs(2147) <= not b or a;
    layer0_outputs(2148) <= not a or b;
    layer0_outputs(2149) <= b and not a;
    layer0_outputs(2150) <= not a;
    layer0_outputs(2151) <= a or b;
    layer0_outputs(2152) <= not a or b;
    layer0_outputs(2153) <= not b;
    layer0_outputs(2154) <= not (a or b);
    layer0_outputs(2155) <= a xor b;
    layer0_outputs(2156) <= not (a or b);
    layer0_outputs(2157) <= not (a or b);
    layer0_outputs(2158) <= not b or a;
    layer0_outputs(2159) <= b;
    layer0_outputs(2160) <= a or b;
    layer0_outputs(2161) <= a and not b;
    layer0_outputs(2162) <= not a or b;
    layer0_outputs(2163) <= not (a or b);
    layer0_outputs(2164) <= not (a or b);
    layer0_outputs(2165) <= a xor b;
    layer0_outputs(2166) <= not b;
    layer0_outputs(2167) <= not (a or b);
    layer0_outputs(2168) <= a xor b;
    layer0_outputs(2169) <= not (a or b);
    layer0_outputs(2170) <= not b or a;
    layer0_outputs(2171) <= not a;
    layer0_outputs(2172) <= not b or a;
    layer0_outputs(2173) <= a and not b;
    layer0_outputs(2174) <= a or b;
    layer0_outputs(2175) <= a or b;
    layer0_outputs(2176) <= a or b;
    layer0_outputs(2177) <= a;
    layer0_outputs(2178) <= a;
    layer0_outputs(2179) <= not (a xor b);
    layer0_outputs(2180) <= a xor b;
    layer0_outputs(2181) <= b;
    layer0_outputs(2182) <= not b;
    layer0_outputs(2183) <= not (a and b);
    layer0_outputs(2184) <= not (a xor b);
    layer0_outputs(2185) <= not b or a;
    layer0_outputs(2186) <= not a;
    layer0_outputs(2187) <= b and not a;
    layer0_outputs(2188) <= a xor b;
    layer0_outputs(2189) <= b;
    layer0_outputs(2190) <= not (a xor b);
    layer0_outputs(2191) <= a xor b;
    layer0_outputs(2192) <= not (a or b);
    layer0_outputs(2193) <= a and not b;
    layer0_outputs(2194) <= b;
    layer0_outputs(2195) <= 1'b0;
    layer0_outputs(2196) <= b and not a;
    layer0_outputs(2197) <= not b;
    layer0_outputs(2198) <= a or b;
    layer0_outputs(2199) <= a or b;
    layer0_outputs(2200) <= a;
    layer0_outputs(2201) <= a or b;
    layer0_outputs(2202) <= not (a or b);
    layer0_outputs(2203) <= not (a or b);
    layer0_outputs(2204) <= a or b;
    layer0_outputs(2205) <= a and b;
    layer0_outputs(2206) <= not (a or b);
    layer0_outputs(2207) <= not (a or b);
    layer0_outputs(2208) <= not (a or b);
    layer0_outputs(2209) <= not (a or b);
    layer0_outputs(2210) <= not (a and b);
    layer0_outputs(2211) <= not (a or b);
    layer0_outputs(2212) <= a or b;
    layer0_outputs(2213) <= a or b;
    layer0_outputs(2214) <= a or b;
    layer0_outputs(2215) <= not a or b;
    layer0_outputs(2216) <= not b or a;
    layer0_outputs(2217) <= not b;
    layer0_outputs(2218) <= a and not b;
    layer0_outputs(2219) <= not b;
    layer0_outputs(2220) <= b;
    layer0_outputs(2221) <= a and not b;
    layer0_outputs(2222) <= 1'b1;
    layer0_outputs(2223) <= a;
    layer0_outputs(2224) <= 1'b0;
    layer0_outputs(2225) <= b and not a;
    layer0_outputs(2226) <= a xor b;
    layer0_outputs(2227) <= a or b;
    layer0_outputs(2228) <= not (a and b);
    layer0_outputs(2229) <= not (a or b);
    layer0_outputs(2230) <= not b or a;
    layer0_outputs(2231) <= a and not b;
    layer0_outputs(2232) <= a or b;
    layer0_outputs(2233) <= not (a or b);
    layer0_outputs(2234) <= a and not b;
    layer0_outputs(2235) <= a;
    layer0_outputs(2236) <= b;
    layer0_outputs(2237) <= b;
    layer0_outputs(2238) <= not (a or b);
    layer0_outputs(2239) <= a and b;
    layer0_outputs(2240) <= not (a and b);
    layer0_outputs(2241) <= not b;
    layer0_outputs(2242) <= not (a or b);
    layer0_outputs(2243) <= not (a or b);
    layer0_outputs(2244) <= not (a or b);
    layer0_outputs(2245) <= not (a xor b);
    layer0_outputs(2246) <= not b or a;
    layer0_outputs(2247) <= b and not a;
    layer0_outputs(2248) <= a or b;
    layer0_outputs(2249) <= not b;
    layer0_outputs(2250) <= not (a or b);
    layer0_outputs(2251) <= 1'b1;
    layer0_outputs(2252) <= not a or b;
    layer0_outputs(2253) <= not (a or b);
    layer0_outputs(2254) <= b;
    layer0_outputs(2255) <= a or b;
    layer0_outputs(2256) <= not (a or b);
    layer0_outputs(2257) <= a or b;
    layer0_outputs(2258) <= not a or b;
    layer0_outputs(2259) <= b;
    layer0_outputs(2260) <= a or b;
    layer0_outputs(2261) <= a or b;
    layer0_outputs(2262) <= b;
    layer0_outputs(2263) <= a or b;
    layer0_outputs(2264) <= a xor b;
    layer0_outputs(2265) <= a or b;
    layer0_outputs(2266) <= 1'b1;
    layer0_outputs(2267) <= not b;
    layer0_outputs(2268) <= a or b;
    layer0_outputs(2269) <= a xor b;
    layer0_outputs(2270) <= not a or b;
    layer0_outputs(2271) <= not (a or b);
    layer0_outputs(2272) <= not (a xor b);
    layer0_outputs(2273) <= not (a xor b);
    layer0_outputs(2274) <= a or b;
    layer0_outputs(2275) <= not (a or b);
    layer0_outputs(2276) <= a or b;
    layer0_outputs(2277) <= a xor b;
    layer0_outputs(2278) <= a;
    layer0_outputs(2279) <= not a or b;
    layer0_outputs(2280) <= not a;
    layer0_outputs(2281) <= not (a or b);
    layer0_outputs(2282) <= a xor b;
    layer0_outputs(2283) <= b;
    layer0_outputs(2284) <= a or b;
    layer0_outputs(2285) <= not b;
    layer0_outputs(2286) <= not a or b;
    layer0_outputs(2287) <= not (a or b);
    layer0_outputs(2288) <= not (a or b);
    layer0_outputs(2289) <= not a or b;
    layer0_outputs(2290) <= b;
    layer0_outputs(2291) <= a xor b;
    layer0_outputs(2292) <= not (a xor b);
    layer0_outputs(2293) <= a or b;
    layer0_outputs(2294) <= not a;
    layer0_outputs(2295) <= not b;
    layer0_outputs(2296) <= not (a or b);
    layer0_outputs(2297) <= a or b;
    layer0_outputs(2298) <= a or b;
    layer0_outputs(2299) <= a or b;
    layer0_outputs(2300) <= not a;
    layer0_outputs(2301) <= not (a or b);
    layer0_outputs(2302) <= a or b;
    layer0_outputs(2303) <= not (a xor b);
    layer0_outputs(2304) <= not (a xor b);
    layer0_outputs(2305) <= b;
    layer0_outputs(2306) <= b;
    layer0_outputs(2307) <= a;
    layer0_outputs(2308) <= not (a or b);
    layer0_outputs(2309) <= not (a or b);
    layer0_outputs(2310) <= b and not a;
    layer0_outputs(2311) <= a xor b;
    layer0_outputs(2312) <= not b or a;
    layer0_outputs(2313) <= b;
    layer0_outputs(2314) <= not (a or b);
    layer0_outputs(2315) <= b;
    layer0_outputs(2316) <= a or b;
    layer0_outputs(2317) <= not (a or b);
    layer0_outputs(2318) <= a xor b;
    layer0_outputs(2319) <= 1'b1;
    layer0_outputs(2320) <= a;
    layer0_outputs(2321) <= not b or a;
    layer0_outputs(2322) <= a or b;
    layer0_outputs(2323) <= not a;
    layer0_outputs(2324) <= a xor b;
    layer0_outputs(2325) <= a;
    layer0_outputs(2326) <= a;
    layer0_outputs(2327) <= a or b;
    layer0_outputs(2328) <= 1'b0;
    layer0_outputs(2329) <= b and not a;
    layer0_outputs(2330) <= not (a or b);
    layer0_outputs(2331) <= a;
    layer0_outputs(2332) <= not (a and b);
    layer0_outputs(2333) <= not a or b;
    layer0_outputs(2334) <= a xor b;
    layer0_outputs(2335) <= a or b;
    layer0_outputs(2336) <= a;
    layer0_outputs(2337) <= not b or a;
    layer0_outputs(2338) <= not b or a;
    layer0_outputs(2339) <= a xor b;
    layer0_outputs(2340) <= not b;
    layer0_outputs(2341) <= not a;
    layer0_outputs(2342) <= a;
    layer0_outputs(2343) <= not a;
    layer0_outputs(2344) <= a and not b;
    layer0_outputs(2345) <= not a or b;
    layer0_outputs(2346) <= b;
    layer0_outputs(2347) <= not a;
    layer0_outputs(2348) <= b and not a;
    layer0_outputs(2349) <= not b;
    layer0_outputs(2350) <= a xor b;
    layer0_outputs(2351) <= a or b;
    layer0_outputs(2352) <= not (a or b);
    layer0_outputs(2353) <= a xor b;
    layer0_outputs(2354) <= not a;
    layer0_outputs(2355) <= a and not b;
    layer0_outputs(2356) <= not b;
    layer0_outputs(2357) <= b;
    layer0_outputs(2358) <= not a;
    layer0_outputs(2359) <= not (a xor b);
    layer0_outputs(2360) <= a or b;
    layer0_outputs(2361) <= a xor b;
    layer0_outputs(2362) <= not b;
    layer0_outputs(2363) <= a or b;
    layer0_outputs(2364) <= a;
    layer0_outputs(2365) <= a or b;
    layer0_outputs(2366) <= a and b;
    layer0_outputs(2367) <= not (a or b);
    layer0_outputs(2368) <= a;
    layer0_outputs(2369) <= not b;
    layer0_outputs(2370) <= not b or a;
    layer0_outputs(2371) <= not b or a;
    layer0_outputs(2372) <= a xor b;
    layer0_outputs(2373) <= not a;
    layer0_outputs(2374) <= a xor b;
    layer0_outputs(2375) <= b;
    layer0_outputs(2376) <= a or b;
    layer0_outputs(2377) <= a;
    layer0_outputs(2378) <= 1'b1;
    layer0_outputs(2379) <= a;
    layer0_outputs(2380) <= a or b;
    layer0_outputs(2381) <= a and not b;
    layer0_outputs(2382) <= not (a or b);
    layer0_outputs(2383) <= a xor b;
    layer0_outputs(2384) <= a or b;
    layer0_outputs(2385) <= a or b;
    layer0_outputs(2386) <= not a or b;
    layer0_outputs(2387) <= a xor b;
    layer0_outputs(2388) <= not (a xor b);
    layer0_outputs(2389) <= not (a and b);
    layer0_outputs(2390) <= a or b;
    layer0_outputs(2391) <= not (a or b);
    layer0_outputs(2392) <= not b;
    layer0_outputs(2393) <= b and not a;
    layer0_outputs(2394) <= a and not b;
    layer0_outputs(2395) <= not (a or b);
    layer0_outputs(2396) <= a xor b;
    layer0_outputs(2397) <= not (a or b);
    layer0_outputs(2398) <= b;
    layer0_outputs(2399) <= a;
    layer0_outputs(2400) <= a or b;
    layer0_outputs(2401) <= b;
    layer0_outputs(2402) <= not (a or b);
    layer0_outputs(2403) <= a or b;
    layer0_outputs(2404) <= not (a xor b);
    layer0_outputs(2405) <= not a or b;
    layer0_outputs(2406) <= a and not b;
    layer0_outputs(2407) <= a or b;
    layer0_outputs(2408) <= not a or b;
    layer0_outputs(2409) <= not a;
    layer0_outputs(2410) <= b;
    layer0_outputs(2411) <= not a;
    layer0_outputs(2412) <= not (a xor b);
    layer0_outputs(2413) <= a and not b;
    layer0_outputs(2414) <= a or b;
    layer0_outputs(2415) <= not (a xor b);
    layer0_outputs(2416) <= not b;
    layer0_outputs(2417) <= not a;
    layer0_outputs(2418) <= b;
    layer0_outputs(2419) <= not (a xor b);
    layer0_outputs(2420) <= not (a xor b);
    layer0_outputs(2421) <= a xor b;
    layer0_outputs(2422) <= not b;
    layer0_outputs(2423) <= a and not b;
    layer0_outputs(2424) <= a xor b;
    layer0_outputs(2425) <= b;
    layer0_outputs(2426) <= not a or b;
    layer0_outputs(2427) <= a or b;
    layer0_outputs(2428) <= b;
    layer0_outputs(2429) <= not (a or b);
    layer0_outputs(2430) <= a;
    layer0_outputs(2431) <= not b;
    layer0_outputs(2432) <= not a;
    layer0_outputs(2433) <= a or b;
    layer0_outputs(2434) <= a or b;
    layer0_outputs(2435) <= not b;
    layer0_outputs(2436) <= a and b;
    layer0_outputs(2437) <= 1'b0;
    layer0_outputs(2438) <= not (a xor b);
    layer0_outputs(2439) <= not a;
    layer0_outputs(2440) <= b and not a;
    layer0_outputs(2441) <= a xor b;
    layer0_outputs(2442) <= b and not a;
    layer0_outputs(2443) <= a or b;
    layer0_outputs(2444) <= not (a or b);
    layer0_outputs(2445) <= not (a or b);
    layer0_outputs(2446) <= a xor b;
    layer0_outputs(2447) <= a and not b;
    layer0_outputs(2448) <= b;
    layer0_outputs(2449) <= a or b;
    layer0_outputs(2450) <= not (a or b);
    layer0_outputs(2451) <= not (a or b);
    layer0_outputs(2452) <= not (a xor b);
    layer0_outputs(2453) <= not (a or b);
    layer0_outputs(2454) <= 1'b0;
    layer0_outputs(2455) <= not (a xor b);
    layer0_outputs(2456) <= a and not b;
    layer0_outputs(2457) <= b and not a;
    layer0_outputs(2458) <= b and not a;
    layer0_outputs(2459) <= not b;
    layer0_outputs(2460) <= not (a or b);
    layer0_outputs(2461) <= not (a or b);
    layer0_outputs(2462) <= a or b;
    layer0_outputs(2463) <= not b;
    layer0_outputs(2464) <= not b;
    layer0_outputs(2465) <= b and not a;
    layer0_outputs(2466) <= b;
    layer0_outputs(2467) <= not b or a;
    layer0_outputs(2468) <= not (a or b);
    layer0_outputs(2469) <= not b or a;
    layer0_outputs(2470) <= a or b;
    layer0_outputs(2471) <= not (a or b);
    layer0_outputs(2472) <= a;
    layer0_outputs(2473) <= b;
    layer0_outputs(2474) <= a or b;
    layer0_outputs(2475) <= b and not a;
    layer0_outputs(2476) <= b;
    layer0_outputs(2477) <= a and not b;
    layer0_outputs(2478) <= a xor b;
    layer0_outputs(2479) <= not (a or b);
    layer0_outputs(2480) <= a;
    layer0_outputs(2481) <= a or b;
    layer0_outputs(2482) <= a or b;
    layer0_outputs(2483) <= not b;
    layer0_outputs(2484) <= not b or a;
    layer0_outputs(2485) <= not b or a;
    layer0_outputs(2486) <= b and not a;
    layer0_outputs(2487) <= a or b;
    layer0_outputs(2488) <= a and not b;
    layer0_outputs(2489) <= b and not a;
    layer0_outputs(2490) <= not (a xor b);
    layer0_outputs(2491) <= b;
    layer0_outputs(2492) <= not b or a;
    layer0_outputs(2493) <= not (a xor b);
    layer0_outputs(2494) <= a or b;
    layer0_outputs(2495) <= not b;
    layer0_outputs(2496) <= a and not b;
    layer0_outputs(2497) <= a or b;
    layer0_outputs(2498) <= not (a or b);
    layer0_outputs(2499) <= a;
    layer0_outputs(2500) <= not b or a;
    layer0_outputs(2501) <= not a or b;
    layer0_outputs(2502) <= b;
    layer0_outputs(2503) <= not (a xor b);
    layer0_outputs(2504) <= not b;
    layer0_outputs(2505) <= not (a xor b);
    layer0_outputs(2506) <= not (a or b);
    layer0_outputs(2507) <= b and not a;
    layer0_outputs(2508) <= b;
    layer0_outputs(2509) <= not b or a;
    layer0_outputs(2510) <= a or b;
    layer0_outputs(2511) <= a xor b;
    layer0_outputs(2512) <= not (a xor b);
    layer0_outputs(2513) <= a;
    layer0_outputs(2514) <= not (a or b);
    layer0_outputs(2515) <= a xor b;
    layer0_outputs(2516) <= a;
    layer0_outputs(2517) <= a or b;
    layer0_outputs(2518) <= not b or a;
    layer0_outputs(2519) <= 1'b1;
    layer0_outputs(2520) <= a and not b;
    layer0_outputs(2521) <= not (a or b);
    layer0_outputs(2522) <= a or b;
    layer0_outputs(2523) <= a or b;
    layer0_outputs(2524) <= b;
    layer0_outputs(2525) <= not (a xor b);
    layer0_outputs(2526) <= not b or a;
    layer0_outputs(2527) <= a;
    layer0_outputs(2528) <= b;
    layer0_outputs(2529) <= a;
    layer0_outputs(2530) <= a xor b;
    layer0_outputs(2531) <= not a or b;
    layer0_outputs(2532) <= a;
    layer0_outputs(2533) <= not (a or b);
    layer0_outputs(2534) <= b and not a;
    layer0_outputs(2535) <= a or b;
    layer0_outputs(2536) <= not (a xor b);
    layer0_outputs(2537) <= not a;
    layer0_outputs(2538) <= b and not a;
    layer0_outputs(2539) <= b;
    layer0_outputs(2540) <= a;
    layer0_outputs(2541) <= not (a xor b);
    layer0_outputs(2542) <= not (a or b);
    layer0_outputs(2543) <= not a or b;
    layer0_outputs(2544) <= a or b;
    layer0_outputs(2545) <= b and not a;
    layer0_outputs(2546) <= not (a xor b);
    layer0_outputs(2547) <= not a;
    layer0_outputs(2548) <= not (a xor b);
    layer0_outputs(2549) <= b and not a;
    layer0_outputs(2550) <= a;
    layer0_outputs(2551) <= a xor b;
    layer0_outputs(2552) <= a or b;
    layer0_outputs(2553) <= a and not b;
    layer0_outputs(2554) <= not a;
    layer0_outputs(2555) <= not b;
    layer0_outputs(2556) <= not a;
    layer0_outputs(2557) <= not b;
    layer0_outputs(2558) <= not b;
    layer0_outputs(2559) <= a and not b;
    outputs(0) <= a;
    outputs(1) <= a and b;
    outputs(2) <= not (a xor b);
    outputs(3) <= not b;
    outputs(4) <= a;
    outputs(5) <= a and not b;
    outputs(6) <= not b or a;
    outputs(7) <= not a or b;
    outputs(8) <= not (a xor b);
    outputs(9) <= not (a xor b);
    outputs(10) <= a;
    outputs(11) <= b;
    outputs(12) <= not (a or b);
    outputs(13) <= b;
    outputs(14) <= b and not a;
    outputs(15) <= not (a and b);
    outputs(16) <= a and b;
    outputs(17) <= b;
    outputs(18) <= not a;
    outputs(19) <= not (a xor b);
    outputs(20) <= not b;
    outputs(21) <= a xor b;
    outputs(22) <= not (a or b);
    outputs(23) <= not a;
    outputs(24) <= b;
    outputs(25) <= a;
    outputs(26) <= b;
    outputs(27) <= a;
    outputs(28) <= a and not b;
    outputs(29) <= not (a or b);
    outputs(30) <= not (a or b);
    outputs(31) <= b;
    outputs(32) <= not b;
    outputs(33) <= b;
    outputs(34) <= not (a xor b);
    outputs(35) <= b and not a;
    outputs(36) <= not b;
    outputs(37) <= a xor b;
    outputs(38) <= a xor b;
    outputs(39) <= not (a and b);
    outputs(40) <= not a;
    outputs(41) <= a;
    outputs(42) <= b;
    outputs(43) <= a xor b;
    outputs(44) <= b and not a;
    outputs(45) <= a;
    outputs(46) <= a and not b;
    outputs(47) <= not a;
    outputs(48) <= a;
    outputs(49) <= a or b;
    outputs(50) <= a and b;
    outputs(51) <= b;
    outputs(52) <= not b or a;
    outputs(53) <= not a;
    outputs(54) <= b;
    outputs(55) <= not b;
    outputs(56) <= a xor b;
    outputs(57) <= a xor b;
    outputs(58) <= a or b;
    outputs(59) <= not (a xor b);
    outputs(60) <= not (a and b);
    outputs(61) <= not (a xor b);
    outputs(62) <= not b;
    outputs(63) <= not (a and b);
    outputs(64) <= not a;
    outputs(65) <= b;
    outputs(66) <= not b;
    outputs(67) <= not b;
    outputs(68) <= not b;
    outputs(69) <= not (a or b);
    outputs(70) <= not b;
    outputs(71) <= b;
    outputs(72) <= b;
    outputs(73) <= not (a or b);
    outputs(74) <= b;
    outputs(75) <= not (a or b);
    outputs(76) <= not b;
    outputs(77) <= a;
    outputs(78) <= b and not a;
    outputs(79) <= not b;
    outputs(80) <= not a;
    outputs(81) <= a and b;
    outputs(82) <= a;
    outputs(83) <= a;
    outputs(84) <= not a or b;
    outputs(85) <= b and not a;
    outputs(86) <= a;
    outputs(87) <= not (a and b);
    outputs(88) <= not b;
    outputs(89) <= a and b;
    outputs(90) <= a and b;
    outputs(91) <= not a;
    outputs(92) <= a and b;
    outputs(93) <= b;
    outputs(94) <= not (a or b);
    outputs(95) <= b;
    outputs(96) <= not (a or b);
    outputs(97) <= not (a or b);
    outputs(98) <= a and b;
    outputs(99) <= a or b;
    outputs(100) <= b;
    outputs(101) <= b and not a;
    outputs(102) <= a;
    outputs(103) <= a;
    outputs(104) <= not (a xor b);
    outputs(105) <= b;
    outputs(106) <= not (a xor b);
    outputs(107) <= not a;
    outputs(108) <= a and b;
    outputs(109) <= a;
    outputs(110) <= a;
    outputs(111) <= a xor b;
    outputs(112) <= a;
    outputs(113) <= not a or b;
    outputs(114) <= a and not b;
    outputs(115) <= not (a and b);
    outputs(116) <= not b or a;
    outputs(117) <= not a;
    outputs(118) <= not (a xor b);
    outputs(119) <= not a;
    outputs(120) <= not (a or b);
    outputs(121) <= not (a and b);
    outputs(122) <= not (a and b);
    outputs(123) <= a;
    outputs(124) <= not a;
    outputs(125) <= not a;
    outputs(126) <= a or b;
    outputs(127) <= a;
    outputs(128) <= not a;
    outputs(129) <= not b;
    outputs(130) <= not (a and b);
    outputs(131) <= a xor b;
    outputs(132) <= b;
    outputs(133) <= a and b;
    outputs(134) <= a and b;
    outputs(135) <= a and not b;
    outputs(136) <= not (a and b);
    outputs(137) <= not b or a;
    outputs(138) <= not (a xor b);
    outputs(139) <= a and not b;
    outputs(140) <= not a or b;
    outputs(141) <= not b;
    outputs(142) <= a;
    outputs(143) <= not (a xor b);
    outputs(144) <= a xor b;
    outputs(145) <= not a;
    outputs(146) <= not b;
    outputs(147) <= a or b;
    outputs(148) <= not a;
    outputs(149) <= a xor b;
    outputs(150) <= a xor b;
    outputs(151) <= a;
    outputs(152) <= b;
    outputs(153) <= not b;
    outputs(154) <= a;
    outputs(155) <= b and not a;
    outputs(156) <= a or b;
    outputs(157) <= a;
    outputs(158) <= not b;
    outputs(159) <= not (a xor b);
    outputs(160) <= a or b;
    outputs(161) <= b and not a;
    outputs(162) <= a;
    outputs(163) <= not b or a;
    outputs(164) <= not (a xor b);
    outputs(165) <= a and b;
    outputs(166) <= a xor b;
    outputs(167) <= a and not b;
    outputs(168) <= a or b;
    outputs(169) <= not (a xor b);
    outputs(170) <= a and not b;
    outputs(171) <= not (a or b);
    outputs(172) <= a xor b;
    outputs(173) <= not a;
    outputs(174) <= a and b;
    outputs(175) <= not b;
    outputs(176) <= b;
    outputs(177) <= a and b;
    outputs(178) <= a;
    outputs(179) <= not (a or b);
    outputs(180) <= b and not a;
    outputs(181) <= a or b;
    outputs(182) <= a and b;
    outputs(183) <= b and not a;
    outputs(184) <= b;
    outputs(185) <= not b;
    outputs(186) <= a and b;
    outputs(187) <= a and not b;
    outputs(188) <= not (a and b);
    outputs(189) <= b and not a;
    outputs(190) <= not (a and b);
    outputs(191) <= not b;
    outputs(192) <= not a or b;
    outputs(193) <= a and not b;
    outputs(194) <= not (a xor b);
    outputs(195) <= a xor b;
    outputs(196) <= a and b;
    outputs(197) <= b;
    outputs(198) <= a;
    outputs(199) <= a;
    outputs(200) <= not (a xor b);
    outputs(201) <= b;
    outputs(202) <= a and b;
    outputs(203) <= b;
    outputs(204) <= not (a or b);
    outputs(205) <= not a;
    outputs(206) <= a;
    outputs(207) <= b and not a;
    outputs(208) <= not b;
    outputs(209) <= a;
    outputs(210) <= not b;
    outputs(211) <= b;
    outputs(212) <= a;
    outputs(213) <= not a or b;
    outputs(214) <= a and b;
    outputs(215) <= b;
    outputs(216) <= a;
    outputs(217) <= b;
    outputs(218) <= b;
    outputs(219) <= a xor b;
    outputs(220) <= a xor b;
    outputs(221) <= a and b;
    outputs(222) <= a and b;
    outputs(223) <= a and b;
    outputs(224) <= a;
    outputs(225) <= not (a or b);
    outputs(226) <= a xor b;
    outputs(227) <= a and b;
    outputs(228) <= b;
    outputs(229) <= not a;
    outputs(230) <= a;
    outputs(231) <= not a or b;
    outputs(232) <= not (a xor b);
    outputs(233) <= not (a and b);
    outputs(234) <= b;
    outputs(235) <= a;
    outputs(236) <= b;
    outputs(237) <= b;
    outputs(238) <= not (a xor b);
    outputs(239) <= not (a xor b);
    outputs(240) <= not (a or b);
    outputs(241) <= b;
    outputs(242) <= b;
    outputs(243) <= a and b;
    outputs(244) <= b;
    outputs(245) <= not b or a;
    outputs(246) <= not (a xor b);
    outputs(247) <= not b;
    outputs(248) <= b;
    outputs(249) <= not a or b;
    outputs(250) <= a;
    outputs(251) <= not a or b;
    outputs(252) <= not a;
    outputs(253) <= a and b;
    outputs(254) <= a;
    outputs(255) <= not (a or b);
    outputs(256) <= a and not b;
    outputs(257) <= b and not a;
    outputs(258) <= a and not b;
    outputs(259) <= a and b;
    outputs(260) <= a and not b;
    outputs(261) <= not (a or b);
    outputs(262) <= a and b;
    outputs(263) <= b and not a;
    outputs(264) <= b and not a;
    outputs(265) <= a and not b;
    outputs(266) <= a and not b;
    outputs(267) <= not b;
    outputs(268) <= a and b;
    outputs(269) <= b;
    outputs(270) <= a and not b;
    outputs(271) <= a and not b;
    outputs(272) <= a and b;
    outputs(273) <= a and b;
    outputs(274) <= b and not a;
    outputs(275) <= not (a or b);
    outputs(276) <= a and not b;
    outputs(277) <= a and not b;
    outputs(278) <= b and not a;
    outputs(279) <= not b;
    outputs(280) <= a and not b;
    outputs(281) <= a;
    outputs(282) <= a;
    outputs(283) <= not a;
    outputs(284) <= a;
    outputs(285) <= a and b;
    outputs(286) <= b;
    outputs(287) <= not b;
    outputs(288) <= a and b;
    outputs(289) <= not (a or b);
    outputs(290) <= not b;
    outputs(291) <= a;
    outputs(292) <= b;
    outputs(293) <= a and not b;
    outputs(294) <= not (a or b);
    outputs(295) <= a and b;
    outputs(296) <= b and not a;
    outputs(297) <= b and not a;
    outputs(298) <= b and not a;
    outputs(299) <= a and not b;
    outputs(300) <= not b;
    outputs(301) <= b and not a;
    outputs(302) <= a;
    outputs(303) <= a and b;
    outputs(304) <= a and b;
    outputs(305) <= a;
    outputs(306) <= a and not b;
    outputs(307) <= b and not a;
    outputs(308) <= not (a or b);
    outputs(309) <= a and not b;
    outputs(310) <= not (a or b);
    outputs(311) <= not b;
    outputs(312) <= a;
    outputs(313) <= a and not b;
    outputs(314) <= not (a or b);
    outputs(315) <= a and not b;
    outputs(316) <= a and b;
    outputs(317) <= not (a or b);
    outputs(318) <= not b or a;
    outputs(319) <= not (a or b);
    outputs(320) <= b and not a;
    outputs(321) <= a and b;
    outputs(322) <= b and not a;
    outputs(323) <= a and b;
    outputs(324) <= a and b;
    outputs(325) <= b and not a;
    outputs(326) <= a and not b;
    outputs(327) <= a and b;
    outputs(328) <= not (a or b);
    outputs(329) <= a;
    outputs(330) <= not (a or b);
    outputs(331) <= not b;
    outputs(332) <= a and not b;
    outputs(333) <= b and not a;
    outputs(334) <= a and not b;
    outputs(335) <= not b;
    outputs(336) <= b and not a;
    outputs(337) <= not (a or b);
    outputs(338) <= a and b;
    outputs(339) <= not (a xor b);
    outputs(340) <= b;
    outputs(341) <= not (a or b);
    outputs(342) <= not (a or b);
    outputs(343) <= b;
    outputs(344) <= b and not a;
    outputs(345) <= a and b;
    outputs(346) <= a and b;
    outputs(347) <= a;
    outputs(348) <= not (a or b);
    outputs(349) <= not (a or b);
    outputs(350) <= a and not b;
    outputs(351) <= a and b;
    outputs(352) <= a xor b;
    outputs(353) <= not (a or b);
    outputs(354) <= not (a or b);
    outputs(355) <= not (a or b);
    outputs(356) <= a and not b;
    outputs(357) <= not (a or b);
    outputs(358) <= a and b;
    outputs(359) <= not (a or b);
    outputs(360) <= a and b;
    outputs(361) <= not b or a;
    outputs(362) <= a and not b;
    outputs(363) <= a and not b;
    outputs(364) <= not a;
    outputs(365) <= not (a or b);
    outputs(366) <= not b;
    outputs(367) <= a and b;
    outputs(368) <= not (a or b);
    outputs(369) <= not b or a;
    outputs(370) <= b and not a;
    outputs(371) <= 1'b0;
    outputs(372) <= not b;
    outputs(373) <= a;
    outputs(374) <= not (a or b);
    outputs(375) <= a and b;
    outputs(376) <= a and not b;
    outputs(377) <= b and not a;
    outputs(378) <= a and not b;
    outputs(379) <= a and b;
    outputs(380) <= 1'b0;
    outputs(381) <= b and not a;
    outputs(382) <= a and b;
    outputs(383) <= b and not a;
    outputs(384) <= b and not a;
    outputs(385) <= a and not b;
    outputs(386) <= a and b;
    outputs(387) <= b and not a;
    outputs(388) <= a and b;
    outputs(389) <= b and not a;
    outputs(390) <= b;
    outputs(391) <= not (a or b);
    outputs(392) <= not (a xor b);
    outputs(393) <= a;
    outputs(394) <= a and not b;
    outputs(395) <= not (a xor b);
    outputs(396) <= a and not b;
    outputs(397) <= a xor b;
    outputs(398) <= a and b;
    outputs(399) <= a and b;
    outputs(400) <= not (a or b);
    outputs(401) <= b and not a;
    outputs(402) <= a xor b;
    outputs(403) <= a and not b;
    outputs(404) <= a and not b;
    outputs(405) <= 1'b0;
    outputs(406) <= a and not b;
    outputs(407) <= not (a xor b);
    outputs(408) <= not (a xor b);
    outputs(409) <= not (a or b);
    outputs(410) <= b and not a;
    outputs(411) <= not (a or b);
    outputs(412) <= a and not b;
    outputs(413) <= not (a or b);
    outputs(414) <= a and b;
    outputs(415) <= b;
    outputs(416) <= a and b;
    outputs(417) <= a and b;
    outputs(418) <= 1'b0;
    outputs(419) <= a and b;
    outputs(420) <= b and not a;
    outputs(421) <= b and not a;
    outputs(422) <= a;
    outputs(423) <= not (a or b);
    outputs(424) <= a and not b;
    outputs(425) <= a and b;
    outputs(426) <= b;
    outputs(427) <= not b;
    outputs(428) <= not (a or b);
    outputs(429) <= not a;
    outputs(430) <= a xor b;
    outputs(431) <= b;
    outputs(432) <= a and b;
    outputs(433) <= not b;
    outputs(434) <= a and not b;
    outputs(435) <= 1'b0;
    outputs(436) <= a and b;
    outputs(437) <= not a;
    outputs(438) <= b and not a;
    outputs(439) <= a and b;
    outputs(440) <= not (a or b);
    outputs(441) <= a;
    outputs(442) <= not (a or b);
    outputs(443) <= 1'b0;
    outputs(444) <= a and not b;
    outputs(445) <= b;
    outputs(446) <= b and not a;
    outputs(447) <= b and not a;
    outputs(448) <= b;
    outputs(449) <= a and not b;
    outputs(450) <= b and not a;
    outputs(451) <= a and b;
    outputs(452) <= a xor b;
    outputs(453) <= not b;
    outputs(454) <= a and b;
    outputs(455) <= not (a xor b);
    outputs(456) <= a and b;
    outputs(457) <= a and b;
    outputs(458) <= a and b;
    outputs(459) <= a or b;
    outputs(460) <= b and not a;
    outputs(461) <= not (a or b);
    outputs(462) <= 1'b0;
    outputs(463) <= a and b;
    outputs(464) <= not a;
    outputs(465) <= not (a or b);
    outputs(466) <= b and not a;
    outputs(467) <= b;
    outputs(468) <= a and b;
    outputs(469) <= b and not a;
    outputs(470) <= not (a or b);
    outputs(471) <= not (a or b);
    outputs(472) <= not (a xor b);
    outputs(473) <= a and not b;
    outputs(474) <= not (a or b);
    outputs(475) <= b and not a;
    outputs(476) <= a and not b;
    outputs(477) <= not (a or b);
    outputs(478) <= a and not b;
    outputs(479) <= a and b;
    outputs(480) <= not (a xor b);
    outputs(481) <= a xor b;
    outputs(482) <= b and not a;
    outputs(483) <= not (a or b);
    outputs(484) <= a and not b;
    outputs(485) <= b and not a;
    outputs(486) <= a and b;
    outputs(487) <= a and b;
    outputs(488) <= a or b;
    outputs(489) <= a and not b;
    outputs(490) <= a and b;
    outputs(491) <= 1'b0;
    outputs(492) <= a and not b;
    outputs(493) <= a xor b;
    outputs(494) <= not (a xor b);
    outputs(495) <= not (a or b);
    outputs(496) <= b;
    outputs(497) <= b and not a;
    outputs(498) <= a and not b;
    outputs(499) <= not a;
    outputs(500) <= a and b;
    outputs(501) <= a and b;
    outputs(502) <= a and not b;
    outputs(503) <= b and not a;
    outputs(504) <= a xor b;
    outputs(505) <= a and not b;
    outputs(506) <= not (a xor b);
    outputs(507) <= b and not a;
    outputs(508) <= a and b;
    outputs(509) <= b;
    outputs(510) <= not (a or b);
    outputs(511) <= a;
    outputs(512) <= b;
    outputs(513) <= b;
    outputs(514) <= not b or a;
    outputs(515) <= a and b;
    outputs(516) <= not (a xor b);
    outputs(517) <= not a or b;
    outputs(518) <= a and b;
    outputs(519) <= a and b;
    outputs(520) <= not a;
    outputs(521) <= not a;
    outputs(522) <= a and not b;
    outputs(523) <= a xor b;
    outputs(524) <= not b;
    outputs(525) <= not b;
    outputs(526) <= a or b;
    outputs(527) <= not (a or b);
    outputs(528) <= a;
    outputs(529) <= a;
    outputs(530) <= not b;
    outputs(531) <= b and not a;
    outputs(532) <= a and b;
    outputs(533) <= a and b;
    outputs(534) <= a xor b;
    outputs(535) <= not (a and b);
    outputs(536) <= a;
    outputs(537) <= not (a or b);
    outputs(538) <= a and not b;
    outputs(539) <= not a;
    outputs(540) <= a;
    outputs(541) <= not (a and b);
    outputs(542) <= not b;
    outputs(543) <= b and not a;
    outputs(544) <= not a;
    outputs(545) <= a or b;
    outputs(546) <= not b;
    outputs(547) <= not (a xor b);
    outputs(548) <= b;
    outputs(549) <= not a or b;
    outputs(550) <= a xor b;
    outputs(551) <= b;
    outputs(552) <= not (a xor b);
    outputs(553) <= not a;
    outputs(554) <= a xor b;
    outputs(555) <= b;
    outputs(556) <= not a or b;
    outputs(557) <= a or b;
    outputs(558) <= b and not a;
    outputs(559) <= b and not a;
    outputs(560) <= a;
    outputs(561) <= not a or b;
    outputs(562) <= not b;
    outputs(563) <= a and b;
    outputs(564) <= not a;
    outputs(565) <= a xor b;
    outputs(566) <= not b or a;
    outputs(567) <= a and not b;
    outputs(568) <= not (a or b);
    outputs(569) <= not a;
    outputs(570) <= not (a xor b);
    outputs(571) <= not b;
    outputs(572) <= a and not b;
    outputs(573) <= b;
    outputs(574) <= not (a and b);
    outputs(575) <= not b;
    outputs(576) <= not (a xor b);
    outputs(577) <= a and b;
    outputs(578) <= not (a xor b);
    outputs(579) <= not a or b;
    outputs(580) <= a xor b;
    outputs(581) <= a or b;
    outputs(582) <= not (a and b);
    outputs(583) <= not (a and b);
    outputs(584) <= a;
    outputs(585) <= not b;
    outputs(586) <= a and not b;
    outputs(587) <= a or b;
    outputs(588) <= not (a and b);
    outputs(589) <= not b or a;
    outputs(590) <= a;
    outputs(591) <= not b;
    outputs(592) <= not b or a;
    outputs(593) <= not b;
    outputs(594) <= a or b;
    outputs(595) <= not a;
    outputs(596) <= not b;
    outputs(597) <= not b or a;
    outputs(598) <= not a or b;
    outputs(599) <= not (a and b);
    outputs(600) <= not (a and b);
    outputs(601) <= not b;
    outputs(602) <= b and not a;
    outputs(603) <= a xor b;
    outputs(604) <= b;
    outputs(605) <= a;
    outputs(606) <= not b;
    outputs(607) <= not (a xor b);
    outputs(608) <= b;
    outputs(609) <= a and b;
    outputs(610) <= not b or a;
    outputs(611) <= not b;
    outputs(612) <= not b;
    outputs(613) <= not (a xor b);
    outputs(614) <= not b or a;
    outputs(615) <= not a or b;
    outputs(616) <= not b or a;
    outputs(617) <= b and not a;
    outputs(618) <= b;
    outputs(619) <= not b or a;
    outputs(620) <= b and not a;
    outputs(621) <= not b or a;
    outputs(622) <= a or b;
    outputs(623) <= b;
    outputs(624) <= not b or a;
    outputs(625) <= not b or a;
    outputs(626) <= not b or a;
    outputs(627) <= not (a xor b);
    outputs(628) <= b;
    outputs(629) <= a or b;
    outputs(630) <= b;
    outputs(631) <= not (a and b);
    outputs(632) <= a;
    outputs(633) <= b;
    outputs(634) <= not b;
    outputs(635) <= a;
    outputs(636) <= a or b;
    outputs(637) <= not (a and b);
    outputs(638) <= not (a xor b);
    outputs(639) <= a and b;
    outputs(640) <= a;
    outputs(641) <= not b or a;
    outputs(642) <= not b;
    outputs(643) <= not (a and b);
    outputs(644) <= not a;
    outputs(645) <= not a or b;
    outputs(646) <= not (a xor b);
    outputs(647) <= not a;
    outputs(648) <= not b;
    outputs(649) <= not (a and b);
    outputs(650) <= a or b;
    outputs(651) <= a or b;
    outputs(652) <= a and b;
    outputs(653) <= not b or a;
    outputs(654) <= a and b;
    outputs(655) <= not a or b;
    outputs(656) <= not b or a;
    outputs(657) <= a;
    outputs(658) <= not a or b;
    outputs(659) <= a or b;
    outputs(660) <= not (a xor b);
    outputs(661) <= a xor b;
    outputs(662) <= b and not a;
    outputs(663) <= b;
    outputs(664) <= not a or b;
    outputs(665) <= b and not a;
    outputs(666) <= a and b;
    outputs(667) <= not a;
    outputs(668) <= not b or a;
    outputs(669) <= not b or a;
    outputs(670) <= not a or b;
    outputs(671) <= a;
    outputs(672) <= a;
    outputs(673) <= not b;
    outputs(674) <= a;
    outputs(675) <= not b or a;
    outputs(676) <= not b or a;
    outputs(677) <= a and b;
    outputs(678) <= not b;
    outputs(679) <= b and not a;
    outputs(680) <= a xor b;
    outputs(681) <= a xor b;
    outputs(682) <= b;
    outputs(683) <= not (a and b);
    outputs(684) <= a;
    outputs(685) <= b;
    outputs(686) <= not a;
    outputs(687) <= a or b;
    outputs(688) <= not a or b;
    outputs(689) <= not a;
    outputs(690) <= a;
    outputs(691) <= a and not b;
    outputs(692) <= not a;
    outputs(693) <= b;
    outputs(694) <= a;
    outputs(695) <= not a;
    outputs(696) <= not a;
    outputs(697) <= not b;
    outputs(698) <= not b;
    outputs(699) <= not a;
    outputs(700) <= not b or a;
    outputs(701) <= not a;
    outputs(702) <= not a;
    outputs(703) <= not b or a;
    outputs(704) <= not b or a;
    outputs(705) <= a xor b;
    outputs(706) <= not b;
    outputs(707) <= not (a or b);
    outputs(708) <= not a;
    outputs(709) <= a and not b;
    outputs(710) <= a and b;
    outputs(711) <= a xor b;
    outputs(712) <= not (a and b);
    outputs(713) <= b and not a;
    outputs(714) <= not a or b;
    outputs(715) <= not a or b;
    outputs(716) <= not b;
    outputs(717) <= not (a or b);
    outputs(718) <= not b;
    outputs(719) <= a or b;
    outputs(720) <= a;
    outputs(721) <= not (a xor b);
    outputs(722) <= b;
    outputs(723) <= b;
    outputs(724) <= not b;
    outputs(725) <= a;
    outputs(726) <= not b;
    outputs(727) <= not b;
    outputs(728) <= a and b;
    outputs(729) <= a and not b;
    outputs(730) <= b and not a;
    outputs(731) <= a;
    outputs(732) <= not a;
    outputs(733) <= not b;
    outputs(734) <= not (a or b);
    outputs(735) <= not (a xor b);
    outputs(736) <= not a;
    outputs(737) <= not (a xor b);
    outputs(738) <= a;
    outputs(739) <= not a;
    outputs(740) <= not (a xor b);
    outputs(741) <= not b;
    outputs(742) <= a;
    outputs(743) <= b and not a;
    outputs(744) <= b;
    outputs(745) <= not (a and b);
    outputs(746) <= not b;
    outputs(747) <= b and not a;
    outputs(748) <= a and b;
    outputs(749) <= a and not b;
    outputs(750) <= a or b;
    outputs(751) <= not a;
    outputs(752) <= a;
    outputs(753) <= not (a xor b);
    outputs(754) <= a and b;
    outputs(755) <= not (a or b);
    outputs(756) <= not b;
    outputs(757) <= b and not a;
    outputs(758) <= not b or a;
    outputs(759) <= a;
    outputs(760) <= a and b;
    outputs(761) <= not (a and b);
    outputs(762) <= a or b;
    outputs(763) <= a;
    outputs(764) <= not a;
    outputs(765) <= a and not b;
    outputs(766) <= not (a xor b);
    outputs(767) <= b;
    outputs(768) <= a;
    outputs(769) <= b;
    outputs(770) <= a and not b;
    outputs(771) <= not b or a;
    outputs(772) <= not b;
    outputs(773) <= not (a or b);
    outputs(774) <= not (a xor b);
    outputs(775) <= a;
    outputs(776) <= a or b;
    outputs(777) <= b and not a;
    outputs(778) <= a and not b;
    outputs(779) <= a or b;
    outputs(780) <= not a;
    outputs(781) <= b;
    outputs(782) <= not (a or b);
    outputs(783) <= not b;
    outputs(784) <= a;
    outputs(785) <= a and b;
    outputs(786) <= a xor b;
    outputs(787) <= a xor b;
    outputs(788) <= a and b;
    outputs(789) <= not b or a;
    outputs(790) <= not b or a;
    outputs(791) <= b and not a;
    outputs(792) <= not b or a;
    outputs(793) <= not a;
    outputs(794) <= a;
    outputs(795) <= not (a or b);
    outputs(796) <= a and not b;
    outputs(797) <= not b;
    outputs(798) <= a;
    outputs(799) <= a and b;
    outputs(800) <= a and b;
    outputs(801) <= a;
    outputs(802) <= b and not a;
    outputs(803) <= a and not b;
    outputs(804) <= a;
    outputs(805) <= not (a and b);
    outputs(806) <= b and not a;
    outputs(807) <= a;
    outputs(808) <= a xor b;
    outputs(809) <= not a;
    outputs(810) <= not b;
    outputs(811) <= a;
    outputs(812) <= b;
    outputs(813) <= b;
    outputs(814) <= a and b;
    outputs(815) <= not b;
    outputs(816) <= not (a or b);
    outputs(817) <= a;
    outputs(818) <= a and not b;
    outputs(819) <= a and not b;
    outputs(820) <= not a;
    outputs(821) <= not a;
    outputs(822) <= a and b;
    outputs(823) <= a xor b;
    outputs(824) <= not a;
    outputs(825) <= a or b;
    outputs(826) <= a xor b;
    outputs(827) <= a;
    outputs(828) <= a xor b;
    outputs(829) <= b;
    outputs(830) <= a and not b;
    outputs(831) <= a xor b;
    outputs(832) <= not (a and b);
    outputs(833) <= not (a or b);
    outputs(834) <= a and not b;
    outputs(835) <= a or b;
    outputs(836) <= not a;
    outputs(837) <= not b or a;
    outputs(838) <= a;
    outputs(839) <= a and not b;
    outputs(840) <= b;
    outputs(841) <= b;
    outputs(842) <= not a;
    outputs(843) <= a and b;
    outputs(844) <= a;
    outputs(845) <= not (a xor b);
    outputs(846) <= a and b;
    outputs(847) <= a and not b;
    outputs(848) <= a and not b;
    outputs(849) <= a and b;
    outputs(850) <= a and b;
    outputs(851) <= not a;
    outputs(852) <= a;
    outputs(853) <= not (a and b);
    outputs(854) <= a and not b;
    outputs(855) <= a xor b;
    outputs(856) <= not a or b;
    outputs(857) <= a and not b;
    outputs(858) <= b;
    outputs(859) <= a and b;
    outputs(860) <= a and b;
    outputs(861) <= a and b;
    outputs(862) <= a or b;
    outputs(863) <= not (a or b);
    outputs(864) <= not a or b;
    outputs(865) <= not (a xor b);
    outputs(866) <= a xor b;
    outputs(867) <= a xor b;
    outputs(868) <= a and not b;
    outputs(869) <= b;
    outputs(870) <= not a;
    outputs(871) <= a;
    outputs(872) <= a xor b;
    outputs(873) <= a and not b;
    outputs(874) <= b;
    outputs(875) <= a;
    outputs(876) <= not (a or b);
    outputs(877) <= a and b;
    outputs(878) <= a and b;
    outputs(879) <= not (a or b);
    outputs(880) <= b and not a;
    outputs(881) <= a and b;
    outputs(882) <= a;
    outputs(883) <= not a;
    outputs(884) <= b and not a;
    outputs(885) <= not a or b;
    outputs(886) <= a xor b;
    outputs(887) <= not (a or b);
    outputs(888) <= b;
    outputs(889) <= not (a or b);
    outputs(890) <= a;
    outputs(891) <= a or b;
    outputs(892) <= not a or b;
    outputs(893) <= a xor b;
    outputs(894) <= a;
    outputs(895) <= not a;
    outputs(896) <= a and b;
    outputs(897) <= b;
    outputs(898) <= a;
    outputs(899) <= not (a xor b);
    outputs(900) <= b;
    outputs(901) <= a;
    outputs(902) <= a;
    outputs(903) <= not b;
    outputs(904) <= b;
    outputs(905) <= a and not b;
    outputs(906) <= b;
    outputs(907) <= a and not b;
    outputs(908) <= not b;
    outputs(909) <= a and b;
    outputs(910) <= not a;
    outputs(911) <= b;
    outputs(912) <= a and not b;
    outputs(913) <= b;
    outputs(914) <= not b;
    outputs(915) <= not b;
    outputs(916) <= not (a xor b);
    outputs(917) <= a and not b;
    outputs(918) <= not (a and b);
    outputs(919) <= not b;
    outputs(920) <= not (a xor b);
    outputs(921) <= a xor b;
    outputs(922) <= not a;
    outputs(923) <= not b;
    outputs(924) <= not (a or b);
    outputs(925) <= not (a xor b);
    outputs(926) <= b;
    outputs(927) <= not (a or b);
    outputs(928) <= not b;
    outputs(929) <= b and not a;
    outputs(930) <= not b;
    outputs(931) <= a or b;
    outputs(932) <= not (a and b);
    outputs(933) <= b;
    outputs(934) <= not (a and b);
    outputs(935) <= a and not b;
    outputs(936) <= a;
    outputs(937) <= b;
    outputs(938) <= not a;
    outputs(939) <= a xor b;
    outputs(940) <= a and not b;
    outputs(941) <= not a or b;
    outputs(942) <= not a or b;
    outputs(943) <= b;
    outputs(944) <= a;
    outputs(945) <= not b;
    outputs(946) <= b and not a;
    outputs(947) <= a and not b;
    outputs(948) <= b;
    outputs(949) <= not (a or b);
    outputs(950) <= a xor b;
    outputs(951) <= b;
    outputs(952) <= not (a or b);
    outputs(953) <= a or b;
    outputs(954) <= b and not a;
    outputs(955) <= a xor b;
    outputs(956) <= b and not a;
    outputs(957) <= not a;
    outputs(958) <= a and b;
    outputs(959) <= not (a or b);
    outputs(960) <= not (a or b);
    outputs(961) <= not b;
    outputs(962) <= not a;
    outputs(963) <= not (a or b);
    outputs(964) <= b;
    outputs(965) <= a and b;
    outputs(966) <= not a or b;
    outputs(967) <= not (a and b);
    outputs(968) <= not b;
    outputs(969) <= b and not a;
    outputs(970) <= b and not a;
    outputs(971) <= b and not a;
    outputs(972) <= not (a xor b);
    outputs(973) <= not a;
    outputs(974) <= a and not b;
    outputs(975) <= a and b;
    outputs(976) <= not (a or b);
    outputs(977) <= a;
    outputs(978) <= not b;
    outputs(979) <= a xor b;
    outputs(980) <= a xor b;
    outputs(981) <= a and not b;
    outputs(982) <= a and b;
    outputs(983) <= not b or a;
    outputs(984) <= a and b;
    outputs(985) <= not b;
    outputs(986) <= a and not b;
    outputs(987) <= not (a or b);
    outputs(988) <= not b;
    outputs(989) <= b and not a;
    outputs(990) <= b;
    outputs(991) <= b;
    outputs(992) <= b and not a;
    outputs(993) <= a and not b;
    outputs(994) <= not a;
    outputs(995) <= not b;
    outputs(996) <= b and not a;
    outputs(997) <= a and b;
    outputs(998) <= a;
    outputs(999) <= a;
    outputs(1000) <= a and b;
    outputs(1001) <= b and not a;
    outputs(1002) <= not a;
    outputs(1003) <= not b or a;
    outputs(1004) <= a xor b;
    outputs(1005) <= not a;
    outputs(1006) <= a or b;
    outputs(1007) <= b;
    outputs(1008) <= a and not b;
    outputs(1009) <= b and not a;
    outputs(1010) <= a and not b;
    outputs(1011) <= not a;
    outputs(1012) <= b;
    outputs(1013) <= not a;
    outputs(1014) <= a and b;
    outputs(1015) <= not (a or b);
    outputs(1016) <= not (a or b);
    outputs(1017) <= a and not b;
    outputs(1018) <= a and b;
    outputs(1019) <= a and not b;
    outputs(1020) <= not b;
    outputs(1021) <= a or b;
    outputs(1022) <= not b or a;
    outputs(1023) <= a xor b;
    outputs(1024) <= b and not a;
    outputs(1025) <= a and not b;
    outputs(1026) <= not b;
    outputs(1027) <= a and b;
    outputs(1028) <= not b;
    outputs(1029) <= a xor b;
    outputs(1030) <= b;
    outputs(1031) <= b and not a;
    outputs(1032) <= a xor b;
    outputs(1033) <= not b;
    outputs(1034) <= b and not a;
    outputs(1035) <= not a;
    outputs(1036) <= not b;
    outputs(1037) <= b and not a;
    outputs(1038) <= not b;
    outputs(1039) <= b;
    outputs(1040) <= not b;
    outputs(1041) <= not b;
    outputs(1042) <= a and not b;
    outputs(1043) <= not (a xor b);
    outputs(1044) <= a and not b;
    outputs(1045) <= b;
    outputs(1046) <= b;
    outputs(1047) <= b and not a;
    outputs(1048) <= not b;
    outputs(1049) <= not (a or b);
    outputs(1050) <= not (a xor b);
    outputs(1051) <= not (a xor b);
    outputs(1052) <= a and not b;
    outputs(1053) <= b and not a;
    outputs(1054) <= not (a and b);
    outputs(1055) <= a and not b;
    outputs(1056) <= not b or a;
    outputs(1057) <= a and b;
    outputs(1058) <= a xor b;
    outputs(1059) <= a and b;
    outputs(1060) <= a and b;
    outputs(1061) <= b;
    outputs(1062) <= b and not a;
    outputs(1063) <= b and not a;
    outputs(1064) <= not (a xor b);
    outputs(1065) <= a or b;
    outputs(1066) <= a;
    outputs(1067) <= a;
    outputs(1068) <= not b;
    outputs(1069) <= a;
    outputs(1070) <= not (a xor b);
    outputs(1071) <= b;
    outputs(1072) <= b and not a;
    outputs(1073) <= a and not b;
    outputs(1074) <= b;
    outputs(1075) <= not (a xor b);
    outputs(1076) <= a and not b;
    outputs(1077) <= a and not b;
    outputs(1078) <= a;
    outputs(1079) <= not (a xor b);
    outputs(1080) <= a xor b;
    outputs(1081) <= a and b;
    outputs(1082) <= a and b;
    outputs(1083) <= not a;
    outputs(1084) <= a and b;
    outputs(1085) <= not a;
    outputs(1086) <= b;
    outputs(1087) <= not (a xor b);
    outputs(1088) <= not b;
    outputs(1089) <= a and not b;
    outputs(1090) <= not b;
    outputs(1091) <= a and b;
    outputs(1092) <= b and not a;
    outputs(1093) <= a and not b;
    outputs(1094) <= not a or b;
    outputs(1095) <= a and not b;
    outputs(1096) <= not b;
    outputs(1097) <= b;
    outputs(1098) <= a xor b;
    outputs(1099) <= b;
    outputs(1100) <= a and not b;
    outputs(1101) <= not b;
    outputs(1102) <= b and not a;
    outputs(1103) <= b and not a;
    outputs(1104) <= a and b;
    outputs(1105) <= not b;
    outputs(1106) <= not b;
    outputs(1107) <= not (a xor b);
    outputs(1108) <= b;
    outputs(1109) <= not (a or b);
    outputs(1110) <= a and not b;
    outputs(1111) <= a and not b;
    outputs(1112) <= b and not a;
    outputs(1113) <= a;
    outputs(1114) <= not (a or b);
    outputs(1115) <= not (a and b);
    outputs(1116) <= a and not b;
    outputs(1117) <= a and b;
    outputs(1118) <= a xor b;
    outputs(1119) <= not a;
    outputs(1120) <= not (a xor b);
    outputs(1121) <= a and not b;
    outputs(1122) <= a;
    outputs(1123) <= a and not b;
    outputs(1124) <= not (a or b);
    outputs(1125) <= b and not a;
    outputs(1126) <= a xor b;
    outputs(1127) <= not (a or b);
    outputs(1128) <= a and b;
    outputs(1129) <= a and not b;
    outputs(1130) <= a and not b;
    outputs(1131) <= not a;
    outputs(1132) <= not a;
    outputs(1133) <= not b;
    outputs(1134) <= not a or b;
    outputs(1135) <= not b or a;
    outputs(1136) <= a and b;
    outputs(1137) <= not (a or b);
    outputs(1138) <= b and not a;
    outputs(1139) <= not (a xor b);
    outputs(1140) <= a and b;
    outputs(1141) <= a and not b;
    outputs(1142) <= not b;
    outputs(1143) <= a xor b;
    outputs(1144) <= not b or a;
    outputs(1145) <= not a;
    outputs(1146) <= a xor b;
    outputs(1147) <= a;
    outputs(1148) <= a xor b;
    outputs(1149) <= not a;
    outputs(1150) <= not a;
    outputs(1151) <= not a;
    outputs(1152) <= not (a or b);
    outputs(1153) <= b and not a;
    outputs(1154) <= not (a xor b);
    outputs(1155) <= b;
    outputs(1156) <= not (a xor b);
    outputs(1157) <= b and not a;
    outputs(1158) <= not b;
    outputs(1159) <= a and b;
    outputs(1160) <= b and not a;
    outputs(1161) <= a xor b;
    outputs(1162) <= a and not b;
    outputs(1163) <= b;
    outputs(1164) <= not (a xor b);
    outputs(1165) <= b and not a;
    outputs(1166) <= a and not b;
    outputs(1167) <= not (a or b);
    outputs(1168) <= b;
    outputs(1169) <= a and b;
    outputs(1170) <= not b;
    outputs(1171) <= a and b;
    outputs(1172) <= b;
    outputs(1173) <= b;
    outputs(1174) <= b;
    outputs(1175) <= not b;
    outputs(1176) <= not (a xor b);
    outputs(1177) <= b and not a;
    outputs(1178) <= not (a or b);
    outputs(1179) <= b and not a;
    outputs(1180) <= b and not a;
    outputs(1181) <= not (a and b);
    outputs(1182) <= not a;
    outputs(1183) <= b and not a;
    outputs(1184) <= b;
    outputs(1185) <= not (a or b);
    outputs(1186) <= a and b;
    outputs(1187) <= a;
    outputs(1188) <= a xor b;
    outputs(1189) <= a and not b;
    outputs(1190) <= not a;
    outputs(1191) <= a xor b;
    outputs(1192) <= not a;
    outputs(1193) <= not a;
    outputs(1194) <= a;
    outputs(1195) <= not a;
    outputs(1196) <= not a;
    outputs(1197) <= a and b;
    outputs(1198) <= a and b;
    outputs(1199) <= a and b;
    outputs(1200) <= b and not a;
    outputs(1201) <= b and not a;
    outputs(1202) <= not (a or b);
    outputs(1203) <= not b;
    outputs(1204) <= not a;
    outputs(1205) <= a and not b;
    outputs(1206) <= not b;
    outputs(1207) <= a and b;
    outputs(1208) <= a and not b;
    outputs(1209) <= not b;
    outputs(1210) <= a xor b;
    outputs(1211) <= not (a xor b);
    outputs(1212) <= not b or a;
    outputs(1213) <= b and not a;
    outputs(1214) <= not (a xor b);
    outputs(1215) <= a;
    outputs(1216) <= a and b;
    outputs(1217) <= a and not b;
    outputs(1218) <= not (a or b);
    outputs(1219) <= not a or b;
    outputs(1220) <= b and not a;
    outputs(1221) <= not (a xor b);
    outputs(1222) <= b and not a;
    outputs(1223) <= b and not a;
    outputs(1224) <= b;
    outputs(1225) <= b and not a;
    outputs(1226) <= not b;
    outputs(1227) <= a and not b;
    outputs(1228) <= not (a or b);
    outputs(1229) <= b;
    outputs(1230) <= not a;
    outputs(1231) <= not a;
    outputs(1232) <= a xor b;
    outputs(1233) <= b and not a;
    outputs(1234) <= a and not b;
    outputs(1235) <= a and b;
    outputs(1236) <= a and b;
    outputs(1237) <= b and not a;
    outputs(1238) <= not a;
    outputs(1239) <= not a;
    outputs(1240) <= not b;
    outputs(1241) <= not (a xor b);
    outputs(1242) <= not (a xor b);
    outputs(1243) <= b and not a;
    outputs(1244) <= b;
    outputs(1245) <= not b;
    outputs(1246) <= b;
    outputs(1247) <= a and b;
    outputs(1248) <= b;
    outputs(1249) <= a and not b;
    outputs(1250) <= a xor b;
    outputs(1251) <= not (a and b);
    outputs(1252) <= b and not a;
    outputs(1253) <= not a;
    outputs(1254) <= b;
    outputs(1255) <= b and not a;
    outputs(1256) <= not b;
    outputs(1257) <= a and not b;
    outputs(1258) <= a or b;
    outputs(1259) <= not a;
    outputs(1260) <= a and not b;
    outputs(1261) <= not a;
    outputs(1262) <= not b;
    outputs(1263) <= a;
    outputs(1264) <= not (a xor b);
    outputs(1265) <= b;
    outputs(1266) <= a and b;
    outputs(1267) <= not b;
    outputs(1268) <= a;
    outputs(1269) <= not b;
    outputs(1270) <= b and not a;
    outputs(1271) <= a and b;
    outputs(1272) <= not b;
    outputs(1273) <= b;
    outputs(1274) <= a and b;
    outputs(1275) <= a xor b;
    outputs(1276) <= not (a xor b);
    outputs(1277) <= a;
    outputs(1278) <= b;
    outputs(1279) <= not a;
    outputs(1280) <= not b;
    outputs(1281) <= b and not a;
    outputs(1282) <= a and not b;
    outputs(1283) <= not (a xor b);
    outputs(1284) <= not b;
    outputs(1285) <= not b;
    outputs(1286) <= a xor b;
    outputs(1287) <= b;
    outputs(1288) <= b;
    outputs(1289) <= a or b;
    outputs(1290) <= a and b;
    outputs(1291) <= not (a xor b);
    outputs(1292) <= not (a or b);
    outputs(1293) <= a;
    outputs(1294) <= a and not b;
    outputs(1295) <= a and b;
    outputs(1296) <= b and not a;
    outputs(1297) <= not b or a;
    outputs(1298) <= a and b;
    outputs(1299) <= not a or b;
    outputs(1300) <= not (a or b);
    outputs(1301) <= b;
    outputs(1302) <= not (a or b);
    outputs(1303) <= a and not b;
    outputs(1304) <= b and not a;
    outputs(1305) <= a and b;
    outputs(1306) <= not a;
    outputs(1307) <= not (a or b);
    outputs(1308) <= not a;
    outputs(1309) <= a;
    outputs(1310) <= a and b;
    outputs(1311) <= b and not a;
    outputs(1312) <= b and not a;
    outputs(1313) <= not (a xor b);
    outputs(1314) <= a;
    outputs(1315) <= a xor b;
    outputs(1316) <= b;
    outputs(1317) <= a and b;
    outputs(1318) <= not a;
    outputs(1319) <= a;
    outputs(1320) <= not a;
    outputs(1321) <= b;
    outputs(1322) <= a xor b;
    outputs(1323) <= a;
    outputs(1324) <= not (a or b);
    outputs(1325) <= not a;
    outputs(1326) <= a xor b;
    outputs(1327) <= b;
    outputs(1328) <= not (a or b);
    outputs(1329) <= a and b;
    outputs(1330) <= not b or a;
    outputs(1331) <= not b or a;
    outputs(1332) <= not b;
    outputs(1333) <= not (a or b);
    outputs(1334) <= not (a or b);
    outputs(1335) <= not a;
    outputs(1336) <= a xor b;
    outputs(1337) <= a;
    outputs(1338) <= b;
    outputs(1339) <= a and not b;
    outputs(1340) <= a;
    outputs(1341) <= not (a xor b);
    outputs(1342) <= a and b;
    outputs(1343) <= a and not b;
    outputs(1344) <= not b;
    outputs(1345) <= not b;
    outputs(1346) <= not a or b;
    outputs(1347) <= a xor b;
    outputs(1348) <= b;
    outputs(1349) <= a and b;
    outputs(1350) <= not b;
    outputs(1351) <= a xor b;
    outputs(1352) <= not b;
    outputs(1353) <= b and not a;
    outputs(1354) <= a and b;
    outputs(1355) <= a and not b;
    outputs(1356) <= not a;
    outputs(1357) <= a and b;
    outputs(1358) <= not a or b;
    outputs(1359) <= a and not b;
    outputs(1360) <= not b or a;
    outputs(1361) <= a xor b;
    outputs(1362) <= b;
    outputs(1363) <= a;
    outputs(1364) <= not a;
    outputs(1365) <= not a;
    outputs(1366) <= a xor b;
    outputs(1367) <= a;
    outputs(1368) <= not a or b;
    outputs(1369) <= not (a xor b);
    outputs(1370) <= b and not a;
    outputs(1371) <= not a;
    outputs(1372) <= b and not a;
    outputs(1373) <= b;
    outputs(1374) <= not a;
    outputs(1375) <= not a;
    outputs(1376) <= a and not b;
    outputs(1377) <= not a or b;
    outputs(1378) <= a xor b;
    outputs(1379) <= a;
    outputs(1380) <= a;
    outputs(1381) <= b;
    outputs(1382) <= not a;
    outputs(1383) <= a;
    outputs(1384) <= not a or b;
    outputs(1385) <= not a;
    outputs(1386) <= not (a or b);
    outputs(1387) <= b and not a;
    outputs(1388) <= b and not a;
    outputs(1389) <= b;
    outputs(1390) <= a and b;
    outputs(1391) <= b and not a;
    outputs(1392) <= a and b;
    outputs(1393) <= not (a xor b);
    outputs(1394) <= a;
    outputs(1395) <= a and not b;
    outputs(1396) <= not b;
    outputs(1397) <= a and not b;
    outputs(1398) <= a or b;
    outputs(1399) <= not a or b;
    outputs(1400) <= not b or a;
    outputs(1401) <= not (a xor b);
    outputs(1402) <= not b;
    outputs(1403) <= a and b;
    outputs(1404) <= b and not a;
    outputs(1405) <= not (a or b);
    outputs(1406) <= not (a xor b);
    outputs(1407) <= a and b;
    outputs(1408) <= b;
    outputs(1409) <= not (a or b);
    outputs(1410) <= a and not b;
    outputs(1411) <= a and not b;
    outputs(1412) <= not (a or b);
    outputs(1413) <= not (a xor b);
    outputs(1414) <= a and not b;
    outputs(1415) <= a and not b;
    outputs(1416) <= not b;
    outputs(1417) <= 1'b0;
    outputs(1418) <= b and not a;
    outputs(1419) <= not b;
    outputs(1420) <= a;
    outputs(1421) <= b and not a;
    outputs(1422) <= a and b;
    outputs(1423) <= not (a xor b);
    outputs(1424) <= a;
    outputs(1425) <= a;
    outputs(1426) <= b;
    outputs(1427) <= not (a or b);
    outputs(1428) <= a xor b;
    outputs(1429) <= not b;
    outputs(1430) <= b and not a;
    outputs(1431) <= not (a or b);
    outputs(1432) <= a;
    outputs(1433) <= b and not a;
    outputs(1434) <= a xor b;
    outputs(1435) <= not (a and b);
    outputs(1436) <= not a;
    outputs(1437) <= not (a xor b);
    outputs(1438) <= not b or a;
    outputs(1439) <= not (a xor b);
    outputs(1440) <= not (a and b);
    outputs(1441) <= not a or b;
    outputs(1442) <= a xor b;
    outputs(1443) <= a xor b;
    outputs(1444) <= not (a and b);
    outputs(1445) <= a xor b;
    outputs(1446) <= b;
    outputs(1447) <= a;
    outputs(1448) <= a xor b;
    outputs(1449) <= b;
    outputs(1450) <= a xor b;
    outputs(1451) <= not b or a;
    outputs(1452) <= not b;
    outputs(1453) <= a xor b;
    outputs(1454) <= a or b;
    outputs(1455) <= a;
    outputs(1456) <= b and not a;
    outputs(1457) <= a or b;
    outputs(1458) <= not (a xor b);
    outputs(1459) <= not (a or b);
    outputs(1460) <= not (a and b);
    outputs(1461) <= a and b;
    outputs(1462) <= not b or a;
    outputs(1463) <= b;
    outputs(1464) <= a and b;
    outputs(1465) <= b;
    outputs(1466) <= b and not a;
    outputs(1467) <= a xor b;
    outputs(1468) <= a or b;
    outputs(1469) <= not (a and b);
    outputs(1470) <= not b;
    outputs(1471) <= b and not a;
    outputs(1472) <= a;
    outputs(1473) <= not (a xor b);
    outputs(1474) <= a and not b;
    outputs(1475) <= b and not a;
    outputs(1476) <= a xor b;
    outputs(1477) <= not (a or b);
    outputs(1478) <= a;
    outputs(1479) <= a and not b;
    outputs(1480) <= not b or a;
    outputs(1481) <= a;
    outputs(1482) <= not (a xor b);
    outputs(1483) <= not (a or b);
    outputs(1484) <= a and b;
    outputs(1485) <= a xor b;
    outputs(1486) <= not b;
    outputs(1487) <= b and not a;
    outputs(1488) <= not (a or b);
    outputs(1489) <= b;
    outputs(1490) <= a and not b;
    outputs(1491) <= a xor b;
    outputs(1492) <= a and b;
    outputs(1493) <= not (a xor b);
    outputs(1494) <= not (a and b);
    outputs(1495) <= not (a xor b);
    outputs(1496) <= not b or a;
    outputs(1497) <= not (a xor b);
    outputs(1498) <= a and b;
    outputs(1499) <= a xor b;
    outputs(1500) <= b;
    outputs(1501) <= a;
    outputs(1502) <= b and not a;
    outputs(1503) <= a and not b;
    outputs(1504) <= not (a or b);
    outputs(1505) <= not a or b;
    outputs(1506) <= not b or a;
    outputs(1507) <= not a;
    outputs(1508) <= a and b;
    outputs(1509) <= a and not b;
    outputs(1510) <= a and not b;
    outputs(1511) <= not (a xor b);
    outputs(1512) <= not (a or b);
    outputs(1513) <= a;
    outputs(1514) <= not (a or b);
    outputs(1515) <= a and not b;
    outputs(1516) <= b;
    outputs(1517) <= a and b;
    outputs(1518) <= not a;
    outputs(1519) <= a and not b;
    outputs(1520) <= b and not a;
    outputs(1521) <= a and b;
    outputs(1522) <= not b or a;
    outputs(1523) <= not b;
    outputs(1524) <= a and b;
    outputs(1525) <= a;
    outputs(1526) <= a or b;
    outputs(1527) <= b;
    outputs(1528) <= b;
    outputs(1529) <= not b;
    outputs(1530) <= b and not a;
    outputs(1531) <= a xor b;
    outputs(1532) <= not (a or b);
    outputs(1533) <= not a;
    outputs(1534) <= not (a xor b);
    outputs(1535) <= a and b;
    outputs(1536) <= a and b;
    outputs(1537) <= a;
    outputs(1538) <= not a;
    outputs(1539) <= not a;
    outputs(1540) <= not b;
    outputs(1541) <= a or b;
    outputs(1542) <= a;
    outputs(1543) <= not b;
    outputs(1544) <= not (a and b);
    outputs(1545) <= a xor b;
    outputs(1546) <= b and not a;
    outputs(1547) <= b;
    outputs(1548) <= not b;
    outputs(1549) <= a and not b;
    outputs(1550) <= not a;
    outputs(1551) <= not a;
    outputs(1552) <= b;
    outputs(1553) <= a or b;
    outputs(1554) <= a and b;
    outputs(1555) <= b;
    outputs(1556) <= a xor b;
    outputs(1557) <= b;
    outputs(1558) <= a and b;
    outputs(1559) <= not b;
    outputs(1560) <= b;
    outputs(1561) <= a;
    outputs(1562) <= a;
    outputs(1563) <= not (a xor b);
    outputs(1564) <= b and not a;
    outputs(1565) <= not b;
    outputs(1566) <= a;
    outputs(1567) <= a and not b;
    outputs(1568) <= b and not a;
    outputs(1569) <= a and b;
    outputs(1570) <= a or b;
    outputs(1571) <= not a or b;
    outputs(1572) <= a and not b;
    outputs(1573) <= not (a xor b);
    outputs(1574) <= not a;
    outputs(1575) <= b and not a;
    outputs(1576) <= b and not a;
    outputs(1577) <= not a;
    outputs(1578) <= not a;
    outputs(1579) <= a xor b;
    outputs(1580) <= a or b;
    outputs(1581) <= b;
    outputs(1582) <= a and b;
    outputs(1583) <= not b;
    outputs(1584) <= not b;
    outputs(1585) <= not (a or b);
    outputs(1586) <= a and not b;
    outputs(1587) <= a;
    outputs(1588) <= a and b;
    outputs(1589) <= a;
    outputs(1590) <= b and not a;
    outputs(1591) <= not (a or b);
    outputs(1592) <= not a;
    outputs(1593) <= b;
    outputs(1594) <= b and not a;
    outputs(1595) <= b;
    outputs(1596) <= not b;
    outputs(1597) <= b and not a;
    outputs(1598) <= not a;
    outputs(1599) <= not (a or b);
    outputs(1600) <= a xor b;
    outputs(1601) <= not a or b;
    outputs(1602) <= not (a or b);
    outputs(1603) <= not (a or b);
    outputs(1604) <= not a;
    outputs(1605) <= not b;
    outputs(1606) <= not b;
    outputs(1607) <= a;
    outputs(1608) <= a and b;
    outputs(1609) <= a xor b;
    outputs(1610) <= b and not a;
    outputs(1611) <= not (a or b);
    outputs(1612) <= b and not a;
    outputs(1613) <= not (a or b);
    outputs(1614) <= b and not a;
    outputs(1615) <= not a;
    outputs(1616) <= not b;
    outputs(1617) <= b;
    outputs(1618) <= not (a or b);
    outputs(1619) <= b and not a;
    outputs(1620) <= not (a xor b);
    outputs(1621) <= a and b;
    outputs(1622) <= not b;
    outputs(1623) <= a and not b;
    outputs(1624) <= a xor b;
    outputs(1625) <= b;
    outputs(1626) <= a;
    outputs(1627) <= a and not b;
    outputs(1628) <= not (a xor b);
    outputs(1629) <= not (a xor b);
    outputs(1630) <= a and b;
    outputs(1631) <= a and b;
    outputs(1632) <= not a or b;
    outputs(1633) <= not (a or b);
    outputs(1634) <= a and not b;
    outputs(1635) <= a xor b;
    outputs(1636) <= b and not a;
    outputs(1637) <= b and not a;
    outputs(1638) <= b;
    outputs(1639) <= a and not b;
    outputs(1640) <= b;
    outputs(1641) <= not (a or b);
    outputs(1642) <= a;
    outputs(1643) <= not (a xor b);
    outputs(1644) <= a;
    outputs(1645) <= not (a xor b);
    outputs(1646) <= a;
    outputs(1647) <= not a;
    outputs(1648) <= b;
    outputs(1649) <= a and not b;
    outputs(1650) <= not a;
    outputs(1651) <= b;
    outputs(1652) <= a and b;
    outputs(1653) <= not (a xor b);
    outputs(1654) <= a and b;
    outputs(1655) <= a and b;
    outputs(1656) <= not b;
    outputs(1657) <= a xor b;
    outputs(1658) <= not a;
    outputs(1659) <= b;
    outputs(1660) <= not (a xor b);
    outputs(1661) <= not b;
    outputs(1662) <= b;
    outputs(1663) <= not b or a;
    outputs(1664) <= a xor b;
    outputs(1665) <= a and not b;
    outputs(1666) <= b and not a;
    outputs(1667) <= a and b;
    outputs(1668) <= b and not a;
    outputs(1669) <= not a or b;
    outputs(1670) <= not (a and b);
    outputs(1671) <= a and b;
    outputs(1672) <= not (a xor b);
    outputs(1673) <= not a;
    outputs(1674) <= not b;
    outputs(1675) <= b;
    outputs(1676) <= a and not b;
    outputs(1677) <= a xor b;
    outputs(1678) <= not b;
    outputs(1679) <= not (a or b);
    outputs(1680) <= not (a or b);
    outputs(1681) <= not (a xor b);
    outputs(1682) <= not (a or b);
    outputs(1683) <= not b;
    outputs(1684) <= a xor b;
    outputs(1685) <= not (a xor b);
    outputs(1686) <= a and not b;
    outputs(1687) <= a and b;
    outputs(1688) <= not a;
    outputs(1689) <= a and b;
    outputs(1690) <= a and not b;
    outputs(1691) <= not b;
    outputs(1692) <= not (a xor b);
    outputs(1693) <= not (a xor b);
    outputs(1694) <= not b or a;
    outputs(1695) <= b;
    outputs(1696) <= a and b;
    outputs(1697) <= not b;
    outputs(1698) <= not a or b;
    outputs(1699) <= b and not a;
    outputs(1700) <= not b;
    outputs(1701) <= not b or a;
    outputs(1702) <= a xor b;
    outputs(1703) <= b and not a;
    outputs(1704) <= not a or b;
    outputs(1705) <= b;
    outputs(1706) <= not b or a;
    outputs(1707) <= a and b;
    outputs(1708) <= a and b;
    outputs(1709) <= not b;
    outputs(1710) <= b;
    outputs(1711) <= a;
    outputs(1712) <= not b or a;
    outputs(1713) <= not a or b;
    outputs(1714) <= not (a xor b);
    outputs(1715) <= not (a or b);
    outputs(1716) <= not (a or b);
    outputs(1717) <= not (a or b);
    outputs(1718) <= b;
    outputs(1719) <= b;
    outputs(1720) <= not (a or b);
    outputs(1721) <= not a;
    outputs(1722) <= a;
    outputs(1723) <= a and b;
    outputs(1724) <= a and not b;
    outputs(1725) <= not (a or b);
    outputs(1726) <= not b;
    outputs(1727) <= not b;
    outputs(1728) <= b;
    outputs(1729) <= a and not b;
    outputs(1730) <= not (a or b);
    outputs(1731) <= not a;
    outputs(1732) <= not (a or b);
    outputs(1733) <= a or b;
    outputs(1734) <= a;
    outputs(1735) <= not (a and b);
    outputs(1736) <= a and b;
    outputs(1737) <= a and not b;
    outputs(1738) <= b;
    outputs(1739) <= b and not a;
    outputs(1740) <= not (a or b);
    outputs(1741) <= not (a xor b);
    outputs(1742) <= a and b;
    outputs(1743) <= a xor b;
    outputs(1744) <= not b;
    outputs(1745) <= not (a or b);
    outputs(1746) <= a and not b;
    outputs(1747) <= a and not b;
    outputs(1748) <= not a;
    outputs(1749) <= b and not a;
    outputs(1750) <= b;
    outputs(1751) <= not (a or b);
    outputs(1752) <= not a;
    outputs(1753) <= not b;
    outputs(1754) <= a xor b;
    outputs(1755) <= not a;
    outputs(1756) <= not (a xor b);
    outputs(1757) <= b and not a;
    outputs(1758) <= a;
    outputs(1759) <= not b or a;
    outputs(1760) <= b and not a;
    outputs(1761) <= not b;
    outputs(1762) <= a or b;
    outputs(1763) <= not (a and b);
    outputs(1764) <= not a;
    outputs(1765) <= not a;
    outputs(1766) <= b and not a;
    outputs(1767) <= not (a or b);
    outputs(1768) <= a xor b;
    outputs(1769) <= not a;
    outputs(1770) <= b;
    outputs(1771) <= not (a xor b);
    outputs(1772) <= a and not b;
    outputs(1773) <= b and not a;
    outputs(1774) <= a or b;
    outputs(1775) <= a and not b;
    outputs(1776) <= a;
    outputs(1777) <= b;
    outputs(1778) <= a and b;
    outputs(1779) <= b and not a;
    outputs(1780) <= b and not a;
    outputs(1781) <= not (a or b);
    outputs(1782) <= not b or a;
    outputs(1783) <= not (a or b);
    outputs(1784) <= a and b;
    outputs(1785) <= not (a or b);
    outputs(1786) <= a xor b;
    outputs(1787) <= b;
    outputs(1788) <= a xor b;
    outputs(1789) <= a;
    outputs(1790) <= not b;
    outputs(1791) <= a;
    outputs(1792) <= not (a xor b);
    outputs(1793) <= a xor b;
    outputs(1794) <= b;
    outputs(1795) <= a and b;
    outputs(1796) <= not b;
    outputs(1797) <= a and b;
    outputs(1798) <= not b;
    outputs(1799) <= not b or a;
    outputs(1800) <= not a or b;
    outputs(1801) <= not b;
    outputs(1802) <= a;
    outputs(1803) <= a and b;
    outputs(1804) <= a and b;
    outputs(1805) <= a and b;
    outputs(1806) <= a or b;
    outputs(1807) <= not b or a;
    outputs(1808) <= not a;
    outputs(1809) <= b and not a;
    outputs(1810) <= b and not a;
    outputs(1811) <= b;
    outputs(1812) <= not (a or b);
    outputs(1813) <= a and b;
    outputs(1814) <= not (a xor b);
    outputs(1815) <= a and b;
    outputs(1816) <= not (a or b);
    outputs(1817) <= a and b;
    outputs(1818) <= b and not a;
    outputs(1819) <= b;
    outputs(1820) <= a and b;
    outputs(1821) <= a and b;
    outputs(1822) <= not a;
    outputs(1823) <= b;
    outputs(1824) <= not b;
    outputs(1825) <= not a or b;
    outputs(1826) <= a and not b;
    outputs(1827) <= a and not b;
    outputs(1828) <= a and b;
    outputs(1829) <= a and b;
    outputs(1830) <= not a;
    outputs(1831) <= a or b;
    outputs(1832) <= a and not b;
    outputs(1833) <= a and b;
    outputs(1834) <= a;
    outputs(1835) <= a and b;
    outputs(1836) <= not a;
    outputs(1837) <= b and not a;
    outputs(1838) <= a xor b;
    outputs(1839) <= b and not a;
    outputs(1840) <= b and not a;
    outputs(1841) <= a and b;
    outputs(1842) <= b and not a;
    outputs(1843) <= a and b;
    outputs(1844) <= not (a xor b);
    outputs(1845) <= not b;
    outputs(1846) <= not (a xor b);
    outputs(1847) <= a and not b;
    outputs(1848) <= a;
    outputs(1849) <= not b or a;
    outputs(1850) <= not b;
    outputs(1851) <= a xor b;
    outputs(1852) <= a xor b;
    outputs(1853) <= not (a and b);
    outputs(1854) <= b;
    outputs(1855) <= b;
    outputs(1856) <= a and b;
    outputs(1857) <= b and not a;
    outputs(1858) <= a and not b;
    outputs(1859) <= a and b;
    outputs(1860) <= a and not b;
    outputs(1861) <= a xor b;
    outputs(1862) <= a and not b;
    outputs(1863) <= not (a or b);
    outputs(1864) <= a;
    outputs(1865) <= a and b;
    outputs(1866) <= a and b;
    outputs(1867) <= a and not b;
    outputs(1868) <= a;
    outputs(1869) <= a and b;
    outputs(1870) <= a;
    outputs(1871) <= a;
    outputs(1872) <= a and not b;
    outputs(1873) <= not b or a;
    outputs(1874) <= a and b;
    outputs(1875) <= a;
    outputs(1876) <= not b;
    outputs(1877) <= a and not b;
    outputs(1878) <= b;
    outputs(1879) <= not b;
    outputs(1880) <= not b;
    outputs(1881) <= not a or b;
    outputs(1882) <= not (a or b);
    outputs(1883) <= b and not a;
    outputs(1884) <= not (a or b);
    outputs(1885) <= not b or a;
    outputs(1886) <= b and not a;
    outputs(1887) <= not (a or b);
    outputs(1888) <= a or b;
    outputs(1889) <= not (a or b);
    outputs(1890) <= a and not b;
    outputs(1891) <= a;
    outputs(1892) <= a and not b;
    outputs(1893) <= b;
    outputs(1894) <= a and b;
    outputs(1895) <= not a;
    outputs(1896) <= not (a and b);
    outputs(1897) <= a and b;
    outputs(1898) <= not (a and b);
    outputs(1899) <= not (a or b);
    outputs(1900) <= b and not a;
    outputs(1901) <= not (a xor b);
    outputs(1902) <= not a;
    outputs(1903) <= not (a or b);
    outputs(1904) <= b and not a;
    outputs(1905) <= b and not a;
    outputs(1906) <= b and not a;
    outputs(1907) <= a and b;
    outputs(1908) <= a;
    outputs(1909) <= not b;
    outputs(1910) <= a xor b;
    outputs(1911) <= b;
    outputs(1912) <= a and not b;
    outputs(1913) <= not (a and b);
    outputs(1914) <= not a;
    outputs(1915) <= not a;
    outputs(1916) <= b and not a;
    outputs(1917) <= not a;
    outputs(1918) <= b and not a;
    outputs(1919) <= b and not a;
    outputs(1920) <= a and not b;
    outputs(1921) <= not (a or b);
    outputs(1922) <= not b or a;
    outputs(1923) <= a;
    outputs(1924) <= a;
    outputs(1925) <= b and not a;
    outputs(1926) <= not a or b;
    outputs(1927) <= b;
    outputs(1928) <= b and not a;
    outputs(1929) <= not b;
    outputs(1930) <= b and not a;
    outputs(1931) <= a and not b;
    outputs(1932) <= a xor b;
    outputs(1933) <= not (a or b);
    outputs(1934) <= a and not b;
    outputs(1935) <= not b;
    outputs(1936) <= not a;
    outputs(1937) <= a and b;
    outputs(1938) <= not (a and b);
    outputs(1939) <= a;
    outputs(1940) <= not (a or b);
    outputs(1941) <= a or b;
    outputs(1942) <= not a;
    outputs(1943) <= a and b;
    outputs(1944) <= not (a or b);
    outputs(1945) <= a xor b;
    outputs(1946) <= b and not a;
    outputs(1947) <= a and b;
    outputs(1948) <= not (a or b);
    outputs(1949) <= a and b;
    outputs(1950) <= b;
    outputs(1951) <= not b;
    outputs(1952) <= not b;
    outputs(1953) <= b and not a;
    outputs(1954) <= a and b;
    outputs(1955) <= b;
    outputs(1956) <= a xor b;
    outputs(1957) <= not b;
    outputs(1958) <= b and not a;
    outputs(1959) <= not (a xor b);
    outputs(1960) <= not (a or b);
    outputs(1961) <= a;
    outputs(1962) <= a xor b;
    outputs(1963) <= b;
    outputs(1964) <= a;
    outputs(1965) <= a and not b;
    outputs(1966) <= a and b;
    outputs(1967) <= not a;
    outputs(1968) <= a and not b;
    outputs(1969) <= not b;
    outputs(1970) <= not (a or b);
    outputs(1971) <= b and not a;
    outputs(1972) <= not a;
    outputs(1973) <= a and b;
    outputs(1974) <= not b;
    outputs(1975) <= a xor b;
    outputs(1976) <= a and b;
    outputs(1977) <= not b;
    outputs(1978) <= not a;
    outputs(1979) <= not (a or b);
    outputs(1980) <= not b or a;
    outputs(1981) <= b;
    outputs(1982) <= a or b;
    outputs(1983) <= not b;
    outputs(1984) <= not (a or b);
    outputs(1985) <= not (a xor b);
    outputs(1986) <= b;
    outputs(1987) <= not (a or b);
    outputs(1988) <= a;
    outputs(1989) <= a and not b;
    outputs(1990) <= b;
    outputs(1991) <= not b;
    outputs(1992) <= a and not b;
    outputs(1993) <= a and not b;
    outputs(1994) <= a or b;
    outputs(1995) <= b;
    outputs(1996) <= a and b;
    outputs(1997) <= a xor b;
    outputs(1998) <= b and not a;
    outputs(1999) <= a and b;
    outputs(2000) <= a and not b;
    outputs(2001) <= not b;
    outputs(2002) <= not a;
    outputs(2003) <= b;
    outputs(2004) <= not (a or b);
    outputs(2005) <= a and b;
    outputs(2006) <= not (a or b);
    outputs(2007) <= a and not b;
    outputs(2008) <= not a;
    outputs(2009) <= not (a or b);
    outputs(2010) <= not b;
    outputs(2011) <= not a or b;
    outputs(2012) <= a;
    outputs(2013) <= not b;
    outputs(2014) <= b and not a;
    outputs(2015) <= b;
    outputs(2016) <= not a;
    outputs(2017) <= b and not a;
    outputs(2018) <= a and b;
    outputs(2019) <= not (a or b);
    outputs(2020) <= b and not a;
    outputs(2021) <= a xor b;
    outputs(2022) <= not (a xor b);
    outputs(2023) <= b;
    outputs(2024) <= not a;
    outputs(2025) <= not (a xor b);
    outputs(2026) <= a and not b;
    outputs(2027) <= b;
    outputs(2028) <= a and not b;
    outputs(2029) <= not a;
    outputs(2030) <= a and b;
    outputs(2031) <= b and not a;
    outputs(2032) <= not (a or b);
    outputs(2033) <= not (a xor b);
    outputs(2034) <= b;
    outputs(2035) <= b;
    outputs(2036) <= a and not b;
    outputs(2037) <= not (a xor b);
    outputs(2038) <= a xor b;
    outputs(2039) <= a or b;
    outputs(2040) <= not a;
    outputs(2041) <= not a or b;
    outputs(2042) <= a and not b;
    outputs(2043) <= a and not b;
    outputs(2044) <= a and not b;
    outputs(2045) <= b and not a;
    outputs(2046) <= not (a xor b);
    outputs(2047) <= a;
    outputs(2048) <= a and b;
    outputs(2049) <= a xor b;
    outputs(2050) <= a xor b;
    outputs(2051) <= not (a xor b);
    outputs(2052) <= not (a xor b);
    outputs(2053) <= not a;
    outputs(2054) <= b;
    outputs(2055) <= not (a xor b);
    outputs(2056) <= not a;
    outputs(2057) <= a and b;
    outputs(2058) <= b;
    outputs(2059) <= not (a or b);
    outputs(2060) <= b and not a;
    outputs(2061) <= not (a or b);
    outputs(2062) <= not b or a;
    outputs(2063) <= a and not b;
    outputs(2064) <= not b or a;
    outputs(2065) <= not b;
    outputs(2066) <= not a;
    outputs(2067) <= b and not a;
    outputs(2068) <= not (a or b);
    outputs(2069) <= b and not a;
    outputs(2070) <= b and not a;
    outputs(2071) <= not b;
    outputs(2072) <= not b;
    outputs(2073) <= b and not a;
    outputs(2074) <= a;
    outputs(2075) <= not b;
    outputs(2076) <= not (a and b);
    outputs(2077) <= not b or a;
    outputs(2078) <= b and not a;
    outputs(2079) <= a;
    outputs(2080) <= not b;
    outputs(2081) <= not (a or b);
    outputs(2082) <= not (a xor b);
    outputs(2083) <= not b;
    outputs(2084) <= not b or a;
    outputs(2085) <= not (a xor b);
    outputs(2086) <= a and not b;
    outputs(2087) <= not (a or b);
    outputs(2088) <= b and not a;
    outputs(2089) <= not b;
    outputs(2090) <= not a or b;
    outputs(2091) <= a xor b;
    outputs(2092) <= not (a xor b);
    outputs(2093) <= not b;
    outputs(2094) <= not b;
    outputs(2095) <= b;
    outputs(2096) <= a and b;
    outputs(2097) <= not (a or b);
    outputs(2098) <= a and not b;
    outputs(2099) <= a xor b;
    outputs(2100) <= a;
    outputs(2101) <= b;
    outputs(2102) <= not (a or b);
    outputs(2103) <= a and not b;
    outputs(2104) <= a and b;
    outputs(2105) <= a and b;
    outputs(2106) <= not a;
    outputs(2107) <= b;
    outputs(2108) <= a xor b;
    outputs(2109) <= not a or b;
    outputs(2110) <= b;
    outputs(2111) <= a and b;
    outputs(2112) <= b;
    outputs(2113) <= a xor b;
    outputs(2114) <= not (a xor b);
    outputs(2115) <= not b or a;
    outputs(2116) <= not (a xor b);
    outputs(2117) <= not (a xor b);
    outputs(2118) <= b;
    outputs(2119) <= b;
    outputs(2120) <= a;
    outputs(2121) <= b and not a;
    outputs(2122) <= not a;
    outputs(2123) <= b and not a;
    outputs(2124) <= not b;
    outputs(2125) <= a or b;
    outputs(2126) <= not (a xor b);
    outputs(2127) <= not (a or b);
    outputs(2128) <= a and b;
    outputs(2129) <= not (a xor b);
    outputs(2130) <= a and not b;
    outputs(2131) <= not b;
    outputs(2132) <= not (a and b);
    outputs(2133) <= a;
    outputs(2134) <= not b or a;
    outputs(2135) <= b and not a;
    outputs(2136) <= not a;
    outputs(2137) <= not b;
    outputs(2138) <= b;
    outputs(2139) <= not a;
    outputs(2140) <= a xor b;
    outputs(2141) <= not (a or b);
    outputs(2142) <= b;
    outputs(2143) <= a and not b;
    outputs(2144) <= a and not b;
    outputs(2145) <= a and b;
    outputs(2146) <= not a;
    outputs(2147) <= not (a or b);
    outputs(2148) <= a xor b;
    outputs(2149) <= not (a xor b);
    outputs(2150) <= b;
    outputs(2151) <= a or b;
    outputs(2152) <= b and not a;
    outputs(2153) <= a and not b;
    outputs(2154) <= not b;
    outputs(2155) <= not b;
    outputs(2156) <= not (a and b);
    outputs(2157) <= a xor b;
    outputs(2158) <= not a;
    outputs(2159) <= a and not b;
    outputs(2160) <= not (a or b);
    outputs(2161) <= a;
    outputs(2162) <= b and not a;
    outputs(2163) <= not b;
    outputs(2164) <= not (a xor b);
    outputs(2165) <= b;
    outputs(2166) <= not a or b;
    outputs(2167) <= a and b;
    outputs(2168) <= b;
    outputs(2169) <= not (a xor b);
    outputs(2170) <= not a or b;
    outputs(2171) <= not (a xor b);
    outputs(2172) <= not (a xor b);
    outputs(2173) <= not b;
    outputs(2174) <= a and not b;
    outputs(2175) <= b and not a;
    outputs(2176) <= a and b;
    outputs(2177) <= not a;
    outputs(2178) <= not (a or b);
    outputs(2179) <= a and not b;
    outputs(2180) <= not (a or b);
    outputs(2181) <= b and not a;
    outputs(2182) <= b and not a;
    outputs(2183) <= not a;
    outputs(2184) <= not b;
    outputs(2185) <= a;
    outputs(2186) <= b and not a;
    outputs(2187) <= not b;
    outputs(2188) <= not (a xor b);
    outputs(2189) <= not b;
    outputs(2190) <= not (a and b);
    outputs(2191) <= a or b;
    outputs(2192) <= not a;
    outputs(2193) <= a;
    outputs(2194) <= not (a and b);
    outputs(2195) <= not b;
    outputs(2196) <= a;
    outputs(2197) <= a and not b;
    outputs(2198) <= a or b;
    outputs(2199) <= b and not a;
    outputs(2200) <= not a;
    outputs(2201) <= b;
    outputs(2202) <= not a;
    outputs(2203) <= a;
    outputs(2204) <= b and not a;
    outputs(2205) <= b and not a;
    outputs(2206) <= a and not b;
    outputs(2207) <= not (a xor b);
    outputs(2208) <= a and b;
    outputs(2209) <= not (a or b);
    outputs(2210) <= not (a xor b);
    outputs(2211) <= b and not a;
    outputs(2212) <= a or b;
    outputs(2213) <= a and b;
    outputs(2214) <= a and b;
    outputs(2215) <= not (a or b);
    outputs(2216) <= not (a and b);
    outputs(2217) <= not (a xor b);
    outputs(2218) <= a;
    outputs(2219) <= not a;
    outputs(2220) <= not b or a;
    outputs(2221) <= not (a or b);
    outputs(2222) <= b and not a;
    outputs(2223) <= b;
    outputs(2224) <= a;
    outputs(2225) <= not a;
    outputs(2226) <= b and not a;
    outputs(2227) <= not a or b;
    outputs(2228) <= a xor b;
    outputs(2229) <= not a;
    outputs(2230) <= b and not a;
    outputs(2231) <= b;
    outputs(2232) <= not a;
    outputs(2233) <= b and not a;
    outputs(2234) <= a and not b;
    outputs(2235) <= not (a or b);
    outputs(2236) <= not (a or b);
    outputs(2237) <= a;
    outputs(2238) <= a xor b;
    outputs(2239) <= not b;
    outputs(2240) <= a;
    outputs(2241) <= not a;
    outputs(2242) <= a;
    outputs(2243) <= not a or b;
    outputs(2244) <= not a or b;
    outputs(2245) <= not a;
    outputs(2246) <= b;
    outputs(2247) <= b and not a;
    outputs(2248) <= not b;
    outputs(2249) <= not a;
    outputs(2250) <= not a;
    outputs(2251) <= b;
    outputs(2252) <= not (a xor b);
    outputs(2253) <= a and not b;
    outputs(2254) <= a;
    outputs(2255) <= not a;
    outputs(2256) <= a xor b;
    outputs(2257) <= not (a or b);
    outputs(2258) <= a and b;
    outputs(2259) <= b and not a;
    outputs(2260) <= a and b;
    outputs(2261) <= not a;
    outputs(2262) <= a;
    outputs(2263) <= a xor b;
    outputs(2264) <= a;
    outputs(2265) <= b;
    outputs(2266) <= b and not a;
    outputs(2267) <= a xor b;
    outputs(2268) <= b;
    outputs(2269) <= not b;
    outputs(2270) <= a or b;
    outputs(2271) <= a xor b;
    outputs(2272) <= b and not a;
    outputs(2273) <= b and not a;
    outputs(2274) <= b and not a;
    outputs(2275) <= b and not a;
    outputs(2276) <= not a;
    outputs(2277) <= b and not a;
    outputs(2278) <= not a;
    outputs(2279) <= b and not a;
    outputs(2280) <= a xor b;
    outputs(2281) <= a and not b;
    outputs(2282) <= not (a and b);
    outputs(2283) <= not (a or b);
    outputs(2284) <= not a or b;
    outputs(2285) <= not (a or b);
    outputs(2286) <= a and b;
    outputs(2287) <= not (a or b);
    outputs(2288) <= not b;
    outputs(2289) <= b;
    outputs(2290) <= a and not b;
    outputs(2291) <= not (a or b);
    outputs(2292) <= not (a or b);
    outputs(2293) <= a and not b;
    outputs(2294) <= not (a xor b);
    outputs(2295) <= a and b;
    outputs(2296) <= b;
    outputs(2297) <= not b;
    outputs(2298) <= not (a xor b);
    outputs(2299) <= b and not a;
    outputs(2300) <= b;
    outputs(2301) <= not (a xor b);
    outputs(2302) <= not b or a;
    outputs(2303) <= b and not a;
    outputs(2304) <= a xor b;
    outputs(2305) <= not a or b;
    outputs(2306) <= not (a and b);
    outputs(2307) <= not a;
    outputs(2308) <= a xor b;
    outputs(2309) <= a or b;
    outputs(2310) <= a;
    outputs(2311) <= a xor b;
    outputs(2312) <= not (a xor b);
    outputs(2313) <= a and b;
    outputs(2314) <= not (a or b);
    outputs(2315) <= not b;
    outputs(2316) <= b and not a;
    outputs(2317) <= not b or a;
    outputs(2318) <= b and not a;
    outputs(2319) <= not (a or b);
    outputs(2320) <= not b;
    outputs(2321) <= b and not a;
    outputs(2322) <= a and not b;
    outputs(2323) <= not (a xor b);
    outputs(2324) <= b and not a;
    outputs(2325) <= not (a or b);
    outputs(2326) <= b;
    outputs(2327) <= not (a or b);
    outputs(2328) <= a and not b;
    outputs(2329) <= not (a xor b);
    outputs(2330) <= a and b;
    outputs(2331) <= a and not b;
    outputs(2332) <= a or b;
    outputs(2333) <= b and not a;
    outputs(2334) <= not a;
    outputs(2335) <= b and not a;
    outputs(2336) <= a xor b;
    outputs(2337) <= a and not b;
    outputs(2338) <= b;
    outputs(2339) <= not (a or b);
    outputs(2340) <= not b;
    outputs(2341) <= a and b;
    outputs(2342) <= not b or a;
    outputs(2343) <= not (a or b);
    outputs(2344) <= not (a or b);
    outputs(2345) <= b and not a;
    outputs(2346) <= not (a or b);
    outputs(2347) <= a and b;
    outputs(2348) <= not a;
    outputs(2349) <= not a;
    outputs(2350) <= not b;
    outputs(2351) <= b and not a;
    outputs(2352) <= b and not a;
    outputs(2353) <= not a;
    outputs(2354) <= a xor b;
    outputs(2355) <= a xor b;
    outputs(2356) <= a and b;
    outputs(2357) <= b and not a;
    outputs(2358) <= not (a or b);
    outputs(2359) <= b and not a;
    outputs(2360) <= a and b;
    outputs(2361) <= b and not a;
    outputs(2362) <= not a;
    outputs(2363) <= b;
    outputs(2364) <= not a;
    outputs(2365) <= a and not b;
    outputs(2366) <= a;
    outputs(2367) <= not (a or b);
    outputs(2368) <= a xor b;
    outputs(2369) <= not b;
    outputs(2370) <= b and not a;
    outputs(2371) <= not b;
    outputs(2372) <= a and b;
    outputs(2373) <= not a;
    outputs(2374) <= not b;
    outputs(2375) <= a and b;
    outputs(2376) <= not (a or b);
    outputs(2377) <= b and not a;
    outputs(2378) <= a and b;
    outputs(2379) <= not (a or b);
    outputs(2380) <= not a or b;
    outputs(2381) <= a and b;
    outputs(2382) <= a and b;
    outputs(2383) <= not a;
    outputs(2384) <= b and not a;
    outputs(2385) <= not (a xor b);
    outputs(2386) <= b and not a;
    outputs(2387) <= not a;
    outputs(2388) <= b and not a;
    outputs(2389) <= b and not a;
    outputs(2390) <= a and b;
    outputs(2391) <= not a or b;
    outputs(2392) <= not (a or b);
    outputs(2393) <= a and b;
    outputs(2394) <= not (a or b);
    outputs(2395) <= a and b;
    outputs(2396) <= a and not b;
    outputs(2397) <= not (a or b);
    outputs(2398) <= not b;
    outputs(2399) <= a and not b;
    outputs(2400) <= not a;
    outputs(2401) <= not b;
    outputs(2402) <= a and b;
    outputs(2403) <= a;
    outputs(2404) <= a and b;
    outputs(2405) <= not (a or b);
    outputs(2406) <= a and not b;
    outputs(2407) <= a and b;
    outputs(2408) <= a and not b;
    outputs(2409) <= a and b;
    outputs(2410) <= a and b;
    outputs(2411) <= b and not a;
    outputs(2412) <= a;
    outputs(2413) <= a;
    outputs(2414) <= a;
    outputs(2415) <= not b;
    outputs(2416) <= b;
    outputs(2417) <= not (a or b);
    outputs(2418) <= a xor b;
    outputs(2419) <= not (a or b);
    outputs(2420) <= a;
    outputs(2421) <= b and not a;
    outputs(2422) <= a and not b;
    outputs(2423) <= b and not a;
    outputs(2424) <= not a;
    outputs(2425) <= a and not b;
    outputs(2426) <= not b;
    outputs(2427) <= not (a xor b);
    outputs(2428) <= a;
    outputs(2429) <= a;
    outputs(2430) <= a and b;
    outputs(2431) <= a and b;
    outputs(2432) <= b;
    outputs(2433) <= not b;
    outputs(2434) <= a and not b;
    outputs(2435) <= b;
    outputs(2436) <= b;
    outputs(2437) <= a and not b;
    outputs(2438) <= a xor b;
    outputs(2439) <= a and b;
    outputs(2440) <= b and not a;
    outputs(2441) <= a and b;
    outputs(2442) <= not (a and b);
    outputs(2443) <= b;
    outputs(2444) <= not (a or b);
    outputs(2445) <= a and not b;
    outputs(2446) <= not (a xor b);
    outputs(2447) <= not a;
    outputs(2448) <= b;
    outputs(2449) <= b and not a;
    outputs(2450) <= b;
    outputs(2451) <= a and b;
    outputs(2452) <= b and not a;
    outputs(2453) <= a and not b;
    outputs(2454) <= not (a or b);
    outputs(2455) <= not a;
    outputs(2456) <= b and not a;
    outputs(2457) <= a and not b;
    outputs(2458) <= not a;
    outputs(2459) <= not (a xor b);
    outputs(2460) <= a and b;
    outputs(2461) <= b and not a;
    outputs(2462) <= a and b;
    outputs(2463) <= b and not a;
    outputs(2464) <= a xor b;
    outputs(2465) <= b;
    outputs(2466) <= a and not b;
    outputs(2467) <= a and b;
    outputs(2468) <= not (a or b);
    outputs(2469) <= a and not b;
    outputs(2470) <= a and b;
    outputs(2471) <= a and not b;
    outputs(2472) <= not a;
    outputs(2473) <= a xor b;
    outputs(2474) <= b;
    outputs(2475) <= not (a and b);
    outputs(2476) <= b and not a;
    outputs(2477) <= a and not b;
    outputs(2478) <= not a;
    outputs(2479) <= not (a or b);
    outputs(2480) <= a and not b;
    outputs(2481) <= not b;
    outputs(2482) <= not b;
    outputs(2483) <= a;
    outputs(2484) <= a;
    outputs(2485) <= not b;
    outputs(2486) <= a and b;
    outputs(2487) <= not b;
    outputs(2488) <= not b;
    outputs(2489) <= not (a or b);
    outputs(2490) <= a and b;
    outputs(2491) <= a;
    outputs(2492) <= a and not b;
    outputs(2493) <= b;
    outputs(2494) <= b and not a;
    outputs(2495) <= not a;
    outputs(2496) <= a;
    outputs(2497) <= b and not a;
    outputs(2498) <= b and not a;
    outputs(2499) <= not a;
    outputs(2500) <= not (a or b);
    outputs(2501) <= not (a or b);
    outputs(2502) <= not a;
    outputs(2503) <= not a;
    outputs(2504) <= not a;
    outputs(2505) <= a xor b;
    outputs(2506) <= a and not b;
    outputs(2507) <= a and b;
    outputs(2508) <= a and b;
    outputs(2509) <= not (a xor b);
    outputs(2510) <= not a;
    outputs(2511) <= b and not a;
    outputs(2512) <= not a;
    outputs(2513) <= not a or b;
    outputs(2514) <= a or b;
    outputs(2515) <= not (a or b);
    outputs(2516) <= a;
    outputs(2517) <= not a;
    outputs(2518) <= a and b;
    outputs(2519) <= not (a xor b);
    outputs(2520) <= a and not b;
    outputs(2521) <= a and b;
    outputs(2522) <= not b;
    outputs(2523) <= not a;
    outputs(2524) <= not b;
    outputs(2525) <= a or b;
    outputs(2526) <= not (a xor b);
    outputs(2527) <= not b;
    outputs(2528) <= a and b;
    outputs(2529) <= a xor b;
    outputs(2530) <= a and b;
    outputs(2531) <= not a;
    outputs(2532) <= not (a or b);
    outputs(2533) <= a and not b;
    outputs(2534) <= b and not a;
    outputs(2535) <= a and not b;
    outputs(2536) <= a or b;
    outputs(2537) <= b and not a;
    outputs(2538) <= not b;
    outputs(2539) <= b and not a;
    outputs(2540) <= b;
    outputs(2541) <= not a;
    outputs(2542) <= not (a and b);
    outputs(2543) <= a xor b;
    outputs(2544) <= not (a or b);
    outputs(2545) <= not (a or b);
    outputs(2546) <= a and b;
    outputs(2547) <= a and b;
    outputs(2548) <= not (a xor b);
    outputs(2549) <= b and not a;
    outputs(2550) <= not (a xor b);
    outputs(2551) <= a and not b;
    outputs(2552) <= a;
    outputs(2553) <= a and not b;
    outputs(2554) <= a;
    outputs(2555) <= a and not b;
    outputs(2556) <= not (a or b);
    outputs(2557) <= a and not b;
    outputs(2558) <= not (a or b);
    outputs(2559) <= not (a or b);
end Behavioral;
