module logic_network(
    input wire [1023:0] inputs,
    output wire [9:0] outputs
);

    wire [2559:0] layer0_outputs;
    wire [2559:0] layer1_outputs;
    wire [2559:0] layer2_outputs;
    wire [2559:0] layer3_outputs;
    wire [2559:0] layer4_outputs;

    assign layer0_outputs[0] = ~(inputs[374]) | (inputs[830]);
    assign layer0_outputs[1] = (inputs[899]) & (inputs[643]);
    assign layer0_outputs[2] = ~((inputs[590]) ^ (inputs[564]));
    assign layer0_outputs[3] = inputs[528];
    assign layer0_outputs[4] = ~((inputs[571]) | (inputs[994]));
    assign layer0_outputs[5] = ~(inputs[72]);
    assign layer0_outputs[6] = (inputs[97]) | (inputs[732]);
    assign layer0_outputs[7] = ~(inputs[719]);
    assign layer0_outputs[8] = inputs[517];
    assign layer0_outputs[9] = ~(inputs[46]) | (inputs[323]);
    assign layer0_outputs[10] = (inputs[305]) | (inputs[1000]);
    assign layer0_outputs[11] = (inputs[147]) ^ (inputs[670]);
    assign layer0_outputs[12] = ~(inputs[853]);
    assign layer0_outputs[13] = ~(inputs[967]) | (inputs[147]);
    assign layer0_outputs[14] = (inputs[752]) & (inputs[454]);
    assign layer0_outputs[15] = ~((inputs[475]) & (inputs[35]));
    assign layer0_outputs[16] = (inputs[107]) ^ (inputs[626]);
    assign layer0_outputs[17] = ~((inputs[744]) ^ (inputs[932]));
    assign layer0_outputs[18] = ~(inputs[876]) | (inputs[543]);
    assign layer0_outputs[19] = ~((inputs[842]) & (inputs[713]));
    assign layer0_outputs[20] = ~((inputs[53]) & (inputs[318]));
    assign layer0_outputs[21] = ~(inputs[713]) | (inputs[234]);
    assign layer0_outputs[22] = inputs[594];
    assign layer0_outputs[23] = ~(inputs[270]) | (inputs[554]);
    assign layer0_outputs[24] = ~((inputs[976]) | (inputs[913]));
    assign layer0_outputs[25] = (inputs[717]) & ~(inputs[196]);
    assign layer0_outputs[26] = (inputs[824]) & ~(inputs[823]);
    assign layer0_outputs[27] = 1'b1;
    assign layer0_outputs[28] = ~(inputs[970]);
    assign layer0_outputs[29] = (inputs[338]) | (inputs[802]);
    assign layer0_outputs[30] = 1'b1;
    assign layer0_outputs[31] = ~(inputs[889]);
    assign layer0_outputs[32] = 1'b1;
    assign layer0_outputs[33] = ~((inputs[170]) | (inputs[503]));
    assign layer0_outputs[34] = 1'b0;
    assign layer0_outputs[35] = ~((inputs[655]) | (inputs[80]));
    assign layer0_outputs[36] = (inputs[481]) | (inputs[1021]);
    assign layer0_outputs[37] = (inputs[767]) | (inputs[887]);
    assign layer0_outputs[38] = ~(inputs[773]) | (inputs[30]);
    assign layer0_outputs[39] = 1'b1;
    assign layer0_outputs[40] = ~(inputs[392]) | (inputs[401]);
    assign layer0_outputs[41] = 1'b0;
    assign layer0_outputs[42] = ~(inputs[966]);
    assign layer0_outputs[43] = (inputs[758]) | (inputs[439]);
    assign layer0_outputs[44] = inputs[434];
    assign layer0_outputs[45] = (inputs[894]) & ~(inputs[161]);
    assign layer0_outputs[46] = ~(inputs[873]);
    assign layer0_outputs[47] = (inputs[553]) & ~(inputs[638]);
    assign layer0_outputs[48] = (inputs[312]) ^ (inputs[546]);
    assign layer0_outputs[49] = (inputs[192]) ^ (inputs[840]);
    assign layer0_outputs[50] = ~(inputs[950]) | (inputs[605]);
    assign layer0_outputs[51] = (inputs[504]) | (inputs[650]);
    assign layer0_outputs[52] = ~(inputs[374]) | (inputs[139]);
    assign layer0_outputs[53] = inputs[814];
    assign layer0_outputs[54] = ~(inputs[325]);
    assign layer0_outputs[55] = (inputs[682]) & ~(inputs[647]);
    assign layer0_outputs[56] = ~(inputs[740]);
    assign layer0_outputs[57] = ~(inputs[258]) | (inputs[881]);
    assign layer0_outputs[58] = 1'b1;
    assign layer0_outputs[59] = ~(inputs[946]) | (inputs[469]);
    assign layer0_outputs[60] = inputs[332];
    assign layer0_outputs[61] = 1'b1;
    assign layer0_outputs[62] = (inputs[560]) | (inputs[711]);
    assign layer0_outputs[63] = (inputs[660]) & (inputs[719]);
    assign layer0_outputs[64] = (inputs[462]) & ~(inputs[17]);
    assign layer0_outputs[65] = ~((inputs[877]) ^ (inputs[225]));
    assign layer0_outputs[66] = inputs[976];
    assign layer0_outputs[67] = (inputs[642]) & ~(inputs[442]);
    assign layer0_outputs[68] = (inputs[968]) ^ (inputs[523]);
    assign layer0_outputs[69] = ~((inputs[18]) | (inputs[384]));
    assign layer0_outputs[70] = inputs[974];
    assign layer0_outputs[71] = (inputs[520]) | (inputs[545]);
    assign layer0_outputs[72] = (inputs[660]) ^ (inputs[197]);
    assign layer0_outputs[73] = inputs[303];
    assign layer0_outputs[74] = ~(inputs[526]) | (inputs[513]);
    assign layer0_outputs[75] = ~((inputs[564]) | (inputs[79]));
    assign layer0_outputs[76] = ~((inputs[407]) | (inputs[668]));
    assign layer0_outputs[77] = ~((inputs[157]) ^ (inputs[654]));
    assign layer0_outputs[78] = ~((inputs[258]) | (inputs[653]));
    assign layer0_outputs[79] = ~((inputs[12]) | (inputs[619]));
    assign layer0_outputs[80] = ~(inputs[861]);
    assign layer0_outputs[81] = (inputs[462]) & (inputs[28]);
    assign layer0_outputs[82] = (inputs[283]) | (inputs[939]);
    assign layer0_outputs[83] = ~(inputs[938]);
    assign layer0_outputs[84] = ~((inputs[656]) | (inputs[453]));
    assign layer0_outputs[85] = (inputs[646]) & ~(inputs[334]);
    assign layer0_outputs[86] = ~((inputs[84]) ^ (inputs[203]));
    assign layer0_outputs[87] = ~((inputs[975]) & (inputs[291]));
    assign layer0_outputs[88] = inputs[314];
    assign layer0_outputs[89] = 1'b1;
    assign layer0_outputs[90] = (inputs[317]) & (inputs[785]);
    assign layer0_outputs[91] = inputs[918];
    assign layer0_outputs[92] = ~(inputs[514]) | (inputs[451]);
    assign layer0_outputs[93] = ~(inputs[374]) | (inputs[905]);
    assign layer0_outputs[94] = 1'b0;
    assign layer0_outputs[95] = ~(inputs[663]);
    assign layer0_outputs[96] = (inputs[858]) & ~(inputs[825]);
    assign layer0_outputs[97] = (inputs[177]) | (inputs[665]);
    assign layer0_outputs[98] = ~(inputs[1001]);
    assign layer0_outputs[99] = (inputs[860]) | (inputs[266]);
    assign layer0_outputs[100] = (inputs[470]) & ~(inputs[427]);
    assign layer0_outputs[101] = inputs[274];
    assign layer0_outputs[102] = (inputs[540]) | (inputs[587]);
    assign layer0_outputs[103] = (inputs[958]) & ~(inputs[952]);
    assign layer0_outputs[104] = ~((inputs[205]) ^ (inputs[289]));
    assign layer0_outputs[105] = ~(inputs[962]);
    assign layer0_outputs[106] = 1'b0;
    assign layer0_outputs[107] = (inputs[16]) & ~(inputs[573]);
    assign layer0_outputs[108] = 1'b0;
    assign layer0_outputs[109] = ~(inputs[202]) | (inputs[1012]);
    assign layer0_outputs[110] = ~(inputs[1007]) | (inputs[947]);
    assign layer0_outputs[111] = ~(inputs[204]);
    assign layer0_outputs[112] = inputs[492];
    assign layer0_outputs[113] = (inputs[89]) ^ (inputs[803]);
    assign layer0_outputs[114] = ~(inputs[840]) | (inputs[288]);
    assign layer0_outputs[115] = ~(inputs[618]);
    assign layer0_outputs[116] = ~(inputs[846]);
    assign layer0_outputs[117] = ~((inputs[573]) | (inputs[95]));
    assign layer0_outputs[118] = ~(inputs[93]);
    assign layer0_outputs[119] = (inputs[499]) & ~(inputs[25]);
    assign layer0_outputs[120] = ~(inputs[609]);
    assign layer0_outputs[121] = 1'b0;
    assign layer0_outputs[122] = (inputs[817]) & ~(inputs[1009]);
    assign layer0_outputs[123] = (inputs[466]) | (inputs[163]);
    assign layer0_outputs[124] = inputs[189];
    assign layer0_outputs[125] = inputs[811];
    assign layer0_outputs[126] = ~(inputs[560]);
    assign layer0_outputs[127] = (inputs[734]) ^ (inputs[111]);
    assign layer0_outputs[128] = (inputs[143]) & ~(inputs[894]);
    assign layer0_outputs[129] = (inputs[386]) & (inputs[91]);
    assign layer0_outputs[130] = ~(inputs[60]) | (inputs[244]);
    assign layer0_outputs[131] = ~((inputs[260]) | (inputs[259]));
    assign layer0_outputs[132] = ~((inputs[37]) | (inputs[691]));
    assign layer0_outputs[133] = inputs[593];
    assign layer0_outputs[134] = ~(inputs[357]);
    assign layer0_outputs[135] = ~((inputs[236]) ^ (inputs[451]));
    assign layer0_outputs[136] = 1'b1;
    assign layer0_outputs[137] = ~((inputs[325]) & (inputs[164]));
    assign layer0_outputs[138] = ~((inputs[935]) | (inputs[230]));
    assign layer0_outputs[139] = (inputs[805]) | (inputs[167]);
    assign layer0_outputs[140] = inputs[968];
    assign layer0_outputs[141] = (inputs[402]) & (inputs[1017]);
    assign layer0_outputs[142] = (inputs[836]) | (inputs[313]);
    assign layer0_outputs[143] = ~((inputs[280]) | (inputs[31]));
    assign layer0_outputs[144] = ~(inputs[227]) | (inputs[801]);
    assign layer0_outputs[145] = ~(inputs[365]) | (inputs[980]);
    assign layer0_outputs[146] = 1'b0;
    assign layer0_outputs[147] = ~((inputs[261]) | (inputs[29]));
    assign layer0_outputs[148] = ~((inputs[676]) & (inputs[419]));
    assign layer0_outputs[149] = 1'b0;
    assign layer0_outputs[150] = inputs[372];
    assign layer0_outputs[151] = ~(inputs[219]);
    assign layer0_outputs[152] = (inputs[870]) | (inputs[377]);
    assign layer0_outputs[153] = 1'b1;
    assign layer0_outputs[154] = 1'b0;
    assign layer0_outputs[155] = (inputs[910]) & ~(inputs[30]);
    assign layer0_outputs[156] = (inputs[200]) & (inputs[966]);
    assign layer0_outputs[157] = (inputs[212]) | (inputs[103]);
    assign layer0_outputs[158] = (inputs[598]) & ~(inputs[977]);
    assign layer0_outputs[159] = 1'b1;
    assign layer0_outputs[160] = ~(inputs[749]);
    assign layer0_outputs[161] = ~(inputs[117]);
    assign layer0_outputs[162] = ~(inputs[166]);
    assign layer0_outputs[163] = (inputs[902]) | (inputs[962]);
    assign layer0_outputs[164] = (inputs[763]) | (inputs[358]);
    assign layer0_outputs[165] = inputs[334];
    assign layer0_outputs[166] = (inputs[813]) & ~(inputs[39]);
    assign layer0_outputs[167] = (inputs[272]) & ~(inputs[149]);
    assign layer0_outputs[168] = ~((inputs[49]) | (inputs[573]));
    assign layer0_outputs[169] = 1'b0;
    assign layer0_outputs[170] = 1'b1;
    assign layer0_outputs[171] = ~(inputs[77]);
    assign layer0_outputs[172] = 1'b0;
    assign layer0_outputs[173] = ~(inputs[922]);
    assign layer0_outputs[174] = 1'b1;
    assign layer0_outputs[175] = ~((inputs[172]) | (inputs[698]));
    assign layer0_outputs[176] = ~(inputs[608]) | (inputs[108]);
    assign layer0_outputs[177] = inputs[265];
    assign layer0_outputs[178] = ~(inputs[850]);
    assign layer0_outputs[179] = inputs[419];
    assign layer0_outputs[180] = ~(inputs[529]) | (inputs[1011]);
    assign layer0_outputs[181] = (inputs[942]) & ~(inputs[159]);
    assign layer0_outputs[182] = inputs[243];
    assign layer0_outputs[183] = (inputs[790]) | (inputs[441]);
    assign layer0_outputs[184] = ~(inputs[275]) | (inputs[152]);
    assign layer0_outputs[185] = inputs[497];
    assign layer0_outputs[186] = 1'b1;
    assign layer0_outputs[187] = inputs[240];
    assign layer0_outputs[188] = 1'b1;
    assign layer0_outputs[189] = ~((inputs[597]) | (inputs[87]));
    assign layer0_outputs[190] = (inputs[255]) & ~(inputs[984]);
    assign layer0_outputs[191] = ~((inputs[49]) | (inputs[105]));
    assign layer0_outputs[192] = (inputs[772]) & (inputs[838]);
    assign layer0_outputs[193] = ~(inputs[759]);
    assign layer0_outputs[194] = 1'b0;
    assign layer0_outputs[195] = (inputs[476]) | (inputs[509]);
    assign layer0_outputs[196] = ~(inputs[728]);
    assign layer0_outputs[197] = ~((inputs[626]) | (inputs[951]));
    assign layer0_outputs[198] = (inputs[89]) & ~(inputs[997]);
    assign layer0_outputs[199] = (inputs[513]) ^ (inputs[649]);
    assign layer0_outputs[200] = ~(inputs[244]) | (inputs[832]);
    assign layer0_outputs[201] = inputs[112];
    assign layer0_outputs[202] = ~(inputs[940]);
    assign layer0_outputs[203] = (inputs[202]) & ~(inputs[393]);
    assign layer0_outputs[204] = ~(inputs[475]) | (inputs[356]);
    assign layer0_outputs[205] = ~(inputs[728]) | (inputs[474]);
    assign layer0_outputs[206] = ~(inputs[210]) | (inputs[955]);
    assign layer0_outputs[207] = (inputs[204]) | (inputs[712]);
    assign layer0_outputs[208] = (inputs[448]) & ~(inputs[166]);
    assign layer0_outputs[209] = ~(inputs[623]) | (inputs[468]);
    assign layer0_outputs[210] = 1'b1;
    assign layer0_outputs[211] = ~((inputs[777]) ^ (inputs[24]));
    assign layer0_outputs[212] = inputs[311];
    assign layer0_outputs[213] = ~(inputs[559]);
    assign layer0_outputs[214] = inputs[76];
    assign layer0_outputs[215] = inputs[468];
    assign layer0_outputs[216] = ~((inputs[927]) & (inputs[637]));
    assign layer0_outputs[217] = ~((inputs[328]) ^ (inputs[80]));
    assign layer0_outputs[218] = (inputs[337]) & (inputs[802]);
    assign layer0_outputs[219] = ~(inputs[336]) | (inputs[762]);
    assign layer0_outputs[220] = inputs[641];
    assign layer0_outputs[221] = ~(inputs[332]) | (inputs[675]);
    assign layer0_outputs[222] = (inputs[681]) & ~(inputs[701]);
    assign layer0_outputs[223] = 1'b0;
    assign layer0_outputs[224] = (inputs[221]) & ~(inputs[929]);
    assign layer0_outputs[225] = ~((inputs[978]) | (inputs[755]));
    assign layer0_outputs[226] = (inputs[873]) & (inputs[263]);
    assign layer0_outputs[227] = inputs[983];
    assign layer0_outputs[228] = (inputs[102]) & ~(inputs[926]);
    assign layer0_outputs[229] = ~((inputs[768]) & (inputs[1004]));
    assign layer0_outputs[230] = (inputs[507]) ^ (inputs[1018]);
    assign layer0_outputs[231] = (inputs[621]) | (inputs[521]);
    assign layer0_outputs[232] = ~((inputs[938]) ^ (inputs[121]));
    assign layer0_outputs[233] = ~((inputs[208]) | (inputs[480]));
    assign layer0_outputs[234] = inputs[567];
    assign layer0_outputs[235] = (inputs[370]) & ~(inputs[797]);
    assign layer0_outputs[236] = ~(inputs[692]) | (inputs[916]);
    assign layer0_outputs[237] = ~((inputs[717]) & (inputs[133]));
    assign layer0_outputs[238] = (inputs[408]) | (inputs[312]);
    assign layer0_outputs[239] = ~(inputs[635]);
    assign layer0_outputs[240] = ~(inputs[623]) | (inputs[877]);
    assign layer0_outputs[241] = ~((inputs[909]) | (inputs[566]));
    assign layer0_outputs[242] = 1'b0;
    assign layer0_outputs[243] = 1'b1;
    assign layer0_outputs[244] = (inputs[639]) & (inputs[1006]);
    assign layer0_outputs[245] = (inputs[356]) & (inputs[218]);
    assign layer0_outputs[246] = (inputs[97]) | (inputs[376]);
    assign layer0_outputs[247] = ~((inputs[1020]) ^ (inputs[293]));
    assign layer0_outputs[248] = ~(inputs[793]);
    assign layer0_outputs[249] = 1'b1;
    assign layer0_outputs[250] = 1'b0;
    assign layer0_outputs[251] = inputs[971];
    assign layer0_outputs[252] = ~((inputs[983]) | (inputs[855]));
    assign layer0_outputs[253] = (inputs[78]) & ~(inputs[215]);
    assign layer0_outputs[254] = ~(inputs[984]) | (inputs[842]);
    assign layer0_outputs[255] = ~((inputs[262]) ^ (inputs[257]));
    assign layer0_outputs[256] = ~(inputs[702]);
    assign layer0_outputs[257] = 1'b0;
    assign layer0_outputs[258] = ~(inputs[574]);
    assign layer0_outputs[259] = ~(inputs[636]);
    assign layer0_outputs[260] = (inputs[530]) & (inputs[722]);
    assign layer0_outputs[261] = ~(inputs[34]);
    assign layer0_outputs[262] = (inputs[562]) | (inputs[26]);
    assign layer0_outputs[263] = (inputs[823]) | (inputs[772]);
    assign layer0_outputs[264] = ~(inputs[936]);
    assign layer0_outputs[265] = ~(inputs[897]) | (inputs[661]);
    assign layer0_outputs[266] = inputs[422];
    assign layer0_outputs[267] = ~(inputs[21]);
    assign layer0_outputs[268] = ~((inputs[120]) | (inputs[179]));
    assign layer0_outputs[269] = (inputs[413]) | (inputs[942]);
    assign layer0_outputs[270] = inputs[594];
    assign layer0_outputs[271] = ~((inputs[988]) ^ (inputs[438]));
    assign layer0_outputs[272] = (inputs[858]) & ~(inputs[599]);
    assign layer0_outputs[273] = ~((inputs[296]) ^ (inputs[544]));
    assign layer0_outputs[274] = 1'b1;
    assign layer0_outputs[275] = inputs[687];
    assign layer0_outputs[276] = (inputs[937]) & (inputs[498]);
    assign layer0_outputs[277] = ~((inputs[342]) | (inputs[844]));
    assign layer0_outputs[278] = 1'b1;
    assign layer0_outputs[279] = ~((inputs[376]) | (inputs[334]));
    assign layer0_outputs[280] = ~(inputs[113]) | (inputs[832]);
    assign layer0_outputs[281] = ~(inputs[286]);
    assign layer0_outputs[282] = ~(inputs[29]) | (inputs[256]);
    assign layer0_outputs[283] = 1'b1;
    assign layer0_outputs[284] = inputs[947];
    assign layer0_outputs[285] = inputs[490];
    assign layer0_outputs[286] = inputs[961];
    assign layer0_outputs[287] = (inputs[571]) & ~(inputs[643]);
    assign layer0_outputs[288] = ~((inputs[378]) | (inputs[155]));
    assign layer0_outputs[289] = ~(inputs[815]);
    assign layer0_outputs[290] = ~(inputs[748]);
    assign layer0_outputs[291] = ~((inputs[451]) ^ (inputs[535]));
    assign layer0_outputs[292] = ~(inputs[17]) | (inputs[642]);
    assign layer0_outputs[293] = (inputs[1019]) & ~(inputs[492]);
    assign layer0_outputs[294] = ~(inputs[12]);
    assign layer0_outputs[295] = (inputs[447]) & ~(inputs[3]);
    assign layer0_outputs[296] = ~(inputs[421]);
    assign layer0_outputs[297] = 1'b0;
    assign layer0_outputs[298] = ~((inputs[391]) | (inputs[737]));
    assign layer0_outputs[299] = ~(inputs[837]) | (inputs[479]);
    assign layer0_outputs[300] = (inputs[338]) & ~(inputs[697]);
    assign layer0_outputs[301] = (inputs[204]) | (inputs[481]);
    assign layer0_outputs[302] = ~((inputs[209]) & (inputs[591]));
    assign layer0_outputs[303] = ~(inputs[440]);
    assign layer0_outputs[304] = (inputs[124]) & (inputs[521]);
    assign layer0_outputs[305] = inputs[893];
    assign layer0_outputs[306] = (inputs[686]) & (inputs[277]);
    assign layer0_outputs[307] = (inputs[910]) | (inputs[813]);
    assign layer0_outputs[308] = ~((inputs[120]) | (inputs[812]));
    assign layer0_outputs[309] = ~(inputs[979]);
    assign layer0_outputs[310] = ~(inputs[427]) | (inputs[460]);
    assign layer0_outputs[311] = ~((inputs[800]) ^ (inputs[912]));
    assign layer0_outputs[312] = (inputs[850]) & ~(inputs[796]);
    assign layer0_outputs[313] = ~(inputs[569]) | (inputs[126]);
    assign layer0_outputs[314] = ~((inputs[404]) | (inputs[612]));
    assign layer0_outputs[315] = inputs[359];
    assign layer0_outputs[316] = (inputs[89]) & ~(inputs[671]);
    assign layer0_outputs[317] = ~((inputs[1019]) ^ (inputs[154]));
    assign layer0_outputs[318] = (inputs[180]) & ~(inputs[448]);
    assign layer0_outputs[319] = inputs[219];
    assign layer0_outputs[320] = (inputs[688]) & ~(inputs[45]);
    assign layer0_outputs[321] = ~(inputs[135]);
    assign layer0_outputs[322] = (inputs[772]) & ~(inputs[375]);
    assign layer0_outputs[323] = (inputs[55]) & (inputs[671]);
    assign layer0_outputs[324] = ~(inputs[565]);
    assign layer0_outputs[325] = inputs[78];
    assign layer0_outputs[326] = ~(inputs[582]);
    assign layer0_outputs[327] = ~(inputs[307]);
    assign layer0_outputs[328] = inputs[915];
    assign layer0_outputs[329] = (inputs[51]) & (inputs[879]);
    assign layer0_outputs[330] = ~(inputs[231]);
    assign layer0_outputs[331] = (inputs[779]) ^ (inputs[126]);
    assign layer0_outputs[332] = 1'b0;
    assign layer0_outputs[333] = inputs[211];
    assign layer0_outputs[334] = (inputs[420]) & ~(inputs[652]);
    assign layer0_outputs[335] = (inputs[216]) & (inputs[228]);
    assign layer0_outputs[336] = (inputs[511]) | (inputs[322]);
    assign layer0_outputs[337] = 1'b0;
    assign layer0_outputs[338] = inputs[781];
    assign layer0_outputs[339] = (inputs[97]) | (inputs[90]);
    assign layer0_outputs[340] = 1'b1;
    assign layer0_outputs[341] = (inputs[658]) & ~(inputs[747]);
    assign layer0_outputs[342] = inputs[261];
    assign layer0_outputs[343] = inputs[654];
    assign layer0_outputs[344] = ~(inputs[2]) | (inputs[609]);
    assign layer0_outputs[345] = (inputs[872]) & ~(inputs[461]);
    assign layer0_outputs[346] = ~((inputs[317]) ^ (inputs[240]));
    assign layer0_outputs[347] = ~(inputs[462]) | (inputs[685]);
    assign layer0_outputs[348] = inputs[905];
    assign layer0_outputs[349] = ~(inputs[653]) | (inputs[981]);
    assign layer0_outputs[350] = inputs[127];
    assign layer0_outputs[351] = 1'b0;
    assign layer0_outputs[352] = ~(inputs[717]);
    assign layer0_outputs[353] = ~((inputs[924]) | (inputs[692]));
    assign layer0_outputs[354] = (inputs[512]) ^ (inputs[85]);
    assign layer0_outputs[355] = inputs[186];
    assign layer0_outputs[356] = 1'b1;
    assign layer0_outputs[357] = ~((inputs[782]) & (inputs[590]));
    assign layer0_outputs[358] = ~(inputs[590]);
    assign layer0_outputs[359] = inputs[477];
    assign layer0_outputs[360] = inputs[239];
    assign layer0_outputs[361] = ~(inputs[955]);
    assign layer0_outputs[362] = ~(inputs[459]);
    assign layer0_outputs[363] = (inputs[713]) & (inputs[174]);
    assign layer0_outputs[364] = (inputs[501]) & ~(inputs[606]);
    assign layer0_outputs[365] = (inputs[391]) ^ (inputs[133]);
    assign layer0_outputs[366] = ~(inputs[18]) | (inputs[69]);
    assign layer0_outputs[367] = ~(inputs[381]) | (inputs[862]);
    assign layer0_outputs[368] = (inputs[55]) & ~(inputs[990]);
    assign layer0_outputs[369] = (inputs[872]) & ~(inputs[786]);
    assign layer0_outputs[370] = 1'b0;
    assign layer0_outputs[371] = ~(inputs[397]);
    assign layer0_outputs[372] = ~((inputs[661]) | (inputs[992]));
    assign layer0_outputs[373] = 1'b1;
    assign layer0_outputs[374] = ~((inputs[679]) & (inputs[222]));
    assign layer0_outputs[375] = (inputs[302]) | (inputs[57]);
    assign layer0_outputs[376] = inputs[62];
    assign layer0_outputs[377] = inputs[218];
    assign layer0_outputs[378] = inputs[593];
    assign layer0_outputs[379] = ~(inputs[333]) | (inputs[367]);
    assign layer0_outputs[380] = ~(inputs[527]);
    assign layer0_outputs[381] = ~((inputs[773]) | (inputs[709]));
    assign layer0_outputs[382] = 1'b0;
    assign layer0_outputs[383] = inputs[491];
    assign layer0_outputs[384] = ~(inputs[544]) | (inputs[930]);
    assign layer0_outputs[385] = 1'b1;
    assign layer0_outputs[386] = (inputs[969]) | (inputs[34]);
    assign layer0_outputs[387] = ~(inputs[847]) | (inputs[142]);
    assign layer0_outputs[388] = 1'b0;
    assign layer0_outputs[389] = ~(inputs[200]);
    assign layer0_outputs[390] = ~(inputs[815]);
    assign layer0_outputs[391] = ~((inputs[268]) & (inputs[790]));
    assign layer0_outputs[392] = ~(inputs[544]) | (inputs[664]);
    assign layer0_outputs[393] = 1'b1;
    assign layer0_outputs[394] = 1'b1;
    assign layer0_outputs[395] = ~((inputs[579]) ^ (inputs[410]));
    assign layer0_outputs[396] = (inputs[395]) & (inputs[875]);
    assign layer0_outputs[397] = ~((inputs[1017]) & (inputs[992]));
    assign layer0_outputs[398] = ~((inputs[1007]) | (inputs[251]));
    assign layer0_outputs[399] = ~(inputs[960]);
    assign layer0_outputs[400] = inputs[708];
    assign layer0_outputs[401] = (inputs[796]) ^ (inputs[252]);
    assign layer0_outputs[402] = ~(inputs[197]);
    assign layer0_outputs[403] = ~(inputs[680]);
    assign layer0_outputs[404] = (inputs[564]) & ~(inputs[458]);
    assign layer0_outputs[405] = ~((inputs[970]) | (inputs[861]));
    assign layer0_outputs[406] = 1'b1;
    assign layer0_outputs[407] = ~(inputs[562]);
    assign layer0_outputs[408] = ~(inputs[414]) | (inputs[265]);
    assign layer0_outputs[409] = inputs[621];
    assign layer0_outputs[410] = ~(inputs[987]) | (inputs[180]);
    assign layer0_outputs[411] = (inputs[748]) | (inputs[354]);
    assign layer0_outputs[412] = (inputs[698]) & (inputs[214]);
    assign layer0_outputs[413] = ~(inputs[34]) | (inputs[190]);
    assign layer0_outputs[414] = inputs[963];
    assign layer0_outputs[415] = (inputs[224]) | (inputs[29]);
    assign layer0_outputs[416] = inputs[684];
    assign layer0_outputs[417] = ~(inputs[628]);
    assign layer0_outputs[418] = inputs[185];
    assign layer0_outputs[419] = (inputs[689]) & ~(inputs[287]);
    assign layer0_outputs[420] = ~(inputs[758]) | (inputs[885]);
    assign layer0_outputs[421] = (inputs[349]) & ~(inputs[20]);
    assign layer0_outputs[422] = ~((inputs[354]) ^ (inputs[416]));
    assign layer0_outputs[423] = inputs[213];
    assign layer0_outputs[424] = (inputs[245]) & ~(inputs[978]);
    assign layer0_outputs[425] = ~(inputs[682]) | (inputs[923]);
    assign layer0_outputs[426] = (inputs[382]) & (inputs[292]);
    assign layer0_outputs[427] = ~((inputs[710]) & (inputs[76]));
    assign layer0_outputs[428] = ~(inputs[685]);
    assign layer0_outputs[429] = ~((inputs[457]) | (inputs[912]));
    assign layer0_outputs[430] = inputs[668];
    assign layer0_outputs[431] = (inputs[343]) & ~(inputs[81]);
    assign layer0_outputs[432] = ~((inputs[795]) | (inputs[606]));
    assign layer0_outputs[433] = ~(inputs[928]) | (inputs[350]);
    assign layer0_outputs[434] = ~(inputs[460]);
    assign layer0_outputs[435] = (inputs[501]) & ~(inputs[281]);
    assign layer0_outputs[436] = 1'b0;
    assign layer0_outputs[437] = ~((inputs[841]) & (inputs[514]));
    assign layer0_outputs[438] = ~(inputs[998]) | (inputs[324]);
    assign layer0_outputs[439] = (inputs[435]) & ~(inputs[450]);
    assign layer0_outputs[440] = ~((inputs[714]) ^ (inputs[4]));
    assign layer0_outputs[441] = 1'b1;
    assign layer0_outputs[442] = (inputs[829]) ^ (inputs[727]);
    assign layer0_outputs[443] = ~(inputs[709]) | (inputs[925]);
    assign layer0_outputs[444] = ~(inputs[742]) | (inputs[121]);
    assign layer0_outputs[445] = (inputs[269]) & ~(inputs[42]);
    assign layer0_outputs[446] = inputs[56];
    assign layer0_outputs[447] = ~(inputs[306]);
    assign layer0_outputs[448] = ~(inputs[522]);
    assign layer0_outputs[449] = ~((inputs[37]) ^ (inputs[143]));
    assign layer0_outputs[450] = ~((inputs[971]) | (inputs[301]));
    assign layer0_outputs[451] = ~(inputs[164]) | (inputs[322]);
    assign layer0_outputs[452] = 1'b1;
    assign layer0_outputs[453] = (inputs[472]) & ~(inputs[983]);
    assign layer0_outputs[454] = (inputs[804]) & ~(inputs[444]);
    assign layer0_outputs[455] = 1'b0;
    assign layer0_outputs[456] = inputs[667];
    assign layer0_outputs[457] = inputs[525];
    assign layer0_outputs[458] = inputs[400];
    assign layer0_outputs[459] = ~(inputs[679]) | (inputs[102]);
    assign layer0_outputs[460] = ~(inputs[718]);
    assign layer0_outputs[461] = (inputs[620]) | (inputs[153]);
    assign layer0_outputs[462] = 1'b1;
    assign layer0_outputs[463] = inputs[764];
    assign layer0_outputs[464] = ~(inputs[778]);
    assign layer0_outputs[465] = ~(inputs[594]);
    assign layer0_outputs[466] = ~((inputs[101]) | (inputs[136]));
    assign layer0_outputs[467] = ~((inputs[589]) ^ (inputs[17]));
    assign layer0_outputs[468] = inputs[503];
    assign layer0_outputs[469] = ~(inputs[264]);
    assign layer0_outputs[470] = ~((inputs[353]) & (inputs[504]));
    assign layer0_outputs[471] = 1'b0;
    assign layer0_outputs[472] = (inputs[139]) & (inputs[133]);
    assign layer0_outputs[473] = (inputs[526]) | (inputs[698]);
    assign layer0_outputs[474] = ~((inputs[295]) | (inputs[699]));
    assign layer0_outputs[475] = (inputs[439]) & ~(inputs[770]);
    assign layer0_outputs[476] = ~(inputs[415]) | (inputs[504]);
    assign layer0_outputs[477] = inputs[285];
    assign layer0_outputs[478] = inputs[237];
    assign layer0_outputs[479] = ~((inputs[159]) | (inputs[474]));
    assign layer0_outputs[480] = ~(inputs[830]);
    assign layer0_outputs[481] = 1'b0;
    assign layer0_outputs[482] = (inputs[549]) | (inputs[317]);
    assign layer0_outputs[483] = (inputs[987]) & ~(inputs[21]);
    assign layer0_outputs[484] = inputs[902];
    assign layer0_outputs[485] = ~(inputs[431]);
    assign layer0_outputs[486] = inputs[591];
    assign layer0_outputs[487] = (inputs[282]) | (inputs[251]);
    assign layer0_outputs[488] = (inputs[780]) ^ (inputs[959]);
    assign layer0_outputs[489] = 1'b0;
    assign layer0_outputs[490] = ~((inputs[1004]) & (inputs[236]));
    assign layer0_outputs[491] = ~((inputs[323]) | (inputs[337]));
    assign layer0_outputs[492] = inputs[310];
    assign layer0_outputs[493] = 1'b0;
    assign layer0_outputs[494] = ~(inputs[241]) | (inputs[870]);
    assign layer0_outputs[495] = inputs[519];
    assign layer0_outputs[496] = (inputs[362]) | (inputs[134]);
    assign layer0_outputs[497] = (inputs[595]) & ~(inputs[87]);
    assign layer0_outputs[498] = inputs[439];
    assign layer0_outputs[499] = ~(inputs[599]);
    assign layer0_outputs[500] = (inputs[640]) | (inputs[725]);
    assign layer0_outputs[501] = ~((inputs[842]) | (inputs[819]));
    assign layer0_outputs[502] = (inputs[878]) & ~(inputs[440]);
    assign layer0_outputs[503] = 1'b0;
    assign layer0_outputs[504] = ~((inputs[538]) | (inputs[24]));
    assign layer0_outputs[505] = 1'b0;
    assign layer0_outputs[506] = inputs[894];
    assign layer0_outputs[507] = ~(inputs[246]) | (inputs[196]);
    assign layer0_outputs[508] = ~(inputs[238]);
    assign layer0_outputs[509] = (inputs[316]) | (inputs[872]);
    assign layer0_outputs[510] = (inputs[983]) & (inputs[884]);
    assign layer0_outputs[511] = (inputs[82]) ^ (inputs[240]);
    assign layer0_outputs[512] = (inputs[750]) & (inputs[109]);
    assign layer0_outputs[513] = ~(inputs[615]) | (inputs[869]);
    assign layer0_outputs[514] = ~(inputs[60]) | (inputs[1005]);
    assign layer0_outputs[515] = 1'b1;
    assign layer0_outputs[516] = (inputs[781]) | (inputs[296]);
    assign layer0_outputs[517] = 1'b0;
    assign layer0_outputs[518] = ~((inputs[849]) & (inputs[443]));
    assign layer0_outputs[519] = (inputs[198]) & ~(inputs[434]);
    assign layer0_outputs[520] = inputs[726];
    assign layer0_outputs[521] = 1'b0;
    assign layer0_outputs[522] = ~(inputs[491]);
    assign layer0_outputs[523] = (inputs[227]) & (inputs[551]);
    assign layer0_outputs[524] = ~(inputs[490]);
    assign layer0_outputs[525] = (inputs[316]) | (inputs[945]);
    assign layer0_outputs[526] = ~(inputs[914]);
    assign layer0_outputs[527] = ~((inputs[908]) | (inputs[85]));
    assign layer0_outputs[528] = (inputs[556]) & ~(inputs[388]);
    assign layer0_outputs[529] = (inputs[391]) & ~(inputs[49]);
    assign layer0_outputs[530] = (inputs[868]) | (inputs[523]);
    assign layer0_outputs[531] = ~(inputs[282]);
    assign layer0_outputs[532] = (inputs[430]) | (inputs[575]);
    assign layer0_outputs[533] = ~((inputs[495]) | (inputs[314]));
    assign layer0_outputs[534] = (inputs[592]) & ~(inputs[895]);
    assign layer0_outputs[535] = ~((inputs[105]) ^ (inputs[348]));
    assign layer0_outputs[536] = ~(inputs[823]) | (inputs[448]);
    assign layer0_outputs[537] = (inputs[954]) & ~(inputs[380]);
    assign layer0_outputs[538] = (inputs[201]) & (inputs[247]);
    assign layer0_outputs[539] = ~(inputs[557]) | (inputs[203]);
    assign layer0_outputs[540] = (inputs[37]) & ~(inputs[833]);
    assign layer0_outputs[541] = ~((inputs[794]) | (inputs[755]));
    assign layer0_outputs[542] = 1'b0;
    assign layer0_outputs[543] = (inputs[292]) | (inputs[79]);
    assign layer0_outputs[544] = ~(inputs[991]);
    assign layer0_outputs[545] = (inputs[638]) & (inputs[738]);
    assign layer0_outputs[546] = ~((inputs[645]) & (inputs[27]));
    assign layer0_outputs[547] = 1'b1;
    assign layer0_outputs[548] = (inputs[904]) & (inputs[233]);
    assign layer0_outputs[549] = inputs[807];
    assign layer0_outputs[550] = ~(inputs[656]);
    assign layer0_outputs[551] = ~((inputs[207]) | (inputs[229]));
    assign layer0_outputs[552] = (inputs[973]) & ~(inputs[135]);
    assign layer0_outputs[553] = ~(inputs[83]);
    assign layer0_outputs[554] = (inputs[668]) | (inputs[238]);
    assign layer0_outputs[555] = (inputs[535]) & ~(inputs[535]);
    assign layer0_outputs[556] = ~((inputs[715]) | (inputs[79]));
    assign layer0_outputs[557] = ~(inputs[989]) | (inputs[633]);
    assign layer0_outputs[558] = ~(inputs[438]);
    assign layer0_outputs[559] = ~(inputs[930]);
    assign layer0_outputs[560] = ~((inputs[143]) & (inputs[965]));
    assign layer0_outputs[561] = 1'b1;
    assign layer0_outputs[562] = (inputs[247]) & ~(inputs[403]);
    assign layer0_outputs[563] = 1'b0;
    assign layer0_outputs[564] = inputs[547];
    assign layer0_outputs[565] = (inputs[216]) & ~(inputs[959]);
    assign layer0_outputs[566] = ~(inputs[296]) | (inputs[925]);
    assign layer0_outputs[567] = ~(inputs[972]) | (inputs[681]);
    assign layer0_outputs[568] = ~((inputs[685]) & (inputs[707]));
    assign layer0_outputs[569] = (inputs[549]) | (inputs[112]);
    assign layer0_outputs[570] = ~(inputs[631]);
    assign layer0_outputs[571] = ~(inputs[131]);
    assign layer0_outputs[572] = (inputs[237]) & ~(inputs[548]);
    assign layer0_outputs[573] = (inputs[118]) | (inputs[607]);
    assign layer0_outputs[574] = ~(inputs[116]);
    assign layer0_outputs[575] = inputs[210];
    assign layer0_outputs[576] = ~(inputs[492]);
    assign layer0_outputs[577] = ~(inputs[239]) | (inputs[146]);
    assign layer0_outputs[578] = ~(inputs[426]);
    assign layer0_outputs[579] = (inputs[123]) | (inputs[306]);
    assign layer0_outputs[580] = (inputs[651]) & (inputs[310]);
    assign layer0_outputs[581] = inputs[686];
    assign layer0_outputs[582] = 1'b0;
    assign layer0_outputs[583] = (inputs[793]) & ~(inputs[293]);
    assign layer0_outputs[584] = (inputs[264]) ^ (inputs[280]);
    assign layer0_outputs[585] = ~((inputs[106]) | (inputs[751]));
    assign layer0_outputs[586] = ~(inputs[491]) | (inputs[484]);
    assign layer0_outputs[587] = 1'b0;
    assign layer0_outputs[588] = 1'b0;
    assign layer0_outputs[589] = ~((inputs[517]) | (inputs[347]));
    assign layer0_outputs[590] = ~(inputs[627]) | (inputs[586]);
    assign layer0_outputs[591] = inputs[788];
    assign layer0_outputs[592] = ~((inputs[908]) | (inputs[923]));
    assign layer0_outputs[593] = (inputs[373]) & ~(inputs[36]);
    assign layer0_outputs[594] = ~(inputs[878]);
    assign layer0_outputs[595] = 1'b1;
    assign layer0_outputs[596] = inputs[397];
    assign layer0_outputs[597] = 1'b1;
    assign layer0_outputs[598] = (inputs[493]) | (inputs[326]);
    assign layer0_outputs[599] = ~((inputs[377]) | (inputs[260]));
    assign layer0_outputs[600] = ~(inputs[65]) | (inputs[985]);
    assign layer0_outputs[601] = ~(inputs[939]);
    assign layer0_outputs[602] = 1'b0;
    assign layer0_outputs[603] = ~((inputs[387]) | (inputs[804]));
    assign layer0_outputs[604] = (inputs[484]) | (inputs[880]);
    assign layer0_outputs[605] = (inputs[522]) & ~(inputs[351]);
    assign layer0_outputs[606] = ~(inputs[656]);
    assign layer0_outputs[607] = ~((inputs[132]) & (inputs[298]));
    assign layer0_outputs[608] = (inputs[229]) & (inputs[532]);
    assign layer0_outputs[609] = ~(inputs[655]);
    assign layer0_outputs[610] = inputs[496];
    assign layer0_outputs[611] = (inputs[414]) & (inputs[776]);
    assign layer0_outputs[612] = ~((inputs[929]) & (inputs[493]));
    assign layer0_outputs[613] = ~((inputs[637]) | (inputs[137]));
    assign layer0_outputs[614] = ~((inputs[63]) | (inputs[630]));
    assign layer0_outputs[615] = (inputs[159]) & ~(inputs[54]);
    assign layer0_outputs[616] = (inputs[138]) ^ (inputs[657]);
    assign layer0_outputs[617] = ~(inputs[27]);
    assign layer0_outputs[618] = 1'b1;
    assign layer0_outputs[619] = (inputs[364]) & ~(inputs[165]);
    assign layer0_outputs[620] = ~(inputs[35]) | (inputs[738]);
    assign layer0_outputs[621] = 1'b1;
    assign layer0_outputs[622] = (inputs[737]) & ~(inputs[692]);
    assign layer0_outputs[623] = (inputs[100]) ^ (inputs[206]);
    assign layer0_outputs[624] = (inputs[274]) & ~(inputs[177]);
    assign layer0_outputs[625] = inputs[884];
    assign layer0_outputs[626] = ~((inputs[883]) & (inputs[411]));
    assign layer0_outputs[627] = ~((inputs[188]) | (inputs[688]));
    assign layer0_outputs[628] = 1'b1;
    assign layer0_outputs[629] = inputs[554];
    assign layer0_outputs[630] = inputs[388];
    assign layer0_outputs[631] = ~(inputs[300]);
    assign layer0_outputs[632] = 1'b1;
    assign layer0_outputs[633] = ~((inputs[863]) | (inputs[140]));
    assign layer0_outputs[634] = (inputs[977]) | (inputs[533]);
    assign layer0_outputs[635] = ~(inputs[988]);
    assign layer0_outputs[636] = (inputs[83]) & (inputs[423]);
    assign layer0_outputs[637] = ~(inputs[446]);
    assign layer0_outputs[638] = 1'b0;
    assign layer0_outputs[639] = ~(inputs[407]);
    assign layer0_outputs[640] = ~((inputs[886]) | (inputs[486]));
    assign layer0_outputs[641] = 1'b1;
    assign layer0_outputs[642] = ~((inputs[406]) | (inputs[9]));
    assign layer0_outputs[643] = ~((inputs[682]) ^ (inputs[57]));
    assign layer0_outputs[644] = inputs[621];
    assign layer0_outputs[645] = inputs[78];
    assign layer0_outputs[646] = (inputs[694]) & ~(inputs[898]);
    assign layer0_outputs[647] = ~(inputs[332]);
    assign layer0_outputs[648] = inputs[454];
    assign layer0_outputs[649] = (inputs[40]) | (inputs[705]);
    assign layer0_outputs[650] = inputs[378];
    assign layer0_outputs[651] = ~(inputs[815]) | (inputs[761]);
    assign layer0_outputs[652] = (inputs[270]) | (inputs[54]);
    assign layer0_outputs[653] = (inputs[950]) & ~(inputs[253]);
    assign layer0_outputs[654] = (inputs[154]) | (inputs[582]);
    assign layer0_outputs[655] = (inputs[740]) | (inputs[93]);
    assign layer0_outputs[656] = ~((inputs[603]) ^ (inputs[381]));
    assign layer0_outputs[657] = (inputs[478]) ^ (inputs[940]);
    assign layer0_outputs[658] = inputs[843];
    assign layer0_outputs[659] = inputs[865];
    assign layer0_outputs[660] = 1'b0;
    assign layer0_outputs[661] = ~(inputs[444]) | (inputs[383]);
    assign layer0_outputs[662] = (inputs[348]) & (inputs[773]);
    assign layer0_outputs[663] = inputs[584];
    assign layer0_outputs[664] = (inputs[341]) | (inputs[611]);
    assign layer0_outputs[665] = ~(inputs[700]) | (inputs[973]);
    assign layer0_outputs[666] = 1'b1;
    assign layer0_outputs[667] = ~((inputs[789]) ^ (inputs[578]));
    assign layer0_outputs[668] = ~(inputs[376]);
    assign layer0_outputs[669] = ~(inputs[528]);
    assign layer0_outputs[670] = ~(inputs[336]) | (inputs[543]);
    assign layer0_outputs[671] = inputs[464];
    assign layer0_outputs[672] = (inputs[763]) & (inputs[247]);
    assign layer0_outputs[673] = inputs[366];
    assign layer0_outputs[674] = ~(inputs[856]);
    assign layer0_outputs[675] = ~(inputs[206]) | (inputs[284]);
    assign layer0_outputs[676] = inputs[62];
    assign layer0_outputs[677] = (inputs[775]) | (inputs[828]);
    assign layer0_outputs[678] = (inputs[791]) & (inputs[580]);
    assign layer0_outputs[679] = (inputs[789]) ^ (inputs[225]);
    assign layer0_outputs[680] = ~((inputs[350]) & (inputs[928]));
    assign layer0_outputs[681] = (inputs[160]) & (inputs[91]);
    assign layer0_outputs[682] = (inputs[361]) | (inputs[522]);
    assign layer0_outputs[683] = ~(inputs[583]) | (inputs[494]);
    assign layer0_outputs[684] = ~(inputs[767]);
    assign layer0_outputs[685] = (inputs[584]) & ~(inputs[641]);
    assign layer0_outputs[686] = ~((inputs[102]) | (inputs[840]));
    assign layer0_outputs[687] = ~(inputs[187]) | (inputs[482]);
    assign layer0_outputs[688] = (inputs[558]) & (inputs[421]);
    assign layer0_outputs[689] = ~(inputs[40]);
    assign layer0_outputs[690] = ~(inputs[635]);
    assign layer0_outputs[691] = ~((inputs[343]) | (inputs[379]));
    assign layer0_outputs[692] = (inputs[7]) | (inputs[1018]);
    assign layer0_outputs[693] = ~((inputs[736]) & (inputs[223]));
    assign layer0_outputs[694] = (inputs[768]) ^ (inputs[439]);
    assign layer0_outputs[695] = inputs[378];
    assign layer0_outputs[696] = ~(inputs[233]);
    assign layer0_outputs[697] = inputs[787];
    assign layer0_outputs[698] = ~(inputs[1001]);
    assign layer0_outputs[699] = ~(inputs[581]);
    assign layer0_outputs[700] = ~((inputs[30]) & (inputs[119]));
    assign layer0_outputs[701] = (inputs[876]) ^ (inputs[979]);
    assign layer0_outputs[702] = ~(inputs[342]) | (inputs[52]);
    assign layer0_outputs[703] = 1'b1;
    assign layer0_outputs[704] = ~(inputs[901]);
    assign layer0_outputs[705] = ~((inputs[707]) | (inputs[965]));
    assign layer0_outputs[706] = ~((inputs[724]) | (inputs[676]));
    assign layer0_outputs[707] = (inputs[603]) ^ (inputs[315]);
    assign layer0_outputs[708] = ~(inputs[224]) | (inputs[220]);
    assign layer0_outputs[709] = (inputs[926]) & ~(inputs[961]);
    assign layer0_outputs[710] = (inputs[619]) & ~(inputs[780]);
    assign layer0_outputs[711] = 1'b1;
    assign layer0_outputs[712] = ~(inputs[57]);
    assign layer0_outputs[713] = (inputs[967]) & ~(inputs[710]);
    assign layer0_outputs[714] = ~((inputs[252]) ^ (inputs[831]));
    assign layer0_outputs[715] = (inputs[150]) | (inputs[554]);
    assign layer0_outputs[716] = (inputs[792]) & ~(inputs[90]);
    assign layer0_outputs[717] = 1'b0;
    assign layer0_outputs[718] = ~((inputs[794]) | (inputs[682]));
    assign layer0_outputs[719] = ~(inputs[624]) | (inputs[426]);
    assign layer0_outputs[720] = ~(inputs[178]) | (inputs[633]);
    assign layer0_outputs[721] = ~(inputs[778]);
    assign layer0_outputs[722] = (inputs[723]) ^ (inputs[853]);
    assign layer0_outputs[723] = (inputs[697]) & ~(inputs[916]);
    assign layer0_outputs[724] = (inputs[287]) & (inputs[925]);
    assign layer0_outputs[725] = (inputs[156]) | (inputs[754]);
    assign layer0_outputs[726] = ~((inputs[308]) ^ (inputs[796]));
    assign layer0_outputs[727] = (inputs[921]) | (inputs[589]);
    assign layer0_outputs[728] = ~(inputs[984]) | (inputs[925]);
    assign layer0_outputs[729] = (inputs[702]) & (inputs[413]);
    assign layer0_outputs[730] = inputs[797];
    assign layer0_outputs[731] = inputs[524];
    assign layer0_outputs[732] = (inputs[200]) | (inputs[371]);
    assign layer0_outputs[733] = ~(inputs[819]);
    assign layer0_outputs[734] = ~(inputs[678]);
    assign layer0_outputs[735] = ~(inputs[247]);
    assign layer0_outputs[736] = ~((inputs[437]) | (inputs[195]));
    assign layer0_outputs[737] = 1'b1;
    assign layer0_outputs[738] = (inputs[583]) | (inputs[341]);
    assign layer0_outputs[739] = inputs[816];
    assign layer0_outputs[740] = ~(inputs[287]);
    assign layer0_outputs[741] = (inputs[1023]) & ~(inputs[532]);
    assign layer0_outputs[742] = ~(inputs[1000]) | (inputs[255]);
    assign layer0_outputs[743] = (inputs[380]) & ~(inputs[217]);
    assign layer0_outputs[744] = ~(inputs[147]) | (inputs[198]);
    assign layer0_outputs[745] = ~(inputs[824]) | (inputs[820]);
    assign layer0_outputs[746] = ~(inputs[982]) | (inputs[916]);
    assign layer0_outputs[747] = 1'b0;
    assign layer0_outputs[748] = (inputs[290]) ^ (inputs[208]);
    assign layer0_outputs[749] = ~(inputs[259]);
    assign layer0_outputs[750] = (inputs[403]) | (inputs[99]);
    assign layer0_outputs[751] = (inputs[393]) ^ (inputs[10]);
    assign layer0_outputs[752] = (inputs[641]) | (inputs[969]);
    assign layer0_outputs[753] = (inputs[288]) & ~(inputs[855]);
    assign layer0_outputs[754] = ~(inputs[192]) | (inputs[422]);
    assign layer0_outputs[755] = (inputs[962]) & (inputs[576]);
    assign layer0_outputs[756] = ~(inputs[821]) | (inputs[894]);
    assign layer0_outputs[757] = (inputs[484]) & ~(inputs[19]);
    assign layer0_outputs[758] = (inputs[162]) | (inputs[973]);
    assign layer0_outputs[759] = (inputs[964]) & ~(inputs[19]);
    assign layer0_outputs[760] = 1'b0;
    assign layer0_outputs[761] = inputs[186];
    assign layer0_outputs[762] = ~(inputs[725]) | (inputs[1022]);
    assign layer0_outputs[763] = 1'b0;
    assign layer0_outputs[764] = ~(inputs[75]);
    assign layer0_outputs[765] = inputs[283];
    assign layer0_outputs[766] = ~(inputs[142]);
    assign layer0_outputs[767] = 1'b0;
    assign layer0_outputs[768] = (inputs[322]) & (inputs[896]);
    assign layer0_outputs[769] = ~((inputs[18]) ^ (inputs[750]));
    assign layer0_outputs[770] = (inputs[368]) & (inputs[197]);
    assign layer0_outputs[771] = (inputs[644]) & ~(inputs[474]);
    assign layer0_outputs[772] = inputs[247];
    assign layer0_outputs[773] = ~((inputs[117]) ^ (inputs[672]));
    assign layer0_outputs[774] = ~((inputs[541]) & (inputs[302]));
    assign layer0_outputs[775] = ~((inputs[966]) | (inputs[703]));
    assign layer0_outputs[776] = ~(inputs[255]) | (inputs[502]);
    assign layer0_outputs[777] = (inputs[923]) & ~(inputs[757]);
    assign layer0_outputs[778] = ~((inputs[118]) | (inputs[720]));
    assign layer0_outputs[779] = inputs[648];
    assign layer0_outputs[780] = ~((inputs[378]) | (inputs[854]));
    assign layer0_outputs[781] = ~(inputs[435]) | (inputs[495]);
    assign layer0_outputs[782] = ~(inputs[769]) | (inputs[709]);
    assign layer0_outputs[783] = (inputs[503]) | (inputs[617]);
    assign layer0_outputs[784] = (inputs[673]) ^ (inputs[285]);
    assign layer0_outputs[785] = ~((inputs[796]) & (inputs[857]));
    assign layer0_outputs[786] = ~(inputs[180]);
    assign layer0_outputs[787] = ~((inputs[628]) | (inputs[251]));
    assign layer0_outputs[788] = (inputs[760]) ^ (inputs[412]);
    assign layer0_outputs[789] = (inputs[113]) | (inputs[149]);
    assign layer0_outputs[790] = (inputs[610]) ^ (inputs[24]);
    assign layer0_outputs[791] = (inputs[80]) | (inputs[747]);
    assign layer0_outputs[792] = ~((inputs[549]) & (inputs[223]));
    assign layer0_outputs[793] = (inputs[667]) & ~(inputs[1002]);
    assign layer0_outputs[794] = (inputs[114]) & ~(inputs[379]);
    assign layer0_outputs[795] = ~((inputs[368]) & (inputs[493]));
    assign layer0_outputs[796] = ~(inputs[587]) | (inputs[317]);
    assign layer0_outputs[797] = inputs[802];
    assign layer0_outputs[798] = ~(inputs[222]);
    assign layer0_outputs[799] = ~(inputs[1000]);
    assign layer0_outputs[800] = ~(inputs[127]);
    assign layer0_outputs[801] = ~(inputs[932]) | (inputs[360]);
    assign layer0_outputs[802] = (inputs[442]) & (inputs[837]);
    assign layer0_outputs[803] = inputs[847];
    assign layer0_outputs[804] = ~((inputs[543]) ^ (inputs[404]));
    assign layer0_outputs[805] = ~((inputs[891]) ^ (inputs[706]));
    assign layer0_outputs[806] = (inputs[83]) & ~(inputs[196]);
    assign layer0_outputs[807] = ~(inputs[185]);
    assign layer0_outputs[808] = (inputs[924]) ^ (inputs[562]);
    assign layer0_outputs[809] = ~(inputs[667]);
    assign layer0_outputs[810] = (inputs[533]) & ~(inputs[850]);
    assign layer0_outputs[811] = (inputs[45]) & (inputs[1003]);
    assign layer0_outputs[812] = inputs[719];
    assign layer0_outputs[813] = (inputs[531]) & ~(inputs[575]);
    assign layer0_outputs[814] = (inputs[903]) & ~(inputs[215]);
    assign layer0_outputs[815] = (inputs[358]) ^ (inputs[857]);
    assign layer0_outputs[816] = (inputs[134]) ^ (inputs[23]);
    assign layer0_outputs[817] = ~(inputs[729]) | (inputs[917]);
    assign layer0_outputs[818] = 1'b0;
    assign layer0_outputs[819] = inputs[829];
    assign layer0_outputs[820] = ~(inputs[799]) | (inputs[1015]);
    assign layer0_outputs[821] = (inputs[902]) ^ (inputs[389]);
    assign layer0_outputs[822] = (inputs[669]) | (inputs[784]);
    assign layer0_outputs[823] = (inputs[284]) | (inputs[589]);
    assign layer0_outputs[824] = ~((inputs[99]) | (inputs[134]));
    assign layer0_outputs[825] = ~((inputs[2]) ^ (inputs[155]));
    assign layer0_outputs[826] = (inputs[761]) ^ (inputs[827]);
    assign layer0_outputs[827] = (inputs[319]) | (inputs[617]);
    assign layer0_outputs[828] = ~(inputs[316]);
    assign layer0_outputs[829] = (inputs[111]) | (inputs[793]);
    assign layer0_outputs[830] = (inputs[134]) & (inputs[816]);
    assign layer0_outputs[831] = inputs[583];
    assign layer0_outputs[832] = (inputs[332]) ^ (inputs[835]);
    assign layer0_outputs[833] = inputs[2];
    assign layer0_outputs[834] = inputs[975];
    assign layer0_outputs[835] = ~(inputs[631]);
    assign layer0_outputs[836] = (inputs[797]) | (inputs[158]);
    assign layer0_outputs[837] = (inputs[551]) | (inputs[583]);
    assign layer0_outputs[838] = (inputs[990]) & ~(inputs[801]);
    assign layer0_outputs[839] = ~(inputs[622]);
    assign layer0_outputs[840] = ~(inputs[900]) | (inputs[156]);
    assign layer0_outputs[841] = ~((inputs[1021]) | (inputs[996]));
    assign layer0_outputs[842] = ~(inputs[859]);
    assign layer0_outputs[843] = ~(inputs[377]) | (inputs[453]);
    assign layer0_outputs[844] = 1'b0;
    assign layer0_outputs[845] = (inputs[33]) ^ (inputs[9]);
    assign layer0_outputs[846] = ~(inputs[495]);
    assign layer0_outputs[847] = (inputs[107]) & ~(inputs[1023]);
    assign layer0_outputs[848] = (inputs[509]) & ~(inputs[503]);
    assign layer0_outputs[849] = inputs[945];
    assign layer0_outputs[850] = (inputs[494]) | (inputs[899]);
    assign layer0_outputs[851] = (inputs[468]) | (inputs[27]);
    assign layer0_outputs[852] = (inputs[755]) ^ (inputs[10]);
    assign layer0_outputs[853] = (inputs[521]) & ~(inputs[805]);
    assign layer0_outputs[854] = (inputs[541]) & (inputs[899]);
    assign layer0_outputs[855] = ~(inputs[536]);
    assign layer0_outputs[856] = (inputs[635]) & (inputs[184]);
    assign layer0_outputs[857] = ~((inputs[749]) ^ (inputs[774]));
    assign layer0_outputs[858] = ~(inputs[704]);
    assign layer0_outputs[859] = 1'b1;
    assign layer0_outputs[860] = (inputs[892]) & (inputs[903]);
    assign layer0_outputs[861] = (inputs[1020]) ^ (inputs[473]);
    assign layer0_outputs[862] = ~(inputs[424]) | (inputs[37]);
    assign layer0_outputs[863] = ~((inputs[11]) ^ (inputs[56]));
    assign layer0_outputs[864] = ~(inputs[683]) | (inputs[339]);
    assign layer0_outputs[865] = (inputs[941]) & ~(inputs[538]);
    assign layer0_outputs[866] = 1'b0;
    assign layer0_outputs[867] = (inputs[852]) | (inputs[661]);
    assign layer0_outputs[868] = 1'b1;
    assign layer0_outputs[869] = ~((inputs[398]) & (inputs[193]));
    assign layer0_outputs[870] = inputs[200];
    assign layer0_outputs[871] = 1'b1;
    assign layer0_outputs[872] = inputs[586];
    assign layer0_outputs[873] = 1'b0;
    assign layer0_outputs[874] = ~(inputs[762]) | (inputs[892]);
    assign layer0_outputs[875] = (inputs[330]) & ~(inputs[145]);
    assign layer0_outputs[876] = ~((inputs[593]) | (inputs[355]));
    assign layer0_outputs[877] = inputs[318];
    assign layer0_outputs[878] = inputs[701];
    assign layer0_outputs[879] = ~(inputs[600]) | (inputs[997]);
    assign layer0_outputs[880] = (inputs[631]) ^ (inputs[1022]);
    assign layer0_outputs[881] = inputs[409];
    assign layer0_outputs[882] = ~(inputs[290]);
    assign layer0_outputs[883] = inputs[906];
    assign layer0_outputs[884] = ~((inputs[924]) & (inputs[854]));
    assign layer0_outputs[885] = (inputs[229]) & ~(inputs[261]);
    assign layer0_outputs[886] = (inputs[270]) | (inputs[443]);
    assign layer0_outputs[887] = ~(inputs[235]);
    assign layer0_outputs[888] = ~(inputs[812]);
    assign layer0_outputs[889] = (inputs[61]) & (inputs[670]);
    assign layer0_outputs[890] = (inputs[892]) & ~(inputs[98]);
    assign layer0_outputs[891] = ~((inputs[224]) | (inputs[348]));
    assign layer0_outputs[892] = ~((inputs[10]) & (inputs[119]));
    assign layer0_outputs[893] = ~((inputs[997]) | (inputs[538]));
    assign layer0_outputs[894] = ~(inputs[248]);
    assign layer0_outputs[895] = ~(inputs[762]) | (inputs[439]);
    assign layer0_outputs[896] = 1'b1;
    assign layer0_outputs[897] = 1'b0;
    assign layer0_outputs[898] = (inputs[73]) | (inputs[177]);
    assign layer0_outputs[899] = 1'b1;
    assign layer0_outputs[900] = (inputs[433]) & ~(inputs[188]);
    assign layer0_outputs[901] = (inputs[922]) ^ (inputs[380]);
    assign layer0_outputs[902] = ~((inputs[218]) | (inputs[332]));
    assign layer0_outputs[903] = 1'b1;
    assign layer0_outputs[904] = ~((inputs[642]) ^ (inputs[399]));
    assign layer0_outputs[905] = ~((inputs[474]) | (inputs[757]));
    assign layer0_outputs[906] = inputs[178];
    assign layer0_outputs[907] = (inputs[534]) | (inputs[81]);
    assign layer0_outputs[908] = (inputs[971]) & ~(inputs[35]);
    assign layer0_outputs[909] = inputs[610];
    assign layer0_outputs[910] = ~(inputs[989]);
    assign layer0_outputs[911] = ~((inputs[1017]) ^ (inputs[648]));
    assign layer0_outputs[912] = ~((inputs[625]) & (inputs[228]));
    assign layer0_outputs[913] = inputs[44];
    assign layer0_outputs[914] = ~((inputs[467]) | (inputs[885]));
    assign layer0_outputs[915] = ~((inputs[850]) | (inputs[245]));
    assign layer0_outputs[916] = (inputs[869]) ^ (inputs[69]);
    assign layer0_outputs[917] = 1'b0;
    assign layer0_outputs[918] = (inputs[142]) & ~(inputs[219]);
    assign layer0_outputs[919] = (inputs[907]) & (inputs[981]);
    assign layer0_outputs[920] = ~(inputs[846]) | (inputs[445]);
    assign layer0_outputs[921] = 1'b0;
    assign layer0_outputs[922] = ~((inputs[329]) | (inputs[193]));
    assign layer0_outputs[923] = (inputs[265]) & ~(inputs[896]);
    assign layer0_outputs[924] = ~(inputs[162]);
    assign layer0_outputs[925] = (inputs[53]) & ~(inputs[2]);
    assign layer0_outputs[926] = ~(inputs[616]) | (inputs[504]);
    assign layer0_outputs[927] = (inputs[33]) & ~(inputs[727]);
    assign layer0_outputs[928] = (inputs[943]) ^ (inputs[291]);
    assign layer0_outputs[929] = 1'b1;
    assign layer0_outputs[930] = (inputs[233]) & ~(inputs[392]);
    assign layer0_outputs[931] = ~(inputs[461]) | (inputs[982]);
    assign layer0_outputs[932] = 1'b1;
    assign layer0_outputs[933] = ~(inputs[142]);
    assign layer0_outputs[934] = ~((inputs[1004]) ^ (inputs[225]));
    assign layer0_outputs[935] = ~((inputs[175]) | (inputs[643]));
    assign layer0_outputs[936] = ~((inputs[226]) | (inputs[355]));
    assign layer0_outputs[937] = (inputs[896]) & ~(inputs[293]);
    assign layer0_outputs[938] = 1'b1;
    assign layer0_outputs[939] = inputs[569];
    assign layer0_outputs[940] = ~(inputs[496]) | (inputs[53]);
    assign layer0_outputs[941] = 1'b1;
    assign layer0_outputs[942] = ~(inputs[694]);
    assign layer0_outputs[943] = ~(inputs[989]);
    assign layer0_outputs[944] = ~((inputs[930]) & (inputs[244]));
    assign layer0_outputs[945] = 1'b1;
    assign layer0_outputs[946] = inputs[714];
    assign layer0_outputs[947] = ~(inputs[969]) | (inputs[677]);
    assign layer0_outputs[948] = ~(inputs[601]) | (inputs[920]);
    assign layer0_outputs[949] = ~(inputs[657]);
    assign layer0_outputs[950] = (inputs[2]) ^ (inputs[245]);
    assign layer0_outputs[951] = ~(inputs[677]);
    assign layer0_outputs[952] = ~(inputs[304]) | (inputs[744]);
    assign layer0_outputs[953] = ~((inputs[899]) ^ (inputs[483]));
    assign layer0_outputs[954] = inputs[490];
    assign layer0_outputs[955] = (inputs[335]) & ~(inputs[756]);
    assign layer0_outputs[956] = inputs[848];
    assign layer0_outputs[957] = 1'b0;
    assign layer0_outputs[958] = (inputs[869]) & ~(inputs[207]);
    assign layer0_outputs[959] = ~(inputs[443]) | (inputs[1001]);
    assign layer0_outputs[960] = 1'b0;
    assign layer0_outputs[961] = ~(inputs[257]) | (inputs[922]);
    assign layer0_outputs[962] = ~((inputs[386]) & (inputs[933]));
    assign layer0_outputs[963] = (inputs[623]) | (inputs[911]);
    assign layer0_outputs[964] = inputs[274];
    assign layer0_outputs[965] = inputs[58];
    assign layer0_outputs[966] = ~((inputs[140]) & (inputs[260]));
    assign layer0_outputs[967] = inputs[277];
    assign layer0_outputs[968] = (inputs[114]) ^ (inputs[528]);
    assign layer0_outputs[969] = ~(inputs[512]) | (inputs[693]);
    assign layer0_outputs[970] = ~(inputs[668]) | (inputs[682]);
    assign layer0_outputs[971] = ~(inputs[94]);
    assign layer0_outputs[972] = inputs[124];
    assign layer0_outputs[973] = ~((inputs[856]) & (inputs[976]));
    assign layer0_outputs[974] = ~(inputs[160]) | (inputs[809]);
    assign layer0_outputs[975] = 1'b0;
    assign layer0_outputs[976] = ~(inputs[394]) | (inputs[492]);
    assign layer0_outputs[977] = (inputs[900]) & (inputs[66]);
    assign layer0_outputs[978] = ~((inputs[839]) | (inputs[169]));
    assign layer0_outputs[979] = 1'b1;
    assign layer0_outputs[980] = (inputs[104]) ^ (inputs[496]);
    assign layer0_outputs[981] = (inputs[735]) & ~(inputs[85]);
    assign layer0_outputs[982] = (inputs[162]) | (inputs[1005]);
    assign layer0_outputs[983] = ~((inputs[434]) & (inputs[927]));
    assign layer0_outputs[984] = inputs[429];
    assign layer0_outputs[985] = ~((inputs[236]) ^ (inputs[317]));
    assign layer0_outputs[986] = (inputs[457]) | (inputs[949]);
    assign layer0_outputs[987] = (inputs[206]) ^ (inputs[786]);
    assign layer0_outputs[988] = (inputs[868]) | (inputs[875]);
    assign layer0_outputs[989] = (inputs[424]) | (inputs[47]);
    assign layer0_outputs[990] = ~((inputs[963]) & (inputs[952]));
    assign layer0_outputs[991] = ~((inputs[100]) | (inputs[5]));
    assign layer0_outputs[992] = 1'b0;
    assign layer0_outputs[993] = ~((inputs[69]) ^ (inputs[931]));
    assign layer0_outputs[994] = (inputs[732]) & ~(inputs[592]);
    assign layer0_outputs[995] = ~(inputs[520]) | (inputs[149]);
    assign layer0_outputs[996] = ~(inputs[913]);
    assign layer0_outputs[997] = (inputs[651]) | (inputs[786]);
    assign layer0_outputs[998] = (inputs[498]) & ~(inputs[722]);
    assign layer0_outputs[999] = ~((inputs[441]) ^ (inputs[155]));
    assign layer0_outputs[1000] = inputs[617];
    assign layer0_outputs[1001] = (inputs[464]) & (inputs[949]);
    assign layer0_outputs[1002] = (inputs[617]) | (inputs[1005]);
    assign layer0_outputs[1003] = (inputs[1023]) & ~(inputs[327]);
    assign layer0_outputs[1004] = ~((inputs[297]) | (inputs[564]));
    assign layer0_outputs[1005] = inputs[972];
    assign layer0_outputs[1006] = (inputs[558]) | (inputs[58]);
    assign layer0_outputs[1007] = (inputs[156]) & (inputs[919]);
    assign layer0_outputs[1008] = (inputs[153]) ^ (inputs[588]);
    assign layer0_outputs[1009] = (inputs[300]) | (inputs[664]);
    assign layer0_outputs[1010] = 1'b1;
    assign layer0_outputs[1011] = ~((inputs[992]) ^ (inputs[328]));
    assign layer0_outputs[1012] = ~(inputs[529]);
    assign layer0_outputs[1013] = ~(inputs[809]) | (inputs[598]);
    assign layer0_outputs[1014] = ~(inputs[783]) | (inputs[833]);
    assign layer0_outputs[1015] = (inputs[450]) ^ (inputs[146]);
    assign layer0_outputs[1016] = (inputs[914]) ^ (inputs[856]);
    assign layer0_outputs[1017] = (inputs[956]) ^ (inputs[21]);
    assign layer0_outputs[1018] = (inputs[883]) ^ (inputs[26]);
    assign layer0_outputs[1019] = (inputs[643]) ^ (inputs[425]);
    assign layer0_outputs[1020] = ~((inputs[996]) | (inputs[673]));
    assign layer0_outputs[1021] = inputs[370];
    assign layer0_outputs[1022] = ~(inputs[315]) | (inputs[534]);
    assign layer0_outputs[1023] = ~((inputs[582]) & (inputs[397]));
    assign layer0_outputs[1024] = ~(inputs[743]);
    assign layer0_outputs[1025] = (inputs[208]) | (inputs[148]);
    assign layer0_outputs[1026] = (inputs[78]) ^ (inputs[118]);
    assign layer0_outputs[1027] = (inputs[250]) | (inputs[281]);
    assign layer0_outputs[1028] = (inputs[194]) & ~(inputs[291]);
    assign layer0_outputs[1029] = ~(inputs[203]);
    assign layer0_outputs[1030] = (inputs[817]) | (inputs[38]);
    assign layer0_outputs[1031] = 1'b1;
    assign layer0_outputs[1032] = 1'b0;
    assign layer0_outputs[1033] = inputs[209];
    assign layer0_outputs[1034] = inputs[748];
    assign layer0_outputs[1035] = (inputs[938]) | (inputs[894]);
    assign layer0_outputs[1036] = ~(inputs[905]);
    assign layer0_outputs[1037] = (inputs[31]) ^ (inputs[455]);
    assign layer0_outputs[1038] = (inputs[384]) & (inputs[821]);
    assign layer0_outputs[1039] = (inputs[266]) & (inputs[457]);
    assign layer0_outputs[1040] = (inputs[341]) | (inputs[677]);
    assign layer0_outputs[1041] = (inputs[158]) ^ (inputs[521]);
    assign layer0_outputs[1042] = (inputs[813]) | (inputs[245]);
    assign layer0_outputs[1043] = ~((inputs[305]) ^ (inputs[157]));
    assign layer0_outputs[1044] = 1'b1;
    assign layer0_outputs[1045] = (inputs[319]) ^ (inputs[77]);
    assign layer0_outputs[1046] = ~(inputs[825]) | (inputs[229]);
    assign layer0_outputs[1047] = inputs[681];
    assign layer0_outputs[1048] = (inputs[735]) & ~(inputs[786]);
    assign layer0_outputs[1049] = ~((inputs[726]) & (inputs[800]));
    assign layer0_outputs[1050] = (inputs[845]) | (inputs[1012]);
    assign layer0_outputs[1051] = inputs[738];
    assign layer0_outputs[1052] = ~(inputs[489]);
    assign layer0_outputs[1053] = inputs[576];
    assign layer0_outputs[1054] = inputs[707];
    assign layer0_outputs[1055] = ~(inputs[587]);
    assign layer0_outputs[1056] = ~(inputs[86]) | (inputs[952]);
    assign layer0_outputs[1057] = ~(inputs[453]);
    assign layer0_outputs[1058] = 1'b1;
    assign layer0_outputs[1059] = ~(inputs[662]) | (inputs[14]);
    assign layer0_outputs[1060] = inputs[362];
    assign layer0_outputs[1061] = 1'b0;
    assign layer0_outputs[1062] = ~(inputs[125]);
    assign layer0_outputs[1063] = (inputs[481]) & (inputs[507]);
    assign layer0_outputs[1064] = ~(inputs[98]);
    assign layer0_outputs[1065] = 1'b0;
    assign layer0_outputs[1066] = ~((inputs[672]) & (inputs[981]));
    assign layer0_outputs[1067] = ~((inputs[910]) & (inputs[113]));
    assign layer0_outputs[1068] = ~((inputs[93]) | (inputs[589]));
    assign layer0_outputs[1069] = 1'b1;
    assign layer0_outputs[1070] = (inputs[817]) & ~(inputs[353]);
    assign layer0_outputs[1071] = (inputs[200]) & ~(inputs[86]);
    assign layer0_outputs[1072] = (inputs[8]) | (inputs[857]);
    assign layer0_outputs[1073] = inputs[470];
    assign layer0_outputs[1074] = (inputs[943]) ^ (inputs[935]);
    assign layer0_outputs[1075] = 1'b1;
    assign layer0_outputs[1076] = inputs[743];
    assign layer0_outputs[1077] = ~((inputs[214]) & (inputs[286]));
    assign layer0_outputs[1078] = ~((inputs[489]) | (inputs[415]));
    assign layer0_outputs[1079] = inputs[381];
    assign layer0_outputs[1080] = ~((inputs[955]) | (inputs[1]));
    assign layer0_outputs[1081] = (inputs[456]) | (inputs[978]);
    assign layer0_outputs[1082] = inputs[12];
    assign layer0_outputs[1083] = (inputs[264]) ^ (inputs[347]);
    assign layer0_outputs[1084] = ~(inputs[789]) | (inputs[889]);
    assign layer0_outputs[1085] = (inputs[139]) | (inputs[946]);
    assign layer0_outputs[1086] = (inputs[795]) | (inputs[455]);
    assign layer0_outputs[1087] = ~((inputs[798]) ^ (inputs[252]));
    assign layer0_outputs[1088] = ~((inputs[778]) | (inputs[790]));
    assign layer0_outputs[1089] = ~(inputs[32]);
    assign layer0_outputs[1090] = inputs[920];
    assign layer0_outputs[1091] = ~((inputs[526]) | (inputs[234]));
    assign layer0_outputs[1092] = ~(inputs[726]) | (inputs[992]);
    assign layer0_outputs[1093] = (inputs[720]) & (inputs[884]);
    assign layer0_outputs[1094] = 1'b1;
    assign layer0_outputs[1095] = inputs[907];
    assign layer0_outputs[1096] = ~((inputs[991]) & (inputs[635]));
    assign layer0_outputs[1097] = ~((inputs[475]) | (inputs[851]));
    assign layer0_outputs[1098] = inputs[747];
    assign layer0_outputs[1099] = (inputs[1018]) & ~(inputs[440]);
    assign layer0_outputs[1100] = (inputs[52]) & ~(inputs[328]);
    assign layer0_outputs[1101] = (inputs[249]) & ~(inputs[1014]);
    assign layer0_outputs[1102] = ~(inputs[556]);
    assign layer0_outputs[1103] = ~(inputs[12]) | (inputs[736]);
    assign layer0_outputs[1104] = 1'b1;
    assign layer0_outputs[1105] = ~((inputs[94]) | (inputs[234]));
    assign layer0_outputs[1106] = (inputs[555]) & (inputs[107]);
    assign layer0_outputs[1107] = (inputs[393]) & ~(inputs[498]);
    assign layer0_outputs[1108] = (inputs[523]) & ~(inputs[607]);
    assign layer0_outputs[1109] = ~(inputs[23]) | (inputs[217]);
    assign layer0_outputs[1110] = (inputs[717]) | (inputs[250]);
    assign layer0_outputs[1111] = ~((inputs[862]) | (inputs[5]));
    assign layer0_outputs[1112] = inputs[428];
    assign layer0_outputs[1113] = ~(inputs[273]) | (inputs[243]);
    assign layer0_outputs[1114] = inputs[40];
    assign layer0_outputs[1115] = ~((inputs[550]) | (inputs[55]));
    assign layer0_outputs[1116] = (inputs[829]) & ~(inputs[551]);
    assign layer0_outputs[1117] = 1'b0;
    assign layer0_outputs[1118] = (inputs[602]) & (inputs[769]);
    assign layer0_outputs[1119] = ~(inputs[308]) | (inputs[61]);
    assign layer0_outputs[1120] = inputs[378];
    assign layer0_outputs[1121] = ~(inputs[304]) | (inputs[685]);
    assign layer0_outputs[1122] = ~((inputs[39]) & (inputs[812]));
    assign layer0_outputs[1123] = (inputs[206]) | (inputs[920]);
    assign layer0_outputs[1124] = (inputs[944]) | (inputs[85]);
    assign layer0_outputs[1125] = inputs[713];
    assign layer0_outputs[1126] = 1'b0;
    assign layer0_outputs[1127] = inputs[399];
    assign layer0_outputs[1128] = ~(inputs[605]) | (inputs[934]);
    assign layer0_outputs[1129] = ~((inputs[234]) & (inputs[232]));
    assign layer0_outputs[1130] = ~(inputs[414]);
    assign layer0_outputs[1131] = (inputs[143]) ^ (inputs[109]);
    assign layer0_outputs[1132] = ~(inputs[213]);
    assign layer0_outputs[1133] = 1'b0;
    assign layer0_outputs[1134] = (inputs[985]) ^ (inputs[506]);
    assign layer0_outputs[1135] = ~((inputs[715]) | (inputs[103]));
    assign layer0_outputs[1136] = ~(inputs[768]);
    assign layer0_outputs[1137] = (inputs[123]) & (inputs[293]);
    assign layer0_outputs[1138] = ~(inputs[980]);
    assign layer0_outputs[1139] = ~(inputs[408]);
    assign layer0_outputs[1140] = (inputs[596]) & (inputs[860]);
    assign layer0_outputs[1141] = ~(inputs[597]);
    assign layer0_outputs[1142] = 1'b1;
    assign layer0_outputs[1143] = inputs[686];
    assign layer0_outputs[1144] = ~(inputs[753]);
    assign layer0_outputs[1145] = (inputs[473]) & ~(inputs[60]);
    assign layer0_outputs[1146] = inputs[218];
    assign layer0_outputs[1147] = ~(inputs[222]);
    assign layer0_outputs[1148] = ~(inputs[572]);
    assign layer0_outputs[1149] = ~((inputs[864]) | (inputs[581]));
    assign layer0_outputs[1150] = (inputs[722]) & (inputs[1021]);
    assign layer0_outputs[1151] = ~(inputs[373]);
    assign layer0_outputs[1152] = ~(inputs[218]) | (inputs[446]);
    assign layer0_outputs[1153] = (inputs[734]) ^ (inputs[986]);
    assign layer0_outputs[1154] = inputs[761];
    assign layer0_outputs[1155] = (inputs[951]) & ~(inputs[470]);
    assign layer0_outputs[1156] = (inputs[822]) ^ (inputs[895]);
    assign layer0_outputs[1157] = 1'b1;
    assign layer0_outputs[1158] = (inputs[124]) | (inputs[117]);
    assign layer0_outputs[1159] = 1'b0;
    assign layer0_outputs[1160] = inputs[560];
    assign layer0_outputs[1161] = (inputs[516]) & (inputs[890]);
    assign layer0_outputs[1162] = 1'b1;
    assign layer0_outputs[1163] = ~(inputs[146]);
    assign layer0_outputs[1164] = (inputs[177]) & ~(inputs[841]);
    assign layer0_outputs[1165] = 1'b0;
    assign layer0_outputs[1166] = (inputs[6]) & ~(inputs[565]);
    assign layer0_outputs[1167] = (inputs[811]) & (inputs[31]);
    assign layer0_outputs[1168] = ~(inputs[795]);
    assign layer0_outputs[1169] = ~((inputs[223]) ^ (inputs[373]));
    assign layer0_outputs[1170] = ~((inputs[982]) & (inputs[187]));
    assign layer0_outputs[1171] = inputs[842];
    assign layer0_outputs[1172] = 1'b0;
    assign layer0_outputs[1173] = (inputs[626]) & (inputs[646]);
    assign layer0_outputs[1174] = (inputs[695]) & ~(inputs[361]);
    assign layer0_outputs[1175] = 1'b0;
    assign layer0_outputs[1176] = 1'b0;
    assign layer0_outputs[1177] = (inputs[663]) | (inputs[648]);
    assign layer0_outputs[1178] = ~(inputs[683]) | (inputs[835]);
    assign layer0_outputs[1179] = inputs[465];
    assign layer0_outputs[1180] = inputs[651];
    assign layer0_outputs[1181] = (inputs[295]) ^ (inputs[106]);
    assign layer0_outputs[1182] = ~((inputs[652]) | (inputs[373]));
    assign layer0_outputs[1183] = ~((inputs[237]) | (inputs[511]));
    assign layer0_outputs[1184] = 1'b0;
    assign layer0_outputs[1185] = ~(inputs[152]);
    assign layer0_outputs[1186] = (inputs[764]) | (inputs[778]);
    assign layer0_outputs[1187] = 1'b0;
    assign layer0_outputs[1188] = (inputs[78]) | (inputs[445]);
    assign layer0_outputs[1189] = 1'b0;
    assign layer0_outputs[1190] = ~(inputs[445]);
    assign layer0_outputs[1191] = (inputs[974]) & (inputs[23]);
    assign layer0_outputs[1192] = 1'b1;
    assign layer0_outputs[1193] = (inputs[596]) & ~(inputs[371]);
    assign layer0_outputs[1194] = ~((inputs[215]) ^ (inputs[821]));
    assign layer0_outputs[1195] = (inputs[744]) & ~(inputs[64]);
    assign layer0_outputs[1196] = 1'b0;
    assign layer0_outputs[1197] = (inputs[172]) & ~(inputs[550]);
    assign layer0_outputs[1198] = inputs[0];
    assign layer0_outputs[1199] = (inputs[110]) & ~(inputs[916]);
    assign layer0_outputs[1200] = 1'b0;
    assign layer0_outputs[1201] = (inputs[592]) & ~(inputs[425]);
    assign layer0_outputs[1202] = ~(inputs[658]) | (inputs[289]);
    assign layer0_outputs[1203] = ~((inputs[96]) & (inputs[276]));
    assign layer0_outputs[1204] = (inputs[684]) & ~(inputs[192]);
    assign layer0_outputs[1205] = 1'b1;
    assign layer0_outputs[1206] = ~(inputs[160]);
    assign layer0_outputs[1207] = ~(inputs[544]);
    assign layer0_outputs[1208] = inputs[1017];
    assign layer0_outputs[1209] = (inputs[1013]) & ~(inputs[735]);
    assign layer0_outputs[1210] = (inputs[933]) ^ (inputs[508]);
    assign layer0_outputs[1211] = (inputs[909]) & ~(inputs[129]);
    assign layer0_outputs[1212] = ~((inputs[169]) | (inputs[843]));
    assign layer0_outputs[1213] = ~(inputs[760]) | (inputs[819]);
    assign layer0_outputs[1214] = ~(inputs[168]);
    assign layer0_outputs[1215] = ~((inputs[849]) | (inputs[655]));
    assign layer0_outputs[1216] = (inputs[934]) ^ (inputs[210]);
    assign layer0_outputs[1217] = inputs[723];
    assign layer0_outputs[1218] = (inputs[739]) & (inputs[350]);
    assign layer0_outputs[1219] = (inputs[828]) & (inputs[465]);
    assign layer0_outputs[1220] = ~(inputs[836]);
    assign layer0_outputs[1221] = ~(inputs[618]);
    assign layer0_outputs[1222] = (inputs[751]) | (inputs[430]);
    assign layer0_outputs[1223] = ~(inputs[164]) | (inputs[488]);
    assign layer0_outputs[1224] = ~((inputs[562]) ^ (inputs[857]));
    assign layer0_outputs[1225] = (inputs[334]) | (inputs[331]);
    assign layer0_outputs[1226] = (inputs[217]) ^ (inputs[45]);
    assign layer0_outputs[1227] = (inputs[520]) & ~(inputs[384]);
    assign layer0_outputs[1228] = (inputs[944]) | (inputs[206]);
    assign layer0_outputs[1229] = (inputs[607]) | (inputs[463]);
    assign layer0_outputs[1230] = 1'b0;
    assign layer0_outputs[1231] = (inputs[301]) | (inputs[278]);
    assign layer0_outputs[1232] = ~((inputs[904]) ^ (inputs[404]));
    assign layer0_outputs[1233] = (inputs[497]) & ~(inputs[710]);
    assign layer0_outputs[1234] = 1'b0;
    assign layer0_outputs[1235] = ~((inputs[748]) | (inputs[849]));
    assign layer0_outputs[1236] = (inputs[409]) | (inputs[687]);
    assign layer0_outputs[1237] = 1'b0;
    assign layer0_outputs[1238] = (inputs[411]) ^ (inputs[337]);
    assign layer0_outputs[1239] = 1'b0;
    assign layer0_outputs[1240] = ~((inputs[259]) ^ (inputs[574]));
    assign layer0_outputs[1241] = 1'b1;
    assign layer0_outputs[1242] = (inputs[500]) & ~(inputs[602]);
    assign layer0_outputs[1243] = inputs[66];
    assign layer0_outputs[1244] = ~(inputs[511]);
    assign layer0_outputs[1245] = ~(inputs[800]) | (inputs[112]);
    assign layer0_outputs[1246] = ~(inputs[716]) | (inputs[174]);
    assign layer0_outputs[1247] = ~(inputs[433]);
    assign layer0_outputs[1248] = (inputs[171]) & (inputs[458]);
    assign layer0_outputs[1249] = (inputs[727]) | (inputs[776]);
    assign layer0_outputs[1250] = ~(inputs[355]);
    assign layer0_outputs[1251] = ~(inputs[953]) | (inputs[612]);
    assign layer0_outputs[1252] = ~(inputs[838]) | (inputs[963]);
    assign layer0_outputs[1253] = ~(inputs[188]);
    assign layer0_outputs[1254] = 1'b1;
    assign layer0_outputs[1255] = ~((inputs[795]) ^ (inputs[996]));
    assign layer0_outputs[1256] = ~(inputs[383]);
    assign layer0_outputs[1257] = (inputs[43]) ^ (inputs[483]);
    assign layer0_outputs[1258] = ~((inputs[801]) & (inputs[45]));
    assign layer0_outputs[1259] = inputs[775];
    assign layer0_outputs[1260] = inputs[101];
    assign layer0_outputs[1261] = ~((inputs[875]) ^ (inputs[154]));
    assign layer0_outputs[1262] = ~(inputs[72]) | (inputs[105]);
    assign layer0_outputs[1263] = (inputs[121]) & ~(inputs[999]);
    assign layer0_outputs[1264] = ~(inputs[609]);
    assign layer0_outputs[1265] = 1'b0;
    assign layer0_outputs[1266] = 1'b0;
    assign layer0_outputs[1267] = (inputs[313]) ^ (inputs[482]);
    assign layer0_outputs[1268] = ~((inputs[494]) ^ (inputs[172]));
    assign layer0_outputs[1269] = ~((inputs[115]) & (inputs[309]));
    assign layer0_outputs[1270] = 1'b0;
    assign layer0_outputs[1271] = inputs[731];
    assign layer0_outputs[1272] = (inputs[634]) & ~(inputs[630]);
    assign layer0_outputs[1273] = ~((inputs[273]) & (inputs[295]));
    assign layer0_outputs[1274] = ~(inputs[699]);
    assign layer0_outputs[1275] = 1'b0;
    assign layer0_outputs[1276] = (inputs[231]) & ~(inputs[510]);
    assign layer0_outputs[1277] = (inputs[766]) & ~(inputs[178]);
    assign layer0_outputs[1278] = ~(inputs[1003]) | (inputs[501]);
    assign layer0_outputs[1279] = (inputs[946]) & ~(inputs[941]);
    assign layer0_outputs[1280] = ~(inputs[583]);
    assign layer0_outputs[1281] = ~(inputs[63]);
    assign layer0_outputs[1282] = ~(inputs[84]);
    assign layer0_outputs[1283] = (inputs[282]) ^ (inputs[739]);
    assign layer0_outputs[1284] = ~(inputs[865]);
    assign layer0_outputs[1285] = inputs[753];
    assign layer0_outputs[1286] = ~(inputs[376]) | (inputs[593]);
    assign layer0_outputs[1287] = inputs[927];
    assign layer0_outputs[1288] = ~((inputs[868]) | (inputs[772]));
    assign layer0_outputs[1289] = ~(inputs[684]) | (inputs[485]);
    assign layer0_outputs[1290] = inputs[859];
    assign layer0_outputs[1291] = inputs[705];
    assign layer0_outputs[1292] = ~(inputs[4]) | (inputs[785]);
    assign layer0_outputs[1293] = (inputs[558]) & (inputs[766]);
    assign layer0_outputs[1294] = ~(inputs[126]) | (inputs[201]);
    assign layer0_outputs[1295] = (inputs[843]) | (inputs[711]);
    assign layer0_outputs[1296] = (inputs[743]) | (inputs[173]);
    assign layer0_outputs[1297] = inputs[947];
    assign layer0_outputs[1298] = (inputs[887]) | (inputs[733]);
    assign layer0_outputs[1299] = (inputs[506]) & ~(inputs[5]);
    assign layer0_outputs[1300] = (inputs[812]) ^ (inputs[6]);
    assign layer0_outputs[1301] = inputs[158];
    assign layer0_outputs[1302] = ~((inputs[764]) ^ (inputs[453]));
    assign layer0_outputs[1303] = inputs[176];
    assign layer0_outputs[1304] = inputs[50];
    assign layer0_outputs[1305] = (inputs[232]) & (inputs[568]);
    assign layer0_outputs[1306] = ~(inputs[1010]) | (inputs[705]);
    assign layer0_outputs[1307] = ~((inputs[990]) ^ (inputs[273]));
    assign layer0_outputs[1308] = inputs[463];
    assign layer0_outputs[1309] = ~(inputs[275]);
    assign layer0_outputs[1310] = 1'b0;
    assign layer0_outputs[1311] = 1'b1;
    assign layer0_outputs[1312] = (inputs[364]) & ~(inputs[950]);
    assign layer0_outputs[1313] = ~(inputs[271]) | (inputs[210]);
    assign layer0_outputs[1314] = ~(inputs[201]);
    assign layer0_outputs[1315] = ~(inputs[805]);
    assign layer0_outputs[1316] = inputs[152];
    assign layer0_outputs[1317] = ~((inputs[161]) & (inputs[435]));
    assign layer0_outputs[1318] = ~((inputs[605]) & (inputs[773]));
    assign layer0_outputs[1319] = (inputs[193]) & ~(inputs[149]);
    assign layer0_outputs[1320] = ~((inputs[508]) | (inputs[205]));
    assign layer0_outputs[1321] = (inputs[716]) & (inputs[51]);
    assign layer0_outputs[1322] = ~((inputs[917]) | (inputs[129]));
    assign layer0_outputs[1323] = (inputs[753]) & ~(inputs[536]);
    assign layer0_outputs[1324] = ~((inputs[518]) ^ (inputs[881]));
    assign layer0_outputs[1325] = (inputs[5]) ^ (inputs[608]);
    assign layer0_outputs[1326] = ~(inputs[373]) | (inputs[383]);
    assign layer0_outputs[1327] = ~(inputs[72]);
    assign layer0_outputs[1328] = ~(inputs[706]);
    assign layer0_outputs[1329] = ~(inputs[99]) | (inputs[19]);
    assign layer0_outputs[1330] = ~((inputs[25]) | (inputs[301]));
    assign layer0_outputs[1331] = 1'b1;
    assign layer0_outputs[1332] = (inputs[349]) & (inputs[1006]);
    assign layer0_outputs[1333] = ~((inputs[465]) ^ (inputs[82]));
    assign layer0_outputs[1334] = (inputs[831]) & ~(inputs[1014]);
    assign layer0_outputs[1335] = ~(inputs[463]) | (inputs[970]);
    assign layer0_outputs[1336] = ~((inputs[671]) ^ (inputs[1003]));
    assign layer0_outputs[1337] = (inputs[550]) & (inputs[644]);
    assign layer0_outputs[1338] = (inputs[703]) | (inputs[999]);
    assign layer0_outputs[1339] = inputs[146];
    assign layer0_outputs[1340] = inputs[516];
    assign layer0_outputs[1341] = (inputs[514]) ^ (inputs[701]);
    assign layer0_outputs[1342] = ~((inputs[454]) ^ (inputs[452]));
    assign layer0_outputs[1343] = (inputs[58]) & (inputs[14]);
    assign layer0_outputs[1344] = 1'b1;
    assign layer0_outputs[1345] = 1'b1;
    assign layer0_outputs[1346] = (inputs[489]) | (inputs[519]);
    assign layer0_outputs[1347] = ~(inputs[493]);
    assign layer0_outputs[1348] = 1'b1;
    assign layer0_outputs[1349] = ~((inputs[724]) ^ (inputs[883]));
    assign layer0_outputs[1350] = (inputs[598]) | (inputs[96]);
    assign layer0_outputs[1351] = ~((inputs[250]) & (inputs[1006]));
    assign layer0_outputs[1352] = (inputs[941]) | (inputs[446]);
    assign layer0_outputs[1353] = 1'b0;
    assign layer0_outputs[1354] = inputs[809];
    assign layer0_outputs[1355] = (inputs[429]) | (inputs[116]);
    assign layer0_outputs[1356] = inputs[437];
    assign layer0_outputs[1357] = (inputs[516]) ^ (inputs[735]);
    assign layer0_outputs[1358] = (inputs[138]) ^ (inputs[151]);
    assign layer0_outputs[1359] = (inputs[417]) ^ (inputs[84]);
    assign layer0_outputs[1360] = ~((inputs[165]) ^ (inputs[309]));
    assign layer0_outputs[1361] = (inputs[134]) | (inputs[807]);
    assign layer0_outputs[1362] = (inputs[587]) & ~(inputs[923]);
    assign layer0_outputs[1363] = (inputs[501]) | (inputs[254]);
    assign layer0_outputs[1364] = (inputs[102]) & (inputs[31]);
    assign layer0_outputs[1365] = 1'b0;
    assign layer0_outputs[1366] = (inputs[193]) | (inputs[433]);
    assign layer0_outputs[1367] = ~((inputs[32]) | (inputs[518]));
    assign layer0_outputs[1368] = ~(inputs[395]) | (inputs[695]);
    assign layer0_outputs[1369] = ~((inputs[183]) | (inputs[749]));
    assign layer0_outputs[1370] = 1'b0;
    assign layer0_outputs[1371] = ~((inputs[269]) ^ (inputs[189]));
    assign layer0_outputs[1372] = inputs[530];
    assign layer0_outputs[1373] = ~((inputs[0]) ^ (inputs[716]));
    assign layer0_outputs[1374] = (inputs[524]) & ~(inputs[1009]);
    assign layer0_outputs[1375] = ~((inputs[81]) ^ (inputs[137]));
    assign layer0_outputs[1376] = (inputs[151]) ^ (inputs[38]);
    assign layer0_outputs[1377] = ~(inputs[548]);
    assign layer0_outputs[1378] = ~((inputs[157]) ^ (inputs[614]));
    assign layer0_outputs[1379] = inputs[195];
    assign layer0_outputs[1380] = inputs[38];
    assign layer0_outputs[1381] = ~(inputs[759]);
    assign layer0_outputs[1382] = ~(inputs[997]);
    assign layer0_outputs[1383] = ~(inputs[975]) | (inputs[680]);
    assign layer0_outputs[1384] = (inputs[578]) | (inputs[159]);
    assign layer0_outputs[1385] = ~(inputs[220]) | (inputs[402]);
    assign layer0_outputs[1386] = (inputs[429]) | (inputs[114]);
    assign layer0_outputs[1387] = ~((inputs[273]) ^ (inputs[320]));
    assign layer0_outputs[1388] = (inputs[424]) & (inputs[869]);
    assign layer0_outputs[1389] = ~(inputs[275]);
    assign layer0_outputs[1390] = (inputs[234]) & (inputs[64]);
    assign layer0_outputs[1391] = ~((inputs[731]) ^ (inputs[890]));
    assign layer0_outputs[1392] = ~((inputs[863]) | (inputs[122]));
    assign layer0_outputs[1393] = (inputs[833]) ^ (inputs[892]);
    assign layer0_outputs[1394] = ~((inputs[843]) | (inputs[65]));
    assign layer0_outputs[1395] = inputs[344];
    assign layer0_outputs[1396] = (inputs[868]) ^ (inputs[80]);
    assign layer0_outputs[1397] = (inputs[126]) & ~(inputs[800]);
    assign layer0_outputs[1398] = ~((inputs[810]) ^ (inputs[973]));
    assign layer0_outputs[1399] = ~(inputs[34]);
    assign layer0_outputs[1400] = ~(inputs[285]);
    assign layer0_outputs[1401] = ~(inputs[880]);
    assign layer0_outputs[1402] = inputs[244];
    assign layer0_outputs[1403] = ~((inputs[127]) ^ (inputs[777]));
    assign layer0_outputs[1404] = (inputs[45]) | (inputs[570]);
    assign layer0_outputs[1405] = inputs[478];
    assign layer0_outputs[1406] = inputs[876];
    assign layer0_outputs[1407] = ~(inputs[599]) | (inputs[1018]);
    assign layer0_outputs[1408] = 1'b1;
    assign layer0_outputs[1409] = (inputs[44]) | (inputs[937]);
    assign layer0_outputs[1410] = ~(inputs[586]);
    assign layer0_outputs[1411] = ~(inputs[246]) | (inputs[940]);
    assign layer0_outputs[1412] = 1'b1;
    assign layer0_outputs[1413] = ~((inputs[741]) | (inputs[190]));
    assign layer0_outputs[1414] = (inputs[82]) & ~(inputs[627]);
    assign layer0_outputs[1415] = ~(inputs[960]);
    assign layer0_outputs[1416] = 1'b1;
    assign layer0_outputs[1417] = ~((inputs[101]) & (inputs[949]));
    assign layer0_outputs[1418] = inputs[995];
    assign layer0_outputs[1419] = 1'b0;
    assign layer0_outputs[1420] = (inputs[76]) | (inputs[838]);
    assign layer0_outputs[1421] = (inputs[96]) | (inputs[636]);
    assign layer0_outputs[1422] = (inputs[857]) & ~(inputs[708]);
    assign layer0_outputs[1423] = (inputs[977]) & ~(inputs[1007]);
    assign layer0_outputs[1424] = ~((inputs[685]) | (inputs[623]));
    assign layer0_outputs[1425] = (inputs[719]) ^ (inputs[705]);
    assign layer0_outputs[1426] = (inputs[860]) ^ (inputs[340]);
    assign layer0_outputs[1427] = 1'b1;
    assign layer0_outputs[1428] = (inputs[359]) & ~(inputs[1002]);
    assign layer0_outputs[1429] = ~((inputs[792]) | (inputs[788]));
    assign layer0_outputs[1430] = (inputs[919]) & ~(inputs[336]);
    assign layer0_outputs[1431] = (inputs[25]) & ~(inputs[353]);
    assign layer0_outputs[1432] = (inputs[304]) | (inputs[100]);
    assign layer0_outputs[1433] = (inputs[483]) & (inputs[622]);
    assign layer0_outputs[1434] = ~(inputs[75]) | (inputs[183]);
    assign layer0_outputs[1435] = ~(inputs[351]) | (inputs[39]);
    assign layer0_outputs[1436] = ~(inputs[202]);
    assign layer0_outputs[1437] = inputs[852];
    assign layer0_outputs[1438] = (inputs[810]) & ~(inputs[367]);
    assign layer0_outputs[1439] = (inputs[590]) & ~(inputs[706]);
    assign layer0_outputs[1440] = 1'b1;
    assign layer0_outputs[1441] = ~((inputs[929]) & (inputs[130]));
    assign layer0_outputs[1442] = inputs[604];
    assign layer0_outputs[1443] = ~((inputs[232]) & (inputs[446]));
    assign layer0_outputs[1444] = (inputs[497]) & ~(inputs[789]);
    assign layer0_outputs[1445] = ~((inputs[921]) ^ (inputs[513]));
    assign layer0_outputs[1446] = 1'b0;
    assign layer0_outputs[1447] = (inputs[663]) | (inputs[831]);
    assign layer0_outputs[1448] = inputs[553];
    assign layer0_outputs[1449] = ~(inputs[304]) | (inputs[738]);
    assign layer0_outputs[1450] = 1'b1;
    assign layer0_outputs[1451] = ~(inputs[1002]) | (inputs[173]);
    assign layer0_outputs[1452] = ~(inputs[264]) | (inputs[91]);
    assign layer0_outputs[1453] = (inputs[504]) & (inputs[423]);
    assign layer0_outputs[1454] = (inputs[611]) | (inputs[1013]);
    assign layer0_outputs[1455] = ~(inputs[463]) | (inputs[488]);
    assign layer0_outputs[1456] = (inputs[557]) | (inputs[212]);
    assign layer0_outputs[1457] = (inputs[950]) & ~(inputs[607]);
    assign layer0_outputs[1458] = (inputs[988]) & ~(inputs[162]);
    assign layer0_outputs[1459] = (inputs[418]) & (inputs[745]);
    assign layer0_outputs[1460] = 1'b0;
    assign layer0_outputs[1461] = (inputs[640]) ^ (inputs[18]);
    assign layer0_outputs[1462] = inputs[712];
    assign layer0_outputs[1463] = ~((inputs[377]) | (inputs[845]));
    assign layer0_outputs[1464] = inputs[461];
    assign layer0_outputs[1465] = ~(inputs[49]);
    assign layer0_outputs[1466] = ~((inputs[387]) & (inputs[25]));
    assign layer0_outputs[1467] = ~((inputs[375]) | (inputs[476]));
    assign layer0_outputs[1468] = inputs[204];
    assign layer0_outputs[1469] = ~(inputs[344]) | (inputs[357]);
    assign layer0_outputs[1470] = (inputs[526]) & (inputs[396]);
    assign layer0_outputs[1471] = ~(inputs[369]);
    assign layer0_outputs[1472] = 1'b0;
    assign layer0_outputs[1473] = (inputs[882]) & ~(inputs[616]);
    assign layer0_outputs[1474] = ~((inputs[541]) | (inputs[486]));
    assign layer0_outputs[1475] = (inputs[267]) & ~(inputs[322]);
    assign layer0_outputs[1476] = ~((inputs[251]) | (inputs[931]));
    assign layer0_outputs[1477] = ~(inputs[212]);
    assign layer0_outputs[1478] = ~((inputs[711]) | (inputs[730]));
    assign layer0_outputs[1479] = 1'b1;
    assign layer0_outputs[1480] = inputs[835];
    assign layer0_outputs[1481] = (inputs[68]) & (inputs[324]);
    assign layer0_outputs[1482] = ~(inputs[622]) | (inputs[14]);
    assign layer0_outputs[1483] = ~(inputs[880]);
    assign layer0_outputs[1484] = inputs[232];
    assign layer0_outputs[1485] = ~(inputs[392]);
    assign layer0_outputs[1486] = ~((inputs[595]) | (inputs[945]));
    assign layer0_outputs[1487] = inputs[22];
    assign layer0_outputs[1488] = ~(inputs[47]);
    assign layer0_outputs[1489] = 1'b1;
    assign layer0_outputs[1490] = ~(inputs[799]) | (inputs[756]);
    assign layer0_outputs[1491] = ~((inputs[891]) & (inputs[123]));
    assign layer0_outputs[1492] = ~(inputs[1006]);
    assign layer0_outputs[1493] = ~((inputs[861]) ^ (inputs[555]));
    assign layer0_outputs[1494] = ~(inputs[714]) | (inputs[229]);
    assign layer0_outputs[1495] = (inputs[755]) & ~(inputs[364]);
    assign layer0_outputs[1496] = ~(inputs[108]) | (inputs[514]);
    assign layer0_outputs[1497] = (inputs[259]) & ~(inputs[417]);
    assign layer0_outputs[1498] = (inputs[298]) & (inputs[239]);
    assign layer0_outputs[1499] = (inputs[71]) | (inputs[903]);
    assign layer0_outputs[1500] = 1'b0;
    assign layer0_outputs[1501] = (inputs[644]) & (inputs[263]);
    assign layer0_outputs[1502] = ~((inputs[570]) | (inputs[185]));
    assign layer0_outputs[1503] = ~(inputs[291]) | (inputs[345]);
    assign layer0_outputs[1504] = (inputs[47]) ^ (inputs[531]);
    assign layer0_outputs[1505] = (inputs[143]) & ~(inputs[867]);
    assign layer0_outputs[1506] = (inputs[376]) & ~(inputs[26]);
    assign layer0_outputs[1507] = (inputs[524]) & ~(inputs[224]);
    assign layer0_outputs[1508] = ~(inputs[452]) | (inputs[305]);
    assign layer0_outputs[1509] = ~((inputs[683]) | (inputs[731]));
    assign layer0_outputs[1510] = inputs[137];
    assign layer0_outputs[1511] = (inputs[246]) ^ (inputs[289]);
    assign layer0_outputs[1512] = (inputs[721]) | (inputs[84]);
    assign layer0_outputs[1513] = ~(inputs[942]);
    assign layer0_outputs[1514] = ~(inputs[759]);
    assign layer0_outputs[1515] = (inputs[129]) & ~(inputs[341]);
    assign layer0_outputs[1516] = ~(inputs[1004]);
    assign layer0_outputs[1517] = ~(inputs[351]);
    assign layer0_outputs[1518] = ~((inputs[174]) ^ (inputs[637]));
    assign layer0_outputs[1519] = 1'b1;
    assign layer0_outputs[1520] = 1'b1;
    assign layer0_outputs[1521] = ~((inputs[729]) | (inputs[217]));
    assign layer0_outputs[1522] = ~(inputs[442]) | (inputs[956]);
    assign layer0_outputs[1523] = ~(inputs[138]) | (inputs[283]);
    assign layer0_outputs[1524] = 1'b0;
    assign layer0_outputs[1525] = ~(inputs[552]) | (inputs[132]);
    assign layer0_outputs[1526] = (inputs[603]) & ~(inputs[384]);
    assign layer0_outputs[1527] = ~(inputs[329]);
    assign layer0_outputs[1528] = ~((inputs[533]) | (inputs[586]));
    assign layer0_outputs[1529] = inputs[340];
    assign layer0_outputs[1530] = ~((inputs[528]) | (inputs[864]));
    assign layer0_outputs[1531] = (inputs[395]) | (inputs[327]);
    assign layer0_outputs[1532] = (inputs[426]) & ~(inputs[838]);
    assign layer0_outputs[1533] = (inputs[129]) ^ (inputs[965]);
    assign layer0_outputs[1534] = ~(inputs[506]);
    assign layer0_outputs[1535] = ~(inputs[554]) | (inputs[100]);
    assign layer0_outputs[1536] = ~(inputs[459]);
    assign layer0_outputs[1537] = ~((inputs[297]) & (inputs[29]));
    assign layer0_outputs[1538] = ~(inputs[845]) | (inputs[970]);
    assign layer0_outputs[1539] = ~((inputs[106]) | (inputs[254]));
    assign layer0_outputs[1540] = ~(inputs[622]);
    assign layer0_outputs[1541] = ~(inputs[619]);
    assign layer0_outputs[1542] = inputs[43];
    assign layer0_outputs[1543] = (inputs[125]) | (inputs[58]);
    assign layer0_outputs[1544] = (inputs[342]) & ~(inputs[946]);
    assign layer0_outputs[1545] = ~(inputs[746]) | (inputs[352]);
    assign layer0_outputs[1546] = (inputs[730]) & (inputs[516]);
    assign layer0_outputs[1547] = (inputs[411]) | (inputs[95]);
    assign layer0_outputs[1548] = ~(inputs[522]) | (inputs[742]);
    assign layer0_outputs[1549] = (inputs[729]) | (inputs[294]);
    assign layer0_outputs[1550] = 1'b0;
    assign layer0_outputs[1551] = (inputs[547]) & ~(inputs[132]);
    assign layer0_outputs[1552] = (inputs[318]) | (inputs[834]);
    assign layer0_outputs[1553] = inputs[671];
    assign layer0_outputs[1554] = ~((inputs[996]) | (inputs[616]));
    assign layer0_outputs[1555] = ~((inputs[516]) | (inputs[233]));
    assign layer0_outputs[1556] = (inputs[443]) & ~(inputs[182]);
    assign layer0_outputs[1557] = (inputs[712]) & ~(inputs[915]);
    assign layer0_outputs[1558] = ~(inputs[57]);
    assign layer0_outputs[1559] = ~(inputs[832]);
    assign layer0_outputs[1560] = ~(inputs[20]) | (inputs[791]);
    assign layer0_outputs[1561] = ~((inputs[691]) | (inputs[570]));
    assign layer0_outputs[1562] = (inputs[907]) & ~(inputs[359]);
    assign layer0_outputs[1563] = ~((inputs[80]) | (inputs[170]));
    assign layer0_outputs[1564] = ~(inputs[67]);
    assign layer0_outputs[1565] = 1'b0;
    assign layer0_outputs[1566] = (inputs[861]) & (inputs[552]);
    assign layer0_outputs[1567] = (inputs[895]) | (inputs[254]);
    assign layer0_outputs[1568] = ~((inputs[124]) ^ (inputs[416]));
    assign layer0_outputs[1569] = inputs[1019];
    assign layer0_outputs[1570] = ~((inputs[71]) | (inputs[497]));
    assign layer0_outputs[1571] = ~((inputs[547]) & (inputs[479]));
    assign layer0_outputs[1572] = (inputs[864]) ^ (inputs[73]);
    assign layer0_outputs[1573] = ~(inputs[697]) | (inputs[611]);
    assign layer0_outputs[1574] = (inputs[780]) & ~(inputs[464]);
    assign layer0_outputs[1575] = (inputs[202]) & ~(inputs[42]);
    assign layer0_outputs[1576] = inputs[11];
    assign layer0_outputs[1577] = ~((inputs[480]) | (inputs[901]));
    assign layer0_outputs[1578] = (inputs[618]) ^ (inputs[909]);
    assign layer0_outputs[1579] = (inputs[437]) | (inputs[499]);
    assign layer0_outputs[1580] = ~(inputs[960]);
    assign layer0_outputs[1581] = ~((inputs[348]) | (inputs[703]));
    assign layer0_outputs[1582] = ~(inputs[818]);
    assign layer0_outputs[1583] = ~(inputs[24]) | (inputs[547]);
    assign layer0_outputs[1584] = ~((inputs[699]) & (inputs[630]));
    assign layer0_outputs[1585] = (inputs[482]) & ~(inputs[408]);
    assign layer0_outputs[1586] = ~((inputs[662]) | (inputs[54]));
    assign layer0_outputs[1587] = ~((inputs[250]) | (inputs[911]));
    assign layer0_outputs[1588] = ~((inputs[420]) & (inputs[676]));
    assign layer0_outputs[1589] = (inputs[267]) & ~(inputs[870]);
    assign layer0_outputs[1590] = inputs[750];
    assign layer0_outputs[1591] = (inputs[88]) & ~(inputs[594]);
    assign layer0_outputs[1592] = ~(inputs[21]) | (inputs[580]);
    assign layer0_outputs[1593] = (inputs[1012]) & (inputs[404]);
    assign layer0_outputs[1594] = ~(inputs[908]);
    assign layer0_outputs[1595] = (inputs[67]) | (inputs[830]);
    assign layer0_outputs[1596] = inputs[531];
    assign layer0_outputs[1597] = (inputs[683]) | (inputs[430]);
    assign layer0_outputs[1598] = ~(inputs[302]);
    assign layer0_outputs[1599] = (inputs[834]) ^ (inputs[714]);
    assign layer0_outputs[1600] = (inputs[726]) | (inputs[739]);
    assign layer0_outputs[1601] = (inputs[987]) ^ (inputs[23]);
    assign layer0_outputs[1602] = (inputs[1015]) ^ (inputs[900]);
    assign layer0_outputs[1603] = ~((inputs[264]) & (inputs[820]));
    assign layer0_outputs[1604] = 1'b1;
    assign layer0_outputs[1605] = ~(inputs[216]) | (inputs[308]);
    assign layer0_outputs[1606] = inputs[649];
    assign layer0_outputs[1607] = ~(inputs[788]);
    assign layer0_outputs[1608] = (inputs[1014]) & ~(inputs[51]);
    assign layer0_outputs[1609] = (inputs[381]) | (inputs[405]);
    assign layer0_outputs[1610] = (inputs[105]) & (inputs[314]);
    assign layer0_outputs[1611] = ~(inputs[330]) | (inputs[59]);
    assign layer0_outputs[1612] = ~(inputs[263]);
    assign layer0_outputs[1613] = ~(inputs[1012]) | (inputs[775]);
    assign layer0_outputs[1614] = ~((inputs[783]) | (inputs[902]));
    assign layer0_outputs[1615] = (inputs[811]) | (inputs[74]);
    assign layer0_outputs[1616] = ~(inputs[885]) | (inputs[469]);
    assign layer0_outputs[1617] = ~(inputs[523]);
    assign layer0_outputs[1618] = ~((inputs[1008]) | (inputs[851]));
    assign layer0_outputs[1619] = (inputs[68]) & (inputs[1007]);
    assign layer0_outputs[1620] = (inputs[738]) & (inputs[783]);
    assign layer0_outputs[1621] = ~(inputs[237]) | (inputs[982]);
    assign layer0_outputs[1622] = (inputs[688]) & ~(inputs[98]);
    assign layer0_outputs[1623] = (inputs[22]) | (inputs[16]);
    assign layer0_outputs[1624] = 1'b0;
    assign layer0_outputs[1625] = (inputs[695]) | (inputs[74]);
    assign layer0_outputs[1626] = (inputs[957]) & (inputs[893]);
    assign layer0_outputs[1627] = (inputs[160]) & ~(inputs[707]);
    assign layer0_outputs[1628] = ~((inputs[115]) & (inputs[445]));
    assign layer0_outputs[1629] = ~(inputs[848]);
    assign layer0_outputs[1630] = (inputs[178]) | (inputs[487]);
    assign layer0_outputs[1631] = inputs[716];
    assign layer0_outputs[1632] = ~((inputs[602]) | (inputs[46]));
    assign layer0_outputs[1633] = (inputs[351]) ^ (inputs[407]);
    assign layer0_outputs[1634] = (inputs[844]) & ~(inputs[839]);
    assign layer0_outputs[1635] = 1'b1;
    assign layer0_outputs[1636] = (inputs[765]) | (inputs[724]);
    assign layer0_outputs[1637] = inputs[296];
    assign layer0_outputs[1638] = (inputs[770]) & ~(inputs[646]);
    assign layer0_outputs[1639] = ~(inputs[389]) | (inputs[286]);
    assign layer0_outputs[1640] = ~((inputs[256]) | (inputs[3]));
    assign layer0_outputs[1641] = ~(inputs[917]);
    assign layer0_outputs[1642] = ~(inputs[278]) | (inputs[64]);
    assign layer0_outputs[1643] = ~(inputs[56]);
    assign layer0_outputs[1644] = inputs[400];
    assign layer0_outputs[1645] = 1'b0;
    assign layer0_outputs[1646] = ~((inputs[387]) & (inputs[208]));
    assign layer0_outputs[1647] = ~(inputs[630]) | (inputs[1010]);
    assign layer0_outputs[1648] = ~(inputs[368]) | (inputs[207]);
    assign layer0_outputs[1649] = inputs[520];
    assign layer0_outputs[1650] = (inputs[1001]) | (inputs[649]);
    assign layer0_outputs[1651] = (inputs[553]) & ~(inputs[578]);
    assign layer0_outputs[1652] = (inputs[778]) & ~(inputs[261]);
    assign layer0_outputs[1653] = (inputs[914]) & ~(inputs[542]);
    assign layer0_outputs[1654] = inputs[186];
    assign layer0_outputs[1655] = (inputs[595]) | (inputs[548]);
    assign layer0_outputs[1656] = 1'b1;
    assign layer0_outputs[1657] = ~(inputs[874]);
    assign layer0_outputs[1658] = ~(inputs[6]) | (inputs[432]);
    assign layer0_outputs[1659] = ~(inputs[124]) | (inputs[16]);
    assign layer0_outputs[1660] = ~(inputs[846]) | (inputs[372]);
    assign layer0_outputs[1661] = ~((inputs[967]) & (inputs[109]));
    assign layer0_outputs[1662] = ~(inputs[614]) | (inputs[125]);
    assign layer0_outputs[1663] = (inputs[75]) | (inputs[214]);
    assign layer0_outputs[1664] = ~((inputs[323]) ^ (inputs[172]));
    assign layer0_outputs[1665] = (inputs[230]) & ~(inputs[509]);
    assign layer0_outputs[1666] = 1'b1;
    assign layer0_outputs[1667] = inputs[1004];
    assign layer0_outputs[1668] = inputs[154];
    assign layer0_outputs[1669] = ~(inputs[925]) | (inputs[563]);
    assign layer0_outputs[1670] = ~((inputs[860]) | (inputs[278]));
    assign layer0_outputs[1671] = ~(inputs[284]);
    assign layer0_outputs[1672] = (inputs[856]) ^ (inputs[937]);
    assign layer0_outputs[1673] = (inputs[510]) & ~(inputs[88]);
    assign layer0_outputs[1674] = ~((inputs[615]) | (inputs[110]));
    assign layer0_outputs[1675] = inputs[886];
    assign layer0_outputs[1676] = ~((inputs[211]) | (inputs[822]));
    assign layer0_outputs[1677] = 1'b1;
    assign layer0_outputs[1678] = ~((inputs[411]) | (inputs[239]));
    assign layer0_outputs[1679] = ~((inputs[675]) | (inputs[277]));
    assign layer0_outputs[1680] = ~(inputs[237]) | (inputs[701]);
    assign layer0_outputs[1681] = ~(inputs[417]) | (inputs[68]);
    assign layer0_outputs[1682] = (inputs[728]) & ~(inputs[766]);
    assign layer0_outputs[1683] = ~(inputs[688]) | (inputs[541]);
    assign layer0_outputs[1684] = (inputs[814]) | (inputs[71]);
    assign layer0_outputs[1685] = ~((inputs[140]) & (inputs[240]));
    assign layer0_outputs[1686] = (inputs[389]) & ~(inputs[62]);
    assign layer0_outputs[1687] = inputs[494];
    assign layer0_outputs[1688] = ~((inputs[900]) | (inputs[879]));
    assign layer0_outputs[1689] = 1'b1;
    assign layer0_outputs[1690] = (inputs[412]) & ~(inputs[74]);
    assign layer0_outputs[1691] = inputs[754];
    assign layer0_outputs[1692] = inputs[458];
    assign layer0_outputs[1693] = (inputs[906]) & (inputs[893]);
    assign layer0_outputs[1694] = ~((inputs[910]) ^ (inputs[674]));
    assign layer0_outputs[1695] = ~((inputs[603]) & (inputs[929]));
    assign layer0_outputs[1696] = inputs[490];
    assign layer0_outputs[1697] = (inputs[364]) & ~(inputs[452]);
    assign layer0_outputs[1698] = ~((inputs[308]) ^ (inputs[4]));
    assign layer0_outputs[1699] = (inputs[398]) ^ (inputs[672]);
    assign layer0_outputs[1700] = 1'b0;
    assign layer0_outputs[1701] = (inputs[253]) ^ (inputs[266]);
    assign layer0_outputs[1702] = (inputs[48]) | (inputs[367]);
    assign layer0_outputs[1703] = (inputs[794]) ^ (inputs[540]);
    assign layer0_outputs[1704] = ~((inputs[1017]) & (inputs[852]));
    assign layer0_outputs[1705] = ~((inputs[1022]) & (inputs[372]));
    assign layer0_outputs[1706] = (inputs[449]) | (inputs[300]);
    assign layer0_outputs[1707] = ~(inputs[152]) | (inputs[761]);
    assign layer0_outputs[1708] = ~((inputs[512]) & (inputs[187]));
    assign layer0_outputs[1709] = ~((inputs[614]) ^ (inputs[49]));
    assign layer0_outputs[1710] = 1'b1;
    assign layer0_outputs[1711] = ~(inputs[845]) | (inputs[175]);
    assign layer0_outputs[1712] = (inputs[557]) & ~(inputs[632]);
    assign layer0_outputs[1713] = ~((inputs[635]) & (inputs[136]));
    assign layer0_outputs[1714] = 1'b1;
    assign layer0_outputs[1715] = ~(inputs[519]) | (inputs[657]);
    assign layer0_outputs[1716] = (inputs[711]) & ~(inputs[994]);
    assign layer0_outputs[1717] = ~((inputs[642]) & (inputs[69]));
    assign layer0_outputs[1718] = (inputs[532]) ^ (inputs[24]);
    assign layer0_outputs[1719] = ~(inputs[592]);
    assign layer0_outputs[1720] = inputs[309];
    assign layer0_outputs[1721] = (inputs[492]) & ~(inputs[262]);
    assign layer0_outputs[1722] = 1'b1;
    assign layer0_outputs[1723] = ~(inputs[587]);
    assign layer0_outputs[1724] = ~((inputs[693]) | (inputs[212]));
    assign layer0_outputs[1725] = (inputs[125]) ^ (inputs[743]);
    assign layer0_outputs[1726] = 1'b0;
    assign layer0_outputs[1727] = (inputs[602]) & (inputs[981]);
    assign layer0_outputs[1728] = inputs[303];
    assign layer0_outputs[1729] = inputs[468];
    assign layer0_outputs[1730] = ~(inputs[94]) | (inputs[408]);
    assign layer0_outputs[1731] = inputs[650];
    assign layer0_outputs[1732] = ~(inputs[652]);
    assign layer0_outputs[1733] = (inputs[333]) & ~(inputs[536]);
    assign layer0_outputs[1734] = inputs[628];
    assign layer0_outputs[1735] = ~(inputs[604]) | (inputs[806]);
    assign layer0_outputs[1736] = (inputs[777]) & ~(inputs[995]);
    assign layer0_outputs[1737] = inputs[640];
    assign layer0_outputs[1738] = ~(inputs[944]);
    assign layer0_outputs[1739] = ~(inputs[95]);
    assign layer0_outputs[1740] = ~((inputs[340]) | (inputs[294]));
    assign layer0_outputs[1741] = ~(inputs[931]) | (inputs[885]);
    assign layer0_outputs[1742] = ~(inputs[148]) | (inputs[510]);
    assign layer0_outputs[1743] = ~(inputs[806]) | (inputs[131]);
    assign layer0_outputs[1744] = ~((inputs[810]) | (inputs[412]));
    assign layer0_outputs[1745] = (inputs[560]) | (inputs[99]);
    assign layer0_outputs[1746] = ~((inputs[581]) & (inputs[1003]));
    assign layer0_outputs[1747] = inputs[810];
    assign layer0_outputs[1748] = (inputs[292]) & (inputs[948]);
    assign layer0_outputs[1749] = (inputs[0]) | (inputs[948]);
    assign layer0_outputs[1750] = ~(inputs[436]);
    assign layer0_outputs[1751] = inputs[665];
    assign layer0_outputs[1752] = 1'b1;
    assign layer0_outputs[1753] = ~((inputs[225]) | (inputs[887]));
    assign layer0_outputs[1754] = 1'b0;
    assign layer0_outputs[1755] = ~((inputs[678]) | (inputs[610]));
    assign layer0_outputs[1756] = ~(inputs[1019]) | (inputs[808]);
    assign layer0_outputs[1757] = ~((inputs[674]) & (inputs[488]));
    assign layer0_outputs[1758] = inputs[945];
    assign layer0_outputs[1759] = 1'b1;
    assign layer0_outputs[1760] = inputs[918];
    assign layer0_outputs[1761] = (inputs[75]) & ~(inputs[736]);
    assign layer0_outputs[1762] = ~((inputs[953]) & (inputs[36]));
    assign layer0_outputs[1763] = inputs[318];
    assign layer0_outputs[1764] = (inputs[414]) | (inputs[60]);
    assign layer0_outputs[1765] = 1'b0;
    assign layer0_outputs[1766] = ~(inputs[196]);
    assign layer0_outputs[1767] = ~(inputs[432]);
    assign layer0_outputs[1768] = (inputs[101]) | (inputs[446]);
    assign layer0_outputs[1769] = (inputs[433]) ^ (inputs[798]);
    assign layer0_outputs[1770] = (inputs[480]) & ~(inputs[36]);
    assign layer0_outputs[1771] = ~((inputs[864]) & (inputs[918]));
    assign layer0_outputs[1772] = (inputs[37]) & ~(inputs[440]);
    assign layer0_outputs[1773] = ~((inputs[797]) & (inputs[508]));
    assign layer0_outputs[1774] = ~((inputs[934]) ^ (inputs[108]));
    assign layer0_outputs[1775] = ~((inputs[177]) | (inputs[179]));
    assign layer0_outputs[1776] = (inputs[130]) & (inputs[491]);
    assign layer0_outputs[1777] = ~((inputs[974]) & (inputs[645]));
    assign layer0_outputs[1778] = inputs[1014];
    assign layer0_outputs[1779] = ~(inputs[128]) | (inputs[502]);
    assign layer0_outputs[1780] = ~(inputs[467]);
    assign layer0_outputs[1781] = (inputs[258]) & ~(inputs[577]);
    assign layer0_outputs[1782] = ~(inputs[230]);
    assign layer0_outputs[1783] = 1'b1;
    assign layer0_outputs[1784] = ~(inputs[813]) | (inputs[81]);
    assign layer0_outputs[1785] = (inputs[601]) | (inputs[871]);
    assign layer0_outputs[1786] = inputs[495];
    assign layer0_outputs[1787] = 1'b0;
    assign layer0_outputs[1788] = inputs[170];
    assign layer0_outputs[1789] = ~(inputs[820]);
    assign layer0_outputs[1790] = ~((inputs[826]) | (inputs[905]));
    assign layer0_outputs[1791] = (inputs[1018]) | (inputs[723]);
    assign layer0_outputs[1792] = inputs[983];
    assign layer0_outputs[1793] = ~(inputs[320]);
    assign layer0_outputs[1794] = ~((inputs[835]) & (inputs[721]));
    assign layer0_outputs[1795] = inputs[551];
    assign layer0_outputs[1796] = (inputs[806]) & (inputs[546]);
    assign layer0_outputs[1797] = 1'b0;
    assign layer0_outputs[1798] = (inputs[589]) ^ (inputs[97]);
    assign layer0_outputs[1799] = ~((inputs[235]) | (inputs[774]));
    assign layer0_outputs[1800] = (inputs[875]) | (inputs[733]);
    assign layer0_outputs[1801] = ~(inputs[818]);
    assign layer0_outputs[1802] = 1'b1;
    assign layer0_outputs[1803] = 1'b0;
    assign layer0_outputs[1804] = ~((inputs[792]) | (inputs[811]));
    assign layer0_outputs[1805] = (inputs[329]) & ~(inputs[116]);
    assign layer0_outputs[1806] = 1'b0;
    assign layer0_outputs[1807] = inputs[537];
    assign layer0_outputs[1808] = (inputs[834]) & ~(inputs[1008]);
    assign layer0_outputs[1809] = 1'b0;
    assign layer0_outputs[1810] = (inputs[191]) & ~(inputs[889]);
    assign layer0_outputs[1811] = ~((inputs[988]) ^ (inputs[163]));
    assign layer0_outputs[1812] = ~(inputs[393]) | (inputs[1008]);
    assign layer0_outputs[1813] = 1'b0;
    assign layer0_outputs[1814] = ~((inputs[957]) & (inputs[848]));
    assign layer0_outputs[1815] = (inputs[370]) & ~(inputs[1023]);
    assign layer0_outputs[1816] = (inputs[17]) ^ (inputs[681]);
    assign layer0_outputs[1817] = (inputs[66]) & ~(inputs[781]);
    assign layer0_outputs[1818] = (inputs[706]) | (inputs[281]);
    assign layer0_outputs[1819] = ~(inputs[396]);
    assign layer0_outputs[1820] = ~(inputs[449]) | (inputs[56]);
    assign layer0_outputs[1821] = ~((inputs[961]) & (inputs[686]));
    assign layer0_outputs[1822] = ~((inputs[186]) | (inputs[614]));
    assign layer0_outputs[1823] = (inputs[747]) & (inputs[361]);
    assign layer0_outputs[1824] = inputs[431];
    assign layer0_outputs[1825] = 1'b1;
    assign layer0_outputs[1826] = (inputs[722]) | (inputs[307]);
    assign layer0_outputs[1827] = (inputs[732]) & (inputs[911]);
    assign layer0_outputs[1828] = ~(inputs[696]);
    assign layer0_outputs[1829] = ~(inputs[565]);
    assign layer0_outputs[1830] = (inputs[515]) & ~(inputs[840]);
    assign layer0_outputs[1831] = ~(inputs[613]);
    assign layer0_outputs[1832] = 1'b1;
    assign layer0_outputs[1833] = (inputs[6]) | (inputs[889]);
    assign layer0_outputs[1834] = ~(inputs[71]);
    assign layer0_outputs[1835] = ~((inputs[847]) | (inputs[852]));
    assign layer0_outputs[1836] = ~(inputs[179]);
    assign layer0_outputs[1837] = 1'b1;
    assign layer0_outputs[1838] = inputs[555];
    assign layer0_outputs[1839] = (inputs[815]) | (inputs[704]);
    assign layer0_outputs[1840] = ~(inputs[678]);
    assign layer0_outputs[1841] = (inputs[593]) ^ (inputs[126]);
    assign layer0_outputs[1842] = ~(inputs[993]);
    assign layer0_outputs[1843] = ~((inputs[469]) | (inputs[764]));
    assign layer0_outputs[1844] = ~(inputs[620]);
    assign layer0_outputs[1845] = ~(inputs[141]) | (inputs[745]);
    assign layer0_outputs[1846] = (inputs[1011]) | (inputs[339]);
    assign layer0_outputs[1847] = inputs[895];
    assign layer0_outputs[1848] = (inputs[414]) & ~(inputs[837]);
    assign layer0_outputs[1849] = ~((inputs[303]) ^ (inputs[712]));
    assign layer0_outputs[1850] = (inputs[420]) & ~(inputs[422]);
    assign layer0_outputs[1851] = (inputs[827]) & ~(inputs[754]);
    assign layer0_outputs[1852] = inputs[83];
    assign layer0_outputs[1853] = 1'b1;
    assign layer0_outputs[1854] = (inputs[50]) ^ (inputs[923]);
    assign layer0_outputs[1855] = 1'b1;
    assign layer0_outputs[1856] = (inputs[771]) & ~(inputs[926]);
    assign layer0_outputs[1857] = ~(inputs[806]);
    assign layer0_outputs[1858] = (inputs[660]) | (inputs[665]);
    assign layer0_outputs[1859] = (inputs[76]) & (inputs[383]);
    assign layer0_outputs[1860] = 1'b1;
    assign layer0_outputs[1861] = (inputs[957]) ^ (inputs[898]);
    assign layer0_outputs[1862] = ~(inputs[539]);
    assign layer0_outputs[1863] = ~(inputs[808]) | (inputs[339]);
    assign layer0_outputs[1864] = 1'b0;
    assign layer0_outputs[1865] = ~(inputs[938]);
    assign layer0_outputs[1866] = (inputs[546]) & ~(inputs[515]);
    assign layer0_outputs[1867] = ~(inputs[465]);
    assign layer0_outputs[1868] = inputs[698];
    assign layer0_outputs[1869] = (inputs[717]) & ~(inputs[188]);
    assign layer0_outputs[1870] = ~((inputs[571]) | (inputs[467]));
    assign layer0_outputs[1871] = inputs[877];
    assign layer0_outputs[1872] = (inputs[118]) & ~(inputs[775]);
    assign layer0_outputs[1873] = (inputs[362]) & ~(inputs[839]);
    assign layer0_outputs[1874] = ~((inputs[634]) | (inputs[236]));
    assign layer0_outputs[1875] = ~((inputs[343]) | (inputs[1010]));
    assign layer0_outputs[1876] = ~(inputs[831]) | (inputs[128]);
    assign layer0_outputs[1877] = 1'b0;
    assign layer0_outputs[1878] = ~(inputs[144]) | (inputs[365]);
    assign layer0_outputs[1879] = ~(inputs[436]);
    assign layer0_outputs[1880] = ~((inputs[835]) | (inputs[469]));
    assign layer0_outputs[1881] = (inputs[363]) | (inputs[873]);
    assign layer0_outputs[1882] = (inputs[226]) & (inputs[267]);
    assign layer0_outputs[1883] = ~(inputs[226]) | (inputs[554]);
    assign layer0_outputs[1884] = ~((inputs[413]) | (inputs[848]));
    assign layer0_outputs[1885] = (inputs[104]) & (inputs[972]);
    assign layer0_outputs[1886] = ~(inputs[397]);
    assign layer0_outputs[1887] = ~(inputs[525]) | (inputs[715]);
    assign layer0_outputs[1888] = (inputs[242]) ^ (inputs[371]);
    assign layer0_outputs[1889] = ~((inputs[400]) | (inputs[741]));
    assign layer0_outputs[1890] = (inputs[808]) | (inputs[809]);
    assign layer0_outputs[1891] = ~(inputs[563]);
    assign layer0_outputs[1892] = (inputs[84]) | (inputs[821]);
    assign layer0_outputs[1893] = ~(inputs[458]);
    assign layer0_outputs[1894] = (inputs[392]) | (inputs[689]);
    assign layer0_outputs[1895] = 1'b0;
    assign layer0_outputs[1896] = ~((inputs[566]) | (inputs[141]));
    assign layer0_outputs[1897] = inputs[527];
    assign layer0_outputs[1898] = ~((inputs[915]) | (inputs[992]));
    assign layer0_outputs[1899] = (inputs[273]) & ~(inputs[882]);
    assign layer0_outputs[1900] = (inputs[625]) & ~(inputs[235]);
    assign layer0_outputs[1901] = 1'b0;
    assign layer0_outputs[1902] = ~(inputs[681]);
    assign layer0_outputs[1903] = (inputs[287]) ^ (inputs[1013]);
    assign layer0_outputs[1904] = inputs[605];
    assign layer0_outputs[1905] = 1'b0;
    assign layer0_outputs[1906] = ~(inputs[190]);
    assign layer0_outputs[1907] = ~((inputs[65]) | (inputs[68]));
    assign layer0_outputs[1908] = ~(inputs[207]) | (inputs[385]);
    assign layer0_outputs[1909] = ~(inputs[52]) | (inputs[548]);
    assign layer0_outputs[1910] = ~((inputs[233]) | (inputs[705]));
    assign layer0_outputs[1911] = (inputs[116]) & ~(inputs[344]);
    assign layer0_outputs[1912] = inputs[240];
    assign layer0_outputs[1913] = ~(inputs[518]) | (inputs[922]);
    assign layer0_outputs[1914] = (inputs[974]) | (inputs[724]);
    assign layer0_outputs[1915] = (inputs[826]) & (inputs[47]);
    assign layer0_outputs[1916] = 1'b1;
    assign layer0_outputs[1917] = (inputs[513]) ^ (inputs[591]);
    assign layer0_outputs[1918] = (inputs[254]) & (inputs[939]);
    assign layer0_outputs[1919] = 1'b1;
    assign layer0_outputs[1920] = (inputs[280]) ^ (inputs[1010]);
    assign layer0_outputs[1921] = (inputs[527]) & ~(inputs[397]);
    assign layer0_outputs[1922] = 1'b1;
    assign layer0_outputs[1923] = (inputs[565]) & (inputs[984]);
    assign layer0_outputs[1924] = ~((inputs[128]) ^ (inputs[574]));
    assign layer0_outputs[1925] = (inputs[315]) | (inputs[345]);
    assign layer0_outputs[1926] = 1'b0;
    assign layer0_outputs[1927] = 1'b1;
    assign layer0_outputs[1928] = ~((inputs[426]) & (inputs[743]));
    assign layer0_outputs[1929] = ~(inputs[115]) | (inputs[1016]);
    assign layer0_outputs[1930] = 1'b0;
    assign layer0_outputs[1931] = (inputs[137]) & ~(inputs[391]);
    assign layer0_outputs[1932] = inputs[208];
    assign layer0_outputs[1933] = (inputs[643]) & (inputs[442]);
    assign layer0_outputs[1934] = 1'b0;
    assign layer0_outputs[1935] = (inputs[29]) | (inputs[636]);
    assign layer0_outputs[1936] = ~(inputs[280]);
    assign layer0_outputs[1937] = (inputs[833]) & ~(inputs[508]);
    assign layer0_outputs[1938] = 1'b1;
    assign layer0_outputs[1939] = ~(inputs[537]) | (inputs[151]);
    assign layer0_outputs[1940] = ~(inputs[166]);
    assign layer0_outputs[1941] = (inputs[147]) & ~(inputs[168]);
    assign layer0_outputs[1942] = inputs[312];
    assign layer0_outputs[1943] = ~(inputs[400]) | (inputs[509]);
    assign layer0_outputs[1944] = (inputs[939]) | (inputs[920]);
    assign layer0_outputs[1945] = inputs[460];
    assign layer0_outputs[1946] = (inputs[380]) & ~(inputs[943]);
    assign layer0_outputs[1947] = 1'b0;
    assign layer0_outputs[1948] = (inputs[588]) | (inputs[67]);
    assign layer0_outputs[1949] = inputs[104];
    assign layer0_outputs[1950] = (inputs[167]) | (inputs[893]);
    assign layer0_outputs[1951] = ~(inputs[525]);
    assign layer0_outputs[1952] = ~(inputs[524]);
    assign layer0_outputs[1953] = ~(inputs[807]) | (inputs[390]);
    assign layer0_outputs[1954] = ~((inputs[783]) & (inputs[670]));
    assign layer0_outputs[1955] = ~(inputs[393]) | (inputs[221]);
    assign layer0_outputs[1956] = (inputs[619]) | (inputs[133]);
    assign layer0_outputs[1957] = ~((inputs[488]) | (inputs[534]));
    assign layer0_outputs[1958] = ~((inputs[248]) ^ (inputs[475]));
    assign layer0_outputs[1959] = ~(inputs[919]);
    assign layer0_outputs[1960] = 1'b1;
    assign layer0_outputs[1961] = (inputs[859]) & ~(inputs[279]);
    assign layer0_outputs[1962] = ~((inputs[327]) & (inputs[382]));
    assign layer0_outputs[1963] = inputs[370];
    assign layer0_outputs[1964] = ~(inputs[696]);
    assign layer0_outputs[1965] = 1'b0;
    assign layer0_outputs[1966] = ~((inputs[885]) | (inputs[428]));
    assign layer0_outputs[1967] = (inputs[551]) ^ (inputs[984]);
    assign layer0_outputs[1968] = 1'b0;
    assign layer0_outputs[1969] = ~((inputs[540]) | (inputs[651]));
    assign layer0_outputs[1970] = (inputs[596]) & ~(inputs[43]);
    assign layer0_outputs[1971] = 1'b1;
    assign layer0_outputs[1972] = ~(inputs[415]) | (inputs[628]);
    assign layer0_outputs[1973] = 1'b1;
    assign layer0_outputs[1974] = inputs[702];
    assign layer0_outputs[1975] = 1'b1;
    assign layer0_outputs[1976] = (inputs[375]) & ~(inputs[939]);
    assign layer0_outputs[1977] = ~(inputs[275]);
    assign layer0_outputs[1978] = (inputs[355]) & ~(inputs[613]);
    assign layer0_outputs[1979] = inputs[394];
    assign layer0_outputs[1980] = ~((inputs[521]) | (inputs[730]));
    assign layer0_outputs[1981] = ~((inputs[52]) ^ (inputs[890]));
    assign layer0_outputs[1982] = ~(inputs[641]) | (inputs[606]);
    assign layer0_outputs[1983] = ~(inputs[706]) | (inputs[201]);
    assign layer0_outputs[1984] = (inputs[194]) & ~(inputs[933]);
    assign layer0_outputs[1985] = ~(inputs[478]) | (inputs[32]);
    assign layer0_outputs[1986] = (inputs[328]) & ~(inputs[1]);
    assign layer0_outputs[1987] = ~((inputs[765]) | (inputs[103]));
    assign layer0_outputs[1988] = (inputs[86]) | (inputs[3]);
    assign layer0_outputs[1989] = ~(inputs[357]) | (inputs[215]);
    assign layer0_outputs[1990] = (inputs[836]) | (inputs[647]);
    assign layer0_outputs[1991] = ~(inputs[941]);
    assign layer0_outputs[1992] = 1'b1;
    assign layer0_outputs[1993] = 1'b0;
    assign layer0_outputs[1994] = ~(inputs[900]) | (inputs[1005]);
    assign layer0_outputs[1995] = ~((inputs[718]) | (inputs[186]));
    assign layer0_outputs[1996] = (inputs[487]) | (inputs[510]);
    assign layer0_outputs[1997] = (inputs[223]) ^ (inputs[616]);
    assign layer0_outputs[1998] = (inputs[427]) & ~(inputs[960]);
    assign layer0_outputs[1999] = ~((inputs[454]) | (inputs[596]));
    assign layer0_outputs[2000] = ~(inputs[165]);
    assign layer0_outputs[2001] = ~(inputs[746]) | (inputs[488]);
    assign layer0_outputs[2002] = (inputs[22]) | (inputs[266]);
    assign layer0_outputs[2003] = inputs[203];
    assign layer0_outputs[2004] = (inputs[676]) | (inputs[403]);
    assign layer0_outputs[2005] = (inputs[539]) | (inputs[765]);
    assign layer0_outputs[2006] = 1'b1;
    assign layer0_outputs[2007] = (inputs[150]) & (inputs[855]);
    assign layer0_outputs[2008] = (inputs[708]) ^ (inputs[70]);
    assign layer0_outputs[2009] = ~(inputs[715]);
    assign layer0_outputs[2010] = (inputs[755]) ^ (inputs[291]);
    assign layer0_outputs[2011] = (inputs[955]) & ~(inputs[986]);
    assign layer0_outputs[2012] = ~(inputs[524]);
    assign layer0_outputs[2013] = (inputs[672]) | (inputs[467]);
    assign layer0_outputs[2014] = ~((inputs[388]) | (inputs[997]));
    assign layer0_outputs[2015] = (inputs[921]) ^ (inputs[770]);
    assign layer0_outputs[2016] = (inputs[410]) & ~(inputs[568]);
    assign layer0_outputs[2017] = ~((inputs[538]) | (inputs[210]));
    assign layer0_outputs[2018] = ~((inputs[256]) | (inputs[298]));
    assign layer0_outputs[2019] = 1'b1;
    assign layer0_outputs[2020] = ~((inputs[231]) & (inputs[452]));
    assign layer0_outputs[2021] = inputs[633];
    assign layer0_outputs[2022] = ~(inputs[657]) | (inputs[509]);
    assign layer0_outputs[2023] = (inputs[181]) | (inputs[663]);
    assign layer0_outputs[2024] = 1'b0;
    assign layer0_outputs[2025] = (inputs[473]) | (inputs[366]);
    assign layer0_outputs[2026] = ~((inputs[482]) | (inputs[808]));
    assign layer0_outputs[2027] = 1'b1;
    assign layer0_outputs[2028] = ~(inputs[599]);
    assign layer0_outputs[2029] = inputs[329];
    assign layer0_outputs[2030] = ~((inputs[165]) | (inputs[1020]));
    assign layer0_outputs[2031] = (inputs[517]) & ~(inputs[479]);
    assign layer0_outputs[2032] = ~((inputs[450]) | (inputs[624]));
    assign layer0_outputs[2033] = 1'b1;
    assign layer0_outputs[2034] = 1'b1;
    assign layer0_outputs[2035] = inputs[782];
    assign layer0_outputs[2036] = inputs[715];
    assign layer0_outputs[2037] = ~(inputs[666]) | (inputs[1015]);
    assign layer0_outputs[2038] = 1'b0;
    assign layer0_outputs[2039] = (inputs[213]) | (inputs[444]);
    assign layer0_outputs[2040] = (inputs[269]) & ~(inputs[531]);
    assign layer0_outputs[2041] = inputs[957];
    assign layer0_outputs[2042] = ~(inputs[979]) | (inputs[60]);
    assign layer0_outputs[2043] = ~(inputs[7]);
    assign layer0_outputs[2044] = (inputs[335]) & ~(inputs[546]);
    assign layer0_outputs[2045] = ~((inputs[881]) | (inputs[450]));
    assign layer0_outputs[2046] = ~((inputs[604]) | (inputs[10]));
    assign layer0_outputs[2047] = ~(inputs[741]) | (inputs[911]);
    assign layer0_outputs[2048] = inputs[403];
    assign layer0_outputs[2049] = ~(inputs[582]) | (inputs[181]);
    assign layer0_outputs[2050] = ~(inputs[221]) | (inputs[830]);
    assign layer0_outputs[2051] = ~(inputs[478]) | (inputs[391]);
    assign layer0_outputs[2052] = (inputs[50]) & ~(inputs[680]);
    assign layer0_outputs[2053] = ~(inputs[144]) | (inputs[363]);
    assign layer0_outputs[2054] = inputs[92];
    assign layer0_outputs[2055] = ~(inputs[618]);
    assign layer0_outputs[2056] = 1'b1;
    assign layer0_outputs[2057] = 1'b0;
    assign layer0_outputs[2058] = inputs[892];
    assign layer0_outputs[2059] = ~(inputs[979]);
    assign layer0_outputs[2060] = ~((inputs[299]) ^ (inputs[1012]));
    assign layer0_outputs[2061] = (inputs[690]) | (inputs[867]);
    assign layer0_outputs[2062] = 1'b0;
    assign layer0_outputs[2063] = inputs[728];
    assign layer0_outputs[2064] = inputs[374];
    assign layer0_outputs[2065] = ~((inputs[231]) | (inputs[763]));
    assign layer0_outputs[2066] = ~((inputs[185]) | (inputs[161]));
    assign layer0_outputs[2067] = (inputs[822]) | (inputs[209]);
    assign layer0_outputs[2068] = ~(inputs[238]);
    assign layer0_outputs[2069] = ~((inputs[479]) & (inputs[979]));
    assign layer0_outputs[2070] = ~((inputs[545]) | (inputs[442]));
    assign layer0_outputs[2071] = (inputs[171]) & ~(inputs[800]);
    assign layer0_outputs[2072] = ~(inputs[615]) | (inputs[136]);
    assign layer0_outputs[2073] = 1'b1;
    assign layer0_outputs[2074] = (inputs[14]) & ~(inputs[978]);
    assign layer0_outputs[2075] = (inputs[182]) & ~(inputs[191]);
    assign layer0_outputs[2076] = (inputs[19]) & (inputs[560]);
    assign layer0_outputs[2077] = (inputs[262]) & ~(inputs[660]);
    assign layer0_outputs[2078] = ~((inputs[572]) | (inputs[998]));
    assign layer0_outputs[2079] = (inputs[398]) & (inputs[769]);
    assign layer0_outputs[2080] = (inputs[1013]) & (inputs[89]);
    assign layer0_outputs[2081] = (inputs[503]) | (inputs[556]);
    assign layer0_outputs[2082] = (inputs[765]) & ~(inputs[915]);
    assign layer0_outputs[2083] = ~(inputs[368]);
    assign layer0_outputs[2084] = inputs[258];
    assign layer0_outputs[2085] = ~((inputs[988]) | (inputs[647]));
    assign layer0_outputs[2086] = (inputs[912]) & ~(inputs[841]);
    assign layer0_outputs[2087] = ~((inputs[47]) | (inputs[315]));
    assign layer0_outputs[2088] = inputs[370];
    assign layer0_outputs[2089] = inputs[9];
    assign layer0_outputs[2090] = inputs[434];
    assign layer0_outputs[2091] = (inputs[314]) | (inputs[942]);
    assign layer0_outputs[2092] = 1'b0;
    assign layer0_outputs[2093] = ~(inputs[995]);
    assign layer0_outputs[2094] = inputs[455];
    assign layer0_outputs[2095] = ~(inputs[432]);
    assign layer0_outputs[2096] = ~((inputs[352]) & (inputs[853]));
    assign layer0_outputs[2097] = ~(inputs[71]) | (inputs[980]);
    assign layer0_outputs[2098] = ~(inputs[471]);
    assign layer0_outputs[2099] = (inputs[986]) & ~(inputs[855]);
    assign layer0_outputs[2100] = (inputs[66]) & (inputs[758]);
    assign layer0_outputs[2101] = ~((inputs[530]) | (inputs[79]));
    assign layer0_outputs[2102] = ~(inputs[815]);
    assign layer0_outputs[2103] = (inputs[928]) & (inputs[187]);
    assign layer0_outputs[2104] = ~(inputs[629]);
    assign layer0_outputs[2105] = inputs[539];
    assign layer0_outputs[2106] = inputs[990];
    assign layer0_outputs[2107] = inputs[804];
    assign layer0_outputs[2108] = inputs[808];
    assign layer0_outputs[2109] = 1'b0;
    assign layer0_outputs[2110] = (inputs[364]) & ~(inputs[670]);
    assign layer0_outputs[2111] = ~((inputs[72]) & (inputs[976]));
    assign layer0_outputs[2112] = (inputs[228]) & (inputs[829]);
    assign layer0_outputs[2113] = inputs[807];
    assign layer0_outputs[2114] = ~(inputs[625]);
    assign layer0_outputs[2115] = ~(inputs[230]);
    assign layer0_outputs[2116] = ~(inputs[620]);
    assign layer0_outputs[2117] = (inputs[444]) ^ (inputs[334]);
    assign layer0_outputs[2118] = ~(inputs[472]);
    assign layer0_outputs[2119] = (inputs[700]) | (inputs[575]);
    assign layer0_outputs[2120] = inputs[295];
    assign layer0_outputs[2121] = (inputs[877]) & (inputs[145]);
    assign layer0_outputs[2122] = ~(inputs[345]) | (inputs[559]);
    assign layer0_outputs[2123] = (inputs[747]) & (inputs[254]);
    assign layer0_outputs[2124] = (inputs[5]) & ~(inputs[601]);
    assign layer0_outputs[2125] = ~((inputs[953]) | (inputs[346]));
    assign layer0_outputs[2126] = ~(inputs[97]) | (inputs[816]);
    assign layer0_outputs[2127] = ~((inputs[1007]) & (inputs[556]));
    assign layer0_outputs[2128] = 1'b1;
    assign layer0_outputs[2129] = (inputs[729]) | (inputs[1009]);
    assign layer0_outputs[2130] = ~(inputs[828]);
    assign layer0_outputs[2131] = ~((inputs[552]) | (inputs[966]));
    assign layer0_outputs[2132] = 1'b1;
    assign layer0_outputs[2133] = ~((inputs[224]) & (inputs[173]));
    assign layer0_outputs[2134] = ~(inputs[82]);
    assign layer0_outputs[2135] = ~(inputs[461]);
    assign layer0_outputs[2136] = inputs[552];
    assign layer0_outputs[2137] = inputs[654];
    assign layer0_outputs[2138] = ~((inputs[632]) | (inputs[493]));
    assign layer0_outputs[2139] = ~(inputs[276]) | (inputs[650]);
    assign layer0_outputs[2140] = ~(inputs[991]);
    assign layer0_outputs[2141] = (inputs[294]) | (inputs[921]);
    assign layer0_outputs[2142] = (inputs[828]) | (inputs[930]);
    assign layer0_outputs[2143] = ~(inputs[451]) | (inputs[735]);
    assign layer0_outputs[2144] = ~(inputs[568]) | (inputs[883]);
    assign layer0_outputs[2145] = (inputs[76]) | (inputs[559]);
    assign layer0_outputs[2146] = (inputs[827]) & (inputs[661]);
    assign layer0_outputs[2147] = (inputs[1016]) | (inputs[787]);
    assign layer0_outputs[2148] = ~(inputs[242]);
    assign layer0_outputs[2149] = ~(inputs[686]);
    assign layer0_outputs[2150] = (inputs[865]) & ~(inputs[879]);
    assign layer0_outputs[2151] = ~((inputs[416]) ^ (inputs[711]));
    assign layer0_outputs[2152] = inputs[741];
    assign layer0_outputs[2153] = 1'b0;
    assign layer0_outputs[2154] = ~(inputs[16]);
    assign layer0_outputs[2155] = (inputs[352]) | (inputs[703]);
    assign layer0_outputs[2156] = (inputs[702]) & (inputs[836]);
    assign layer0_outputs[2157] = ~((inputs[269]) & (inputs[221]));
    assign layer0_outputs[2158] = ~((inputs[669]) | (inputs[244]));
    assign layer0_outputs[2159] = (inputs[667]) | (inputs[107]);
    assign layer0_outputs[2160] = ~(inputs[784]);
    assign layer0_outputs[2161] = ~((inputs[684]) & (inputs[489]));
    assign layer0_outputs[2162] = ~((inputs[611]) & (inputs[959]));
    assign layer0_outputs[2163] = ~(inputs[510]) | (inputs[987]);
    assign layer0_outputs[2164] = (inputs[288]) ^ (inputs[958]);
    assign layer0_outputs[2165] = (inputs[175]) & (inputs[8]);
    assign layer0_outputs[2166] = ~(inputs[385]);
    assign layer0_outputs[2167] = inputs[646];
    assign layer0_outputs[2168] = ~(inputs[556]);
    assign layer0_outputs[2169] = ~(inputs[266]) | (inputs[505]);
    assign layer0_outputs[2170] = inputs[943];
    assign layer0_outputs[2171] = (inputs[213]) | (inputs[561]);
    assign layer0_outputs[2172] = (inputs[35]) & ~(inputs[310]);
    assign layer0_outputs[2173] = (inputs[107]) & ~(inputs[961]);
    assign layer0_outputs[2174] = (inputs[1016]) & ~(inputs[347]);
    assign layer0_outputs[2175] = (inputs[787]) | (inputs[649]);
    assign layer0_outputs[2176] = ~((inputs[591]) | (inputs[991]));
    assign layer0_outputs[2177] = (inputs[172]) | (inputs[42]);
    assign layer0_outputs[2178] = (inputs[585]) | (inputs[531]);
    assign layer0_outputs[2179] = (inputs[184]) & (inputs[155]);
    assign layer0_outputs[2180] = inputs[211];
    assign layer0_outputs[2181] = (inputs[222]) & ~(inputs[746]);
    assign layer0_outputs[2182] = (inputs[141]) & (inputs[539]);
    assign layer0_outputs[2183] = (inputs[396]) & ~(inputs[199]);
    assign layer0_outputs[2184] = 1'b1;
    assign layer0_outputs[2185] = (inputs[561]) | (inputs[837]);
    assign layer0_outputs[2186] = ~(inputs[817]) | (inputs[157]);
    assign layer0_outputs[2187] = ~(inputs[781]);
    assign layer0_outputs[2188] = ~(inputs[562]);
    assign layer0_outputs[2189] = (inputs[754]) & ~(inputs[350]);
    assign layer0_outputs[2190] = 1'b1;
    assign layer0_outputs[2191] = ~((inputs[502]) & (inputs[579]));
    assign layer0_outputs[2192] = (inputs[958]) ^ (inputs[720]);
    assign layer0_outputs[2193] = 1'b1;
    assign layer0_outputs[2194] = (inputs[145]) & ~(inputs[219]);
    assign layer0_outputs[2195] = 1'b1;
    assign layer0_outputs[2196] = ~((inputs[238]) | (inputs[170]));
    assign layer0_outputs[2197] = ~(inputs[633]);
    assign layer0_outputs[2198] = ~((inputs[272]) | (inputs[799]));
    assign layer0_outputs[2199] = ~(inputs[936]);
    assign layer0_outputs[2200] = (inputs[430]) ^ (inputs[505]);
    assign layer0_outputs[2201] = ~(inputs[15]);
    assign layer0_outputs[2202] = (inputs[170]) | (inputs[117]);
    assign layer0_outputs[2203] = (inputs[242]) & (inputs[756]);
    assign layer0_outputs[2204] = 1'b1;
    assign layer0_outputs[2205] = (inputs[1020]) & (inputs[380]);
    assign layer0_outputs[2206] = ~(inputs[627]) | (inputs[577]);
    assign layer0_outputs[2207] = ~(inputs[832]);
    assign layer0_outputs[2208] = (inputs[297]) & (inputs[420]);
    assign layer0_outputs[2209] = inputs[1006];
    assign layer0_outputs[2210] = ~(inputs[260]) | (inputs[41]);
    assign layer0_outputs[2211] = inputs[673];
    assign layer0_outputs[2212] = (inputs[197]) & ~(inputs[308]);
    assign layer0_outputs[2213] = (inputs[792]) & ~(inputs[121]);
    assign layer0_outputs[2214] = ~((inputs[13]) & (inputs[262]));
    assign layer0_outputs[2215] = (inputs[448]) | (inputs[508]);
    assign layer0_outputs[2216] = (inputs[588]) | (inputs[46]);
    assign layer0_outputs[2217] = ~((inputs[382]) ^ (inputs[826]));
    assign layer0_outputs[2218] = ~((inputs[379]) ^ (inputs[239]));
    assign layer0_outputs[2219] = ~((inputs[550]) | (inputs[663]));
    assign layer0_outputs[2220] = inputs[624];
    assign layer0_outputs[2221] = ~(inputs[282]) | (inputs[153]);
    assign layer0_outputs[2222] = ~((inputs[791]) | (inputs[388]));
    assign layer0_outputs[2223] = (inputs[612]) & ~(inputs[602]);
    assign layer0_outputs[2224] = (inputs[549]) & (inputs[132]);
    assign layer0_outputs[2225] = (inputs[28]) | (inputs[199]);
    assign layer0_outputs[2226] = (inputs[600]) | (inputs[232]);
    assign layer0_outputs[2227] = (inputs[91]) & (inputs[825]);
    assign layer0_outputs[2228] = ~(inputs[768]);
    assign layer0_outputs[2229] = (inputs[495]) | (inputs[680]);
    assign layer0_outputs[2230] = (inputs[926]) | (inputs[242]);
    assign layer0_outputs[2231] = ~(inputs[476]);
    assign layer0_outputs[2232] = (inputs[954]) | (inputs[862]);
    assign layer0_outputs[2233] = (inputs[634]) & ~(inputs[369]);
    assign layer0_outputs[2234] = (inputs[926]) & ~(inputs[352]);
    assign layer0_outputs[2235] = (inputs[385]) & ~(inputs[125]);
    assign layer0_outputs[2236] = (inputs[951]) | (inputs[421]);
    assign layer0_outputs[2237] = ~(inputs[529]) | (inputs[537]);
    assign layer0_outputs[2238] = (inputs[64]) & ~(inputs[851]);
    assign layer0_outputs[2239] = (inputs[20]) & ~(inputs[111]);
    assign layer0_outputs[2240] = (inputs[68]) | (inputs[534]);
    assign layer0_outputs[2241] = ~(inputs[745]);
    assign layer0_outputs[2242] = 1'b0;
    assign layer0_outputs[2243] = (inputs[462]) | (inputs[40]);
    assign layer0_outputs[2244] = inputs[687];
    assign layer0_outputs[2245] = inputs[936];
    assign layer0_outputs[2246] = 1'b0;
    assign layer0_outputs[2247] = (inputs[103]) | (inputs[389]);
    assign layer0_outputs[2248] = inputs[586];
    assign layer0_outputs[2249] = ~(inputs[371]);
    assign layer0_outputs[2250] = inputs[881];
    assign layer0_outputs[2251] = (inputs[326]) | (inputs[363]);
    assign layer0_outputs[2252] = (inputs[651]) ^ (inputs[230]);
    assign layer0_outputs[2253] = ~(inputs[846]);
    assign layer0_outputs[2254] = (inputs[546]) | (inputs[662]);
    assign layer0_outputs[2255] = (inputs[43]) & (inputs[90]);
    assign layer0_outputs[2256] = (inputs[653]) & ~(inputs[220]);
    assign layer0_outputs[2257] = ~(inputs[733]);
    assign layer0_outputs[2258] = inputs[652];
    assign layer0_outputs[2259] = 1'b0;
    assign layer0_outputs[2260] = (inputs[438]) & ~(inputs[698]);
    assign layer0_outputs[2261] = inputs[620];
    assign layer0_outputs[2262] = inputs[148];
    assign layer0_outputs[2263] = (inputs[946]) ^ (inputs[679]);
    assign layer0_outputs[2264] = ~((inputs[732]) | (inputs[166]));
    assign layer0_outputs[2265] = inputs[710];
    assign layer0_outputs[2266] = ~(inputs[401]);
    assign layer0_outputs[2267] = 1'b0;
    assign layer0_outputs[2268] = ~((inputs[757]) | (inputs[867]));
    assign layer0_outputs[2269] = (inputs[658]) & ~(inputs[216]);
    assign layer0_outputs[2270] = ~((inputs[603]) & (inputs[499]));
    assign layer0_outputs[2271] = ~((inputs[365]) | (inputs[377]));
    assign layer0_outputs[2272] = ~((inputs[953]) & (inputs[251]));
    assign layer0_outputs[2273] = ~(inputs[236]) | (inputs[540]);
    assign layer0_outputs[2274] = 1'b1;
    assign layer0_outputs[2275] = ~((inputs[3]) | (inputs[863]));
    assign layer0_outputs[2276] = ~((inputs[669]) ^ (inputs[727]));
    assign layer0_outputs[2277] = ~((inputs[693]) | (inputs[202]));
    assign layer0_outputs[2278] = ~((inputs[87]) ^ (inputs[290]));
    assign layer0_outputs[2279] = inputs[906];
    assign layer0_outputs[2280] = ~(inputs[629]);
    assign layer0_outputs[2281] = ~((inputs[455]) ^ (inputs[197]));
    assign layer0_outputs[2282] = (inputs[863]) ^ (inputs[59]);
    assign layer0_outputs[2283] = (inputs[960]) & ~(inputs[570]);
    assign layer0_outputs[2284] = inputs[941];
    assign layer0_outputs[2285] = 1'b1;
    assign layer0_outputs[2286] = 1'b0;
    assign layer0_outputs[2287] = ~(inputs[437]) | (inputs[511]);
    assign layer0_outputs[2288] = 1'b0;
    assign layer0_outputs[2289] = 1'b0;
    assign layer0_outputs[2290] = (inputs[922]) ^ (inputs[886]);
    assign layer0_outputs[2291] = inputs[702];
    assign layer0_outputs[2292] = 1'b1;
    assign layer0_outputs[2293] = ~((inputs[363]) ^ (inputs[25]));
    assign layer0_outputs[2294] = inputs[35];
    assign layer0_outputs[2295] = (inputs[156]) ^ (inputs[136]);
    assign layer0_outputs[2296] = ~((inputs[379]) | (inputs[301]));
    assign layer0_outputs[2297] = (inputs[476]) & ~(inputs[798]);
    assign layer0_outputs[2298] = (inputs[506]) | (inputs[779]);
    assign layer0_outputs[2299] = (inputs[679]) | (inputs[410]);
    assign layer0_outputs[2300] = inputs[410];
    assign layer0_outputs[2301] = 1'b1;
    assign layer0_outputs[2302] = inputs[272];
    assign layer0_outputs[2303] = 1'b1;
    assign layer0_outputs[2304] = inputs[776];
    assign layer0_outputs[2305] = ~(inputs[567]) | (inputs[873]);
    assign layer0_outputs[2306] = inputs[83];
    assign layer0_outputs[2307] = ~(inputs[578]);
    assign layer0_outputs[2308] = inputs[253];
    assign layer0_outputs[2309] = inputs[211];
    assign layer0_outputs[2310] = inputs[718];
    assign layer0_outputs[2311] = (inputs[909]) ^ (inputs[801]);
    assign layer0_outputs[2312] = (inputs[687]) & ~(inputs[456]);
    assign layer0_outputs[2313] = (inputs[173]) & ~(inputs[666]);
    assign layer0_outputs[2314] = ~(inputs[147]);
    assign layer0_outputs[2315] = (inputs[48]) & (inputs[246]);
    assign layer0_outputs[2316] = ~(inputs[360]);
    assign layer0_outputs[2317] = (inputs[359]) & ~(inputs[119]);
    assign layer0_outputs[2318] = ~((inputs[829]) ^ (inputs[283]));
    assign layer0_outputs[2319] = ~((inputs[441]) | (inputs[178]));
    assign layer0_outputs[2320] = ~(inputs[459]);
    assign layer0_outputs[2321] = 1'b1;
    assign layer0_outputs[2322] = ~((inputs[263]) | (inputs[745]));
    assign layer0_outputs[2323] = (inputs[505]) & ~(inputs[627]);
    assign layer0_outputs[2324] = (inputs[323]) & ~(inputs[733]);
    assign layer0_outputs[2325] = 1'b1;
    assign layer0_outputs[2326] = ~((inputs[70]) ^ (inputs[918]));
    assign layer0_outputs[2327] = ~(inputs[783]) | (inputs[693]);
    assign layer0_outputs[2328] = 1'b0;
    assign layer0_outputs[2329] = (inputs[199]) ^ (inputs[62]);
    assign layer0_outputs[2330] = ~((inputs[842]) | (inputs[411]));
    assign layer0_outputs[2331] = ~(inputs[195]);
    assign layer0_outputs[2332] = ~(inputs[518]) | (inputs[104]);
    assign layer0_outputs[2333] = ~((inputs[227]) | (inputs[163]));
    assign layer0_outputs[2334] = 1'b0;
    assign layer0_outputs[2335] = ~((inputs[936]) | (inputs[818]));
    assign layer0_outputs[2336] = (inputs[0]) & (inputs[897]);
    assign layer0_outputs[2337] = (inputs[998]) & ~(inputs[974]);
    assign layer0_outputs[2338] = ~(inputs[405]) | (inputs[584]);
    assign layer0_outputs[2339] = (inputs[670]) & (inputs[559]);
    assign layer0_outputs[2340] = ~((inputs[571]) | (inputs[417]));
    assign layer0_outputs[2341] = 1'b1;
    assign layer0_outputs[2342] = ~(inputs[540]);
    assign layer0_outputs[2343] = (inputs[527]) & (inputs[795]);
    assign layer0_outputs[2344] = inputs[876];
    assign layer0_outputs[2345] = ~(inputs[465]) | (inputs[324]);
    assign layer0_outputs[2346] = ~((inputs[690]) | (inputs[998]));
    assign layer0_outputs[2347] = ~(inputs[505]);
    assign layer0_outputs[2348] = ~((inputs[888]) ^ (inputs[34]));
    assign layer0_outputs[2349] = inputs[526];
    assign layer0_outputs[2350] = ~((inputs[417]) ^ (inputs[123]));
    assign layer0_outputs[2351] = ~(inputs[491]);
    assign layer0_outputs[2352] = ~(inputs[456]) | (inputs[26]);
    assign layer0_outputs[2353] = (inputs[896]) ^ (inputs[428]);
    assign layer0_outputs[2354] = (inputs[151]) | (inputs[752]);
    assign layer0_outputs[2355] = inputs[188];
    assign layer0_outputs[2356] = 1'b1;
    assign layer0_outputs[2357] = ~(inputs[564]) | (inputs[419]);
    assign layer0_outputs[2358] = inputs[746];
    assign layer0_outputs[2359] = ~((inputs[774]) | (inputs[871]));
    assign layer0_outputs[2360] = (inputs[889]) & ~(inputs[677]);
    assign layer0_outputs[2361] = ~(inputs[139]) | (inputs[782]);
    assign layer0_outputs[2362] = ~(inputs[869]) | (inputs[879]);
    assign layer0_outputs[2363] = ~(inputs[784]);
    assign layer0_outputs[2364] = (inputs[909]) & (inputs[719]);
    assign layer0_outputs[2365] = inputs[596];
    assign layer0_outputs[2366] = (inputs[450]) & ~(inputs[226]);
    assign layer0_outputs[2367] = ~(inputs[563]);
    assign layer0_outputs[2368] = ~(inputs[149]);
    assign layer0_outputs[2369] = 1'b1;
    assign layer0_outputs[2370] = (inputs[387]) & ~(inputs[111]);
    assign layer0_outputs[2371] = ~(inputs[362]) | (inputs[739]);
    assign layer0_outputs[2372] = 1'b1;
    assign layer0_outputs[2373] = 1'b1;
    assign layer0_outputs[2374] = ~((inputs[98]) | (inputs[7]));
    assign layer0_outputs[2375] = ~(inputs[543]);
    assign layer0_outputs[2376] = 1'b1;
    assign layer0_outputs[2377] = (inputs[722]) ^ (inputs[11]);
    assign layer0_outputs[2378] = ~((inputs[854]) | (inputs[406]));
    assign layer0_outputs[2379] = ~(inputs[645]);
    assign layer0_outputs[2380] = inputs[312];
    assign layer0_outputs[2381] = (inputs[592]) ^ (inputs[163]);
    assign layer0_outputs[2382] = ~((inputs[477]) | (inputs[772]));
    assign layer0_outputs[2383] = (inputs[297]) | (inputs[965]);
    assign layer0_outputs[2384] = inputs[947];
    assign layer0_outputs[2385] = ~(inputs[435]);
    assign layer0_outputs[2386] = ~(inputs[945]) | (inputs[477]);
    assign layer0_outputs[2387] = ~(inputs[572]);
    assign layer0_outputs[2388] = ~(inputs[921]);
    assign layer0_outputs[2389] = inputs[1009];
    assign layer0_outputs[2390] = ~(inputs[173]);
    assign layer0_outputs[2391] = (inputs[694]) | (inputs[733]);
    assign layer0_outputs[2392] = ~(inputs[191]) | (inputs[356]);
    assign layer0_outputs[2393] = inputs[292];
    assign layer0_outputs[2394] = ~(inputs[858]) | (inputs[822]);
    assign layer0_outputs[2395] = (inputs[181]) & ~(inputs[164]);
    assign layer0_outputs[2396] = ~((inputs[993]) | (inputs[620]));
    assign layer0_outputs[2397] = 1'b1;
    assign layer0_outputs[2398] = (inputs[144]) | (inputs[1015]);
    assign layer0_outputs[2399] = inputs[409];
    assign layer0_outputs[2400] = ~((inputs[573]) & (inputs[952]));
    assign layer0_outputs[2401] = (inputs[653]) | (inputs[180]);
    assign layer0_outputs[2402] = inputs[57];
    assign layer0_outputs[2403] = ~((inputs[819]) | (inputs[866]));
    assign layer0_outputs[2404] = ~((inputs[336]) ^ (inputs[96]));
    assign layer0_outputs[2405] = ~((inputs[90]) | (inputs[871]));
    assign layer0_outputs[2406] = ~(inputs[253]) | (inputs[638]);
    assign layer0_outputs[2407] = ~(inputs[346]);
    assign layer0_outputs[2408] = (inputs[399]) & (inputs[106]);
    assign layer0_outputs[2409] = inputs[563];
    assign layer0_outputs[2410] = ~((inputs[401]) | (inputs[732]));
    assign layer0_outputs[2411] = ~(inputs[659]) | (inputs[782]);
    assign layer0_outputs[2412] = (inputs[827]) & ~(inputs[301]);
    assign layer0_outputs[2413] = (inputs[360]) ^ (inputs[385]);
    assign layer0_outputs[2414] = (inputs[796]) | (inputs[528]);
    assign layer0_outputs[2415] = inputs[379];
    assign layer0_outputs[2416] = (inputs[718]) | (inputs[381]);
    assign layer0_outputs[2417] = ~(inputs[486]) | (inputs[601]);
    assign layer0_outputs[2418] = ~((inputs[410]) | (inputs[175]));
    assign layer0_outputs[2419] = (inputs[142]) & ~(inputs[844]);
    assign layer0_outputs[2420] = ~(inputs[135]) | (inputs[585]);
    assign layer0_outputs[2421] = (inputs[302]) & ~(inputs[737]);
    assign layer0_outputs[2422] = (inputs[110]) | (inputs[436]);
    assign layer0_outputs[2423] = 1'b0;
    assign layer0_outputs[2424] = (inputs[64]) & (inputs[7]);
    assign layer0_outputs[2425] = ~(inputs[87]) | (inputs[669]);
    assign layer0_outputs[2426] = ~((inputs[903]) | (inputs[316]));
    assign layer0_outputs[2427] = ~(inputs[333]);
    assign layer0_outputs[2428] = (inputs[54]) & ~(inputs[327]);
    assign layer0_outputs[2429] = ~((inputs[116]) & (inputs[249]));
    assign layer0_outputs[2430] = ~(inputs[675]) | (inputs[199]);
    assign layer0_outputs[2431] = ~(inputs[20]);
    assign layer0_outputs[2432] = (inputs[386]) ^ (inputs[866]);
    assign layer0_outputs[2433] = ~((inputs[205]) & (inputs[191]));
    assign layer0_outputs[2434] = ~(inputs[533]) | (inputs[585]);
    assign layer0_outputs[2435] = ~(inputs[897]) | (inputs[785]);
    assign layer0_outputs[2436] = ~(inputs[309]);
    assign layer0_outputs[2437] = (inputs[401]) & ~(inputs[235]);
    assign layer0_outputs[2438] = inputs[38];
    assign layer0_outputs[2439] = ~(inputs[115]);
    assign layer0_outputs[2440] = (inputs[422]) | (inputs[426]);
    assign layer0_outputs[2441] = ~(inputs[691]) | (inputs[1022]);
    assign layer0_outputs[2442] = ~((inputs[714]) | (inputs[85]));
    assign layer0_outputs[2443] = inputs[954];
    assign layer0_outputs[2444] = inputs[48];
    assign layer0_outputs[2445] = ~(inputs[458]) | (inputs[951]);
    assign layer0_outputs[2446] = 1'b0;
    assign layer0_outputs[2447] = ~((inputs[600]) | (inputs[409]));
    assign layer0_outputs[2448] = (inputs[917]) | (inputs[324]);
    assign layer0_outputs[2449] = inputs[568];
    assign layer0_outputs[2450] = ~(inputs[891]) | (inputs[918]);
    assign layer0_outputs[2451] = inputs[148];
    assign layer0_outputs[2452] = (inputs[862]) & ~(inputs[342]);
    assign layer0_outputs[2453] = 1'b1;
    assign layer0_outputs[2454] = inputs[150];
    assign layer0_outputs[2455] = ~(inputs[563]);
    assign layer0_outputs[2456] = ~(inputs[63]);
    assign layer0_outputs[2457] = inputs[1011];
    assign layer0_outputs[2458] = ~(inputs[956]) | (inputs[986]);
    assign layer0_outputs[2459] = (inputs[664]) & (inputs[112]);
    assign layer0_outputs[2460] = (inputs[189]) | (inputs[517]);
    assign layer0_outputs[2461] = ~(inputs[184]);
    assign layer0_outputs[2462] = ~((inputs[416]) & (inputs[849]));
    assign layer0_outputs[2463] = ~(inputs[145]);
    assign layer0_outputs[2464] = inputs[285];
    assign layer0_outputs[2465] = (inputs[423]) ^ (inputs[1020]);
    assign layer0_outputs[2466] = (inputs[852]) & ~(inputs[759]);
    assign layer0_outputs[2467] = ~((inputs[878]) ^ (inputs[158]));
    assign layer0_outputs[2468] = ~(inputs[314]);
    assign layer0_outputs[2469] = ~((inputs[730]) | (inputs[625]));
    assign layer0_outputs[2470] = (inputs[58]) & (inputs[67]);
    assign layer0_outputs[2471] = ~(inputs[574]);
    assign layer0_outputs[2472] = (inputs[744]) & ~(inputs[119]);
    assign layer0_outputs[2473] = ~(inputs[999]) | (inputs[487]);
    assign layer0_outputs[2474] = ~((inputs[770]) ^ (inputs[348]));
    assign layer0_outputs[2475] = ~((inputs[920]) & (inputs[490]));
    assign layer0_outputs[2476] = ~(inputs[615]) | (inputs[94]);
    assign layer0_outputs[2477] = ~(inputs[371]) | (inputs[413]);
    assign layer0_outputs[2478] = ~(inputs[878]);
    assign layer0_outputs[2479] = inputs[487];
    assign layer0_outputs[2480] = ~((inputs[467]) ^ (inputs[769]));
    assign layer0_outputs[2481] = (inputs[296]) ^ (inputs[418]);
    assign layer0_outputs[2482] = ~((inputs[529]) & (inputs[962]));
    assign layer0_outputs[2483] = ~((inputs[346]) | (inputs[716]));
    assign layer0_outputs[2484] = ~(inputs[987]) | (inputs[709]);
    assign layer0_outputs[2485] = ~((inputs[427]) ^ (inputs[46]));
    assign layer0_outputs[2486] = ~((inputs[213]) & (inputs[854]));
    assign layer0_outputs[2487] = ~(inputs[199]) | (inputs[485]);
    assign layer0_outputs[2488] = ~((inputs[496]) ^ (inputs[1]));
    assign layer0_outputs[2489] = (inputs[507]) & (inputs[709]);
    assign layer0_outputs[2490] = ~((inputs[390]) | (inputs[791]));
    assign layer0_outputs[2491] = (inputs[874]) & ~(inputs[447]);
    assign layer0_outputs[2492] = (inputs[629]) ^ (inputs[343]);
    assign layer0_outputs[2493] = ~(inputs[519]);
    assign layer0_outputs[2494] = 1'b0;
    assign layer0_outputs[2495] = (inputs[775]) ^ (inputs[990]);
    assign layer0_outputs[2496] = ~(inputs[8]) | (inputs[250]);
    assign layer0_outputs[2497] = ~(inputs[727]);
    assign layer0_outputs[2498] = ~(inputs[859]);
    assign layer0_outputs[2499] = (inputs[176]) | (inputs[777]);
    assign layer0_outputs[2500] = (inputs[365]) | (inputs[659]);
    assign layer0_outputs[2501] = ~(inputs[366]) | (inputs[955]);
    assign layer0_outputs[2502] = ~((inputs[153]) | (inputs[692]));
    assign layer0_outputs[2503] = 1'b1;
    assign layer0_outputs[2504] = ~((inputs[365]) | (inputs[384]));
    assign layer0_outputs[2505] = (inputs[855]) | (inputs[760]);
    assign layer0_outputs[2506] = (inputs[744]) ^ (inputs[65]);
    assign layer0_outputs[2507] = ~(inputs[460]);
    assign layer0_outputs[2508] = (inputs[678]) & ~(inputs[758]);
    assign layer0_outputs[2509] = ~((inputs[345]) | (inputs[459]));
    assign layer0_outputs[2510] = ~((inputs[144]) | (inputs[837]));
    assign layer0_outputs[2511] = (inputs[522]) | (inputs[537]);
    assign layer0_outputs[2512] = ~(inputs[953]) | (inputs[302]);
    assign layer0_outputs[2513] = ~(inputs[248]);
    assign layer0_outputs[2514] = inputs[320];
    assign layer0_outputs[2515] = ~(inputs[38]);
    assign layer0_outputs[2516] = (inputs[631]) ^ (inputs[10]);
    assign layer0_outputs[2517] = (inputs[699]) & (inputs[425]);
    assign layer0_outputs[2518] = ~((inputs[948]) | (inputs[335]));
    assign layer0_outputs[2519] = 1'b0;
    assign layer0_outputs[2520] = 1'b0;
    assign layer0_outputs[2521] = inputs[552];
    assign layer0_outputs[2522] = ~(inputs[41]) | (inputs[896]);
    assign layer0_outputs[2523] = 1'b0;
    assign layer0_outputs[2524] = ~(inputs[6]);
    assign layer0_outputs[2525] = ~((inputs[575]) | (inputs[141]));
    assign layer0_outputs[2526] = ~(inputs[931]) | (inputs[231]);
    assign layer0_outputs[2527] = (inputs[382]) | (inputs[741]);
    assign layer0_outputs[2528] = (inputs[530]) | (inputs[977]);
    assign layer0_outputs[2529] = 1'b0;
    assign layer0_outputs[2530] = ~(inputs[845]);
    assign layer0_outputs[2531] = ~(inputs[179]) | (inputs[307]);
    assign layer0_outputs[2532] = inputs[774];
    assign layer0_outputs[2533] = inputs[658];
    assign layer0_outputs[2534] = ~(inputs[877]);
    assign layer0_outputs[2535] = inputs[22];
    assign layer0_outputs[2536] = ~(inputs[823]) | (inputs[506]);
    assign layer0_outputs[2537] = (inputs[150]) | (inputs[194]);
    assign layer0_outputs[2538] = ~((inputs[115]) & (inputs[356]));
    assign layer0_outputs[2539] = ~(inputs[145]);
    assign layer0_outputs[2540] = (inputs[820]) & ~(inputs[648]);
    assign layer0_outputs[2541] = (inputs[333]) | (inputs[103]);
    assign layer0_outputs[2542] = (inputs[39]) & ~(inputs[818]);
    assign layer0_outputs[2543] = 1'b1;
    assign layer0_outputs[2544] = 1'b1;
    assign layer0_outputs[2545] = ~((inputs[683]) | (inputs[882]));
    assign layer0_outputs[2546] = 1'b0;
    assign layer0_outputs[2547] = ~(inputs[936]) | (inputs[958]);
    assign layer0_outputs[2548] = 1'b1;
    assign layer0_outputs[2549] = (inputs[736]) | (inputs[110]);
    assign layer0_outputs[2550] = ~(inputs[303]);
    assign layer0_outputs[2551] = (inputs[994]) | (inputs[323]);
    assign layer0_outputs[2552] = ~(inputs[525]);
    assign layer0_outputs[2553] = ~((inputs[399]) & (inputs[771]));
    assign layer0_outputs[2554] = inputs[940];
    assign layer0_outputs[2555] = ~(inputs[640]);
    assign layer0_outputs[2556] = (inputs[52]) & (inputs[92]);
    assign layer0_outputs[2557] = (inputs[449]) | (inputs[30]);
    assign layer0_outputs[2558] = 1'b0;
    assign layer0_outputs[2559] = (inputs[519]) | (inputs[816]);
    assign layer1_outputs[0] = (layer0_outputs[624]) & ~(layer0_outputs[658]);
    assign layer1_outputs[1] = ~((layer0_outputs[575]) | (layer0_outputs[1988]));
    assign layer1_outputs[2] = ~((layer0_outputs[2315]) | (layer0_outputs[1828]));
    assign layer1_outputs[3] = ~(layer0_outputs[660]);
    assign layer1_outputs[4] = (layer0_outputs[775]) & (layer0_outputs[2211]);
    assign layer1_outputs[5] = 1'b0;
    assign layer1_outputs[6] = ~(layer0_outputs[35]);
    assign layer1_outputs[7] = (layer0_outputs[1685]) ^ (layer0_outputs[1335]);
    assign layer1_outputs[8] = (layer0_outputs[2144]) & ~(layer0_outputs[1807]);
    assign layer1_outputs[9] = ~((layer0_outputs[90]) | (layer0_outputs[736]));
    assign layer1_outputs[10] = ~(layer0_outputs[809]);
    assign layer1_outputs[11] = (layer0_outputs[626]) & ~(layer0_outputs[1391]);
    assign layer1_outputs[12] = ~(layer0_outputs[1985]);
    assign layer1_outputs[13] = layer0_outputs[1027];
    assign layer1_outputs[14] = ~((layer0_outputs[1945]) & (layer0_outputs[264]));
    assign layer1_outputs[15] = ~(layer0_outputs[1312]);
    assign layer1_outputs[16] = (layer0_outputs[1170]) ^ (layer0_outputs[1908]);
    assign layer1_outputs[17] = (layer0_outputs[1290]) | (layer0_outputs[178]);
    assign layer1_outputs[18] = (layer0_outputs[55]) & ~(layer0_outputs[665]);
    assign layer1_outputs[19] = ~(layer0_outputs[2042]);
    assign layer1_outputs[20] = ~(layer0_outputs[1838]);
    assign layer1_outputs[21] = ~(layer0_outputs[125]);
    assign layer1_outputs[22] = ~(layer0_outputs[322]) | (layer0_outputs[138]);
    assign layer1_outputs[23] = (layer0_outputs[567]) | (layer0_outputs[1205]);
    assign layer1_outputs[24] = layer0_outputs[1778];
    assign layer1_outputs[25] = (layer0_outputs[1578]) & (layer0_outputs[1392]);
    assign layer1_outputs[26] = layer0_outputs[1914];
    assign layer1_outputs[27] = layer0_outputs[2340];
    assign layer1_outputs[28] = (layer0_outputs[239]) & (layer0_outputs[624]);
    assign layer1_outputs[29] = ~(layer0_outputs[1997]);
    assign layer1_outputs[30] = (layer0_outputs[255]) & (layer0_outputs[122]);
    assign layer1_outputs[31] = layer0_outputs[1779];
    assign layer1_outputs[32] = ~((layer0_outputs[422]) | (layer0_outputs[1262]));
    assign layer1_outputs[33] = 1'b1;
    assign layer1_outputs[34] = 1'b1;
    assign layer1_outputs[35] = ~(layer0_outputs[684]);
    assign layer1_outputs[36] = (layer0_outputs[2074]) & ~(layer0_outputs[384]);
    assign layer1_outputs[37] = ~(layer0_outputs[2243]);
    assign layer1_outputs[38] = ~(layer0_outputs[172]) | (layer0_outputs[249]);
    assign layer1_outputs[39] = 1'b1;
    assign layer1_outputs[40] = ~(layer0_outputs[491]);
    assign layer1_outputs[41] = (layer0_outputs[2178]) & ~(layer0_outputs[543]);
    assign layer1_outputs[42] = 1'b1;
    assign layer1_outputs[43] = ~((layer0_outputs[2524]) | (layer0_outputs[2284]));
    assign layer1_outputs[44] = ~((layer0_outputs[930]) | (layer0_outputs[821]));
    assign layer1_outputs[45] = (layer0_outputs[212]) | (layer0_outputs[943]);
    assign layer1_outputs[46] = (layer0_outputs[1413]) & ~(layer0_outputs[1996]);
    assign layer1_outputs[47] = layer0_outputs[1180];
    assign layer1_outputs[48] = layer0_outputs[2198];
    assign layer1_outputs[49] = layer0_outputs[830];
    assign layer1_outputs[50] = (layer0_outputs[2378]) & (layer0_outputs[24]);
    assign layer1_outputs[51] = layer0_outputs[1816];
    assign layer1_outputs[52] = (layer0_outputs[436]) & (layer0_outputs[2165]);
    assign layer1_outputs[53] = ~(layer0_outputs[1727]) | (layer0_outputs[826]);
    assign layer1_outputs[54] = ~(layer0_outputs[995]);
    assign layer1_outputs[55] = layer0_outputs[457];
    assign layer1_outputs[56] = layer0_outputs[240];
    assign layer1_outputs[57] = (layer0_outputs[1464]) ^ (layer0_outputs[1913]);
    assign layer1_outputs[58] = (layer0_outputs[1280]) & ~(layer0_outputs[463]);
    assign layer1_outputs[59] = (layer0_outputs[672]) & ~(layer0_outputs[2006]);
    assign layer1_outputs[60] = ~(layer0_outputs[2421]);
    assign layer1_outputs[61] = layer0_outputs[1105];
    assign layer1_outputs[62] = 1'b0;
    assign layer1_outputs[63] = ~(layer0_outputs[501]) | (layer0_outputs[699]);
    assign layer1_outputs[64] = 1'b0;
    assign layer1_outputs[65] = layer0_outputs[762];
    assign layer1_outputs[66] = (layer0_outputs[1775]) & ~(layer0_outputs[1617]);
    assign layer1_outputs[67] = 1'b0;
    assign layer1_outputs[68] = layer0_outputs[2349];
    assign layer1_outputs[69] = ~(layer0_outputs[1257]) | (layer0_outputs[2141]);
    assign layer1_outputs[70] = ~(layer0_outputs[2013]) | (layer0_outputs[1044]);
    assign layer1_outputs[71] = ~(layer0_outputs[1625]);
    assign layer1_outputs[72] = (layer0_outputs[1152]) & ~(layer0_outputs[1984]);
    assign layer1_outputs[73] = ~(layer0_outputs[2048]);
    assign layer1_outputs[74] = 1'b1;
    assign layer1_outputs[75] = ~(layer0_outputs[1836]);
    assign layer1_outputs[76] = (layer0_outputs[2164]) | (layer0_outputs[142]);
    assign layer1_outputs[77] = layer0_outputs[1694];
    assign layer1_outputs[78] = layer0_outputs[2177];
    assign layer1_outputs[79] = 1'b1;
    assign layer1_outputs[80] = layer0_outputs[429];
    assign layer1_outputs[81] = ~(layer0_outputs[876]);
    assign layer1_outputs[82] = ~(layer0_outputs[578]) | (layer0_outputs[1760]);
    assign layer1_outputs[83] = (layer0_outputs[730]) & ~(layer0_outputs[843]);
    assign layer1_outputs[84] = layer0_outputs[1587];
    assign layer1_outputs[85] = ~((layer0_outputs[1349]) ^ (layer0_outputs[927]));
    assign layer1_outputs[86] = ~((layer0_outputs[1407]) | (layer0_outputs[2269]));
    assign layer1_outputs[87] = (layer0_outputs[706]) & ~(layer0_outputs[1915]);
    assign layer1_outputs[88] = (layer0_outputs[310]) & ~(layer0_outputs[168]);
    assign layer1_outputs[89] = (layer0_outputs[423]) ^ (layer0_outputs[1510]);
    assign layer1_outputs[90] = 1'b1;
    assign layer1_outputs[91] = (layer0_outputs[1413]) & (layer0_outputs[211]);
    assign layer1_outputs[92] = (layer0_outputs[1925]) | (layer0_outputs[2160]);
    assign layer1_outputs[93] = ~(layer0_outputs[1151]);
    assign layer1_outputs[94] = (layer0_outputs[754]) & ~(layer0_outputs[609]);
    assign layer1_outputs[95] = 1'b1;
    assign layer1_outputs[96] = ~((layer0_outputs[2272]) | (layer0_outputs[555]));
    assign layer1_outputs[97] = ~(layer0_outputs[2208]) | (layer0_outputs[693]);
    assign layer1_outputs[98] = 1'b1;
    assign layer1_outputs[99] = ~(layer0_outputs[157]);
    assign layer1_outputs[100] = layer0_outputs[9];
    assign layer1_outputs[101] = ~(layer0_outputs[439]) | (layer0_outputs[1272]);
    assign layer1_outputs[102] = layer0_outputs[592];
    assign layer1_outputs[103] = ~(layer0_outputs[1242]) | (layer0_outputs[2029]);
    assign layer1_outputs[104] = (layer0_outputs[1053]) & ~(layer0_outputs[1284]);
    assign layer1_outputs[105] = (layer0_outputs[2150]) & ~(layer0_outputs[2456]);
    assign layer1_outputs[106] = 1'b1;
    assign layer1_outputs[107] = 1'b1;
    assign layer1_outputs[108] = (layer0_outputs[2268]) & (layer0_outputs[1397]);
    assign layer1_outputs[109] = 1'b1;
    assign layer1_outputs[110] = (layer0_outputs[505]) & ~(layer0_outputs[1252]);
    assign layer1_outputs[111] = (layer0_outputs[622]) & ~(layer0_outputs[1971]);
    assign layer1_outputs[112] = layer0_outputs[2102];
    assign layer1_outputs[113] = ~(layer0_outputs[2145]);
    assign layer1_outputs[114] = (layer0_outputs[931]) | (layer0_outputs[1007]);
    assign layer1_outputs[115] = layer0_outputs[2513];
    assign layer1_outputs[116] = (layer0_outputs[1559]) & ~(layer0_outputs[273]);
    assign layer1_outputs[117] = ~(layer0_outputs[323]);
    assign layer1_outputs[118] = ~((layer0_outputs[738]) & (layer0_outputs[1958]));
    assign layer1_outputs[119] = ~((layer0_outputs[1631]) | (layer0_outputs[41]));
    assign layer1_outputs[120] = layer0_outputs[1632];
    assign layer1_outputs[121] = 1'b0;
    assign layer1_outputs[122] = 1'b1;
    assign layer1_outputs[123] = ~(layer0_outputs[1646]) | (layer0_outputs[2101]);
    assign layer1_outputs[124] = layer0_outputs[2504];
    assign layer1_outputs[125] = (layer0_outputs[555]) & ~(layer0_outputs[335]);
    assign layer1_outputs[126] = layer0_outputs[465];
    assign layer1_outputs[127] = ~(layer0_outputs[1787]);
    assign layer1_outputs[128] = (layer0_outputs[567]) | (layer0_outputs[1519]);
    assign layer1_outputs[129] = layer0_outputs[1705];
    assign layer1_outputs[130] = layer0_outputs[519];
    assign layer1_outputs[131] = (layer0_outputs[2264]) & (layer0_outputs[1764]);
    assign layer1_outputs[132] = (layer0_outputs[7]) & ~(layer0_outputs[1942]);
    assign layer1_outputs[133] = (layer0_outputs[1315]) & ~(layer0_outputs[1224]);
    assign layer1_outputs[134] = layer0_outputs[247];
    assign layer1_outputs[135] = ~(layer0_outputs[1375]);
    assign layer1_outputs[136] = ~(layer0_outputs[263]);
    assign layer1_outputs[137] = ~(layer0_outputs[1885]) | (layer0_outputs[800]);
    assign layer1_outputs[138] = layer0_outputs[215];
    assign layer1_outputs[139] = ~(layer0_outputs[1494]) | (layer0_outputs[1912]);
    assign layer1_outputs[140] = 1'b0;
    assign layer1_outputs[141] = ~((layer0_outputs[178]) | (layer0_outputs[2313]));
    assign layer1_outputs[142] = 1'b1;
    assign layer1_outputs[143] = (layer0_outputs[594]) & (layer0_outputs[737]);
    assign layer1_outputs[144] = 1'b1;
    assign layer1_outputs[145] = ~(layer0_outputs[107]) | (layer0_outputs[1959]);
    assign layer1_outputs[146] = ~((layer0_outputs[2155]) | (layer0_outputs[875]));
    assign layer1_outputs[147] = layer0_outputs[1060];
    assign layer1_outputs[148] = ~((layer0_outputs[442]) & (layer0_outputs[2493]));
    assign layer1_outputs[149] = (layer0_outputs[466]) & ~(layer0_outputs[2036]);
    assign layer1_outputs[150] = ~(layer0_outputs[2387]) | (layer0_outputs[825]);
    assign layer1_outputs[151] = (layer0_outputs[548]) & ~(layer0_outputs[437]);
    assign layer1_outputs[152] = ~(layer0_outputs[1653]) | (layer0_outputs[510]);
    assign layer1_outputs[153] = (layer0_outputs[33]) & ~(layer0_outputs[261]);
    assign layer1_outputs[154] = ~(layer0_outputs[1889]);
    assign layer1_outputs[155] = ~(layer0_outputs[123]);
    assign layer1_outputs[156] = ~((layer0_outputs[235]) & (layer0_outputs[2087]));
    assign layer1_outputs[157] = (layer0_outputs[1897]) & ~(layer0_outputs[939]);
    assign layer1_outputs[158] = layer0_outputs[1858];
    assign layer1_outputs[159] = ~((layer0_outputs[1723]) | (layer0_outputs[198]));
    assign layer1_outputs[160] = ~(layer0_outputs[2075]) | (layer0_outputs[192]);
    assign layer1_outputs[161] = 1'b1;
    assign layer1_outputs[162] = ~(layer0_outputs[357]) | (layer0_outputs[785]);
    assign layer1_outputs[163] = 1'b1;
    assign layer1_outputs[164] = ~(layer0_outputs[2353]) | (layer0_outputs[772]);
    assign layer1_outputs[165] = ~(layer0_outputs[1429]) | (layer0_outputs[697]);
    assign layer1_outputs[166] = (layer0_outputs[1999]) & ~(layer0_outputs[213]);
    assign layer1_outputs[167] = ~(layer0_outputs[179]);
    assign layer1_outputs[168] = ~(layer0_outputs[2485]) | (layer0_outputs[1047]);
    assign layer1_outputs[169] = (layer0_outputs[1059]) | (layer0_outputs[2229]);
    assign layer1_outputs[170] = ~((layer0_outputs[525]) | (layer0_outputs[1410]));
    assign layer1_outputs[171] = layer0_outputs[1711];
    assign layer1_outputs[172] = layer0_outputs[93];
    assign layer1_outputs[173] = ~(layer0_outputs[370]) | (layer0_outputs[1073]);
    assign layer1_outputs[174] = ~(layer0_outputs[2293]);
    assign layer1_outputs[175] = ~(layer0_outputs[1163]);
    assign layer1_outputs[176] = (layer0_outputs[2543]) & ~(layer0_outputs[52]);
    assign layer1_outputs[177] = ~((layer0_outputs[1759]) | (layer0_outputs[1983]));
    assign layer1_outputs[178] = layer0_outputs[2310];
    assign layer1_outputs[179] = layer0_outputs[732];
    assign layer1_outputs[180] = (layer0_outputs[27]) | (layer0_outputs[2539]);
    assign layer1_outputs[181] = layer0_outputs[1098];
    assign layer1_outputs[182] = 1'b0;
    assign layer1_outputs[183] = layer0_outputs[915];
    assign layer1_outputs[184] = (layer0_outputs[1166]) | (layer0_outputs[1956]);
    assign layer1_outputs[185] = ~((layer0_outputs[49]) | (layer0_outputs[1338]));
    assign layer1_outputs[186] = ~(layer0_outputs[1219]) | (layer0_outputs[985]);
    assign layer1_outputs[187] = ~(layer0_outputs[898]) | (layer0_outputs[1033]);
    assign layer1_outputs[188] = layer0_outputs[1531];
    assign layer1_outputs[189] = ~(layer0_outputs[1397]);
    assign layer1_outputs[190] = layer0_outputs[2374];
    assign layer1_outputs[191] = (layer0_outputs[1840]) & (layer0_outputs[1542]);
    assign layer1_outputs[192] = layer0_outputs[1320];
    assign layer1_outputs[193] = layer0_outputs[547];
    assign layer1_outputs[194] = layer0_outputs[38];
    assign layer1_outputs[195] = ~((layer0_outputs[357]) | (layer0_outputs[401]));
    assign layer1_outputs[196] = ~(layer0_outputs[1078]);
    assign layer1_outputs[197] = ~(layer0_outputs[51]);
    assign layer1_outputs[198] = (layer0_outputs[373]) | (layer0_outputs[627]);
    assign layer1_outputs[199] = (layer0_outputs[2267]) & ~(layer0_outputs[1334]);
    assign layer1_outputs[200] = ~((layer0_outputs[2322]) & (layer0_outputs[656]));
    assign layer1_outputs[201] = (layer0_outputs[2072]) | (layer0_outputs[1218]);
    assign layer1_outputs[202] = ~(layer0_outputs[2390]);
    assign layer1_outputs[203] = ~(layer0_outputs[1448]) | (layer0_outputs[126]);
    assign layer1_outputs[204] = (layer0_outputs[475]) & (layer0_outputs[1511]);
    assign layer1_outputs[205] = 1'b1;
    assign layer1_outputs[206] = ~((layer0_outputs[1793]) & (layer0_outputs[725]));
    assign layer1_outputs[207] = ~(layer0_outputs[2448]);
    assign layer1_outputs[208] = layer0_outputs[185];
    assign layer1_outputs[209] = layer0_outputs[2350];
    assign layer1_outputs[210] = 1'b1;
    assign layer1_outputs[211] = ~((layer0_outputs[483]) ^ (layer0_outputs[1661]));
    assign layer1_outputs[212] = ~(layer0_outputs[404]) | (layer0_outputs[1946]);
    assign layer1_outputs[213] = layer0_outputs[291];
    assign layer1_outputs[214] = ~((layer0_outputs[86]) & (layer0_outputs[1621]));
    assign layer1_outputs[215] = (layer0_outputs[2249]) & (layer0_outputs[2344]);
    assign layer1_outputs[216] = layer0_outputs[479];
    assign layer1_outputs[217] = 1'b0;
    assign layer1_outputs[218] = (layer0_outputs[954]) & ~(layer0_outputs[2343]);
    assign layer1_outputs[219] = ~(layer0_outputs[735]);
    assign layer1_outputs[220] = layer0_outputs[2297];
    assign layer1_outputs[221] = (layer0_outputs[2209]) ^ (layer0_outputs[933]);
    assign layer1_outputs[222] = ~(layer0_outputs[1773]);
    assign layer1_outputs[223] = layer0_outputs[1144];
    assign layer1_outputs[224] = ~(layer0_outputs[1158]) | (layer0_outputs[729]);
    assign layer1_outputs[225] = ~((layer0_outputs[2164]) & (layer0_outputs[1177]));
    assign layer1_outputs[226] = ~(layer0_outputs[1804]);
    assign layer1_outputs[227] = ~(layer0_outputs[85]);
    assign layer1_outputs[228] = 1'b1;
    assign layer1_outputs[229] = 1'b1;
    assign layer1_outputs[230] = (layer0_outputs[1713]) | (layer0_outputs[43]);
    assign layer1_outputs[231] = 1'b0;
    assign layer1_outputs[232] = ~((layer0_outputs[1598]) & (layer0_outputs[1991]));
    assign layer1_outputs[233] = (layer0_outputs[358]) & ~(layer0_outputs[41]);
    assign layer1_outputs[234] = layer0_outputs[2048];
    assign layer1_outputs[235] = ~(layer0_outputs[1238]) | (layer0_outputs[2262]);
    assign layer1_outputs[236] = 1'b1;
    assign layer1_outputs[237] = (layer0_outputs[2019]) & (layer0_outputs[1804]);
    assign layer1_outputs[238] = (layer0_outputs[1958]) | (layer0_outputs[1695]);
    assign layer1_outputs[239] = ~(layer0_outputs[2338]);
    assign layer1_outputs[240] = ~(layer0_outputs[570]) | (layer0_outputs[1689]);
    assign layer1_outputs[241] = 1'b1;
    assign layer1_outputs[242] = ~(layer0_outputs[1633]) | (layer0_outputs[325]);
    assign layer1_outputs[243] = ~(layer0_outputs[1217]);
    assign layer1_outputs[244] = ~(layer0_outputs[2166]) | (layer0_outputs[1745]);
    assign layer1_outputs[245] = ~((layer0_outputs[1346]) | (layer0_outputs[1900]));
    assign layer1_outputs[246] = ~((layer0_outputs[1582]) | (layer0_outputs[622]));
    assign layer1_outputs[247] = ~(layer0_outputs[1134]);
    assign layer1_outputs[248] = 1'b0;
    assign layer1_outputs[249] = layer0_outputs[983];
    assign layer1_outputs[250] = ~(layer0_outputs[2202]) | (layer0_outputs[2093]);
    assign layer1_outputs[251] = ~((layer0_outputs[841]) | (layer0_outputs[514]));
    assign layer1_outputs[252] = ~(layer0_outputs[1676]);
    assign layer1_outputs[253] = layer0_outputs[77];
    assign layer1_outputs[254] = 1'b1;
    assign layer1_outputs[255] = ~(layer0_outputs[242]) | (layer0_outputs[636]);
    assign layer1_outputs[256] = 1'b1;
    assign layer1_outputs[257] = ~((layer0_outputs[2009]) ^ (layer0_outputs[456]));
    assign layer1_outputs[258] = layer0_outputs[327];
    assign layer1_outputs[259] = (layer0_outputs[2037]) & (layer0_outputs[1029]);
    assign layer1_outputs[260] = (layer0_outputs[164]) ^ (layer0_outputs[2551]);
    assign layer1_outputs[261] = ~(layer0_outputs[409]);
    assign layer1_outputs[262] = ~(layer0_outputs[570]) | (layer0_outputs[2298]);
    assign layer1_outputs[263] = ~(layer0_outputs[2271]);
    assign layer1_outputs[264] = (layer0_outputs[1261]) | (layer0_outputs[620]);
    assign layer1_outputs[265] = ~((layer0_outputs[1375]) & (layer0_outputs[152]));
    assign layer1_outputs[266] = ~((layer0_outputs[197]) | (layer0_outputs[400]));
    assign layer1_outputs[267] = 1'b0;
    assign layer1_outputs[268] = layer0_outputs[1721];
    assign layer1_outputs[269] = ~(layer0_outputs[1253]) | (layer0_outputs[3]);
    assign layer1_outputs[270] = (layer0_outputs[342]) & ~(layer0_outputs[373]);
    assign layer1_outputs[271] = ~(layer0_outputs[1729]);
    assign layer1_outputs[272] = (layer0_outputs[1177]) & ~(layer0_outputs[648]);
    assign layer1_outputs[273] = layer0_outputs[2493];
    assign layer1_outputs[274] = ~(layer0_outputs[1324]) | (layer0_outputs[2091]);
    assign layer1_outputs[275] = (layer0_outputs[1510]) | (layer0_outputs[1788]);
    assign layer1_outputs[276] = (layer0_outputs[667]) & (layer0_outputs[1462]);
    assign layer1_outputs[277] = (layer0_outputs[1766]) & (layer0_outputs[269]);
    assign layer1_outputs[278] = (layer0_outputs[1915]) | (layer0_outputs[2090]);
    assign layer1_outputs[279] = ~(layer0_outputs[372]);
    assign layer1_outputs[280] = ~(layer0_outputs[2426]) | (layer0_outputs[482]);
    assign layer1_outputs[281] = 1'b1;
    assign layer1_outputs[282] = (layer0_outputs[192]) & (layer0_outputs[784]);
    assign layer1_outputs[283] = ~((layer0_outputs[839]) | (layer0_outputs[2129]));
    assign layer1_outputs[284] = (layer0_outputs[1977]) | (layer0_outputs[1034]);
    assign layer1_outputs[285] = (layer0_outputs[105]) | (layer0_outputs[175]);
    assign layer1_outputs[286] = ~((layer0_outputs[1109]) & (layer0_outputs[1481]));
    assign layer1_outputs[287] = ~(layer0_outputs[1865]);
    assign layer1_outputs[288] = ~(layer0_outputs[1415]) | (layer0_outputs[1371]);
    assign layer1_outputs[289] = 1'b1;
    assign layer1_outputs[290] = layer0_outputs[2476];
    assign layer1_outputs[291] = (layer0_outputs[705]) | (layer0_outputs[293]);
    assign layer1_outputs[292] = ~(layer0_outputs[1125]);
    assign layer1_outputs[293] = layer0_outputs[377];
    assign layer1_outputs[294] = ~(layer0_outputs[1740]);
    assign layer1_outputs[295] = (layer0_outputs[1878]) & (layer0_outputs[23]);
    assign layer1_outputs[296] = layer0_outputs[233];
    assign layer1_outputs[297] = ~((layer0_outputs[1658]) | (layer0_outputs[399]));
    assign layer1_outputs[298] = ~(layer0_outputs[2117]) | (layer0_outputs[532]);
    assign layer1_outputs[299] = ~(layer0_outputs[702]);
    assign layer1_outputs[300] = ~(layer0_outputs[378]) | (layer0_outputs[2535]);
    assign layer1_outputs[301] = layer0_outputs[2138];
    assign layer1_outputs[302] = 1'b1;
    assign layer1_outputs[303] = layer0_outputs[556];
    assign layer1_outputs[304] = (layer0_outputs[183]) & ~(layer0_outputs[492]);
    assign layer1_outputs[305] = ~(layer0_outputs[12]);
    assign layer1_outputs[306] = ~(layer0_outputs[2253]);
    assign layer1_outputs[307] = layer0_outputs[2234];
    assign layer1_outputs[308] = (layer0_outputs[1647]) & (layer0_outputs[1887]);
    assign layer1_outputs[309] = 1'b1;
    assign layer1_outputs[310] = 1'b1;
    assign layer1_outputs[311] = 1'b1;
    assign layer1_outputs[312] = ~((layer0_outputs[1871]) | (layer0_outputs[97]));
    assign layer1_outputs[313] = (layer0_outputs[657]) & (layer0_outputs[760]);
    assign layer1_outputs[314] = layer0_outputs[1493];
    assign layer1_outputs[315] = ~(layer0_outputs[1408]);
    assign layer1_outputs[316] = layer0_outputs[73];
    assign layer1_outputs[317] = (layer0_outputs[48]) & (layer0_outputs[633]);
    assign layer1_outputs[318] = 1'b1;
    assign layer1_outputs[319] = ~((layer0_outputs[1628]) | (layer0_outputs[2056]));
    assign layer1_outputs[320] = (layer0_outputs[308]) & (layer0_outputs[105]);
    assign layer1_outputs[321] = layer0_outputs[183];
    assign layer1_outputs[322] = 1'b1;
    assign layer1_outputs[323] = ~((layer0_outputs[1896]) | (layer0_outputs[583]));
    assign layer1_outputs[324] = ~(layer0_outputs[1424]);
    assign layer1_outputs[325] = layer0_outputs[2283];
    assign layer1_outputs[326] = (layer0_outputs[821]) | (layer0_outputs[2226]);
    assign layer1_outputs[327] = 1'b1;
    assign layer1_outputs[328] = (layer0_outputs[739]) | (layer0_outputs[1083]);
    assign layer1_outputs[329] = layer0_outputs[1978];
    assign layer1_outputs[330] = (layer0_outputs[238]) | (layer0_outputs[270]);
    assign layer1_outputs[331] = ~(layer0_outputs[295]);
    assign layer1_outputs[332] = 1'b0;
    assign layer1_outputs[333] = (layer0_outputs[466]) & ~(layer0_outputs[2245]);
    assign layer1_outputs[334] = ~((layer0_outputs[809]) | (layer0_outputs[1246]));
    assign layer1_outputs[335] = (layer0_outputs[1953]) & (layer0_outputs[1637]);
    assign layer1_outputs[336] = (layer0_outputs[1076]) & ~(layer0_outputs[1569]);
    assign layer1_outputs[337] = ~(layer0_outputs[421]) | (layer0_outputs[2336]);
    assign layer1_outputs[338] = ~(layer0_outputs[934]);
    assign layer1_outputs[339] = layer0_outputs[781];
    assign layer1_outputs[340] = ~(layer0_outputs[1871]);
    assign layer1_outputs[341] = layer0_outputs[207];
    assign layer1_outputs[342] = layer0_outputs[1169];
    assign layer1_outputs[343] = ~(layer0_outputs[312]);
    assign layer1_outputs[344] = ~(layer0_outputs[744]) | (layer0_outputs[253]);
    assign layer1_outputs[345] = (layer0_outputs[2220]) & ~(layer0_outputs[1095]);
    assign layer1_outputs[346] = (layer0_outputs[398]) & ~(layer0_outputs[1874]);
    assign layer1_outputs[347] = layer0_outputs[2485];
    assign layer1_outputs[348] = layer0_outputs[531];
    assign layer1_outputs[349] = ~(layer0_outputs[2003]);
    assign layer1_outputs[350] = ~(layer0_outputs[1976]) | (layer0_outputs[334]);
    assign layer1_outputs[351] = ~(layer0_outputs[2151]);
    assign layer1_outputs[352] = ~(layer0_outputs[367]);
    assign layer1_outputs[353] = ~((layer0_outputs[1387]) ^ (layer0_outputs[2543]));
    assign layer1_outputs[354] = (layer0_outputs[566]) & (layer0_outputs[2254]);
    assign layer1_outputs[355] = (layer0_outputs[799]) & ~(layer0_outputs[2275]);
    assign layer1_outputs[356] = (layer0_outputs[355]) & ~(layer0_outputs[2338]);
    assign layer1_outputs[357] = ~((layer0_outputs[80]) | (layer0_outputs[158]));
    assign layer1_outputs[358] = layer0_outputs[2067];
    assign layer1_outputs[359] = (layer0_outputs[941]) & (layer0_outputs[1984]);
    assign layer1_outputs[360] = (layer0_outputs[1473]) | (layer0_outputs[956]);
    assign layer1_outputs[361] = 1'b0;
    assign layer1_outputs[362] = (layer0_outputs[2023]) & ~(layer0_outputs[588]);
    assign layer1_outputs[363] = ~((layer0_outputs[2434]) & (layer0_outputs[1347]));
    assign layer1_outputs[364] = 1'b1;
    assign layer1_outputs[365] = layer0_outputs[2073];
    assign layer1_outputs[366] = (layer0_outputs[1624]) & ~(layer0_outputs[478]);
    assign layer1_outputs[367] = ~((layer0_outputs[743]) & (layer0_outputs[1484]));
    assign layer1_outputs[368] = 1'b1;
    assign layer1_outputs[369] = (layer0_outputs[1733]) & ~(layer0_outputs[26]);
    assign layer1_outputs[370] = layer0_outputs[1232];
    assign layer1_outputs[371] = (layer0_outputs[1856]) & ~(layer0_outputs[320]);
    assign layer1_outputs[372] = ~(layer0_outputs[923]) | (layer0_outputs[700]);
    assign layer1_outputs[373] = ~(layer0_outputs[1902]) | (layer0_outputs[621]);
    assign layer1_outputs[374] = 1'b0;
    assign layer1_outputs[375] = (layer0_outputs[1264]) | (layer0_outputs[1623]);
    assign layer1_outputs[376] = ~((layer0_outputs[2469]) & (layer0_outputs[153]));
    assign layer1_outputs[377] = ~((layer0_outputs[2066]) & (layer0_outputs[813]));
    assign layer1_outputs[378] = (layer0_outputs[250]) & ~(layer0_outputs[1111]);
    assign layer1_outputs[379] = ~(layer0_outputs[1648]);
    assign layer1_outputs[380] = layer0_outputs[252];
    assign layer1_outputs[381] = layer0_outputs[562];
    assign layer1_outputs[382] = ~(layer0_outputs[1128]);
    assign layer1_outputs[383] = (layer0_outputs[1967]) | (layer0_outputs[1724]);
    assign layer1_outputs[384] = ~(layer0_outputs[1559]) | (layer0_outputs[2187]);
    assign layer1_outputs[385] = ~((layer0_outputs[779]) & (layer0_outputs[251]));
    assign layer1_outputs[386] = ~(layer0_outputs[1917]);
    assign layer1_outputs[387] = ~(layer0_outputs[2300]) | (layer0_outputs[1862]);
    assign layer1_outputs[388] = ~(layer0_outputs[1719]);
    assign layer1_outputs[389] = ~(layer0_outputs[2324]) | (layer0_outputs[1727]);
    assign layer1_outputs[390] = layer0_outputs[1964];
    assign layer1_outputs[391] = (layer0_outputs[1417]) | (layer0_outputs[2000]);
    assign layer1_outputs[392] = (layer0_outputs[387]) ^ (layer0_outputs[1905]);
    assign layer1_outputs[393] = ~(layer0_outputs[2028]);
    assign layer1_outputs[394] = ~((layer0_outputs[861]) | (layer0_outputs[2532]));
    assign layer1_outputs[395] = ~(layer0_outputs[2047]) | (layer0_outputs[2414]);
    assign layer1_outputs[396] = ~(layer0_outputs[49]) | (layer0_outputs[545]);
    assign layer1_outputs[397] = 1'b0;
    assign layer1_outputs[398] = layer0_outputs[2244];
    assign layer1_outputs[399] = ~((layer0_outputs[476]) | (layer0_outputs[2292]));
    assign layer1_outputs[400] = (layer0_outputs[2089]) & ~(layer0_outputs[1739]);
    assign layer1_outputs[401] = ~(layer0_outputs[1322]) | (layer0_outputs[1042]);
    assign layer1_outputs[402] = ~(layer0_outputs[1225]);
    assign layer1_outputs[403] = (layer0_outputs[773]) & ~(layer0_outputs[889]);
    assign layer1_outputs[404] = layer0_outputs[132];
    assign layer1_outputs[405] = (layer0_outputs[1107]) & ~(layer0_outputs[651]);
    assign layer1_outputs[406] = (layer0_outputs[753]) & (layer0_outputs[2061]);
    assign layer1_outputs[407] = ~((layer0_outputs[1149]) | (layer0_outputs[1270]));
    assign layer1_outputs[408] = ~((layer0_outputs[1164]) ^ (layer0_outputs[2003]));
    assign layer1_outputs[409] = layer0_outputs[191];
    assign layer1_outputs[410] = ~((layer0_outputs[1599]) & (layer0_outputs[640]));
    assign layer1_outputs[411] = layer0_outputs[1551];
    assign layer1_outputs[412] = layer0_outputs[966];
    assign layer1_outputs[413] = layer0_outputs[2276];
    assign layer1_outputs[414] = (layer0_outputs[483]) | (layer0_outputs[2352]);
    assign layer1_outputs[415] = ~(layer0_outputs[575]);
    assign layer1_outputs[416] = ~(layer0_outputs[189]);
    assign layer1_outputs[417] = layer0_outputs[2516];
    assign layer1_outputs[418] = (layer0_outputs[1075]) & ~(layer0_outputs[608]);
    assign layer1_outputs[419] = ~(layer0_outputs[1411]);
    assign layer1_outputs[420] = 1'b0;
    assign layer1_outputs[421] = ~(layer0_outputs[1326]);
    assign layer1_outputs[422] = layer0_outputs[928];
    assign layer1_outputs[423] = (layer0_outputs[2060]) & ~(layer0_outputs[1405]);
    assign layer1_outputs[424] = 1'b1;
    assign layer1_outputs[425] = layer0_outputs[113];
    assign layer1_outputs[426] = ~(layer0_outputs[303]) | (layer0_outputs[2149]);
    assign layer1_outputs[427] = ~((layer0_outputs[485]) & (layer0_outputs[306]));
    assign layer1_outputs[428] = ~((layer0_outputs[1651]) & (layer0_outputs[1811]));
    assign layer1_outputs[429] = (layer0_outputs[874]) & ~(layer0_outputs[198]);
    assign layer1_outputs[430] = ~(layer0_outputs[1145]) | (layer0_outputs[964]);
    assign layer1_outputs[431] = (layer0_outputs[697]) & ~(layer0_outputs[2529]);
    assign layer1_outputs[432] = ~(layer0_outputs[968]);
    assign layer1_outputs[433] = ~(layer0_outputs[213]);
    assign layer1_outputs[434] = ~((layer0_outputs[325]) | (layer0_outputs[1358]));
    assign layer1_outputs[435] = 1'b1;
    assign layer1_outputs[436] = ~(layer0_outputs[81]);
    assign layer1_outputs[437] = ~((layer0_outputs[714]) & (layer0_outputs[2293]));
    assign layer1_outputs[438] = ~(layer0_outputs[1186]);
    assign layer1_outputs[439] = layer0_outputs[1366];
    assign layer1_outputs[440] = ~(layer0_outputs[1006]);
    assign layer1_outputs[441] = ~(layer0_outputs[2093]) | (layer0_outputs[2369]);
    assign layer1_outputs[442] = ~(layer0_outputs[1049]) | (layer0_outputs[837]);
    assign layer1_outputs[443] = ~(layer0_outputs[1368]) | (layer0_outputs[659]);
    assign layer1_outputs[444] = layer0_outputs[1970];
    assign layer1_outputs[445] = ~((layer0_outputs[114]) ^ (layer0_outputs[517]));
    assign layer1_outputs[446] = ~(layer0_outputs[2463]);
    assign layer1_outputs[447] = (layer0_outputs[1168]) & ~(layer0_outputs[203]);
    assign layer1_outputs[448] = layer0_outputs[1908];
    assign layer1_outputs[449] = ~(layer0_outputs[2556]) | (layer0_outputs[1077]);
    assign layer1_outputs[450] = layer0_outputs[2379];
    assign layer1_outputs[451] = (layer0_outputs[224]) ^ (layer0_outputs[1448]);
    assign layer1_outputs[452] = (layer0_outputs[2359]) | (layer0_outputs[1250]);
    assign layer1_outputs[453] = (layer0_outputs[308]) & ~(layer0_outputs[777]);
    assign layer1_outputs[454] = layer0_outputs[668];
    assign layer1_outputs[455] = 1'b1;
    assign layer1_outputs[456] = ~(layer0_outputs[479]);
    assign layer1_outputs[457] = layer0_outputs[1744];
    assign layer1_outputs[458] = layer0_outputs[2217];
    assign layer1_outputs[459] = ~(layer0_outputs[1644]) | (layer0_outputs[508]);
    assign layer1_outputs[460] = 1'b0;
    assign layer1_outputs[461] = ~(layer0_outputs[2527]);
    assign layer1_outputs[462] = ~(layer0_outputs[76]);
    assign layer1_outputs[463] = layer0_outputs[2309];
    assign layer1_outputs[464] = ~((layer0_outputs[1636]) | (layer0_outputs[2430]));
    assign layer1_outputs[465] = 1'b0;
    assign layer1_outputs[466] = layer0_outputs[1218];
    assign layer1_outputs[467] = ~((layer0_outputs[830]) & (layer0_outputs[2546]));
    assign layer1_outputs[468] = ~(layer0_outputs[360]) | (layer0_outputs[1911]);
    assign layer1_outputs[469] = ~((layer0_outputs[2163]) & (layer0_outputs[2222]));
    assign layer1_outputs[470] = layer0_outputs[1683];
    assign layer1_outputs[471] = ~(layer0_outputs[474]) | (layer0_outputs[562]);
    assign layer1_outputs[472] = (layer0_outputs[1602]) & (layer0_outputs[689]);
    assign layer1_outputs[473] = ~((layer0_outputs[1455]) | (layer0_outputs[2297]));
    assign layer1_outputs[474] = layer0_outputs[1586];
    assign layer1_outputs[475] = 1'b1;
    assign layer1_outputs[476] = ~((layer0_outputs[1099]) | (layer0_outputs[551]));
    assign layer1_outputs[477] = ~(layer0_outputs[2240]) | (layer0_outputs[942]);
    assign layer1_outputs[478] = (layer0_outputs[354]) & (layer0_outputs[683]);
    assign layer1_outputs[479] = layer0_outputs[491];
    assign layer1_outputs[480] = ~((layer0_outputs[2464]) & (layer0_outputs[867]));
    assign layer1_outputs[481] = ~(layer0_outputs[331]) | (layer0_outputs[1695]);
    assign layer1_outputs[482] = layer0_outputs[1619];
    assign layer1_outputs[483] = (layer0_outputs[298]) & ~(layer0_outputs[2154]);
    assign layer1_outputs[484] = 1'b0;
    assign layer1_outputs[485] = ~(layer0_outputs[120]) | (layer0_outputs[2177]);
    assign layer1_outputs[486] = 1'b1;
    assign layer1_outputs[487] = ~((layer0_outputs[1485]) & (layer0_outputs[1597]));
    assign layer1_outputs[488] = (layer0_outputs[2478]) & ~(layer0_outputs[2372]);
    assign layer1_outputs[489] = (layer0_outputs[717]) & ~(layer0_outputs[776]);
    assign layer1_outputs[490] = ~((layer0_outputs[2227]) | (layer0_outputs[1660]));
    assign layer1_outputs[491] = ~(layer0_outputs[448]);
    assign layer1_outputs[492] = ~(layer0_outputs[46]) | (layer0_outputs[1373]);
    assign layer1_outputs[493] = layer0_outputs[390];
    assign layer1_outputs[494] = layer0_outputs[2229];
    assign layer1_outputs[495] = ~((layer0_outputs[1421]) | (layer0_outputs[22]));
    assign layer1_outputs[496] = ~(layer0_outputs[2325]);
    assign layer1_outputs[497] = (layer0_outputs[1281]) | (layer0_outputs[612]);
    assign layer1_outputs[498] = ~((layer0_outputs[669]) & (layer0_outputs[17]));
    assign layer1_outputs[499] = (layer0_outputs[1354]) & ~(layer0_outputs[1937]);
    assign layer1_outputs[500] = ~((layer0_outputs[392]) & (layer0_outputs[1143]));
    assign layer1_outputs[501] = layer0_outputs[230];
    assign layer1_outputs[502] = layer0_outputs[1255];
    assign layer1_outputs[503] = (layer0_outputs[264]) & ~(layer0_outputs[2247]);
    assign layer1_outputs[504] = ~(layer0_outputs[1761]);
    assign layer1_outputs[505] = ~((layer0_outputs[1333]) & (layer0_outputs[1943]));
    assign layer1_outputs[506] = ~((layer0_outputs[1960]) | (layer0_outputs[1298]));
    assign layer1_outputs[507] = (layer0_outputs[655]) | (layer0_outputs[2367]);
    assign layer1_outputs[508] = ~(layer0_outputs[1736]);
    assign layer1_outputs[509] = (layer0_outputs[928]) & (layer0_outputs[2079]);
    assign layer1_outputs[510] = (layer0_outputs[2370]) & (layer0_outputs[499]);
    assign layer1_outputs[511] = ~((layer0_outputs[728]) ^ (layer0_outputs[2270]));
    assign layer1_outputs[512] = (layer0_outputs[546]) & (layer0_outputs[1608]);
    assign layer1_outputs[513] = layer0_outputs[643];
    assign layer1_outputs[514] = (layer0_outputs[828]) & (layer0_outputs[1704]);
    assign layer1_outputs[515] = ~(layer0_outputs[1457]) | (layer0_outputs[523]);
    assign layer1_outputs[516] = ~((layer0_outputs[300]) ^ (layer0_outputs[1862]));
    assign layer1_outputs[517] = (layer0_outputs[91]) | (layer0_outputs[1456]);
    assign layer1_outputs[518] = (layer0_outputs[2084]) & (layer0_outputs[1310]);
    assign layer1_outputs[519] = 1'b1;
    assign layer1_outputs[520] = (layer0_outputs[1102]) & ~(layer0_outputs[654]);
    assign layer1_outputs[521] = (layer0_outputs[1480]) & (layer0_outputs[2415]);
    assign layer1_outputs[522] = ~(layer0_outputs[2159]);
    assign layer1_outputs[523] = ~((layer0_outputs[654]) ^ (layer0_outputs[2535]));
    assign layer1_outputs[524] = (layer0_outputs[2398]) | (layer0_outputs[246]);
    assign layer1_outputs[525] = layer0_outputs[877];
    assign layer1_outputs[526] = ~((layer0_outputs[1082]) | (layer0_outputs[932]));
    assign layer1_outputs[527] = (layer0_outputs[223]) & ~(layer0_outputs[395]);
    assign layer1_outputs[528] = (layer0_outputs[822]) | (layer0_outputs[2432]);
    assign layer1_outputs[529] = ~(layer0_outputs[1844]) | (layer0_outputs[1439]);
    assign layer1_outputs[530] = layer0_outputs[727];
    assign layer1_outputs[531] = ~((layer0_outputs[140]) | (layer0_outputs[2405]));
    assign layer1_outputs[532] = (layer0_outputs[324]) & ~(layer0_outputs[2255]);
    assign layer1_outputs[533] = (layer0_outputs[309]) & ~(layer0_outputs[1378]);
    assign layer1_outputs[534] = ~(layer0_outputs[2548]);
    assign layer1_outputs[535] = (layer0_outputs[1054]) | (layer0_outputs[1753]);
    assign layer1_outputs[536] = (layer0_outputs[2239]) ^ (layer0_outputs[1148]);
    assign layer1_outputs[537] = ~(layer0_outputs[2025]);
    assign layer1_outputs[538] = ~((layer0_outputs[2294]) ^ (layer0_outputs[1982]));
    assign layer1_outputs[539] = 1'b0;
    assign layer1_outputs[540] = layer0_outputs[1740];
    assign layer1_outputs[541] = 1'b1;
    assign layer1_outputs[542] = ~(layer0_outputs[1430]);
    assign layer1_outputs[543] = layer0_outputs[2424];
    assign layer1_outputs[544] = 1'b1;
    assign layer1_outputs[545] = (layer0_outputs[826]) & ~(layer0_outputs[948]);
    assign layer1_outputs[546] = ~((layer0_outputs[998]) | (layer0_outputs[277]));
    assign layer1_outputs[547] = (layer0_outputs[2515]) | (layer0_outputs[1853]);
    assign layer1_outputs[548] = 1'b0;
    assign layer1_outputs[549] = (layer0_outputs[1381]) | (layer0_outputs[2324]);
    assign layer1_outputs[550] = (layer0_outputs[572]) ^ (layer0_outputs[5]);
    assign layer1_outputs[551] = ~(layer0_outputs[1812]) | (layer0_outputs[1532]);
    assign layer1_outputs[552] = ~((layer0_outputs[2540]) & (layer0_outputs[803]));
    assign layer1_outputs[553] = 1'b1;
    assign layer1_outputs[554] = 1'b0;
    assign layer1_outputs[555] = (layer0_outputs[1278]) & ~(layer0_outputs[1738]);
    assign layer1_outputs[556] = ~(layer0_outputs[1884]);
    assign layer1_outputs[557] = (layer0_outputs[1953]) ^ (layer0_outputs[2481]);
    assign layer1_outputs[558] = ~((layer0_outputs[967]) | (layer0_outputs[1295]));
    assign layer1_outputs[559] = ~((layer0_outputs[1219]) ^ (layer0_outputs[1969]));
    assign layer1_outputs[560] = ~((layer0_outputs[1225]) | (layer0_outputs[829]));
    assign layer1_outputs[561] = ~((layer0_outputs[1003]) ^ (layer0_outputs[21]));
    assign layer1_outputs[562] = (layer0_outputs[521]) & ~(layer0_outputs[2228]);
    assign layer1_outputs[563] = layer0_outputs[461];
    assign layer1_outputs[564] = ~(layer0_outputs[382]);
    assign layer1_outputs[565] = ~(layer0_outputs[1363]) | (layer0_outputs[244]);
    assign layer1_outputs[566] = (layer0_outputs[750]) & (layer0_outputs[977]);
    assign layer1_outputs[567] = (layer0_outputs[1941]) & ~(layer0_outputs[1438]);
    assign layer1_outputs[568] = layer0_outputs[1717];
    assign layer1_outputs[569] = ~(layer0_outputs[1717]);
    assign layer1_outputs[570] = layer0_outputs[1762];
    assign layer1_outputs[571] = 1'b1;
    assign layer1_outputs[572] = (layer0_outputs[1803]) & ~(layer0_outputs[1855]);
    assign layer1_outputs[573] = (layer0_outputs[613]) ^ (layer0_outputs[872]);
    assign layer1_outputs[574] = (layer0_outputs[759]) | (layer0_outputs[1914]);
    assign layer1_outputs[575] = ~(layer0_outputs[1667]);
    assign layer1_outputs[576] = (layer0_outputs[1647]) & ~(layer0_outputs[265]);
    assign layer1_outputs[577] = (layer0_outputs[2295]) | (layer0_outputs[1303]);
    assign layer1_outputs[578] = 1'b1;
    assign layer1_outputs[579] = ~((layer0_outputs[561]) & (layer0_outputs[1595]));
    assign layer1_outputs[580] = layer0_outputs[1939];
    assign layer1_outputs[581] = (layer0_outputs[1827]) & ~(layer0_outputs[820]);
    assign layer1_outputs[582] = (layer0_outputs[1869]) | (layer0_outputs[1180]);
    assign layer1_outputs[583] = (layer0_outputs[722]) & ~(layer0_outputs[237]);
    assign layer1_outputs[584] = ~(layer0_outputs[893]) | (layer0_outputs[1220]);
    assign layer1_outputs[585] = ~(layer0_outputs[1749]);
    assign layer1_outputs[586] = ~((layer0_outputs[397]) & (layer0_outputs[744]));
    assign layer1_outputs[587] = 1'b1;
    assign layer1_outputs[588] = ~(layer0_outputs[1611]) | (layer0_outputs[1196]);
    assign layer1_outputs[589] = layer0_outputs[1561];
    assign layer1_outputs[590] = ~(layer0_outputs[421]);
    assign layer1_outputs[591] = ~(layer0_outputs[2476]) | (layer0_outputs[2106]);
    assign layer1_outputs[592] = layer0_outputs[2221];
    assign layer1_outputs[593] = layer0_outputs[2345];
    assign layer1_outputs[594] = ~(layer0_outputs[1183]);
    assign layer1_outputs[595] = ~((layer0_outputs[1621]) & (layer0_outputs[20]));
    assign layer1_outputs[596] = ~(layer0_outputs[1274]) | (layer0_outputs[2233]);
    assign layer1_outputs[597] = (layer0_outputs[2392]) | (layer0_outputs[1779]);
    assign layer1_outputs[598] = ~(layer0_outputs[1562]);
    assign layer1_outputs[599] = ~(layer0_outputs[2294]);
    assign layer1_outputs[600] = ~((layer0_outputs[2479]) | (layer0_outputs[2348]));
    assign layer1_outputs[601] = ~(layer0_outputs[1450]) | (layer0_outputs[643]);
    assign layer1_outputs[602] = layer0_outputs[2468];
    assign layer1_outputs[603] = (layer0_outputs[26]) | (layer0_outputs[2173]);
    assign layer1_outputs[604] = ~(layer0_outputs[1165]) | (layer0_outputs[34]);
    assign layer1_outputs[605] = layer0_outputs[1099];
    assign layer1_outputs[606] = (layer0_outputs[2318]) & ~(layer0_outputs[1437]);
    assign layer1_outputs[607] = 1'b0;
    assign layer1_outputs[608] = 1'b0;
    assign layer1_outputs[609] = (layer0_outputs[2368]) & (layer0_outputs[88]);
    assign layer1_outputs[610] = ~(layer0_outputs[1809]) | (layer0_outputs[842]);
    assign layer1_outputs[611] = ~(layer0_outputs[872]);
    assign layer1_outputs[612] = (layer0_outputs[385]) | (layer0_outputs[1737]);
    assign layer1_outputs[613] = ~((layer0_outputs[2220]) & (layer0_outputs[1314]));
    assign layer1_outputs[614] = (layer0_outputs[1446]) | (layer0_outputs[764]);
    assign layer1_outputs[615] = (layer0_outputs[734]) & (layer0_outputs[1429]);
    assign layer1_outputs[616] = ~(layer0_outputs[1629]) | (layer0_outputs[1684]);
    assign layer1_outputs[617] = ~(layer0_outputs[101]) | (layer0_outputs[581]);
    assign layer1_outputs[618] = ~((layer0_outputs[913]) & (layer0_outputs[755]));
    assign layer1_outputs[619] = ~(layer0_outputs[1898]);
    assign layer1_outputs[620] = 1'b1;
    assign layer1_outputs[621] = layer0_outputs[1181];
    assign layer1_outputs[622] = ~(layer0_outputs[1134]);
    assign layer1_outputs[623] = layer0_outputs[207];
    assign layer1_outputs[624] = (layer0_outputs[1116]) & ~(layer0_outputs[2388]);
    assign layer1_outputs[625] = (layer0_outputs[2308]) & (layer0_outputs[1501]);
    assign layer1_outputs[626] = (layer0_outputs[1386]) | (layer0_outputs[2114]);
    assign layer1_outputs[627] = ~((layer0_outputs[1682]) | (layer0_outputs[1852]));
    assign layer1_outputs[628] = 1'b0;
    assign layer1_outputs[629] = 1'b1;
    assign layer1_outputs[630] = (layer0_outputs[1282]) & (layer0_outputs[1579]);
    assign layer1_outputs[631] = layer0_outputs[2122];
    assign layer1_outputs[632] = ~((layer0_outputs[2351]) & (layer0_outputs[381]));
    assign layer1_outputs[633] = 1'b1;
    assign layer1_outputs[634] = ~(layer0_outputs[275]);
    assign layer1_outputs[635] = layer0_outputs[1833];
    assign layer1_outputs[636] = ~((layer0_outputs[1679]) & (layer0_outputs[1894]));
    assign layer1_outputs[637] = ~(layer0_outputs[2418]);
    assign layer1_outputs[638] = ~((layer0_outputs[2482]) ^ (layer0_outputs[259]));
    assign layer1_outputs[639] = layer0_outputs[991];
    assign layer1_outputs[640] = (layer0_outputs[2281]) & (layer0_outputs[1738]);
    assign layer1_outputs[641] = ~(layer0_outputs[2026]) | (layer0_outputs[1605]);
    assign layer1_outputs[642] = (layer0_outputs[1435]) & (layer0_outputs[412]);
    assign layer1_outputs[643] = ~((layer0_outputs[12]) & (layer0_outputs[143]));
    assign layer1_outputs[644] = layer0_outputs[1775];
    assign layer1_outputs[645] = ~(layer0_outputs[1548]);
    assign layer1_outputs[646] = ~(layer0_outputs[282]) | (layer0_outputs[664]);
    assign layer1_outputs[647] = (layer0_outputs[1224]) & ~(layer0_outputs[906]);
    assign layer1_outputs[648] = ~(layer0_outputs[972]);
    assign layer1_outputs[649] = layer0_outputs[2365];
    assign layer1_outputs[650] = layer0_outputs[2541];
    assign layer1_outputs[651] = layer0_outputs[2118];
    assign layer1_outputs[652] = ~(layer0_outputs[404]);
    assign layer1_outputs[653] = ~(layer0_outputs[1300]) | (layer0_outputs[145]);
    assign layer1_outputs[654] = layer0_outputs[180];
    assign layer1_outputs[655] = (layer0_outputs[2454]) & (layer0_outputs[2307]);
    assign layer1_outputs[656] = 1'b0;
    assign layer1_outputs[657] = ~(layer0_outputs[1360]);
    assign layer1_outputs[658] = (layer0_outputs[2269]) & (layer0_outputs[1383]);
    assign layer1_outputs[659] = layer0_outputs[807];
    assign layer1_outputs[660] = 1'b1;
    assign layer1_outputs[661] = (layer0_outputs[1202]) & (layer0_outputs[1535]);
    assign layer1_outputs[662] = ~(layer0_outputs[327]);
    assign layer1_outputs[663] = (layer0_outputs[1088]) & (layer0_outputs[361]);
    assign layer1_outputs[664] = (layer0_outputs[1428]) | (layer0_outputs[2377]);
    assign layer1_outputs[665] = layer0_outputs[1528];
    assign layer1_outputs[666] = layer0_outputs[509];
    assign layer1_outputs[667] = (layer0_outputs[314]) & ~(layer0_outputs[2112]);
    assign layer1_outputs[668] = ~((layer0_outputs[2383]) | (layer0_outputs[1792]));
    assign layer1_outputs[669] = ~((layer0_outputs[285]) | (layer0_outputs[70]));
    assign layer1_outputs[670] = ~((layer0_outputs[388]) ^ (layer0_outputs[2547]));
    assign layer1_outputs[671] = ~(layer0_outputs[1890]) | (layer0_outputs[783]);
    assign layer1_outputs[672] = (layer0_outputs[1362]) & (layer0_outputs[632]);
    assign layer1_outputs[673] = (layer0_outputs[1960]) & (layer0_outputs[1325]);
    assign layer1_outputs[674] = ~(layer0_outputs[1287]) | (layer0_outputs[970]);
    assign layer1_outputs[675] = ~((layer0_outputs[2392]) & (layer0_outputs[656]));
    assign layer1_outputs[676] = ~(layer0_outputs[551]);
    assign layer1_outputs[677] = ~((layer0_outputs[372]) & (layer0_outputs[236]));
    assign layer1_outputs[678] = ~(layer0_outputs[900]);
    assign layer1_outputs[679] = (layer0_outputs[1940]) & ~(layer0_outputs[1807]);
    assign layer1_outputs[680] = (layer0_outputs[1904]) | (layer0_outputs[522]);
    assign layer1_outputs[681] = ~(layer0_outputs[502]);
    assign layer1_outputs[682] = ~(layer0_outputs[681]);
    assign layer1_outputs[683] = (layer0_outputs[2160]) & ~(layer0_outputs[573]);
    assign layer1_outputs[684] = layer0_outputs[2480];
    assign layer1_outputs[685] = layer0_outputs[1570];
    assign layer1_outputs[686] = (layer0_outputs[2417]) & (layer0_outputs[646]);
    assign layer1_outputs[687] = ~((layer0_outputs[1572]) | (layer0_outputs[2506]));
    assign layer1_outputs[688] = 1'b1;
    assign layer1_outputs[689] = ~(layer0_outputs[1335]);
    assign layer1_outputs[690] = (layer0_outputs[495]) | (layer0_outputs[2440]);
    assign layer1_outputs[691] = (layer0_outputs[1496]) & ~(layer0_outputs[1121]);
    assign layer1_outputs[692] = ~(layer0_outputs[454]);
    assign layer1_outputs[693] = ~((layer0_outputs[607]) | (layer0_outputs[2162]));
    assign layer1_outputs[694] = layer0_outputs[2290];
    assign layer1_outputs[695] = ~(layer0_outputs[586]) | (layer0_outputs[285]);
    assign layer1_outputs[696] = (layer0_outputs[720]) & ~(layer0_outputs[1649]);
    assign layer1_outputs[697] = layer0_outputs[1525];
    assign layer1_outputs[698] = ~(layer0_outputs[162]) | (layer0_outputs[2198]);
    assign layer1_outputs[699] = layer0_outputs[2549];
    assign layer1_outputs[700] = (layer0_outputs[1022]) & ~(layer0_outputs[1221]);
    assign layer1_outputs[701] = layer0_outputs[1137];
    assign layer1_outputs[702] = (layer0_outputs[600]) & (layer0_outputs[1771]);
    assign layer1_outputs[703] = ~(layer0_outputs[1306]) | (layer0_outputs[10]);
    assign layer1_outputs[704] = ~(layer0_outputs[2049]) | (layer0_outputs[1483]);
    assign layer1_outputs[705] = 1'b0;
    assign layer1_outputs[706] = layer0_outputs[77];
    assign layer1_outputs[707] = ~(layer0_outputs[321]);
    assign layer1_outputs[708] = ~(layer0_outputs[1675]) | (layer0_outputs[1918]);
    assign layer1_outputs[709] = ~(layer0_outputs[2521]);
    assign layer1_outputs[710] = 1'b1;
    assign layer1_outputs[711] = ~(layer0_outputs[2085]) | (layer0_outputs[1879]);
    assign layer1_outputs[712] = (layer0_outputs[2042]) | (layer0_outputs[1316]);
    assign layer1_outputs[713] = (layer0_outputs[745]) & ~(layer0_outputs[91]);
    assign layer1_outputs[714] = ~(layer0_outputs[387]) | (layer0_outputs[2111]);
    assign layer1_outputs[715] = layer0_outputs[187];
    assign layer1_outputs[716] = ~(layer0_outputs[930]);
    assign layer1_outputs[717] = layer0_outputs[289];
    assign layer1_outputs[718] = (layer0_outputs[1778]) | (layer0_outputs[109]);
    assign layer1_outputs[719] = layer0_outputs[1632];
    assign layer1_outputs[720] = ~(layer0_outputs[256]);
    assign layer1_outputs[721] = (layer0_outputs[1253]) & ~(layer0_outputs[2116]);
    assign layer1_outputs[722] = ~((layer0_outputs[336]) ^ (layer0_outputs[1504]));
    assign layer1_outputs[723] = layer0_outputs[2510];
    assign layer1_outputs[724] = ~(layer0_outputs[538]);
    assign layer1_outputs[725] = layer0_outputs[185];
    assign layer1_outputs[726] = (layer0_outputs[695]) & ~(layer0_outputs[672]);
    assign layer1_outputs[727] = (layer0_outputs[2470]) ^ (layer0_outputs[1110]);
    assign layer1_outputs[728] = layer0_outputs[1336];
    assign layer1_outputs[729] = 1'b0;
    assign layer1_outputs[730] = ~(layer0_outputs[407]) | (layer0_outputs[450]);
    assign layer1_outputs[731] = ~(layer0_outputs[1502]) | (layer0_outputs[2192]);
    assign layer1_outputs[732] = ~((layer0_outputs[2425]) & (layer0_outputs[1012]));
    assign layer1_outputs[733] = ~(layer0_outputs[1640]) | (layer0_outputs[1088]);
    assign layer1_outputs[734] = 1'b0;
    assign layer1_outputs[735] = 1'b1;
    assign layer1_outputs[736] = ~((layer0_outputs[2147]) ^ (layer0_outputs[896]));
    assign layer1_outputs[737] = ~(layer0_outputs[1553]);
    assign layer1_outputs[738] = (layer0_outputs[1472]) & ~(layer0_outputs[1919]);
    assign layer1_outputs[739] = layer0_outputs[417];
    assign layer1_outputs[740] = layer0_outputs[831];
    assign layer1_outputs[741] = (layer0_outputs[1321]) & ~(layer0_outputs[917]);
    assign layer1_outputs[742] = layer0_outputs[594];
    assign layer1_outputs[743] = layer0_outputs[1002];
    assign layer1_outputs[744] = layer0_outputs[866];
    assign layer1_outputs[745] = ~((layer0_outputs[1281]) | (layer0_outputs[2319]));
    assign layer1_outputs[746] = 1'b1;
    assign layer1_outputs[747] = ~((layer0_outputs[1256]) | (layer0_outputs[141]));
    assign layer1_outputs[748] = ~((layer0_outputs[1191]) & (layer0_outputs[1547]));
    assign layer1_outputs[749] = (layer0_outputs[125]) & ~(layer0_outputs[1051]);
    assign layer1_outputs[750] = (layer0_outputs[1052]) & ~(layer0_outputs[665]);
    assign layer1_outputs[751] = (layer0_outputs[1860]) & ~(layer0_outputs[658]);
    assign layer1_outputs[752] = ~(layer0_outputs[835]);
    assign layer1_outputs[753] = ~(layer0_outputs[2201]);
    assign layer1_outputs[754] = (layer0_outputs[1124]) & ~(layer0_outputs[333]);
    assign layer1_outputs[755] = (layer0_outputs[1669]) | (layer0_outputs[259]);
    assign layer1_outputs[756] = ~((layer0_outputs[73]) & (layer0_outputs[1906]));
    assign layer1_outputs[757] = layer0_outputs[653];
    assign layer1_outputs[758] = ~(layer0_outputs[957]) | (layer0_outputs[1478]);
    assign layer1_outputs[759] = ~(layer0_outputs[1839]);
    assign layer1_outputs[760] = 1'b1;
    assign layer1_outputs[761] = layer0_outputs[801];
    assign layer1_outputs[762] = (layer0_outputs[1016]) | (layer0_outputs[2487]);
    assign layer1_outputs[763] = ~((layer0_outputs[1114]) & (layer0_outputs[1186]));
    assign layer1_outputs[764] = (layer0_outputs[2018]) & (layer0_outputs[57]);
    assign layer1_outputs[765] = ~((layer0_outputs[2278]) | (layer0_outputs[2156]));
    assign layer1_outputs[766] = (layer0_outputs[124]) & (layer0_outputs[634]);
    assign layer1_outputs[767] = ~((layer0_outputs[28]) & (layer0_outputs[1145]));
    assign layer1_outputs[768] = layer0_outputs[416];
    assign layer1_outputs[769] = (layer0_outputs[1123]) | (layer0_outputs[1178]);
    assign layer1_outputs[770] = ~(layer0_outputs[111]) | (layer0_outputs[2358]);
    assign layer1_outputs[771] = (layer0_outputs[1758]) & ~(layer0_outputs[402]);
    assign layer1_outputs[772] = ~((layer0_outputs[931]) & (layer0_outputs[2061]));
    assign layer1_outputs[773] = (layer0_outputs[2382]) & ~(layer0_outputs[533]);
    assign layer1_outputs[774] = layer0_outputs[1423];
    assign layer1_outputs[775] = (layer0_outputs[1403]) & ~(layer0_outputs[1805]);
    assign layer1_outputs[776] = ~((layer0_outputs[1766]) & (layer0_outputs[311]));
    assign layer1_outputs[777] = layer0_outputs[2080];
    assign layer1_outputs[778] = ~((layer0_outputs[195]) | (layer0_outputs[1936]));
    assign layer1_outputs[779] = ~((layer0_outputs[2181]) | (layer0_outputs[796]));
    assign layer1_outputs[780] = (layer0_outputs[403]) & ~(layer0_outputs[1481]);
    assign layer1_outputs[781] = (layer0_outputs[1508]) & ~(layer0_outputs[1105]);
    assign layer1_outputs[782] = (layer0_outputs[2446]) & (layer0_outputs[1706]);
    assign layer1_outputs[783] = ~((layer0_outputs[1601]) & (layer0_outputs[1818]));
    assign layer1_outputs[784] = layer0_outputs[743];
    assign layer1_outputs[785] = (layer0_outputs[1844]) & (layer0_outputs[2075]);
    assign layer1_outputs[786] = ~((layer0_outputs[1882]) | (layer0_outputs[48]));
    assign layer1_outputs[787] = ~(layer0_outputs[1929]);
    assign layer1_outputs[788] = ~(layer0_outputs[1460]) | (layer0_outputs[1613]);
    assign layer1_outputs[789] = (layer0_outputs[1940]) & (layer0_outputs[1030]);
    assign layer1_outputs[790] = (layer0_outputs[1350]) ^ (layer0_outputs[1278]);
    assign layer1_outputs[791] = layer0_outputs[984];
    assign layer1_outputs[792] = (layer0_outputs[231]) | (layer0_outputs[119]);
    assign layer1_outputs[793] = (layer0_outputs[2045]) | (layer0_outputs[354]);
    assign layer1_outputs[794] = ~(layer0_outputs[366]) | (layer0_outputs[1455]);
    assign layer1_outputs[795] = (layer0_outputs[2223]) | (layer0_outputs[1524]);
    assign layer1_outputs[796] = (layer0_outputs[1470]) & ~(layer0_outputs[304]);
    assign layer1_outputs[797] = (layer0_outputs[438]) & ~(layer0_outputs[1955]);
    assign layer1_outputs[798] = (layer0_outputs[1538]) & (layer0_outputs[449]);
    assign layer1_outputs[799] = ~(layer0_outputs[2127]) | (layer0_outputs[256]);
    assign layer1_outputs[800] = 1'b0;
    assign layer1_outputs[801] = ~(layer0_outputs[780]);
    assign layer1_outputs[802] = ~((layer0_outputs[2461]) | (layer0_outputs[1585]));
    assign layer1_outputs[803] = ~(layer0_outputs[677]);
    assign layer1_outputs[804] = layer0_outputs[2488];
    assign layer1_outputs[805] = ~(layer0_outputs[1676]);
    assign layer1_outputs[806] = ~((layer0_outputs[652]) | (layer0_outputs[1820]));
    assign layer1_outputs[807] = ~((layer0_outputs[1612]) | (layer0_outputs[1320]));
    assign layer1_outputs[808] = (layer0_outputs[679]) & (layer0_outputs[1039]);
    assign layer1_outputs[809] = 1'b0;
    assign layer1_outputs[810] = 1'b1;
    assign layer1_outputs[811] = layer0_outputs[968];
    assign layer1_outputs[812] = ~(layer0_outputs[1214]);
    assign layer1_outputs[813] = (layer0_outputs[1762]) ^ (layer0_outputs[2279]);
    assign layer1_outputs[814] = (layer0_outputs[2279]) ^ (layer0_outputs[1257]);
    assign layer1_outputs[815] = (layer0_outputs[309]) & ~(layer0_outputs[2210]);
    assign layer1_outputs[816] = ~(layer0_outputs[1135]);
    assign layer1_outputs[817] = layer0_outputs[1119];
    assign layer1_outputs[818] = (layer0_outputs[2065]) & (layer0_outputs[132]);
    assign layer1_outputs[819] = 1'b0;
    assign layer1_outputs[820] = (layer0_outputs[2015]) & ~(layer0_outputs[2385]);
    assign layer1_outputs[821] = (layer0_outputs[1745]) & ~(layer0_outputs[1883]);
    assign layer1_outputs[822] = ~(layer0_outputs[362]) | (layer0_outputs[910]);
    assign layer1_outputs[823] = (layer0_outputs[2323]) & (layer0_outputs[1739]);
    assign layer1_outputs[824] = ~((layer0_outputs[1352]) | (layer0_outputs[1935]));
    assign layer1_outputs[825] = ~(layer0_outputs[764]) | (layer0_outputs[416]);
    assign layer1_outputs[826] = layer0_outputs[2342];
    assign layer1_outputs[827] = (layer0_outputs[338]) | (layer0_outputs[646]);
    assign layer1_outputs[828] = 1'b0;
    assign layer1_outputs[829] = (layer0_outputs[1033]) ^ (layer0_outputs[2482]);
    assign layer1_outputs[830] = ~(layer0_outputs[808]);
    assign layer1_outputs[831] = ~(layer0_outputs[499]) | (layer0_outputs[629]);
    assign layer1_outputs[832] = ~(layer0_outputs[2467]) | (layer0_outputs[1079]);
    assign layer1_outputs[833] = 1'b1;
    assign layer1_outputs[834] = layer0_outputs[1682];
    assign layer1_outputs[835] = ~(layer0_outputs[1948]) | (layer0_outputs[1050]);
    assign layer1_outputs[836] = 1'b1;
    assign layer1_outputs[837] = ~(layer0_outputs[1059]);
    assign layer1_outputs[838] = layer0_outputs[1356];
    assign layer1_outputs[839] = (layer0_outputs[1048]) & (layer0_outputs[2282]);
    assign layer1_outputs[840] = 1'b1;
    assign layer1_outputs[841] = ~((layer0_outputs[2337]) & (layer0_outputs[110]));
    assign layer1_outputs[842] = (layer0_outputs[2262]) & ~(layer0_outputs[615]);
    assign layer1_outputs[843] = layer0_outputs[2533];
    assign layer1_outputs[844] = 1'b0;
    assign layer1_outputs[845] = ~(layer0_outputs[2238]) | (layer0_outputs[2462]);
    assign layer1_outputs[846] = layer0_outputs[2129];
    assign layer1_outputs[847] = ~((layer0_outputs[406]) & (layer0_outputs[2315]));
    assign layer1_outputs[848] = (layer0_outputs[35]) | (layer0_outputs[1458]);
    assign layer1_outputs[849] = layer0_outputs[610];
    assign layer1_outputs[850] = layer0_outputs[1404];
    assign layer1_outputs[851] = layer0_outputs[706];
    assign layer1_outputs[852] = ~(layer0_outputs[789]) | (layer0_outputs[190]);
    assign layer1_outputs[853] = ~(layer0_outputs[2481]) | (layer0_outputs[1996]);
    assign layer1_outputs[854] = ~(layer0_outputs[1983]);
    assign layer1_outputs[855] = ~((layer0_outputs[1417]) ^ (layer0_outputs[1071]));
    assign layer1_outputs[856] = ~((layer0_outputs[882]) | (layer0_outputs[253]));
    assign layer1_outputs[857] = ~((layer0_outputs[2135]) & (layer0_outputs[2504]));
    assign layer1_outputs[858] = ~((layer0_outputs[1244]) & (layer0_outputs[459]));
    assign layer1_outputs[859] = ~(layer0_outputs[962]);
    assign layer1_outputs[860] = (layer0_outputs[543]) & ~(layer0_outputs[1351]);
    assign layer1_outputs[861] = 1'b0;
    assign layer1_outputs[862] = 1'b0;
    assign layer1_outputs[863] = 1'b0;
    assign layer1_outputs[864] = ~(layer0_outputs[1288]);
    assign layer1_outputs[865] = (layer0_outputs[291]) & ~(layer0_outputs[2362]);
    assign layer1_outputs[866] = 1'b0;
    assign layer1_outputs[867] = (layer0_outputs[1678]) & (layer0_outputs[234]);
    assign layer1_outputs[868] = (layer0_outputs[2553]) | (layer0_outputs[1560]);
    assign layer1_outputs[869] = ~(layer0_outputs[925]) | (layer0_outputs[498]);
    assign layer1_outputs[870] = layer0_outputs[1628];
    assign layer1_outputs[871] = 1'b1;
    assign layer1_outputs[872] = ~(layer0_outputs[1554]) | (layer0_outputs[2421]);
    assign layer1_outputs[873] = ~(layer0_outputs[2381]);
    assign layer1_outputs[874] = ~((layer0_outputs[1828]) | (layer0_outputs[1039]));
    assign layer1_outputs[875] = layer0_outputs[1830];
    assign layer1_outputs[876] = ~(layer0_outputs[187]) | (layer0_outputs[484]);
    assign layer1_outputs[877] = layer0_outputs[488];
    assign layer1_outputs[878] = layer0_outputs[1482];
    assign layer1_outputs[879] = ~((layer0_outputs[52]) | (layer0_outputs[15]));
    assign layer1_outputs[880] = (layer0_outputs[2383]) & ~(layer0_outputs[1922]);
    assign layer1_outputs[881] = ~(layer0_outputs[652]);
    assign layer1_outputs[882] = layer0_outputs[1476];
    assign layer1_outputs[883] = (layer0_outputs[1372]) | (layer0_outputs[1768]);
    assign layer1_outputs[884] = (layer0_outputs[2328]) & ~(layer0_outputs[1141]);
    assign layer1_outputs[885] = ~((layer0_outputs[2499]) & (layer0_outputs[911]));
    assign layer1_outputs[886] = (layer0_outputs[208]) & (layer0_outputs[1657]);
    assign layer1_outputs[887] = (layer0_outputs[603]) & ~(layer0_outputs[988]);
    assign layer1_outputs[888] = 1'b1;
    assign layer1_outputs[889] = ~(layer0_outputs[1950]);
    assign layer1_outputs[890] = ~(layer0_outputs[1625]);
    assign layer1_outputs[891] = layer0_outputs[79];
    assign layer1_outputs[892] = ~(layer0_outputs[307]) | (layer0_outputs[1654]);
    assign layer1_outputs[893] = layer0_outputs[1503];
    assign layer1_outputs[894] = ~(layer0_outputs[1952]);
    assign layer1_outputs[895] = 1'b0;
    assign layer1_outputs[896] = ~((layer0_outputs[681]) & (layer0_outputs[181]));
    assign layer1_outputs[897] = (layer0_outputs[1297]) & ~(layer0_outputs[1359]);
    assign layer1_outputs[898] = (layer0_outputs[2500]) | (layer0_outputs[2327]);
    assign layer1_outputs[899] = ~(layer0_outputs[1680]);
    assign layer1_outputs[900] = layer0_outputs[1161];
    assign layer1_outputs[901] = 1'b0;
    assign layer1_outputs[902] = ~((layer0_outputs[1854]) & (layer0_outputs[666]));
    assign layer1_outputs[903] = ~(layer0_outputs[222]);
    assign layer1_outputs[904] = ~(layer0_outputs[2298]);
    assign layer1_outputs[905] = 1'b0;
    assign layer1_outputs[906] = ~(layer0_outputs[182]);
    assign layer1_outputs[907] = ~(layer0_outputs[2490]) | (layer0_outputs[698]);
    assign layer1_outputs[908] = ~(layer0_outputs[881]) | (layer0_outputs[1336]);
    assign layer1_outputs[909] = layer0_outputs[2175];
    assign layer1_outputs[910] = layer0_outputs[1509];
    assign layer1_outputs[911] = ~((layer0_outputs[1283]) & (layer0_outputs[2089]));
    assign layer1_outputs[912] = 1'b1;
    assign layer1_outputs[913] = layer0_outputs[349];
    assign layer1_outputs[914] = ~(layer0_outputs[1308]);
    assign layer1_outputs[915] = ~(layer0_outputs[558]);
    assign layer1_outputs[916] = ~((layer0_outputs[1355]) | (layer0_outputs[1041]));
    assign layer1_outputs[917] = ~((layer0_outputs[1337]) | (layer0_outputs[1535]));
    assign layer1_outputs[918] = ~((layer0_outputs[288]) & (layer0_outputs[1141]));
    assign layer1_outputs[919] = ~(layer0_outputs[1398]);
    assign layer1_outputs[920] = ~((layer0_outputs[1741]) | (layer0_outputs[2544]));
    assign layer1_outputs[921] = ~(layer0_outputs[1663]);
    assign layer1_outputs[922] = (layer0_outputs[451]) & (layer0_outputs[2409]);
    assign layer1_outputs[923] = ~((layer0_outputs[687]) & (layer0_outputs[1731]));
    assign layer1_outputs[924] = ~((layer0_outputs[1271]) & (layer0_outputs[299]));
    assign layer1_outputs[925] = (layer0_outputs[89]) & ~(layer0_outputs[1240]);
    assign layer1_outputs[926] = ~((layer0_outputs[350]) ^ (layer0_outputs[1791]));
    assign layer1_outputs[927] = (layer0_outputs[2213]) & (layer0_outputs[858]);
    assign layer1_outputs[928] = ~(layer0_outputs[391]) | (layer0_outputs[864]);
    assign layer1_outputs[929] = ~(layer0_outputs[1064]) | (layer0_outputs[1998]);
    assign layer1_outputs[930] = layer0_outputs[710];
    assign layer1_outputs[931] = ~((layer0_outputs[2102]) | (layer0_outputs[301]));
    assign layer1_outputs[932] = ~(layer0_outputs[1586]) | (layer0_outputs[2495]);
    assign layer1_outputs[933] = (layer0_outputs[2337]) & (layer0_outputs[1277]);
    assign layer1_outputs[934] = (layer0_outputs[2134]) & ~(layer0_outputs[1921]);
    assign layer1_outputs[935] = ~(layer0_outputs[593]) | (layer0_outputs[2355]);
    assign layer1_outputs[936] = ~(layer0_outputs[527]) | (layer0_outputs[808]);
    assign layer1_outputs[937] = ~(layer0_outputs[529]);
    assign layer1_outputs[938] = ~((layer0_outputs[1210]) | (layer0_outputs[1167]));
    assign layer1_outputs[939] = 1'b0;
    assign layer1_outputs[940] = ~(layer0_outputs[1653]) | (layer0_outputs[20]);
    assign layer1_outputs[941] = ~(layer0_outputs[2039]);
    assign layer1_outputs[942] = ~((layer0_outputs[765]) & (layer0_outputs[1949]));
    assign layer1_outputs[943] = layer0_outputs[2330];
    assign layer1_outputs[944] = ~(layer0_outputs[530]) | (layer0_outputs[8]);
    assign layer1_outputs[945] = (layer0_outputs[2437]) & (layer0_outputs[1926]);
    assign layer1_outputs[946] = 1'b1;
    assign layer1_outputs[947] = ~((layer0_outputs[284]) ^ (layer0_outputs[13]));
    assign layer1_outputs[948] = ~((layer0_outputs[751]) | (layer0_outputs[1270]));
    assign layer1_outputs[949] = layer0_outputs[1655];
    assign layer1_outputs[950] = ~(layer0_outputs[1463]);
    assign layer1_outputs[951] = (layer0_outputs[1001]) & ~(layer0_outputs[1571]);
    assign layer1_outputs[952] = 1'b1;
    assign layer1_outputs[953] = layer0_outputs[1092];
    assign layer1_outputs[954] = layer0_outputs[2555];
    assign layer1_outputs[955] = 1'b0;
    assign layer1_outputs[956] = ~(layer0_outputs[2186]);
    assign layer1_outputs[957] = ~(layer0_outputs[146]) | (layer0_outputs[1245]);
    assign layer1_outputs[958] = ~((layer0_outputs[1550]) ^ (layer0_outputs[986]));
    assign layer1_outputs[959] = ~(layer0_outputs[162]) | (layer0_outputs[1116]);
    assign layer1_outputs[960] = (layer0_outputs[1234]) & ~(layer0_outputs[584]);
    assign layer1_outputs[961] = ~((layer0_outputs[1789]) ^ (layer0_outputs[1863]));
    assign layer1_outputs[962] = (layer0_outputs[854]) & ~(layer0_outputs[2081]);
    assign layer1_outputs[963] = layer0_outputs[440];
    assign layer1_outputs[964] = 1'b0;
    assign layer1_outputs[965] = 1'b1;
    assign layer1_outputs[966] = (layer0_outputs[2435]) & ~(layer0_outputs[1687]);
    assign layer1_outputs[967] = ~(layer0_outputs[298]);
    assign layer1_outputs[968] = ~(layer0_outputs[275]);
    assign layer1_outputs[969] = layer0_outputs[1998];
    assign layer1_outputs[970] = 1'b1;
    assign layer1_outputs[971] = 1'b0;
    assign layer1_outputs[972] = (layer0_outputs[1047]) & (layer0_outputs[2550]);
    assign layer1_outputs[973] = layer0_outputs[1924];
    assign layer1_outputs[974] = (layer0_outputs[235]) & ~(layer0_outputs[128]);
    assign layer1_outputs[975] = (layer0_outputs[785]) & ~(layer0_outputs[1406]);
    assign layer1_outputs[976] = ~((layer0_outputs[688]) | (layer0_outputs[425]));
    assign layer1_outputs[977] = ~((layer0_outputs[1279]) & (layer0_outputs[2234]));
    assign layer1_outputs[978] = ~(layer0_outputs[435]) | (layer0_outputs[1285]);
    assign layer1_outputs[979] = ~(layer0_outputs[210]) | (layer0_outputs[1426]);
    assign layer1_outputs[980] = ~(layer0_outputs[2386]);
    assign layer1_outputs[981] = ~((layer0_outputs[2088]) & (layer0_outputs[151]));
    assign layer1_outputs[982] = ~(layer0_outputs[704]);
    assign layer1_outputs[983] = 1'b1;
    assign layer1_outputs[984] = layer0_outputs[1295];
    assign layer1_outputs[985] = 1'b0;
    assign layer1_outputs[986] = ~(layer0_outputs[884]) | (layer0_outputs[996]);
    assign layer1_outputs[987] = ~(layer0_outputs[1465]);
    assign layer1_outputs[988] = 1'b0;
    assign layer1_outputs[989] = ~((layer0_outputs[1015]) | (layer0_outputs[2045]));
    assign layer1_outputs[990] = (layer0_outputs[1212]) & (layer0_outputs[1190]);
    assign layer1_outputs[991] = 1'b0;
    assign layer1_outputs[992] = ~((layer0_outputs[597]) & (layer0_outputs[104]));
    assign layer1_outputs[993] = ~(layer0_outputs[2138]);
    assign layer1_outputs[994] = ~((layer0_outputs[25]) & (layer0_outputs[0]));
    assign layer1_outputs[995] = layer0_outputs[863];
    assign layer1_outputs[996] = 1'b0;
    assign layer1_outputs[997] = ~(layer0_outputs[1907]);
    assign layer1_outputs[998] = (layer0_outputs[2490]) & ~(layer0_outputs[827]);
    assign layer1_outputs[999] = layer0_outputs[1930];
    assign layer1_outputs[1000] = 1'b0;
    assign layer1_outputs[1001] = ~((layer0_outputs[897]) | (layer0_outputs[2287]));
    assign layer1_outputs[1002] = ~(layer0_outputs[1466]) | (layer0_outputs[1652]);
    assign layer1_outputs[1003] = layer0_outputs[2522];
    assign layer1_outputs[1004] = (layer0_outputs[2471]) & ~(layer0_outputs[8]);
    assign layer1_outputs[1005] = 1'b0;
    assign layer1_outputs[1006] = ~(layer0_outputs[313]);
    assign layer1_outputs[1007] = ~(layer0_outputs[2066]) | (layer0_outputs[83]);
    assign layer1_outputs[1008] = (layer0_outputs[216]) | (layer0_outputs[926]);
    assign layer1_outputs[1009] = ~(layer0_outputs[781]) | (layer0_outputs[946]);
    assign layer1_outputs[1010] = ~(layer0_outputs[380]);
    assign layer1_outputs[1011] = (layer0_outputs[2107]) | (layer0_outputs[363]);
    assign layer1_outputs[1012] = (layer0_outputs[1435]) ^ (layer0_outputs[1156]);
    assign layer1_outputs[1013] = ~((layer0_outputs[1935]) & (layer0_outputs[2474]));
    assign layer1_outputs[1014] = (layer0_outputs[626]) & ~(layer0_outputs[50]);
    assign layer1_outputs[1015] = ~((layer0_outputs[541]) | (layer0_outputs[2197]));
    assign layer1_outputs[1016] = (layer0_outputs[2235]) & ~(layer0_outputs[1967]);
    assign layer1_outputs[1017] = layer0_outputs[1028];
    assign layer1_outputs[1018] = ~(layer0_outputs[1726]) | (layer0_outputs[1129]);
    assign layer1_outputs[1019] = ~(layer0_outputs[1506]);
    assign layer1_outputs[1020] = ~(layer0_outputs[553]) | (layer0_outputs[516]);
    assign layer1_outputs[1021] = ~(layer0_outputs[1865]) | (layer0_outputs[502]);
    assign layer1_outputs[1022] = layer0_outputs[1903];
    assign layer1_outputs[1023] = (layer0_outputs[843]) & (layer0_outputs[784]);
    assign layer1_outputs[1024] = 1'b0;
    assign layer1_outputs[1025] = layer0_outputs[78];
    assign layer1_outputs[1026] = (layer0_outputs[1836]) ^ (layer0_outputs[967]);
    assign layer1_outputs[1027] = (layer0_outputs[469]) & (layer0_outputs[2280]);
    assign layer1_outputs[1028] = ~(layer0_outputs[1340]) | (layer0_outputs[2257]);
    assign layer1_outputs[1029] = ~(layer0_outputs[1325]) | (layer0_outputs[484]);
    assign layer1_outputs[1030] = (layer0_outputs[1016]) ^ (layer0_outputs[202]);
    assign layer1_outputs[1031] = (layer0_outputs[510]) & (layer0_outputs[1208]);
    assign layer1_outputs[1032] = (layer0_outputs[592]) & (layer0_outputs[447]);
    assign layer1_outputs[1033] = layer0_outputs[2047];
    assign layer1_outputs[1034] = ~(layer0_outputs[1011]);
    assign layer1_outputs[1035] = 1'b1;
    assign layer1_outputs[1036] = ~(layer0_outputs[2411]);
    assign layer1_outputs[1037] = ~(layer0_outputs[2057]) | (layer0_outputs[397]);
    assign layer1_outputs[1038] = (layer0_outputs[1616]) & ~(layer0_outputs[225]);
    assign layer1_outputs[1039] = ~(layer0_outputs[1702]);
    assign layer1_outputs[1040] = ~(layer0_outputs[1916]);
    assign layer1_outputs[1041] = layer0_outputs[2500];
    assign layer1_outputs[1042] = layer0_outputs[1407];
    assign layer1_outputs[1043] = 1'b0;
    assign layer1_outputs[1044] = ~(layer0_outputs[1973]);
    assign layer1_outputs[1045] = ~(layer0_outputs[2518]);
    assign layer1_outputs[1046] = layer0_outputs[1815];
    assign layer1_outputs[1047] = ~(layer0_outputs[1179]) | (layer0_outputs[1795]);
    assign layer1_outputs[1048] = (layer0_outputs[2113]) | (layer0_outputs[1594]);
    assign layer1_outputs[1049] = (layer0_outputs[934]) ^ (layer0_outputs[557]);
    assign layer1_outputs[1050] = 1'b0;
    assign layer1_outputs[1051] = (layer0_outputs[749]) & ~(layer0_outputs[852]);
    assign layer1_outputs[1052] = ~((layer0_outputs[1520]) & (layer0_outputs[958]));
    assign layer1_outputs[1053] = layer0_outputs[1426];
    assign layer1_outputs[1054] = ~(layer0_outputs[758]);
    assign layer1_outputs[1055] = ~(layer0_outputs[2483]) | (layer0_outputs[834]);
    assign layer1_outputs[1056] = 1'b0;
    assign layer1_outputs[1057] = (layer0_outputs[1542]) & ~(layer0_outputs[2397]);
    assign layer1_outputs[1058] = (layer0_outputs[2007]) & (layer0_outputs[1848]);
    assign layer1_outputs[1059] = ~((layer0_outputs[965]) & (layer0_outputs[2288]));
    assign layer1_outputs[1060] = ~(layer0_outputs[1612]) | (layer0_outputs[810]);
    assign layer1_outputs[1061] = ~(layer0_outputs[565]);
    assign layer1_outputs[1062] = (layer0_outputs[1505]) & (layer0_outputs[2440]);
    assign layer1_outputs[1063] = (layer0_outputs[239]) & ~(layer0_outputs[1548]);
    assign layer1_outputs[1064] = ~((layer0_outputs[2519]) | (layer0_outputs[2012]));
    assign layer1_outputs[1065] = (layer0_outputs[1464]) | (layer0_outputs[134]);
    assign layer1_outputs[1066] = layer0_outputs[2347];
    assign layer1_outputs[1067] = layer0_outputs[2016];
    assign layer1_outputs[1068] = ~((layer0_outputs[2373]) ^ (layer0_outputs[603]));
    assign layer1_outputs[1069] = 1'b1;
    assign layer1_outputs[1070] = (layer0_outputs[1995]) & ~(layer0_outputs[623]);
    assign layer1_outputs[1071] = ~((layer0_outputs[1931]) ^ (layer0_outputs[1342]));
    assign layer1_outputs[1072] = (layer0_outputs[2179]) & (layer0_outputs[1130]);
    assign layer1_outputs[1073] = ~(layer0_outputs[1563]) | (layer0_outputs[1600]);
    assign layer1_outputs[1074] = ~(layer0_outputs[1694]) | (layer0_outputs[969]);
    assign layer1_outputs[1075] = ~(layer0_outputs[2027]) | (layer0_outputs[2368]);
    assign layer1_outputs[1076] = (layer0_outputs[444]) & (layer0_outputs[248]);
    assign layer1_outputs[1077] = (layer0_outputs[856]) & ~(layer0_outputs[1492]);
    assign layer1_outputs[1078] = 1'b0;
    assign layer1_outputs[1079] = layer0_outputs[17];
    assign layer1_outputs[1080] = (layer0_outputs[1101]) | (layer0_outputs[816]);
    assign layer1_outputs[1081] = layer0_outputs[1009];
    assign layer1_outputs[1082] = (layer0_outputs[1511]) & (layer0_outputs[637]);
    assign layer1_outputs[1083] = ~(layer0_outputs[196]);
    assign layer1_outputs[1084] = ~(layer0_outputs[2153]) | (layer0_outputs[1356]);
    assign layer1_outputs[1085] = ~(layer0_outputs[2534]);
    assign layer1_outputs[1086] = layer0_outputs[1891];
    assign layer1_outputs[1087] = ~(layer0_outputs[1966]);
    assign layer1_outputs[1088] = ~((layer0_outputs[95]) & (layer0_outputs[188]));
    assign layer1_outputs[1089] = ~((layer0_outputs[801]) & (layer0_outputs[673]));
    assign layer1_outputs[1090] = ~(layer0_outputs[205]) | (layer0_outputs[409]);
    assign layer1_outputs[1091] = (layer0_outputs[961]) ^ (layer0_outputs[1383]);
    assign layer1_outputs[1092] = ~(layer0_outputs[2218]);
    assign layer1_outputs[1093] = ~((layer0_outputs[2332]) | (layer0_outputs[734]));
    assign layer1_outputs[1094] = (layer0_outputs[1834]) ^ (layer0_outputs[2238]);
    assign layer1_outputs[1095] = ~(layer0_outputs[960]) | (layer0_outputs[1104]);
    assign layer1_outputs[1096] = layer0_outputs[1801];
    assign layer1_outputs[1097] = layer0_outputs[2479];
    assign layer1_outputs[1098] = ~(layer0_outputs[914]);
    assign layer1_outputs[1099] = ~(layer0_outputs[1794]) | (layer0_outputs[1233]);
    assign layer1_outputs[1100] = (layer0_outputs[1956]) & (layer0_outputs[1821]);
    assign layer1_outputs[1101] = layer0_outputs[2280];
    assign layer1_outputs[1102] = (layer0_outputs[14]) & (layer0_outputs[208]);
    assign layer1_outputs[1103] = ~(layer0_outputs[766]) | (layer0_outputs[1367]);
    assign layer1_outputs[1104] = ~(layer0_outputs[428]);
    assign layer1_outputs[1105] = (layer0_outputs[1957]) & (layer0_outputs[1056]);
    assign layer1_outputs[1106] = layer0_outputs[1969];
    assign layer1_outputs[1107] = ~((layer0_outputs[870]) | (layer0_outputs[494]));
    assign layer1_outputs[1108] = ~(layer0_outputs[394]) | (layer0_outputs[2367]);
    assign layer1_outputs[1109] = 1'b0;
    assign layer1_outputs[1110] = layer0_outputs[2530];
    assign layer1_outputs[1111] = ~((layer0_outputs[1332]) | (layer0_outputs[2430]));
    assign layer1_outputs[1112] = ~(layer0_outputs[1346]);
    assign layer1_outputs[1113] = (layer0_outputs[1505]) & (layer0_outputs[1388]);
    assign layer1_outputs[1114] = 1'b1;
    assign layer1_outputs[1115] = ~(layer0_outputs[272]);
    assign layer1_outputs[1116] = 1'b0;
    assign layer1_outputs[1117] = layer0_outputs[345];
    assign layer1_outputs[1118] = ~(layer0_outputs[1810]) | (layer0_outputs[254]);
    assign layer1_outputs[1119] = 1'b0;
    assign layer1_outputs[1120] = layer0_outputs[1354];
    assign layer1_outputs[1121] = (layer0_outputs[1751]) & ~(layer0_outputs[1153]);
    assign layer1_outputs[1122] = (layer0_outputs[1401]) & (layer0_outputs[651]);
    assign layer1_outputs[1123] = ~(layer0_outputs[964]);
    assign layer1_outputs[1124] = (layer0_outputs[807]) | (layer0_outputs[2451]);
    assign layer1_outputs[1125] = ~(layer0_outputs[270]);
    assign layer1_outputs[1126] = (layer0_outputs[2441]) & ~(layer0_outputs[2556]);
    assign layer1_outputs[1127] = ~((layer0_outputs[2040]) | (layer0_outputs[389]));
    assign layer1_outputs[1128] = (layer0_outputs[2539]) & ~(layer0_outputs[2395]);
    assign layer1_outputs[1129] = ~(layer0_outputs[1881]);
    assign layer1_outputs[1130] = 1'b1;
    assign layer1_outputs[1131] = 1'b1;
    assign layer1_outputs[1132] = layer0_outputs[554];
    assign layer1_outputs[1133] = (layer0_outputs[1630]) & ~(layer0_outputs[1851]);
    assign layer1_outputs[1134] = ~(layer0_outputs[1696]);
    assign layer1_outputs[1135] = (layer0_outputs[2257]) & (layer0_outputs[481]);
    assign layer1_outputs[1136] = ~(layer0_outputs[2052]);
    assign layer1_outputs[1137] = layer0_outputs[576];
    assign layer1_outputs[1138] = ~((layer0_outputs[2201]) ^ (layer0_outputs[1615]));
    assign layer1_outputs[1139] = ~((layer0_outputs[1693]) ^ (layer0_outputs[2108]));
    assign layer1_outputs[1140] = layer0_outputs[1030];
    assign layer1_outputs[1141] = 1'b1;
    assign layer1_outputs[1142] = ~(layer0_outputs[1290]) | (layer0_outputs[1376]);
    assign layer1_outputs[1143] = ~(layer0_outputs[2414]);
    assign layer1_outputs[1144] = (layer0_outputs[1003]) & (layer0_outputs[661]);
    assign layer1_outputs[1145] = 1'b1;
    assign layer1_outputs[1146] = ~(layer0_outputs[1554]);
    assign layer1_outputs[1147] = ~(layer0_outputs[1573]) | (layer0_outputs[463]);
    assign layer1_outputs[1148] = ~(layer0_outputs[1425]);
    assign layer1_outputs[1149] = (layer0_outputs[1968]) & ~(layer0_outputs[1517]);
    assign layer1_outputs[1150] = ~((layer0_outputs[44]) | (layer0_outputs[1117]));
    assign layer1_outputs[1151] = layer0_outputs[1636];
    assign layer1_outputs[1152] = (layer0_outputs[98]) & ~(layer0_outputs[1708]);
    assign layer1_outputs[1153] = ~(layer0_outputs[1622]);
    assign layer1_outputs[1154] = ~((layer0_outputs[1987]) & (layer0_outputs[1131]));
    assign layer1_outputs[1155] = ~(layer0_outputs[1829]) | (layer0_outputs[63]);
    assign layer1_outputs[1156] = ~(layer0_outputs[1316]) | (layer0_outputs[319]);
    assign layer1_outputs[1157] = (layer0_outputs[556]) & ~(layer0_outputs[1543]);
    assign layer1_outputs[1158] = (layer0_outputs[1697]) | (layer0_outputs[2185]);
    assign layer1_outputs[1159] = layer0_outputs[1304];
    assign layer1_outputs[1160] = ~(layer0_outputs[1662]) | (layer0_outputs[1944]);
    assign layer1_outputs[1161] = ~((layer0_outputs[228]) & (layer0_outputs[1663]));
    assign layer1_outputs[1162] = 1'b1;
    assign layer1_outputs[1163] = ~(layer0_outputs[1728]);
    assign layer1_outputs[1164] = layer0_outputs[371];
    assign layer1_outputs[1165] = (layer0_outputs[2021]) & ~(layer0_outputs[1734]);
    assign layer1_outputs[1166] = ~(layer0_outputs[2266]);
    assign layer1_outputs[1167] = 1'b0;
    assign layer1_outputs[1168] = ~(layer0_outputs[487]);
    assign layer1_outputs[1169] = layer0_outputs[2445];
    assign layer1_outputs[1170] = ~((layer0_outputs[589]) & (layer0_outputs[2022]));
    assign layer1_outputs[1171] = (layer0_outputs[862]) & ~(layer0_outputs[2492]);
    assign layer1_outputs[1172] = (layer0_outputs[2098]) & ~(layer0_outputs[2052]);
    assign layer1_outputs[1173] = (layer0_outputs[692]) & ~(layer0_outputs[876]);
    assign layer1_outputs[1174] = ~(layer0_outputs[1846]);
    assign layer1_outputs[1175] = ~((layer0_outputs[1307]) & (layer0_outputs[1513]));
    assign layer1_outputs[1176] = ~(layer0_outputs[1773]) | (layer0_outputs[1512]);
    assign layer1_outputs[1177] = layer0_outputs[628];
    assign layer1_outputs[1178] = ~(layer0_outputs[1024]) | (layer0_outputs[1484]);
    assign layer1_outputs[1179] = layer0_outputs[2150];
    assign layer1_outputs[1180] = ~(layer0_outputs[1317]);
    assign layer1_outputs[1181] = 1'b1;
    assign layer1_outputs[1182] = ~((layer0_outputs[2558]) & (layer0_outputs[1012]));
    assign layer1_outputs[1183] = (layer0_outputs[1605]) & (layer0_outputs[907]);
    assign layer1_outputs[1184] = ~(layer0_outputs[980]);
    assign layer1_outputs[1185] = 1'b0;
    assign layer1_outputs[1186] = ~(layer0_outputs[2254]) | (layer0_outputs[2501]);
    assign layer1_outputs[1187] = ~(layer0_outputs[4]);
    assign layer1_outputs[1188] = ~(layer0_outputs[469]);
    assign layer1_outputs[1189] = ~((layer0_outputs[1858]) & (layer0_outputs[1229]));
    assign layer1_outputs[1190] = layer0_outputs[2251];
    assign layer1_outputs[1191] = ~(layer0_outputs[611]) | (layer0_outputs[828]);
    assign layer1_outputs[1192] = ~(layer0_outputs[1780]);
    assign layer1_outputs[1193] = ~(layer0_outputs[19]);
    assign layer1_outputs[1194] = (layer0_outputs[1743]) ^ (layer0_outputs[1206]);
    assign layer1_outputs[1195] = ~((layer0_outputs[707]) | (layer0_outputs[287]));
    assign layer1_outputs[1196] = (layer0_outputs[2144]) & ~(layer0_outputs[359]);
    assign layer1_outputs[1197] = (layer0_outputs[747]) & (layer0_outputs[2076]);
    assign layer1_outputs[1198] = (layer0_outputs[1641]) & (layer0_outputs[453]);
    assign layer1_outputs[1199] = (layer0_outputs[528]) & ~(layer0_outputs[1577]);
    assign layer1_outputs[1200] = (layer0_outputs[431]) | (layer0_outputs[61]);
    assign layer1_outputs[1201] = (layer0_outputs[2363]) & ~(layer0_outputs[932]);
    assign layer1_outputs[1202] = layer0_outputs[1447];
    assign layer1_outputs[1203] = (layer0_outputs[174]) | (layer0_outputs[1521]);
    assign layer1_outputs[1204] = (layer0_outputs[920]) & ~(layer0_outputs[1498]);
    assign layer1_outputs[1205] = (layer0_outputs[267]) & (layer0_outputs[2466]);
    assign layer1_outputs[1206] = (layer0_outputs[288]) & (layer0_outputs[1183]);
    assign layer1_outputs[1207] = ~(layer0_outputs[860]) | (layer0_outputs[2277]);
    assign layer1_outputs[1208] = ~(layer0_outputs[1361]);
    assign layer1_outputs[1209] = ~((layer0_outputs[536]) & (layer0_outputs[2552]));
    assign layer1_outputs[1210] = ~(layer0_outputs[99]);
    assign layer1_outputs[1211] = ~(layer0_outputs[1361]);
    assign layer1_outputs[1212] = ~(layer0_outputs[2064]) | (layer0_outputs[1950]);
    assign layer1_outputs[1213] = 1'b0;
    assign layer1_outputs[1214] = ~(layer0_outputs[411]) | (layer0_outputs[71]);
    assign layer1_outputs[1215] = ~((layer0_outputs[884]) ^ (layer0_outputs[1900]));
    assign layer1_outputs[1216] = (layer0_outputs[584]) | (layer0_outputs[344]);
    assign layer1_outputs[1217] = ~((layer0_outputs[1120]) ^ (layer0_outputs[386]));
    assign layer1_outputs[1218] = 1'b0;
    assign layer1_outputs[1219] = (layer0_outputs[2253]) & ~(layer0_outputs[1608]);
    assign layer1_outputs[1220] = ~(layer0_outputs[32]) | (layer0_outputs[534]);
    assign layer1_outputs[1221] = ~(layer0_outputs[2364]) | (layer0_outputs[1826]);
    assign layer1_outputs[1222] = ~(layer0_outputs[2117]);
    assign layer1_outputs[1223] = (layer0_outputs[1973]) & (layer0_outputs[286]);
    assign layer1_outputs[1224] = 1'b1;
    assign layer1_outputs[1225] = layer0_outputs[2243];
    assign layer1_outputs[1226] = (layer0_outputs[515]) & ~(layer0_outputs[791]);
    assign layer1_outputs[1227] = ~(layer0_outputs[2455]) | (layer0_outputs[2549]);
    assign layer1_outputs[1228] = ~(layer0_outputs[649]);
    assign layer1_outputs[1229] = ~((layer0_outputs[344]) ^ (layer0_outputs[206]));
    assign layer1_outputs[1230] = (layer0_outputs[729]) & ~(layer0_outputs[1638]);
    assign layer1_outputs[1231] = layer0_outputs[1913];
    assign layer1_outputs[1232] = ~((layer0_outputs[1567]) | (layer0_outputs[1427]));
    assign layer1_outputs[1233] = 1'b0;
    assign layer1_outputs[1234] = (layer0_outputs[711]) & ~(layer0_outputs[1901]);
    assign layer1_outputs[1235] = (layer0_outputs[328]) & ~(layer0_outputs[817]);
    assign layer1_outputs[1236] = (layer0_outputs[1365]) & ~(layer0_outputs[824]);
    assign layer1_outputs[1237] = ~(layer0_outputs[2067]);
    assign layer1_outputs[1238] = ~(layer0_outputs[2480]);
    assign layer1_outputs[1239] = ~(layer0_outputs[1139]);
    assign layer1_outputs[1240] = layer0_outputs[2511];
    assign layer1_outputs[1241] = (layer0_outputs[1471]) & ~(layer0_outputs[1051]);
    assign layer1_outputs[1242] = ~(layer0_outputs[2051]) | (layer0_outputs[84]);
    assign layer1_outputs[1243] = layer0_outputs[1549];
    assign layer1_outputs[1244] = ~(layer0_outputs[301]);
    assign layer1_outputs[1245] = layer0_outputs[262];
    assign layer1_outputs[1246] = (layer0_outputs[500]) ^ (layer0_outputs[568]);
    assign layer1_outputs[1247] = ~(layer0_outputs[2031]) | (layer0_outputs[590]);
    assign layer1_outputs[1248] = layer0_outputs[2335];
    assign layer1_outputs[1249] = (layer0_outputs[990]) | (layer0_outputs[1883]);
    assign layer1_outputs[1250] = (layer0_outputs[840]) & ~(layer0_outputs[379]);
    assign layer1_outputs[1251] = 1'b1;
    assign layer1_outputs[1252] = ~(layer0_outputs[1817]) | (layer0_outputs[1268]);
    assign layer1_outputs[1253] = ~((layer0_outputs[2020]) | (layer0_outputs[559]));
    assign layer1_outputs[1254] = (layer0_outputs[2258]) & (layer0_outputs[2348]);
    assign layer1_outputs[1255] = (layer0_outputs[1884]) & ~(layer0_outputs[2100]);
    assign layer1_outputs[1256] = ~(layer0_outputs[726]) | (layer0_outputs[209]);
    assign layer1_outputs[1257] = 1'b1;
    assign layer1_outputs[1258] = (layer0_outputs[638]) & ~(layer0_outputs[892]);
    assign layer1_outputs[1259] = ~((layer0_outputs[2231]) & (layer0_outputs[1289]));
    assign layer1_outputs[1260] = ~(layer0_outputs[135]) | (layer0_outputs[987]);
    assign layer1_outputs[1261] = ~(layer0_outputs[1981]) | (layer0_outputs[173]);
    assign layer1_outputs[1262] = ~(layer0_outputs[528]) | (layer0_outputs[460]);
    assign layer1_outputs[1263] = 1'b1;
    assign layer1_outputs[1264] = (layer0_outputs[2205]) & (layer0_outputs[2457]);
    assign layer1_outputs[1265] = (layer0_outputs[1666]) & (layer0_outputs[464]);
    assign layer1_outputs[1266] = ~(layer0_outputs[1698]) | (layer0_outputs[771]);
    assign layer1_outputs[1267] = layer0_outputs[475];
    assign layer1_outputs[1268] = 1'b0;
    assign layer1_outputs[1269] = ~(layer0_outputs[701]) | (layer0_outputs[1487]);
    assign layer1_outputs[1270] = ~(layer0_outputs[1277]);
    assign layer1_outputs[1271] = (layer0_outputs[1567]) | (layer0_outputs[1008]);
    assign layer1_outputs[1272] = ~(layer0_outputs[1910]);
    assign layer1_outputs[1273] = ~(layer0_outputs[1454]) | (layer0_outputs[792]);
    assign layer1_outputs[1274] = layer0_outputs[364];
    assign layer1_outputs[1275] = ~(layer0_outputs[2452]);
    assign layer1_outputs[1276] = 1'b1;
    assign layer1_outputs[1277] = (layer0_outputs[1236]) & ~(layer0_outputs[158]);
    assign layer1_outputs[1278] = ~((layer0_outputs[2521]) & (layer0_outputs[1169]));
    assign layer1_outputs[1279] = 1'b0;
    assign layer1_outputs[1280] = ~(layer0_outputs[1899]) | (layer0_outputs[1722]);
    assign layer1_outputs[1281] = ~((layer0_outputs[405]) ^ (layer0_outputs[768]));
    assign layer1_outputs[1282] = 1'b0;
    assign layer1_outputs[1283] = (layer0_outputs[2188]) & ~(layer0_outputs[641]);
    assign layer1_outputs[1284] = (layer0_outputs[1558]) | (layer0_outputs[1818]);
    assign layer1_outputs[1285] = (layer0_outputs[1231]) & (layer0_outputs[350]);
    assign layer1_outputs[1286] = ~((layer0_outputs[1050]) | (layer0_outputs[1074]));
    assign layer1_outputs[1287] = ~((layer0_outputs[857]) & (layer0_outputs[1477]));
    assign layer1_outputs[1288] = (layer0_outputs[1398]) | (layer0_outputs[2142]);
    assign layer1_outputs[1289] = 1'b0;
    assign layer1_outputs[1290] = ~((layer0_outputs[220]) | (layer0_outputs[2395]));
    assign layer1_outputs[1291] = ~((layer0_outputs[1204]) | (layer0_outputs[269]));
    assign layer1_outputs[1292] = ~(layer0_outputs[467]) | (layer0_outputs[1592]);
    assign layer1_outputs[1293] = ~((layer0_outputs[2439]) & (layer0_outputs[1249]));
    assign layer1_outputs[1294] = ~(layer0_outputs[1368]);
    assign layer1_outputs[1295] = ~(layer0_outputs[232]);
    assign layer1_outputs[1296] = ~((layer0_outputs[1311]) | (layer0_outputs[364]));
    assign layer1_outputs[1297] = ~(layer0_outputs[2296]);
    assign layer1_outputs[1298] = (layer0_outputs[701]) & ~(layer0_outputs[2464]);
    assign layer1_outputs[1299] = ~(layer0_outputs[2391]);
    assign layer1_outputs[1300] = 1'b0;
    assign layer1_outputs[1301] = ~((layer0_outputs[1506]) ^ (layer0_outputs[750]));
    assign layer1_outputs[1302] = ~(layer0_outputs[834]) | (layer0_outputs[617]);
    assign layer1_outputs[1303] = (layer0_outputs[129]) & ~(layer0_outputs[42]);
    assign layer1_outputs[1304] = 1'b0;
    assign layer1_outputs[1305] = 1'b1;
    assign layer1_outputs[1306] = ~(layer0_outputs[1875]) | (layer0_outputs[1061]);
    assign layer1_outputs[1307] = layer0_outputs[2499];
    assign layer1_outputs[1308] = ~((layer0_outputs[1164]) | (layer0_outputs[803]));
    assign layer1_outputs[1309] = (layer0_outputs[2305]) & ~(layer0_outputs[1507]);
    assign layer1_outputs[1310] = ~((layer0_outputs[2065]) & (layer0_outputs[2525]));
    assign layer1_outputs[1311] = (layer0_outputs[1812]) ^ (layer0_outputs[693]);
    assign layer1_outputs[1312] = ~(layer0_outputs[944]) | (layer0_outputs[1540]);
    assign layer1_outputs[1313] = ~((layer0_outputs[1474]) & (layer0_outputs[883]));
    assign layer1_outputs[1314] = ~((layer0_outputs[1995]) & (layer0_outputs[1707]));
    assign layer1_outputs[1315] = 1'b0;
    assign layer1_outputs[1316] = (layer0_outputs[1657]) & ~(layer0_outputs[2110]);
    assign layer1_outputs[1317] = ~((layer0_outputs[415]) ^ (layer0_outputs[1359]));
    assign layer1_outputs[1318] = ~(layer0_outputs[1986]) | (layer0_outputs[2202]);
    assign layer1_outputs[1319] = ~((layer0_outputs[2557]) | (layer0_outputs[1103]));
    assign layer1_outputs[1320] = ~((layer0_outputs[775]) & (layer0_outputs[201]));
    assign layer1_outputs[1321] = 1'b1;
    assign layer1_outputs[1322] = ~(layer0_outputs[977]) | (layer0_outputs[1240]);
    assign layer1_outputs[1323] = ~(layer0_outputs[67]) | (layer0_outputs[2133]);
    assign layer1_outputs[1324] = (layer0_outputs[1293]) & ~(layer0_outputs[1880]);
    assign layer1_outputs[1325] = layer0_outputs[835];
    assign layer1_outputs[1326] = ~(layer0_outputs[1607]) | (layer0_outputs[72]);
    assign layer1_outputs[1327] = ~(layer0_outputs[1744]);
    assign layer1_outputs[1328] = ~((layer0_outputs[493]) & (layer0_outputs[1692]));
    assign layer1_outputs[1329] = (layer0_outputs[1604]) | (layer0_outputs[205]);
    assign layer1_outputs[1330] = layer0_outputs[181];
    assign layer1_outputs[1331] = ~(layer0_outputs[580]) | (layer0_outputs[169]);
    assign layer1_outputs[1332] = ~(layer0_outputs[2196]) | (layer0_outputs[1195]);
    assign layer1_outputs[1333] = (layer0_outputs[526]) | (layer0_outputs[540]);
    assign layer1_outputs[1334] = ~(layer0_outputs[58]) | (layer0_outputs[1128]);
    assign layer1_outputs[1335] = layer0_outputs[1583];
    assign layer1_outputs[1336] = layer0_outputs[2105];
    assign layer1_outputs[1337] = (layer0_outputs[763]) & ~(layer0_outputs[1677]);
    assign layer1_outputs[1338] = layer0_outputs[160];
    assign layer1_outputs[1339] = (layer0_outputs[2012]) & ~(layer0_outputs[1304]);
    assign layer1_outputs[1340] = (layer0_outputs[402]) & (layer0_outputs[115]);
    assign layer1_outputs[1341] = (layer0_outputs[1171]) | (layer0_outputs[1060]);
    assign layer1_outputs[1342] = 1'b0;
    assign layer1_outputs[1343] = (layer0_outputs[800]) | (layer0_outputs[130]);
    assign layer1_outputs[1344] = ~(layer0_outputs[454]) | (layer0_outputs[2242]);
    assign layer1_outputs[1345] = ~(layer0_outputs[2197]);
    assign layer1_outputs[1346] = (layer0_outputs[2035]) & ~(layer0_outputs[1736]);
    assign layer1_outputs[1347] = (layer0_outputs[2256]) & (layer0_outputs[221]);
    assign layer1_outputs[1348] = ~(layer0_outputs[516]) | (layer0_outputs[1434]);
    assign layer1_outputs[1349] = ~((layer0_outputs[2224]) & (layer0_outputs[1201]));
    assign layer1_outputs[1350] = layer0_outputs[1840];
    assign layer1_outputs[1351] = ~((layer0_outputs[601]) & (layer0_outputs[1976]));
    assign layer1_outputs[1352] = (layer0_outputs[414]) & ~(layer0_outputs[1232]);
    assign layer1_outputs[1353] = (layer0_outputs[2168]) & (layer0_outputs[2136]);
    assign layer1_outputs[1354] = (layer0_outputs[1315]) | (layer0_outputs[797]);
    assign layer1_outputs[1355] = ~(layer0_outputs[1280]);
    assign layer1_outputs[1356] = (layer0_outputs[2359]) & ~(layer0_outputs[2137]);
    assign layer1_outputs[1357] = layer0_outputs[2380];
    assign layer1_outputs[1358] = (layer0_outputs[445]) & ~(layer0_outputs[916]);
    assign layer1_outputs[1359] = ~((layer0_outputs[1918]) & (layer0_outputs[2329]));
    assign layer1_outputs[1360] = (layer0_outputs[583]) & ~(layer0_outputs[568]);
    assign layer1_outputs[1361] = ~((layer0_outputs[274]) | (layer0_outputs[1010]));
    assign layer1_outputs[1362] = 1'b1;
    assign layer1_outputs[1363] = (layer0_outputs[1572]) ^ (layer0_outputs[1966]);
    assign layer1_outputs[1364] = ~(layer0_outputs[1416]) | (layer0_outputs[2127]);
    assign layer1_outputs[1365] = ~(layer0_outputs[900]);
    assign layer1_outputs[1366] = 1'b1;
    assign layer1_outputs[1367] = ~(layer0_outputs[2074]) | (layer0_outputs[280]);
    assign layer1_outputs[1368] = layer0_outputs[2547];
    assign layer1_outputs[1369] = ~((layer0_outputs[894]) & (layer0_outputs[2158]));
    assign layer1_outputs[1370] = ~(layer0_outputs[1671]);
    assign layer1_outputs[1371] = ~(layer0_outputs[1895]) | (layer0_outputs[438]);
    assign layer1_outputs[1372] = ~(layer0_outputs[2287]);
    assign layer1_outputs[1373] = 1'b0;
    assign layer1_outputs[1374] = (layer0_outputs[2333]) & ~(layer0_outputs[313]);
    assign layer1_outputs[1375] = ~(layer0_outputs[1402]) | (layer0_outputs[1565]);
    assign layer1_outputs[1376] = layer0_outputs[1078];
    assign layer1_outputs[1377] = ~((layer0_outputs[833]) | (layer0_outputs[432]));
    assign layer1_outputs[1378] = (layer0_outputs[1526]) & ~(layer0_outputs[2514]);
    assign layer1_outputs[1379] = 1'b0;
    assign layer1_outputs[1380] = (layer0_outputs[1086]) ^ (layer0_outputs[1819]);
    assign layer1_outputs[1381] = ~(layer0_outputs[1673]) | (layer0_outputs[337]);
    assign layer1_outputs[1382] = ~((layer0_outputs[424]) | (layer0_outputs[2134]));
    assign layer1_outputs[1383] = (layer0_outputs[1390]) & (layer0_outputs[471]);
    assign layer1_outputs[1384] = ~(layer0_outputs[629]);
    assign layer1_outputs[1385] = (layer0_outputs[1892]) & ~(layer0_outputs[973]);
    assign layer1_outputs[1386] = (layer0_outputs[2206]) & (layer0_outputs[2242]);
    assign layer1_outputs[1387] = layer0_outputs[147];
    assign layer1_outputs[1388] = (layer0_outputs[1831]) ^ (layer0_outputs[520]);
    assign layer1_outputs[1389] = layer0_outputs[1555];
    assign layer1_outputs[1390] = ~((layer0_outputs[2221]) & (layer0_outputs[1306]));
    assign layer1_outputs[1391] = layer0_outputs[995];
    assign layer1_outputs[1392] = (layer0_outputs[2375]) ^ (layer0_outputs[1530]);
    assign layer1_outputs[1393] = (layer0_outputs[103]) | (layer0_outputs[334]);
    assign layer1_outputs[1394] = layer0_outputs[116];
    assign layer1_outputs[1395] = ~(layer0_outputs[2304]) | (layer0_outputs[838]);
    assign layer1_outputs[1396] = 1'b0;
    assign layer1_outputs[1397] = layer0_outputs[1813];
    assign layer1_outputs[1398] = ~((layer0_outputs[2189]) & (layer0_outputs[1313]));
    assign layer1_outputs[1399] = (layer0_outputs[1390]) | (layer0_outputs[1541]);
    assign layer1_outputs[1400] = (layer0_outputs[598]) & (layer0_outputs[1450]);
    assign layer1_outputs[1401] = (layer0_outputs[696]) & ~(layer0_outputs[2449]);
    assign layer1_outputs[1402] = layer0_outputs[447];
    assign layer1_outputs[1403] = (layer0_outputs[1790]) & (layer0_outputs[605]);
    assign layer1_outputs[1404] = ~((layer0_outputs[1596]) ^ (layer0_outputs[2331]));
    assign layer1_outputs[1405] = ~((layer0_outputs[139]) & (layer0_outputs[1200]));
    assign layer1_outputs[1406] = (layer0_outputs[441]) ^ (layer0_outputs[981]);
    assign layer1_outputs[1407] = (layer0_outputs[217]) | (layer0_outputs[93]);
    assign layer1_outputs[1408] = (layer0_outputs[1737]) | (layer0_outputs[391]);
    assign layer1_outputs[1409] = layer0_outputs[320];
    assign layer1_outputs[1410] = (layer0_outputs[1011]) | (layer0_outputs[2420]);
    assign layer1_outputs[1411] = (layer0_outputs[2313]) | (layer0_outputs[1231]);
    assign layer1_outputs[1412] = (layer0_outputs[2106]) & ~(layer0_outputs[518]);
    assign layer1_outputs[1413] = 1'b1;
    assign layer1_outputs[1414] = ~((layer0_outputs[759]) ^ (layer0_outputs[40]));
    assign layer1_outputs[1415] = ~(layer0_outputs[695]) | (layer0_outputs[1412]);
    assign layer1_outputs[1416] = ~((layer0_outputs[770]) & (layer0_outputs[2131]));
    assign layer1_outputs[1417] = layer0_outputs[333];
    assign layer1_outputs[1418] = (layer0_outputs[1143]) & ~(layer0_outputs[236]);
    assign layer1_outputs[1419] = 1'b0;
    assign layer1_outputs[1420] = layer0_outputs[2511];
    assign layer1_outputs[1421] = ~((layer0_outputs[1974]) ^ (layer0_outputs[2264]));
    assign layer1_outputs[1422] = layer0_outputs[1085];
    assign layer1_outputs[1423] = ~(layer0_outputs[2410]) | (layer0_outputs[787]);
    assign layer1_outputs[1424] = layer0_outputs[109];
    assign layer1_outputs[1425] = 1'b1;
    assign layer1_outputs[1426] = (layer0_outputs[2355]) | (layer0_outputs[2209]);
    assign layer1_outputs[1427] = (layer0_outputs[1515]) & ~(layer0_outputs[1469]);
    assign layer1_outputs[1428] = layer0_outputs[486];
    assign layer1_outputs[1429] = ~(layer0_outputs[2386]);
    assign layer1_outputs[1430] = (layer0_outputs[1399]) & ~(layer0_outputs[2533]);
    assign layer1_outputs[1431] = ~(layer0_outputs[842]);
    assign layer1_outputs[1432] = ~(layer0_outputs[1179]);
    assign layer1_outputs[1433] = ~(layer0_outputs[413]);
    assign layer1_outputs[1434] = (layer0_outputs[2491]) & ~(layer0_outputs[707]);
    assign layer1_outputs[1435] = (layer0_outputs[1276]) & (layer0_outputs[1020]);
    assign layer1_outputs[1436] = (layer0_outputs[1173]) & ~(layer0_outputs[2126]);
    assign layer1_outputs[1437] = ~((layer0_outputs[1449]) & (layer0_outputs[1057]));
    assign layer1_outputs[1438] = ~(layer0_outputs[1590]) | (layer0_outputs[2304]);
    assign layer1_outputs[1439] = ~((layer0_outputs[173]) & (layer0_outputs[1108]));
    assign layer1_outputs[1440] = ~(layer0_outputs[255]) | (layer0_outputs[1188]);
    assign layer1_outputs[1441] = 1'b0;
    assign layer1_outputs[1442] = (layer0_outputs[1247]) & ~(layer0_outputs[1758]);
    assign layer1_outputs[1443] = ~((layer0_outputs[2037]) | (layer0_outputs[2207]));
    assign layer1_outputs[1444] = layer0_outputs[403];
    assign layer1_outputs[1445] = ~((layer0_outputs[925]) & (layer0_outputs[554]));
    assign layer1_outputs[1446] = (layer0_outputs[922]) & (layer0_outputs[136]);
    assign layer1_outputs[1447] = (layer0_outputs[949]) ^ (layer0_outputs[1343]);
    assign layer1_outputs[1448] = layer0_outputs[1909];
    assign layer1_outputs[1449] = (layer0_outputs[1886]) ^ (layer0_outputs[1353]);
    assign layer1_outputs[1450] = ~((layer0_outputs[223]) | (layer0_outputs[314]));
    assign layer1_outputs[1451] = ~(layer0_outputs[647]) | (layer0_outputs[955]);
    assign layer1_outputs[1452] = ~((layer0_outputs[1019]) | (layer0_outputs[1249]));
    assign layer1_outputs[1453] = (layer0_outputs[2013]) | (layer0_outputs[2466]);
    assign layer1_outputs[1454] = ~(layer0_outputs[1857]) | (layer0_outputs[2407]);
    assign layer1_outputs[1455] = 1'b1;
    assign layer1_outputs[1456] = (layer0_outputs[2301]) & ~(layer0_outputs[978]);
    assign layer1_outputs[1457] = ~(layer0_outputs[1115]) | (layer0_outputs[650]);
    assign layer1_outputs[1458] = (layer0_outputs[369]) & (layer0_outputs[1968]);
    assign layer1_outputs[1459] = ~((layer0_outputs[1861]) | (layer0_outputs[1522]));
    assign layer1_outputs[1460] = (layer0_outputs[2207]) | (layer0_outputs[1954]);
    assign layer1_outputs[1461] = ~((layer0_outputs[723]) & (layer0_outputs[2498]));
    assign layer1_outputs[1462] = ~(layer0_outputs[588]) | (layer0_outputs[929]);
    assign layer1_outputs[1463] = ~(layer0_outputs[1854]) | (layer0_outputs[614]);
    assign layer1_outputs[1464] = ~(layer0_outputs[18]);
    assign layer1_outputs[1465] = 1'b0;
    assign layer1_outputs[1466] = ~((layer0_outputs[1338]) ^ (layer0_outputs[640]));
    assign layer1_outputs[1467] = layer0_outputs[2192];
    assign layer1_outputs[1468] = ~(layer0_outputs[2475]);
    assign layer1_outputs[1469] = (layer0_outputs[152]) | (layer0_outputs[1889]);
    assign layer1_outputs[1470] = (layer0_outputs[1207]) | (layer0_outputs[283]);
    assign layer1_outputs[1471] = ~(layer0_outputs[126]);
    assign layer1_outputs[1472] = ~((layer0_outputs[53]) & (layer0_outputs[30]));
    assign layer1_outputs[1473] = (layer0_outputs[1842]) ^ (layer0_outputs[1540]);
    assign layer1_outputs[1474] = 1'b1;
    assign layer1_outputs[1475] = layer0_outputs[1856];
    assign layer1_outputs[1476] = ~(layer0_outputs[1784]);
    assign layer1_outputs[1477] = ~((layer0_outputs[316]) ^ (layer0_outputs[375]));
    assign layer1_outputs[1478] = 1'b0;
    assign layer1_outputs[1479] = ~(layer0_outputs[1433]) | (layer0_outputs[1794]);
    assign layer1_outputs[1480] = ~(layer0_outputs[316]) | (layer0_outputs[1539]);
    assign layer1_outputs[1481] = ~(layer0_outputs[106]) | (layer0_outputs[34]);
    assign layer1_outputs[1482] = 1'b0;
    assign layer1_outputs[1483] = ~(layer0_outputs[2373]) | (layer0_outputs[738]);
    assign layer1_outputs[1484] = layer0_outputs[2425];
    assign layer1_outputs[1485] = (layer0_outputs[2020]) & ~(layer0_outputs[600]);
    assign layer1_outputs[1486] = ~(layer0_outputs[844]) | (layer0_outputs[1711]);
    assign layer1_outputs[1487] = layer0_outputs[1769];
    assign layer1_outputs[1488] = ~(layer0_outputs[1851]) | (layer0_outputs[2216]);
    assign layer1_outputs[1489] = (layer0_outputs[1906]) & ~(layer0_outputs[577]);
    assign layer1_outputs[1490] = (layer0_outputs[60]) | (layer0_outputs[619]);
    assign layer1_outputs[1491] = 1'b1;
    assign layer1_outputs[1492] = layer0_outputs[888];
    assign layer1_outputs[1493] = 1'b0;
    assign layer1_outputs[1494] = ~(layer0_outputs[1395]) | (layer0_outputs[1173]);
    assign layer1_outputs[1495] = ~((layer0_outputs[545]) & (layer0_outputs[1115]));
    assign layer1_outputs[1496] = ~((layer0_outputs[318]) | (layer0_outputs[1997]));
    assign layer1_outputs[1497] = (layer0_outputs[2534]) & ~(layer0_outputs[163]);
    assign layer1_outputs[1498] = ~(layer0_outputs[62]) | (layer0_outputs[988]);
    assign layer1_outputs[1499] = 1'b1;
    assign layer1_outputs[1500] = ~(layer0_outputs[1037]) | (layer0_outputs[1198]);
    assign layer1_outputs[1501] = ~(layer0_outputs[1394]);
    assign layer1_outputs[1502] = layer0_outputs[2063];
    assign layer1_outputs[1503] = (layer0_outputs[323]) & ~(layer0_outputs[1023]);
    assign layer1_outputs[1504] = (layer0_outputs[2145]) & ~(layer0_outputs[472]);
    assign layer1_outputs[1505] = layer0_outputs[6];
    assign layer1_outputs[1506] = (layer0_outputs[1556]) & ~(layer0_outputs[2288]);
    assign layer1_outputs[1507] = 1'b0;
    assign layer1_outputs[1508] = 1'b1;
    assign layer1_outputs[1509] = ~((layer0_outputs[1769]) & (layer0_outputs[1468]));
    assign layer1_outputs[1510] = ~((layer0_outputs[2211]) ^ (layer0_outputs[2378]));
    assign layer1_outputs[1511] = layer0_outputs[1378];
    assign layer1_outputs[1512] = ~(layer0_outputs[644]);
    assign layer1_outputs[1513] = (layer0_outputs[2085]) ^ (layer0_outputs[1237]);
    assign layer1_outputs[1514] = (layer0_outputs[2212]) & ~(layer0_outputs[1722]);
    assign layer1_outputs[1515] = ~(layer0_outputs[2083]) | (layer0_outputs[425]);
    assign layer1_outputs[1516] = layer0_outputs[1309];
    assign layer1_outputs[1517] = ~(layer0_outputs[2502]);
    assign layer1_outputs[1518] = ~(layer0_outputs[2295]) | (layer0_outputs[918]);
    assign layer1_outputs[1519] = ~((layer0_outputs[978]) | (layer0_outputs[1106]));
    assign layer1_outputs[1520] = (layer0_outputs[1720]) & ~(layer0_outputs[2222]);
    assign layer1_outputs[1521] = (layer0_outputs[2449]) & ~(layer0_outputs[470]);
    assign layer1_outputs[1522] = layer0_outputs[1668];
    assign layer1_outputs[1523] = ~((layer0_outputs[2178]) | (layer0_outputs[1235]));
    assign layer1_outputs[1524] = (layer0_outputs[2555]) & ~(layer0_outputs[1534]);
    assign layer1_outputs[1525] = 1'b0;
    assign layer1_outputs[1526] = layer0_outputs[305];
    assign layer1_outputs[1527] = ~(layer0_outputs[266]) | (layer0_outputs[2250]);
    assign layer1_outputs[1528] = 1'b0;
    assign layer1_outputs[1529] = (layer0_outputs[2389]) ^ (layer0_outputs[1459]);
    assign layer1_outputs[1530] = ~((layer0_outputs[1832]) ^ (layer0_outputs[1230]));
    assign layer1_outputs[1531] = ~(layer0_outputs[137]) | (layer0_outputs[1132]);
    assign layer1_outputs[1532] = ~((layer0_outputs[11]) & (layer0_outputs[232]));
    assign layer1_outputs[1533] = ~((layer0_outputs[2474]) & (layer0_outputs[1268]));
    assign layer1_outputs[1534] = (layer0_outputs[881]) & (layer0_outputs[1236]);
    assign layer1_outputs[1535] = (layer0_outputs[2399]) & ~(layer0_outputs[413]);
    assign layer1_outputs[1536] = ~((layer0_outputs[1182]) & (layer0_outputs[855]));
    assign layer1_outputs[1537] = (layer0_outputs[410]) & ~(layer0_outputs[966]);
    assign layer1_outputs[1538] = ~(layer0_outputs[2364]) | (layer0_outputs[1296]);
    assign layer1_outputs[1539] = 1'b0;
    assign layer1_outputs[1540] = (layer0_outputs[204]) & ~(layer0_outputs[2]);
    assign layer1_outputs[1541] = ~(layer0_outputs[176]) | (layer0_outputs[1868]);
    assign layer1_outputs[1542] = ~(layer0_outputs[1289]);
    assign layer1_outputs[1543] = ~((layer0_outputs[200]) | (layer0_outputs[2179]));
    assign layer1_outputs[1544] = ~((layer0_outputs[82]) ^ (layer0_outputs[2152]));
    assign layer1_outputs[1545] = ~(layer0_outputs[111]);
    assign layer1_outputs[1546] = 1'b1;
    assign layer1_outputs[1547] = layer0_outputs[1418];
    assign layer1_outputs[1548] = (layer0_outputs[850]) & ~(layer0_outputs[1198]);
    assign layer1_outputs[1549] = ~(layer0_outputs[1052]) | (layer0_outputs[2416]);
    assign layer1_outputs[1550] = 1'b1;
    assign layer1_outputs[1551] = ~(layer0_outputs[1753]) | (layer0_outputs[2018]);
    assign layer1_outputs[1552] = (layer0_outputs[1135]) & ~(layer0_outputs[127]);
    assign layer1_outputs[1553] = (layer0_outputs[1419]) & ~(layer0_outputs[1465]);
    assign layer1_outputs[1554] = layer0_outputs[1125];
    assign layer1_outputs[1555] = 1'b1;
    assign layer1_outputs[1556] = layer0_outputs[302];
    assign layer1_outputs[1557] = ~((layer0_outputs[1329]) & (layer0_outputs[905]));
    assign layer1_outputs[1558] = layer0_outputs[1392];
    assign layer1_outputs[1559] = (layer0_outputs[121]) | (layer0_outputs[1400]);
    assign layer1_outputs[1560] = ~(layer0_outputs[2161]) | (layer0_outputs[1503]);
    assign layer1_outputs[1561] = 1'b0;
    assign layer1_outputs[1562] = ~((layer0_outputs[1688]) & (layer0_outputs[46]));
    assign layer1_outputs[1563] = ~((layer0_outputs[2413]) | (layer0_outputs[1767]));
    assign layer1_outputs[1564] = (layer0_outputs[2321]) & (layer0_outputs[1665]);
    assign layer1_outputs[1565] = layer0_outputs[794];
    assign layer1_outputs[1566] = (layer0_outputs[1763]) | (layer0_outputs[1853]);
    assign layer1_outputs[1567] = (layer0_outputs[2043]) | (layer0_outputs[2043]);
    assign layer1_outputs[1568] = ~(layer0_outputs[2171]) | (layer0_outputs[550]);
    assign layer1_outputs[1569] = ~(layer0_outputs[2101]) | (layer0_outputs[133]);
    assign layer1_outputs[1570] = ~((layer0_outputs[2453]) ^ (layer0_outputs[1690]));
    assign layer1_outputs[1571] = (layer0_outputs[1474]) & ~(layer0_outputs[806]);
    assign layer1_outputs[1572] = layer0_outputs[812];
    assign layer1_outputs[1573] = 1'b0;
    assign layer1_outputs[1574] = (layer0_outputs[241]) & ~(layer0_outputs[989]);
    assign layer1_outputs[1575] = layer0_outputs[857];
    assign layer1_outputs[1576] = 1'b0;
    assign layer1_outputs[1577] = ~(layer0_outputs[511]);
    assign layer1_outputs[1578] = layer0_outputs[645];
    assign layer1_outputs[1579] = ~((layer0_outputs[50]) ^ (layer0_outputs[1643]));
    assign layer1_outputs[1580] = layer0_outputs[690];
    assign layer1_outputs[1581] = ~(layer0_outputs[1303]);
    assign layer1_outputs[1582] = (layer0_outputs[247]) & ~(layer0_outputs[1668]);
    assign layer1_outputs[1583] = layer0_outputs[480];
    assign layer1_outputs[1584] = ~((layer0_outputs[1798]) & (layer0_outputs[1488]));
    assign layer1_outputs[1585] = 1'b0;
    assign layer1_outputs[1586] = ~(layer0_outputs[230]) | (layer0_outputs[2069]);
    assign layer1_outputs[1587] = ~(layer0_outputs[340]) | (layer0_outputs[2388]);
    assign layer1_outputs[1588] = (layer0_outputs[606]) & ~(layer0_outputs[420]);
    assign layer1_outputs[1589] = ~((layer0_outputs[2252]) | (layer0_outputs[1805]));
    assign layer1_outputs[1590] = 1'b1;
    assign layer1_outputs[1591] = (layer0_outputs[167]) & ~(layer0_outputs[1990]);
    assign layer1_outputs[1592] = layer0_outputs[783];
    assign layer1_outputs[1593] = layer0_outputs[2433];
    assign layer1_outputs[1594] = (layer0_outputs[2311]) | (layer0_outputs[1728]);
    assign layer1_outputs[1595] = 1'b0;
    assign layer1_outputs[1596] = 1'b1;
    assign layer1_outputs[1597] = (layer0_outputs[1168]) & ~(layer0_outputs[1606]);
    assign layer1_outputs[1598] = ~((layer0_outputs[2044]) | (layer0_outputs[2366]));
    assign layer1_outputs[1599] = (layer0_outputs[193]) | (layer0_outputs[1471]);
    assign layer1_outputs[1600] = (layer0_outputs[2241]) & (layer0_outputs[2325]);
    assign layer1_outputs[1601] = 1'b0;
    assign layer1_outputs[1602] = layer0_outputs[2329];
    assign layer1_outputs[1603] = layer0_outputs[1686];
    assign layer1_outputs[1604] = layer0_outputs[755];
    assign layer1_outputs[1605] = 1'b1;
    assign layer1_outputs[1606] = (layer0_outputs[1138]) & ~(layer0_outputs[1557]);
    assign layer1_outputs[1607] = ~(layer0_outputs[1196]) | (layer0_outputs[59]);
    assign layer1_outputs[1608] = (layer0_outputs[172]) & ~(layer0_outputs[1832]);
    assign layer1_outputs[1609] = ~(layer0_outputs[2303]) | (layer0_outputs[1948]);
    assign layer1_outputs[1610] = layer0_outputs[1686];
    assign layer1_outputs[1611] = ~(layer0_outputs[776]) | (layer0_outputs[1149]);
    assign layer1_outputs[1612] = (layer0_outputs[507]) | (layer0_outputs[2008]);
    assign layer1_outputs[1613] = ~(layer0_outputs[2135]);
    assign layer1_outputs[1614] = layer0_outputs[2104];
    assign layer1_outputs[1615] = ~((layer0_outputs[969]) | (layer0_outputs[2199]));
    assign layer1_outputs[1616] = layer0_outputs[1490];
    assign layer1_outputs[1617] = 1'b1;
    assign layer1_outputs[1618] = ~(layer0_outputs[197]) | (layer0_outputs[1867]);
    assign layer1_outputs[1619] = layer0_outputs[2442];
    assign layer1_outputs[1620] = ~(layer0_outputs[2507]) | (layer0_outputs[837]);
    assign layer1_outputs[1621] = layer0_outputs[504];
    assign layer1_outputs[1622] = ~((layer0_outputs[2103]) | (layer0_outputs[2091]));
    assign layer1_outputs[1623] = layer0_outputs[839];
    assign layer1_outputs[1624] = ~((layer0_outputs[1649]) & (layer0_outputs[1749]));
    assign layer1_outputs[1625] = ~(layer0_outputs[1482]);
    assign layer1_outputs[1626] = (layer0_outputs[507]) & (layer0_outputs[200]);
    assign layer1_outputs[1627] = ~(layer0_outputs[1409]) | (layer0_outputs[243]);
    assign layer1_outputs[1628] = ~(layer0_outputs[756]);
    assign layer1_outputs[1629] = ~(layer0_outputs[2193]) | (layer0_outputs[879]);
    assign layer1_outputs[1630] = ~((layer0_outputs[433]) ^ (layer0_outputs[2306]));
    assign layer1_outputs[1631] = (layer0_outputs[1430]) & (layer0_outputs[1927]);
    assign layer1_outputs[1632] = (layer0_outputs[43]) & ~(layer0_outputs[65]);
    assign layer1_outputs[1633] = (layer0_outputs[168]) ^ (layer0_outputs[1026]);
    assign layer1_outputs[1634] = layer0_outputs[2004];
    assign layer1_outputs[1635] = (layer0_outputs[367]) & ~(layer0_outputs[1994]);
    assign layer1_outputs[1636] = (layer0_outputs[2545]) ^ (layer0_outputs[1923]);
    assign layer1_outputs[1637] = ~(layer0_outputs[147]);
    assign layer1_outputs[1638] = layer0_outputs[731];
    assign layer1_outputs[1639] = (layer0_outputs[1288]) & ~(layer0_outputs[779]);
    assign layer1_outputs[1640] = 1'b0;
    assign layer1_outputs[1641] = (layer0_outputs[229]) ^ (layer0_outputs[495]);
    assign layer1_outputs[1642] = ~(layer0_outputs[625]);
    assign layer1_outputs[1643] = 1'b1;
    assign layer1_outputs[1644] = (layer0_outputs[1070]) | (layer0_outputs[825]);
    assign layer1_outputs[1645] = (layer0_outputs[1475]) & (layer0_outputs[885]);
    assign layer1_outputs[1646] = layer0_outputs[2540];
    assign layer1_outputs[1647] = ~(layer0_outputs[362]);
    assign layer1_outputs[1648] = layer0_outputs[678];
    assign layer1_outputs[1649] = (layer0_outputs[9]) & ~(layer0_outputs[55]);
    assign layer1_outputs[1650] = layer0_outputs[1199];
    assign layer1_outputs[1651] = (layer0_outputs[1302]) & (layer0_outputs[1573]);
    assign layer1_outputs[1652] = ~(layer0_outputs[1469]) | (layer0_outputs[585]);
    assign layer1_outputs[1653] = layer0_outputs[520];
    assign layer1_outputs[1654] = ~(layer0_outputs[1475]);
    assign layer1_outputs[1655] = layer0_outputs[531];
    assign layer1_outputs[1656] = ~((layer0_outputs[1229]) & (layer0_outputs[728]));
    assign layer1_outputs[1657] = ~(layer0_outputs[2183]);
    assign layer1_outputs[1658] = 1'b1;
    assign layer1_outputs[1659] = 1'b0;
    assign layer1_outputs[1660] = ~(layer0_outputs[1631]);
    assign layer1_outputs[1661] = ~((layer0_outputs[945]) & (layer0_outputs[790]));
    assign layer1_outputs[1662] = layer0_outputs[1651];
    assign layer1_outputs[1663] = ~((layer0_outputs[2263]) ^ (layer0_outputs[2496]));
    assign layer1_outputs[1664] = (layer0_outputs[1157]) & ~(layer0_outputs[2484]);
    assign layer1_outputs[1665] = (layer0_outputs[2212]) & (layer0_outputs[1267]);
    assign layer1_outputs[1666] = ~((layer0_outputs[2358]) | (layer0_outputs[617]));
    assign layer1_outputs[1667] = ~(layer0_outputs[559]) | (layer0_outputs[2009]);
    assign layer1_outputs[1668] = 1'b1;
    assign layer1_outputs[1669] = ~((layer0_outputs[16]) | (layer0_outputs[1339]));
    assign layer1_outputs[1670] = (layer0_outputs[2261]) | (layer0_outputs[1931]);
    assign layer1_outputs[1671] = (layer0_outputs[1491]) ^ (layer0_outputs[1977]);
    assign layer1_outputs[1672] = (layer0_outputs[1534]) | (layer0_outputs[1118]);
    assign layer1_outputs[1673] = (layer0_outputs[1593]) | (layer0_outputs[1843]);
    assign layer1_outputs[1674] = (layer0_outputs[445]) | (layer0_outputs[365]);
    assign layer1_outputs[1675] = ~(layer0_outputs[2468]);
    assign layer1_outputs[1676] = ~(layer0_outputs[1148]);
    assign layer1_outputs[1677] = (layer0_outputs[1330]) & ~(layer0_outputs[1357]);
    assign layer1_outputs[1678] = ~(layer0_outputs[596]) | (layer0_outputs[1193]);
    assign layer1_outputs[1679] = (layer0_outputs[1386]) & ~(layer0_outputs[1776]);
    assign layer1_outputs[1680] = (layer0_outputs[2230]) & (layer0_outputs[1476]);
    assign layer1_outputs[1681] = 1'b1;
    assign layer1_outputs[1682] = ~(layer0_outputs[1808]);
    assign layer1_outputs[1683] = (layer0_outputs[1222]) & ~(layer0_outputs[1282]);
    assign layer1_outputs[1684] = (layer0_outputs[1190]) | (layer0_outputs[908]);
    assign layer1_outputs[1685] = ~(layer0_outputs[2274]);
    assign layer1_outputs[1686] = ~(layer0_outputs[1275]);
    assign layer1_outputs[1687] = (layer0_outputs[668]) | (layer0_outputs[1445]);
    assign layer1_outputs[1688] = (layer0_outputs[1848]) ^ (layer0_outputs[1374]);
    assign layer1_outputs[1689] = 1'b0;
    assign layer1_outputs[1690] = layer0_outputs[206];
    assign layer1_outputs[1691] = layer0_outputs[1729];
    assign layer1_outputs[1692] = layer0_outputs[715];
    assign layer1_outputs[1693] = ~((layer0_outputs[1531]) & (layer0_outputs[1291]));
    assign layer1_outputs[1694] = layer0_outputs[715];
    assign layer1_outputs[1695] = (layer0_outputs[2182]) & ~(layer0_outputs[1382]);
    assign layer1_outputs[1696] = layer0_outputs[609];
    assign layer1_outputs[1697] = ~((layer0_outputs[1962]) & (layer0_outputs[1411]));
    assign layer1_outputs[1698] = ~(layer0_outputs[2099]) | (layer0_outputs[302]);
    assign layer1_outputs[1699] = ~(layer0_outputs[2542]) | (layer0_outputs[851]);
    assign layer1_outputs[1700] = 1'b1;
    assign layer1_outputs[1701] = ~(layer0_outputs[2199]) | (layer0_outputs[840]);
    assign layer1_outputs[1702] = ~(layer0_outputs[1537]) | (layer0_outputs[699]);
    assign layer1_outputs[1703] = (layer0_outputs[820]) & (layer0_outputs[1849]);
    assign layer1_outputs[1704] = 1'b0;
    assign layer1_outputs[1705] = (layer0_outputs[1604]) & ~(layer0_outputs[18]);
    assign layer1_outputs[1706] = 1'b1;
    assign layer1_outputs[1707] = (layer0_outputs[1870]) & (layer0_outputs[380]);
    assign layer1_outputs[1708] = layer0_outputs[935];
    assign layer1_outputs[1709] = ~(layer0_outputs[1461]);
    assign layer1_outputs[1710] = ~((layer0_outputs[2334]) | (layer0_outputs[1488]));
    assign layer1_outputs[1711] = ~((layer0_outputs[1919]) | (layer0_outputs[263]));
    assign layer1_outputs[1712] = ~(layer0_outputs[1202]) | (layer0_outputs[2413]);
    assign layer1_outputs[1713] = ~(layer0_outputs[281]) | (layer0_outputs[558]);
    assign layer1_outputs[1714] = ~(layer0_outputs[664]) | (layer0_outputs[1358]);
    assign layer1_outputs[1715] = layer0_outputs[2354];
    assign layer1_outputs[1716] = ~((layer0_outputs[1597]) & (layer0_outputs[1256]));
    assign layer1_outputs[1717] = layer0_outputs[1719];
    assign layer1_outputs[1718] = 1'b0;
    assign layer1_outputs[1719] = ~(layer0_outputs[2226]);
    assign layer1_outputs[1720] = 1'b0;
    assign layer1_outputs[1721] = layer0_outputs[2002];
    assign layer1_outputs[1722] = layer0_outputs[674];
    assign layer1_outputs[1723] = ~(layer0_outputs[1369]) | (layer0_outputs[1213]);
    assign layer1_outputs[1724] = ~(layer0_outputs[165]);
    assign layer1_outputs[1725] = ~(layer0_outputs[450]) | (layer0_outputs[383]);
    assign layer1_outputs[1726] = 1'b0;
    assign layer1_outputs[1727] = (layer0_outputs[897]) & (layer0_outputs[2558]);
    assign layer1_outputs[1728] = ~(layer0_outputs[1819]);
    assign layer1_outputs[1729] = 1'b1;
    assign layer1_outputs[1730] = ~((layer0_outputs[1437]) & (layer0_outputs[937]));
    assign layer1_outputs[1731] = (layer0_outputs[1821]) | (layer0_outputs[433]);
    assign layer1_outputs[1732] = ~(layer0_outputs[2011]);
    assign layer1_outputs[1733] = 1'b1;
    assign layer1_outputs[1734] = (layer0_outputs[2248]) & ~(layer0_outputs[1044]);
    assign layer1_outputs[1735] = ~(layer0_outputs[137]) | (layer0_outputs[161]);
    assign layer1_outputs[1736] = ~((layer0_outputs[773]) ^ (layer0_outputs[1228]));
    assign layer1_outputs[1737] = ~(layer0_outputs[694]);
    assign layer1_outputs[1738] = ~((layer0_outputs[1136]) | (layer0_outputs[798]));
    assign layer1_outputs[1739] = 1'b1;
    assign layer1_outputs[1740] = (layer0_outputs[456]) ^ (layer0_outputs[1886]);
    assign layer1_outputs[1741] = ~((layer0_outputs[1814]) | (layer0_outputs[281]));
    assign layer1_outputs[1742] = 1'b0;
    assign layer1_outputs[1743] = ~((layer0_outputs[718]) | (layer0_outputs[1305]));
    assign layer1_outputs[1744] = (layer0_outputs[1331]) & (layer0_outputs[2194]);
    assign layer1_outputs[1745] = (layer0_outputs[1690]) & ~(layer0_outputs[669]);
    assign layer1_outputs[1746] = layer0_outputs[486];
    assign layer1_outputs[1747] = ~((layer0_outputs[268]) & (layer0_outputs[1496]));
    assign layer1_outputs[1748] = (layer0_outputs[1929]) & ~(layer0_outputs[2472]);
    assign layer1_outputs[1749] = layer0_outputs[542];
    assign layer1_outputs[1750] = ~(layer0_outputs[865]);
    assign layer1_outputs[1751] = (layer0_outputs[1817]) | (layer0_outputs[1347]);
    assign layer1_outputs[1752] = (layer0_outputs[2146]) & ~(layer0_outputs[1058]);
    assign layer1_outputs[1753] = ~((layer0_outputs[1993]) & (layer0_outputs[307]));
    assign layer1_outputs[1754] = (layer0_outputs[1027]) & ~(layer0_outputs[42]);
    assign layer1_outputs[1755] = ~((layer0_outputs[1723]) & (layer0_outputs[1272]));
    assign layer1_outputs[1756] = (layer0_outputs[240]) & ~(layer0_outputs[768]);
    assign layer1_outputs[1757] = (layer0_outputs[1747]) ^ (layer0_outputs[490]);
    assign layer1_outputs[1758] = (layer0_outputs[2393]) & ~(layer0_outputs[1420]);
    assign layer1_outputs[1759] = layer0_outputs[1897];
    assign layer1_outputs[1760] = (layer0_outputs[1588]) | (layer0_outputs[2361]);
    assign layer1_outputs[1761] = (layer0_outputs[1553]) & ~(layer0_outputs[799]);
    assign layer1_outputs[1762] = (layer0_outputs[1473]) & ~(layer0_outputs[2420]);
    assign layer1_outputs[1763] = layer0_outputs[1872];
    assign layer1_outputs[1764] = ~(layer0_outputs[2371]);
    assign layer1_outputs[1765] = layer0_outputs[501];
    assign layer1_outputs[1766] = ~((layer0_outputs[1795]) & (layer0_outputs[713]));
    assign layer1_outputs[1767] = 1'b1;
    assign layer1_outputs[1768] = 1'b0;
    assign layer1_outputs[1769] = 1'b0;
    assign layer1_outputs[1770] = ~(layer0_outputs[348]);
    assign layer1_outputs[1771] = ~((layer0_outputs[1327]) | (layer0_outputs[184]));
    assign layer1_outputs[1772] = (layer0_outputs[2053]) & ~(layer0_outputs[1071]);
    assign layer1_outputs[1773] = layer0_outputs[1493];
    assign layer1_outputs[1774] = ~(layer0_outputs[102]) | (layer0_outputs[88]);
    assign layer1_outputs[1775] = ~(layer0_outputs[1454]) | (layer0_outputs[1566]);
    assign layer1_outputs[1776] = (layer0_outputs[2439]) & (layer0_outputs[586]);
    assign layer1_outputs[1777] = ~(layer0_outputs[817]) | (layer0_outputs[1606]);
    assign layer1_outputs[1778] = ~((layer0_outputs[887]) & (layer0_outputs[2407]));
    assign layer1_outputs[1779] = layer0_outputs[1081];
    assign layer1_outputs[1780] = ~(layer0_outputs[1654]) | (layer0_outputs[1096]);
    assign layer1_outputs[1781] = 1'b0;
    assign layer1_outputs[1782] = (layer0_outputs[392]) | (layer0_outputs[1305]);
    assign layer1_outputs[1783] = 1'b0;
    assign layer1_outputs[1784] = 1'b0;
    assign layer1_outputs[1785] = (layer0_outputs[2542]) & ~(layer0_outputs[1122]);
    assign layer1_outputs[1786] = ~((layer0_outputs[1102]) & (layer0_outputs[245]));
    assign layer1_outputs[1787] = (layer0_outputs[2291]) & ~(layer0_outputs[452]);
    assign layer1_outputs[1788] = ~(layer0_outputs[1146]) | (layer0_outputs[795]);
    assign layer1_outputs[1789] = layer0_outputs[1841];
    assign layer1_outputs[1790] = (layer0_outputs[1893]) & (layer0_outputs[31]);
    assign layer1_outputs[1791] = (layer0_outputs[396]) | (layer0_outputs[1888]);
    assign layer1_outputs[1792] = ~(layer0_outputs[2352]);
    assign layer1_outputs[1793] = ~((layer0_outputs[2428]) | (layer0_outputs[2072]));
    assign layer1_outputs[1794] = (layer0_outputs[2228]) & ~(layer0_outputs[1596]);
    assign layer1_outputs[1795] = layer0_outputs[805];
    assign layer1_outputs[1796] = ~(layer0_outputs[659]);
    assign layer1_outputs[1797] = (layer0_outputs[1667]) & ~(layer0_outputs[1746]);
    assign layer1_outputs[1798] = ~(layer0_outputs[1536]);
    assign layer1_outputs[1799] = (layer0_outputs[1683]) & (layer0_outputs[796]);
    assign layer1_outputs[1800] = layer0_outputs[62];
    assign layer1_outputs[1801] = ~(layer0_outputs[303]);
    assign layer1_outputs[1802] = (layer0_outputs[1142]) & (layer0_outputs[1701]);
    assign layer1_outputs[1803] = (layer0_outputs[1420]) | (layer0_outputs[112]);
    assign layer1_outputs[1804] = ~(layer0_outputs[1715]);
    assign layer1_outputs[1805] = ~(layer0_outputs[2237]);
    assign layer1_outputs[1806] = ~(layer0_outputs[393]) | (layer0_outputs[452]);
    assign layer1_outputs[1807] = layer0_outputs[1565];
    assign layer1_outputs[1808] = layer0_outputs[530];
    assign layer1_outputs[1809] = ~((layer0_outputs[1577]) ^ (layer0_outputs[1747]));
    assign layer1_outputs[1810] = (layer0_outputs[1959]) | (layer0_outputs[1443]);
    assign layer1_outputs[1811] = ~(layer0_outputs[1563]);
    assign layer1_outputs[1812] = ~(layer0_outputs[2044]) | (layer0_outputs[1432]);
    assign layer1_outputs[1813] = ~(layer0_outputs[1701]) | (layer0_outputs[1698]);
    assign layer1_outputs[1814] = ~(layer0_outputs[829]) | (layer0_outputs[2159]);
    assign layer1_outputs[1815] = ~(layer0_outputs[1147]) | (layer0_outputs[1574]);
    assign layer1_outputs[1816] = ~(layer0_outputs[888]) | (layer0_outputs[572]);
    assign layer1_outputs[1817] = layer0_outputs[1709];
    assign layer1_outputs[1818] = ~((layer0_outputs[1674]) & (layer0_outputs[933]));
    assign layer1_outputs[1819] = ~(layer0_outputs[2236]) | (layer0_outputs[1868]);
    assign layer1_outputs[1820] = 1'b0;
    assign layer1_outputs[1821] = ~(layer0_outputs[1932]);
    assign layer1_outputs[1822] = layer0_outputs[1444];
    assign layer1_outputs[1823] = ~((layer0_outputs[2030]) & (layer0_outputs[1724]));
    assign layer1_outputs[1824] = (layer0_outputs[2147]) & (layer0_outputs[1117]);
    assign layer1_outputs[1825] = layer0_outputs[1946];
    assign layer1_outputs[1826] = ~((layer0_outputs[959]) & (layer0_outputs[2050]));
    assign layer1_outputs[1827] = 1'b1;
    assign layer1_outputs[1828] = 1'b0;
    assign layer1_outputs[1829] = (layer0_outputs[1013]) & ~(layer0_outputs[2419]);
    assign layer1_outputs[1830] = ~((layer0_outputs[1587]) | (layer0_outputs[2206]));
    assign layer1_outputs[1831] = (layer0_outputs[1980]) & ~(layer0_outputs[2200]);
    assign layer1_outputs[1832] = (layer0_outputs[859]) | (layer0_outputs[427]);
    assign layer1_outputs[1833] = (layer0_outputs[1389]) & (layer0_outputs[1607]);
    assign layer1_outputs[1834] = ~(layer0_outputs[1735]);
    assign layer1_outputs[1835] = (layer0_outputs[1580]) & ~(layer0_outputs[1046]);
    assign layer1_outputs[1836] = layer0_outputs[312];
    assign layer1_outputs[1837] = 1'b0;
    assign layer1_outputs[1838] = ~(layer0_outputs[16]);
    assign layer1_outputs[1839] = layer0_outputs[279];
    assign layer1_outputs[1840] = ~((layer0_outputs[798]) | (layer0_outputs[2400]));
    assign layer1_outputs[1841] = (layer0_outputs[2316]) & ~(layer0_outputs[1097]);
    assign layer1_outputs[1842] = layer0_outputs[1847];
    assign layer1_outputs[1843] = (layer0_outputs[2506]) & ~(layer0_outputs[1986]);
    assign layer1_outputs[1844] = (layer0_outputs[2400]) | (layer0_outputs[940]);
    assign layer1_outputs[1845] = 1'b0;
    assign layer1_outputs[1846] = ~((layer0_outputs[1230]) & (layer0_outputs[614]));
    assign layer1_outputs[1847] = ~(layer0_outputs[905]);
    assign layer1_outputs[1848] = (layer0_outputs[1517]) & ~(layer0_outputs[2522]);
    assign layer1_outputs[1849] = ~(layer0_outputs[64]);
    assign layer1_outputs[1850] = ~((layer0_outputs[1750]) | (layer0_outputs[1599]));
    assign layer1_outputs[1851] = 1'b0;
    assign layer1_outputs[1852] = ~((layer0_outputs[1954]) & (layer0_outputs[167]));
    assign layer1_outputs[1853] = ~((layer0_outputs[587]) & (layer0_outputs[2423]));
    assign layer1_outputs[1854] = (layer0_outputs[1521]) & ~(layer0_outputs[2010]);
    assign layer1_outputs[1855] = (layer0_outputs[431]) | (layer0_outputs[71]);
    assign layer1_outputs[1856] = (layer0_outputs[54]) ^ (layer0_outputs[2032]);
    assign layer1_outputs[1857] = ~(layer0_outputs[1802]) | (layer0_outputs[1574]);
    assign layer1_outputs[1858] = ~((layer0_outputs[84]) & (layer0_outputs[1041]));
    assign layer1_outputs[1859] = layer0_outputs[1896];
    assign layer1_outputs[1860] = ~(layer0_outputs[1005]) | (layer0_outputs[641]);
    assign layer1_outputs[1861] = 1'b1;
    assign layer1_outputs[1862] = 1'b1;
    assign layer1_outputs[1863] = (layer0_outputs[1203]) | (layer0_outputs[1989]);
    assign layer1_outputs[1864] = (layer0_outputs[716]) ^ (layer0_outputs[2158]);
    assign layer1_outputs[1865] = (layer0_outputs[1829]) & ~(layer0_outputs[57]);
    assign layer1_outputs[1866] = layer0_outputs[1876];
    assign layer1_outputs[1867] = (layer0_outputs[2195]) | (layer0_outputs[2219]);
    assign layer1_outputs[1868] = 1'b0;
    assign layer1_outputs[1869] = ~(layer0_outputs[2401]);
    assign layer1_outputs[1870] = ~((layer0_outputs[2441]) & (layer0_outputs[891]));
    assign layer1_outputs[1871] = (layer0_outputs[1934]) & ~(layer0_outputs[2087]);
    assign layer1_outputs[1872] = ~(layer0_outputs[1699]);
    assign layer1_outputs[1873] = (layer0_outputs[2376]) | (layer0_outputs[1646]);
    assign layer1_outputs[1874] = ~((layer0_outputs[2334]) | (layer0_outputs[1252]));
    assign layer1_outputs[1875] = ~((layer0_outputs[2512]) & (layer0_outputs[1127]));
    assign layer1_outputs[1876] = (layer0_outputs[631]) | (layer0_outputs[886]);
    assign layer1_outputs[1877] = layer0_outputs[667];
    assign layer1_outputs[1878] = 1'b1;
    assign layer1_outputs[1879] = ~(layer0_outputs[371]) | (layer0_outputs[228]);
    assign layer1_outputs[1880] = ~(layer0_outputs[1156]) | (layer0_outputs[2233]);
    assign layer1_outputs[1881] = (layer0_outputs[680]) & ~(layer0_outputs[999]);
    assign layer1_outputs[1882] = layer0_outputs[1055];
    assign layer1_outputs[1883] = (layer0_outputs[2357]) & ~(layer0_outputs[1957]);
    assign layer1_outputs[1884] = ~((layer0_outputs[1165]) | (layer0_outputs[436]));
    assign layer1_outputs[1885] = (layer0_outputs[999]) & ~(layer0_outputs[140]);
    assign layer1_outputs[1886] = ~(layer0_outputs[1691]);
    assign layer1_outputs[1887] = ~((layer0_outputs[2444]) ^ (layer0_outputs[1617]));
    assign layer1_outputs[1888] = ~((layer0_outputs[374]) | (layer0_outputs[2278]));
    assign layer1_outputs[1889] = (layer0_outputs[1053]) & (layer0_outputs[459]);
    assign layer1_outputs[1890] = ~(layer0_outputs[271]);
    assign layer1_outputs[1891] = ~(layer0_outputs[751]) | (layer0_outputs[329]);
    assign layer1_outputs[1892] = 1'b1;
    assign layer1_outputs[1893] = (layer0_outputs[1627]) & (layer0_outputs[1645]);
    assign layer1_outputs[1894] = ~((layer0_outputs[419]) | (layer0_outputs[1005]));
    assign layer1_outputs[1895] = layer0_outputs[1823];
    assign layer1_outputs[1896] = (layer0_outputs[2099]) & (layer0_outputs[2271]);
    assign layer1_outputs[1897] = (layer0_outputs[2131]) & (layer0_outputs[478]);
    assign layer1_outputs[1898] = 1'b0;
    assign layer1_outputs[1899] = (layer0_outputs[24]) & (layer0_outputs[1579]);
    assign layer1_outputs[1900] = ~((layer0_outputs[1332]) & (layer0_outputs[332]));
    assign layer1_outputs[1901] = ~((layer0_outputs[2130]) | (layer0_outputs[87]));
    assign layer1_outputs[1902] = layer0_outputs[1495];
    assign layer1_outputs[1903] = (layer0_outputs[865]) & (layer0_outputs[100]);
    assign layer1_outputs[1904] = (layer0_outputs[374]) & (layer0_outputs[1578]);
    assign layer1_outputs[1905] = ~(layer0_outputs[300]);
    assign layer1_outputs[1906] = layer0_outputs[2029];
    assign layer1_outputs[1907] = 1'b1;
    assign layer1_outputs[1908] = (layer0_outputs[171]) & (layer0_outputs[467]);
    assign layer1_outputs[1909] = ~(layer0_outputs[2071]) | (layer0_outputs[990]);
    assign layer1_outputs[1910] = 1'b0;
    assign layer1_outputs[1911] = (layer0_outputs[802]) & ~(layer0_outputs[2462]);
    assign layer1_outputs[1912] = (layer0_outputs[698]) & (layer0_outputs[123]);
    assign layer1_outputs[1913] = ~((layer0_outputs[601]) ^ (layer0_outputs[1048]));
    assign layer1_outputs[1914] = (layer0_outputs[194]) & ~(layer0_outputs[2105]);
    assign layer1_outputs[1915] = (layer0_outputs[1562]) & (layer0_outputs[2036]);
    assign layer1_outputs[1916] = (layer0_outputs[222]) & (layer0_outputs[1204]);
    assign layer1_outputs[1917] = (layer0_outputs[949]) | (layer0_outputs[1269]);
    assign layer1_outputs[1918] = ~(layer0_outputs[2140]) | (layer0_outputs[219]);
    assign layer1_outputs[1919] = (layer0_outputs[687]) & ~(layer0_outputs[2081]);
    assign layer1_outputs[1920] = ~(layer0_outputs[1627]) | (layer0_outputs[1584]);
    assign layer1_outputs[1921] = ~(layer0_outputs[1905]);
    assign layer1_outputs[1922] = (layer0_outputs[1571]) & (layer0_outputs[923]);
    assign layer1_outputs[1923] = layer0_outputs[782];
    assign layer1_outputs[1924] = (layer0_outputs[444]) & ~(layer0_outputs[635]);
    assign layer1_outputs[1925] = 1'b0;
    assign layer1_outputs[1926] = 1'b1;
    assign layer1_outputs[1927] = (layer0_outputs[703]) & (layer0_outputs[2152]);
    assign layer1_outputs[1928] = layer0_outputs[2258];
    assign layer1_outputs[1929] = layer0_outputs[604];
    assign layer1_outputs[1930] = layer0_outputs[1609];
    assign layer1_outputs[1931] = (layer0_outputs[2309]) | (layer0_outputs[2344]);
    assign layer1_outputs[1932] = ~((layer0_outputs[440]) & (layer0_outputs[1279]));
    assign layer1_outputs[1933] = (layer0_outputs[690]) & ~(layer0_outputs[950]);
    assign layer1_outputs[1934] = (layer0_outputs[488]) | (layer0_outputs[2213]);
    assign layer1_outputs[1935] = layer0_outputs[612];
    assign layer1_outputs[1936] = (layer0_outputs[1917]) & (layer0_outputs[1222]);
    assign layer1_outputs[1937] = ~((layer0_outputs[1193]) | (layer0_outputs[793]));
    assign layer1_outputs[1938] = ~((layer0_outputs[2377]) & (layer0_outputs[1199]));
    assign layer1_outputs[1939] = (layer0_outputs[893]) & (layer0_outputs[1680]);
    assign layer1_outputs[1940] = (layer0_outputs[848]) & ~(layer0_outputs[2014]);
    assign layer1_outputs[1941] = (layer0_outputs[1838]) & ~(layer0_outputs[946]);
    assign layer1_outputs[1942] = ~((layer0_outputs[1187]) | (layer0_outputs[795]));
    assign layer1_outputs[1943] = ~(layer0_outputs[1834]);
    assign layer1_outputs[1944] = ~((layer0_outputs[1685]) | (layer0_outputs[1032]));
    assign layer1_outputs[1945] = ~((layer0_outputs[709]) ^ (layer0_outputs[2305]));
    assign layer1_outputs[1946] = layer0_outputs[1063];
    assign layer1_outputs[1947] = layer0_outputs[1339];
    assign layer1_outputs[1948] = (layer0_outputs[2119]) | (layer0_outputs[1570]);
    assign layer1_outputs[1949] = layer0_outputs[1569];
    assign layer1_outputs[1950] = (layer0_outputs[2423]) & (layer0_outputs[1989]);
    assign layer1_outputs[1951] = ~(layer0_outputs[797]);
    assign layer1_outputs[1952] = ~(layer0_outputs[2231]);
    assign layer1_outputs[1953] = ~(layer0_outputs[448]);
    assign layer1_outputs[1954] = ~((layer0_outputs[1707]) ^ (layer0_outputs[534]));
    assign layer1_outputs[1955] = ~((layer0_outputs[566]) & (layer0_outputs[1639]));
    assign layer1_outputs[1956] = 1'b0;
    assign layer1_outputs[1957] = (layer0_outputs[273]) & (layer0_outputs[879]);
    assign layer1_outputs[1958] = (layer0_outputs[2143]) & ~(layer0_outputs[2025]);
    assign layer1_outputs[1959] = ~(layer0_outputs[855]) | (layer0_outputs[2488]);
    assign layer1_outputs[1960] = ~(layer0_outputs[524]) | (layer0_outputs[260]);
    assign layer1_outputs[1961] = (layer0_outputs[1933]) & ~(layer0_outputs[2019]);
    assign layer1_outputs[1962] = layer0_outputs[1526];
    assign layer1_outputs[1963] = ~(layer0_outputs[868]);
    assign layer1_outputs[1964] = ~((layer0_outputs[1436]) | (layer0_outputs[1258]));
    assign layer1_outputs[1965] = layer0_outputs[1226];
    assign layer1_outputs[1966] = layer0_outputs[2235];
    assign layer1_outputs[1967] = ~(layer0_outputs[914]);
    assign layer1_outputs[1968] = layer0_outputs[238];
    assign layer1_outputs[1969] = ~((layer0_outputs[982]) & (layer0_outputs[2495]));
    assign layer1_outputs[1970] = ~(layer0_outputs[69]);
    assign layer1_outputs[1971] = layer0_outputs[1912];
    assign layer1_outputs[1972] = (layer0_outputs[2384]) | (layer0_outputs[2095]);
    assign layer1_outputs[1973] = (layer0_outputs[2371]) ^ (layer0_outputs[1550]);
    assign layer1_outputs[1974] = ~(layer0_outputs[186]);
    assign layer1_outputs[1975] = 1'b0;
    assign layer1_outputs[1976] = (layer0_outputs[2237]) & (layer0_outputs[804]);
    assign layer1_outputs[1977] = (layer0_outputs[317]) ^ (layer0_outputs[1366]);
    assign layer1_outputs[1978] = (layer0_outputs[924]) & (layer0_outputs[53]);
    assign layer1_outputs[1979] = (layer0_outputs[1442]) | (layer0_outputs[663]);
    assign layer1_outputs[1980] = layer0_outputs[1734];
    assign layer1_outputs[1981] = layer0_outputs[472];
    assign layer1_outputs[1982] = ~(layer0_outputs[873]) | (layer0_outputs[1523]);
    assign layer1_outputs[1983] = (layer0_outputs[1371]) | (layer0_outputs[347]);
    assign layer1_outputs[1984] = ~((layer0_outputs[220]) & (layer0_outputs[14]));
    assign layer1_outputs[1985] = ~((layer0_outputs[1811]) ^ (layer0_outputs[1502]));
    assign layer1_outputs[1986] = ~(layer0_outputs[2125]) | (layer0_outputs[166]);
    assign layer1_outputs[1987] = layer0_outputs[585];
    assign layer1_outputs[1988] = ~((layer0_outputs[297]) & (layer0_outputs[2239]));
    assign layer1_outputs[1989] = (layer0_outputs[996]) & ~(layer0_outputs[1147]);
    assign layer1_outputs[1990] = (layer0_outputs[770]) & (layer0_outputs[1210]);
    assign layer1_outputs[1991] = ~(layer0_outputs[1979]);
    assign layer1_outputs[1992] = ~(layer0_outputs[465]);
    assign layer1_outputs[1993] = layer0_outputs[982];
    assign layer1_outputs[1994] = ~(layer0_outputs[2108]) | (layer0_outputs[1990]);
    assign layer1_outputs[1995] = ~((layer0_outputs[1635]) & (layer0_outputs[2532]));
    assign layer1_outputs[1996] = (layer0_outputs[315]) | (layer0_outputs[2345]);
    assign layer1_outputs[1997] = 1'b1;
    assign layer1_outputs[1998] = layer0_outputs[1395];
    assign layer1_outputs[1999] = ~((layer0_outputs[688]) & (layer0_outputs[127]));
    assign layer1_outputs[2000] = (layer0_outputs[2005]) & ~(layer0_outputs[1824]);
    assign layer1_outputs[2001] = ~(layer0_outputs[748]);
    assign layer1_outputs[2002] = layer0_outputs[2176];
    assign layer1_outputs[2003] = (layer0_outputs[774]) & ~(layer0_outputs[2157]);
    assign layer1_outputs[2004] = (layer0_outputs[45]) & (layer0_outputs[1993]);
    assign layer1_outputs[2005] = (layer0_outputs[512]) & (layer0_outputs[2546]);
    assign layer1_outputs[2006] = 1'b0;
    assign layer1_outputs[2007] = ~((layer0_outputs[1611]) ^ (layer0_outputs[1036]));
    assign layer1_outputs[2008] = ~(layer0_outputs[2310]) | (layer0_outputs[2082]);
    assign layer1_outputs[2009] = ~((layer0_outputs[29]) & (layer0_outputs[671]));
    assign layer1_outputs[2010] = ~(layer0_outputs[850]);
    assign layer1_outputs[2011] = ~(layer0_outputs[296]) | (layer0_outputs[1720]);
    assign layer1_outputs[2012] = 1'b0;
    assign layer1_outputs[2013] = (layer0_outputs[1547]) & (layer0_outputs[2382]);
    assign layer1_outputs[2014] = ~(layer0_outputs[1974]) | (layer0_outputs[1241]);
    assign layer1_outputs[2015] = ~((layer0_outputs[1478]) & (layer0_outputs[76]));
    assign layer1_outputs[2016] = (layer0_outputs[1385]) & ~(layer0_outputs[428]);
    assign layer1_outputs[2017] = ~(layer0_outputs[1981]) | (layer0_outputs[2312]);
    assign layer1_outputs[2018] = 1'b1;
    assign layer1_outputs[2019] = ~(layer0_outputs[2501]);
    assign layer1_outputs[2020] = 1'b0;
    assign layer1_outputs[2021] = ~((layer0_outputs[2422]) | (layer0_outputs[1242]));
    assign layer1_outputs[2022] = ~((layer0_outputs[1084]) & (layer0_outputs[1004]));
    assign layer1_outputs[2023] = ~(layer0_outputs[1877]) | (layer0_outputs[176]);
    assign layer1_outputs[2024] = (layer0_outputs[2070]) | (layer0_outputs[1121]);
    assign layer1_outputs[2025] = ~(layer0_outputs[175]) | (layer0_outputs[102]);
    assign layer1_outputs[2026] = ~((layer0_outputs[1206]) & (layer0_outputs[1835]));
    assign layer1_outputs[2027] = 1'b1;
    assign layer1_outputs[2028] = ~(layer0_outputs[487]) | (layer0_outputs[2526]);
    assign layer1_outputs[2029] = ~((layer0_outputs[1799]) & (layer0_outputs[1815]));
    assign layer1_outputs[2030] = ~((layer0_outputs[2215]) ^ (layer0_outputs[887]));
    assign layer1_outputs[2031] = (layer0_outputs[1501]) & ~(layer0_outputs[441]);
    assign layer1_outputs[2032] = ~((layer0_outputs[1037]) & (layer0_outputs[118]));
    assign layer1_outputs[2033] = ~((layer0_outputs[353]) ^ (layer0_outputs[1095]));
    assign layer1_outputs[2034] = ~(layer0_outputs[2396]);
    assign layer1_outputs[2035] = 1'b0;
    assign layer1_outputs[2036] = layer0_outputs[434];
    assign layer1_outputs[2037] = layer0_outputs[1890];
    assign layer1_outputs[2038] = 1'b1;
    assign layer1_outputs[2039] = (layer0_outputs[218]) | (layer0_outputs[2125]);
    assign layer1_outputs[2040] = (layer0_outputs[1215]) & ~(layer0_outputs[1045]);
    assign layer1_outputs[2041] = ~((layer0_outputs[224]) | (layer0_outputs[1283]));
    assign layer1_outputs[2042] = ~(layer0_outputs[1928]);
    assign layer1_outputs[2043] = 1'b0;
    assign layer1_outputs[2044] = (layer0_outputs[907]) ^ (layer0_outputs[2002]);
    assign layer1_outputs[2045] = ~((layer0_outputs[92]) | (layer0_outputs[1415]));
    assign layer1_outputs[2046] = 1'b1;
    assign layer1_outputs[2047] = layer0_outputs[2302];
    assign layer1_outputs[2048] = ~(layer0_outputs[1961]) | (layer0_outputs[2024]);
    assign layer1_outputs[2049] = layer0_outputs[382];
    assign layer1_outputs[2050] = layer0_outputs[719];
    assign layer1_outputs[2051] = ~(layer0_outputs[723]);
    assign layer1_outputs[2052] = (layer0_outputs[953]) | (layer0_outputs[1639]);
    assign layer1_outputs[2053] = layer0_outputs[2429];
    assign layer1_outputs[2054] = (layer0_outputs[78]) & (layer0_outputs[1139]);
    assign layer1_outputs[2055] = (layer0_outputs[1009]) | (layer0_outputs[1718]);
    assign layer1_outputs[2056] = 1'b0;
    assign layer1_outputs[2057] = (layer0_outputs[2098]) & ~(layer0_outputs[435]);
    assign layer1_outputs[2058] = ~(layer0_outputs[155]) | (layer0_outputs[1267]);
    assign layer1_outputs[2059] = ~(layer0_outputs[891]) | (layer0_outputs[1880]);
    assign layer1_outputs[2060] = ~(layer0_outputs[610]);
    assign layer1_outputs[2061] = (layer0_outputs[1673]) | (layer0_outputs[2513]);
    assign layer1_outputs[2062] = (layer0_outputs[1492]) & ~(layer0_outputs[2467]);
    assign layer1_outputs[2063] = (layer0_outputs[174]) & (layer0_outputs[2046]);
    assign layer1_outputs[2064] = ~(layer0_outputs[2458]) | (layer0_outputs[880]);
    assign layer1_outputs[2065] = (layer0_outputs[1757]) & ~(layer0_outputs[2274]);
    assign layer1_outputs[2066] = (layer0_outputs[576]) & ~(layer0_outputs[939]);
    assign layer1_outputs[2067] = 1'b0;
    assign layer1_outputs[2068] = ~(layer0_outputs[2302]);
    assign layer1_outputs[2069] = layer0_outputs[2320];
    assign layer1_outputs[2070] = (layer0_outputs[1087]) & (layer0_outputs[901]);
    assign layer1_outputs[2071] = ~((layer0_outputs[782]) ^ (layer0_outputs[1925]));
    assign layer1_outputs[2072] = ~(layer0_outputs[2326]);
    assign layer1_outputs[2073] = (layer0_outputs[678]) & ~(layer0_outputs[2431]);
    assign layer1_outputs[2074] = layer0_outputs[675];
    assign layer1_outputs[2075] = (layer0_outputs[1431]) ^ (layer0_outputs[2086]);
    assign layer1_outputs[2076] = ~(layer0_outputs[746]) | (layer0_outputs[30]);
    assign layer1_outputs[2077] = 1'b1;
    assign layer1_outputs[2078] = ~(layer0_outputs[1975]) | (layer0_outputs[1112]);
    assign layer1_outputs[2079] = (layer0_outputs[901]) | (layer0_outputs[29]);
    assign layer1_outputs[2080] = ~(layer0_outputs[477]);
    assign layer1_outputs[2081] = layer0_outputs[980];
    assign layer1_outputs[2082] = (layer0_outputs[1093]) & ~(layer0_outputs[1094]);
    assign layer1_outputs[2083] = ~(layer0_outputs[2323]) | (layer0_outputs[2223]);
    assign layer1_outputs[2084] = 1'b1;
    assign layer1_outputs[2085] = ~(layer0_outputs[1409]);
    assign layer1_outputs[2086] = (layer0_outputs[1263]) | (layer0_outputs[1963]);
    assign layer1_outputs[2087] = (layer0_outputs[218]) & ~(layer0_outputs[2453]);
    assign layer1_outputs[2088] = layer0_outputs[1557];
    assign layer1_outputs[2089] = ~((layer0_outputs[720]) ^ (layer0_outputs[938]));
    assign layer1_outputs[2090] = 1'b1;
    assign layer1_outputs[2091] = ~(layer0_outputs[1921]) | (layer0_outputs[284]);
    assign layer1_outputs[2092] = (layer0_outputs[1480]) ^ (layer0_outputs[951]);
    assign layer1_outputs[2093] = ~(layer0_outputs[2443]);
    assign layer1_outputs[2094] = ~((layer0_outputs[204]) & (layer0_outputs[2384]));
    assign layer1_outputs[2095] = (layer0_outputs[332]) & ~(layer0_outputs[330]);
    assign layer1_outputs[2096] = layer0_outputs[2314];
    assign layer1_outputs[2097] = (layer0_outputs[356]) & ~(layer0_outputs[1785]);
    assign layer1_outputs[2098] = ~(layer0_outputs[691]);
    assign layer1_outputs[2099] = layer0_outputs[114];
    assign layer1_outputs[2100] = (layer0_outputs[1533]) & ~(layer0_outputs[1872]);
    assign layer1_outputs[2101] = (layer0_outputs[1329]) ^ (layer0_outputs[375]);
    assign layer1_outputs[2102] = layer0_outputs[1576];
    assign layer1_outputs[2103] = ~(layer0_outputs[1025]);
    assign layer1_outputs[2104] = (layer0_outputs[358]) & ~(layer0_outputs[2381]);
    assign layer1_outputs[2105] = (layer0_outputs[199]) ^ (layer0_outputs[186]);
    assign layer1_outputs[2106] = ~((layer0_outputs[638]) | (layer0_outputs[1598]));
    assign layer1_outputs[2107] = (layer0_outputs[847]) & ~(layer0_outputs[2508]);
    assign layer1_outputs[2108] = ~(layer0_outputs[599]) | (layer0_outputs[377]);
    assign layer1_outputs[2109] = layer0_outputs[203];
    assign layer1_outputs[2110] = ~(layer0_outputs[2073]) | (layer0_outputs[2124]);
    assign layer1_outputs[2111] = ~((layer0_outputs[1008]) | (layer0_outputs[150]));
    assign layer1_outputs[2112] = (layer0_outputs[1385]) | (layer0_outputs[411]);
    assign layer1_outputs[2113] = 1'b0;
    assign layer1_outputs[2114] = ~((layer0_outputs[322]) & (layer0_outputs[324]));
    assign layer1_outputs[2115] = layer0_outputs[489];
    assign layer1_outputs[2116] = ~((layer0_outputs[657]) ^ (layer0_outputs[2059]));
    assign layer1_outputs[2117] = (layer0_outputs[1881]) & ~(layer0_outputs[1396]);
    assign layer1_outputs[2118] = (layer0_outputs[2175]) | (layer0_outputs[1215]);
    assign layer1_outputs[2119] = ~(layer0_outputs[1108]);
    assign layer1_outputs[2120] = layer0_outputs[1873];
    assign layer1_outputs[2121] = ~((layer0_outputs[2092]) | (layer0_outputs[2115]));
    assign layer1_outputs[2122] = layer0_outputs[2068];
    assign layer1_outputs[2123] = layer0_outputs[791];
    assign layer1_outputs[2124] = (layer0_outputs[2412]) & (layer0_outputs[2454]);
    assign layer1_outputs[2125] = 1'b1;
    assign layer1_outputs[2126] = 1'b1;
    assign layer1_outputs[2127] = 1'b1;
    assign layer1_outputs[2128] = ~(layer0_outputs[112]);
    assign layer1_outputs[2129] = layer0_outputs[2188];
    assign layer1_outputs[2130] = layer0_outputs[677];
    assign layer1_outputs[2131] = ~((layer0_outputs[1111]) | (layer0_outputs[340]));
    assign layer1_outputs[2132] = ~((layer0_outputs[878]) | (layer0_outputs[1251]));
    assign layer1_outputs[2133] = (layer0_outputs[2249]) & ~(layer0_outputs[655]);
    assign layer1_outputs[2134] = (layer0_outputs[406]) | (layer0_outputs[774]);
    assign layer1_outputs[2135] = ~(layer0_outputs[1000]);
    assign layer1_outputs[2136] = 1'b0;
    assign layer1_outputs[2137] = (layer0_outputs[2335]) & ~(layer0_outputs[209]);
    assign layer1_outputs[2138] = ~((layer0_outputs[217]) & (layer0_outputs[2116]));
    assign layer1_outputs[2139] = (layer0_outputs[2402]) & (layer0_outputs[1885]);
    assign layer1_outputs[2140] = ~((layer0_outputs[2545]) ^ (layer0_outputs[890]));
    assign layer1_outputs[2141] = layer0_outputs[851];
    assign layer1_outputs[2142] = ~(layer0_outputs[940]);
    assign layer1_outputs[2143] = ~(layer0_outputs[2402]) | (layer0_outputs[2486]);
    assign layer1_outputs[2144] = ~(layer0_outputs[1084]);
    assign layer1_outputs[2145] = (layer0_outputs[685]) | (layer0_outputs[2465]);
    assign layer1_outputs[2146] = ~(layer0_outputs[1161]) | (layer0_outputs[2022]);
    assign layer1_outputs[2147] = ~((layer0_outputs[1814]) & (layer0_outputs[2447]));
    assign layer1_outputs[2148] = ~((layer0_outputs[1589]) & (layer0_outputs[2404]));
    assign layer1_outputs[2149] = 1'b1;
    assign layer1_outputs[2150] = ~(layer0_outputs[1675]);
    assign layer1_outputs[2151] = (layer0_outputs[1845]) & (layer0_outputs[1870]);
    assign layer1_outputs[2152] = layer0_outputs[131];
    assign layer1_outputs[2153] = ~(layer0_outputs[992]) | (layer0_outputs[1178]);
    assign layer1_outputs[2154] = ~(layer0_outputs[788]);
    assign layer1_outputs[2155] = ~(layer0_outputs[673]);
    assign layer1_outputs[2156] = (layer0_outputs[74]) | (layer0_outputs[1904]);
    assign layer1_outputs[2157] = 1'b0;
    assign layer1_outputs[2158] = 1'b1;
    assign layer1_outputs[2159] = ~(layer0_outputs[1622]) | (layer0_outputs[177]);
    assign layer1_outputs[2160] = ~((layer0_outputs[1382]) | (layer0_outputs[1194]));
    assign layer1_outputs[2161] = ~((layer0_outputs[1019]) & (layer0_outputs[918]));
    assign layer1_outputs[2162] = 1'b1;
    assign layer1_outputs[2163] = 1'b1;
    assign layer1_outputs[2164] = ~(layer0_outputs[267]) | (layer0_outputs[544]);
    assign layer1_outputs[2165] = layer0_outputs[473];
    assign layer1_outputs[2166] = ~(layer0_outputs[1424]);
    assign layer1_outputs[2167] = 1'b0;
    assign layer1_outputs[2168] = layer0_outputs[211];
    assign layer1_outputs[2169] = ~(layer0_outputs[1497]);
    assign layer1_outputs[2170] = ~((layer0_outputs[2450]) ^ (layer0_outputs[1731]));
    assign layer1_outputs[2171] = ~(layer0_outputs[1576]) | (layer0_outputs[1399]);
    assign layer1_outputs[2172] = layer0_outputs[246];
    assign layer1_outputs[2173] = (layer0_outputs[1499]) & ~(layer0_outputs[1777]);
    assign layer1_outputs[2174] = ~(layer0_outputs[2450]);
    assign layer1_outputs[2175] = ~(layer0_outputs[2240]);
    assign layer1_outputs[2176] = ~(layer0_outputs[32]);
    assign layer1_outputs[2177] = ~((layer0_outputs[1650]) & (layer0_outputs[2217]));
    assign layer1_outputs[2178] = ~(layer0_outputs[2225]);
    assign layer1_outputs[2179] = (layer0_outputs[66]) & ~(layer0_outputs[1241]);
    assign layer1_outputs[2180] = (layer0_outputs[407]) | (layer0_outputs[2123]);
    assign layer1_outputs[2181] = ~((layer0_outputs[1348]) ^ (layer0_outputs[1068]));
    assign layer1_outputs[2182] = 1'b0;
    assign layer1_outputs[2183] = ~((layer0_outputs[214]) | (layer0_outputs[157]));
    assign layer1_outputs[2184] = layer0_outputs[1987];
    assign layer1_outputs[2185] = (layer0_outputs[1453]) & ~(layer0_outputs[700]);
    assign layer1_outputs[2186] = ~((layer0_outputs[993]) | (layer0_outputs[1489]));
    assign layer1_outputs[2187] = (layer0_outputs[2477]) & (layer0_outputs[144]);
    assign layer1_outputs[2188] = ~(layer0_outputs[1861]) | (layer0_outputs[2078]);
    assign layer1_outputs[2189] = 1'b1;
    assign layer1_outputs[2190] = layer0_outputs[1692];
    assign layer1_outputs[2191] = (layer0_outputs[1580]) & (layer0_outputs[1716]);
    assign layer1_outputs[2192] = ~(layer0_outputs[2]);
    assign layer1_outputs[2193] = ~(layer0_outputs[2083]);
    assign layer1_outputs[2194] = ~(layer0_outputs[165]);
    assign layer1_outputs[2195] = (layer0_outputs[1583]) ^ (layer0_outputs[2277]);
    assign layer1_outputs[2196] = (layer0_outputs[234]) | (layer0_outputs[824]);
    assign layer1_outputs[2197] = ~(layer0_outputs[2068]);
    assign layer1_outputs[2198] = (layer0_outputs[1251]) | (layer0_outputs[1911]);
    assign layer1_outputs[2199] = 1'b0;
    assign layer1_outputs[2200] = 1'b0;
    assign layer1_outputs[2201] = (layer0_outputs[1070]) & ~(layer0_outputs[412]);
    assign layer1_outputs[2202] = (layer0_outputs[2122]) & ~(layer0_outputs[1822]);
    assign layer1_outputs[2203] = ~((layer0_outputs[686]) & (layer0_outputs[661]));
    assign layer1_outputs[2204] = layer0_outputs[343];
    assign layer1_outputs[2205] = ~((layer0_outputs[1504]) | (layer0_outputs[139]));
    assign layer1_outputs[2206] = ~((layer0_outputs[1703]) & (layer0_outputs[343]));
    assign layer1_outputs[2207] = 1'b1;
    assign layer1_outputs[2208] = (layer0_outputs[1377]) & ~(layer0_outputs[326]);
    assign layer1_outputs[2209] = (layer0_outputs[2196]) & (layer0_outputs[1452]);
    assign layer1_outputs[2210] = (layer0_outputs[1944]) & ~(layer0_outputs[335]);
    assign layer1_outputs[2211] = 1'b0;
    assign layer1_outputs[2212] = ~(layer0_outputs[942]);
    assign layer1_outputs[2213] = ~(layer0_outputs[1101]) | (layer0_outputs[2272]);
    assign layer1_outputs[2214] = ~(layer0_outputs[490]);
    assign layer1_outputs[2215] = ~((layer0_outputs[2055]) | (layer0_outputs[190]));
    assign layer1_outputs[2216] = (layer0_outputs[2038]) & ~(layer0_outputs[903]);
    assign layer1_outputs[2217] = (layer0_outputs[241]) & ~(layer0_outputs[679]);
    assign layer1_outputs[2218] = 1'b1;
    assign layer1_outputs[2219] = layer0_outputs[44];
    assign layer1_outputs[2220] = ~(layer0_outputs[191]) | (layer0_outputs[2169]);
    assign layer1_outputs[2221] = ~(layer0_outputs[4]);
    assign layer1_outputs[2222] = ~(layer0_outputs[1826]);
    assign layer1_outputs[2223] = (layer0_outputs[1025]) | (layer0_outputs[1154]);
    assign layer1_outputs[2224] = ~(layer0_outputs[1721]) | (layer0_outputs[1341]);
    assign layer1_outputs[2225] = layer0_outputs[215];
    assign layer1_outputs[2226] = ~(layer0_outputs[443]) | (layer0_outputs[260]);
    assign layer1_outputs[2227] = layer0_outputs[1730];
    assign layer1_outputs[2228] = ~((layer0_outputs[2005]) | (layer0_outputs[619]));
    assign layer1_outputs[2229] = (layer0_outputs[368]) & ~(layer0_outputs[2520]);
    assign layer1_outputs[2230] = layer0_outputs[2416];
    assign layer1_outputs[2231] = ~(layer0_outputs[685]);
    assign layer1_outputs[2232] = ~(layer0_outputs[2232]);
    assign layer1_outputs[2233] = ~((layer0_outputs[2528]) | (layer0_outputs[227]));
    assign layer1_outputs[2234] = (layer0_outputs[904]) & (layer0_outputs[2063]);
    assign layer1_outputs[2235] = ~(layer0_outputs[164]);
    assign layer1_outputs[2236] = ~(layer0_outputs[573]) | (layer0_outputs[315]);
    assign layer1_outputs[2237] = (layer0_outputs[184]) & ~(layer0_outputs[1693]);
    assign layer1_outputs[2238] = 1'b0;
    assign layer1_outputs[2239] = ~(layer0_outputs[79]);
    assign layer1_outputs[2240] = (layer0_outputs[1863]) | (layer0_outputs[1010]);
    assign layer1_outputs[2241] = layer0_outputs[2286];
    assign layer1_outputs[2242] = ~(layer0_outputs[2559]);
    assign layer1_outputs[2243] = ~(layer0_outputs[2375]);
    assign layer1_outputs[2244] = 1'b0;
    assign layer1_outputs[2245] = 1'b1;
    assign layer1_outputs[2246] = 1'b1;
    assign layer1_outputs[2247] = layer0_outputs[277];
    assign layer1_outputs[2248] = ~(layer0_outputs[2032]);
    assign layer1_outputs[2249] = ~(layer0_outputs[2115]) | (layer0_outputs[1831]);
    assign layer1_outputs[2250] = ~((layer0_outputs[2194]) | (layer0_outputs[1869]));
    assign layer1_outputs[2251] = ~((layer0_outputs[381]) | (layer0_outputs[1301]));
    assign layer1_outputs[2252] = ~(layer0_outputs[196]);
    assign layer1_outputs[2253] = ~(layer0_outputs[131]);
    assign layer1_outputs[2254] = (layer0_outputs[1185]) & ~(layer0_outputs[251]);
    assign layer1_outputs[2255] = ~((layer0_outputs[890]) | (layer0_outputs[361]));
    assign layer1_outputs[2256] = ~(layer0_outputs[1490]);
    assign layer1_outputs[2257] = ~(layer0_outputs[64]) | (layer0_outputs[266]);
    assign layer1_outputs[2258] = layer0_outputs[1367];
    assign layer1_outputs[2259] = layer0_outputs[2064];
    assign layer1_outputs[2260] = layer0_outputs[1244];
    assign layer1_outputs[2261] = 1'b0;
    assign layer1_outputs[2262] = ~(layer0_outputs[1227]) | (layer0_outputs[2203]);
    assign layer1_outputs[2263] = (layer0_outputs[134]) | (layer0_outputs[1130]);
    assign layer1_outputs[2264] = ~((layer0_outputs[338]) | (layer0_outputs[11]));
    assign layer1_outputs[2265] = ~(layer0_outputs[2406]);
    assign layer1_outputs[2266] = (layer0_outputs[1706]) & ~(layer0_outputs[1187]);
    assign layer1_outputs[2267] = ~(layer0_outputs[2128]) | (layer0_outputs[1518]);
    assign layer1_outputs[2268] = (layer0_outputs[921]) & ~(layer0_outputs[1508]);
    assign layer1_outputs[2269] = ~(layer0_outputs[1054]);
    assign layer1_outputs[2270] = layer0_outputs[1543];
    assign layer1_outputs[2271] = (layer0_outputs[511]) ^ (layer0_outputs[282]);
    assign layer1_outputs[2272] = (layer0_outputs[1544]) & ~(layer0_outputs[786]);
    assign layer1_outputs[2273] = ~((layer0_outputs[2356]) & (layer0_outputs[1209]));
    assign layer1_outputs[2274] = ~(layer0_outputs[2030]);
    assign layer1_outputs[2275] = ~(layer0_outputs[671]);
    assign layer1_outputs[2276] = (layer0_outputs[2497]) & (layer0_outputs[2241]);
    assign layer1_outputs[2277] = ~(layer0_outputs[1532]);
    assign layer1_outputs[2278] = ~(layer0_outputs[2149]);
    assign layer1_outputs[2279] = (layer0_outputs[432]) & (layer0_outputs[1678]);
    assign layer1_outputs[2280] = ~((layer0_outputs[1472]) & (layer0_outputs[471]));
    assign layer1_outputs[2281] = ~(layer0_outputs[1629]) | (layer0_outputs[818]);
    assign layer1_outputs[2282] = 1'b0;
    assign layer1_outputs[2283] = layer0_outputs[718];
    assign layer1_outputs[2284] = (layer0_outputs[2322]) & ~(layer0_outputs[2554]);
    assign layer1_outputs[2285] = (layer0_outputs[929]) | (layer0_outputs[2404]);
    assign layer1_outputs[2286] = 1'b0;
    assign layer1_outputs[2287] = ~(layer0_outputs[2527]);
    assign layer1_outputs[2288] = ~(layer0_outputs[1184]) | (layer0_outputs[535]);
    assign layer1_outputs[2289] = (layer0_outputs[822]) & ~(layer0_outputs[2282]);
    assign layer1_outputs[2290] = (layer0_outputs[892]) & (layer0_outputs[832]);
    assign layer1_outputs[2291] = (layer0_outputs[1774]) & ~(layer0_outputs[1530]);
    assign layer1_outputs[2292] = ~(layer0_outputs[526]) | (layer0_outputs[951]);
    assign layer1_outputs[2293] = 1'b1;
    assign layer1_outputs[2294] = ~(layer0_outputs[1581]);
    assign layer1_outputs[2295] = ~((layer0_outputs[1344]) & (layer0_outputs[1895]));
    assign layer1_outputs[2296] = ~(layer0_outputs[1436]);
    assign layer1_outputs[2297] = 1'b1;
    assign layer1_outputs[2298] = ~(layer0_outputs[160]);
    assign layer1_outputs[2299] = ~((layer0_outputs[676]) & (layer0_outputs[2062]));
    assign layer1_outputs[2300] = ~((layer0_outputs[2168]) & (layer0_outputs[1223]));
    assign layer1_outputs[2301] = ~(layer0_outputs[2180]);
    assign layer1_outputs[2302] = (layer0_outputs[2515]) | (layer0_outputs[1519]);
    assign layer1_outputs[2303] = layer0_outputs[716];
    assign layer1_outputs[2304] = ~(layer0_outputs[2219]) | (layer0_outputs[727]);
    assign layer1_outputs[2305] = ~((layer0_outputs[1322]) | (layer0_outputs[2341]));
    assign layer1_outputs[2306] = (layer0_outputs[2442]) & (layer0_outputs[1265]);
    assign layer1_outputs[2307] = ~(layer0_outputs[935]);
    assign layer1_outputs[2308] = ~(layer0_outputs[1835]) | (layer0_outputs[405]);
    assign layer1_outputs[2309] = ~((layer0_outputs[2185]) ^ (layer0_outputs[1842]));
    assign layer1_outputs[2310] = ~(layer0_outputs[1360]);
    assign layer1_outputs[2311] = ~(layer0_outputs[462]);
    assign layer1_outputs[2312] = ~((layer0_outputs[1446]) & (layer0_outputs[1866]));
    assign layer1_outputs[2313] = ~((layer0_outputs[615]) & (layer0_outputs[2289]));
    assign layer1_outputs[2314] = ~(layer0_outputs[1486]) | (layer0_outputs[2451]);
    assign layer1_outputs[2315] = layer0_outputs[330];
    assign layer1_outputs[2316] = (layer0_outputs[2436]) | (layer0_outputs[1864]);
    assign layer1_outputs[2317] = ~((layer0_outputs[3]) | (layer0_outputs[1160]));
    assign layer1_outputs[2318] = (layer0_outputs[1432]) | (layer0_outputs[458]);
    assign layer1_outputs[2319] = layer0_outputs[1081];
    assign layer1_outputs[2320] = layer0_outputs[608];
    assign layer1_outputs[2321] = ~(layer0_outputs[65]);
    assign layer1_outputs[2322] = ~((layer0_outputs[1243]) ^ (layer0_outputs[252]));
    assign layer1_outputs[2323] = ~(layer0_outputs[853]);
    assign layer1_outputs[2324] = ~(layer0_outputs[1072]);
    assign layer1_outputs[2325] = layer0_outputs[644];
    assign layer1_outputs[2326] = ~(layer0_outputs[1014]);
    assign layer1_outputs[2327] = (layer0_outputs[1961]) & ~(layer0_outputs[599]);
    assign layer1_outputs[2328] = (layer0_outputs[287]) & (layer0_outputs[81]);
    assign layer1_outputs[2329] = (layer0_outputs[2225]) ^ (layer0_outputs[1221]);
    assign layer1_outputs[2330] = ~(layer0_outputs[22]) | (layer0_outputs[2011]);
    assign layer1_outputs[2331] = layer0_outputs[2347];
    assign layer1_outputs[2332] = ~((layer0_outputs[460]) & (layer0_outputs[1093]));
    assign layer1_outputs[2333] = ~((layer0_outputs[422]) & (layer0_outputs[2427]));
    assign layer1_outputs[2334] = ~(layer0_outputs[722]);
    assign layer1_outputs[2335] = (layer0_outputs[1085]) ^ (layer0_outputs[339]);
    assign layer1_outputs[2336] = ~(layer0_outputs[752]) | (layer0_outputs[2224]);
    assign layer1_outputs[2337] = ~(layer0_outputs[639]);
    assign layer1_outputs[2338] = (layer0_outputs[579]) & ~(layer0_outputs[1892]);
    assign layer1_outputs[2339] = (layer0_outputs[2346]) & ~(layer0_outputs[1891]);
    assign layer1_outputs[2340] = (layer0_outputs[1978]) & ~(layer0_outputs[870]);
    assign layer1_outputs[2341] = ~(layer0_outputs[815]);
    assign layer1_outputs[2342] = (layer0_outputs[2268]) | (layer0_outputs[1772]);
    assign layer1_outputs[2343] = ~(layer0_outputs[2537]);
    assign layer1_outputs[2344] = layer0_outputs[47];
    assign layer1_outputs[2345] = ~(layer0_outputs[1353]);
    assign layer1_outputs[2346] = ~((layer0_outputs[75]) ^ (layer0_outputs[2333]));
    assign layer1_outputs[2347] = ~((layer0_outputs[265]) & (layer0_outputs[682]));
    assign layer1_outputs[2348] = (layer0_outputs[2541]) & (layer0_outputs[1755]);
    assign layer1_outputs[2349] = ~((layer0_outputs[1864]) & (layer0_outputs[39]));
    assign layer1_outputs[2350] = ~(layer0_outputs[2491]) | (layer0_outputs[1643]);
    assign layer1_outputs[2351] = (layer0_outputs[761]) | (layer0_outputs[1040]);
    assign layer1_outputs[2352] = 1'b1;
    assign layer1_outputs[2353] = ~((layer0_outputs[262]) ^ (layer0_outputs[295]));
    assign layer1_outputs[2354] = 1'b1;
    assign layer1_outputs[2355] = layer0_outputs[68];
    assign layer1_outputs[2356] = ~((layer0_outputs[2082]) ^ (layer0_outputs[1463]));
    assign layer1_outputs[2357] = layer0_outputs[2120];
    assign layer1_outputs[2358] = layer0_outputs[1920];
    assign layer1_outputs[2359] = ~((layer0_outputs[1396]) | (layer0_outputs[675]));
    assign layer1_outputs[2360] = ~(layer0_outputs[355]) | (layer0_outputs[537]);
    assign layer1_outputs[2361] = layer0_outputs[1716];
    assign layer1_outputs[2362] = (layer0_outputs[1609]) | (layer0_outputs[2141]);
    assign layer1_outputs[2363] = ~(layer0_outputs[635]) | (layer0_outputs[2266]);
    assign layer1_outputs[2364] = layer0_outputs[271];
    assign layer1_outputs[2365] = (layer0_outputs[867]) | (layer0_outputs[591]);
    assign layer1_outputs[2366] = ~((layer0_outputs[1063]) & (layer0_outputs[51]));
    assign layer1_outputs[2367] = ~((layer0_outputs[1345]) | (layer0_outputs[2275]));
    assign layer1_outputs[2368] = ~(layer0_outputs[861]);
    assign layer1_outputs[2369] = ~(layer0_outputs[536]);
    assign layer1_outputs[2370] = (layer0_outputs[1064]) & (layer0_outputs[2424]);
    assign layer1_outputs[2371] = layer0_outputs[778];
    assign layer1_outputs[2372] = (layer0_outputs[56]) & (layer0_outputs[1951]);
    assign layer1_outputs[2373] = ~((layer0_outputs[941]) & (layer0_outputs[37]));
    assign layer1_outputs[2374] = (layer0_outputs[1770]) & ~(layer0_outputs[2151]);
    assign layer1_outputs[2375] = (layer0_outputs[1924]) ^ (layer0_outputs[710]);
    assign layer1_outputs[2376] = ~((layer0_outputs[294]) & (layer0_outputs[2410]));
    assign layer1_outputs[2377] = ~(layer0_outputs[1308]);
    assign layer1_outputs[2378] = ~((layer0_outputs[1394]) | (layer0_outputs[254]));
    assign layer1_outputs[2379] = ~(layer0_outputs[948]);
    assign layer1_outputs[2380] = (layer0_outputs[1209]) & ~(layer0_outputs[171]);
    assign layer1_outputs[2381] = 1'b0;
    assign layer1_outputs[2382] = ~(layer0_outputs[611]) | (layer0_outputs[1018]);
    assign layer1_outputs[2383] = (layer0_outputs[1642]) | (layer0_outputs[494]);
    assign layer1_outputs[2384] = ~((layer0_outputs[846]) | (layer0_outputs[1797]));
    assign layer1_outputs[2385] = ~(layer0_outputs[1159]) | (layer0_outputs[2000]);
    assign layer1_outputs[2386] = ~((layer0_outputs[1470]) | (layer0_outputs[2436]));
    assign layer1_outputs[2387] = (layer0_outputs[823]) & ~(layer0_outputs[2001]);
    assign layer1_outputs[2388] = (layer0_outputs[141]) & ~(layer0_outputs[620]);
    assign layer1_outputs[2389] = ~(layer0_outputs[713]);
    assign layer1_outputs[2390] = layer0_outputs[2434];
    assign layer1_outputs[2391] = ~((layer0_outputs[193]) & (layer0_outputs[443]));
    assign layer1_outputs[2392] = ~(layer0_outputs[1902]) | (layer0_outputs[318]);
    assign layer1_outputs[2393] = (layer0_outputs[1591]) & (layer0_outputs[757]);
    assign layer1_outputs[2394] = ~(layer0_outputs[1387]);
    assign layer1_outputs[2395] = ~((layer0_outputs[2292]) & (layer0_outputs[290]));
    assign layer1_outputs[2396] = ~((layer0_outputs[2550]) & (layer0_outputs[1516]));
    assign layer1_outputs[2397] = (layer0_outputs[1898]) & (layer0_outputs[163]);
    assign layer1_outputs[2398] = ~((layer0_outputs[1191]) & (layer0_outputs[418]));
    assign layer1_outputs[2399] = (layer0_outputs[541]) | (layer0_outputs[564]);
    assign layer1_outputs[2400] = ~(layer0_outputs[2038]) | (layer0_outputs[1031]);
    assign layer1_outputs[2401] = layer0_outputs[1525];
    assign layer1_outputs[2402] = (layer0_outputs[849]) & (layer0_outputs[708]);
    assign layer1_outputs[2403] = ~(layer0_outputs[2431]);
    assign layer1_outputs[2404] = ~(layer0_outputs[1545]);
    assign layer1_outputs[2405] = ~(layer0_outputs[1374]) | (layer0_outputs[1181]);
    assign layer1_outputs[2406] = ~((layer0_outputs[2411]) | (layer0_outputs[2484]));
    assign layer1_outputs[2407] = layer0_outputs[1575];
    assign layer1_outputs[2408] = ~((layer0_outputs[1963]) | (layer0_outputs[1641]));
    assign layer1_outputs[2409] = layer0_outputs[1153];
    assign layer1_outputs[2410] = layer0_outputs[1089];
    assign layer1_outputs[2411] = layer0_outputs[2403];
    assign layer1_outputs[2412] = (layer0_outputs[419]) & ~(layer0_outputs[518]);
    assign layer1_outputs[2413] = ~(layer0_outputs[569]) | (layer0_outputs[482]);
    assign layer1_outputs[2414] = (layer0_outputs[2143]) | (layer0_outputs[1551]);
    assign layer1_outputs[2415] = ~(layer0_outputs[1462]);
    assign layer1_outputs[2416] = ~(layer0_outputs[1022]);
    assign layer1_outputs[2417] = layer0_outputs[613];
    assign layer1_outputs[2418] = (layer0_outputs[2357]) | (layer0_outputs[1195]);
    assign layer1_outputs[2419] = ~(layer0_outputs[2161]) | (layer0_outputs[417]);
    assign layer1_outputs[2420] = ~((layer0_outputs[2307]) | (layer0_outputs[1994]));
    assign layer1_outputs[2421] = ~((layer0_outputs[1026]) | (layer0_outputs[1133]));
    assign layer1_outputs[2422] = layer0_outputs[1699];
    assign layer1_outputs[2423] = (layer0_outputs[2385]) & ~(layer0_outputs[1468]);
    assign layer1_outputs[2424] = ~((layer0_outputs[2121]) ^ (layer0_outputs[258]));
    assign layer1_outputs[2425] = ~(layer0_outputs[1237]) | (layer0_outputs[21]);
    assign layer1_outputs[2426] = (layer0_outputs[823]) & (layer0_outputs[1351]);
    assign layer1_outputs[2427] = 1'b1;
    assign layer1_outputs[2428] = layer0_outputs[1760];
    assign layer1_outputs[2429] = layer0_outputs[1260];
    assign layer1_outputs[2430] = ~(layer0_outputs[1614]);
    assign layer1_outputs[2431] = layer0_outputs[2251];
    assign layer1_outputs[2432] = (layer0_outputs[0]) & ~(layer0_outputs[739]);
    assign layer1_outputs[2433] = ~((layer0_outputs[1319]) | (layer0_outputs[745]));
    assign layer1_outputs[2434] = (layer0_outputs[437]) | (layer0_outputs[845]);
    assign layer1_outputs[2435] = ~((layer0_outputs[874]) | (layer0_outputs[1938]));
    assign layer1_outputs[2436] = ~(layer0_outputs[2017]);
    assign layer1_outputs[2437] = ~(layer0_outputs[1208]) | (layer0_outputs[632]);
    assign layer1_outputs[2438] = layer0_outputs[2319];
    assign layer1_outputs[2439] = ~(layer0_outputs[1512]);
    assign layer1_outputs[2440] = ~(layer0_outputs[1328]) | (layer0_outputs[2463]);
    assign layer1_outputs[2441] = layer0_outputs[1509];
    assign layer1_outputs[2442] = (layer0_outputs[2284]) | (layer0_outputs[1888]);
    assign layer1_outputs[2443] = (layer0_outputs[2008]) | (layer0_outputs[1536]);
    assign layer1_outputs[2444] = 1'b0;
    assign layer1_outputs[2445] = ~(layer0_outputs[2317]) | (layer0_outputs[1661]);
    assign layer1_outputs[2446] = ~((layer0_outputs[1404]) | (layer0_outputs[1350]));
    assign layer1_outputs[2447] = (layer0_outputs[1438]) & ~(layer0_outputs[1333]);
    assign layer1_outputs[2448] = ~(layer0_outputs[415]) | (layer0_outputs[604]);
    assign layer1_outputs[2449] = ~(layer0_outputs[2148]) | (layer0_outputs[552]);
    assign layer1_outputs[2450] = ~(layer0_outputs[2109]) | (layer0_outputs[1927]);
    assign layer1_outputs[2451] = layer0_outputs[2218];
    assign layer1_outputs[2452] = (layer0_outputs[1459]) & ~(layer0_outputs[1344]);
    assign layer1_outputs[2453] = ~(layer0_outputs[54]) | (layer0_outputs[2409]);
    assign layer1_outputs[2454] = (layer0_outputs[150]) & ~(layer0_outputs[1079]);
    assign layer1_outputs[2455] = ~((layer0_outputs[2023]) & (layer0_outputs[1618]));
    assign layer1_outputs[2456] = 1'b0;
    assign layer1_outputs[2457] = 1'b0;
    assign layer1_outputs[2458] = (layer0_outputs[1660]) & ~(layer0_outputs[336]);
    assign layer1_outputs[2459] = ~((layer0_outputs[276]) | (layer0_outputs[634]));
    assign layer1_outputs[2460] = ~((layer0_outputs[845]) & (layer0_outputs[1558]));
    assign layer1_outputs[2461] = 1'b0;
    assign layer1_outputs[2462] = ~(layer0_outputs[1486]);
    assign layer1_outputs[2463] = ~((layer0_outputs[1941]) | (layer0_outputs[2273]));
    assign layer1_outputs[2464] = (layer0_outputs[75]) & (layer0_outputs[936]);
    assign layer1_outputs[2465] = ~(layer0_outputs[2370]) | (layer0_outputs[1269]);
    assign layer1_outputs[2466] = ~((layer0_outputs[280]) & (layer0_outputs[2497]));
    assign layer1_outputs[2467] = ~((layer0_outputs[2538]) | (layer0_outputs[1447]));
    assign layer1_outputs[2468] = ~(layer0_outputs[1477]) | (layer0_outputs[721]);
    assign layer1_outputs[2469] = ~(layer0_outputs[595]) | (layer0_outputs[805]);
    assign layer1_outputs[2470] = ~(layer0_outputs[880]);
    assign layer1_outputs[2471] = (layer0_outputs[748]) & ~(layer0_outputs[1781]);
    assign layer1_outputs[2472] = ~(layer0_outputs[1823]) | (layer0_outputs[1211]);
    assign layer1_outputs[2473] = ~((layer0_outputs[1001]) & (layer0_outputs[540]));
    assign layer1_outputs[2474] = ~(layer0_outputs[424]) | (layer0_outputs[2396]);
    assign layer1_outputs[2475] = ~(layer0_outputs[1552]);
    assign layer1_outputs[2476] = ~((layer0_outputs[2523]) ^ (layer0_outputs[245]));
    assign layer1_outputs[2477] = (layer0_outputs[1799]) & (layer0_outputs[2050]);
    assign layer1_outputs[2478] = 1'b0;
    assign layer1_outputs[2479] = layer0_outputs[2078];
    assign layer1_outputs[2480] = ~(layer0_outputs[1035]) | (layer0_outputs[1866]);
    assign layer1_outputs[2481] = ~(layer0_outputs[1080]) | (layer0_outputs[2232]);
    assign layer1_outputs[2482] = ~(layer0_outputs[1712]) | (layer0_outputs[1703]);
    assign layer1_outputs[2483] = (layer0_outputs[1786]) & ~(layer0_outputs[648]);
    assign layer1_outputs[2484] = ~((layer0_outputs[458]) | (layer0_outputs[642]));
    assign layer1_outputs[2485] = layer0_outputs[1697];
    assign layer1_outputs[2486] = (layer0_outputs[399]) | (layer0_outputs[514]);
    assign layer1_outputs[2487] = ~(layer0_outputs[1670]);
    assign layer1_outputs[2488] = ~(layer0_outputs[101]);
    assign layer1_outputs[2489] = layer0_outputs[1442];
    assign layer1_outputs[2490] = layer0_outputs[2203];
    assign layer1_outputs[2491] = (layer0_outputs[2100]) & ~(layer0_outputs[1074]);
    assign layer1_outputs[2492] = (layer0_outputs[2494]) & ~(layer0_outputs[836]);
    assign layer1_outputs[2493] = ~((layer0_outputs[2092]) ^ (layer0_outputs[2046]));
    assign layer1_outputs[2494] = layer0_outputs[769];
    assign layer1_outputs[2495] = (layer0_outputs[752]) & ~(layer0_outputs[1568]);
    assign layer1_outputs[2496] = ~(layer0_outputs[365]);
    assign layer1_outputs[2497] = ~(layer0_outputs[1800]) | (layer0_outputs[305]);
    assign layer1_outputs[2498] = layer0_outputs[473];
    assign layer1_outputs[2499] = layer0_outputs[2531];
    assign layer1_outputs[2500] = ~(layer0_outputs[2247]) | (layer0_outputs[1545]);
    assign layer1_outputs[2501] = ~(layer0_outputs[1259]);
    assign layer1_outputs[2502] = (layer0_outputs[920]) & ~(layer0_outputs[159]);
    assign layer1_outputs[2503] = ~(layer0_outputs[2156]) | (layer0_outputs[1972]);
    assign layer1_outputs[2504] = (layer0_outputs[1800]) & ~(layer0_outputs[1782]);
    assign layer1_outputs[2505] = 1'b0;
    assign layer1_outputs[2506] = layer0_outputs[2183];
    assign layer1_outputs[2507] = ~((layer0_outputs[1644]) & (layer0_outputs[2060]));
    assign layer1_outputs[2508] = (layer0_outputs[1933]) & (layer0_outputs[2443]);
    assign layer1_outputs[2509] = layer0_outputs[513];
    assign layer1_outputs[2510] = ~(layer0_outputs[1402]);
    assign layer1_outputs[2511] = ~(layer0_outputs[2255]);
    assign layer1_outputs[2512] = ~(layer0_outputs[1951]) | (layer0_outputs[219]);
    assign layer1_outputs[2513] = ~(layer0_outputs[1539]) | (layer0_outputs[2505]);
    assign layer1_outputs[2514] = (layer0_outputs[994]) & (layer0_outputs[1806]);
    assign layer1_outputs[2515] = 1'b0;
    assign layer1_outputs[2516] = (layer0_outputs[1428]) | (layer0_outputs[670]);
    assign layer1_outputs[2517] = (layer0_outputs[2460]) & ~(layer0_outputs[818]);
    assign layer1_outputs[2518] = (layer0_outputs[1300]) & ~(layer0_outputs[2077]);
    assign layer1_outputs[2519] = 1'b0;
    assign layer1_outputs[2520] = (layer0_outputs[221]) & ~(layer0_outputs[1090]);
    assign layer1_outputs[2521] = (layer0_outputs[243]) | (layer0_outputs[1774]);
    assign layer1_outputs[2522] = ~((layer0_outputs[2191]) | (layer0_outputs[2379]));
    assign layer1_outputs[2523] = ~(layer0_outputs[60]) | (layer0_outputs[1422]);
    assign layer1_outputs[2524] = (layer0_outputs[1768]) ^ (layer0_outputs[1457]);
    assign layer1_outputs[2525] = (layer0_outputs[535]) ^ (layer0_outputs[299]);
    assign layer1_outputs[2526] = (layer0_outputs[813]) & ~(layer0_outputs[1725]);
    assign layer1_outputs[2527] = ~((layer0_outputs[714]) | (layer0_outputs[2195]));
    assign layer1_outputs[2528] = ~((layer0_outputs[2380]) | (layer0_outputs[2107]));
    assign layer1_outputs[2529] = ~(layer0_outputs[1152]);
    assign layer1_outputs[2530] = ~((layer0_outputs[2111]) | (layer0_outputs[973]));
    assign layer1_outputs[2531] = layer0_outputs[119];
    assign layer1_outputs[2532] = ~(layer0_outputs[189]);
    assign layer1_outputs[2533] = ~(layer0_outputs[504]);
    assign layer1_outputs[2534] = ~(layer0_outputs[1467]) | (layer0_outputs[2216]);
    assign layer1_outputs[2535] = ~(layer0_outputs[1979]) | (layer0_outputs[1793]);
    assign layer1_outputs[2536] = 1'b0;
    assign layer1_outputs[2537] = 1'b1;
    assign layer1_outputs[2538] = ~(layer0_outputs[1516]) | (layer0_outputs[1733]);
    assign layer1_outputs[2539] = (layer0_outputs[468]) | (layer0_outputs[496]);
    assign layer1_outputs[2540] = ~(layer0_outputs[2010]);
    assign layer1_outputs[2541] = ~(layer0_outputs[497]) | (layer0_outputs[2554]);
    assign layer1_outputs[2542] = (layer0_outputs[1175]) & (layer0_outputs[2148]);
    assign layer1_outputs[2543] = layer0_outputs[1857];
    assign layer1_outputs[2544] = ~((layer0_outputs[434]) ^ (layer0_outputs[85]));
    assign layer1_outputs[2545] = layer0_outputs[2503];
    assign layer1_outputs[2546] = (layer0_outputs[758]) & ~(layer0_outputs[1318]);
    assign layer1_outputs[2547] = 1'b1;
    assign layer1_outputs[2548] = ~(layer0_outputs[1541]);
    assign layer1_outputs[2549] = 1'b0;
    assign layer1_outputs[2550] = ~((layer0_outputs[261]) ^ (layer0_outputs[1126]));
    assign layer1_outputs[2551] = (layer0_outputs[983]) | (layer0_outputs[2133]);
    assign layer1_outputs[2552] = 1'b1;
    assign layer1_outputs[2553] = ~(layer0_outputs[1658]) | (layer0_outputs[1023]);
    assign layer1_outputs[2554] = ~(layer0_outputs[628]);
    assign layer1_outputs[2555] = (layer0_outputs[128]) | (layer0_outputs[2401]);
    assign layer1_outputs[2556] = ~(layer0_outputs[1783]);
    assign layer1_outputs[2557] = (layer0_outputs[1806]) & ~(layer0_outputs[1412]);
    assign layer1_outputs[2558] = ~(layer0_outputs[1494]);
    assign layer1_outputs[2559] = ~(layer0_outputs[1839]);
    assign layer2_outputs[0] = 1'b1;
    assign layer2_outputs[1] = (layer1_outputs[1214]) | (layer1_outputs[586]);
    assign layer2_outputs[2] = ~(layer1_outputs[2072]);
    assign layer2_outputs[3] = (layer1_outputs[242]) | (layer1_outputs[1106]);
    assign layer2_outputs[4] = layer1_outputs[260];
    assign layer2_outputs[5] = ~((layer1_outputs[8]) & (layer1_outputs[1862]));
    assign layer2_outputs[6] = layer1_outputs[1897];
    assign layer2_outputs[7] = layer1_outputs[1330];
    assign layer2_outputs[8] = ~(layer1_outputs[2386]) | (layer1_outputs[642]);
    assign layer2_outputs[9] = layer1_outputs[797];
    assign layer2_outputs[10] = layer1_outputs[1821];
    assign layer2_outputs[11] = ~(layer1_outputs[1930]);
    assign layer2_outputs[12] = ~((layer1_outputs[1857]) | (layer1_outputs[717]));
    assign layer2_outputs[13] = (layer1_outputs[1553]) & ~(layer1_outputs[429]);
    assign layer2_outputs[14] = layer1_outputs[540];
    assign layer2_outputs[15] = ~(layer1_outputs[32]);
    assign layer2_outputs[16] = (layer1_outputs[2179]) & ~(layer1_outputs[2189]);
    assign layer2_outputs[17] = ~((layer1_outputs[1829]) | (layer1_outputs[215]));
    assign layer2_outputs[18] = layer1_outputs[950];
    assign layer2_outputs[19] = 1'b1;
    assign layer2_outputs[20] = ~(layer1_outputs[2255]) | (layer1_outputs[2158]);
    assign layer2_outputs[21] = (layer1_outputs[718]) & ~(layer1_outputs[158]);
    assign layer2_outputs[22] = (layer1_outputs[506]) & ~(layer1_outputs[1474]);
    assign layer2_outputs[23] = ~((layer1_outputs[835]) ^ (layer1_outputs[11]));
    assign layer2_outputs[24] = ~((layer1_outputs[1262]) | (layer1_outputs[1124]));
    assign layer2_outputs[25] = ~((layer1_outputs[2391]) & (layer1_outputs[2137]));
    assign layer2_outputs[26] = ~((layer1_outputs[974]) & (layer1_outputs[1354]));
    assign layer2_outputs[27] = (layer1_outputs[2116]) & (layer1_outputs[1]);
    assign layer2_outputs[28] = ~(layer1_outputs[333]) | (layer1_outputs[2504]);
    assign layer2_outputs[29] = ~((layer1_outputs[938]) ^ (layer1_outputs[2292]));
    assign layer2_outputs[30] = layer1_outputs[1900];
    assign layer2_outputs[31] = layer1_outputs[1503];
    assign layer2_outputs[32] = ~(layer1_outputs[2541]);
    assign layer2_outputs[33] = ~(layer1_outputs[2108]);
    assign layer2_outputs[34] = ~(layer1_outputs[127]) | (layer1_outputs[508]);
    assign layer2_outputs[35] = ~(layer1_outputs[1606]) | (layer1_outputs[594]);
    assign layer2_outputs[36] = ~(layer1_outputs[2506]);
    assign layer2_outputs[37] = 1'b0;
    assign layer2_outputs[38] = ~(layer1_outputs[846]) | (layer1_outputs[2474]);
    assign layer2_outputs[39] = (layer1_outputs[703]) | (layer1_outputs[1027]);
    assign layer2_outputs[40] = 1'b0;
    assign layer2_outputs[41] = ~(layer1_outputs[986]) | (layer1_outputs[362]);
    assign layer2_outputs[42] = ~(layer1_outputs[1146]);
    assign layer2_outputs[43] = 1'b0;
    assign layer2_outputs[44] = 1'b0;
    assign layer2_outputs[45] = ~(layer1_outputs[1864]);
    assign layer2_outputs[46] = ~(layer1_outputs[2501]) | (layer1_outputs[994]);
    assign layer2_outputs[47] = 1'b1;
    assign layer2_outputs[48] = ~(layer1_outputs[2526]);
    assign layer2_outputs[49] = (layer1_outputs[47]) ^ (layer1_outputs[1185]);
    assign layer2_outputs[50] = ~((layer1_outputs[118]) | (layer1_outputs[1752]));
    assign layer2_outputs[51] = 1'b1;
    assign layer2_outputs[52] = ~((layer1_outputs[803]) & (layer1_outputs[710]));
    assign layer2_outputs[53] = (layer1_outputs[1408]) | (layer1_outputs[906]);
    assign layer2_outputs[54] = layer1_outputs[1979];
    assign layer2_outputs[55] = 1'b0;
    assign layer2_outputs[56] = layer1_outputs[2364];
    assign layer2_outputs[57] = ~(layer1_outputs[1290]);
    assign layer2_outputs[58] = ~(layer1_outputs[2017]) | (layer1_outputs[501]);
    assign layer2_outputs[59] = ~((layer1_outputs[2090]) ^ (layer1_outputs[1713]));
    assign layer2_outputs[60] = (layer1_outputs[1848]) & ~(layer1_outputs[1837]);
    assign layer2_outputs[61] = ~(layer1_outputs[2245]);
    assign layer2_outputs[62] = (layer1_outputs[2239]) & ~(layer1_outputs[1650]);
    assign layer2_outputs[63] = layer1_outputs[513];
    assign layer2_outputs[64] = layer1_outputs[1582];
    assign layer2_outputs[65] = (layer1_outputs[4]) & (layer1_outputs[2491]);
    assign layer2_outputs[66] = 1'b1;
    assign layer2_outputs[67] = layer1_outputs[779];
    assign layer2_outputs[68] = 1'b0;
    assign layer2_outputs[69] = ~(layer1_outputs[72]);
    assign layer2_outputs[70] = ~(layer1_outputs[2353]) | (layer1_outputs[2409]);
    assign layer2_outputs[71] = layer1_outputs[1453];
    assign layer2_outputs[72] = layer1_outputs[2117];
    assign layer2_outputs[73] = 1'b1;
    assign layer2_outputs[74] = ~(layer1_outputs[1285]) | (layer1_outputs[94]);
    assign layer2_outputs[75] = 1'b0;
    assign layer2_outputs[76] = (layer1_outputs[1550]) & (layer1_outputs[1418]);
    assign layer2_outputs[77] = ~(layer1_outputs[1440]);
    assign layer2_outputs[78] = ~((layer1_outputs[190]) | (layer1_outputs[1233]));
    assign layer2_outputs[79] = ~((layer1_outputs[1756]) | (layer1_outputs[2478]));
    assign layer2_outputs[80] = ~((layer1_outputs[781]) | (layer1_outputs[2118]));
    assign layer2_outputs[81] = ~(layer1_outputs[832]);
    assign layer2_outputs[82] = (layer1_outputs[1959]) & ~(layer1_outputs[420]);
    assign layer2_outputs[83] = ~(layer1_outputs[2103]) | (layer1_outputs[68]);
    assign layer2_outputs[84] = ~(layer1_outputs[457]);
    assign layer2_outputs[85] = ~(layer1_outputs[2250]);
    assign layer2_outputs[86] = (layer1_outputs[964]) & ~(layer1_outputs[1776]);
    assign layer2_outputs[87] = ~(layer1_outputs[467]) | (layer1_outputs[1651]);
    assign layer2_outputs[88] = layer1_outputs[1476];
    assign layer2_outputs[89] = ~((layer1_outputs[1682]) | (layer1_outputs[1590]));
    assign layer2_outputs[90] = layer1_outputs[1643];
    assign layer2_outputs[91] = ~(layer1_outputs[2228]) | (layer1_outputs[2070]);
    assign layer2_outputs[92] = (layer1_outputs[305]) & ~(layer1_outputs[277]);
    assign layer2_outputs[93] = ~(layer1_outputs[1516]);
    assign layer2_outputs[94] = layer1_outputs[410];
    assign layer2_outputs[95] = ~(layer1_outputs[41]) | (layer1_outputs[1347]);
    assign layer2_outputs[96] = 1'b0;
    assign layer2_outputs[97] = 1'b1;
    assign layer2_outputs[98] = layer1_outputs[270];
    assign layer2_outputs[99] = 1'b1;
    assign layer2_outputs[100] = 1'b1;
    assign layer2_outputs[101] = layer1_outputs[2175];
    assign layer2_outputs[102] = 1'b1;
    assign layer2_outputs[103] = (layer1_outputs[1387]) & (layer1_outputs[349]);
    assign layer2_outputs[104] = layer1_outputs[1696];
    assign layer2_outputs[105] = 1'b1;
    assign layer2_outputs[106] = (layer1_outputs[1136]) & (layer1_outputs[1833]);
    assign layer2_outputs[107] = 1'b0;
    assign layer2_outputs[108] = (layer1_outputs[1902]) | (layer1_outputs[2456]);
    assign layer2_outputs[109] = (layer1_outputs[1951]) & (layer1_outputs[530]);
    assign layer2_outputs[110] = layer1_outputs[1075];
    assign layer2_outputs[111] = ~(layer1_outputs[1747]);
    assign layer2_outputs[112] = layer1_outputs[440];
    assign layer2_outputs[113] = layer1_outputs[2414];
    assign layer2_outputs[114] = (layer1_outputs[444]) ^ (layer1_outputs[1323]);
    assign layer2_outputs[115] = ~(layer1_outputs[306]) | (layer1_outputs[567]);
    assign layer2_outputs[116] = (layer1_outputs[206]) & (layer1_outputs[1877]);
    assign layer2_outputs[117] = (layer1_outputs[937]) & ~(layer1_outputs[2538]);
    assign layer2_outputs[118] = ~(layer1_outputs[226]);
    assign layer2_outputs[119] = layer1_outputs[2363];
    assign layer2_outputs[120] = ~(layer1_outputs[1039]) | (layer1_outputs[91]);
    assign layer2_outputs[121] = ~((layer1_outputs[1112]) ^ (layer1_outputs[1486]));
    assign layer2_outputs[122] = ~((layer1_outputs[870]) ^ (layer1_outputs[1279]));
    assign layer2_outputs[123] = ~((layer1_outputs[142]) | (layer1_outputs[1858]));
    assign layer2_outputs[124] = (layer1_outputs[358]) & ~(layer1_outputs[1871]);
    assign layer2_outputs[125] = ~(layer1_outputs[1431]) | (layer1_outputs[2313]);
    assign layer2_outputs[126] = ~(layer1_outputs[681]);
    assign layer2_outputs[127] = ~(layer1_outputs[1404]);
    assign layer2_outputs[128] = 1'b1;
    assign layer2_outputs[129] = ~((layer1_outputs[1220]) | (layer1_outputs[1925]));
    assign layer2_outputs[130] = ~((layer1_outputs[1134]) & (layer1_outputs[1727]));
    assign layer2_outputs[131] = ~(layer1_outputs[1647]);
    assign layer2_outputs[132] = layer1_outputs[1081];
    assign layer2_outputs[133] = ~((layer1_outputs[2001]) & (layer1_outputs[313]));
    assign layer2_outputs[134] = ~(layer1_outputs[2110]);
    assign layer2_outputs[135] = (layer1_outputs[2480]) & ~(layer1_outputs[592]);
    assign layer2_outputs[136] = ~(layer1_outputs[1012]) | (layer1_outputs[984]);
    assign layer2_outputs[137] = 1'b0;
    assign layer2_outputs[138] = (layer1_outputs[1863]) ^ (layer1_outputs[1196]);
    assign layer2_outputs[139] = (layer1_outputs[2399]) & (layer1_outputs[2010]);
    assign layer2_outputs[140] = ~(layer1_outputs[917]);
    assign layer2_outputs[141] = layer1_outputs[963];
    assign layer2_outputs[142] = ~(layer1_outputs[803]);
    assign layer2_outputs[143] = ~((layer1_outputs[1092]) ^ (layer1_outputs[741]));
    assign layer2_outputs[144] = (layer1_outputs[2184]) & ~(layer1_outputs[521]);
    assign layer2_outputs[145] = ~((layer1_outputs[2346]) & (layer1_outputs[589]));
    assign layer2_outputs[146] = ~(layer1_outputs[2217]) | (layer1_outputs[632]);
    assign layer2_outputs[147] = layer1_outputs[1469];
    assign layer2_outputs[148] = 1'b0;
    assign layer2_outputs[149] = ~(layer1_outputs[581]) | (layer1_outputs[2092]);
    assign layer2_outputs[150] = (layer1_outputs[325]) & ~(layer1_outputs[1778]);
    assign layer2_outputs[151] = layer1_outputs[2002];
    assign layer2_outputs[152] = ~((layer1_outputs[1643]) | (layer1_outputs[1736]));
    assign layer2_outputs[153] = (layer1_outputs[2002]) | (layer1_outputs[314]);
    assign layer2_outputs[154] = (layer1_outputs[444]) | (layer1_outputs[920]);
    assign layer2_outputs[155] = (layer1_outputs[297]) & (layer1_outputs[607]);
    assign layer2_outputs[156] = ~(layer1_outputs[1987]);
    assign layer2_outputs[157] = layer1_outputs[1099];
    assign layer2_outputs[158] = ~((layer1_outputs[2251]) | (layer1_outputs[1155]));
    assign layer2_outputs[159] = ~(layer1_outputs[838]);
    assign layer2_outputs[160] = ~(layer1_outputs[2369]);
    assign layer2_outputs[161] = ~((layer1_outputs[358]) & (layer1_outputs[2157]));
    assign layer2_outputs[162] = layer1_outputs[2151];
    assign layer2_outputs[163] = layer1_outputs[724];
    assign layer2_outputs[164] = (layer1_outputs[526]) & ~(layer1_outputs[986]);
    assign layer2_outputs[165] = layer1_outputs[265];
    assign layer2_outputs[166] = (layer1_outputs[1076]) & ~(layer1_outputs[1859]);
    assign layer2_outputs[167] = (layer1_outputs[640]) & (layer1_outputs[2058]);
    assign layer2_outputs[168] = ~((layer1_outputs[1825]) | (layer1_outputs[680]));
    assign layer2_outputs[169] = (layer1_outputs[1102]) & ~(layer1_outputs[2497]);
    assign layer2_outputs[170] = ~(layer1_outputs[323]);
    assign layer2_outputs[171] = 1'b0;
    assign layer2_outputs[172] = layer1_outputs[2064];
    assign layer2_outputs[173] = ~(layer1_outputs[2288]);
    assign layer2_outputs[174] = layer1_outputs[1296];
    assign layer2_outputs[175] = ~(layer1_outputs[2233]);
    assign layer2_outputs[176] = ~(layer1_outputs[2384]);
    assign layer2_outputs[177] = 1'b0;
    assign layer2_outputs[178] = (layer1_outputs[2287]) & ~(layer1_outputs[749]);
    assign layer2_outputs[179] = layer1_outputs[1809];
    assign layer2_outputs[180] = ~(layer1_outputs[273]) | (layer1_outputs[220]);
    assign layer2_outputs[181] = (layer1_outputs[1137]) ^ (layer1_outputs[977]);
    assign layer2_outputs[182] = (layer1_outputs[1177]) & ~(layer1_outputs[1808]);
    assign layer2_outputs[183] = ~(layer1_outputs[2264]);
    assign layer2_outputs[184] = (layer1_outputs[762]) ^ (layer1_outputs[411]);
    assign layer2_outputs[185] = layer1_outputs[258];
    assign layer2_outputs[186] = layer1_outputs[681];
    assign layer2_outputs[187] = (layer1_outputs[504]) & ~(layer1_outputs[932]);
    assign layer2_outputs[188] = ~(layer1_outputs[903]) | (layer1_outputs[2023]);
    assign layer2_outputs[189] = 1'b1;
    assign layer2_outputs[190] = ~(layer1_outputs[1840]);
    assign layer2_outputs[191] = (layer1_outputs[1509]) & ~(layer1_outputs[1138]);
    assign layer2_outputs[192] = ~(layer1_outputs[1456]) | (layer1_outputs[808]);
    assign layer2_outputs[193] = ~(layer1_outputs[2062]);
    assign layer2_outputs[194] = (layer1_outputs[279]) & ~(layer1_outputs[1567]);
    assign layer2_outputs[195] = 1'b1;
    assign layer2_outputs[196] = ~(layer1_outputs[306]);
    assign layer2_outputs[197] = ~(layer1_outputs[2542]);
    assign layer2_outputs[198] = (layer1_outputs[1918]) & ~(layer1_outputs[814]);
    assign layer2_outputs[199] = (layer1_outputs[2300]) | (layer1_outputs[1578]);
    assign layer2_outputs[200] = ~((layer1_outputs[2408]) & (layer1_outputs[1263]));
    assign layer2_outputs[201] = ~((layer1_outputs[590]) ^ (layer1_outputs[850]));
    assign layer2_outputs[202] = layer1_outputs[80];
    assign layer2_outputs[203] = ~(layer1_outputs[1390]);
    assign layer2_outputs[204] = 1'b0;
    assign layer2_outputs[205] = layer1_outputs[829];
    assign layer2_outputs[206] = ~(layer1_outputs[120]);
    assign layer2_outputs[207] = (layer1_outputs[796]) & ~(layer1_outputs[871]);
    assign layer2_outputs[208] = (layer1_outputs[840]) | (layer1_outputs[1114]);
    assign layer2_outputs[209] = ~((layer1_outputs[2328]) & (layer1_outputs[1720]));
    assign layer2_outputs[210] = (layer1_outputs[1195]) & ~(layer1_outputs[1146]);
    assign layer2_outputs[211] = (layer1_outputs[1856]) & ~(layer1_outputs[2363]);
    assign layer2_outputs[212] = ~(layer1_outputs[149]);
    assign layer2_outputs[213] = ~(layer1_outputs[1082]) | (layer1_outputs[46]);
    assign layer2_outputs[214] = ~(layer1_outputs[359]);
    assign layer2_outputs[215] = ~(layer1_outputs[1444]);
    assign layer2_outputs[216] = ~(layer1_outputs[2330]);
    assign layer2_outputs[217] = 1'b1;
    assign layer2_outputs[218] = (layer1_outputs[89]) & ~(layer1_outputs[1946]);
    assign layer2_outputs[219] = (layer1_outputs[1943]) & ~(layer1_outputs[109]);
    assign layer2_outputs[220] = ~(layer1_outputs[225]) | (layer1_outputs[1256]);
    assign layer2_outputs[221] = 1'b1;
    assign layer2_outputs[222] = 1'b1;
    assign layer2_outputs[223] = ~(layer1_outputs[1001]);
    assign layer2_outputs[224] = layer1_outputs[580];
    assign layer2_outputs[225] = layer1_outputs[934];
    assign layer2_outputs[226] = layer1_outputs[1808];
    assign layer2_outputs[227] = 1'b1;
    assign layer2_outputs[228] = 1'b1;
    assign layer2_outputs[229] = ~((layer1_outputs[1295]) | (layer1_outputs[1492]));
    assign layer2_outputs[230] = ~(layer1_outputs[1972]);
    assign layer2_outputs[231] = (layer1_outputs[1180]) & (layer1_outputs[771]);
    assign layer2_outputs[232] = layer1_outputs[393];
    assign layer2_outputs[233] = layer1_outputs[2559];
    assign layer2_outputs[234] = layer1_outputs[2496];
    assign layer2_outputs[235] = layer1_outputs[517];
    assign layer2_outputs[236] = (layer1_outputs[463]) | (layer1_outputs[1489]);
    assign layer2_outputs[237] = ~((layer1_outputs[2252]) | (layer1_outputs[2030]));
    assign layer2_outputs[238] = ~(layer1_outputs[1952]) | (layer1_outputs[826]);
    assign layer2_outputs[239] = ~((layer1_outputs[1122]) & (layer1_outputs[1625]));
    assign layer2_outputs[240] = ~(layer1_outputs[963]);
    assign layer2_outputs[241] = layer1_outputs[1442];
    assign layer2_outputs[242] = ~(layer1_outputs[1568]) | (layer1_outputs[184]);
    assign layer2_outputs[243] = ~((layer1_outputs[2333]) & (layer1_outputs[845]));
    assign layer2_outputs[244] = ~((layer1_outputs[1938]) ^ (layer1_outputs[1759]));
    assign layer2_outputs[245] = ~(layer1_outputs[1490]);
    assign layer2_outputs[246] = ~(layer1_outputs[914]);
    assign layer2_outputs[247] = ~(layer1_outputs[2380]);
    assign layer2_outputs[248] = (layer1_outputs[2152]) & (layer1_outputs[2558]);
    assign layer2_outputs[249] = ~(layer1_outputs[1390]);
    assign layer2_outputs[250] = layer1_outputs[1246];
    assign layer2_outputs[251] = ~((layer1_outputs[603]) ^ (layer1_outputs[1906]));
    assign layer2_outputs[252] = (layer1_outputs[1676]) & ~(layer1_outputs[1127]);
    assign layer2_outputs[253] = 1'b1;
    assign layer2_outputs[254] = layer1_outputs[15];
    assign layer2_outputs[255] = layer1_outputs[193];
    assign layer2_outputs[256] = (layer1_outputs[1077]) & ~(layer1_outputs[1207]);
    assign layer2_outputs[257] = (layer1_outputs[2254]) & (layer1_outputs[2506]);
    assign layer2_outputs[258] = 1'b1;
    assign layer2_outputs[259] = layer1_outputs[2283];
    assign layer2_outputs[260] = ~(layer1_outputs[1190]);
    assign layer2_outputs[261] = ~(layer1_outputs[967]);
    assign layer2_outputs[262] = (layer1_outputs[2099]) & ~(layer1_outputs[1993]);
    assign layer2_outputs[263] = ~(layer1_outputs[1955]);
    assign layer2_outputs[264] = ~(layer1_outputs[1936]) | (layer1_outputs[1691]);
    assign layer2_outputs[265] = layer1_outputs[156];
    assign layer2_outputs[266] = (layer1_outputs[2547]) & ~(layer1_outputs[1660]);
    assign layer2_outputs[267] = layer1_outputs[2317];
    assign layer2_outputs[268] = (layer1_outputs[2397]) & ~(layer1_outputs[1469]);
    assign layer2_outputs[269] = ~(layer1_outputs[2]) | (layer1_outputs[636]);
    assign layer2_outputs[270] = 1'b0;
    assign layer2_outputs[271] = (layer1_outputs[1856]) & ~(layer1_outputs[815]);
    assign layer2_outputs[272] = 1'b1;
    assign layer2_outputs[273] = (layer1_outputs[2052]) & ~(layer1_outputs[2459]);
    assign layer2_outputs[274] = layer1_outputs[2425];
    assign layer2_outputs[275] = (layer1_outputs[2220]) & ~(layer1_outputs[2135]);
    assign layer2_outputs[276] = layer1_outputs[2368];
    assign layer2_outputs[277] = (layer1_outputs[2372]) & ~(layer1_outputs[120]);
    assign layer2_outputs[278] = ~((layer1_outputs[712]) & (layer1_outputs[1105]));
    assign layer2_outputs[279] = (layer1_outputs[971]) & (layer1_outputs[2068]);
    assign layer2_outputs[280] = ~(layer1_outputs[2125]);
    assign layer2_outputs[281] = ~(layer1_outputs[327]);
    assign layer2_outputs[282] = layer1_outputs[239];
    assign layer2_outputs[283] = (layer1_outputs[1851]) & ~(layer1_outputs[648]);
    assign layer2_outputs[284] = ~(layer1_outputs[1178]);
    assign layer2_outputs[285] = (layer1_outputs[1066]) | (layer1_outputs[1035]);
    assign layer2_outputs[286] = ~(layer1_outputs[352]);
    assign layer2_outputs[287] = (layer1_outputs[1667]) & ~(layer1_outputs[1770]);
    assign layer2_outputs[288] = ~(layer1_outputs[1379]);
    assign layer2_outputs[289] = layer1_outputs[1103];
    assign layer2_outputs[290] = layer1_outputs[1898];
    assign layer2_outputs[291] = layer1_outputs[684];
    assign layer2_outputs[292] = (layer1_outputs[1644]) & (layer1_outputs[977]);
    assign layer2_outputs[293] = layer1_outputs[314];
    assign layer2_outputs[294] = ~(layer1_outputs[299]);
    assign layer2_outputs[295] = ~(layer1_outputs[194]);
    assign layer2_outputs[296] = (layer1_outputs[2076]) & (layer1_outputs[1815]);
    assign layer2_outputs[297] = ~(layer1_outputs[1629]);
    assign layer2_outputs[298] = (layer1_outputs[1868]) & ~(layer1_outputs[599]);
    assign layer2_outputs[299] = (layer1_outputs[1127]) & ~(layer1_outputs[1734]);
    assign layer2_outputs[300] = (layer1_outputs[296]) & ~(layer1_outputs[1592]);
    assign layer2_outputs[301] = 1'b1;
    assign layer2_outputs[302] = 1'b1;
    assign layer2_outputs[303] = ~(layer1_outputs[2208]);
    assign layer2_outputs[304] = (layer1_outputs[653]) & (layer1_outputs[1806]);
    assign layer2_outputs[305] = (layer1_outputs[1684]) | (layer1_outputs[1194]);
    assign layer2_outputs[306] = ~((layer1_outputs[2093]) & (layer1_outputs[2129]));
    assign layer2_outputs[307] = layer1_outputs[1391];
    assign layer2_outputs[308] = 1'b1;
    assign layer2_outputs[309] = layer1_outputs[2380];
    assign layer2_outputs[310] = 1'b1;
    assign layer2_outputs[311] = ~(layer1_outputs[101]);
    assign layer2_outputs[312] = (layer1_outputs[334]) & ~(layer1_outputs[1454]);
    assign layer2_outputs[313] = (layer1_outputs[1542]) | (layer1_outputs[1271]);
    assign layer2_outputs[314] = ~((layer1_outputs[1865]) & (layer1_outputs[2166]));
    assign layer2_outputs[315] = (layer1_outputs[1072]) | (layer1_outputs[1368]);
    assign layer2_outputs[316] = ~((layer1_outputs[722]) & (layer1_outputs[2032]));
    assign layer2_outputs[317] = (layer1_outputs[1799]) & ~(layer1_outputs[2475]);
    assign layer2_outputs[318] = 1'b1;
    assign layer2_outputs[319] = ~(layer1_outputs[1874]);
    assign layer2_outputs[320] = ~(layer1_outputs[827]) | (layer1_outputs[774]);
    assign layer2_outputs[321] = (layer1_outputs[1367]) & ~(layer1_outputs[825]);
    assign layer2_outputs[322] = layer1_outputs[2555];
    assign layer2_outputs[323] = ~(layer1_outputs[1818]) | (layer1_outputs[908]);
    assign layer2_outputs[324] = (layer1_outputs[2448]) & ~(layer1_outputs[2389]);
    assign layer2_outputs[325] = ~(layer1_outputs[2221]);
    assign layer2_outputs[326] = layer1_outputs[1698];
    assign layer2_outputs[327] = (layer1_outputs[1508]) & ~(layer1_outputs[2418]);
    assign layer2_outputs[328] = ~(layer1_outputs[181]);
    assign layer2_outputs[329] = (layer1_outputs[1156]) ^ (layer1_outputs[2047]);
    assign layer2_outputs[330] = ~(layer1_outputs[529]);
    assign layer2_outputs[331] = layer1_outputs[2209];
    assign layer2_outputs[332] = (layer1_outputs[1032]) | (layer1_outputs[493]);
    assign layer2_outputs[333] = ~((layer1_outputs[1545]) | (layer1_outputs[1095]));
    assign layer2_outputs[334] = ~(layer1_outputs[1855]);
    assign layer2_outputs[335] = (layer1_outputs[1626]) | (layer1_outputs[293]);
    assign layer2_outputs[336] = ~((layer1_outputs[1754]) | (layer1_outputs[33]));
    assign layer2_outputs[337] = layer1_outputs[1649];
    assign layer2_outputs[338] = 1'b1;
    assign layer2_outputs[339] = layer1_outputs[673];
    assign layer2_outputs[340] = (layer1_outputs[290]) & (layer1_outputs[328]);
    assign layer2_outputs[341] = (layer1_outputs[1679]) & ~(layer1_outputs[1022]);
    assign layer2_outputs[342] = layer1_outputs[1423];
    assign layer2_outputs[343] = layer1_outputs[1212];
    assign layer2_outputs[344] = ~(layer1_outputs[852]);
    assign layer2_outputs[345] = ~(layer1_outputs[2528]) | (layer1_outputs[2067]);
    assign layer2_outputs[346] = ~((layer1_outputs[1131]) | (layer1_outputs[737]));
    assign layer2_outputs[347] = layer1_outputs[2027];
    assign layer2_outputs[348] = 1'b1;
    assign layer2_outputs[349] = ~(layer1_outputs[151]) | (layer1_outputs[2146]);
    assign layer2_outputs[350] = 1'b1;
    assign layer2_outputs[351] = layer1_outputs[219];
    assign layer2_outputs[352] = ~(layer1_outputs[2059]);
    assign layer2_outputs[353] = (layer1_outputs[1655]) & ~(layer1_outputs[1628]);
    assign layer2_outputs[354] = ~((layer1_outputs[837]) & (layer1_outputs[702]));
    assign layer2_outputs[355] = layer1_outputs[172];
    assign layer2_outputs[356] = 1'b1;
    assign layer2_outputs[357] = (layer1_outputs[1520]) | (layer1_outputs[1796]);
    assign layer2_outputs[358] = layer1_outputs[2361];
    assign layer2_outputs[359] = ~(layer1_outputs[1245]);
    assign layer2_outputs[360] = ~(layer1_outputs[1997]);
    assign layer2_outputs[361] = ~((layer1_outputs[2098]) | (layer1_outputs[1505]));
    assign layer2_outputs[362] = ~((layer1_outputs[212]) & (layer1_outputs[1801]));
    assign layer2_outputs[363] = layer1_outputs[2231];
    assign layer2_outputs[364] = ~(layer1_outputs[1097]);
    assign layer2_outputs[365] = ~((layer1_outputs[1664]) | (layer1_outputs[2193]));
    assign layer2_outputs[366] = ~(layer1_outputs[1169]) | (layer1_outputs[1623]);
    assign layer2_outputs[367] = layer1_outputs[795];
    assign layer2_outputs[368] = ~((layer1_outputs[471]) | (layer1_outputs[812]));
    assign layer2_outputs[369] = 1'b0;
    assign layer2_outputs[370] = (layer1_outputs[1211]) & (layer1_outputs[1620]);
    assign layer2_outputs[371] = ~(layer1_outputs[1143]) | (layer1_outputs[922]);
    assign layer2_outputs[372] = ~((layer1_outputs[1334]) ^ (layer1_outputs[1949]));
    assign layer2_outputs[373] = layer1_outputs[116];
    assign layer2_outputs[374] = 1'b1;
    assign layer2_outputs[375] = ~(layer1_outputs[304]);
    assign layer2_outputs[376] = ~((layer1_outputs[2301]) | (layer1_outputs[2282]));
    assign layer2_outputs[377] = ~(layer1_outputs[891]);
    assign layer2_outputs[378] = ~(layer1_outputs[2370]);
    assign layer2_outputs[379] = layer1_outputs[1446];
    assign layer2_outputs[380] = (layer1_outputs[2372]) & ~(layer1_outputs[694]);
    assign layer2_outputs[381] = 1'b0;
    assign layer2_outputs[382] = ~(layer1_outputs[1208]);
    assign layer2_outputs[383] = ~((layer1_outputs[34]) & (layer1_outputs[1572]));
    assign layer2_outputs[384] = layer1_outputs[2173];
    assign layer2_outputs[385] = (layer1_outputs[2521]) & ~(layer1_outputs[635]);
    assign layer2_outputs[386] = ~(layer1_outputs[2007]) | (layer1_outputs[1294]);
    assign layer2_outputs[387] = ~(layer1_outputs[347]);
    assign layer2_outputs[388] = ~(layer1_outputs[1910]) | (layer1_outputs[869]);
    assign layer2_outputs[389] = (layer1_outputs[87]) & ~(layer1_outputs[188]);
    assign layer2_outputs[390] = (layer1_outputs[466]) & ~(layer1_outputs[416]);
    assign layer2_outputs[391] = ~(layer1_outputs[2242]) | (layer1_outputs[1523]);
    assign layer2_outputs[392] = ~(layer1_outputs[1544]) | (layer1_outputs[1332]);
    assign layer2_outputs[393] = (layer1_outputs[641]) & ~(layer1_outputs[2323]);
    assign layer2_outputs[394] = layer1_outputs[1901];
    assign layer2_outputs[395] = (layer1_outputs[1630]) & ~(layer1_outputs[2160]);
    assign layer2_outputs[396] = ~(layer1_outputs[2137]) | (layer1_outputs[1144]);
    assign layer2_outputs[397] = ~(layer1_outputs[2424]);
    assign layer2_outputs[398] = layer1_outputs[488];
    assign layer2_outputs[399] = (layer1_outputs[640]) & (layer1_outputs[2274]);
    assign layer2_outputs[400] = layer1_outputs[1255];
    assign layer2_outputs[401] = (layer1_outputs[1831]) & ~(layer1_outputs[1870]);
    assign layer2_outputs[402] = (layer1_outputs[478]) & ~(layer1_outputs[2183]);
    assign layer2_outputs[403] = ~(layer1_outputs[1575]);
    assign layer2_outputs[404] = layer1_outputs[1408];
    assign layer2_outputs[405] = ~((layer1_outputs[945]) & (layer1_outputs[1609]));
    assign layer2_outputs[406] = ~(layer1_outputs[696]);
    assign layer2_outputs[407] = ~(layer1_outputs[2183]) | (layer1_outputs[2253]);
    assign layer2_outputs[408] = ~(layer1_outputs[114]);
    assign layer2_outputs[409] = ~((layer1_outputs[599]) ^ (layer1_outputs[495]));
    assign layer2_outputs[410] = ~((layer1_outputs[2379]) & (layer1_outputs[566]));
    assign layer2_outputs[411] = ~(layer1_outputs[538]) | (layer1_outputs[1551]);
    assign layer2_outputs[412] = layer1_outputs[113];
    assign layer2_outputs[413] = layer1_outputs[1310];
    assign layer2_outputs[414] = (layer1_outputs[1113]) & ~(layer1_outputs[762]);
    assign layer2_outputs[415] = ~(layer1_outputs[180]) | (layer1_outputs[59]);
    assign layer2_outputs[416] = layer1_outputs[2068];
    assign layer2_outputs[417] = (layer1_outputs[592]) & (layer1_outputs[171]);
    assign layer2_outputs[418] = layer1_outputs[727];
    assign layer2_outputs[419] = layer1_outputs[879];
    assign layer2_outputs[420] = ~(layer1_outputs[852]) | (layer1_outputs[1384]);
    assign layer2_outputs[421] = (layer1_outputs[2198]) | (layer1_outputs[1004]);
    assign layer2_outputs[422] = layer1_outputs[1675];
    assign layer2_outputs[423] = ~(layer1_outputs[171]) | (layer1_outputs[1225]);
    assign layer2_outputs[424] = (layer1_outputs[1800]) & ~(layer1_outputs[943]);
    assign layer2_outputs[425] = ~((layer1_outputs[52]) & (layer1_outputs[224]));
    assign layer2_outputs[426] = (layer1_outputs[1267]) & ~(layer1_outputs[493]);
    assign layer2_outputs[427] = ~((layer1_outputs[1016]) & (layer1_outputs[1932]));
    assign layer2_outputs[428] = ~(layer1_outputs[1533]);
    assign layer2_outputs[429] = (layer1_outputs[2327]) & ~(layer1_outputs[1585]);
    assign layer2_outputs[430] = layer1_outputs[2200];
    assign layer2_outputs[431] = (layer1_outputs[1526]) & (layer1_outputs[2305]);
    assign layer2_outputs[432] = ~(layer1_outputs[40]);
    assign layer2_outputs[433] = (layer1_outputs[1344]) | (layer1_outputs[1555]);
    assign layer2_outputs[434] = (layer1_outputs[1224]) & (layer1_outputs[2434]);
    assign layer2_outputs[435] = layer1_outputs[1500];
    assign layer2_outputs[436] = layer1_outputs[13];
    assign layer2_outputs[437] = ~(layer1_outputs[1265]);
    assign layer2_outputs[438] = ~(layer1_outputs[1619]) | (layer1_outputs[1966]);
    assign layer2_outputs[439] = (layer1_outputs[487]) | (layer1_outputs[1116]);
    assign layer2_outputs[440] = layer1_outputs[1842];
    assign layer2_outputs[441] = layer1_outputs[1598];
    assign layer2_outputs[442] = ~(layer1_outputs[689]);
    assign layer2_outputs[443] = 1'b0;
    assign layer2_outputs[444] = layer1_outputs[580];
    assign layer2_outputs[445] = ~(layer1_outputs[1518]);
    assign layer2_outputs[446] = ~((layer1_outputs[167]) ^ (layer1_outputs[2336]));
    assign layer2_outputs[447] = (layer1_outputs[390]) & (layer1_outputs[2001]);
    assign layer2_outputs[448] = ~((layer1_outputs[280]) | (layer1_outputs[132]));
    assign layer2_outputs[449] = ~(layer1_outputs[1813]) | (layer1_outputs[2309]);
    assign layer2_outputs[450] = ~(layer1_outputs[1338]);
    assign layer2_outputs[451] = 1'b0;
    assign layer2_outputs[452] = ~(layer1_outputs[1882]);
    assign layer2_outputs[453] = (layer1_outputs[418]) & (layer1_outputs[172]);
    assign layer2_outputs[454] = ~(layer1_outputs[790]);
    assign layer2_outputs[455] = layer1_outputs[112];
    assign layer2_outputs[456] = ~(layer1_outputs[370]);
    assign layer2_outputs[457] = layer1_outputs[1625];
    assign layer2_outputs[458] = (layer1_outputs[616]) & ~(layer1_outputs[812]);
    assign layer2_outputs[459] = (layer1_outputs[987]) & (layer1_outputs[1693]);
    assign layer2_outputs[460] = ~(layer1_outputs[953]);
    assign layer2_outputs[461] = ~((layer1_outputs[595]) | (layer1_outputs[2404]));
    assign layer2_outputs[462] = ~((layer1_outputs[156]) & (layer1_outputs[810]));
    assign layer2_outputs[463] = ~(layer1_outputs[1746]) | (layer1_outputs[1741]);
    assign layer2_outputs[464] = (layer1_outputs[2133]) | (layer1_outputs[352]);
    assign layer2_outputs[465] = ~((layer1_outputs[1071]) & (layer1_outputs[288]));
    assign layer2_outputs[466] = (layer1_outputs[245]) & ~(layer1_outputs[1158]);
    assign layer2_outputs[467] = layer1_outputs[2103];
    assign layer2_outputs[468] = ~(layer1_outputs[1013]);
    assign layer2_outputs[469] = ~(layer1_outputs[1350]) | (layer1_outputs[1663]);
    assign layer2_outputs[470] = 1'b1;
    assign layer2_outputs[471] = 1'b1;
    assign layer2_outputs[472] = (layer1_outputs[1875]) ^ (layer1_outputs[346]);
    assign layer2_outputs[473] = ~(layer1_outputs[958]);
    assign layer2_outputs[474] = ~(layer1_outputs[903]);
    assign layer2_outputs[475] = ~(layer1_outputs[126]);
    assign layer2_outputs[476] = ~((layer1_outputs[95]) & (layer1_outputs[283]));
    assign layer2_outputs[477] = (layer1_outputs[824]) & ~(layer1_outputs[1694]);
    assign layer2_outputs[478] = ~((layer1_outputs[268]) | (layer1_outputs[2078]));
    assign layer2_outputs[479] = ~(layer1_outputs[1549]) | (layer1_outputs[766]);
    assign layer2_outputs[480] = (layer1_outputs[1152]) & (layer1_outputs[140]);
    assign layer2_outputs[481] = (layer1_outputs[1862]) & ~(layer1_outputs[1239]);
    assign layer2_outputs[482] = ~(layer1_outputs[1835]);
    assign layer2_outputs[483] = ~((layer1_outputs[568]) | (layer1_outputs[1635]));
    assign layer2_outputs[484] = layer1_outputs[1715];
    assign layer2_outputs[485] = ~(layer1_outputs[1137]);
    assign layer2_outputs[486] = ~(layer1_outputs[112]);
    assign layer2_outputs[487] = layer1_outputs[1118];
    assign layer2_outputs[488] = 1'b1;
    assign layer2_outputs[489] = (layer1_outputs[1459]) & ~(layer1_outputs[152]);
    assign layer2_outputs[490] = layer1_outputs[1330];
    assign layer2_outputs[491] = layer1_outputs[308];
    assign layer2_outputs[492] = (layer1_outputs[713]) | (layer1_outputs[1135]);
    assign layer2_outputs[493] = layer1_outputs[906];
    assign layer2_outputs[494] = ~(layer1_outputs[1295]) | (layer1_outputs[2168]);
    assign layer2_outputs[495] = ~(layer1_outputs[2128]);
    assign layer2_outputs[496] = ~(layer1_outputs[1651]);
    assign layer2_outputs[497] = 1'b0;
    assign layer2_outputs[498] = (layer1_outputs[455]) & (layer1_outputs[1341]);
    assign layer2_outputs[499] = ~(layer1_outputs[217]);
    assign layer2_outputs[500] = 1'b1;
    assign layer2_outputs[501] = (layer1_outputs[1925]) & ~(layer1_outputs[122]);
    assign layer2_outputs[502] = layer1_outputs[1372];
    assign layer2_outputs[503] = ~(layer1_outputs[223]) | (layer1_outputs[195]);
    assign layer2_outputs[504] = (layer1_outputs[348]) & (layer1_outputs[686]);
    assign layer2_outputs[505] = layer1_outputs[1172];
    assign layer2_outputs[506] = (layer1_outputs[204]) ^ (layer1_outputs[2393]);
    assign layer2_outputs[507] = ~((layer1_outputs[456]) ^ (layer1_outputs[777]));
    assign layer2_outputs[508] = 1'b1;
    assign layer2_outputs[509] = layer1_outputs[687];
    assign layer2_outputs[510] = 1'b1;
    assign layer2_outputs[511] = ~((layer1_outputs[1993]) | (layer1_outputs[776]));
    assign layer2_outputs[512] = (layer1_outputs[1928]) & (layer1_outputs[2081]);
    assign layer2_outputs[513] = ~(layer1_outputs[2406]) | (layer1_outputs[2094]);
    assign layer2_outputs[514] = ~(layer1_outputs[2249]);
    assign layer2_outputs[515] = ~(layer1_outputs[1210]);
    assign layer2_outputs[516] = ~(layer1_outputs[1795]);
    assign layer2_outputs[517] = (layer1_outputs[1740]) & ~(layer1_outputs[2558]);
    assign layer2_outputs[518] = ~((layer1_outputs[1294]) & (layer1_outputs[1513]));
    assign layer2_outputs[519] = layer1_outputs[1788];
    assign layer2_outputs[520] = (layer1_outputs[2199]) & ~(layer1_outputs[449]);
    assign layer2_outputs[521] = layer1_outputs[1355];
    assign layer2_outputs[522] = ~((layer1_outputs[1286]) | (layer1_outputs[2216]));
    assign layer2_outputs[523] = layer1_outputs[296];
    assign layer2_outputs[524] = layer1_outputs[791];
    assign layer2_outputs[525] = ~(layer1_outputs[330]) | (layer1_outputs[647]);
    assign layer2_outputs[526] = (layer1_outputs[2257]) & ~(layer1_outputs[1838]);
    assign layer2_outputs[527] = layer1_outputs[1851];
    assign layer2_outputs[528] = ~(layer1_outputs[1087]);
    assign layer2_outputs[529] = layer1_outputs[979];
    assign layer2_outputs[530] = ~(layer1_outputs[1791]);
    assign layer2_outputs[531] = (layer1_outputs[775]) & ~(layer1_outputs[2487]);
    assign layer2_outputs[532] = ~(layer1_outputs[1735]) | (layer1_outputs[611]);
    assign layer2_outputs[533] = ~(layer1_outputs[1090]);
    assign layer2_outputs[534] = 1'b0;
    assign layer2_outputs[535] = layer1_outputs[1818];
    assign layer2_outputs[536] = (layer1_outputs[1409]) & ~(layer1_outputs[501]);
    assign layer2_outputs[537] = ~(layer1_outputs[1115]);
    assign layer2_outputs[538] = (layer1_outputs[409]) | (layer1_outputs[448]);
    assign layer2_outputs[539] = layer1_outputs[1184];
    assign layer2_outputs[540] = 1'b0;
    assign layer2_outputs[541] = ~(layer1_outputs[1822]) | (layer1_outputs[105]);
    assign layer2_outputs[542] = ~(layer1_outputs[2484]);
    assign layer2_outputs[543] = ~((layer1_outputs[2168]) | (layer1_outputs[2517]));
    assign layer2_outputs[544] = layer1_outputs[221];
    assign layer2_outputs[545] = (layer1_outputs[2521]) & ~(layer1_outputs[841]);
    assign layer2_outputs[546] = (layer1_outputs[939]) & ~(layer1_outputs[163]);
    assign layer2_outputs[547] = (layer1_outputs[331]) ^ (layer1_outputs[1843]);
    assign layer2_outputs[548] = ~(layer1_outputs[634]);
    assign layer2_outputs[549] = ~(layer1_outputs[1685]) | (layer1_outputs[670]);
    assign layer2_outputs[550] = layer1_outputs[1971];
    assign layer2_outputs[551] = ~(layer1_outputs[1313]);
    assign layer2_outputs[552] = (layer1_outputs[1011]) ^ (layer1_outputs[1668]);
    assign layer2_outputs[553] = (layer1_outputs[1750]) & ~(layer1_outputs[1154]);
    assign layer2_outputs[554] = layer1_outputs[145];
    assign layer2_outputs[555] = ~((layer1_outputs[420]) | (layer1_outputs[2144]));
    assign layer2_outputs[556] = layer1_outputs[80];
    assign layer2_outputs[557] = layer1_outputs[2557];
    assign layer2_outputs[558] = (layer1_outputs[1407]) | (layer1_outputs[2290]);
    assign layer2_outputs[559] = layer1_outputs[380];
    assign layer2_outputs[560] = (layer1_outputs[652]) & ~(layer1_outputs[2432]);
    assign layer2_outputs[561] = ~(layer1_outputs[2551]) | (layer1_outputs[2430]);
    assign layer2_outputs[562] = 1'b1;
    assign layer2_outputs[563] = (layer1_outputs[158]) | (layer1_outputs[214]);
    assign layer2_outputs[564] = (layer1_outputs[2485]) | (layer1_outputs[1356]);
    assign layer2_outputs[565] = ~(layer1_outputs[350]);
    assign layer2_outputs[566] = ~(layer1_outputs[1027]);
    assign layer2_outputs[567] = layer1_outputs[593];
    assign layer2_outputs[568] = 1'b1;
    assign layer2_outputs[569] = layer1_outputs[1383];
    assign layer2_outputs[570] = (layer1_outputs[1627]) | (layer1_outputs[1984]);
    assign layer2_outputs[571] = (layer1_outputs[1521]) ^ (layer1_outputs[884]);
    assign layer2_outputs[572] = (layer1_outputs[1240]) & ~(layer1_outputs[839]);
    assign layer2_outputs[573] = layer1_outputs[235];
    assign layer2_outputs[574] = (layer1_outputs[554]) & ~(layer1_outputs[239]);
    assign layer2_outputs[575] = (layer1_outputs[103]) | (layer1_outputs[251]);
    assign layer2_outputs[576] = layer1_outputs[87];
    assign layer2_outputs[577] = ~(layer1_outputs[141]);
    assign layer2_outputs[578] = 1'b1;
    assign layer2_outputs[579] = ~(layer1_outputs[1917]) | (layer1_outputs[337]);
    assign layer2_outputs[580] = ~((layer1_outputs[541]) & (layer1_outputs[1697]));
    assign layer2_outputs[581] = ~(layer1_outputs[641]) | (layer1_outputs[645]);
    assign layer2_outputs[582] = ~(layer1_outputs[1757]);
    assign layer2_outputs[583] = ~(layer1_outputs[2279]);
    assign layer2_outputs[584] = (layer1_outputs[1819]) & ~(layer1_outputs[1992]);
    assign layer2_outputs[585] = ~(layer1_outputs[1960]);
    assign layer2_outputs[586] = ~(layer1_outputs[424]);
    assign layer2_outputs[587] = ~((layer1_outputs[1246]) & (layer1_outputs[1269]));
    assign layer2_outputs[588] = ~((layer1_outputs[1872]) & (layer1_outputs[387]));
    assign layer2_outputs[589] = ~(layer1_outputs[416]);
    assign layer2_outputs[590] = ~(layer1_outputs[1890]);
    assign layer2_outputs[591] = 1'b1;
    assign layer2_outputs[592] = (layer1_outputs[93]) & ~(layer1_outputs[768]);
    assign layer2_outputs[593] = ~(layer1_outputs[1673]);
    assign layer2_outputs[594] = (layer1_outputs[2014]) ^ (layer1_outputs[877]);
    assign layer2_outputs[595] = ~(layer1_outputs[99]) | (layer1_outputs[489]);
    assign layer2_outputs[596] = (layer1_outputs[1066]) & ~(layer1_outputs[194]);
    assign layer2_outputs[597] = layer1_outputs[777];
    assign layer2_outputs[598] = (layer1_outputs[2178]) & ~(layer1_outputs[2015]);
    assign layer2_outputs[599] = (layer1_outputs[2113]) & (layer1_outputs[111]);
    assign layer2_outputs[600] = layer1_outputs[451];
    assign layer2_outputs[601] = 1'b1;
    assign layer2_outputs[602] = 1'b1;
    assign layer2_outputs[603] = layer1_outputs[1489];
    assign layer2_outputs[604] = (layer1_outputs[1670]) | (layer1_outputs[470]);
    assign layer2_outputs[605] = ~((layer1_outputs[191]) | (layer1_outputs[1342]));
    assign layer2_outputs[606] = ~((layer1_outputs[793]) & (layer1_outputs[892]));
    assign layer2_outputs[607] = (layer1_outputs[251]) & (layer1_outputs[1536]);
    assign layer2_outputs[608] = ~(layer1_outputs[1639]);
    assign layer2_outputs[609] = (layer1_outputs[632]) | (layer1_outputs[1841]);
    assign layer2_outputs[610] = layer1_outputs[2483];
    assign layer2_outputs[611] = ~(layer1_outputs[1335]) | (layer1_outputs[2014]);
    assign layer2_outputs[612] = 1'b0;
    assign layer2_outputs[613] = ~(layer1_outputs[187]);
    assign layer2_outputs[614] = (layer1_outputs[1171]) & ~(layer1_outputs[1345]);
    assign layer2_outputs[615] = ~((layer1_outputs[1000]) & (layer1_outputs[1635]));
    assign layer2_outputs[616] = ~((layer1_outputs[2311]) & (layer1_outputs[12]));
    assign layer2_outputs[617] = ~(layer1_outputs[49]) | (layer1_outputs[1586]);
    assign layer2_outputs[618] = ~(layer1_outputs[1471]) | (layer1_outputs[472]);
    assign layer2_outputs[619] = (layer1_outputs[79]) & ~(layer1_outputs[1259]);
    assign layer2_outputs[620] = 1'b1;
    assign layer2_outputs[621] = ~(layer1_outputs[232]);
    assign layer2_outputs[622] = layer1_outputs[2357];
    assign layer2_outputs[623] = ~((layer1_outputs[1672]) & (layer1_outputs[492]));
    assign layer2_outputs[624] = ~((layer1_outputs[58]) | (layer1_outputs[111]));
    assign layer2_outputs[625] = 1'b1;
    assign layer2_outputs[626] = (layer1_outputs[1774]) & ~(layer1_outputs[2122]);
    assign layer2_outputs[627] = ~((layer1_outputs[2080]) & (layer1_outputs[1828]));
    assign layer2_outputs[628] = (layer1_outputs[1718]) & (layer1_outputs[1248]);
    assign layer2_outputs[629] = ~(layer1_outputs[1196]);
    assign layer2_outputs[630] = layer1_outputs[1745];
    assign layer2_outputs[631] = ~((layer1_outputs[802]) | (layer1_outputs[2510]));
    assign layer2_outputs[632] = ~(layer1_outputs[498]);
    assign layer2_outputs[633] = ~(layer1_outputs[1054]);
    assign layer2_outputs[634] = (layer1_outputs[1362]) & ~(layer1_outputs[1736]);
    assign layer2_outputs[635] = (layer1_outputs[37]) & ~(layer1_outputs[2120]);
    assign layer2_outputs[636] = (layer1_outputs[1957]) & (layer1_outputs[2446]);
    assign layer2_outputs[637] = ~(layer1_outputs[1047]) | (layer1_outputs[1715]);
    assign layer2_outputs[638] = (layer1_outputs[407]) & (layer1_outputs[254]);
    assign layer2_outputs[639] = layer1_outputs[2529];
    assign layer2_outputs[640] = ~((layer1_outputs[1461]) | (layer1_outputs[1810]));
    assign layer2_outputs[641] = ~(layer1_outputs[1711]) | (layer1_outputs[711]);
    assign layer2_outputs[642] = 1'b0;
    assign layer2_outputs[643] = ~(layer1_outputs[1974]) | (layer1_outputs[95]);
    assign layer2_outputs[644] = (layer1_outputs[763]) | (layer1_outputs[890]);
    assign layer2_outputs[645] = ~(layer1_outputs[1534]);
    assign layer2_outputs[646] = layer1_outputs[725];
    assign layer2_outputs[647] = ~(layer1_outputs[2258]);
    assign layer2_outputs[648] = layer1_outputs[1346];
    assign layer2_outputs[649] = ~((layer1_outputs[56]) & (layer1_outputs[967]));
    assign layer2_outputs[650] = ~(layer1_outputs[716]);
    assign layer2_outputs[651] = 1'b0;
    assign layer2_outputs[652] = (layer1_outputs[1316]) & ~(layer1_outputs[200]);
    assign layer2_outputs[653] = ~((layer1_outputs[1185]) | (layer1_outputs[2210]));
    assign layer2_outputs[654] = (layer1_outputs[266]) & ~(layer1_outputs[355]);
    assign layer2_outputs[655] = layer1_outputs[1340];
    assign layer2_outputs[656] = layer1_outputs[2440];
    assign layer2_outputs[657] = 1'b0;
    assign layer2_outputs[658] = ~(layer1_outputs[499]);
    assign layer2_outputs[659] = ~(layer1_outputs[969]);
    assign layer2_outputs[660] = ~(layer1_outputs[1046]);
    assign layer2_outputs[661] = ~((layer1_outputs[1802]) & (layer1_outputs[1139]));
    assign layer2_outputs[662] = (layer1_outputs[1333]) & ~(layer1_outputs[1510]);
    assign layer2_outputs[663] = ~(layer1_outputs[2204]) | (layer1_outputs[612]);
    assign layer2_outputs[664] = layer1_outputs[2052];
    assign layer2_outputs[665] = ~((layer1_outputs[639]) | (layer1_outputs[709]));
    assign layer2_outputs[666] = layer1_outputs[1011];
    assign layer2_outputs[667] = (layer1_outputs[729]) & ~(layer1_outputs[109]);
    assign layer2_outputs[668] = ~((layer1_outputs[1512]) ^ (layer1_outputs[689]));
    assign layer2_outputs[669] = layer1_outputs[1157];
    assign layer2_outputs[670] = (layer1_outputs[711]) & (layer1_outputs[2229]);
    assign layer2_outputs[671] = layer1_outputs[1588];
    assign layer2_outputs[672] = layer1_outputs[1090];
    assign layer2_outputs[673] = ~(layer1_outputs[619]);
    assign layer2_outputs[674] = ~(layer1_outputs[2142]);
    assign layer2_outputs[675] = ~((layer1_outputs[1591]) & (layer1_outputs[28]));
    assign layer2_outputs[676] = ~(layer1_outputs[2376]);
    assign layer2_outputs[677] = ~((layer1_outputs[755]) ^ (layer1_outputs[1351]));
    assign layer2_outputs[678] = ~(layer1_outputs[577]);
    assign layer2_outputs[679] = ~((layer1_outputs[1048]) & (layer1_outputs[2512]));
    assign layer2_outputs[680] = layer1_outputs[1580];
    assign layer2_outputs[681] = 1'b1;
    assign layer2_outputs[682] = ~(layer1_outputs[983]);
    assign layer2_outputs[683] = ~((layer1_outputs[1130]) & (layer1_outputs[530]));
    assign layer2_outputs[684] = (layer1_outputs[1559]) & ~(layer1_outputs[993]);
    assign layer2_outputs[685] = ~(layer1_outputs[269]);
    assign layer2_outputs[686] = ~((layer1_outputs[1673]) | (layer1_outputs[545]));
    assign layer2_outputs[687] = layer1_outputs[1202];
    assign layer2_outputs[688] = layer1_outputs[873];
    assign layer2_outputs[689] = ~(layer1_outputs[1354]);
    assign layer2_outputs[690] = (layer1_outputs[1150]) ^ (layer1_outputs[441]);
    assign layer2_outputs[691] = (layer1_outputs[657]) | (layer1_outputs[572]);
    assign layer2_outputs[692] = 1'b0;
    assign layer2_outputs[693] = ~(layer1_outputs[1274]);
    assign layer2_outputs[694] = layer1_outputs[1416];
    assign layer2_outputs[695] = ~((layer1_outputs[136]) | (layer1_outputs[436]));
    assign layer2_outputs[696] = (layer1_outputs[1584]) & ~(layer1_outputs[1928]);
    assign layer2_outputs[697] = layer1_outputs[1899];
    assign layer2_outputs[698] = (layer1_outputs[1305]) | (layer1_outputs[256]);
    assign layer2_outputs[699] = (layer1_outputs[1298]) | (layer1_outputs[2250]);
    assign layer2_outputs[700] = layer1_outputs[730];
    assign layer2_outputs[701] = ~(layer1_outputs[2071]);
    assign layer2_outputs[702] = layer1_outputs[997];
    assign layer2_outputs[703] = ~(layer1_outputs[2358]) | (layer1_outputs[292]);
    assign layer2_outputs[704] = ~(layer1_outputs[76]) | (layer1_outputs[568]);
    assign layer2_outputs[705] = (layer1_outputs[810]) | (layer1_outputs[1878]);
    assign layer2_outputs[706] = ~((layer1_outputs[1801]) & (layer1_outputs[1711]));
    assign layer2_outputs[707] = ~((layer1_outputs[2319]) | (layer1_outputs[2290]));
    assign layer2_outputs[708] = 1'b1;
    assign layer2_outputs[709] = (layer1_outputs[429]) & ~(layer1_outputs[582]);
    assign layer2_outputs[710] = ~((layer1_outputs[714]) | (layer1_outputs[1985]));
    assign layer2_outputs[711] = (layer1_outputs[509]) & ~(layer1_outputs[78]);
    assign layer2_outputs[712] = layer1_outputs[910];
    assign layer2_outputs[713] = layer1_outputs[1965];
    assign layer2_outputs[714] = ~(layer1_outputs[2256]) | (layer1_outputs[458]);
    assign layer2_outputs[715] = (layer1_outputs[1953]) & ~(layer1_outputs[1268]);
    assign layer2_outputs[716] = (layer1_outputs[379]) & ~(layer1_outputs[994]);
    assign layer2_outputs[717] = (layer1_outputs[767]) & ~(layer1_outputs[1362]);
    assign layer2_outputs[718] = ~(layer1_outputs[993]);
    assign layer2_outputs[719] = 1'b0;
    assign layer2_outputs[720] = (layer1_outputs[1514]) & (layer1_outputs[2132]);
    assign layer2_outputs[721] = ~((layer1_outputs[867]) | (layer1_outputs[872]));
    assign layer2_outputs[722] = ~((layer1_outputs[1809]) ^ (layer1_outputs[614]));
    assign layer2_outputs[723] = ~(layer1_outputs[1435]);
    assign layer2_outputs[724] = (layer1_outputs[1307]) & (layer1_outputs[128]);
    assign layer2_outputs[725] = ~(layer1_outputs[2104]);
    assign layer2_outputs[726] = ~(layer1_outputs[864]) | (layer1_outputs[1484]);
    assign layer2_outputs[727] = ~(layer1_outputs[213]) | (layer1_outputs[1884]);
    assign layer2_outputs[728] = ~((layer1_outputs[1100]) & (layer1_outputs[1963]));
    assign layer2_outputs[729] = ~(layer1_outputs[2338]) | (layer1_outputs[478]);
    assign layer2_outputs[730] = layer1_outputs[1571];
    assign layer2_outputs[731] = ~(layer1_outputs[200]);
    assign layer2_outputs[732] = layer1_outputs[1484];
    assign layer2_outputs[733] = (layer1_outputs[1129]) | (layer1_outputs[1897]);
    assign layer2_outputs[734] = 1'b0;
    assign layer2_outputs[735] = (layer1_outputs[243]) & ~(layer1_outputs[386]);
    assign layer2_outputs[736] = ~(layer1_outputs[1866]);
    assign layer2_outputs[737] = layer1_outputs[1961];
    assign layer2_outputs[738] = ~(layer1_outputs[801]);
    assign layer2_outputs[739] = (layer1_outputs[1751]) & (layer1_outputs[1672]);
    assign layer2_outputs[740] = ~(layer1_outputs[2188]);
    assign layer2_outputs[741] = (layer1_outputs[52]) & ~(layer1_outputs[571]);
    assign layer2_outputs[742] = (layer1_outputs[1174]) & ~(layer1_outputs[2301]);
    assign layer2_outputs[743] = (layer1_outputs[19]) ^ (layer1_outputs[459]);
    assign layer2_outputs[744] = layer1_outputs[524];
    assign layer2_outputs[745] = ~((layer1_outputs[888]) | (layer1_outputs[1754]));
    assign layer2_outputs[746] = ~(layer1_outputs[475]);
    assign layer2_outputs[747] = ~(layer1_outputs[2407]);
    assign layer2_outputs[748] = layer1_outputs[2065];
    assign layer2_outputs[749] = ~((layer1_outputs[1844]) & (layer1_outputs[757]));
    assign layer2_outputs[750] = (layer1_outputs[1093]) & (layer1_outputs[1940]);
    assign layer2_outputs[751] = (layer1_outputs[1848]) & ~(layer1_outputs[1699]);
    assign layer2_outputs[752] = ~((layer1_outputs[1911]) | (layer1_outputs[2341]));
    assign layer2_outputs[753] = (layer1_outputs[434]) & (layer1_outputs[691]);
    assign layer2_outputs[754] = (layer1_outputs[1405]) | (layer1_outputs[365]);
    assign layer2_outputs[755] = ~(layer1_outputs[14]);
    assign layer2_outputs[756] = ~((layer1_outputs[626]) | (layer1_outputs[1748]));
    assign layer2_outputs[757] = layer1_outputs[1599];
    assign layer2_outputs[758] = (layer1_outputs[1879]) | (layer1_outputs[1368]);
    assign layer2_outputs[759] = ~(layer1_outputs[1376]) | (layer1_outputs[1229]);
    assign layer2_outputs[760] = ~(layer1_outputs[618]) | (layer1_outputs[981]);
    assign layer2_outputs[761] = layer1_outputs[630];
    assign layer2_outputs[762] = 1'b0;
    assign layer2_outputs[763] = ~((layer1_outputs[396]) & (layer1_outputs[60]));
    assign layer2_outputs[764] = ~(layer1_outputs[2302]);
    assign layer2_outputs[765] = layer1_outputs[1123];
    assign layer2_outputs[766] = layer1_outputs[1697];
    assign layer2_outputs[767] = ~(layer1_outputs[2331]);
    assign layer2_outputs[768] = (layer1_outputs[1385]) | (layer1_outputs[124]);
    assign layer2_outputs[769] = ~(layer1_outputs[878]) | (layer1_outputs[2433]);
    assign layer2_outputs[770] = layer1_outputs[1169];
    assign layer2_outputs[771] = layer1_outputs[2224];
    assign layer2_outputs[772] = ~(layer1_outputs[65]);
    assign layer2_outputs[773] = (layer1_outputs[656]) | (layer1_outputs[1055]);
    assign layer2_outputs[774] = (layer1_outputs[1515]) & ~(layer1_outputs[1364]);
    assign layer2_outputs[775] = (layer1_outputs[756]) ^ (layer1_outputs[137]);
    assign layer2_outputs[776] = (layer1_outputs[1195]) ^ (layer1_outputs[1151]);
    assign layer2_outputs[777] = ~(layer1_outputs[2374]) | (layer1_outputs[1328]);
    assign layer2_outputs[778] = ~((layer1_outputs[1226]) | (layer1_outputs[657]));
    assign layer2_outputs[779] = layer1_outputs[290];
    assign layer2_outputs[780] = (layer1_outputs[1819]) & ~(layer1_outputs[1737]);
    assign layer2_outputs[781] = (layer1_outputs[1710]) & ~(layer1_outputs[2038]);
    assign layer2_outputs[782] = (layer1_outputs[2277]) & ~(layer1_outputs[25]);
    assign layer2_outputs[783] = layer1_outputs[426];
    assign layer2_outputs[784] = layer1_outputs[1291];
    assign layer2_outputs[785] = ~((layer1_outputs[389]) | (layer1_outputs[1892]));
    assign layer2_outputs[786] = (layer1_outputs[2244]) & ~(layer1_outputs[708]);
    assign layer2_outputs[787] = ~(layer1_outputs[2113]);
    assign layer2_outputs[788] = layer1_outputs[1598];
    assign layer2_outputs[789] = ~(layer1_outputs[1311]);
    assign layer2_outputs[790] = layer1_outputs[1107];
    assign layer2_outputs[791] = ~(layer1_outputs[1432]);
    assign layer2_outputs[792] = ~(layer1_outputs[742]);
    assign layer2_outputs[793] = layer1_outputs[1370];
    assign layer2_outputs[794] = layer1_outputs[929];
    assign layer2_outputs[795] = (layer1_outputs[1429]) & ~(layer1_outputs[2556]);
    assign layer2_outputs[796] = ~((layer1_outputs[258]) & (layer1_outputs[2015]));
    assign layer2_outputs[797] = ~(layer1_outputs[606]) | (layer1_outputs[2074]);
    assign layer2_outputs[798] = layer1_outputs[2096];
    assign layer2_outputs[799] = ~(layer1_outputs[1188]);
    assign layer2_outputs[800] = ~(layer1_outputs[634]);
    assign layer2_outputs[801] = ~(layer1_outputs[792]);
    assign layer2_outputs[802] = (layer1_outputs[915]) ^ (layer1_outputs[2503]);
    assign layer2_outputs[803] = (layer1_outputs[860]) ^ (layer1_outputs[781]);
    assign layer2_outputs[804] = ~(layer1_outputs[828]);
    assign layer2_outputs[805] = ~(layer1_outputs[1267]);
    assign layer2_outputs[806] = (layer1_outputs[801]) & ~(layer1_outputs[1304]);
    assign layer2_outputs[807] = (layer1_outputs[662]) & ~(layer1_outputs[2531]);
    assign layer2_outputs[808] = ~(layer1_outputs[2195]);
    assign layer2_outputs[809] = ~(layer1_outputs[1204]) | (layer1_outputs[441]);
    assign layer2_outputs[810] = layer1_outputs[1746];
    assign layer2_outputs[811] = layer1_outputs[208];
    assign layer2_outputs[812] = (layer1_outputs[2490]) & ~(layer1_outputs[593]);
    assign layer2_outputs[813] = (layer1_outputs[401]) | (layer1_outputs[1607]);
    assign layer2_outputs[814] = (layer1_outputs[430]) | (layer1_outputs[788]);
    assign layer2_outputs[815] = ~((layer1_outputs[1068]) ^ (layer1_outputs[1898]));
    assign layer2_outputs[816] = (layer1_outputs[2518]) | (layer1_outputs[785]);
    assign layer2_outputs[817] = (layer1_outputs[2163]) ^ (layer1_outputs[2088]);
    assign layer2_outputs[818] = (layer1_outputs[1319]) & ~(layer1_outputs[173]);
    assign layer2_outputs[819] = layer1_outputs[1085];
    assign layer2_outputs[820] = 1'b0;
    assign layer2_outputs[821] = 1'b1;
    assign layer2_outputs[822] = layer1_outputs[354];
    assign layer2_outputs[823] = ~(layer1_outputs[177]) | (layer1_outputs[49]);
    assign layer2_outputs[824] = ~(layer1_outputs[1482]) | (layer1_outputs[1280]);
    assign layer2_outputs[825] = ~(layer1_outputs[1253]) | (layer1_outputs[720]);
    assign layer2_outputs[826] = ~(layer1_outputs[669]);
    assign layer2_outputs[827] = ~((layer1_outputs[2190]) & (layer1_outputs[2064]));
    assign layer2_outputs[828] = ~(layer1_outputs[2451]);
    assign layer2_outputs[829] = (layer1_outputs[378]) & ~(layer1_outputs[228]);
    assign layer2_outputs[830] = (layer1_outputs[1826]) | (layer1_outputs[805]);
    assign layer2_outputs[831] = ~(layer1_outputs[927]) | (layer1_outputs[2111]);
    assign layer2_outputs[832] = ~((layer1_outputs[804]) & (layer1_outputs[391]));
    assign layer2_outputs[833] = ~(layer1_outputs[1351]);
    assign layer2_outputs[834] = ~(layer1_outputs[2249]) | (layer1_outputs[2005]);
    assign layer2_outputs[835] = ~(layer1_outputs[1344]);
    assign layer2_outputs[836] = (layer1_outputs[2512]) & ~(layer1_outputs[2203]);
    assign layer2_outputs[837] = layer1_outputs[425];
    assign layer2_outputs[838] = layer1_outputs[2488];
    assign layer2_outputs[839] = layer1_outputs[2197];
    assign layer2_outputs[840] = (layer1_outputs[928]) & ~(layer1_outputs[2344]);
    assign layer2_outputs[841] = ~((layer1_outputs[1571]) | (layer1_outputs[2022]));
    assign layer2_outputs[842] = ~((layer1_outputs[2094]) & (layer1_outputs[1381]));
    assign layer2_outputs[843] = 1'b1;
    assign layer2_outputs[844] = (layer1_outputs[335]) & ~(layer1_outputs[2400]);
    assign layer2_outputs[845] = ~(layer1_outputs[933]);
    assign layer2_outputs[846] = (layer1_outputs[721]) & ~(layer1_outputs[666]);
    assign layer2_outputs[847] = layer1_outputs[688];
    assign layer2_outputs[848] = 1'b1;
    assign layer2_outputs[849] = (layer1_outputs[1642]) & (layer1_outputs[537]);
    assign layer2_outputs[850] = ~(layer1_outputs[1667]) | (layer1_outputs[2330]);
    assign layer2_outputs[851] = layer1_outputs[2081];
    assign layer2_outputs[852] = ~(layer1_outputs[1917]) | (layer1_outputs[1007]);
    assign layer2_outputs[853] = ~(layer1_outputs[1244]);
    assign layer2_outputs[854] = layer1_outputs[527];
    assign layer2_outputs[855] = ~(layer1_outputs[582]);
    assign layer2_outputs[856] = ~(layer1_outputs[1682]) | (layer1_outputs[353]);
    assign layer2_outputs[857] = layer1_outputs[1821];
    assign layer2_outputs[858] = ~(layer1_outputs[2049]) | (layer1_outputs[1853]);
    assign layer2_outputs[859] = layer1_outputs[961];
    assign layer2_outputs[860] = layer1_outputs[2498];
    assign layer2_outputs[861] = ~(layer1_outputs[2449]);
    assign layer2_outputs[862] = (layer1_outputs[1149]) ^ (layer1_outputs[1910]);
    assign layer2_outputs[863] = layer1_outputs[2025];
    assign layer2_outputs[864] = (layer1_outputs[1441]) ^ (layer1_outputs[1158]);
    assign layer2_outputs[865] = 1'b0;
    assign layer2_outputs[866] = layer1_outputs[15];
    assign layer2_outputs[867] = 1'b1;
    assign layer2_outputs[868] = ~(layer1_outputs[114]);
    assign layer2_outputs[869] = layer1_outputs[905];
    assign layer2_outputs[870] = ~((layer1_outputs[255]) | (layer1_outputs[480]));
    assign layer2_outputs[871] = ~((layer1_outputs[287]) | (layer1_outputs[414]));
    assign layer2_outputs[872] = ~(layer1_outputs[667]);
    assign layer2_outputs[873] = layer1_outputs[958];
    assign layer2_outputs[874] = ~(layer1_outputs[512]) | (layer1_outputs[729]);
    assign layer2_outputs[875] = ~(layer1_outputs[438]);
    assign layer2_outputs[876] = ~(layer1_outputs[1326]);
    assign layer2_outputs[877] = ~(layer1_outputs[345]);
    assign layer2_outputs[878] = layer1_outputs[573];
    assign layer2_outputs[879] = 1'b0;
    assign layer2_outputs[880] = ~((layer1_outputs[2556]) ^ (layer1_outputs[1775]));
    assign layer2_outputs[881] = ~(layer1_outputs[1150]) | (layer1_outputs[1812]);
    assign layer2_outputs[882] = ~(layer1_outputs[804]) | (layer1_outputs[1038]);
    assign layer2_outputs[883] = 1'b0;
    assign layer2_outputs[884] = ~(layer1_outputs[2239]) | (layer1_outputs[174]);
    assign layer2_outputs[885] = (layer1_outputs[84]) | (layer1_outputs[2189]);
    assign layer2_outputs[886] = ~((layer1_outputs[1093]) | (layer1_outputs[2016]));
    assign layer2_outputs[887] = ~(layer1_outputs[1891]) | (layer1_outputs[1325]);
    assign layer2_outputs[888] = (layer1_outputs[26]) & ~(layer1_outputs[981]);
    assign layer2_outputs[889] = ~(layer1_outputs[1757]);
    assign layer2_outputs[890] = ~(layer1_outputs[2200]);
    assign layer2_outputs[891] = ~((layer1_outputs[1047]) | (layer1_outputs[1610]));
    assign layer2_outputs[892] = ~((layer1_outputs[272]) & (layer1_outputs[2437]));
    assign layer2_outputs[893] = (layer1_outputs[297]) & (layer1_outputs[1324]);
    assign layer2_outputs[894] = ~(layer1_outputs[947]);
    assign layer2_outputs[895] = ~(layer1_outputs[1498]) | (layer1_outputs[1676]);
    assign layer2_outputs[896] = ~(layer1_outputs[2123]) | (layer1_outputs[2405]);
    assign layer2_outputs[897] = (layer1_outputs[1654]) & ~(layer1_outputs[2355]);
    assign layer2_outputs[898] = ~(layer1_outputs[390]);
    assign layer2_outputs[899] = (layer1_outputs[1493]) & (layer1_outputs[1401]);
    assign layer2_outputs[900] = ~(layer1_outputs[2402]);
    assign layer2_outputs[901] = (layer1_outputs[1899]) & ~(layer1_outputs[1904]);
    assign layer2_outputs[902] = (layer1_outputs[2024]) | (layer1_outputs[997]);
    assign layer2_outputs[903] = (layer1_outputs[1612]) & (layer1_outputs[1816]);
    assign layer2_outputs[904] = ~((layer1_outputs[838]) & (layer1_outputs[1739]));
    assign layer2_outputs[905] = (layer1_outputs[2085]) & ~(layer1_outputs[300]);
    assign layer2_outputs[906] = ~(layer1_outputs[1219]);
    assign layer2_outputs[907] = ~(layer1_outputs[1222]);
    assign layer2_outputs[908] = (layer1_outputs[1040]) & ~(layer1_outputs[412]);
    assign layer2_outputs[909] = (layer1_outputs[2415]) & (layer1_outputs[2501]);
    assign layer2_outputs[910] = ~(layer1_outputs[1070]);
    assign layer2_outputs[911] = ~(layer1_outputs[741]);
    assign layer2_outputs[912] = (layer1_outputs[1832]) | (layer1_outputs[189]);
    assign layer2_outputs[913] = ~(layer1_outputs[860]) | (layer1_outputs[1329]);
    assign layer2_outputs[914] = ~(layer1_outputs[1231]);
    assign layer2_outputs[915] = ~(layer1_outputs[1543]) | (layer1_outputs[2269]);
    assign layer2_outputs[916] = ~((layer1_outputs[1998]) ^ (layer1_outputs[2505]));
    assign layer2_outputs[917] = (layer1_outputs[1933]) & ~(layer1_outputs[2109]);
    assign layer2_outputs[918] = (layer1_outputs[1045]) | (layer1_outputs[1791]);
    assign layer2_outputs[919] = ~((layer1_outputs[1288]) | (layer1_outputs[115]));
    assign layer2_outputs[920] = layer1_outputs[2523];
    assign layer2_outputs[921] = ~(layer1_outputs[2235]) | (layer1_outputs[1261]);
    assign layer2_outputs[922] = ~((layer1_outputs[538]) & (layer1_outputs[1804]));
    assign layer2_outputs[923] = (layer1_outputs[1681]) & (layer1_outputs[123]);
    assign layer2_outputs[924] = ~(layer1_outputs[2232]);
    assign layer2_outputs[925] = ~((layer1_outputs[2018]) & (layer1_outputs[1631]));
    assign layer2_outputs[926] = ~(layer1_outputs[661]) | (layer1_outputs[1683]);
    assign layer2_outputs[927] = (layer1_outputs[159]) & (layer1_outputs[1179]);
    assign layer2_outputs[928] = ~(layer1_outputs[1039]);
    assign layer2_outputs[929] = layer1_outputs[731];
    assign layer2_outputs[930] = 1'b0;
    assign layer2_outputs[931] = ~(layer1_outputs[654]);
    assign layer2_outputs[932] = ~((layer1_outputs[2059]) ^ (layer1_outputs[1099]));
    assign layer2_outputs[933] = ~(layer1_outputs[559]);
    assign layer2_outputs[934] = layer1_outputs[22];
    assign layer2_outputs[935] = (layer1_outputs[1709]) & ~(layer1_outputs[20]);
    assign layer2_outputs[936] = ~(layer1_outputs[247]);
    assign layer2_outputs[937] = layer1_outputs[2323];
    assign layer2_outputs[938] = 1'b0;
    assign layer2_outputs[939] = ~(layer1_outputs[1979]);
    assign layer2_outputs[940] = layer1_outputs[1744];
    assign layer2_outputs[941] = 1'b1;
    assign layer2_outputs[942] = layer1_outputs[340];
    assign layer2_outputs[943] = ~(layer1_outputs[2101]);
    assign layer2_outputs[944] = layer1_outputs[1220];
    assign layer2_outputs[945] = ~((layer1_outputs[222]) & (layer1_outputs[2438]));
    assign layer2_outputs[946] = ~(layer1_outputs[377]);
    assign layer2_outputs[947] = ~(layer1_outputs[2029]);
    assign layer2_outputs[948] = layer1_outputs[907];
    assign layer2_outputs[949] = (layer1_outputs[863]) & ~(layer1_outputs[614]);
    assign layer2_outputs[950] = ~(layer1_outputs[2261]) | (layer1_outputs[250]);
    assign layer2_outputs[951] = ~(layer1_outputs[1554]);
    assign layer2_outputs[952] = (layer1_outputs[2515]) & (layer1_outputs[1956]);
    assign layer2_outputs[953] = ~(layer1_outputs[2412]) | (layer1_outputs[631]);
    assign layer2_outputs[954] = ~(layer1_outputs[1140]);
    assign layer2_outputs[955] = ~((layer1_outputs[119]) & (layer1_outputs[1257]));
    assign layer2_outputs[956] = layer1_outputs[1134];
    assign layer2_outputs[957] = (layer1_outputs[482]) | (layer1_outputs[160]);
    assign layer2_outputs[958] = (layer1_outputs[1606]) & ~(layer1_outputs[2192]);
    assign layer2_outputs[959] = ~((layer1_outputs[2106]) | (layer1_outputs[548]));
    assign layer2_outputs[960] = layer1_outputs[1931];
    assign layer2_outputs[961] = ~(layer1_outputs[2066]);
    assign layer2_outputs[962] = ~(layer1_outputs[1649]);
    assign layer2_outputs[963] = (layer1_outputs[2265]) & ~(layer1_outputs[2360]);
    assign layer2_outputs[964] = ~(layer1_outputs[1912]);
    assign layer2_outputs[965] = (layer1_outputs[16]) ^ (layer1_outputs[642]);
    assign layer2_outputs[966] = layer1_outputs[1444];
    assign layer2_outputs[967] = ~((layer1_outputs[48]) | (layer1_outputs[1043]));
    assign layer2_outputs[968] = (layer1_outputs[845]) & (layer1_outputs[2439]);
    assign layer2_outputs[969] = 1'b0;
    assign layer2_outputs[970] = (layer1_outputs[88]) & ~(layer1_outputs[71]);
    assign layer2_outputs[971] = (layer1_outputs[2211]) & ~(layer1_outputs[769]);
    assign layer2_outputs[972] = ~((layer1_outputs[466]) & (layer1_outputs[931]));
    assign layer2_outputs[973] = 1'b1;
    assign layer2_outputs[974] = 1'b0;
    assign layer2_outputs[975] = ~(layer1_outputs[133]);
    assign layer2_outputs[976] = ~(layer1_outputs[1638]) | (layer1_outputs[1533]);
    assign layer2_outputs[977] = ~(layer1_outputs[1912]);
    assign layer2_outputs[978] = ~(layer1_outputs[615]);
    assign layer2_outputs[979] = (layer1_outputs[401]) & (layer1_outputs[587]);
    assign layer2_outputs[980] = ~(layer1_outputs[1065]) | (layer1_outputs[992]);
    assign layer2_outputs[981] = (layer1_outputs[754]) | (layer1_outputs[574]);
    assign layer2_outputs[982] = layer1_outputs[185];
    assign layer2_outputs[983] = ~(layer1_outputs[1639]);
    assign layer2_outputs[984] = ~((layer1_outputs[1798]) | (layer1_outputs[2431]));
    assign layer2_outputs[985] = layer1_outputs[2262];
    assign layer2_outputs[986] = ~(layer1_outputs[703]);
    assign layer2_outputs[987] = (layer1_outputs[2557]) | (layer1_outputs[1908]);
    assign layer2_outputs[988] = ~(layer1_outputs[264]);
    assign layer2_outputs[989] = 1'b0;
    assign layer2_outputs[990] = ~(layer1_outputs[748]);
    assign layer2_outputs[991] = ~(layer1_outputs[1538]) | (layer1_outputs[394]);
    assign layer2_outputs[992] = (layer1_outputs[1199]) & (layer1_outputs[2519]);
    assign layer2_outputs[993] = ~(layer1_outputs[1847]);
    assign layer2_outputs[994] = ~(layer1_outputs[2367]) | (layer1_outputs[1463]);
    assign layer2_outputs[995] = layer1_outputs[2223];
    assign layer2_outputs[996] = layer1_outputs[1942];
    assign layer2_outputs[997] = layer1_outputs[794];
    assign layer2_outputs[998] = ~((layer1_outputs[2270]) & (layer1_outputs[1689]));
    assign layer2_outputs[999] = ~((layer1_outputs[1973]) & (layer1_outputs[2472]));
    assign layer2_outputs[1000] = ~(layer1_outputs[2236]) | (layer1_outputs[1383]);
    assign layer2_outputs[1001] = (layer1_outputs[2498]) ^ (layer1_outputs[1873]);
    assign layer2_outputs[1002] = ~((layer1_outputs[2147]) ^ (layer1_outputs[1610]));
    assign layer2_outputs[1003] = ~(layer1_outputs[706]) | (layer1_outputs[552]);
    assign layer2_outputs[1004] = ~((layer1_outputs[2046]) | (layer1_outputs[162]));
    assign layer2_outputs[1005] = layer1_outputs[785];
    assign layer2_outputs[1006] = ~(layer1_outputs[1249]);
    assign layer2_outputs[1007] = ~((layer1_outputs[2225]) | (layer1_outputs[1363]));
    assign layer2_outputs[1008] = (layer1_outputs[1823]) | (layer1_outputs[285]);
    assign layer2_outputs[1009] = 1'b0;
    assign layer2_outputs[1010] = (layer1_outputs[129]) | (layer1_outputs[598]);
    assign layer2_outputs[1011] = (layer1_outputs[1732]) & ~(layer1_outputs[1849]);
    assign layer2_outputs[1012] = ~(layer1_outputs[1379]) | (layer1_outputs[440]);
    assign layer2_outputs[1013] = ~((layer1_outputs[783]) | (layer1_outputs[755]));
    assign layer2_outputs[1014] = layer1_outputs[152];
    assign layer2_outputs[1015] = ~(layer1_outputs[1187]) | (layer1_outputs[2334]);
    assign layer2_outputs[1016] = ~((layer1_outputs[1175]) | (layer1_outputs[1986]));
    assign layer2_outputs[1017] = ~((layer1_outputs[1223]) & (layer1_outputs[602]));
    assign layer2_outputs[1018] = (layer1_outputs[2003]) & ~(layer1_outputs[679]);
    assign layer2_outputs[1019] = ~(layer1_outputs[57]);
    assign layer2_outputs[1020] = layer1_outputs[436];
    assign layer2_outputs[1021] = layer1_outputs[1319];
    assign layer2_outputs[1022] = (layer1_outputs[1954]) & (layer1_outputs[224]);
    assign layer2_outputs[1023] = ~((layer1_outputs[787]) & (layer1_outputs[1173]));
    assign layer2_outputs[1024] = layer1_outputs[654];
    assign layer2_outputs[1025] = (layer1_outputs[2428]) & ~(layer1_outputs[2395]);
    assign layer2_outputs[1026] = ~(layer1_outputs[2291]);
    assign layer2_outputs[1027] = (layer1_outputs[438]) & (layer1_outputs[2354]);
    assign layer2_outputs[1028] = (layer1_outputs[75]) & (layer1_outputs[1573]);
    assign layer2_outputs[1029] = layer1_outputs[286];
    assign layer2_outputs[1030] = ~(layer1_outputs[192]);
    assign layer2_outputs[1031] = ~(layer1_outputs[1831]);
    assign layer2_outputs[1032] = ~(layer1_outputs[1825]) | (layer1_outputs[564]);
    assign layer2_outputs[1033] = layer1_outputs[497];
    assign layer2_outputs[1034] = layer1_outputs[1183];
    assign layer2_outputs[1035] = 1'b0;
    assign layer2_outputs[1036] = ~(layer1_outputs[895]) | (layer1_outputs[519]);
    assign layer2_outputs[1037] = ~(layer1_outputs[2096]) | (layer1_outputs[507]);
    assign layer2_outputs[1038] = 1'b0;
    assign layer2_outputs[1039] = ~(layer1_outputs[820]);
    assign layer2_outputs[1040] = (layer1_outputs[402]) & ~(layer1_outputs[1094]);
    assign layer2_outputs[1041] = ~(layer1_outputs[1031]) | (layer1_outputs[1969]);
    assign layer2_outputs[1042] = 1'b0;
    assign layer2_outputs[1043] = (layer1_outputs[563]) | (layer1_outputs[2416]);
    assign layer2_outputs[1044] = 1'b1;
    assign layer2_outputs[1045] = (layer1_outputs[995]) & (layer1_outputs[2322]);
    assign layer2_outputs[1046] = (layer1_outputs[2219]) & ~(layer1_outputs[381]);
    assign layer2_outputs[1047] = ~((layer1_outputs[2175]) | (layer1_outputs[1496]));
    assign layer2_outputs[1048] = ~(layer1_outputs[1045]);
    assign layer2_outputs[1049] = ~((layer1_outputs[1061]) ^ (layer1_outputs[1032]));
    assign layer2_outputs[1050] = layer1_outputs[491];
    assign layer2_outputs[1051] = (layer1_outputs[517]) & (layer1_outputs[2031]);
    assign layer2_outputs[1052] = layer1_outputs[731];
    assign layer2_outputs[1053] = 1'b0;
    assign layer2_outputs[1054] = 1'b0;
    assign layer2_outputs[1055] = ~((layer1_outputs[2287]) & (layer1_outputs[1919]));
    assign layer2_outputs[1056] = ~(layer1_outputs[1041]) | (layer1_outputs[2237]);
    assign layer2_outputs[1057] = (layer1_outputs[2019]) | (layer1_outputs[426]);
    assign layer2_outputs[1058] = ~((layer1_outputs[1519]) & (layer1_outputs[2036]));
    assign layer2_outputs[1059] = (layer1_outputs[1764]) ^ (layer1_outputs[228]);
    assign layer2_outputs[1060] = (layer1_outputs[3]) | (layer1_outputs[2413]);
    assign layer2_outputs[1061] = ~(layer1_outputs[722]) | (layer1_outputs[897]);
    assign layer2_outputs[1062] = ~(layer1_outputs[2194]) | (layer1_outputs[644]);
    assign layer2_outputs[1063] = (layer1_outputs[502]) | (layer1_outputs[66]);
    assign layer2_outputs[1064] = (layer1_outputs[1907]) & ~(layer1_outputs[1148]);
    assign layer2_outputs[1065] = layer1_outputs[2443];
    assign layer2_outputs[1066] = (layer1_outputs[1083]) | (layer1_outputs[1934]);
    assign layer2_outputs[1067] = (layer1_outputs[1126]) & ~(layer1_outputs[2033]);
    assign layer2_outputs[1068] = ~(layer1_outputs[832]);
    assign layer2_outputs[1069] = ~(layer1_outputs[2522]) | (layer1_outputs[2280]);
    assign layer2_outputs[1070] = ~(layer1_outputs[2361]);
    assign layer2_outputs[1071] = (layer1_outputs[1283]) & (layer1_outputs[1215]);
    assign layer2_outputs[1072] = 1'b1;
    assign layer2_outputs[1073] = ~(layer1_outputs[2260]);
    assign layer2_outputs[1074] = (layer1_outputs[2000]) ^ (layer1_outputs[1712]);
    assign layer2_outputs[1075] = ~(layer1_outputs[252]);
    assign layer2_outputs[1076] = layer1_outputs[386];
    assign layer2_outputs[1077] = ~(layer1_outputs[1850]);
    assign layer2_outputs[1078] = (layer1_outputs[1627]) & ~(layer1_outputs[2198]);
    assign layer2_outputs[1079] = 1'b1;
    assign layer2_outputs[1080] = layer1_outputs[1680];
    assign layer2_outputs[1081] = layer1_outputs[303];
    assign layer2_outputs[1082] = ~(layer1_outputs[2046]);
    assign layer2_outputs[1083] = layer1_outputs[1242];
    assign layer2_outputs[1084] = layer1_outputs[1420];
    assign layer2_outputs[1085] = ~(layer1_outputs[770]);
    assign layer2_outputs[1086] = 1'b1;
    assign layer2_outputs[1087] = (layer1_outputs[2010]) & ~(layer1_outputs[2321]);
    assign layer2_outputs[1088] = ~(layer1_outputs[67]) | (layer1_outputs[1413]);
    assign layer2_outputs[1089] = layer1_outputs[622];
    assign layer2_outputs[1090] = 1'b0;
    assign layer2_outputs[1091] = ~(layer1_outputs[1790]) | (layer1_outputs[138]);
    assign layer2_outputs[1092] = ~(layer1_outputs[1556]);
    assign layer2_outputs[1093] = layer1_outputs[672];
    assign layer2_outputs[1094] = (layer1_outputs[1893]) & ~(layer1_outputs[2024]);
    assign layer2_outputs[1095] = (layer1_outputs[2233]) & ~(layer1_outputs[406]);
    assign layer2_outputs[1096] = ~(layer1_outputs[805]) | (layer1_outputs[576]);
    assign layer2_outputs[1097] = ~(layer1_outputs[1968]);
    assign layer2_outputs[1098] = ~(layer1_outputs[1937]);
    assign layer2_outputs[1099] = (layer1_outputs[546]) & ~(layer1_outputs[2447]);
    assign layer2_outputs[1100] = (layer1_outputs[127]) | (layer1_outputs[1607]);
    assign layer2_outputs[1101] = (layer1_outputs[108]) & ~(layer1_outputs[609]);
    assign layer2_outputs[1102] = ~(layer1_outputs[1583]) | (layer1_outputs[811]);
    assign layer2_outputs[1103] = layer1_outputs[2258];
    assign layer2_outputs[1104] = ~((layer1_outputs[1002]) | (layer1_outputs[414]));
    assign layer2_outputs[1105] = (layer1_outputs[955]) & ~(layer1_outputs[2194]);
    assign layer2_outputs[1106] = ~((layer1_outputs[2461]) | (layer1_outputs[201]));
    assign layer2_outputs[1107] = (layer1_outputs[554]) & ~(layer1_outputs[255]);
    assign layer2_outputs[1108] = ~(layer1_outputs[176]);
    assign layer2_outputs[1109] = layer1_outputs[1209];
    assign layer2_outputs[1110] = layer1_outputs[389];
    assign layer2_outputs[1111] = ~((layer1_outputs[925]) ^ (layer1_outputs[1227]));
    assign layer2_outputs[1112] = layer1_outputs[1502];
    assign layer2_outputs[1113] = ~((layer1_outputs[301]) & (layer1_outputs[2257]));
    assign layer2_outputs[1114] = (layer1_outputs[1238]) | (layer1_outputs[648]);
    assign layer2_outputs[1115] = (layer1_outputs[747]) & ~(layer1_outputs[1336]);
    assign layer2_outputs[1116] = ~(layer1_outputs[2201]);
    assign layer2_outputs[1117] = layer1_outputs[637];
    assign layer2_outputs[1118] = layer1_outputs[244];
    assign layer2_outputs[1119] = layer1_outputs[1900];
    assign layer2_outputs[1120] = layer1_outputs[1115];
    assign layer2_outputs[1121] = ~((layer1_outputs[1975]) & (layer1_outputs[62]));
    assign layer2_outputs[1122] = (layer1_outputs[2394]) & ~(layer1_outputs[586]);
    assign layer2_outputs[1123] = (layer1_outputs[82]) & (layer1_outputs[1371]);
    assign layer2_outputs[1124] = (layer1_outputs[1784]) & ~(layer1_outputs[2552]);
    assign layer2_outputs[1125] = ~(layer1_outputs[42]);
    assign layer2_outputs[1126] = ~((layer1_outputs[1293]) & (layer1_outputs[831]));
    assign layer2_outputs[1127] = ~(layer1_outputs[1430]);
    assign layer2_outputs[1128] = (layer1_outputs[1077]) & ~(layer1_outputs[545]);
    assign layer2_outputs[1129] = layer1_outputs[2057];
    assign layer2_outputs[1130] = ~((layer1_outputs[1250]) | (layer1_outputs[857]));
    assign layer2_outputs[1131] = (layer1_outputs[2179]) & (layer1_outputs[2140]);
    assign layer2_outputs[1132] = ~(layer1_outputs[2099]) | (layer1_outputs[1902]);
    assign layer2_outputs[1133] = ~(layer1_outputs[2067]) | (layer1_outputs[575]);
    assign layer2_outputs[1134] = (layer1_outputs[477]) ^ (layer1_outputs[2288]);
    assign layer2_outputs[1135] = (layer1_outputs[1661]) & (layer1_outputs[2335]);
    assign layer2_outputs[1136] = ~(layer1_outputs[1959]);
    assign layer2_outputs[1137] = ~(layer1_outputs[1600]);
    assign layer2_outputs[1138] = (layer1_outputs[1104]) & (layer1_outputs[343]);
    assign layer2_outputs[1139] = layer1_outputs[259];
    assign layer2_outputs[1140] = 1'b1;
    assign layer2_outputs[1141] = ~(layer1_outputs[2277]);
    assign layer2_outputs[1142] = layer1_outputs[532];
    assign layer2_outputs[1143] = ~(layer1_outputs[1775]) | (layer1_outputs[2401]);
    assign layer2_outputs[1144] = ~(layer1_outputs[1000]) | (layer1_outputs[1655]);
    assign layer2_outputs[1145] = (layer1_outputs[677]) & ~(layer1_outputs[743]);
    assign layer2_outputs[1146] = (layer1_outputs[1792]) & (layer1_outputs[1532]);
    assign layer2_outputs[1147] = ~(layer1_outputs[1662]);
    assign layer2_outputs[1148] = ~((layer1_outputs[1860]) ^ (layer1_outputs[1245]));
    assign layer2_outputs[1149] = layer1_outputs[1053];
    assign layer2_outputs[1150] = (layer1_outputs[1356]) & ~(layer1_outputs[1224]);
    assign layer2_outputs[1151] = ~((layer1_outputs[237]) | (layer1_outputs[1281]));
    assign layer2_outputs[1152] = ~((layer1_outputs[91]) & (layer1_outputs[1042]));
    assign layer2_outputs[1153] = ~(layer1_outputs[2342]);
    assign layer2_outputs[1154] = (layer1_outputs[942]) | (layer1_outputs[1668]);
    assign layer2_outputs[1155] = (layer1_outputs[1807]) ^ (layer1_outputs[396]);
    assign layer2_outputs[1156] = layer1_outputs[750];
    assign layer2_outputs[1157] = (layer1_outputs[1288]) & ~(layer1_outputs[1113]);
    assign layer2_outputs[1158] = ~(layer1_outputs[439]);
    assign layer2_outputs[1159] = ~((layer1_outputs[491]) | (layer1_outputs[2215]));
    assign layer2_outputs[1160] = ~((layer1_outputs[732]) | (layer1_outputs[1522]));
    assign layer2_outputs[1161] = ~(layer1_outputs[116]);
    assign layer2_outputs[1162] = layer1_outputs[2340];
    assign layer2_outputs[1163] = ~(layer1_outputs[274]);
    assign layer2_outputs[1164] = ~(layer1_outputs[1565]);
    assign layer2_outputs[1165] = 1'b0;
    assign layer2_outputs[1166] = ~((layer1_outputs[2377]) & (layer1_outputs[277]));
    assign layer2_outputs[1167] = ~(layer1_outputs[2343]) | (layer1_outputs[567]);
    assign layer2_outputs[1168] = (layer1_outputs[1670]) & ~(layer1_outputs[1175]);
    assign layer2_outputs[1169] = ~(layer1_outputs[1852]) | (layer1_outputs[1417]);
    assign layer2_outputs[1170] = ~(layer1_outputs[631]) | (layer1_outputs[1075]);
    assign layer2_outputs[1171] = ~((layer1_outputs[1982]) ^ (layer1_outputs[559]));
    assign layer2_outputs[1172] = (layer1_outputs[1335]) ^ (layer1_outputs[913]);
    assign layer2_outputs[1173] = layer1_outputs[697];
    assign layer2_outputs[1174] = ~(layer1_outputs[2267]) | (layer1_outputs[321]);
    assign layer2_outputs[1175] = ~(layer1_outputs[1967]);
    assign layer2_outputs[1176] = layer1_outputs[1515];
    assign layer2_outputs[1177] = ~(layer1_outputs[886]);
    assign layer2_outputs[1178] = 1'b0;
    assign layer2_outputs[1179] = 1'b0;
    assign layer2_outputs[1180] = ~(layer1_outputs[372]);
    assign layer2_outputs[1181] = layer1_outputs[320];
    assign layer2_outputs[1182] = (layer1_outputs[1168]) & (layer1_outputs[2247]);
    assign layer2_outputs[1183] = ~((layer1_outputs[694]) ^ (layer1_outputs[30]));
    assign layer2_outputs[1184] = (layer1_outputs[585]) & ~(layer1_outputs[1872]);
    assign layer2_outputs[1185] = 1'b0;
    assign layer2_outputs[1186] = ~(layer1_outputs[1297]);
    assign layer2_outputs[1187] = layer1_outputs[2050];
    assign layer2_outputs[1188] = ~(layer1_outputs[1338]);
    assign layer2_outputs[1189] = (layer1_outputs[496]) & ~(layer1_outputs[1142]);
    assign layer2_outputs[1190] = (layer1_outputs[248]) & (layer1_outputs[733]);
    assign layer2_outputs[1191] = ~((layer1_outputs[2136]) ^ (layer1_outputs[2510]));
    assign layer2_outputs[1192] = (layer1_outputs[540]) & ~(layer1_outputs[1735]);
    assign layer2_outputs[1193] = 1'b0;
    assign layer2_outputs[1194] = layer1_outputs[1458];
    assign layer2_outputs[1195] = layer1_outputs[300];
    assign layer2_outputs[1196] = ~(layer1_outputs[468]);
    assign layer2_outputs[1197] = layer1_outputs[1942];
    assign layer2_outputs[1198] = ~((layer1_outputs[842]) | (layer1_outputs[2326]));
    assign layer2_outputs[1199] = (layer1_outputs[701]) & (layer1_outputs[1915]);
    assign layer2_outputs[1200] = (layer1_outputs[1798]) | (layer1_outputs[1133]);
    assign layer2_outputs[1201] = ~(layer1_outputs[1813]) | (layer1_outputs[1341]);
    assign layer2_outputs[1202] = ~(layer1_outputs[1527]) | (layer1_outputs[1209]);
    assign layer2_outputs[1203] = layer1_outputs[780];
    assign layer2_outputs[1204] = ~((layer1_outputs[1276]) | (layer1_outputs[924]));
    assign layer2_outputs[1205] = (layer1_outputs[1167]) & (layer1_outputs[1888]);
    assign layer2_outputs[1206] = layer1_outputs[2030];
    assign layer2_outputs[1207] = (layer1_outputs[836]) & ~(layer1_outputs[2541]);
    assign layer2_outputs[1208] = 1'b1;
    assign layer2_outputs[1209] = ~(layer1_outputs[2474]);
    assign layer2_outputs[1210] = layer1_outputs[1577];
    assign layer2_outputs[1211] = ~(layer1_outputs[1163]);
    assign layer2_outputs[1212] = ~(layer1_outputs[1774]) | (layer1_outputs[1811]);
    assign layer2_outputs[1213] = ~((layer1_outputs[1028]) | (layer1_outputs[1118]));
    assign layer2_outputs[1214] = 1'b0;
    assign layer2_outputs[1215] = ~((layer1_outputs[7]) | (layer1_outputs[1318]));
    assign layer2_outputs[1216] = 1'b0;
    assign layer2_outputs[1217] = 1'b0;
    assign layer2_outputs[1218] = (layer1_outputs[1314]) & (layer1_outputs[602]);
    assign layer2_outputs[1219] = ~(layer1_outputs[842]) | (layer1_outputs[1824]);
    assign layer2_outputs[1220] = ~(layer1_outputs[2328]);
    assign layer2_outputs[1221] = ~(layer1_outputs[1062]);
    assign layer2_outputs[1222] = ~((layer1_outputs[2303]) | (layer1_outputs[1575]));
    assign layer2_outputs[1223] = layer1_outputs[1364];
    assign layer2_outputs[1224] = ~((layer1_outputs[242]) & (layer1_outputs[1413]));
    assign layer2_outputs[1225] = ~((layer1_outputs[164]) & (layer1_outputs[2231]));
    assign layer2_outputs[1226] = 1'b0;
    assign layer2_outputs[1227] = ~(layer1_outputs[1122]);
    assign layer2_outputs[1228] = ~(layer1_outputs[1536]);
    assign layer2_outputs[1229] = ~(layer1_outputs[2084]);
    assign layer2_outputs[1230] = (layer1_outputs[2174]) | (layer1_outputs[2136]);
    assign layer2_outputs[1231] = 1'b0;
    assign layer2_outputs[1232] = ~(layer1_outputs[2228]) | (layer1_outputs[1833]);
    assign layer2_outputs[1233] = (layer1_outputs[1671]) & ~(layer1_outputs[379]);
    assign layer2_outputs[1234] = ~((layer1_outputs[2525]) | (layer1_outputs[2090]));
    assign layer2_outputs[1235] = layer1_outputs[1815];
    assign layer2_outputs[1236] = ~(layer1_outputs[1166]) | (layer1_outputs[1283]);
    assign layer2_outputs[1237] = 1'b0;
    assign layer2_outputs[1238] = ~(layer1_outputs[1392]);
    assign layer2_outputs[1239] = (layer1_outputs[428]) & ~(layer1_outputs[778]);
    assign layer2_outputs[1240] = ~(layer1_outputs[1800]) | (layer1_outputs[685]);
    assign layer2_outputs[1241] = layer1_outputs[1339];
    assign layer2_outputs[1242] = 1'b1;
    assign layer2_outputs[1243] = ~(layer1_outputs[949]);
    assign layer2_outputs[1244] = ~(layer1_outputs[292]) | (layer1_outputs[2525]);
    assign layer2_outputs[1245] = ~(layer1_outputs[539]) | (layer1_outputs[129]);
    assign layer2_outputs[1246] = ~(layer1_outputs[1369]);
    assign layer2_outputs[1247] = ~((layer1_outputs[1732]) | (layer1_outputs[2209]));
    assign layer2_outputs[1248] = layer1_outputs[2390];
    assign layer2_outputs[1249] = (layer1_outputs[2303]) | (layer1_outputs[2218]);
    assign layer2_outputs[1250] = (layer1_outputs[2083]) | (layer1_outputs[2462]);
    assign layer2_outputs[1251] = ~(layer1_outputs[686]);
    assign layer2_outputs[1252] = ~(layer1_outputs[1065]) | (layer1_outputs[495]);
    assign layer2_outputs[1253] = layer1_outputs[935];
    assign layer2_outputs[1254] = (layer1_outputs[2417]) & ~(layer1_outputs[1340]);
    assign layer2_outputs[1255] = (layer1_outputs[1105]) & ~(layer1_outputs[1100]);
    assign layer2_outputs[1256] = (layer1_outputs[108]) & (layer1_outputs[1277]);
    assign layer2_outputs[1257] = 1'b1;
    assign layer2_outputs[1258] = layer1_outputs[798];
    assign layer2_outputs[1259] = ~(layer1_outputs[2344]);
    assign layer2_outputs[1260] = (layer1_outputs[1530]) & ~(layer1_outputs[1141]);
    assign layer2_outputs[1261] = ~(layer1_outputs[432]);
    assign layer2_outputs[1262] = (layer1_outputs[1706]) & ~(layer1_outputs[262]);
    assign layer2_outputs[1263] = layer1_outputs[2532];
    assign layer2_outputs[1264] = layer1_outputs[2459];
    assign layer2_outputs[1265] = ~(layer1_outputs[2325]);
    assign layer2_outputs[1266] = (layer1_outputs[368]) & ~(layer1_outputs[893]);
    assign layer2_outputs[1267] = ~(layer1_outputs[1222]);
    assign layer2_outputs[1268] = ~((layer1_outputs[1404]) | (layer1_outputs[649]));
    assign layer2_outputs[1269] = layer1_outputs[1394];
    assign layer2_outputs[1270] = ~((layer1_outputs[2383]) & (layer1_outputs[704]));
    assign layer2_outputs[1271] = ~(layer1_outputs[1172]);
    assign layer2_outputs[1272] = (layer1_outputs[2370]) & (layer1_outputs[2241]);
    assign layer2_outputs[1273] = (layer1_outputs[1657]) & ~(layer1_outputs[468]);
    assign layer2_outputs[1274] = ~(layer1_outputs[1300]) | (layer1_outputs[131]);
    assign layer2_outputs[1275] = layer1_outputs[1126];
    assign layer2_outputs[1276] = ~(layer1_outputs[2371]);
    assign layer2_outputs[1277] = layer1_outputs[1428];
    assign layer2_outputs[1278] = (layer1_outputs[2334]) & (layer1_outputs[166]);
    assign layer2_outputs[1279] = ~(layer1_outputs[552]);
    assign layer2_outputs[1280] = (layer1_outputs[1342]) | (layer1_outputs[233]);
    assign layer2_outputs[1281] = ~(layer1_outputs[1539]) | (layer1_outputs[912]);
    assign layer2_outputs[1282] = 1'b0;
    assign layer2_outputs[1283] = ~(layer1_outputs[1618]);
    assign layer2_outputs[1284] = ~(layer1_outputs[2069]);
    assign layer2_outputs[1285] = ~(layer1_outputs[541]);
    assign layer2_outputs[1286] = (layer1_outputs[1710]) ^ (layer1_outputs[359]);
    assign layer2_outputs[1287] = ~(layer1_outputs[415]);
    assign layer2_outputs[1288] = (layer1_outputs[1839]) & ~(layer1_outputs[170]);
    assign layer2_outputs[1289] = (layer1_outputs[106]) & ~(layer1_outputs[21]);
    assign layer2_outputs[1290] = (layer1_outputs[2416]) & (layer1_outputs[1179]);
    assign layer2_outputs[1291] = ~(layer1_outputs[2398]) | (layer1_outputs[1662]);
    assign layer2_outputs[1292] = ~(layer1_outputs[2464]) | (layer1_outputs[725]);
    assign layer2_outputs[1293] = ~(layer1_outputs[535]);
    assign layer2_outputs[1294] = (layer1_outputs[751]) & ~(layer1_outputs[1776]);
    assign layer2_outputs[1295] = ~(layer1_outputs[1418]) | (layer1_outputs[661]);
    assign layer2_outputs[1296] = ~((layer1_outputs[2177]) & (layer1_outputs[2092]));
    assign layer2_outputs[1297] = layer1_outputs[964];
    assign layer2_outputs[1298] = ~(layer1_outputs[2224]);
    assign layer2_outputs[1299] = ~(layer1_outputs[2544]);
    assign layer2_outputs[1300] = ~(layer1_outputs[1244]);
    assign layer2_outputs[1301] = ~((layer1_outputs[398]) & (layer1_outputs[1154]));
    assign layer2_outputs[1302] = ~(layer1_outputs[2451]);
    assign layer2_outputs[1303] = ~(layer1_outputs[848]);
    assign layer2_outputs[1304] = ~(layer1_outputs[2108]);
    assign layer2_outputs[1305] = 1'b1;
    assign layer2_outputs[1306] = ~((layer1_outputs[919]) ^ (layer1_outputs[833]));
    assign layer2_outputs[1307] = ~(layer1_outputs[789]);
    assign layer2_outputs[1308] = ~(layer1_outputs[2455]);
    assign layer2_outputs[1309] = (layer1_outputs[1197]) ^ (layer1_outputs[2188]);
    assign layer2_outputs[1310] = (layer1_outputs[1965]) & ~(layer1_outputs[688]);
    assign layer2_outputs[1311] = (layer1_outputs[2071]) & ~(layer1_outputs[1966]);
    assign layer2_outputs[1312] = ~((layer1_outputs[1088]) | (layer1_outputs[984]));
    assign layer2_outputs[1313] = 1'b0;
    assign layer2_outputs[1314] = (layer1_outputs[1260]) & ~(layer1_outputs[1981]);
    assign layer2_outputs[1315] = ~(layer1_outputs[139]);
    assign layer2_outputs[1316] = ~(layer1_outputs[923]);
    assign layer2_outputs[1317] = layer1_outputs[2494];
    assign layer2_outputs[1318] = layer1_outputs[202];
    assign layer2_outputs[1319] = ~((layer1_outputs[2036]) & (layer1_outputs[596]));
    assign layer2_outputs[1320] = layer1_outputs[1577];
    assign layer2_outputs[1321] = (layer1_outputs[236]) ^ (layer1_outputs[1704]);
    assign layer2_outputs[1322] = ~(layer1_outputs[2537]) | (layer1_outputs[233]);
    assign layer2_outputs[1323] = 1'b1;
    assign layer2_outputs[1324] = ~(layer1_outputs[2061]) | (layer1_outputs[1333]);
    assign layer2_outputs[1325] = ~(layer1_outputs[1192]);
    assign layer2_outputs[1326] = ~(layer1_outputs[433]);
    assign layer2_outputs[1327] = (layer1_outputs[596]) & ~(layer1_outputs[1166]);
    assign layer2_outputs[1328] = ~(layer1_outputs[708]) | (layer1_outputs[148]);
    assign layer2_outputs[1329] = 1'b0;
    assign layer2_outputs[1330] = ~(layer1_outputs[1742]);
    assign layer2_outputs[1331] = ~(layer1_outputs[617]);
    assign layer2_outputs[1332] = ~((layer1_outputs[1463]) & (layer1_outputs[1384]));
    assign layer2_outputs[1333] = layer1_outputs[615];
    assign layer2_outputs[1334] = ~(layer1_outputs[2130]);
    assign layer2_outputs[1335] = layer1_outputs[597];
    assign layer2_outputs[1336] = (layer1_outputs[365]) & ~(layer1_outputs[1108]);
    assign layer2_outputs[1337] = (layer1_outputs[1455]) | (layer1_outputs[2150]);
    assign layer2_outputs[1338] = layer1_outputs[2422];
    assign layer2_outputs[1339] = (layer1_outputs[76]) & ~(layer1_outputs[505]);
    assign layer2_outputs[1340] = layer1_outputs[1556];
    assign layer2_outputs[1341] = ~(layer1_outputs[2037]);
    assign layer2_outputs[1342] = (layer1_outputs[1274]) & ~(layer1_outputs[548]);
    assign layer2_outputs[1343] = ~((layer1_outputs[1089]) | (layer1_outputs[1779]));
    assign layer2_outputs[1344] = ~(layer1_outputs[780]);
    assign layer2_outputs[1345] = 1'b0;
    assign layer2_outputs[1346] = layer1_outputs[2453];
    assign layer2_outputs[1347] = (layer1_outputs[299]) ^ (layer1_outputs[2413]);
    assign layer2_outputs[1348] = layer1_outputs[1487];
    assign layer2_outputs[1349] = (layer1_outputs[1268]) & ~(layer1_outputs[571]);
    assign layer2_outputs[1350] = ~(layer1_outputs[2499]) | (layer1_outputs[1423]);
    assign layer2_outputs[1351] = layer1_outputs[454];
    assign layer2_outputs[1352] = ~(layer1_outputs[1038]) | (layer1_outputs[551]);
    assign layer2_outputs[1353] = ~(layer1_outputs[1316]);
    assign layer2_outputs[1354] = layer1_outputs[1080];
    assign layer2_outputs[1355] = ~((layer1_outputs[1529]) & (layer1_outputs[2216]));
    assign layer2_outputs[1356] = ~(layer1_outputs[405]) | (layer1_outputs[2349]);
    assign layer2_outputs[1357] = (layer1_outputs[1919]) | (layer1_outputs[1566]);
    assign layer2_outputs[1358] = (layer1_outputs[413]) & (layer1_outputs[775]);
    assign layer2_outputs[1359] = (layer1_outputs[117]) & (layer1_outputs[909]);
    assign layer2_outputs[1360] = ~(layer1_outputs[2470]) | (layer1_outputs[351]);
    assign layer2_outputs[1361] = layer1_outputs[103];
    assign layer2_outputs[1362] = layer1_outputs[1419];
    assign layer2_outputs[1363] = ~((layer1_outputs[543]) ^ (layer1_outputs[1310]));
    assign layer2_outputs[1364] = ~(layer1_outputs[2205]) | (layer1_outputs[1722]);
    assign layer2_outputs[1365] = layer1_outputs[2534];
    assign layer2_outputs[1366] = ~(layer1_outputs[901]);
    assign layer2_outputs[1367] = (layer1_outputs[1580]) & (layer1_outputs[1021]);
    assign layer2_outputs[1368] = ~(layer1_outputs[134]);
    assign layer2_outputs[1369] = (layer1_outputs[398]) & ~(layer1_outputs[1940]);
    assign layer2_outputs[1370] = ~((layer1_outputs[479]) | (layer1_outputs[894]));
    assign layer2_outputs[1371] = 1'b0;
    assign layer2_outputs[1372] = ~((layer1_outputs[2185]) ^ (layer1_outputs[1272]));
    assign layer2_outputs[1373] = ~(layer1_outputs[155]) | (layer1_outputs[2082]);
    assign layer2_outputs[1374] = ~((layer1_outputs[1320]) & (layer1_outputs[474]));
    assign layer2_outputs[1375] = ~(layer1_outputs[395]);
    assign layer2_outputs[1376] = (layer1_outputs[1743]) & ~(layer1_outputs[1608]);
    assign layer2_outputs[1377] = layer1_outputs[1992];
    assign layer2_outputs[1378] = ~(layer1_outputs[1759]);
    assign layer2_outputs[1379] = (layer1_outputs[422]) & ~(layer1_outputs[526]);
    assign layer2_outputs[1380] = 1'b1;
    assign layer2_outputs[1381] = ~(layer1_outputs[2187]);
    assign layer2_outputs[1382] = 1'b1;
    assign layer2_outputs[1383] = (layer1_outputs[1480]) & ~(layer1_outputs[1537]);
    assign layer2_outputs[1384] = 1'b1;
    assign layer2_outputs[1385] = ~(layer1_outputs[492]);
    assign layer2_outputs[1386] = (layer1_outputs[1178]) & (layer1_outputs[2417]);
    assign layer2_outputs[1387] = ~(layer1_outputs[201]);
    assign layer2_outputs[1388] = ~(layer1_outputs[1034]) | (layer1_outputs[2295]);
    assign layer2_outputs[1389] = (layer1_outputs[60]) | (layer1_outputs[1434]);
    assign layer2_outputs[1390] = layer1_outputs[990];
    assign layer2_outputs[1391] = layer1_outputs[868];
    assign layer2_outputs[1392] = ~(layer1_outputs[1552]);
    assign layer2_outputs[1393] = ~(layer1_outputs[2482]);
    assign layer2_outputs[1394] = layer1_outputs[790];
    assign layer2_outputs[1395] = layer1_outputs[1010];
    assign layer2_outputs[1396] = ~(layer1_outputs[1793]);
    assign layer2_outputs[1397] = ~(layer1_outputs[1941]);
    assign layer2_outputs[1398] = ~(layer1_outputs[2165]);
    assign layer2_outputs[1399] = ~(layer1_outputs[2107]);
    assign layer2_outputs[1400] = ~((layer1_outputs[2253]) & (layer1_outputs[2070]));
    assign layer2_outputs[1401] = ~(layer1_outputs[1954]);
    assign layer2_outputs[1402] = ~(layer1_outputs[2141]);
    assign layer2_outputs[1403] = ~(layer1_outputs[1366]) | (layer1_outputs[788]);
    assign layer2_outputs[1404] = ~(layer1_outputs[555]);
    assign layer2_outputs[1405] = ~(layer1_outputs[462]);
    assign layer2_outputs[1406] = ~(layer1_outputs[1165]);
    assign layer2_outputs[1407] = layer1_outputs[1116];
    assign layer2_outputs[1408] = ~(layer1_outputs[607]) | (layer1_outputs[836]);
    assign layer2_outputs[1409] = (layer1_outputs[168]) | (layer1_outputs[772]);
    assign layer2_outputs[1410] = ~(layer1_outputs[646]);
    assign layer2_outputs[1411] = 1'b0;
    assign layer2_outputs[1412] = ~((layer1_outputs[1297]) | (layer1_outputs[1347]));
    assign layer2_outputs[1413] = layer1_outputs[663];
    assign layer2_outputs[1414] = ~(layer1_outputs[1936]);
    assign layer2_outputs[1415] = ~(layer1_outputs[2041]) | (layer1_outputs[816]);
    assign layer2_outputs[1416] = 1'b0;
    assign layer2_outputs[1417] = ~(layer1_outputs[667]);
    assign layer2_outputs[1418] = layer1_outputs[749];
    assign layer2_outputs[1419] = ~((layer1_outputs[2008]) ^ (layer1_outputs[1026]));
    assign layer2_outputs[1420] = (layer1_outputs[769]) & ~(layer1_outputs[415]);
    assign layer2_outputs[1421] = ~((layer1_outputs[570]) & (layer1_outputs[2102]));
    assign layer2_outputs[1422] = ~(layer1_outputs[909]);
    assign layer2_outputs[1423] = (layer1_outputs[707]) | (layer1_outputs[2485]);
    assign layer2_outputs[1424] = ~(layer1_outputs[482]) | (layer1_outputs[2383]);
    assign layer2_outputs[1425] = 1'b0;
    assign layer2_outputs[1426] = (layer1_outputs[2009]) & ~(layer1_outputs[2454]);
    assign layer2_outputs[1427] = ~(layer1_outputs[1789]);
    assign layer2_outputs[1428] = ~((layer1_outputs[1525]) ^ (layer1_outputs[796]));
    assign layer2_outputs[1429] = ~(layer1_outputs[1212]);
    assign layer2_outputs[1430] = ~((layer1_outputs[1570]) & (layer1_outputs[1128]));
    assign layer2_outputs[1431] = layer1_outputs[367];
    assign layer2_outputs[1432] = ~((layer1_outputs[1850]) & (layer1_outputs[1432]));
    assign layer2_outputs[1433] = 1'b1;
    assign layer2_outputs[1434] = ~(layer1_outputs[407]);
    assign layer2_outputs[1435] = ~((layer1_outputs[1930]) ^ (layer1_outputs[2345]));
    assign layer2_outputs[1436] = ~(layer1_outputs[2407]) | (layer1_outputs[827]);
    assign layer2_outputs[1437] = ~(layer1_outputs[1098]);
    assign layer2_outputs[1438] = ~(layer1_outputs[2289]) | (layer1_outputs[131]);
    assign layer2_outputs[1439] = ~(layer1_outputs[2226]);
    assign layer2_outputs[1440] = ~(layer1_outputs[1787]);
    assign layer2_outputs[1441] = (layer1_outputs[560]) & (layer1_outputs[1608]);
    assign layer2_outputs[1442] = (layer1_outputs[183]) & ~(layer1_outputs[556]);
    assign layer2_outputs[1443] = 1'b0;
    assign layer2_outputs[1444] = ~(layer1_outputs[537]);
    assign layer2_outputs[1445] = (layer1_outputs[2140]) & ~(layer1_outputs[325]);
    assign layer2_outputs[1446] = ~((layer1_outputs[674]) ^ (layer1_outputs[2337]));
    assign layer2_outputs[1447] = ~(layer1_outputs[1363]);
    assign layer2_outputs[1448] = ~((layer1_outputs[2269]) & (layer1_outputs[1170]));
    assign layer2_outputs[1449] = layer1_outputs[1985];
    assign layer2_outputs[1450] = ~((layer1_outputs[31]) & (layer1_outputs[1669]));
    assign layer2_outputs[1451] = (layer1_outputs[1614]) | (layer1_outputs[1960]);
    assign layer2_outputs[1452] = layer1_outputs[1108];
    assign layer2_outputs[1453] = (layer1_outputs[339]) & ~(layer1_outputs[175]);
    assign layer2_outputs[1454] = (layer1_outputs[186]) & ~(layer1_outputs[1543]);
    assign layer2_outputs[1455] = layer1_outputs[853];
    assign layer2_outputs[1456] = layer1_outputs[392];
    assign layer2_outputs[1457] = (layer1_outputs[585]) | (layer1_outputs[612]);
    assign layer2_outputs[1458] = (layer1_outputs[1397]) & ~(layer1_outputs[1074]);
    assign layer2_outputs[1459] = ~(layer1_outputs[1254]);
    assign layer2_outputs[1460] = 1'b0;
    assign layer2_outputs[1461] = layer1_outputs[1451];
    assign layer2_outputs[1462] = layer1_outputs[1779];
    assign layer2_outputs[1463] = layer1_outputs[1847];
    assign layer2_outputs[1464] = (layer1_outputs[335]) & (layer1_outputs[1622]);
    assign layer2_outputs[1465] = (layer1_outputs[86]) & ~(layer1_outputs[930]);
    assign layer2_outputs[1466] = ~((layer1_outputs[2532]) | (layer1_outputs[326]));
    assign layer2_outputs[1467] = layer1_outputs[1712];
    assign layer2_outputs[1468] = layer1_outputs[996];
    assign layer2_outputs[1469] = ~(layer1_outputs[849]);
    assign layer2_outputs[1470] = layer1_outputs[551];
    assign layer2_outputs[1471] = (layer1_outputs[1435]) & ~(layer1_outputs[110]);
    assign layer2_outputs[1472] = (layer1_outputs[921]) & (layer1_outputs[1880]);
    assign layer2_outputs[1473] = layer1_outputs[990];
    assign layer2_outputs[1474] = (layer1_outputs[1921]) | (layer1_outputs[1348]);
    assign layer2_outputs[1475] = (layer1_outputs[9]) & ~(layer1_outputs[11]);
    assign layer2_outputs[1476] = layer1_outputs[1719];
    assign layer2_outputs[1477] = ~(layer1_outputs[621]) | (layer1_outputs[779]);
    assign layer2_outputs[1478] = ~((layer1_outputs[1426]) ^ (layer1_outputs[1177]));
    assign layer2_outputs[1479] = ~(layer1_outputs[2275]);
    assign layer2_outputs[1480] = layer1_outputs[1161];
    assign layer2_outputs[1481] = layer1_outputs[1277];
    assign layer2_outputs[1482] = 1'b1;
    assign layer2_outputs[1483] = ~((layer1_outputs[1473]) | (layer1_outputs[1353]));
    assign layer2_outputs[1484] = ~(layer1_outputs[1517]) | (layer1_outputs[726]);
    assign layer2_outputs[1485] = ~(layer1_outputs[1132]);
    assign layer2_outputs[1486] = ~((layer1_outputs[473]) & (layer1_outputs[2349]));
    assign layer2_outputs[1487] = (layer1_outputs[594]) & (layer1_outputs[736]);
    assign layer2_outputs[1488] = (layer1_outputs[46]) & ~(layer1_outputs[874]);
    assign layer2_outputs[1489] = ~(layer1_outputs[1773]) | (layer1_outputs[899]);
    assign layer2_outputs[1490] = ~(layer1_outputs[44]);
    assign layer2_outputs[1491] = ~(layer1_outputs[1248]);
    assign layer2_outputs[1492] = ~((layer1_outputs[876]) | (layer1_outputs[549]));
    assign layer2_outputs[1493] = (layer1_outputs[700]) & ~(layer1_outputs[1705]);
    assign layer2_outputs[1494] = (layer1_outputs[135]) & ~(layer1_outputs[183]);
    assign layer2_outputs[1495] = (layer1_outputs[2156]) | (layer1_outputs[329]);
    assign layer2_outputs[1496] = (layer1_outputs[784]) | (layer1_outputs[1301]);
    assign layer2_outputs[1497] = ~(layer1_outputs[110]);
    assign layer2_outputs[1498] = 1'b1;
    assign layer2_outputs[1499] = (layer1_outputs[862]) ^ (layer1_outputs[1552]);
    assign layer2_outputs[1500] = ~(layer1_outputs[923]);
    assign layer2_outputs[1501] = ~(layer1_outputs[1271]);
    assign layer2_outputs[1502] = (layer1_outputs[705]) & ~(layer1_outputs[1560]);
    assign layer2_outputs[1503] = ~(layer1_outputs[12]) | (layer1_outputs[662]);
    assign layer2_outputs[1504] = ~((layer1_outputs[1109]) & (layer1_outputs[1485]));
    assign layer2_outputs[1505] = layer1_outputs[226];
    assign layer2_outputs[1506] = ~((layer1_outputs[2204]) & (layer1_outputs[1532]));
    assign layer2_outputs[1507] = 1'b1;
    assign layer2_outputs[1508] = ~((layer1_outputs[1760]) & (layer1_outputs[1399]));
    assign layer2_outputs[1509] = layer1_outputs[1411];
    assign layer2_outputs[1510] = (layer1_outputs[704]) & ~(layer1_outputs[2379]);
    assign layer2_outputs[1511] = ~((layer1_outputs[1998]) & (layer1_outputs[610]));
    assign layer2_outputs[1512] = layer1_outputs[858];
    assign layer2_outputs[1513] = layer1_outputs[2537];
    assign layer2_outputs[1514] = (layer1_outputs[675]) & ~(layer1_outputs[2389]);
    assign layer2_outputs[1515] = (layer1_outputs[150]) & ~(layer1_outputs[1240]);
    assign layer2_outputs[1516] = ~(layer1_outputs[425]);
    assign layer2_outputs[1517] = ~(layer1_outputs[2316]);
    assign layer2_outputs[1518] = (layer1_outputs[2004]) & ~(layer1_outputs[298]);
    assign layer2_outputs[1519] = (layer1_outputs[1885]) & ~(layer1_outputs[1466]);
    assign layer2_outputs[1520] = 1'b1;
    assign layer2_outputs[1521] = ~(layer1_outputs[1935]) | (layer1_outputs[1587]);
    assign layer2_outputs[1522] = ~((layer1_outputs[739]) & (layer1_outputs[1920]));
    assign layer2_outputs[1523] = (layer1_outputs[1102]) & ~(layer1_outputs[383]);
    assign layer2_outputs[1524] = ~(layer1_outputs[1041]) | (layer1_outputs[1637]);
    assign layer2_outputs[1525] = layer1_outputs[2488];
    assign layer2_outputs[1526] = ~(layer1_outputs[2293]);
    assign layer2_outputs[1527] = 1'b1;
    assign layer2_outputs[1528] = ~((layer1_outputs[945]) & (layer1_outputs[905]));
    assign layer2_outputs[1529] = ~(layer1_outputs[459]);
    assign layer2_outputs[1530] = (layer1_outputs[1091]) & ~(layer1_outputs[1200]);
    assign layer2_outputs[1531] = layer1_outputs[2494];
    assign layer2_outputs[1532] = ~(layer1_outputs[1228]) | (layer1_outputs[1450]);
    assign layer2_outputs[1533] = layer1_outputs[1913];
    assign layer2_outputs[1534] = (layer1_outputs[2161]) & (layer1_outputs[2419]);
    assign layer2_outputs[1535] = layer1_outputs[1564];
    assign layer2_outputs[1536] = (layer1_outputs[1920]) & ~(layer1_outputs[1061]);
    assign layer2_outputs[1537] = (layer1_outputs[2450]) & (layer1_outputs[630]);
    assign layer2_outputs[1538] = (layer1_outputs[2222]) & (layer1_outputs[1855]);
    assign layer2_outputs[1539] = ~(layer1_outputs[509]) | (layer1_outputs[1003]);
    assign layer2_outputs[1540] = (layer1_outputs[1250]) | (layer1_outputs[1980]);
    assign layer2_outputs[1541] = layer1_outputs[377];
    assign layer2_outputs[1542] = (layer1_outputs[1653]) | (layer1_outputs[1976]);
    assign layer2_outputs[1543] = ~(layer1_outputs[99]);
    assign layer2_outputs[1544] = ~((layer1_outputs[1164]) ^ (layer1_outputs[50]));
    assign layer2_outputs[1545] = (layer1_outputs[1957]) | (layer1_outputs[74]);
    assign layer2_outputs[1546] = ~(layer1_outputs[2343]);
    assign layer2_outputs[1547] = (layer1_outputs[451]) | (layer1_outputs[1216]);
    assign layer2_outputs[1548] = ~((layer1_outputs[437]) | (layer1_outputs[1457]));
    assign layer2_outputs[1549] = ~((layer1_outputs[542]) ^ (layer1_outputs[1785]));
    assign layer2_outputs[1550] = layer1_outputs[1811];
    assign layer2_outputs[1551] = layer1_outputs[1557];
    assign layer2_outputs[1552] = 1'b0;
    assign layer2_outputs[1553] = ~((layer1_outputs[928]) & (layer1_outputs[294]));
    assign layer2_outputs[1554] = ~(layer1_outputs[1778]);
    assign layer2_outputs[1555] = layer1_outputs[1613];
    assign layer2_outputs[1556] = ~((layer1_outputs[848]) & (layer1_outputs[1810]));
    assign layer2_outputs[1557] = 1'b1;
    assign layer2_outputs[1558] = ~((layer1_outputs[2013]) ^ (layer1_outputs[2241]));
    assign layer2_outputs[1559] = (layer1_outputs[976]) | (layer1_outputs[1307]);
    assign layer2_outputs[1560] = ~(layer1_outputs[1690]);
    assign layer2_outputs[1561] = ~(layer1_outputs[2054]);
    assign layer2_outputs[1562] = layer1_outputs[157];
    assign layer2_outputs[1563] = 1'b1;
    assign layer2_outputs[1564] = (layer1_outputs[1457]) & ~(layer1_outputs[2530]);
    assign layer2_outputs[1565] = 1'b0;
    assign layer2_outputs[1566] = layer1_outputs[1909];
    assign layer2_outputs[1567] = layer1_outputs[1452];
    assign layer2_outputs[1568] = (layer1_outputs[759]) | (layer1_outputs[51]);
    assign layer2_outputs[1569] = ~(layer1_outputs[1767]) | (layer1_outputs[2206]);
    assign layer2_outputs[1570] = ~((layer1_outputs[1057]) | (layer1_outputs[1089]));
    assign layer2_outputs[1571] = 1'b0;
    assign layer2_outputs[1572] = ~(layer1_outputs[1990]);
    assign layer2_outputs[1573] = layer1_outputs[1217];
    assign layer2_outputs[1574] = ~((layer1_outputs[2171]) | (layer1_outputs[2079]));
    assign layer2_outputs[1575] = ~(layer1_outputs[2187]);
    assign layer2_outputs[1576] = ~(layer1_outputs[373]);
    assign layer2_outputs[1577] = (layer1_outputs[1048]) & (layer1_outputs[433]);
    assign layer2_outputs[1578] = (layer1_outputs[2161]) & ~(layer1_outputs[765]);
    assign layer2_outputs[1579] = ~(layer1_outputs[1138]);
    assign layer2_outputs[1580] = layer1_outputs[1725];
    assign layer2_outputs[1581] = 1'b0;
    assign layer2_outputs[1582] = (layer1_outputs[1760]) & ~(layer1_outputs[2169]);
    assign layer2_outputs[1583] = ~(layer1_outputs[1799]) | (layer1_outputs[65]);
    assign layer2_outputs[1584] = ~(layer1_outputs[165]);
    assign layer2_outputs[1585] = ~(layer1_outputs[2489]) | (layer1_outputs[1687]);
    assign layer2_outputs[1586] = (layer1_outputs[1730]) ^ (layer1_outputs[1650]);
    assign layer2_outputs[1587] = layer1_outputs[754];
    assign layer2_outputs[1588] = ~((layer1_outputs[1406]) & (layer1_outputs[1377]));
    assign layer2_outputs[1589] = (layer1_outputs[25]) & ~(layer1_outputs[249]);
    assign layer2_outputs[1590] = (layer1_outputs[1885]) & ~(layer1_outputs[320]);
    assign layer2_outputs[1591] = ~((layer1_outputs[1517]) | (layer1_outputs[774]));
    assign layer2_outputs[1592] = (layer1_outputs[1252]) & ~(layer1_outputs[1206]);
    assign layer2_outputs[1593] = ~(layer1_outputs[2401]);
    assign layer2_outputs[1594] = (layer1_outputs[1343]) & ~(layer1_outputs[6]);
    assign layer2_outputs[1595] = layer1_outputs[1929];
    assign layer2_outputs[1596] = ~(layer1_outputs[962]) | (layer1_outputs[1162]);
    assign layer2_outputs[1597] = (layer1_outputs[949]) & ~(layer1_outputs[270]);
    assign layer2_outputs[1598] = ~((layer1_outputs[446]) | (layer1_outputs[623]));
    assign layer2_outputs[1599] = (layer1_outputs[1377]) & ~(layer1_outputs[1857]);
    assign layer2_outputs[1600] = ~(layer1_outputs[1593]) | (layer1_outputs[1756]);
    assign layer2_outputs[1601] = ~(layer1_outputs[1063]) | (layer1_outputs[402]);
    assign layer2_outputs[1602] = (layer1_outputs[2341]) | (layer1_outputs[2023]);
    assign layer2_outputs[1603] = (layer1_outputs[1184]) & (layer1_outputs[1402]);
    assign layer2_outputs[1604] = layer1_outputs[1777];
    assign layer2_outputs[1605] = layer1_outputs[1926];
    assign layer2_outputs[1606] = 1'b0;
    assign layer2_outputs[1607] = layer1_outputs[507];
    assign layer2_outputs[1608] = 1'b1;
    assign layer2_outputs[1609] = ~(layer1_outputs[2307]) | (layer1_outputs[1605]);
    assign layer2_outputs[1610] = (layer1_outputs[1574]) & ~(layer1_outputs[1345]);
    assign layer2_outputs[1611] = (layer1_outputs[2154]) & ~(layer1_outputs[623]);
    assign layer2_outputs[1612] = layer1_outputs[1403];
    assign layer2_outputs[1613] = ~(layer1_outputs[1476]);
    assign layer2_outputs[1614] = ~(layer1_outputs[679]);
    assign layer2_outputs[1615] = (layer1_outputs[1522]) & ~(layer1_outputs[893]);
    assign layer2_outputs[1616] = ~(layer1_outputs[339]) | (layer1_outputs[1036]);
    assign layer2_outputs[1617] = ~((layer1_outputs[2101]) ^ (layer1_outputs[141]));
    assign layer2_outputs[1618] = ~(layer1_outputs[550]);
    assign layer2_outputs[1619] = 1'b1;
    assign layer2_outputs[1620] = layer1_outputs[650];
    assign layer2_outputs[1621] = ~(layer1_outputs[1198]);
    assign layer2_outputs[1622] = ~(layer1_outputs[1604]);
    assign layer2_outputs[1623] = 1'b0;
    assign layer2_outputs[1624] = ~(layer1_outputs[1807]) | (layer1_outputs[241]);
    assign layer2_outputs[1625] = (layer1_outputs[35]) & (layer1_outputs[2312]);
    assign layer2_outputs[1626] = layer1_outputs[934];
    assign layer2_outputs[1627] = (layer1_outputs[2148]) & ~(layer1_outputs[834]);
    assign layer2_outputs[1628] = 1'b0;
    assign layer2_outputs[1629] = (layer1_outputs[247]) & ~(layer1_outputs[1602]);
    assign layer2_outputs[1630] = ~(layer1_outputs[147]);
    assign layer2_outputs[1631] = layer1_outputs[565];
    assign layer2_outputs[1632] = 1'b1;
    assign layer2_outputs[1633] = (layer1_outputs[1160]) & ~(layer1_outputs[2279]);
    assign layer2_outputs[1634] = (layer1_outputs[1382]) & (layer1_outputs[1009]);
    assign layer2_outputs[1635] = (layer1_outputs[1962]) | (layer1_outputs[51]);
    assign layer2_outputs[1636] = layer1_outputs[382];
    assign layer2_outputs[1637] = ~((layer1_outputs[1597]) & (layer1_outputs[126]));
    assign layer2_outputs[1638] = layer1_outputs[484];
    assign layer2_outputs[1639] = (layer1_outputs[1657]) & ~(layer1_outputs[1064]);
    assign layer2_outputs[1640] = 1'b0;
    assign layer2_outputs[1641] = ~((layer1_outputs[2304]) | (layer1_outputs[922]));
    assign layer2_outputs[1642] = (layer1_outputs[1983]) & ~(layer1_outputs[1501]);
    assign layer2_outputs[1643] = ~(layer1_outputs[2248]);
    assign layer2_outputs[1644] = ~((layer1_outputs[1873]) ^ (layer1_outputs[181]));
    assign layer2_outputs[1645] = layer1_outputs[773];
    assign layer2_outputs[1646] = (layer1_outputs[794]) & ~(layer1_outputs[1895]);
    assign layer2_outputs[1647] = ~((layer1_outputs[1745]) & (layer1_outputs[2056]));
    assign layer2_outputs[1648] = ~(layer1_outputs[709]);
    assign layer2_outputs[1649] = (layer1_outputs[1389]) & ~(layer1_outputs[2507]);
    assign layer2_outputs[1650] = layer1_outputs[1581];
    assign layer2_outputs[1651] = layer1_outputs[57];
    assign layer2_outputs[1652] = (layer1_outputs[1002]) & ~(layer1_outputs[2447]);
    assign layer2_outputs[1653] = (layer1_outputs[1700]) & (layer1_outputs[2296]);
    assign layer2_outputs[1654] = (layer1_outputs[1648]) & ~(layer1_outputs[2027]);
    assign layer2_outputs[1655] = (layer1_outputs[1254]) & (layer1_outputs[186]);
    assign layer2_outputs[1656] = ~((layer1_outputs[419]) | (layer1_outputs[391]));
    assign layer2_outputs[1657] = layer1_outputs[146];
    assign layer2_outputs[1658] = 1'b1;
    assign layer2_outputs[1659] = ~((layer1_outputs[2476]) & (layer1_outputs[972]));
    assign layer2_outputs[1660] = layer1_outputs[2191];
    assign layer2_outputs[1661] = ~(layer1_outputs[2426]);
    assign layer2_outputs[1662] = (layer1_outputs[86]) | (layer1_outputs[79]);
    assign layer2_outputs[1663] = layer1_outputs[341];
    assign layer2_outputs[1664] = 1'b0;
    assign layer2_outputs[1665] = ~(layer1_outputs[605]) | (layer1_outputs[1416]);
    assign layer2_outputs[1666] = ~(layer1_outputs[2348]) | (layer1_outputs[34]);
    assign layer2_outputs[1667] = ~(layer1_outputs[2395]) | (layer1_outputs[19]);
    assign layer2_outputs[1668] = ~(layer1_outputs[674]);
    assign layer2_outputs[1669] = ~(layer1_outputs[1487]);
    assign layer2_outputs[1670] = (layer1_outputs[1946]) & ~(layer1_outputs[786]);
    assign layer2_outputs[1671] = ~(layer1_outputs[1253]);
    assign layer2_outputs[1672] = ~((layer1_outputs[1652]) ^ (layer1_outputs[281]));
    assign layer2_outputs[1673] = ~(layer1_outputs[528]);
    assign layer2_outputs[1674] = ~(layer1_outputs[1293]);
    assign layer2_outputs[1675] = ~(layer1_outputs[1241]);
    assign layer2_outputs[1676] = ~(layer1_outputs[626]) | (layer1_outputs[2075]);
    assign layer2_outputs[1677] = (layer1_outputs[2476]) & ~(layer1_outputs[1621]);
    assign layer2_outputs[1678] = ~(layer1_outputs[197]);
    assign layer2_outputs[1679] = layer1_outputs[885];
    assign layer2_outputs[1680] = (layer1_outputs[1074]) & ~(layer1_outputs[1616]);
    assign layer2_outputs[1681] = ~(layer1_outputs[317]) | (layer1_outputs[1695]);
    assign layer2_outputs[1682] = ~((layer1_outputs[2418]) | (layer1_outputs[1945]));
    assign layer2_outputs[1683] = ~((layer1_outputs[1769]) | (layer1_outputs[2021]));
    assign layer2_outputs[1684] = 1'b1;
    assign layer2_outputs[1685] = (layer1_outputs[1832]) & ~(layer1_outputs[2542]);
    assign layer2_outputs[1686] = ~((layer1_outputs[522]) & (layer1_outputs[2333]));
    assign layer2_outputs[1687] = ~(layer1_outputs[941]);
    assign layer2_outputs[1688] = layer1_outputs[936];
    assign layer2_outputs[1689] = layer1_outputs[1939];
    assign layer2_outputs[1690] = (layer1_outputs[1599]) ^ (layer1_outputs[41]);
    assign layer2_outputs[1691] = layer1_outputs[1997];
    assign layer2_outputs[1692] = (layer1_outputs[318]) ^ (layer1_outputs[2388]);
    assign layer2_outputs[1693] = layer1_outputs[353];
    assign layer2_outputs[1694] = ~((layer1_outputs[472]) & (layer1_outputs[525]));
    assign layer2_outputs[1695] = (layer1_outputs[1700]) & ~(layer1_outputs[1448]);
    assign layer2_outputs[1696] = ~((layer1_outputs[1600]) & (layer1_outputs[2051]));
    assign layer2_outputs[1697] = ~(layer1_outputs[1193]) | (layer1_outputs[946]);
    assign layer2_outputs[1698] = ~((layer1_outputs[2326]) | (layer1_outputs[2396]));
    assign layer2_outputs[1699] = ~(layer1_outputs[1069]);
    assign layer2_outputs[1700] = layer1_outputs[1306];
    assign layer2_outputs[1701] = layer1_outputs[221];
    assign layer2_outputs[1702] = layer1_outputs[1070];
    assign layer2_outputs[1703] = ~(layer1_outputs[1410]) | (layer1_outputs[638]);
    assign layer2_outputs[1704] = (layer1_outputs[2039]) & ~(layer1_outputs[132]);
    assign layer2_outputs[1705] = ~((layer1_outputs[293]) | (layer1_outputs[190]));
    assign layer2_outputs[1706] = layer1_outputs[2266];
    assign layer2_outputs[1707] = ~(layer1_outputs[1237]) | (layer1_outputs[1334]);
    assign layer2_outputs[1708] = ~(layer1_outputs[481]) | (layer1_outputs[1462]);
    assign layer2_outputs[1709] = layer1_outputs[219];
    assign layer2_outputs[1710] = ~((layer1_outputs[1072]) ^ (layer1_outputs[1414]));
    assign layer2_outputs[1711] = (layer1_outputs[1513]) & ~(layer1_outputs[2047]);
    assign layer2_outputs[1712] = 1'b0;
    assign layer2_outputs[1713] = ~(layer1_outputs[883]);
    assign layer2_outputs[1714] = ~(layer1_outputs[374]) | (layer1_outputs[1366]);
    assign layer2_outputs[1715] = ~(layer1_outputs[960]) | (layer1_outputs[1035]);
    assign layer2_outputs[1716] = ~((layer1_outputs[212]) & (layer1_outputs[671]));
    assign layer2_outputs[1717] = ~((layer1_outputs[2273]) & (layer1_outputs[2155]));
    assign layer2_outputs[1718] = ~(layer1_outputs[450]) | (layer1_outputs[360]);
    assign layer2_outputs[1719] = ~(layer1_outputs[723]);
    assign layer2_outputs[1720] = ~(layer1_outputs[2539]) | (layer1_outputs[2462]);
    assign layer2_outputs[1721] = 1'b1;
    assign layer2_outputs[1722] = ~((layer1_outputs[2297]) | (layer1_outputs[1393]));
    assign layer2_outputs[1723] = (layer1_outputs[288]) ^ (layer1_outputs[814]);
    assign layer2_outputs[1724] = ~(layer1_outputs[1171]) | (layer1_outputs[54]);
    assign layer2_outputs[1725] = (layer1_outputs[1726]) & ~(layer1_outputs[940]);
    assign layer2_outputs[1726] = ~(layer1_outputs[146]);
    assign layer2_outputs[1727] = ~((layer1_outputs[503]) ^ (layer1_outputs[275]));
    assign layer2_outputs[1728] = ~(layer1_outputs[192]) | (layer1_outputs[1947]);
    assign layer2_outputs[1729] = 1'b1;
    assign layer2_outputs[1730] = (layer1_outputs[2320]) | (layer1_outputs[1646]);
    assign layer2_outputs[1731] = (layer1_outputs[799]) & ~(layer1_outputs[295]);
    assign layer2_outputs[1732] = (layer1_outputs[245]) & ~(layer1_outputs[1771]);
    assign layer2_outputs[1733] = ~((layer1_outputs[490]) | (layer1_outputs[818]));
    assign layer2_outputs[1734] = ~(layer1_outputs[1142]) | (layer1_outputs[1400]);
    assign layer2_outputs[1735] = layer1_outputs[1110];
    assign layer2_outputs[1736] = (layer1_outputs[408]) & (layer1_outputs[1768]);
    assign layer2_outputs[1737] = (layer1_outputs[2408]) & (layer1_outputs[1915]);
    assign layer2_outputs[1738] = layer1_outputs[1365];
    assign layer2_outputs[1739] = ~(layer1_outputs[600]);
    assign layer2_outputs[1740] = ~(layer1_outputs[473]);
    assign layer2_outputs[1741] = (layer1_outputs[637]) | (layer1_outputs[807]);
    assign layer2_outputs[1742] = layer1_outputs[1096];
    assign layer2_outputs[1743] = layer1_outputs[1511];
    assign layer2_outputs[1744] = ~(layer1_outputs[926]);
    assign layer2_outputs[1745] = layer1_outputs[1749];
    assign layer2_outputs[1746] = ~((layer1_outputs[2063]) | (layer1_outputs[2452]));
    assign layer2_outputs[1747] = ~((layer1_outputs[978]) & (layer1_outputs[1620]));
    assign layer2_outputs[1748] = ~(layer1_outputs[1322]);
    assign layer2_outputs[1749] = (layer1_outputs[130]) & ~(layer1_outputs[1621]);
    assign layer2_outputs[1750] = layer1_outputs[1229];
    assign layer2_outputs[1751] = layer1_outputs[980];
    assign layer2_outputs[1752] = (layer1_outputs[1060]) ^ (layer1_outputs[1062]);
    assign layer2_outputs[1753] = ~(layer1_outputs[2390]);
    assign layer2_outputs[1754] = 1'b0;
    assign layer2_outputs[1755] = ~((layer1_outputs[819]) & (layer1_outputs[1665]));
    assign layer2_outputs[1756] = ~(layer1_outputs[1189]);
    assign layer2_outputs[1757] = ~(layer1_outputs[1019]);
    assign layer2_outputs[1758] = (layer1_outputs[2069]) & (layer1_outputs[2293]);
    assign layer2_outputs[1759] = ~((layer1_outputs[165]) & (layer1_outputs[542]));
    assign layer2_outputs[1760] = ~((layer1_outputs[800]) & (layer1_outputs[717]));
    assign layer2_outputs[1761] = ~(layer1_outputs[1251]);
    assign layer2_outputs[1762] = (layer1_outputs[1458]) & ~(layer1_outputs[373]);
    assign layer2_outputs[1763] = ~((layer1_outputs[535]) ^ (layer1_outputs[700]));
    assign layer2_outputs[1764] = layer1_outputs[2316];
    assign layer2_outputs[1765] = layer1_outputs[1905];
    assign layer2_outputs[1766] = ~(layer1_outputs[2172]);
    assign layer2_outputs[1767] = ~(layer1_outputs[1523]) | (layer1_outputs[833]);
    assign layer2_outputs[1768] = (layer1_outputs[1724]) & ~(layer1_outputs[1153]);
    assign layer2_outputs[1769] = (layer1_outputs[374]) & ~(layer1_outputs[117]);
    assign layer2_outputs[1770] = 1'b1;
    assign layer2_outputs[1771] = ~(layer1_outputs[1060]);
    assign layer2_outputs[1772] = layer1_outputs[1948];
    assign layer2_outputs[1773] = layer1_outputs[461];
    assign layer2_outputs[1774] = (layer1_outputs[1978]) & (layer1_outputs[1771]);
    assign layer2_outputs[1775] = layer1_outputs[1653];
    assign layer2_outputs[1776] = ~(layer1_outputs[2080]) | (layer1_outputs[253]);
    assign layer2_outputs[1777] = (layer1_outputs[1547]) & ~(layer1_outputs[1982]);
    assign layer2_outputs[1778] = (layer1_outputs[1317]) & (layer1_outputs[1018]);
    assign layer2_outputs[1779] = ~((layer1_outputs[2272]) & (layer1_outputs[588]));
    assign layer2_outputs[1780] = (layer1_outputs[1008]) & ~(layer1_outputs[1234]);
    assign layer2_outputs[1781] = ~(layer1_outputs[752]);
    assign layer2_outputs[1782] = (layer1_outputs[343]) | (layer1_outputs[710]);
    assign layer2_outputs[1783] = (layer1_outputs[1972]) ^ (layer1_outputs[1478]);
    assign layer2_outputs[1784] = layer1_outputs[1793];
    assign layer2_outputs[1785] = (layer1_outputs[896]) & ~(layer1_outputs[924]);
    assign layer2_outputs[1786] = (layer1_outputs[1360]) & ~(layer1_outputs[203]);
    assign layer2_outputs[1787] = layer1_outputs[271];
    assign layer2_outputs[1788] = (layer1_outputs[2283]) & ~(layer1_outputs[2329]);
    assign layer2_outputs[1789] = ~(layer1_outputs[1157]);
    assign layer2_outputs[1790] = (layer1_outputs[260]) | (layer1_outputs[1420]);
    assign layer2_outputs[1791] = ~((layer1_outputs[66]) & (layer1_outputs[687]));
    assign layer2_outputs[1792] = (layer1_outputs[1014]) & (layer1_outputs[323]);
    assign layer2_outputs[1793] = (layer1_outputs[1707]) | (layer1_outputs[2307]);
    assign layer2_outputs[1794] = 1'b1;
    assign layer2_outputs[1795] = 1'b1;
    assign layer2_outputs[1796] = ~(layer1_outputs[697]);
    assign layer2_outputs[1797] = ~(layer1_outputs[227]);
    assign layer2_outputs[1798] = ~(layer1_outputs[875]);
    assign layer2_outputs[1799] = layer1_outputs[919];
    assign layer2_outputs[1800] = (layer1_outputs[2315]) & ~(layer1_outputs[2206]);
    assign layer2_outputs[1801] = ~(layer1_outputs[1871]);
    assign layer2_outputs[1802] = ~((layer1_outputs[2396]) | (layer1_outputs[670]));
    assign layer2_outputs[1803] = ~(layer1_outputs[2247]) | (layer1_outputs[317]);
    assign layer2_outputs[1804] = layer1_outputs[291];
    assign layer2_outputs[1805] = 1'b0;
    assign layer2_outputs[1806] = layer1_outputs[619];
    assign layer2_outputs[1807] = 1'b0;
    assign layer2_outputs[1808] = layer1_outputs[1];
    assign layer2_outputs[1809] = ~(layer1_outputs[751]);
    assign layer2_outputs[1810] = 1'b0;
    assign layer2_outputs[1811] = ~(layer1_outputs[2105]) | (layer1_outputs[2119]);
    assign layer2_outputs[1812] = ~(layer1_outputs[2463]);
    assign layer2_outputs[1813] = 1'b1;
    assign layer2_outputs[1814] = layer1_outputs[0];
    assign layer2_outputs[1815] = ~((layer1_outputs[419]) | (layer1_outputs[878]));
    assign layer2_outputs[1816] = (layer1_outputs[2411]) & ~(layer1_outputs[1327]);
    assign layer2_outputs[1817] = (layer1_outputs[2148]) & ~(layer1_outputs[1613]);
    assign layer2_outputs[1818] = layer1_outputs[553];
    assign layer2_outputs[1819] = (layer1_outputs[1505]) ^ (layer1_outputs[2495]);
    assign layer2_outputs[1820] = ~(layer1_outputs[776]) | (layer1_outputs[1891]);
    assign layer2_outputs[1821] = ~(layer1_outputs[2213]) | (layer1_outputs[207]);
    assign layer2_outputs[1822] = layer1_outputs[2314];
    assign layer2_outputs[1823] = 1'b1;
    assign layer2_outputs[1824] = layer1_outputs[311];
    assign layer2_outputs[1825] = ~(layer1_outputs[1504]);
    assign layer2_outputs[1826] = layer1_outputs[1299];
    assign layer2_outputs[1827] = (layer1_outputs[1388]) & ~(layer1_outputs[1747]);
    assign layer2_outputs[1828] = layer1_outputs[2087];
    assign layer2_outputs[1829] = ~((layer1_outputs[743]) | (layer1_outputs[1326]));
    assign layer2_outputs[1830] = (layer1_outputs[606]) | (layer1_outputs[975]);
    assign layer2_outputs[1831] = ~((layer1_outputs[234]) & (layer1_outputs[627]));
    assign layer2_outputs[1832] = ~((layer1_outputs[696]) ^ (layer1_outputs[713]));
    assign layer2_outputs[1833] = layer1_outputs[881];
    assign layer2_outputs[1834] = 1'b1;
    assign layer2_outputs[1835] = ~(layer1_outputs[2278]);
    assign layer2_outputs[1836] = (layer1_outputs[1329]) & ~(layer1_outputs[47]);
    assign layer2_outputs[1837] = 1'b1;
    assign layer2_outputs[1838] = ~(layer1_outputs[616]);
    assign layer2_outputs[1839] = (layer1_outputs[1082]) | (layer1_outputs[1922]);
    assign layer2_outputs[1840] = ~(layer1_outputs[1509]);
    assign layer2_outputs[1841] = layer1_outputs[677];
    assign layer2_outputs[1842] = layer1_outputs[54];
    assign layer2_outputs[1843] = layer1_outputs[1875];
    assign layer2_outputs[1844] = layer1_outputs[2230];
    assign layer2_outputs[1845] = layer1_outputs[2553];
    assign layer2_outputs[1846] = ~(layer1_outputs[2394]);
    assign layer2_outputs[1847] = ~(layer1_outputs[1563]) | (layer1_outputs[1272]);
    assign layer2_outputs[1848] = ~(layer1_outputs[1443]);
    assign layer2_outputs[1849] = ~(layer1_outputs[81]);
    assign layer2_outputs[1850] = ~(layer1_outputs[282]) | (layer1_outputs[604]);
    assign layer2_outputs[1851] = (layer1_outputs[1201]) & (layer1_outputs[231]);
    assign layer2_outputs[1852] = layer1_outputs[2392];
    assign layer2_outputs[1853] = ~(layer1_outputs[2440]);
    assign layer2_outputs[1854] = ~(layer1_outputs[295]) | (layer1_outputs[1462]);
    assign layer2_outputs[1855] = ~((layer1_outputs[204]) | (layer1_outputs[2126]));
    assign layer2_outputs[1856] = ~((layer1_outputs[2432]) | (layer1_outputs[1999]));
    assign layer2_outputs[1857] = ~(layer1_outputs[490]) | (layer1_outputs[1506]);
    assign layer2_outputs[1858] = (layer1_outputs[476]) | (layer1_outputs[2466]);
    assign layer2_outputs[1859] = ~(layer1_outputs[2264]) | (layer1_outputs[1802]);
    assign layer2_outputs[1860] = ~(layer1_outputs[972]) | (layer1_outputs[139]);
    assign layer2_outputs[1861] = ~((layer1_outputs[2211]) & (layer1_outputs[823]));
    assign layer2_outputs[1862] = ~(layer1_outputs[1563]);
    assign layer2_outputs[1863] = 1'b0;
    assign layer2_outputs[1864] = ~(layer1_outputs[388]);
    assign layer2_outputs[1865] = (layer1_outputs[1273]) | (layer1_outputs[2518]);
    assign layer2_outputs[1866] = ~((layer1_outputs[1863]) ^ (layer1_outputs[1456]));
    assign layer2_outputs[1867] = ~((layer1_outputs[1562]) | (layer1_outputs[918]));
    assign layer2_outputs[1868] = layer1_outputs[447];
    assign layer2_outputs[1869] = ~((layer1_outputs[1343]) & (layer1_outputs[82]));
    assign layer2_outputs[1870] = ~(layer1_outputs[85]) | (layer1_outputs[1091]);
    assign layer2_outputs[1871] = 1'b1;
    assign layer2_outputs[1872] = layer1_outputs[1679];
    assign layer2_outputs[1873] = ~((layer1_outputs[1790]) | (layer1_outputs[205]));
    assign layer2_outputs[1874] = (layer1_outputs[733]) ^ (layer1_outputs[2373]);
    assign layer2_outputs[1875] = 1'b1;
    assign layer2_outputs[1876] = ~(layer1_outputs[1490]);
    assign layer2_outputs[1877] = ~(layer1_outputs[2364]) | (layer1_outputs[1721]);
    assign layer2_outputs[1878] = ~(layer1_outputs[2531]);
    assign layer2_outputs[1879] = (layer1_outputs[100]) | (layer1_outputs[544]);
    assign layer2_outputs[1880] = ~(layer1_outputs[916]);
    assign layer2_outputs[1881] = ~(layer1_outputs[1933]);
    assign layer2_outputs[1882] = ~(layer1_outputs[1717]);
    assign layer2_outputs[1883] = ~(layer1_outputs[369]);
    assign layer2_outputs[1884] = layer1_outputs[1656];
    assign layer2_outputs[1885] = layer1_outputs[2548];
    assign layer2_outputs[1886] = (layer1_outputs[305]) | (layer1_outputs[2294]);
    assign layer2_outputs[1887] = ~(layer1_outputs[1886]) | (layer1_outputs[369]);
    assign layer2_outputs[1888] = ~(layer1_outputs[2559]) | (layer1_outputs[2062]);
    assign layer2_outputs[1889] = (layer1_outputs[951]) ^ (layer1_outputs[2555]);
    assign layer2_outputs[1890] = ~(layer1_outputs[943]);
    assign layer2_outputs[1891] = layer1_outputs[1439];
    assign layer2_outputs[1892] = ~(layer1_outputs[1421]);
    assign layer2_outputs[1893] = ~((layer1_outputs[936]) | (layer1_outputs[2524]));
    assign layer2_outputs[1894] = ~((layer1_outputs[1860]) ^ (layer1_outputs[1660]));
    assign layer2_outputs[1895] = ~((layer1_outputs[757]) ^ (layer1_outputs[2299]));
    assign layer2_outputs[1896] = layer1_outputs[1480];
    assign layer2_outputs[1897] = (layer1_outputs[2479]) ^ (layer1_outputs[583]);
    assign layer2_outputs[1898] = ~(layer1_outputs[118]) | (layer1_outputs[965]);
    assign layer2_outputs[1899] = layer1_outputs[1299];
    assign layer2_outputs[1900] = layer1_outputs[529];
    assign layer2_outputs[1901] = ~(layer1_outputs[1836]);
    assign layer2_outputs[1902] = layer1_outputs[1869];
    assign layer2_outputs[1903] = layer1_outputs[1401];
    assign layer2_outputs[1904] = layer1_outputs[1976];
    assign layer2_outputs[1905] = layer1_outputs[503];
    assign layer2_outputs[1906] = (layer1_outputs[1494]) & ~(layer1_outputs[505]);
    assign layer2_outputs[1907] = ~((layer1_outputs[1194]) ^ (layer1_outputs[1058]));
    assign layer2_outputs[1908] = layer1_outputs[1301];
    assign layer2_outputs[1909] = layer1_outputs[159];
    assign layer2_outputs[1910] = ~((layer1_outputs[1162]) | (layer1_outputs[702]));
    assign layer2_outputs[1911] = ~(layer1_outputs[267]) | (layer1_outputs[2011]);
    assign layer2_outputs[1912] = layer1_outputs[301];
    assign layer2_outputs[1913] = ~(layer1_outputs[73]) | (layer1_outputs[1977]);
    assign layer2_outputs[1914] = 1'b0;
    assign layer2_outputs[1915] = (layer1_outputs[283]) & ~(layer1_outputs[1943]);
    assign layer2_outputs[1916] = layer1_outputs[2088];
    assign layer2_outputs[1917] = ~(layer1_outputs[1255]);
    assign layer2_outputs[1918] = 1'b0;
    assign layer2_outputs[1919] = layer1_outputs[1468];
    assign layer2_outputs[1920] = ~((layer1_outputs[2008]) & (layer1_outputs[1428]));
    assign layer2_outputs[1921] = (layer1_outputs[1544]) & ~(layer1_outputs[26]);
    assign layer2_outputs[1922] = ~(layer1_outputs[916]);
    assign layer2_outputs[1923] = ~(layer1_outputs[2040]) | (layer1_outputs[561]);
    assign layer2_outputs[1924] = layer1_outputs[1148];
    assign layer2_outputs[1925] = (layer1_outputs[1882]) & ~(layer1_outputs[211]);
    assign layer2_outputs[1926] = ~(layer1_outputs[2325]);
    assign layer2_outputs[1927] = ~(layer1_outputs[1678]) | (layer1_outputs[1357]);
    assign layer2_outputs[1928] = ~(layer1_outputs[770]);
    assign layer2_outputs[1929] = ~(layer1_outputs[1496]) | (layer1_outputs[748]);
    assign layer2_outputs[1930] = (layer1_outputs[1430]) & (layer1_outputs[1761]);
    assign layer2_outputs[1931] = layer1_outputs[2170];
    assign layer2_outputs[1932] = ~((layer1_outputs[2505]) ^ (layer1_outputs[1453]));
    assign layer2_outputs[1933] = (layer1_outputs[2212]) | (layer1_outputs[1421]);
    assign layer2_outputs[1934] = ~(layer1_outputs[874]) | (layer1_outputs[1583]);
    assign layer2_outputs[1935] = ~(layer1_outputs[155]);
    assign layer2_outputs[1936] = (layer1_outputs[1983]) & (layer1_outputs[1243]);
    assign layer2_outputs[1937] = layer1_outputs[2317];
    assign layer2_outputs[1938] = layer1_outputs[1876];
    assign layer2_outputs[1939] = ~(layer1_outputs[1064]);
    assign layer2_outputs[1940] = 1'b0;
    assign layer2_outputs[1941] = layer1_outputs[690];
    assign layer2_outputs[1942] = layer1_outputs[857];
    assign layer2_outputs[1943] = ~(layer1_outputs[1991]);
    assign layer2_outputs[1944] = (layer1_outputs[2315]) & (layer1_outputs[2091]);
    assign layer2_outputs[1945] = (layer1_outputs[850]) & ~(layer1_outputs[1913]);
    assign layer2_outputs[1946] = (layer1_outputs[344]) & ~(layer1_outputs[1595]);
    assign layer2_outputs[1947] = 1'b0;
    assign layer2_outputs[1948] = ~(layer1_outputs[421]);
    assign layer2_outputs[1949] = ~((layer1_outputs[1434]) ^ (layer1_outputs[1944]));
    assign layer2_outputs[1950] = ~(layer1_outputs[397]) | (layer1_outputs[2460]);
    assign layer2_outputs[1951] = layer1_outputs[2434];
    assign layer2_outputs[1952] = ~(layer1_outputs[1132]);
    assign layer2_outputs[1953] = ~(layer1_outputs[830]);
    assign layer2_outputs[1954] = ~(layer1_outputs[2453]);
    assign layer2_outputs[1955] = (layer1_outputs[2110]) & ~(layer1_outputs[798]);
    assign layer2_outputs[1956] = (layer1_outputs[1510]) & ~(layer1_outputs[2107]);
    assign layer2_outputs[1957] = ~((layer1_outputs[1346]) | (layer1_outputs[2331]));
    assign layer2_outputs[1958] = ~(layer1_outputs[636]);
    assign layer2_outputs[1959] = (layer1_outputs[2477]) & (layer1_outputs[1217]);
    assign layer2_outputs[1960] = ~(layer1_outputs[2520]);
    assign layer2_outputs[1961] = (layer1_outputs[1206]) & ~(layer1_outputs[1633]);
    assign layer2_outputs[1962] = ~((layer1_outputs[1425]) | (layer1_outputs[638]));
    assign layer2_outputs[1963] = (layer1_outputs[2544]) & (layer1_outputs[1357]);
    assign layer2_outputs[1964] = ~(layer1_outputs[2042]) | (layer1_outputs[1331]);
    assign layer2_outputs[1965] = layer1_outputs[1901];
    assign layer2_outputs[1966] = (layer1_outputs[1101]) & ~(layer1_outputs[2539]);
    assign layer2_outputs[1967] = layer1_outputs[1436];
    assign layer2_outputs[1968] = 1'b0;
    assign layer2_outputs[1969] = layer1_outputs[718];
    assign layer2_outputs[1970] = ~(layer1_outputs[366]) | (layer1_outputs[385]);
    assign layer2_outputs[1971] = 1'b0;
    assign layer2_outputs[1972] = (layer1_outputs[1566]) & ~(layer1_outputs[1978]);
    assign layer2_outputs[1973] = (layer1_outputs[633]) & ~(layer1_outputs[1308]);
    assign layer2_outputs[1974] = ~((layer1_outputs[806]) & (layer1_outputs[24]));
    assign layer2_outputs[1975] = ~(layer1_outputs[324]);
    assign layer2_outputs[1976] = ~(layer1_outputs[1619]);
    assign layer2_outputs[1977] = ~(layer1_outputs[738]) | (layer1_outputs[1846]);
    assign layer2_outputs[1978] = layer1_outputs[1358];
    assign layer2_outputs[1979] = ~(layer1_outputs[246]);
    assign layer2_outputs[1980] = ~(layer1_outputs[2006]) | (layer1_outputs[1495]);
    assign layer2_outputs[1981] = ~(layer1_outputs[2404]);
    assign layer2_outputs[1982] = (layer1_outputs[1728]) & ~(layer1_outputs[2337]);
    assign layer2_outputs[1983] = ~((layer1_outputs[2377]) | (layer1_outputs[88]));
    assign layer2_outputs[1984] = ~((layer1_outputs[1315]) | (layer1_outputs[1237]));
    assign layer2_outputs[1985] = ~(layer1_outputs[2351]);
    assign layer2_outputs[1986] = 1'b0;
    assign layer2_outputs[1987] = layer1_outputs[94];
    assign layer2_outputs[1988] = ~(layer1_outputs[17]) | (layer1_outputs[280]);
    assign layer2_outputs[1989] = ~((layer1_outputs[403]) & (layer1_outputs[7]));
    assign layer2_outputs[1990] = layer1_outputs[1412];
    assign layer2_outputs[1991] = ~(layer1_outputs[2182]) | (layer1_outputs[1767]);
    assign layer2_outputs[1992] = (layer1_outputs[1547]) & ~(layer1_outputs[1512]);
    assign layer2_outputs[1993] = ~((layer1_outputs[1640]) | (layer1_outputs[349]));
    assign layer2_outputs[1994] = layer1_outputs[969];
    assign layer2_outputs[1995] = 1'b0;
    assign layer2_outputs[1996] = ~((layer1_outputs[1306]) | (layer1_outputs[1406]));
    assign layer2_outputs[1997] = layer1_outputs[692];
    assign layer2_outputs[1998] = layer1_outputs[719];
    assign layer2_outputs[1999] = 1'b1;
    assign layer2_outputs[2000] = (layer1_outputs[946]) | (layer1_outputs[2048]);
    assign layer2_outputs[2001] = (layer1_outputs[61]) & (layer1_outputs[1554]);
    assign layer2_outputs[2002] = ~(layer1_outputs[262]);
    assign layer2_outputs[2003] = ~(layer1_outputs[2145]);
    assign layer2_outputs[2004] = 1'b0;
    assign layer2_outputs[2005] = layer1_outputs[1238];
    assign layer2_outputs[2006] = ~(layer1_outputs[2492]) | (layer1_outputs[846]);
    assign layer2_outputs[2007] = (layer1_outputs[1365]) & ~(layer1_outputs[136]);
    assign layer2_outputs[2008] = layer1_outputs[169];
    assign layer2_outputs[2009] = ~((layer1_outputs[2060]) | (layer1_outputs[2120]));
    assign layer2_outputs[2010] = ~((layer1_outputs[1755]) | (layer1_outputs[394]));
    assign layer2_outputs[2011] = layer1_outputs[170];
    assign layer2_outputs[2012] = 1'b0;
    assign layer2_outputs[2013] = layer1_outputs[384];
    assign layer2_outputs[2014] = layer1_outputs[2225];
    assign layer2_outputs[2015] = ~(layer1_outputs[2054]);
    assign layer2_outputs[2016] = (layer1_outputs[1292]) & (layer1_outputs[2058]);
    assign layer2_outputs[2017] = (layer1_outputs[536]) & ~(layer1_outputs[336]);
    assign layer2_outputs[2018] = layer1_outputs[1804];
    assign layer2_outputs[2019] = layer1_outputs[1350];
    assign layer2_outputs[2020] = (layer1_outputs[952]) & ~(layer1_outputs[2449]);
    assign layer2_outputs[2021] = ~((layer1_outputs[2367]) & (layer1_outputs[399]));
    assign layer2_outputs[2022] = ~(layer1_outputs[1669]);
    assign layer2_outputs[2023] = layer1_outputs[462];
    assign layer2_outputs[2024] = ~(layer1_outputs[1877]);
    assign layer2_outputs[2025] = ~(layer1_outputs[2119]);
    assign layer2_outputs[2026] = ~((layer1_outputs[1665]) & (layer1_outputs[746]));
    assign layer2_outputs[2027] = ~(layer1_outputs[138]);
    assign layer2_outputs[2028] = ~(layer1_outputs[1450]);
    assign layer2_outputs[2029] = layer1_outputs[1249];
    assign layer2_outputs[2030] = 1'b0;
    assign layer2_outputs[2031] = (layer1_outputs[1581]) & (layer1_outputs[996]);
    assign layer2_outputs[2032] = (layer1_outputs[1159]) ^ (layer1_outputs[528]);
    assign layer2_outputs[2033] = 1'b0;
    assign layer2_outputs[2034] = layer1_outputs[768];
    assign layer2_outputs[2035] = layer1_outputs[1323];
    assign layer2_outputs[2036] = ~(layer1_outputs[2513]);
    assign layer2_outputs[2037] = ~(layer1_outputs[38]);
    assign layer2_outputs[2038] = ~(layer1_outputs[930]);
    assign layer2_outputs[2039] = (layer1_outputs[328]) & ~(layer1_outputs[728]);
    assign layer2_outputs[2040] = ~(layer1_outputs[1451]);
    assign layer2_outputs[2041] = layer1_outputs[1437];
    assign layer2_outputs[2042] = 1'b1;
    assign layer2_outputs[2043] = 1'b0;
    assign layer2_outputs[2044] = ~((layer1_outputs[527]) | (layer1_outputs[1339]));
    assign layer2_outputs[2045] = ~(layer1_outputs[330]);
    assign layer2_outputs[2046] = layer1_outputs[61];
    assign layer2_outputs[2047] = ~((layer1_outputs[1948]) & (layer1_outputs[1303]));
    assign layer2_outputs[2048] = (layer1_outputs[484]) & (layer1_outputs[1524]);
    assign layer2_outputs[2049] = layer1_outputs[515];
    assign layer2_outputs[2050] = ~(layer1_outputs[1020]);
    assign layer2_outputs[2051] = 1'b0;
    assign layer2_outputs[2052] = ~(layer1_outputs[2127]);
    assign layer2_outputs[2053] = ~(layer1_outputs[2032]) | (layer1_outputs[308]);
    assign layer2_outputs[2054] = 1'b0;
    assign layer2_outputs[2055] = (layer1_outputs[2527]) & ~(layer1_outputs[452]);
    assign layer2_outputs[2056] = ~(layer1_outputs[2481]);
    assign layer2_outputs[2057] = ~(layer1_outputs[1353]);
    assign layer2_outputs[2058] = layer1_outputs[1675];
    assign layer2_outputs[2059] = ~((layer1_outputs[581]) & (layer1_outputs[1602]));
    assign layer2_outputs[2060] = layer1_outputs[432];
    assign layer2_outputs[2061] = ~(layer1_outputs[873]) | (layer1_outputs[289]);
    assign layer2_outputs[2062] = layer1_outputs[1637];
    assign layer2_outputs[2063] = ~(layer1_outputs[1282]);
    assign layer2_outputs[2064] = (layer1_outputs[1286]) | (layer1_outputs[333]);
    assign layer2_outputs[2065] = ~(layer1_outputs[887]);
    assign layer2_outputs[2066] = ~(layer1_outputs[1232]) | (layer1_outputs[1182]);
    assign layer2_outputs[2067] = ~((layer1_outputs[1405]) | (layer1_outputs[761]));
    assign layer2_outputs[2068] = ~(layer1_outputs[361]);
    assign layer2_outputs[2069] = (layer1_outputs[315]) & ~(layer1_outputs[1617]);
    assign layer2_outputs[2070] = (layer1_outputs[999]) & ~(layer1_outputs[1861]);
    assign layer2_outputs[2071] = 1'b1;
    assign layer2_outputs[2072] = ~(layer1_outputs[1630]);
    assign layer2_outputs[2073] = layer1_outputs[876];
    assign layer2_outputs[2074] = ~(layer1_outputs[452]);
    assign layer2_outputs[2075] = 1'b0;
    assign layer2_outputs[2076] = (layer1_outputs[106]) ^ (layer1_outputs[392]);
    assign layer2_outputs[2077] = (layer1_outputs[357]) | (layer1_outputs[485]);
    assign layer2_outputs[2078] = ~(layer1_outputs[191]) | (layer1_outputs[2475]);
    assign layer2_outputs[2079] = 1'b0;
    assign layer2_outputs[2080] = ~(layer1_outputs[1964]) | (layer1_outputs[264]);
    assign layer2_outputs[2081] = ~(layer1_outputs[601]);
    assign layer2_outputs[2082] = ~((layer1_outputs[1755]) | (layer1_outputs[1540]));
    assign layer2_outputs[2083] = 1'b0;
    assign layer2_outputs[2084] = (layer1_outputs[1387]) | (layer1_outputs[1733]);
    assign layer2_outputs[2085] = layer1_outputs[375];
    assign layer2_outputs[2086] = ~(layer1_outputs[1176]);
    assign layer2_outputs[2087] = (layer1_outputs[2493]) | (layer1_outputs[1318]);
    assign layer2_outputs[2088] = ~((layer1_outputs[1973]) & (layer1_outputs[1394]));
    assign layer2_outputs[2089] = ~(layer1_outputs[1822]);
    assign layer2_outputs[2090] = ~(layer1_outputs[1677]);
    assign layer2_outputs[2091] = 1'b0;
    assign layer2_outputs[2092] = (layer1_outputs[383]) & ~(layer1_outputs[992]);
    assign layer2_outputs[2093] = ~(layer1_outputs[119]);
    assign layer2_outputs[2094] = ~(layer1_outputs[1605]);
    assign layer2_outputs[2095] = layer1_outputs[513];
    assign layer2_outputs[2096] = 1'b0;
    assign layer2_outputs[2097] = (layer1_outputs[75]) | (layer1_outputs[2436]);
    assign layer2_outputs[2098] = ~((layer1_outputs[1591]) & (layer1_outputs[1924]));
    assign layer2_outputs[2099] = (layer1_outputs[1772]) & ~(layer1_outputs[858]);
    assign layer2_outputs[2100] = 1'b0;
    assign layer2_outputs[2101] = (layer1_outputs[1519]) & (layer1_outputs[1996]);
    assign layer2_outputs[2102] = ~(layer1_outputs[443]);
    assign layer2_outputs[2103] = (layer1_outputs[2457]) & ~(layer1_outputs[2201]);
    assign layer2_outputs[2104] = layer1_outputs[2441];
    assign layer2_outputs[2105] = (layer1_outputs[851]) & (layer1_outputs[1019]);
    assign layer2_outputs[2106] = (layer1_outputs[1499]) | (layer1_outputs[2545]);
    assign layer2_outputs[2107] = layer1_outputs[1164];
    assign layer2_outputs[2108] = (layer1_outputs[476]) | (layer1_outputs[1125]);
    assign layer2_outputs[2109] = ~(layer1_outputs[644]) | (layer1_outputs[78]);
    assign layer2_outputs[2110] = (layer1_outputs[1652]) | (layer1_outputs[2479]);
    assign layer2_outputs[2111] = (layer1_outputs[102]) & (layer1_outputs[716]);
    assign layer2_outputs[2112] = (layer1_outputs[2213]) & ~(layer1_outputs[2037]);
    assign layer2_outputs[2113] = layer1_outputs[520];
    assign layer2_outputs[2114] = (layer1_outputs[2276]) & ~(layer1_outputs[1117]);
    assign layer2_outputs[2115] = ~(layer1_outputs[469]) | (layer1_outputs[1989]);
    assign layer2_outputs[2116] = 1'b0;
    assign layer2_outputs[2117] = layer1_outputs[2441];
    assign layer2_outputs[2118] = ~((layer1_outputs[2230]) | (layer1_outputs[2150]));
    assign layer2_outputs[2119] = (layer1_outputs[1803]) & ~(layer1_outputs[1817]);
    assign layer2_outputs[2120] = (layer1_outputs[1701]) & (layer1_outputs[937]);
    assign layer2_outputs[2121] = ~((layer1_outputs[1349]) & (layer1_outputs[1461]));
    assign layer2_outputs[2122] = ~(layer1_outputs[1375]) | (layer1_outputs[671]);
    assign layer2_outputs[2123] = layer1_outputs[48];
    assign layer2_outputs[2124] = ~(layer1_outputs[1805]);
    assign layer2_outputs[2125] = (layer1_outputs[500]) | (layer1_outputs[121]);
    assign layer2_outputs[2126] = ~(layer1_outputs[898]);
    assign layer2_outputs[2127] = ~(layer1_outputs[839]) | (layer1_outputs[250]);
    assign layer2_outputs[2128] = ~((layer1_outputs[2436]) ^ (layer1_outputs[2366]));
    assign layer2_outputs[2129] = ~((layer1_outputs[2286]) & (layer1_outputs[2087]));
    assign layer2_outputs[2130] = ~((layer1_outputs[1269]) ^ (layer1_outputs[2524]));
    assign layer2_outputs[2131] = (layer1_outputs[2105]) & ~(layer1_outputs[825]);
    assign layer2_outputs[2132] = (layer1_outputs[693]) & (layer1_outputs[624]);
    assign layer2_outputs[2133] = ~((layer1_outputs[431]) & (layer1_outputs[1097]));
    assign layer2_outputs[2134] = layer1_outputs[1688];
    assign layer2_outputs[2135] = (layer1_outputs[1908]) & (layer1_outputs[1706]);
    assign layer2_outputs[2136] = ~(layer1_outputs[2318]) | (layer1_outputs[137]);
    assign layer2_outputs[2137] = 1'b0;
    assign layer2_outputs[2138] = (layer1_outputs[1325]) & ~(layer1_outputs[268]);
    assign layer2_outputs[2139] = (layer1_outputs[2005]) & ~(layer1_outputs[1133]);
    assign layer2_outputs[2140] = ~(layer1_outputs[1739]) | (layer1_outputs[2464]);
    assign layer2_outputs[2141] = (layer1_outputs[587]) & ~(layer1_outputs[678]);
    assign layer2_outputs[2142] = (layer1_outputs[2097]) & ~(layer1_outputs[676]);
    assign layer2_outputs[2143] = ~(layer1_outputs[276]);
    assign layer2_outputs[2144] = ~(layer1_outputs[179]) | (layer1_outputs[1743]);
    assign layer2_outputs[2145] = layer1_outputs[168];
    assign layer2_outputs[2146] = (layer1_outputs[744]) & ~(layer1_outputs[1455]);
    assign layer2_outputs[2147] = ~(layer1_outputs[927]) | (layer1_outputs[2196]);
    assign layer2_outputs[2148] = ~((layer1_outputs[1033]) | (layer1_outputs[1296]));
    assign layer2_outputs[2149] = (layer1_outputs[621]) & ~(layer1_outputs[1529]);
    assign layer2_outputs[2150] = layer1_outputs[1923];
    assign layer2_outputs[2151] = ~(layer1_outputs[363]);
    assign layer2_outputs[2152] = layer1_outputs[772];
    assign layer2_outputs[2153] = ~(layer1_outputs[1932]) | (layer1_outputs[792]);
    assign layer2_outputs[2154] = ~(layer1_outputs[2346]);
    assign layer2_outputs[2155] = ~(layer1_outputs[1485]) | (layer1_outputs[1163]);
    assign layer2_outputs[2156] = (layer1_outputs[1228]) ^ (layer1_outputs[2166]);
    assign layer2_outputs[2157] = ~(layer1_outputs[2400]);
    assign layer2_outputs[2158] = layer1_outputs[558];
    assign layer2_outputs[2159] = ~(layer1_outputs[1574]) | (layer1_outputs[2011]);
    assign layer2_outputs[2160] = ~((layer1_outputs[1557]) | (layer1_outputs[494]));
    assign layer2_outputs[2161] = layer1_outputs[932];
    assign layer2_outputs[2162] = 1'b1;
    assign layer2_outputs[2163] = ~(layer1_outputs[658]);
    assign layer2_outputs[2164] = (layer1_outputs[1967]) & ~(layer1_outputs[1632]);
    assign layer2_outputs[2165] = (layer1_outputs[113]) & ~(layer1_outputs[605]);
    assign layer2_outputs[2166] = (layer1_outputs[1587]) ^ (layer1_outputs[835]);
    assign layer2_outputs[2167] = ~(layer1_outputs[1823]);
    assign layer2_outputs[2168] = ~(layer1_outputs[1939]) | (layer1_outputs[2163]);
    assign layer2_outputs[2169] = ~(layer1_outputs[134]);
    assign layer2_outputs[2170] = ~(layer1_outputs[124]) | (layer1_outputs[1834]);
    assign layer2_outputs[2171] = ~(layer1_outputs[1147]);
    assign layer2_outputs[2172] = (layer1_outputs[1121]) & (layer1_outputs[2078]);
    assign layer2_outputs[2173] = (layer1_outputs[422]) & ~(layer1_outputs[1788]);
    assign layer2_outputs[2174] = ~(layer1_outputs[1225]);
    assign layer2_outputs[2175] = (layer1_outputs[1042]) ^ (layer1_outputs[2516]);
    assign layer2_outputs[2176] = ~(layer1_outputs[1031]) | (layer1_outputs[198]);
    assign layer2_outputs[2177] = (layer1_outputs[560]) & ~(layer1_outputs[2304]);
    assign layer2_outputs[2178] = layer1_outputs[1887];
    assign layer2_outputs[2179] = 1'b0;
    assign layer2_outputs[2180] = ~(layer1_outputs[1582]) | (layer1_outputs[1611]);
    assign layer2_outputs[2181] = layer1_outputs[1143];
    assign layer2_outputs[2182] = layer1_outputs[931];
    assign layer2_outputs[2183] = layer1_outputs[764];
    assign layer2_outputs[2184] = ~(layer1_outputs[2022]) | (layer1_outputs[1994]);
    assign layer2_outputs[2185] = ~(layer1_outputs[791]);
    assign layer2_outputs[2186] = layer1_outputs[197];
    assign layer2_outputs[2187] = ~(layer1_outputs[2193]);
    assign layer2_outputs[2188] = ~(layer1_outputs[408]) | (layer1_outputs[1436]);
    assign layer2_outputs[2189] = (layer1_outputs[1634]) & ~(layer1_outputs[2278]);
    assign layer2_outputs[2190] = ~((layer1_outputs[1629]) | (layer1_outputs[2322]));
    assign layer2_outputs[2191] = layer1_outputs[1612];
    assign layer2_outputs[2192] = (layer1_outputs[508]) & (layer1_outputs[520]);
    assign layer2_outputs[2193] = layer1_outputs[557];
    assign layer2_outputs[2194] = (layer1_outputs[1287]) & (layer1_outputs[1590]);
    assign layer2_outputs[2195] = (layer1_outputs[2339]) & ~(layer1_outputs[2021]);
    assign layer2_outputs[2196] = layer1_outputs[2180];
    assign layer2_outputs[2197] = layer1_outputs[1219];
    assign layer2_outputs[2198] = (layer1_outputs[1916]) & ~(layer1_outputs[384]);
    assign layer2_outputs[2199] = (layer1_outputs[2340]) | (layer1_outputs[1634]);
    assign layer2_outputs[2200] = ~(layer1_outputs[2347]);
    assign layer2_outputs[2201] = ~(layer1_outputs[2286]);
    assign layer2_outputs[2202] = (layer1_outputs[2497]) & (layer1_outputs[2458]);
    assign layer2_outputs[2203] = ~(layer1_outputs[1095]) | (layer1_outputs[27]);
    assign layer2_outputs[2204] = layer1_outputs[38];
    assign layer2_outputs[2205] = 1'b1;
    assign layer2_outputs[2206] = (layer1_outputs[44]) & ~(layer1_outputs[1073]);
    assign layer2_outputs[2207] = ~(layer1_outputs[1589]);
    assign layer2_outputs[2208] = (layer1_outputs[917]) & (layer1_outputs[578]);
    assign layer2_outputs[2209] = ~(layer1_outputs[1714]) | (layer1_outputs[643]);
    assign layer2_outputs[2210] = ~((layer1_outputs[966]) | (layer1_outputs[533]));
    assign layer2_outputs[2211] = (layer1_outputs[556]) | (layer1_outputs[334]);
    assign layer2_outputs[2212] = ~((layer1_outputs[2360]) ^ (layer1_outputs[33]));
    assign layer2_outputs[2213] = ~((layer1_outputs[2345]) ^ (layer1_outputs[338]));
    assign layer2_outputs[2214] = ~(layer1_outputs[2086]);
    assign layer2_outputs[2215] = ~(layer1_outputs[882]);
    assign layer2_outputs[2216] = layer1_outputs[447];
    assign layer2_outputs[2217] = ~((layer1_outputs[1153]) | (layer1_outputs[2271]));
    assign layer2_outputs[2218] = (layer1_outputs[1034]) | (layer1_outputs[1025]);
    assign layer2_outputs[2219] = ~(layer1_outputs[724]);
    assign layer2_outputs[2220] = layer1_outputs[914];
    assign layer2_outputs[2221] = ~(layer1_outputs[1690]);
    assign layer2_outputs[2222] = 1'b0;
    assign layer2_outputs[2223] = ~(layer1_outputs[348]) | (layer1_outputs[645]);
    assign layer2_outputs[2224] = ~(layer1_outputs[1391]) | (layer1_outputs[695]);
    assign layer2_outputs[2225] = (layer1_outputs[944]) & ~(layer1_outputs[691]);
    assign layer2_outputs[2226] = ~(layer1_outputs[2125]);
    assign layer2_outputs[2227] = ~(layer1_outputs[178]);
    assign layer2_outputs[2228] = (layer1_outputs[2375]) & ~(layer1_outputs[443]);
    assign layer2_outputs[2229] = ~((layer1_outputs[2151]) ^ (layer1_outputs[2156]));
    assign layer2_outputs[2230] = layer1_outputs[953];
    assign layer2_outputs[2231] = ~((layer1_outputs[1079]) | (layer1_outputs[1988]));
    assign layer2_outputs[2232] = layer1_outputs[1086];
    assign layer2_outputs[2233] = ~(layer1_outputs[90]) | (layer1_outputs[427]);
    assign layer2_outputs[2234] = layer1_outputs[1762];
    assign layer2_outputs[2235] = layer1_outputs[1106];
    assign layer2_outputs[2236] = ~(layer1_outputs[773]) | (layer1_outputs[1422]);
    assign layer2_outputs[2237] = ~((layer1_outputs[2509]) & (layer1_outputs[1501]));
    assign layer2_outputs[2238] = (layer1_outputs[223]) & ~(layer1_outputs[1709]);
    assign layer2_outputs[2239] = ~(layer1_outputs[2214]) | (layer1_outputs[761]);
    assign layer2_outputs[2240] = layer1_outputs[2123];
    assign layer2_outputs[2241] = layer1_outputs[59];
    assign layer2_outputs[2242] = (layer1_outputs[1361]) & ~(layer1_outputs[2114]);
    assign layer2_outputs[2243] = (layer1_outputs[1242]) & ~(layer1_outputs[1445]);
    assign layer2_outputs[2244] = layer1_outputs[885];
    assign layer2_outputs[2245] = ~(layer1_outputs[979]);
    assign layer2_outputs[2246] = (layer1_outputs[162]) | (layer1_outputs[2139]);
    assign layer2_outputs[2247] = ~(layer1_outputs[698]) | (layer1_outputs[2073]);
    assign layer2_outputs[2248] = (layer1_outputs[1409]) & ~(layer1_outputs[1030]);
    assign layer2_outputs[2249] = ~(layer1_outputs[1221]);
    assign layer2_outputs[2250] = (layer1_outputs[1442]) & ~(layer1_outputs[1407]);
    assign layer2_outputs[2251] = ~((layer1_outputs[463]) & (layer1_outputs[1596]));
    assign layer2_outputs[2252] = (layer1_outputs[664]) | (layer1_outputs[214]);
    assign layer2_outputs[2253] = (layer1_outputs[1125]) | (layer1_outputs[2268]);
    assign layer2_outputs[2254] = ~(layer1_outputs[442]);
    assign layer2_outputs[2255] = ~(layer1_outputs[1415]) | (layer1_outputs[322]);
    assign layer2_outputs[2256] = ~((layer1_outputs[2319]) | (layer1_outputs[1764]));
    assign layer2_outputs[2257] = ~((layer1_outputs[897]) & (layer1_outputs[510]));
    assign layer2_outputs[2258] = 1'b0;
    assign layer2_outputs[2259] = (layer1_outputs[2043]) | (layer1_outputs[1782]);
    assign layer2_outputs[2260] = layer1_outputs[2548];
    assign layer2_outputs[2261] = layer1_outputs[1929];
    assign layer2_outputs[2262] = ~(layer1_outputs[2310]);
    assign layer2_outputs[2263] = (layer1_outputs[1692]) & (layer1_outputs[282]);
    assign layer2_outputs[2264] = layer1_outputs[376];
    assign layer2_outputs[2265] = (layer1_outputs[2298]) ^ (layer1_outputs[2471]);
    assign layer2_outputs[2266] = (layer1_outputs[816]) | (layer1_outputs[823]);
    assign layer2_outputs[2267] = ~((layer1_outputs[1506]) | (layer1_outputs[1448]));
    assign layer2_outputs[2268] = ~((layer1_outputs[2482]) & (layer1_outputs[2538]));
    assign layer2_outputs[2269] = layer1_outputs[1202];
    assign layer2_outputs[2270] = (layer1_outputs[2259]) & ~(layer1_outputs[104]);
    assign layer2_outputs[2271] = 1'b1;
    assign layer2_outputs[2272] = (layer1_outputs[2442]) & (layer1_outputs[910]);
    assign layer2_outputs[2273] = ~((layer1_outputs[1349]) & (layer1_outputs[811]));
    assign layer2_outputs[2274] = ~(layer1_outputs[1705]);
    assign layer2_outputs[2275] = ~(layer1_outputs[2365]);
    assign layer2_outputs[2276] = layer1_outputs[182];
    assign layer2_outputs[2277] = (layer1_outputs[89]) & ~(layer1_outputs[1136]);
    assign layer2_outputs[2278] = layer1_outputs[179];
    assign layer2_outputs[2279] = ~(layer1_outputs[1816]);
    assign layer2_outputs[2280] = (layer1_outputs[2339]) & ~(layer1_outputs[235]);
    assign layer2_outputs[2281] = ~(layer1_outputs[2245]);
    assign layer2_outputs[2282] = ~(layer1_outputs[1087]);
    assign layer2_outputs[2283] = (layer1_outputs[629]) & ~(layer1_outputs[678]);
    assign layer2_outputs[2284] = (layer1_outputs[523]) & ~(layer1_outputs[453]);
    assign layer2_outputs[2285] = ~(layer1_outputs[1508]);
    assign layer2_outputs[2286] = (layer1_outputs[900]) & (layer1_outputs[1994]);
    assign layer2_outputs[2287] = layer1_outputs[2281];
    assign layer2_outputs[2288] = layer1_outputs[237];
    assign layer2_outputs[2289] = ~((layer1_outputs[410]) ^ (layer1_outputs[97]));
    assign layer2_outputs[2290] = ~(layer1_outputs[1618]) | (layer1_outputs[1402]);
    assign layer2_outputs[2291] = ~(layer1_outputs[2515]) | (layer1_outputs[1208]);
    assign layer2_outputs[2292] = layer1_outputs[1475];
    assign layer2_outputs[2293] = ~(layer1_outputs[904]) | (layer1_outputs[2272]);
    assign layer2_outputs[2294] = layer1_outputs[1395];
    assign layer2_outputs[2295] = (layer1_outputs[1015]) ^ (layer1_outputs[1683]);
    assign layer2_outputs[2296] = ~(layer1_outputs[1259]);
    assign layer2_outputs[2297] = ~(layer1_outputs[2426]) | (layer1_outputs[584]);
    assign layer2_outputs[2298] = (layer1_outputs[1073]) | (layer1_outputs[2055]);
    assign layer2_outputs[2299] = (layer1_outputs[2308]) & ~(layer1_outputs[1691]);
    assign layer2_outputs[2300] = ~(layer1_outputs[143]);
    assign layer2_outputs[2301] = layer1_outputs[2351];
    assign layer2_outputs[2302] = (layer1_outputs[2075]) & (layer1_outputs[1360]);
    assign layer2_outputs[2303] = (layer1_outputs[1731]) | (layer1_outputs[2202]);
    assign layer2_outputs[2304] = ~((layer1_outputs[758]) | (layer1_outputs[1263]));
    assign layer2_outputs[2305] = ~(layer1_outputs[21]);
    assign layer2_outputs[2306] = ~(layer1_outputs[668]) | (layer1_outputs[1304]);
    assign layer2_outputs[2307] = layer1_outputs[1492];
    assign layer2_outputs[2308] = (layer1_outputs[611]) & ~(layer1_outputs[400]);
    assign layer2_outputs[2309] = (layer1_outputs[1017]) & ~(layer1_outputs[1376]);
    assign layer2_outputs[2310] = ~((layer1_outputs[1328]) | (layer1_outputs[1879]));
    assign layer2_outputs[2311] = ~(layer1_outputs[1204]) | (layer1_outputs[1152]);
    assign layer2_outputs[2312] = layer1_outputs[1313];
    assign layer2_outputs[2313] = layer1_outputs[1454];
    assign layer2_outputs[2314] = layer1_outputs[2165];
    assign layer2_outputs[2315] = ~((layer1_outputs[1674]) | (layer1_outputs[2019]));
    assign layer2_outputs[2316] = (layer1_outputs[1289]) & ~(layer1_outputs[23]);
    assign layer2_outputs[2317] = 1'b1;
    assign layer2_outputs[2318] = layer1_outputs[2392];
    assign layer2_outputs[2319] = layer1_outputs[342];
    assign layer2_outputs[2320] = ~(layer1_outputs[1174]);
    assign layer2_outputs[2321] = (layer1_outputs[207]) & (layer1_outputs[1611]);
    assign layer2_outputs[2322] = ~(layer1_outputs[1374]) | (layer1_outputs[1947]);
    assign layer2_outputs[2323] = ~(layer1_outputs[2243]);
    assign layer2_outputs[2324] = (layer1_outputs[851]) | (layer1_outputs[2543]);
    assign layer2_outputs[2325] = ~(layer1_outputs[446]);
    assign layer2_outputs[2326] = ~(layer1_outputs[272]) | (layer1_outputs[558]);
    assign layer2_outputs[2327] = (layer1_outputs[1894]) & ~(layer1_outputs[699]);
    assign layer2_outputs[2328] = 1'b1;
    assign layer2_outputs[2329] = ~(layer1_outputs[460]) | (layer1_outputs[2232]);
    assign layer2_outputs[2330] = layer1_outputs[2155];
    assign layer2_outputs[2331] = layer1_outputs[975];
    assign layer2_outputs[2332] = ~((layer1_outputs[1471]) & (layer1_outputs[590]));
    assign layer2_outputs[2333] = ~(layer1_outputs[1398]);
    assign layer2_outputs[2334] = (layer1_outputs[583]) & (layer1_outputs[1914]);
    assign layer2_outputs[2335] = (layer1_outputs[1941]) & ~(layer1_outputs[1562]);
    assign layer2_outputs[2336] = 1'b1;
    assign layer2_outputs[2337] = ~((layer1_outputs[2142]) & (layer1_outputs[225]));
    assign layer2_outputs[2338] = ~((layer1_outputs[908]) | (layer1_outputs[1079]));
    assign layer2_outputs[2339] = ~(layer1_outputs[284]);
    assign layer2_outputs[2340] = (layer1_outputs[92]) & ~(layer1_outputs[1564]);
    assign layer2_outputs[2341] = ~(layer1_outputs[2463]) | (layer1_outputs[14]);
    assign layer2_outputs[2342] = (layer1_outputs[515]) & (layer1_outputs[1938]);
    assign layer2_outputs[2343] = ~(layer1_outputs[2026]);
    assign layer2_outputs[2344] = (layer1_outputs[1971]) | (layer1_outputs[1601]);
    assign layer2_outputs[2345] = ~((layer1_outputs[1187]) & (layer1_outputs[1144]));
    assign layer2_outputs[2346] = ~(layer1_outputs[196]);
    assign layer2_outputs[2347] = ~((layer1_outputs[448]) & (layer1_outputs[786]));
    assign layer2_outputs[2348] = ~(layer1_outputs[2035]) | (layer1_outputs[1866]);
    assign layer2_outputs[2349] = (layer1_outputs[405]) ^ (layer1_outputs[1708]);
    assign layer2_outputs[2350] = ~(layer1_outputs[496]) | (layer1_outputs[2444]);
    assign layer2_outputs[2351] = 1'b0;
    assign layer2_outputs[2352] = ~(layer1_outputs[1332]);
    assign layer2_outputs[2353] = ~(layer1_outputs[1449]);
    assign layer2_outputs[2354] = ~(layer1_outputs[1287]) | (layer1_outputs[740]);
    assign layer2_outputs[2355] = ~(layer1_outputs[2215]);
    assign layer2_outputs[2356] = ~(layer1_outputs[1708]) | (layer1_outputs[1193]);
    assign layer2_outputs[2357] = 1'b0;
    assign layer2_outputs[2358] = (layer1_outputs[1927]) | (layer1_outputs[176]);
    assign layer2_outputs[2359] = (layer1_outputs[2540]) ^ (layer1_outputs[1176]);
    assign layer2_outputs[2360] = (layer1_outputs[892]) | (layer1_outputs[2427]);
    assign layer2_outputs[2361] = ~(layer1_outputs[64]) | (layer1_outputs[357]);
    assign layer2_outputs[2362] = ~(layer1_outputs[1717]);
    assign layer2_outputs[2363] = (layer1_outputs[591]) | (layer1_outputs[1497]);
    assign layer2_outputs[2364] = ~(layer1_outputs[715]);
    assign layer2_outputs[2365] = (layer1_outputs[2376]) & ~(layer1_outputs[397]);
    assign layer2_outputs[2366] = (layer1_outputs[1995]) & ~(layer1_outputs[2513]);
    assign layer2_outputs[2367] = (layer1_outputs[1765]) & ~(layer1_outputs[1226]);
    assign layer2_outputs[2368] = ~(layer1_outputs[1996]) | (layer1_outputs[1869]);
    assign layer2_outputs[2369] = (layer1_outputs[1207]) ^ (layer1_outputs[13]);
    assign layer2_outputs[2370] = (layer1_outputs[1465]) & ~(layer1_outputs[2511]);
    assign layer2_outputs[2371] = ~(layer1_outputs[2495]);
    assign layer2_outputs[2372] = 1'b1;
    assign layer2_outputs[2373] = layer1_outputs[1641];
    assign layer2_outputs[2374] = (layer1_outputs[926]) & ~(layer1_outputs[2000]);
    assign layer2_outputs[2375] = ~(layer1_outputs[915]);
    assign layer2_outputs[2376] = ~(layer1_outputs[456]) | (layer1_outputs[659]);
    assign layer2_outputs[2377] = ~((layer1_outputs[1911]) | (layer1_outputs[651]));
    assign layer2_outputs[2378] = ~((layer1_outputs[1849]) & (layer1_outputs[1531]));
    assign layer2_outputs[2379] = ~(layer1_outputs[968]) | (layer1_outputs[562]);
    assign layer2_outputs[2380] = layer1_outputs[683];
    assign layer2_outputs[2381] = (layer1_outputs[813]) & ~(layer1_outputs[516]);
    assign layer2_outputs[2382] = ~(layer1_outputs[1030]);
    assign layer2_outputs[2383] = (layer1_outputs[1439]) & ~(layer1_outputs[218]);
    assign layer2_outputs[2384] = ~((layer1_outputs[698]) | (layer1_outputs[336]));
    assign layer2_outputs[2385] = layer1_outputs[682];
    assign layer2_outputs[2386] = (layer1_outputs[563]) & (layer1_outputs[1051]);
    assign layer2_outputs[2387] = (layer1_outputs[2350]) | (layer1_outputs[72]);
    assign layer2_outputs[2388] = layer1_outputs[1055];
    assign layer2_outputs[2389] = (layer1_outputs[569]) & (layer1_outputs[1514]);
    assign layer2_outputs[2390] = (layer1_outputs[2130]) & (layer1_outputs[1878]);
    assign layer2_outputs[2391] = ~(layer1_outputs[2433]);
    assign layer2_outputs[2392] = 1'b1;
    assign layer2_outputs[2393] = (layer1_outputs[2553]) | (layer1_outputs[690]);
    assign layer2_outputs[2394] = ~(layer1_outputs[1120]);
    assign layer2_outputs[2395] = ~(layer1_outputs[1777]);
    assign layer2_outputs[2396] = ~(layer1_outputs[1231]) | (layer1_outputs[658]);
    assign layer2_outputs[2397] = ~(layer1_outputs[1147]);
    assign layer2_outputs[2398] = ~((layer1_outputs[2411]) & (layer1_outputs[50]));
    assign layer2_outputs[2399] = 1'b1;
    assign layer2_outputs[2400] = (layer1_outputs[1703]) & ~(layer1_outputs[1752]);
    assign layer2_outputs[2401] = layer1_outputs[2284];
    assign layer2_outputs[2402] = (layer1_outputs[1681]) & ~(layer1_outputs[1375]);
    assign layer2_outputs[2403] = ~((layer1_outputs[1107]) ^ (layer1_outputs[387]));
    assign layer2_outputs[2404] = 1'b1;
    assign layer2_outputs[2405] = (layer1_outputs[423]) | (layer1_outputs[561]);
    assign layer2_outputs[2406] = (layer1_outputs[2251]) & ~(layer1_outputs[1223]);
    assign layer2_outputs[2407] = (layer1_outputs[1464]) & (layer1_outputs[523]);
    assign layer2_outputs[2408] = ~((layer1_outputs[1160]) ^ (layer1_outputs[287]));
    assign layer2_outputs[2409] = ~(layer1_outputs[175]) | (layer1_outputs[2350]);
    assign layer2_outputs[2410] = (layer1_outputs[469]) & ~(layer1_outputs[253]);
    assign layer2_outputs[2411] = 1'b0;
    assign layer2_outputs[2412] = (layer1_outputs[889]) | (layer1_outputs[2191]);
    assign layer2_outputs[2413] = (layer1_outputs[338]) & ~(layer1_outputs[995]);
    assign layer2_outputs[2414] = ~(layer1_outputs[787]);
    assign layer2_outputs[2415] = ~((layer1_outputs[2536]) & (layer1_outputs[378]));
    assign layer2_outputs[2416] = (layer1_outputs[1317]) & (layer1_outputs[1378]);
    assign layer2_outputs[2417] = ~(layer1_outputs[911]) | (layer1_outputs[1838]);
    assign layer2_outputs[2418] = ~(layer1_outputs[1646]);
    assign layer2_outputs[2419] = (layer1_outputs[988]) | (layer1_outputs[29]);
    assign layer2_outputs[2420] = (layer1_outputs[307]) & ~(layer1_outputs[1741]);
    assign layer2_outputs[2421] = layer1_outputs[388];
    assign layer2_outputs[2422] = (layer1_outputs[1114]) & ~(layer1_outputs[257]);
    assign layer2_outputs[2423] = ~(layer1_outputs[395]) | (layer1_outputs[39]);
    assign layer2_outputs[2424] = (layer1_outputs[1744]) & ~(layer1_outputs[822]);
    assign layer2_outputs[2425] = ~(layer1_outputs[279]);
    assign layer2_outputs[2426] = ~(layer1_outputs[730]) | (layer1_outputs[265]);
    assign layer2_outputs[2427] = 1'b0;
    assign layer2_outputs[2428] = 1'b1;
    assign layer2_outputs[2429] = ~(layer1_outputs[347]);
    assign layer2_outputs[2430] = (layer1_outputs[2454]) & ~(layer1_outputs[173]);
    assign layer2_outputs[2431] = 1'b1;
    assign layer2_outputs[2432] = layer1_outputs[1794];
    assign layer2_outputs[2433] = layer1_outputs[1120];
    assign layer2_outputs[2434] = ~((layer1_outputs[497]) | (layer1_outputs[834]));
    assign layer2_outputs[2435] = ~(layer1_outputs[1594]);
    assign layer2_outputs[2436] = layer1_outputs[1056];
    assign layer2_outputs[2437] = ~((layer1_outputs[973]) & (layer1_outputs[2034]));
    assign layer2_outputs[2438] = ~(layer1_outputs[2318]);
    assign layer2_outputs[2439] = ~(layer1_outputs[1427]);
    assign layer2_outputs[2440] = (layer1_outputs[2373]) & ~(layer1_outputs[2291]);
    assign layer2_outputs[2441] = (layer1_outputs[2202]) & ~(layer1_outputs[421]);
    assign layer2_outputs[2442] = ~(layer1_outputs[971]) | (layer1_outputs[522]);
    assign layer2_outputs[2443] = layer1_outputs[1040];
    assign layer2_outputs[2444] = 1'b0;
    assign layer2_outputs[2445] = ~(layer1_outputs[2534]);
    assign layer2_outputs[2446] = 1'b1;
    assign layer2_outputs[2447] = layer1_outputs[1403];
    assign layer2_outputs[2448] = (layer1_outputs[2118]) & (layer1_outputs[817]);
    assign layer2_outputs[2449] = ~((layer1_outputs[1944]) ^ (layer1_outputs[1053]));
    assign layer2_outputs[2450] = 1'b1;
    assign layer2_outputs[2451] = ~(layer1_outputs[1438]);
    assign layer2_outputs[2452] = 1'b1;
    assign layer2_outputs[2453] = ~((layer1_outputs[2051]) | (layer1_outputs[1273]));
    assign layer2_outputs[2454] = ~(layer1_outputs[676]) | (layer1_outputs[1950]);
    assign layer2_outputs[2455] = (layer1_outputs[2529]) | (layer1_outputs[727]);
    assign layer2_outputs[2456] = layer1_outputs[2423];
    assign layer2_outputs[2457] = (layer1_outputs[324]) | (layer1_outputs[944]);
    assign layer2_outputs[2458] = layer1_outputs[1380];
    assign layer2_outputs[2459] = (layer1_outputs[68]) & ~(layer1_outputs[2448]);
    assign layer2_outputs[2460] = ~((layer1_outputs[752]) ^ (layer1_outputs[271]));
    assign layer2_outputs[2461] = (layer1_outputs[218]) | (layer1_outputs[196]);
    assign layer2_outputs[2462] = ~((layer1_outputs[2329]) ^ (layer1_outputs[1068]));
    assign layer2_outputs[2463] = (layer1_outputs[2124]) & (layer1_outputs[1758]);
    assign layer2_outputs[2464] = (layer1_outputs[665]) & (layer1_outputs[2399]);
    assign layer2_outputs[2465] = ~(layer1_outputs[263]);
    assign layer2_outputs[2466] = 1'b0;
    assign layer2_outputs[2467] = ~(layer1_outputs[1477]) | (layer1_outputs[989]);
    assign layer2_outputs[2468] = ~(layer1_outputs[2025]) | (layer1_outputs[2422]);
    assign layer2_outputs[2469] = ~(layer1_outputs[1569]);
    assign layer2_outputs[2470] = layer1_outputs[562];
    assign layer2_outputs[2471] = layer1_outputs[37];
    assign layer2_outputs[2472] = (layer1_outputs[1550]) & ~(layer1_outputs[1958]);
    assign layer2_outputs[2473] = (layer1_outputs[1803]) & ~(layer1_outputs[216]);
    assign layer2_outputs[2474] = (layer1_outputs[2122]) & (layer1_outputs[312]);
    assign layer2_outputs[2475] = 1'b1;
    assign layer2_outputs[2476] = (layer1_outputs[767]) & ~(layer1_outputs[1078]);
    assign layer2_outputs[2477] = ~(layer1_outputs[2160]) | (layer1_outputs[1470]);
    assign layer2_outputs[2478] = ~(layer1_outputs[2040]) | (layer1_outputs[1861]);
    assign layer2_outputs[2479] = layer1_outputs[28];
    assign layer2_outputs[2480] = layer1_outputs[1266];
    assign layer2_outputs[2481] = ~((layer1_outputs[248]) ^ (layer1_outputs[1888]));
    assign layer2_outputs[2482] = layer1_outputs[453];
    assign layer2_outputs[2483] = ~(layer1_outputs[344]) | (layer1_outputs[1369]);
    assign layer2_outputs[2484] = ~((layer1_outputs[1024]) ^ (layer1_outputs[2181]));
    assign layer2_outputs[2485] = layer1_outputs[2227];
    assign layer2_outputs[2486] = ~(layer1_outputs[257]);
    assign layer2_outputs[2487] = layer1_outputs[2197];
    assign layer2_outputs[2488] = 1'b0;
    assign layer2_outputs[2489] = layer1_outputs[966];
    assign layer2_outputs[2490] = ~(layer1_outputs[1466]);
    assign layer2_outputs[2491] = ~(layer1_outputs[202]);
    assign layer2_outputs[2492] = (layer1_outputs[1773]) & (layer1_outputs[1795]);
    assign layer2_outputs[2493] = ~(layer1_outputs[890]);
    assign layer2_outputs[2494] = ~((layer1_outputs[1881]) ^ (layer1_outputs[185]));
    assign layer2_outputs[2495] = layer1_outputs[1526];
    assign layer2_outputs[2496] = layer1_outputs[1534];
    assign layer2_outputs[2497] = layer1_outputs[765];
    assign layer2_outputs[2498] = ~((layer1_outputs[655]) & (layer1_outputs[1247]));
    assign layer2_outputs[2499] = ~(layer1_outputs[2149]);
    assign layer2_outputs[2500] = 1'b1;
    assign layer2_outputs[2501] = ~((layer1_outputs[399]) & (layer1_outputs[275]));
    assign layer2_outputs[2502] = ~(layer1_outputs[1548]);
    assign layer2_outputs[2503] = (layer1_outputs[2031]) & ~(layer1_outputs[2146]);
    assign layer2_outputs[2504] = layer1_outputs[1411];
    assign layer2_outputs[2505] = ~(layer1_outputs[2335]);
    assign layer2_outputs[2506] = ~(layer1_outputs[1096]) | (layer1_outputs[1520]);
    assign layer2_outputs[2507] = (layer1_outputs[1441]) & ~(layer1_outputs[2292]);
    assign layer2_outputs[2508] = layer1_outputs[603];
    assign layer2_outputs[2509] = ~(layer1_outputs[458]) | (layer1_outputs[1609]);
    assign layer2_outputs[2510] = ~((layer1_outputs[1980]) & (layer1_outputs[2381]));
    assign layer2_outputs[2511] = layer1_outputs[669];
    assign layer2_outputs[2512] = layer1_outputs[706];
    assign layer2_outputs[2513] = ~(layer1_outputs[1817]);
    assign layer2_outputs[2514] = layer1_outputs[342];
    assign layer2_outputs[2515] = (layer1_outputs[2061]) & ~(layer1_outputs[1291]);
    assign layer2_outputs[2516] = ~((layer1_outputs[22]) ^ (layer1_outputs[1738]));
    assign layer2_outputs[2517] = ~(layer1_outputs[1374]);
    assign layer2_outputs[2518] = (layer1_outputs[1805]) & ~(layer1_outputs[802]);
    assign layer2_outputs[2519] = ~(layer1_outputs[1309]) | (layer1_outputs[2294]);
    assign layer2_outputs[2520] = (layer1_outputs[434]) & ~(layer1_outputs[55]);
    assign layer2_outputs[2521] = ~(layer1_outputs[1921]);
    assign layer2_outputs[2522] = layer1_outputs[85];
    assign layer2_outputs[2523] = 1'b0;
    assign layer2_outputs[2524] = layer1_outputs[266];
    assign layer2_outputs[2525] = ~((layer1_outputs[1025]) | (layer1_outputs[1043]));
    assign layer2_outputs[2526] = layer1_outputs[1243];
    assign layer2_outputs[2527] = (layer1_outputs[595]) & (layer1_outputs[2424]);
    assign layer2_outputs[2528] = layer1_outputs[1792];
    assign layer2_outputs[2529] = (layer1_outputs[940]) | (layer1_outputs[2246]);
    assign layer2_outputs[2530] = 1'b1;
    assign layer2_outputs[2531] = ~(layer1_outputs[154]);
    assign layer2_outputs[2532] = ~(layer1_outputs[1230]) | (layer1_outputs[2083]);
    assign layer2_outputs[2533] = ~(layer1_outputs[261]);
    assign layer2_outputs[2534] = 1'b1;
    assign layer2_outputs[2535] = ~(layer1_outputs[1974]) | (layer1_outputs[896]);
    assign layer2_outputs[2536] = (layer1_outputs[428]) | (layer1_outputs[465]);
    assign layer2_outputs[2537] = layer1_outputs[55];
    assign layer2_outputs[2538] = layer1_outputs[1958];
    assign layer2_outputs[2539] = ~(layer1_outputs[1309]);
    assign layer2_outputs[2540] = layer1_outputs[1086];
    assign layer2_outputs[2541] = ~((layer1_outputs[382]) & (layer1_outputs[345]));
    assign layer2_outputs[2542] = 1'b1;
    assign layer2_outputs[2543] = 1'b0;
    assign layer2_outputs[2544] = layer1_outputs[2016];
    assign layer2_outputs[2545] = layer1_outputs[1864];
    assign layer2_outputs[2546] = layer1_outputs[683];
    assign layer2_outputs[2547] = (layer1_outputs[577]) & ~(layer1_outputs[797]);
    assign layer2_outputs[2548] = ~(layer1_outputs[2526]);
    assign layer2_outputs[2549] = 1'b0;
    assign layer2_outputs[2550] = ~(layer1_outputs[1545]) | (layer1_outputs[1382]);
    assign layer2_outputs[2551] = layer1_outputs[1443];
    assign layer2_outputs[2552] = ~(layer1_outputs[985]) | (layer1_outputs[2063]);
    assign layer2_outputs[2553] = ~((layer1_outputs[2]) & (layer1_outputs[1012]));
    assign layer2_outputs[2554] = ~(layer1_outputs[2234]) | (layer1_outputs[1386]);
    assign layer2_outputs[2555] = (layer1_outputs[337]) & ~(layer1_outputs[1355]);
    assign layer2_outputs[2556] = ~(layer1_outputs[1680]);
    assign layer2_outputs[2557] = ~(layer1_outputs[1546]) | (layer1_outputs[269]);
    assign layer2_outputs[2558] = 1'b0;
    assign layer2_outputs[2559] = ~(layer1_outputs[1728]);
    assign layer3_outputs[0] = ~(layer2_outputs[392]) | (layer2_outputs[1148]);
    assign layer3_outputs[1] = ~(layer2_outputs[2069]);
    assign layer3_outputs[2] = layer2_outputs[951];
    assign layer3_outputs[3] = (layer2_outputs[13]) & (layer2_outputs[2346]);
    assign layer3_outputs[4] = ~(layer2_outputs[1218]);
    assign layer3_outputs[5] = layer2_outputs[250];
    assign layer3_outputs[6] = (layer2_outputs[1871]) | (layer2_outputs[501]);
    assign layer3_outputs[7] = layer2_outputs[2405];
    assign layer3_outputs[8] = (layer2_outputs[2549]) | (layer2_outputs[1184]);
    assign layer3_outputs[9] = (layer2_outputs[79]) | (layer2_outputs[468]);
    assign layer3_outputs[10] = layer2_outputs[1590];
    assign layer3_outputs[11] = ~((layer2_outputs[2246]) ^ (layer2_outputs[920]));
    assign layer3_outputs[12] = layer2_outputs[497];
    assign layer3_outputs[13] = (layer2_outputs[2355]) ^ (layer2_outputs[1710]);
    assign layer3_outputs[14] = (layer2_outputs[1039]) | (layer2_outputs[197]);
    assign layer3_outputs[15] = ~(layer2_outputs[785]);
    assign layer3_outputs[16] = ~(layer2_outputs[1667]);
    assign layer3_outputs[17] = ~(layer2_outputs[2085]);
    assign layer3_outputs[18] = layer2_outputs[2015];
    assign layer3_outputs[19] = ~((layer2_outputs[1907]) ^ (layer2_outputs[184]));
    assign layer3_outputs[20] = layer2_outputs[2417];
    assign layer3_outputs[21] = ~(layer2_outputs[1112]);
    assign layer3_outputs[22] = ~((layer2_outputs[2087]) | (layer2_outputs[1606]));
    assign layer3_outputs[23] = ~(layer2_outputs[1130]);
    assign layer3_outputs[24] = layer2_outputs[937];
    assign layer3_outputs[25] = ~(layer2_outputs[2292]);
    assign layer3_outputs[26] = ~(layer2_outputs[840]);
    assign layer3_outputs[27] = ~(layer2_outputs[2114]);
    assign layer3_outputs[28] = (layer2_outputs[315]) & (layer2_outputs[1886]);
    assign layer3_outputs[29] = ~(layer2_outputs[2290]);
    assign layer3_outputs[30] = ~(layer2_outputs[1095]);
    assign layer3_outputs[31] = (layer2_outputs[2052]) & ~(layer2_outputs[411]);
    assign layer3_outputs[32] = ~(layer2_outputs[636]) | (layer2_outputs[943]);
    assign layer3_outputs[33] = ~(layer2_outputs[1317]);
    assign layer3_outputs[34] = ~(layer2_outputs[1137]);
    assign layer3_outputs[35] = (layer2_outputs[1293]) & ~(layer2_outputs[1368]);
    assign layer3_outputs[36] = layer2_outputs[1858];
    assign layer3_outputs[37] = ~(layer2_outputs[1346]);
    assign layer3_outputs[38] = (layer2_outputs[2131]) & ~(layer2_outputs[2370]);
    assign layer3_outputs[39] = layer2_outputs[1387];
    assign layer3_outputs[40] = ~(layer2_outputs[2117]);
    assign layer3_outputs[41] = (layer2_outputs[2372]) & ~(layer2_outputs[784]);
    assign layer3_outputs[42] = (layer2_outputs[1762]) & ~(layer2_outputs[83]);
    assign layer3_outputs[43] = ~(layer2_outputs[36]);
    assign layer3_outputs[44] = ~((layer2_outputs[243]) & (layer2_outputs[36]));
    assign layer3_outputs[45] = ~(layer2_outputs[2554]);
    assign layer3_outputs[46] = ~(layer2_outputs[1387]);
    assign layer3_outputs[47] = ~(layer2_outputs[1485]);
    assign layer3_outputs[48] = (layer2_outputs[611]) & ~(layer2_outputs[2332]);
    assign layer3_outputs[49] = (layer2_outputs[2012]) | (layer2_outputs[1427]);
    assign layer3_outputs[50] = ~((layer2_outputs[2412]) ^ (layer2_outputs[866]));
    assign layer3_outputs[51] = ~(layer2_outputs[589]);
    assign layer3_outputs[52] = layer2_outputs[1357];
    assign layer3_outputs[53] = ~(layer2_outputs[2288]);
    assign layer3_outputs[54] = ~(layer2_outputs[814]) | (layer2_outputs[162]);
    assign layer3_outputs[55] = (layer2_outputs[1078]) & ~(layer2_outputs[549]);
    assign layer3_outputs[56] = ~((layer2_outputs[1899]) & (layer2_outputs[754]));
    assign layer3_outputs[57] = (layer2_outputs[881]) ^ (layer2_outputs[1279]);
    assign layer3_outputs[58] = ~(layer2_outputs[2218]);
    assign layer3_outputs[59] = ~(layer2_outputs[1]) | (layer2_outputs[1674]);
    assign layer3_outputs[60] = layer2_outputs[1901];
    assign layer3_outputs[61] = ~(layer2_outputs[451]) | (layer2_outputs[388]);
    assign layer3_outputs[62] = ~(layer2_outputs[2484]);
    assign layer3_outputs[63] = ~(layer2_outputs[2200]) | (layer2_outputs[1582]);
    assign layer3_outputs[64] = (layer2_outputs[2102]) | (layer2_outputs[1775]);
    assign layer3_outputs[65] = ~(layer2_outputs[2210]);
    assign layer3_outputs[66] = layer2_outputs[1884];
    assign layer3_outputs[67] = (layer2_outputs[362]) & (layer2_outputs[1880]);
    assign layer3_outputs[68] = ~(layer2_outputs[2188]);
    assign layer3_outputs[69] = ~(layer2_outputs[1842]);
    assign layer3_outputs[70] = ~(layer2_outputs[165]) | (layer2_outputs[1809]);
    assign layer3_outputs[71] = ~(layer2_outputs[379]);
    assign layer3_outputs[72] = ~((layer2_outputs[2489]) ^ (layer2_outputs[1266]));
    assign layer3_outputs[73] = ~(layer2_outputs[609]);
    assign layer3_outputs[74] = ~(layer2_outputs[623]);
    assign layer3_outputs[75] = (layer2_outputs[2123]) & ~(layer2_outputs[2417]);
    assign layer3_outputs[76] = ~(layer2_outputs[26]);
    assign layer3_outputs[77] = ~((layer2_outputs[291]) & (layer2_outputs[869]));
    assign layer3_outputs[78] = (layer2_outputs[660]) | (layer2_outputs[1889]);
    assign layer3_outputs[79] = (layer2_outputs[181]) | (layer2_outputs[504]);
    assign layer3_outputs[80] = ~((layer2_outputs[955]) & (layer2_outputs[896]));
    assign layer3_outputs[81] = (layer2_outputs[41]) | (layer2_outputs[1350]);
    assign layer3_outputs[82] = ~(layer2_outputs[1627]);
    assign layer3_outputs[83] = ~(layer2_outputs[118]) | (layer2_outputs[1536]);
    assign layer3_outputs[84] = (layer2_outputs[281]) ^ (layer2_outputs[2476]);
    assign layer3_outputs[85] = ~(layer2_outputs[1113]);
    assign layer3_outputs[86] = ~(layer2_outputs[1955]) | (layer2_outputs[2457]);
    assign layer3_outputs[87] = (layer2_outputs[1629]) ^ (layer2_outputs[1961]);
    assign layer3_outputs[88] = ~(layer2_outputs[1296]);
    assign layer3_outputs[89] = ~(layer2_outputs[420]) | (layer2_outputs[1891]);
    assign layer3_outputs[90] = ~(layer2_outputs[678]) | (layer2_outputs[965]);
    assign layer3_outputs[91] = ~(layer2_outputs[804]);
    assign layer3_outputs[92] = ~(layer2_outputs[2464]);
    assign layer3_outputs[93] = ~((layer2_outputs[901]) & (layer2_outputs[182]));
    assign layer3_outputs[94] = 1'b0;
    assign layer3_outputs[95] = (layer2_outputs[1791]) & ~(layer2_outputs[2523]);
    assign layer3_outputs[96] = 1'b0;
    assign layer3_outputs[97] = layer2_outputs[242];
    assign layer3_outputs[98] = ~(layer2_outputs[2378]);
    assign layer3_outputs[99] = ~(layer2_outputs[1173]) | (layer2_outputs[2105]);
    assign layer3_outputs[100] = ~(layer2_outputs[555]);
    assign layer3_outputs[101] = layer2_outputs[699];
    assign layer3_outputs[102] = (layer2_outputs[1424]) | (layer2_outputs[1603]);
    assign layer3_outputs[103] = (layer2_outputs[733]) & ~(layer2_outputs[1994]);
    assign layer3_outputs[104] = layer2_outputs[2000];
    assign layer3_outputs[105] = ~(layer2_outputs[1568]) | (layer2_outputs[1252]);
    assign layer3_outputs[106] = (layer2_outputs[1250]) & ~(layer2_outputs[1501]);
    assign layer3_outputs[107] = ~(layer2_outputs[2156]) | (layer2_outputs[750]);
    assign layer3_outputs[108] = ~(layer2_outputs[1631]);
    assign layer3_outputs[109] = ~(layer2_outputs[544]);
    assign layer3_outputs[110] = ~(layer2_outputs[1056]) | (layer2_outputs[1792]);
    assign layer3_outputs[111] = layer2_outputs[1080];
    assign layer3_outputs[112] = layer2_outputs[1413];
    assign layer3_outputs[113] = (layer2_outputs[632]) & ~(layer2_outputs[766]);
    assign layer3_outputs[114] = ~((layer2_outputs[608]) & (layer2_outputs[217]));
    assign layer3_outputs[115] = (layer2_outputs[2177]) & ~(layer2_outputs[2467]);
    assign layer3_outputs[116] = ~(layer2_outputs[361]);
    assign layer3_outputs[117] = 1'b1;
    assign layer3_outputs[118] = (layer2_outputs[622]) & ~(layer2_outputs[963]);
    assign layer3_outputs[119] = 1'b0;
    assign layer3_outputs[120] = (layer2_outputs[778]) & ~(layer2_outputs[16]);
    assign layer3_outputs[121] = ~(layer2_outputs[2379]);
    assign layer3_outputs[122] = 1'b0;
    assign layer3_outputs[123] = ~(layer2_outputs[1613]);
    assign layer3_outputs[124] = ~(layer2_outputs[448]);
    assign layer3_outputs[125] = layer2_outputs[1059];
    assign layer3_outputs[126] = ~((layer2_outputs[2349]) ^ (layer2_outputs[1926]));
    assign layer3_outputs[127] = ~(layer2_outputs[1049]);
    assign layer3_outputs[128] = ~(layer2_outputs[1471]);
    assign layer3_outputs[129] = (layer2_outputs[1060]) & ~(layer2_outputs[101]);
    assign layer3_outputs[130] = (layer2_outputs[1709]) | (layer2_outputs[1287]);
    assign layer3_outputs[131] = 1'b1;
    assign layer3_outputs[132] = layer2_outputs[358];
    assign layer3_outputs[133] = ~(layer2_outputs[1826]);
    assign layer3_outputs[134] = (layer2_outputs[100]) ^ (layer2_outputs[1162]);
    assign layer3_outputs[135] = (layer2_outputs[1494]) | (layer2_outputs[886]);
    assign layer3_outputs[136] = layer2_outputs[619];
    assign layer3_outputs[137] = ~(layer2_outputs[2250]) | (layer2_outputs[1665]);
    assign layer3_outputs[138] = 1'b0;
    assign layer3_outputs[139] = (layer2_outputs[2160]) | (layer2_outputs[856]);
    assign layer3_outputs[140] = (layer2_outputs[2024]) | (layer2_outputs[454]);
    assign layer3_outputs[141] = (layer2_outputs[1334]) & ~(layer2_outputs[2432]);
    assign layer3_outputs[142] = ~(layer2_outputs[509]) | (layer2_outputs[1643]);
    assign layer3_outputs[143] = ~((layer2_outputs[2307]) & (layer2_outputs[915]));
    assign layer3_outputs[144] = (layer2_outputs[1837]) | (layer2_outputs[2118]);
    assign layer3_outputs[145] = ~(layer2_outputs[1553]);
    assign layer3_outputs[146] = (layer2_outputs[407]) & ~(layer2_outputs[1764]);
    assign layer3_outputs[147] = ~((layer2_outputs[1344]) ^ (layer2_outputs[2308]));
    assign layer3_outputs[148] = ~(layer2_outputs[156]) | (layer2_outputs[2402]);
    assign layer3_outputs[149] = ~(layer2_outputs[935]) | (layer2_outputs[2410]);
    assign layer3_outputs[150] = ~((layer2_outputs[1861]) & (layer2_outputs[531]));
    assign layer3_outputs[151] = ~((layer2_outputs[1775]) ^ (layer2_outputs[1854]));
    assign layer3_outputs[152] = (layer2_outputs[1956]) | (layer2_outputs[855]);
    assign layer3_outputs[153] = (layer2_outputs[1890]) & ~(layer2_outputs[124]);
    assign layer3_outputs[154] = 1'b0;
    assign layer3_outputs[155] = (layer2_outputs[857]) & ~(layer2_outputs[2265]);
    assign layer3_outputs[156] = ~(layer2_outputs[1005]) | (layer2_outputs[1236]);
    assign layer3_outputs[157] = ~(layer2_outputs[781]);
    assign layer3_outputs[158] = ~((layer2_outputs[2334]) | (layer2_outputs[552]));
    assign layer3_outputs[159] = layer2_outputs[2141];
    assign layer3_outputs[160] = layer2_outputs[1284];
    assign layer3_outputs[161] = ~((layer2_outputs[727]) ^ (layer2_outputs[1321]));
    assign layer3_outputs[162] = ~(layer2_outputs[2393]);
    assign layer3_outputs[163] = (layer2_outputs[884]) | (layer2_outputs[613]);
    assign layer3_outputs[164] = ~(layer2_outputs[2044]);
    assign layer3_outputs[165] = (layer2_outputs[2165]) | (layer2_outputs[193]);
    assign layer3_outputs[166] = ~(layer2_outputs[944]) | (layer2_outputs[692]);
    assign layer3_outputs[167] = ~(layer2_outputs[67]);
    assign layer3_outputs[168] = ~((layer2_outputs[1888]) ^ (layer2_outputs[1707]));
    assign layer3_outputs[169] = ~(layer2_outputs[1435]);
    assign layer3_outputs[170] = (layer2_outputs[1235]) & ~(layer2_outputs[1100]);
    assign layer3_outputs[171] = ~(layer2_outputs[1158]);
    assign layer3_outputs[172] = ~(layer2_outputs[2303]);
    assign layer3_outputs[173] = 1'b0;
    assign layer3_outputs[174] = (layer2_outputs[2460]) & ~(layer2_outputs[1045]);
    assign layer3_outputs[175] = ~(layer2_outputs[1138]);
    assign layer3_outputs[176] = (layer2_outputs[2018]) | (layer2_outputs[1757]);
    assign layer3_outputs[177] = ~(layer2_outputs[141]);
    assign layer3_outputs[178] = ~(layer2_outputs[528]);
    assign layer3_outputs[179] = 1'b0;
    assign layer3_outputs[180] = ~((layer2_outputs[416]) | (layer2_outputs[2386]));
    assign layer3_outputs[181] = ~(layer2_outputs[1203]) | (layer2_outputs[596]);
    assign layer3_outputs[182] = layer2_outputs[1169];
    assign layer3_outputs[183] = ~((layer2_outputs[1329]) | (layer2_outputs[485]));
    assign layer3_outputs[184] = 1'b1;
    assign layer3_outputs[185] = ~((layer2_outputs[2352]) & (layer2_outputs[1798]));
    assign layer3_outputs[186] = layer2_outputs[844];
    assign layer3_outputs[187] = (layer2_outputs[628]) & ~(layer2_outputs[1269]);
    assign layer3_outputs[188] = ~(layer2_outputs[2362]);
    assign layer3_outputs[189] = ~((layer2_outputs[2488]) ^ (layer2_outputs[1604]));
    assign layer3_outputs[190] = layer2_outputs[2546];
    assign layer3_outputs[191] = ~(layer2_outputs[1064]) | (layer2_outputs[1769]);
    assign layer3_outputs[192] = layer2_outputs[1831];
    assign layer3_outputs[193] = ~(layer2_outputs[1106]);
    assign layer3_outputs[194] = ~(layer2_outputs[997]);
    assign layer3_outputs[195] = (layer2_outputs[1817]) ^ (layer2_outputs[1053]);
    assign layer3_outputs[196] = ~((layer2_outputs[1161]) ^ (layer2_outputs[940]));
    assign layer3_outputs[197] = (layer2_outputs[897]) & (layer2_outputs[2434]);
    assign layer3_outputs[198] = ~(layer2_outputs[270]);
    assign layer3_outputs[199] = 1'b1;
    assign layer3_outputs[200] = 1'b1;
    assign layer3_outputs[201] = ~(layer2_outputs[2116]);
    assign layer3_outputs[202] = 1'b1;
    assign layer3_outputs[203] = ~((layer2_outputs[2360]) | (layer2_outputs[615]));
    assign layer3_outputs[204] = ~(layer2_outputs[1846]);
    assign layer3_outputs[205] = ~(layer2_outputs[8]) | (layer2_outputs[1399]);
    assign layer3_outputs[206] = (layer2_outputs[56]) ^ (layer2_outputs[2411]);
    assign layer3_outputs[207] = ~((layer2_outputs[329]) & (layer2_outputs[1728]));
    assign layer3_outputs[208] = ~(layer2_outputs[1371]) | (layer2_outputs[2068]);
    assign layer3_outputs[209] = ~((layer2_outputs[1334]) & (layer2_outputs[371]));
    assign layer3_outputs[210] = ~(layer2_outputs[1531]) | (layer2_outputs[484]);
    assign layer3_outputs[211] = ~(layer2_outputs[1998]) | (layer2_outputs[302]);
    assign layer3_outputs[212] = layer2_outputs[219];
    assign layer3_outputs[213] = layer2_outputs[37];
    assign layer3_outputs[214] = ~(layer2_outputs[179]);
    assign layer3_outputs[215] = ~((layer2_outputs[1004]) | (layer2_outputs[1379]));
    assign layer3_outputs[216] = ~(layer2_outputs[1834]);
    assign layer3_outputs[217] = ~(layer2_outputs[2498]) | (layer2_outputs[1200]);
    assign layer3_outputs[218] = ~(layer2_outputs[653]);
    assign layer3_outputs[219] = ~(layer2_outputs[2321]);
    assign layer3_outputs[220] = ~((layer2_outputs[2318]) & (layer2_outputs[602]));
    assign layer3_outputs[221] = ~(layer2_outputs[2005]);
    assign layer3_outputs[222] = layer2_outputs[1024];
    assign layer3_outputs[223] = (layer2_outputs[741]) & (layer2_outputs[2076]);
    assign layer3_outputs[224] = (layer2_outputs[51]) & (layer2_outputs[1085]);
    assign layer3_outputs[225] = (layer2_outputs[285]) & (layer2_outputs[537]);
    assign layer3_outputs[226] = ~(layer2_outputs[2137]);
    assign layer3_outputs[227] = ~(layer2_outputs[562]);
    assign layer3_outputs[228] = ~(layer2_outputs[475]);
    assign layer3_outputs[229] = (layer2_outputs[1659]) | (layer2_outputs[225]);
    assign layer3_outputs[230] = (layer2_outputs[1772]) ^ (layer2_outputs[914]);
    assign layer3_outputs[231] = ~((layer2_outputs[387]) | (layer2_outputs[617]));
    assign layer3_outputs[232] = (layer2_outputs[303]) | (layer2_outputs[2090]);
    assign layer3_outputs[233] = (layer2_outputs[64]) & (layer2_outputs[2403]);
    assign layer3_outputs[234] = ~((layer2_outputs[2095]) ^ (layer2_outputs[285]));
    assign layer3_outputs[235] = ~(layer2_outputs[2407]);
    assign layer3_outputs[236] = (layer2_outputs[496]) & ~(layer2_outputs[690]);
    assign layer3_outputs[237] = layer2_outputs[779];
    assign layer3_outputs[238] = (layer2_outputs[1117]) | (layer2_outputs[2240]);
    assign layer3_outputs[239] = 1'b1;
    assign layer3_outputs[240] = ~(layer2_outputs[1223]);
    assign layer3_outputs[241] = ~(layer2_outputs[857]);
    assign layer3_outputs[242] = 1'b0;
    assign layer3_outputs[243] = (layer2_outputs[1799]) & ~(layer2_outputs[1417]);
    assign layer3_outputs[244] = layer2_outputs[2394];
    assign layer3_outputs[245] = ~(layer2_outputs[2299]);
    assign layer3_outputs[246] = layer2_outputs[1601];
    assign layer3_outputs[247] = ~(layer2_outputs[1942]);
    assign layer3_outputs[248] = (layer2_outputs[1729]) & ~(layer2_outputs[1804]);
    assign layer3_outputs[249] = (layer2_outputs[435]) ^ (layer2_outputs[2255]);
    assign layer3_outputs[250] = ~(layer2_outputs[114]) | (layer2_outputs[1124]);
    assign layer3_outputs[251] = (layer2_outputs[880]) | (layer2_outputs[1191]);
    assign layer3_outputs[252] = ~(layer2_outputs[1701]);
    assign layer3_outputs[253] = (layer2_outputs[1348]) | (layer2_outputs[336]);
    assign layer3_outputs[254] = (layer2_outputs[739]) & (layer2_outputs[1188]);
    assign layer3_outputs[255] = ~((layer2_outputs[1967]) ^ (layer2_outputs[853]));
    assign layer3_outputs[256] = layer2_outputs[619];
    assign layer3_outputs[257] = (layer2_outputs[2119]) & ~(layer2_outputs[1374]);
    assign layer3_outputs[258] = (layer2_outputs[653]) & (layer2_outputs[423]);
    assign layer3_outputs[259] = (layer2_outputs[396]) & ~(layer2_outputs[156]);
    assign layer3_outputs[260] = layer2_outputs[1635];
    assign layer3_outputs[261] = (layer2_outputs[1185]) & ~(layer2_outputs[189]);
    assign layer3_outputs[262] = (layer2_outputs[1366]) ^ (layer2_outputs[583]);
    assign layer3_outputs[263] = layer2_outputs[502];
    assign layer3_outputs[264] = layer2_outputs[2347];
    assign layer3_outputs[265] = (layer2_outputs[1300]) & ~(layer2_outputs[1598]);
    assign layer3_outputs[266] = layer2_outputs[1678];
    assign layer3_outputs[267] = 1'b1;
    assign layer3_outputs[268] = layer2_outputs[1187];
    assign layer3_outputs[269] = ~(layer2_outputs[2054]);
    assign layer3_outputs[270] = ~((layer2_outputs[960]) | (layer2_outputs[1318]));
    assign layer3_outputs[271] = layer2_outputs[542];
    assign layer3_outputs[272] = ~(layer2_outputs[1413]) | (layer2_outputs[1308]);
    assign layer3_outputs[273] = layer2_outputs[2343];
    assign layer3_outputs[274] = (layer2_outputs[988]) & ~(layer2_outputs[2220]);
    assign layer3_outputs[275] = (layer2_outputs[2470]) | (layer2_outputs[1336]);
    assign layer3_outputs[276] = ~((layer2_outputs[1341]) & (layer2_outputs[456]));
    assign layer3_outputs[277] = ~(layer2_outputs[2459]) | (layer2_outputs[1766]);
    assign layer3_outputs[278] = ~((layer2_outputs[671]) & (layer2_outputs[2490]));
    assign layer3_outputs[279] = layer2_outputs[159];
    assign layer3_outputs[280] = layer2_outputs[1292];
    assign layer3_outputs[281] = 1'b1;
    assign layer3_outputs[282] = ~(layer2_outputs[1514]);
    assign layer3_outputs[283] = ~(layer2_outputs[626]) | (layer2_outputs[2066]);
    assign layer3_outputs[284] = ~((layer2_outputs[2533]) & (layer2_outputs[2088]));
    assign layer3_outputs[285] = layer2_outputs[1726];
    assign layer3_outputs[286] = ~(layer2_outputs[2461]);
    assign layer3_outputs[287] = ~(layer2_outputs[1515]);
    assign layer3_outputs[288] = ~(layer2_outputs[733]);
    assign layer3_outputs[289] = 1'b1;
    assign layer3_outputs[290] = ~((layer2_outputs[2145]) & (layer2_outputs[2297]));
    assign layer3_outputs[291] = ~((layer2_outputs[734]) & (layer2_outputs[2058]));
    assign layer3_outputs[292] = (layer2_outputs[2112]) & ~(layer2_outputs[1283]);
    assign layer3_outputs[293] = ~((layer2_outputs[367]) & (layer2_outputs[1955]));
    assign layer3_outputs[294] = layer2_outputs[1821];
    assign layer3_outputs[295] = (layer2_outputs[2511]) & ~(layer2_outputs[2060]);
    assign layer3_outputs[296] = layer2_outputs[2330];
    assign layer3_outputs[297] = layer2_outputs[2544];
    assign layer3_outputs[298] = 1'b0;
    assign layer3_outputs[299] = (layer2_outputs[117]) & (layer2_outputs[1197]);
    assign layer3_outputs[300] = ~((layer2_outputs[823]) ^ (layer2_outputs[1705]));
    assign layer3_outputs[301] = ~(layer2_outputs[567]);
    assign layer3_outputs[302] = (layer2_outputs[1990]) ^ (layer2_outputs[2267]);
    assign layer3_outputs[303] = ~(layer2_outputs[2456]);
    assign layer3_outputs[304] = ~(layer2_outputs[20]);
    assign layer3_outputs[305] = ~(layer2_outputs[711]) | (layer2_outputs[1477]);
    assign layer3_outputs[306] = ~(layer2_outputs[1128]) | (layer2_outputs[1328]);
    assign layer3_outputs[307] = (layer2_outputs[2048]) ^ (layer2_outputs[1031]);
    assign layer3_outputs[308] = ~(layer2_outputs[1087]);
    assign layer3_outputs[309] = ~(layer2_outputs[1978]) | (layer2_outputs[466]);
    assign layer3_outputs[310] = (layer2_outputs[2404]) & ~(layer2_outputs[1443]);
    assign layer3_outputs[311] = layer2_outputs[2407];
    assign layer3_outputs[312] = ~(layer2_outputs[591]) | (layer2_outputs[664]);
    assign layer3_outputs[313] = ~(layer2_outputs[1527]) | (layer2_outputs[1242]);
    assign layer3_outputs[314] = layer2_outputs[902];
    assign layer3_outputs[315] = ~(layer2_outputs[1236]) | (layer2_outputs[2356]);
    assign layer3_outputs[316] = ~(layer2_outputs[1711]);
    assign layer3_outputs[317] = layer2_outputs[2216];
    assign layer3_outputs[318] = ~(layer2_outputs[572]);
    assign layer3_outputs[319] = (layer2_outputs[2387]) | (layer2_outputs[1545]);
    assign layer3_outputs[320] = (layer2_outputs[703]) & (layer2_outputs[531]);
    assign layer3_outputs[321] = ~(layer2_outputs[1903]) | (layer2_outputs[2128]);
    assign layer3_outputs[322] = layer2_outputs[2232];
    assign layer3_outputs[323] = layer2_outputs[1758];
    assign layer3_outputs[324] = layer2_outputs[2282];
    assign layer3_outputs[325] = ~(layer2_outputs[893]) | (layer2_outputs[513]);
    assign layer3_outputs[326] = (layer2_outputs[166]) | (layer2_outputs[401]);
    assign layer3_outputs[327] = (layer2_outputs[1299]) & (layer2_outputs[771]);
    assign layer3_outputs[328] = (layer2_outputs[2181]) ^ (layer2_outputs[510]);
    assign layer3_outputs[329] = ~((layer2_outputs[819]) ^ (layer2_outputs[2427]));
    assign layer3_outputs[330] = (layer2_outputs[1823]) & (layer2_outputs[1030]);
    assign layer3_outputs[331] = ~(layer2_outputs[92]) | (layer2_outputs[435]);
    assign layer3_outputs[332] = (layer2_outputs[2069]) & (layer2_outputs[720]);
    assign layer3_outputs[333] = (layer2_outputs[1278]) & (layer2_outputs[1562]);
    assign layer3_outputs[334] = (layer2_outputs[966]) & ~(layer2_outputs[2298]);
    assign layer3_outputs[335] = ~((layer2_outputs[2122]) | (layer2_outputs[1520]));
    assign layer3_outputs[336] = 1'b1;
    assign layer3_outputs[337] = (layer2_outputs[828]) | (layer2_outputs[1287]);
    assign layer3_outputs[338] = ~(layer2_outputs[2351]);
    assign layer3_outputs[339] = (layer2_outputs[129]) | (layer2_outputs[1336]);
    assign layer3_outputs[340] = ~(layer2_outputs[1508]);
    assign layer3_outputs[341] = ~(layer2_outputs[765]);
    assign layer3_outputs[342] = ~(layer2_outputs[1683]);
    assign layer3_outputs[343] = ~(layer2_outputs[1289]);
    assign layer3_outputs[344] = ~((layer2_outputs[1837]) & (layer2_outputs[1941]));
    assign layer3_outputs[345] = ~(layer2_outputs[794]);
    assign layer3_outputs[346] = (layer2_outputs[448]) & (layer2_outputs[1674]);
    assign layer3_outputs[347] = ~(layer2_outputs[2287]);
    assign layer3_outputs[348] = (layer2_outputs[1924]) & ~(layer2_outputs[2013]);
    assign layer3_outputs[349] = ~((layer2_outputs[1335]) & (layer2_outputs[889]));
    assign layer3_outputs[350] = layer2_outputs[2531];
    assign layer3_outputs[351] = ~((layer2_outputs[1305]) | (layer2_outputs[753]));
    assign layer3_outputs[352] = ~(layer2_outputs[463]);
    assign layer3_outputs[353] = layer2_outputs[319];
    assign layer3_outputs[354] = (layer2_outputs[173]) & ~(layer2_outputs[1402]);
    assign layer3_outputs[355] = layer2_outputs[679];
    assign layer3_outputs[356] = ~(layer2_outputs[1077]);
    assign layer3_outputs[357] = (layer2_outputs[1325]) ^ (layer2_outputs[89]);
    assign layer3_outputs[358] = ~(layer2_outputs[1376]) | (layer2_outputs[985]);
    assign layer3_outputs[359] = ~((layer2_outputs[2057]) & (layer2_outputs[185]));
    assign layer3_outputs[360] = ~((layer2_outputs[2246]) & (layer2_outputs[249]));
    assign layer3_outputs[361] = ~(layer2_outputs[469]);
    assign layer3_outputs[362] = layer2_outputs[1859];
    assign layer3_outputs[363] = 1'b1;
    assign layer3_outputs[364] = ~((layer2_outputs[1217]) ^ (layer2_outputs[851]));
    assign layer3_outputs[365] = ~(layer2_outputs[701]) | (layer2_outputs[9]);
    assign layer3_outputs[366] = layer2_outputs[2315];
    assign layer3_outputs[367] = layer2_outputs[1003];
    assign layer3_outputs[368] = ~(layer2_outputs[296]);
    assign layer3_outputs[369] = ~(layer2_outputs[1386]);
    assign layer3_outputs[370] = (layer2_outputs[624]) | (layer2_outputs[1410]);
    assign layer3_outputs[371] = (layer2_outputs[2451]) & (layer2_outputs[1008]);
    assign layer3_outputs[372] = ~(layer2_outputs[1693]);
    assign layer3_outputs[373] = (layer2_outputs[1759]) | (layer2_outputs[1568]);
    assign layer3_outputs[374] = ~((layer2_outputs[147]) & (layer2_outputs[2472]));
    assign layer3_outputs[375] = ~((layer2_outputs[1977]) & (layer2_outputs[426]));
    assign layer3_outputs[376] = ~(layer2_outputs[2357]) | (layer2_outputs[834]);
    assign layer3_outputs[377] = ~(layer2_outputs[1164]) | (layer2_outputs[202]);
    assign layer3_outputs[378] = layer2_outputs[1315];
    assign layer3_outputs[379] = ~(layer2_outputs[1019]);
    assign layer3_outputs[380] = 1'b0;
    assign layer3_outputs[381] = layer2_outputs[372];
    assign layer3_outputs[382] = ~((layer2_outputs[1023]) ^ (layer2_outputs[2168]));
    assign layer3_outputs[383] = layer2_outputs[2041];
    assign layer3_outputs[384] = ~(layer2_outputs[1717]) | (layer2_outputs[2526]);
    assign layer3_outputs[385] = (layer2_outputs[1676]) & ~(layer2_outputs[2081]);
    assign layer3_outputs[386] = (layer2_outputs[842]) | (layer2_outputs[1921]);
    assign layer3_outputs[387] = ~(layer2_outputs[2012]) | (layer2_outputs[1333]);
    assign layer3_outputs[388] = ~((layer2_outputs[521]) | (layer2_outputs[1853]));
    assign layer3_outputs[389] = (layer2_outputs[726]) ^ (layer2_outputs[257]);
    assign layer3_outputs[390] = ~((layer2_outputs[1007]) | (layer2_outputs[2073]));
    assign layer3_outputs[391] = layer2_outputs[715];
    assign layer3_outputs[392] = ~(layer2_outputs[752]);
    assign layer3_outputs[393] = (layer2_outputs[1440]) & (layer2_outputs[754]);
    assign layer3_outputs[394] = ~(layer2_outputs[1493]);
    assign layer3_outputs[395] = ~(layer2_outputs[2461]);
    assign layer3_outputs[396] = ~(layer2_outputs[1472]) | (layer2_outputs[1612]);
    assign layer3_outputs[397] = ~(layer2_outputs[2282]);
    assign layer3_outputs[398] = layer2_outputs[397];
    assign layer3_outputs[399] = layer2_outputs[1126];
    assign layer3_outputs[400] = (layer2_outputs[753]) & ~(layer2_outputs[2547]);
    assign layer3_outputs[401] = (layer2_outputs[1671]) | (layer2_outputs[1569]);
    assign layer3_outputs[402] = ~(layer2_outputs[2009]);
    assign layer3_outputs[403] = layer2_outputs[267];
    assign layer3_outputs[404] = layer2_outputs[2535];
    assign layer3_outputs[405] = layer2_outputs[1360];
    assign layer3_outputs[406] = ~((layer2_outputs[1688]) | (layer2_outputs[1864]));
    assign layer3_outputs[407] = ~(layer2_outputs[78]) | (layer2_outputs[2201]);
    assign layer3_outputs[408] = layer2_outputs[1232];
    assign layer3_outputs[409] = ~(layer2_outputs[155]);
    assign layer3_outputs[410] = ~((layer2_outputs[1550]) | (layer2_outputs[1182]));
    assign layer3_outputs[411] = layer2_outputs[2516];
    assign layer3_outputs[412] = (layer2_outputs[1193]) | (layer2_outputs[1062]);
    assign layer3_outputs[413] = ~(layer2_outputs[824]) | (layer2_outputs[1561]);
    assign layer3_outputs[414] = (layer2_outputs[1114]) & ~(layer2_outputs[2000]);
    assign layer3_outputs[415] = layer2_outputs[1145];
    assign layer3_outputs[416] = layer2_outputs[1002];
    assign layer3_outputs[417] = ~(layer2_outputs[1784]);
    assign layer3_outputs[418] = layer2_outputs[2205];
    assign layer3_outputs[419] = ~(layer2_outputs[1394]) | (layer2_outputs[983]);
    assign layer3_outputs[420] = 1'b0;
    assign layer3_outputs[421] = layer2_outputs[2223];
    assign layer3_outputs[422] = ~((layer2_outputs[2379]) | (layer2_outputs[2142]));
    assign layer3_outputs[423] = (layer2_outputs[2479]) & ~(layer2_outputs[2281]);
    assign layer3_outputs[424] = layer2_outputs[2548];
    assign layer3_outputs[425] = (layer2_outputs[1985]) & ~(layer2_outputs[2473]);
    assign layer3_outputs[426] = 1'b1;
    assign layer3_outputs[427] = layer2_outputs[1652];
    assign layer3_outputs[428] = ~(layer2_outputs[444]) | (layer2_outputs[2010]);
    assign layer3_outputs[429] = 1'b0;
    assign layer3_outputs[430] = layer2_outputs[718];
    assign layer3_outputs[431] = (layer2_outputs[363]) ^ (layer2_outputs[695]);
    assign layer3_outputs[432] = ~(layer2_outputs[1043]);
    assign layer3_outputs[433] = ~(layer2_outputs[2529]);
    assign layer3_outputs[434] = layer2_outputs[337];
    assign layer3_outputs[435] = ~((layer2_outputs[1046]) & (layer2_outputs[1490]));
    assign layer3_outputs[436] = layer2_outputs[280];
    assign layer3_outputs[437] = (layer2_outputs[1081]) | (layer2_outputs[2248]);
    assign layer3_outputs[438] = 1'b1;
    assign layer3_outputs[439] = ~(layer2_outputs[1352]);
    assign layer3_outputs[440] = ~(layer2_outputs[2225]);
    assign layer3_outputs[441] = layer2_outputs[1303];
    assign layer3_outputs[442] = ~((layer2_outputs[2483]) & (layer2_outputs[698]));
    assign layer3_outputs[443] = layer2_outputs[230];
    assign layer3_outputs[444] = (layer2_outputs[1397]) & ~(layer2_outputs[2478]);
    assign layer3_outputs[445] = ~(layer2_outputs[344]);
    assign layer3_outputs[446] = (layer2_outputs[1000]) & ~(layer2_outputs[1766]);
    assign layer3_outputs[447] = ~(layer2_outputs[313]);
    assign layer3_outputs[448] = layer2_outputs[1118];
    assign layer3_outputs[449] = ~((layer2_outputs[2485]) ^ (layer2_outputs[740]));
    assign layer3_outputs[450] = ~(layer2_outputs[1389]);
    assign layer3_outputs[451] = layer2_outputs[2292];
    assign layer3_outputs[452] = ~(layer2_outputs[1414]);
    assign layer3_outputs[453] = (layer2_outputs[771]) & ~(layer2_outputs[772]);
    assign layer3_outputs[454] = ~((layer2_outputs[2390]) | (layer2_outputs[2214]));
    assign layer3_outputs[455] = ~(layer2_outputs[2388]);
    assign layer3_outputs[456] = (layer2_outputs[2303]) | (layer2_outputs[200]);
    assign layer3_outputs[457] = ~(layer2_outputs[333]) | (layer2_outputs[102]);
    assign layer3_outputs[458] = layer2_outputs[1947];
    assign layer3_outputs[459] = ~(layer2_outputs[2326]);
    assign layer3_outputs[460] = (layer2_outputs[1365]) | (layer2_outputs[588]);
    assign layer3_outputs[461] = (layer2_outputs[1173]) & (layer2_outputs[1912]);
    assign layer3_outputs[462] = layer2_outputs[1074];
    assign layer3_outputs[463] = ~((layer2_outputs[981]) | (layer2_outputs[2011]));
    assign layer3_outputs[464] = ~(layer2_outputs[591]);
    assign layer3_outputs[465] = ~(layer2_outputs[1730]);
    assign layer3_outputs[466] = (layer2_outputs[996]) ^ (layer2_outputs[1586]);
    assign layer3_outputs[467] = 1'b0;
    assign layer3_outputs[468] = (layer2_outputs[1579]) & (layer2_outputs[1333]);
    assign layer3_outputs[469] = ~(layer2_outputs[275]) | (layer2_outputs[1075]);
    assign layer3_outputs[470] = ~(layer2_outputs[2406]) | (layer2_outputs[1343]);
    assign layer3_outputs[471] = ~((layer2_outputs[1465]) ^ (layer2_outputs[751]));
    assign layer3_outputs[472] = ~(layer2_outputs[29]);
    assign layer3_outputs[473] = (layer2_outputs[2023]) & (layer2_outputs[1940]);
    assign layer3_outputs[474] = 1'b0;
    assign layer3_outputs[475] = ~(layer2_outputs[1361]) | (layer2_outputs[1271]);
    assign layer3_outputs[476] = ~(layer2_outputs[1184]);
    assign layer3_outputs[477] = ~(layer2_outputs[1706]) | (layer2_outputs[2145]);
    assign layer3_outputs[478] = (layer2_outputs[2184]) | (layer2_outputs[571]);
    assign layer3_outputs[479] = (layer2_outputs[1822]) & ~(layer2_outputs[23]);
    assign layer3_outputs[480] = layer2_outputs[1000];
    assign layer3_outputs[481] = (layer2_outputs[1275]) & ~(layer2_outputs[1691]);
    assign layer3_outputs[482] = ~(layer2_outputs[2338]) | (layer2_outputs[197]);
    assign layer3_outputs[483] = layer2_outputs[2230];
    assign layer3_outputs[484] = ~(layer2_outputs[949]) | (layer2_outputs[506]);
    assign layer3_outputs[485] = ~(layer2_outputs[360]);
    assign layer3_outputs[486] = ~((layer2_outputs[1192]) & (layer2_outputs[1400]));
    assign layer3_outputs[487] = (layer2_outputs[725]) | (layer2_outputs[1972]);
    assign layer3_outputs[488] = ~((layer2_outputs[1364]) ^ (layer2_outputs[1949]));
    assign layer3_outputs[489] = ~(layer2_outputs[1643]) | (layer2_outputs[835]);
    assign layer3_outputs[490] = ~(layer2_outputs[1908]);
    assign layer3_outputs[491] = (layer2_outputs[1725]) & ~(layer2_outputs[498]);
    assign layer3_outputs[492] = ~(layer2_outputs[2221]);
    assign layer3_outputs[493] = (layer2_outputs[1773]) & ~(layer2_outputs[458]);
    assign layer3_outputs[494] = layer2_outputs[2445];
    assign layer3_outputs[495] = (layer2_outputs[1519]) & (layer2_outputs[210]);
    assign layer3_outputs[496] = (layer2_outputs[1550]) ^ (layer2_outputs[1951]);
    assign layer3_outputs[497] = ~((layer2_outputs[2289]) & (layer2_outputs[798]));
    assign layer3_outputs[498] = layer2_outputs[2337];
    assign layer3_outputs[499] = ~(layer2_outputs[1361]);
    assign layer3_outputs[500] = ~((layer2_outputs[123]) & (layer2_outputs[52]));
    assign layer3_outputs[501] = layer2_outputs[1186];
    assign layer3_outputs[502] = (layer2_outputs[1237]) & (layer2_outputs[790]);
    assign layer3_outputs[503] = ~(layer2_outputs[900]);
    assign layer3_outputs[504] = layer2_outputs[755];
    assign layer3_outputs[505] = (layer2_outputs[265]) & ~(layer2_outputs[2426]);
    assign layer3_outputs[506] = ~(layer2_outputs[1396]);
    assign layer3_outputs[507] = ~(layer2_outputs[1278]);
    assign layer3_outputs[508] = ~(layer2_outputs[2278]);
    assign layer3_outputs[509] = ~((layer2_outputs[4]) & (layer2_outputs[1656]));
    assign layer3_outputs[510] = ~(layer2_outputs[2396]);
    assign layer3_outputs[511] = (layer2_outputs[2312]) & ~(layer2_outputs[610]);
    assign layer3_outputs[512] = ~((layer2_outputs[356]) | (layer2_outputs[204]));
    assign layer3_outputs[513] = layer2_outputs[1132];
    assign layer3_outputs[514] = layer2_outputs[2066];
    assign layer3_outputs[515] = (layer2_outputs[1931]) | (layer2_outputs[2273]);
    assign layer3_outputs[516] = layer2_outputs[495];
    assign layer3_outputs[517] = (layer2_outputs[488]) ^ (layer2_outputs[371]);
    assign layer3_outputs[518] = ~(layer2_outputs[2045]);
    assign layer3_outputs[519] = ~((layer2_outputs[1136]) & (layer2_outputs[998]));
    assign layer3_outputs[520] = ~(layer2_outputs[1068]) | (layer2_outputs[1055]);
    assign layer3_outputs[521] = ~(layer2_outputs[832]);
    assign layer3_outputs[522] = (layer2_outputs[1646]) & ~(layer2_outputs[904]);
    assign layer3_outputs[523] = layer2_outputs[1109];
    assign layer3_outputs[524] = layer2_outputs[203];
    assign layer3_outputs[525] = ~((layer2_outputs[599]) ^ (layer2_outputs[903]));
    assign layer3_outputs[526] = layer2_outputs[1881];
    assign layer3_outputs[527] = ~((layer2_outputs[574]) & (layer2_outputs[1055]));
    assign layer3_outputs[528] = layer2_outputs[2060];
    assign layer3_outputs[529] = ~((layer2_outputs[959]) | (layer2_outputs[6]));
    assign layer3_outputs[530] = (layer2_outputs[134]) | (layer2_outputs[1201]);
    assign layer3_outputs[531] = ~((layer2_outputs[22]) & (layer2_outputs[2033]));
    assign layer3_outputs[532] = layer2_outputs[1307];
    assign layer3_outputs[533] = layer2_outputs[1318];
    assign layer3_outputs[534] = ~(layer2_outputs[1255]) | (layer2_outputs[132]);
    assign layer3_outputs[535] = (layer2_outputs[2104]) & (layer2_outputs[2439]);
    assign layer3_outputs[536] = ~(layer2_outputs[2518]);
    assign layer3_outputs[537] = layer2_outputs[724];
    assign layer3_outputs[538] = layer2_outputs[2435];
    assign layer3_outputs[539] = 1'b0;
    assign layer3_outputs[540] = ~(layer2_outputs[1983]);
    assign layer3_outputs[541] = (layer2_outputs[223]) & ~(layer2_outputs[2191]);
    assign layer3_outputs[542] = ~(layer2_outputs[1212]);
    assign layer3_outputs[543] = ~(layer2_outputs[2117]);
    assign layer3_outputs[544] = layer2_outputs[1231];
    assign layer3_outputs[545] = ~((layer2_outputs[27]) | (layer2_outputs[479]));
    assign layer3_outputs[546] = layer2_outputs[1326];
    assign layer3_outputs[547] = ~(layer2_outputs[2512]);
    assign layer3_outputs[548] = (layer2_outputs[2118]) & (layer2_outputs[1680]);
    assign layer3_outputs[549] = 1'b1;
    assign layer3_outputs[550] = layer2_outputs[1846];
    assign layer3_outputs[551] = layer2_outputs[133];
    assign layer3_outputs[552] = ~(layer2_outputs[609]);
    assign layer3_outputs[553] = ~(layer2_outputs[596]) | (layer2_outputs[938]);
    assign layer3_outputs[554] = ~(layer2_outputs[2269]) | (layer2_outputs[1104]);
    assign layer3_outputs[555] = ~(layer2_outputs[822]);
    assign layer3_outputs[556] = (layer2_outputs[638]) & (layer2_outputs[641]);
    assign layer3_outputs[557] = (layer2_outputs[1245]) & ~(layer2_outputs[1542]);
    assign layer3_outputs[558] = ~(layer2_outputs[1235]);
    assign layer3_outputs[559] = ~(layer2_outputs[204]) | (layer2_outputs[2080]);
    assign layer3_outputs[560] = (layer2_outputs[1942]) & ~(layer2_outputs[1471]);
    assign layer3_outputs[561] = ~(layer2_outputs[455]);
    assign layer3_outputs[562] = ~(layer2_outputs[905]);
    assign layer3_outputs[563] = ~((layer2_outputs[1815]) | (layer2_outputs[2438]));
    assign layer3_outputs[564] = ~(layer2_outputs[82]);
    assign layer3_outputs[565] = ~(layer2_outputs[1372]) | (layer2_outputs[2070]);
    assign layer3_outputs[566] = ~((layer2_outputs[1001]) & (layer2_outputs[48]));
    assign layer3_outputs[567] = ~((layer2_outputs[649]) & (layer2_outputs[49]));
    assign layer3_outputs[568] = (layer2_outputs[714]) & (layer2_outputs[229]);
    assign layer3_outputs[569] = layer2_outputs[2314];
    assign layer3_outputs[570] = (layer2_outputs[1391]) & ~(layer2_outputs[428]);
    assign layer3_outputs[571] = ~(layer2_outputs[2076]);
    assign layer3_outputs[572] = ~((layer2_outputs[600]) | (layer2_outputs[404]));
    assign layer3_outputs[573] = (layer2_outputs[1132]) | (layer2_outputs[2161]);
    assign layer3_outputs[574] = ~(layer2_outputs[282]);
    assign layer3_outputs[575] = layer2_outputs[830];
    assign layer3_outputs[576] = 1'b1;
    assign layer3_outputs[577] = (layer2_outputs[701]) & ~(layer2_outputs[688]);
    assign layer3_outputs[578] = ~(layer2_outputs[63]);
    assign layer3_outputs[579] = layer2_outputs[1900];
    assign layer3_outputs[580] = ~(layer2_outputs[1573]);
    assign layer3_outputs[581] = ~(layer2_outputs[2510]) | (layer2_outputs[2159]);
    assign layer3_outputs[582] = ~(layer2_outputs[1758]) | (layer2_outputs[1099]);
    assign layer3_outputs[583] = ~(layer2_outputs[226]);
    assign layer3_outputs[584] = 1'b0;
    assign layer3_outputs[585] = ~(layer2_outputs[576]) | (layer2_outputs[2448]);
    assign layer3_outputs[586] = (layer2_outputs[1893]) ^ (layer2_outputs[837]);
    assign layer3_outputs[587] = ~(layer2_outputs[2354]) | (layer2_outputs[2074]);
    assign layer3_outputs[588] = (layer2_outputs[352]) & ~(layer2_outputs[343]);
    assign layer3_outputs[589] = ~(layer2_outputs[1350]);
    assign layer3_outputs[590] = ~(layer2_outputs[980]);
    assign layer3_outputs[591] = ~(layer2_outputs[2150]) | (layer2_outputs[1728]);
    assign layer3_outputs[592] = (layer2_outputs[206]) & ~(layer2_outputs[2369]);
    assign layer3_outputs[593] = (layer2_outputs[1645]) ^ (layer2_outputs[2096]);
    assign layer3_outputs[594] = (layer2_outputs[1699]) & (layer2_outputs[2470]);
    assign layer3_outputs[595] = (layer2_outputs[2455]) ^ (layer2_outputs[2055]);
    assign layer3_outputs[596] = (layer2_outputs[262]) ^ (layer2_outputs[1089]);
    assign layer3_outputs[597] = ~((layer2_outputs[2217]) & (layer2_outputs[2228]));
    assign layer3_outputs[598] = layer2_outputs[439];
    assign layer3_outputs[599] = ~((layer2_outputs[2116]) ^ (layer2_outputs[108]));
    assign layer3_outputs[600] = ~((layer2_outputs[1844]) | (layer2_outputs[974]));
    assign layer3_outputs[601] = ~((layer2_outputs[900]) & (layer2_outputs[2435]));
    assign layer3_outputs[602] = ~((layer2_outputs[1264]) & (layer2_outputs[349]));
    assign layer3_outputs[603] = (layer2_outputs[827]) & ~(layer2_outputs[2092]);
    assign layer3_outputs[604] = ~(layer2_outputs[2211]);
    assign layer3_outputs[605] = ~((layer2_outputs[2483]) & (layer2_outputs[187]));
    assign layer3_outputs[606] = ~(layer2_outputs[1763]);
    assign layer3_outputs[607] = ~(layer2_outputs[556]);
    assign layer3_outputs[608] = (layer2_outputs[1217]) ^ (layer2_outputs[1293]);
    assign layer3_outputs[609] = (layer2_outputs[1013]) | (layer2_outputs[380]);
    assign layer3_outputs[610] = ~((layer2_outputs[150]) ^ (layer2_outputs[307]));
    assign layer3_outputs[611] = ~((layer2_outputs[183]) | (layer2_outputs[1853]));
    assign layer3_outputs[612] = 1'b0;
    assign layer3_outputs[613] = layer2_outputs[2216];
    assign layer3_outputs[614] = (layer2_outputs[416]) & ~(layer2_outputs[2338]);
    assign layer3_outputs[615] = ~((layer2_outputs[2120]) | (layer2_outputs[1156]));
    assign layer3_outputs[616] = 1'b1;
    assign layer3_outputs[617] = ~(layer2_outputs[1061]);
    assign layer3_outputs[618] = layer2_outputs[792];
    assign layer3_outputs[619] = ~(layer2_outputs[1652]) | (layer2_outputs[1468]);
    assign layer3_outputs[620] = ~(layer2_outputs[95]);
    assign layer3_outputs[621] = (layer2_outputs[768]) | (layer2_outputs[373]);
    assign layer3_outputs[622] = (layer2_outputs[1170]) & ~(layer2_outputs[876]);
    assign layer3_outputs[623] = ~(layer2_outputs[648]);
    assign layer3_outputs[624] = (layer2_outputs[300]) & ~(layer2_outputs[1219]);
    assign layer3_outputs[625] = ~(layer2_outputs[504]);
    assign layer3_outputs[626] = ~(layer2_outputs[2266]);
    assign layer3_outputs[627] = (layer2_outputs[220]) & ~(layer2_outputs[1510]);
    assign layer3_outputs[628] = layer2_outputs[1061];
    assign layer3_outputs[629] = ~((layer2_outputs[158]) & (layer2_outputs[1070]));
    assign layer3_outputs[630] = ~(layer2_outputs[94]);
    assign layer3_outputs[631] = layer2_outputs[460];
    assign layer3_outputs[632] = 1'b0;
    assign layer3_outputs[633] = ~(layer2_outputs[1696]) | (layer2_outputs[317]);
    assign layer3_outputs[634] = ~((layer2_outputs[2545]) & (layer2_outputs[845]));
    assign layer3_outputs[635] = ~(layer2_outputs[2123]);
    assign layer3_outputs[636] = layer2_outputs[1827];
    assign layer3_outputs[637] = ~(layer2_outputs[1882]);
    assign layer3_outputs[638] = ~((layer2_outputs[318]) | (layer2_outputs[1818]));
    assign layer3_outputs[639] = ~(layer2_outputs[2343]);
    assign layer3_outputs[640] = layer2_outputs[1753];
    assign layer3_outputs[641] = (layer2_outputs[2492]) & ~(layer2_outputs[2252]);
    assign layer3_outputs[642] = ~((layer2_outputs[707]) | (layer2_outputs[765]));
    assign layer3_outputs[643] = ~(layer2_outputs[309]) | (layer2_outputs[213]);
    assign layer3_outputs[644] = ~((layer2_outputs[1103]) & (layer2_outputs[14]));
    assign layer3_outputs[645] = ~(layer2_outputs[786]);
    assign layer3_outputs[646] = (layer2_outputs[1805]) | (layer2_outputs[130]);
    assign layer3_outputs[647] = (layer2_outputs[1795]) ^ (layer2_outputs[160]);
    assign layer3_outputs[648] = ~(layer2_outputs[1805]) | (layer2_outputs[87]);
    assign layer3_outputs[649] = (layer2_outputs[140]) & (layer2_outputs[2218]);
    assign layer3_outputs[650] = ~(layer2_outputs[1111]);
    assign layer3_outputs[651] = ~((layer2_outputs[359]) ^ (layer2_outputs[1208]));
    assign layer3_outputs[652] = ~((layer2_outputs[216]) | (layer2_outputs[2022]));
    assign layer3_outputs[653] = layer2_outputs[1611];
    assign layer3_outputs[654] = (layer2_outputs[1180]) | (layer2_outputs[2256]);
    assign layer3_outputs[655] = layer2_outputs[269];
    assign layer3_outputs[656] = (layer2_outputs[2100]) ^ (layer2_outputs[1651]);
    assign layer3_outputs[657] = layer2_outputs[2493];
    assign layer3_outputs[658] = ~(layer2_outputs[1259]);
    assign layer3_outputs[659] = layer2_outputs[473];
    assign layer3_outputs[660] = (layer2_outputs[324]) & ~(layer2_outputs[154]);
    assign layer3_outputs[661] = layer2_outputs[1466];
    assign layer3_outputs[662] = layer2_outputs[232];
    assign layer3_outputs[663] = ~(layer2_outputs[168]);
    assign layer3_outputs[664] = (layer2_outputs[1920]) & ~(layer2_outputs[840]);
    assign layer3_outputs[665] = ~(layer2_outputs[334]);
    assign layer3_outputs[666] = ~((layer2_outputs[1743]) & (layer2_outputs[2065]));
    assign layer3_outputs[667] = (layer2_outputs[1294]) | (layer2_outputs[2519]);
    assign layer3_outputs[668] = 1'b0;
    assign layer3_outputs[669] = ~(layer2_outputs[315]) | (layer2_outputs[1227]);
    assign layer3_outputs[670] = ~((layer2_outputs[0]) | (layer2_outputs[892]));
    assign layer3_outputs[671] = ~(layer2_outputs[964]);
    assign layer3_outputs[672] = ~(layer2_outputs[2539]) | (layer2_outputs[1704]);
    assign layer3_outputs[673] = layer2_outputs[279];
    assign layer3_outputs[674] = ~(layer2_outputs[1353]);
    assign layer3_outputs[675] = ~((layer2_outputs[1721]) | (layer2_outputs[1080]));
    assign layer3_outputs[676] = ~(layer2_outputs[2333]);
    assign layer3_outputs[677] = (layer2_outputs[2280]) | (layer2_outputs[1417]);
    assign layer3_outputs[678] = ~(layer2_outputs[750]) | (layer2_outputs[549]);
    assign layer3_outputs[679] = ~(layer2_outputs[1754]);
    assign layer3_outputs[680] = 1'b1;
    assign layer3_outputs[681] = ~(layer2_outputs[2532]) | (layer2_outputs[48]);
    assign layer3_outputs[682] = ~(layer2_outputs[2437]);
    assign layer3_outputs[683] = ~((layer2_outputs[301]) & (layer2_outputs[1927]));
    assign layer3_outputs[684] = (layer2_outputs[1153]) ^ (layer2_outputs[2365]);
    assign layer3_outputs[685] = layer2_outputs[2138];
    assign layer3_outputs[686] = (layer2_outputs[2355]) & ~(layer2_outputs[863]);
    assign layer3_outputs[687] = layer2_outputs[718];
    assign layer3_outputs[688] = ~(layer2_outputs[138]);
    assign layer3_outputs[689] = ~(layer2_outputs[1878]) | (layer2_outputs[630]);
    assign layer3_outputs[690] = ~(layer2_outputs[1733]);
    assign layer3_outputs[691] = (layer2_outputs[1091]) & (layer2_outputs[861]);
    assign layer3_outputs[692] = ~(layer2_outputs[2275]);
    assign layer3_outputs[693] = layer2_outputs[131];
    assign layer3_outputs[694] = (layer2_outputs[1229]) ^ (layer2_outputs[1040]);
    assign layer3_outputs[695] = (layer2_outputs[548]) & (layer2_outputs[2127]);
    assign layer3_outputs[696] = ~(layer2_outputs[511]) | (layer2_outputs[391]);
    assign layer3_outputs[697] = (layer2_outputs[1459]) & ~(layer2_outputs[256]);
    assign layer3_outputs[698] = layer2_outputs[142];
    assign layer3_outputs[699] = layer2_outputs[2460];
    assign layer3_outputs[700] = layer2_outputs[147];
    assign layer3_outputs[701] = (layer2_outputs[474]) ^ (layer2_outputs[1018]);
    assign layer3_outputs[702] = ~(layer2_outputs[1011]) | (layer2_outputs[486]);
    assign layer3_outputs[703] = ~(layer2_outputs[577]);
    assign layer3_outputs[704] = ~(layer2_outputs[1277]);
    assign layer3_outputs[705] = ~(layer2_outputs[2228]);
    assign layer3_outputs[706] = 1'b1;
    assign layer3_outputs[707] = ~(layer2_outputs[422]);
    assign layer3_outputs[708] = ~(layer2_outputs[2178]);
    assign layer3_outputs[709] = (layer2_outputs[57]) & ~(layer2_outputs[1270]);
    assign layer3_outputs[710] = (layer2_outputs[1351]) | (layer2_outputs[634]);
    assign layer3_outputs[711] = layer2_outputs[1187];
    assign layer3_outputs[712] = layer2_outputs[2081];
    assign layer3_outputs[713] = layer2_outputs[1555];
    assign layer3_outputs[714] = ~(layer2_outputs[971]) | (layer2_outputs[1821]);
    assign layer3_outputs[715] = ~(layer2_outputs[109]);
    assign layer3_outputs[716] = (layer2_outputs[1284]) & ~(layer2_outputs[535]);
    assign layer3_outputs[717] = ~(layer2_outputs[91]);
    assign layer3_outputs[718] = ~(layer2_outputs[2296]);
    assign layer3_outputs[719] = layer2_outputs[452];
    assign layer3_outputs[720] = (layer2_outputs[1214]) & (layer2_outputs[1799]);
    assign layer3_outputs[721] = (layer2_outputs[740]) & (layer2_outputs[1899]);
    assign layer3_outputs[722] = (layer2_outputs[984]) & ~(layer2_outputs[2289]);
    assign layer3_outputs[723] = ~(layer2_outputs[1310]) | (layer2_outputs[3]);
    assign layer3_outputs[724] = ~((layer2_outputs[1077]) | (layer2_outputs[2295]));
    assign layer3_outputs[725] = (layer2_outputs[1662]) | (layer2_outputs[1630]);
    assign layer3_outputs[726] = 1'b0;
    assign layer3_outputs[727] = 1'b1;
    assign layer3_outputs[728] = layer2_outputs[1098];
    assign layer3_outputs[729] = (layer2_outputs[1295]) | (layer2_outputs[896]);
    assign layer3_outputs[730] = (layer2_outputs[167]) | (layer2_outputs[84]);
    assign layer3_outputs[731] = (layer2_outputs[616]) ^ (layer2_outputs[283]);
    assign layer3_outputs[732] = layer2_outputs[175];
    assign layer3_outputs[733] = (layer2_outputs[340]) & (layer2_outputs[979]);
    assign layer3_outputs[734] = ~(layer2_outputs[1988]);
    assign layer3_outputs[735] = layer2_outputs[1166];
    assign layer3_outputs[736] = (layer2_outputs[2205]) & ~(layer2_outputs[1644]);
    assign layer3_outputs[737] = (layer2_outputs[1677]) | (layer2_outputs[475]);
    assign layer3_outputs[738] = ~((layer2_outputs[1679]) & (layer2_outputs[2370]));
    assign layer3_outputs[739] = (layer2_outputs[815]) & (layer2_outputs[472]);
    assign layer3_outputs[740] = ~(layer2_outputs[991]) | (layer2_outputs[1916]);
    assign layer3_outputs[741] = ~(layer2_outputs[1420]);
    assign layer3_outputs[742] = ~(layer2_outputs[1530]) | (layer2_outputs[1069]);
    assign layer3_outputs[743] = 1'b1;
    assign layer3_outputs[744] = (layer2_outputs[2418]) & ~(layer2_outputs[2300]);
    assign layer3_outputs[745] = layer2_outputs[916];
    assign layer3_outputs[746] = 1'b0;
    assign layer3_outputs[747] = (layer2_outputs[260]) & (layer2_outputs[2494]);
    assign layer3_outputs[748] = ~(layer2_outputs[796]);
    assign layer3_outputs[749] = ~((layer2_outputs[2257]) & (layer2_outputs[930]));
    assign layer3_outputs[750] = layer2_outputs[2496];
    assign layer3_outputs[751] = (layer2_outputs[2337]) & (layer2_outputs[618]);
    assign layer3_outputs[752] = layer2_outputs[240];
    assign layer3_outputs[753] = ~(layer2_outputs[1549]);
    assign layer3_outputs[754] = (layer2_outputs[1914]) ^ (layer2_outputs[1531]);
    assign layer3_outputs[755] = ~(layer2_outputs[194]);
    assign layer3_outputs[756] = layer2_outputs[1206];
    assign layer3_outputs[757] = (layer2_outputs[2275]) & (layer2_outputs[2366]);
    assign layer3_outputs[758] = (layer2_outputs[1973]) & ~(layer2_outputs[935]);
    assign layer3_outputs[759] = layer2_outputs[240];
    assign layer3_outputs[760] = layer2_outputs[1261];
    assign layer3_outputs[761] = ~(layer2_outputs[2442]);
    assign layer3_outputs[762] = layer2_outputs[241];
    assign layer3_outputs[763] = ~(layer2_outputs[406]);
    assign layer3_outputs[764] = layer2_outputs[2158];
    assign layer3_outputs[765] = ~(layer2_outputs[1670]) | (layer2_outputs[689]);
    assign layer3_outputs[766] = layer2_outputs[1708];
    assign layer3_outputs[767] = layer2_outputs[172];
    assign layer3_outputs[768] = ~(layer2_outputs[176]);
    assign layer3_outputs[769] = layer2_outputs[39];
    assign layer3_outputs[770] = ~(layer2_outputs[224]) | (layer2_outputs[1811]);
    assign layer3_outputs[771] = (layer2_outputs[32]) ^ (layer2_outputs[1516]);
    assign layer3_outputs[772] = ~(layer2_outputs[2449]) | (layer2_outputs[1677]);
    assign layer3_outputs[773] = layer2_outputs[1198];
    assign layer3_outputs[774] = ~(layer2_outputs[1469]);
    assign layer3_outputs[775] = (layer2_outputs[2452]) | (layer2_outputs[1392]);
    assign layer3_outputs[776] = (layer2_outputs[2133]) ^ (layer2_outputs[1003]);
    assign layer3_outputs[777] = (layer2_outputs[1058]) & ~(layer2_outputs[2038]);
    assign layer3_outputs[778] = ~(layer2_outputs[151]);
    assign layer3_outputs[779] = ~(layer2_outputs[443]);
    assign layer3_outputs[780] = (layer2_outputs[1880]) & (layer2_outputs[105]);
    assign layer3_outputs[781] = ~(layer2_outputs[2310]);
    assign layer3_outputs[782] = layer2_outputs[563];
    assign layer3_outputs[783] = (layer2_outputs[2326]) & ~(layer2_outputs[2403]);
    assign layer3_outputs[784] = ~(layer2_outputs[1290]);
    assign layer3_outputs[785] = ~((layer2_outputs[2202]) & (layer2_outputs[1511]));
    assign layer3_outputs[786] = 1'b1;
    assign layer3_outputs[787] = (layer2_outputs[2132]) & ~(layer2_outputs[712]);
    assign layer3_outputs[788] = ~(layer2_outputs[2177]);
    assign layer3_outputs[789] = ~((layer2_outputs[1133]) & (layer2_outputs[1620]));
    assign layer3_outputs[790] = (layer2_outputs[1874]) & (layer2_outputs[852]);
    assign layer3_outputs[791] = (layer2_outputs[1296]) ^ (layer2_outputs[1144]);
    assign layer3_outputs[792] = (layer2_outputs[428]) & (layer2_outputs[970]);
    assign layer3_outputs[793] = layer2_outputs[593];
    assign layer3_outputs[794] = 1'b0;
    assign layer3_outputs[795] = (layer2_outputs[130]) & (layer2_outputs[476]);
    assign layer3_outputs[796] = ~((layer2_outputs[374]) | (layer2_outputs[1086]));
    assign layer3_outputs[797] = ~(layer2_outputs[1207]) | (layer2_outputs[1373]);
    assign layer3_outputs[798] = ~(layer2_outputs[93]);
    assign layer3_outputs[799] = ~(layer2_outputs[2325]) | (layer2_outputs[1377]);
    assign layer3_outputs[800] = (layer2_outputs[1722]) ^ (layer2_outputs[1915]);
    assign layer3_outputs[801] = (layer2_outputs[1270]) | (layer2_outputs[722]);
    assign layer3_outputs[802] = (layer2_outputs[31]) & ~(layer2_outputs[1425]);
    assign layer3_outputs[803] = ~(layer2_outputs[1725]) | (layer2_outputs[2313]);
    assign layer3_outputs[804] = layer2_outputs[1276];
    assign layer3_outputs[805] = (layer2_outputs[1797]) & ~(layer2_outputs[1997]);
    assign layer3_outputs[806] = ~(layer2_outputs[377]);
    assign layer3_outputs[807] = (layer2_outputs[1101]) & ~(layer2_outputs[943]);
    assign layer3_outputs[808] = (layer2_outputs[1014]) & (layer2_outputs[2274]);
    assign layer3_outputs[809] = ~(layer2_outputs[1844]) | (layer2_outputs[1840]);
    assign layer3_outputs[810] = layer2_outputs[1956];
    assign layer3_outputs[811] = 1'b1;
    assign layer3_outputs[812] = ~(layer2_outputs[259]);
    assign layer3_outputs[813] = ~(layer2_outputs[643]);
    assign layer3_outputs[814] = ~((layer2_outputs[71]) ^ (layer2_outputs[2127]));
    assign layer3_outputs[815] = layer2_outputs[12];
    assign layer3_outputs[816] = ~(layer2_outputs[1735]);
    assign layer3_outputs[817] = (layer2_outputs[230]) & ~(layer2_outputs[1628]);
    assign layer3_outputs[818] = ~(layer2_outputs[237]);
    assign layer3_outputs[819] = ~(layer2_outputs[2436]);
    assign layer3_outputs[820] = (layer2_outputs[1892]) & ~(layer2_outputs[1251]);
    assign layer3_outputs[821] = 1'b1;
    assign layer3_outputs[822] = ~(layer2_outputs[2538]);
    assign layer3_outputs[823] = 1'b0;
    assign layer3_outputs[824] = ~(layer2_outputs[238]) | (layer2_outputs[1575]);
    assign layer3_outputs[825] = layer2_outputs[978];
    assign layer3_outputs[826] = layer2_outputs[1734];
    assign layer3_outputs[827] = 1'b1;
    assign layer3_outputs[828] = ~((layer2_outputs[1232]) & (layer2_outputs[500]));
    assign layer3_outputs[829] = ~(layer2_outputs[2209]);
    assign layer3_outputs[830] = (layer2_outputs[192]) & ~(layer2_outputs[1744]);
    assign layer3_outputs[831] = ~(layer2_outputs[485]);
    assign layer3_outputs[832] = layer2_outputs[1483];
    assign layer3_outputs[833] = ~(layer2_outputs[2079]);
    assign layer3_outputs[834] = ~(layer2_outputs[827]) | (layer2_outputs[426]);
    assign layer3_outputs[835] = ~((layer2_outputs[633]) & (layer2_outputs[1611]));
    assign layer3_outputs[836] = ~(layer2_outputs[1771]);
    assign layer3_outputs[837] = layer2_outputs[2321];
    assign layer3_outputs[838] = layer2_outputs[1393];
    assign layer3_outputs[839] = layer2_outputs[1258];
    assign layer3_outputs[840] = layer2_outputs[1116];
    assign layer3_outputs[841] = layer2_outputs[1059];
    assign layer3_outputs[842] = (layer2_outputs[274]) & ~(layer2_outputs[1439]);
    assign layer3_outputs[843] = ~(layer2_outputs[198]);
    assign layer3_outputs[844] = ~(layer2_outputs[263]);
    assign layer3_outputs[845] = ~(layer2_outputs[1372]);
    assign layer3_outputs[846] = layer2_outputs[2533];
    assign layer3_outputs[847] = ~((layer2_outputs[1817]) ^ (layer2_outputs[1337]));
    assign layer3_outputs[848] = ~(layer2_outputs[1933]);
    assign layer3_outputs[849] = ~(layer2_outputs[1870]);
    assign layer3_outputs[850] = ~(layer2_outputs[1418]);
    assign layer3_outputs[851] = (layer2_outputs[314]) & ~(layer2_outputs[2110]);
    assign layer3_outputs[852] = layer2_outputs[2192];
    assign layer3_outputs[853] = (layer2_outputs[410]) & ~(layer2_outputs[1987]);
    assign layer3_outputs[854] = ~((layer2_outputs[2305]) | (layer2_outputs[1487]));
    assign layer3_outputs[855] = layer2_outputs[2189];
    assign layer3_outputs[856] = ~(layer2_outputs[1757]);
    assign layer3_outputs[857] = ~((layer2_outputs[500]) ^ (layer2_outputs[1442]));
    assign layer3_outputs[858] = ~((layer2_outputs[296]) & (layer2_outputs[979]));
    assign layer3_outputs[859] = layer2_outputs[2520];
    assign layer3_outputs[860] = ~(layer2_outputs[598]);
    assign layer3_outputs[861] = ~(layer2_outputs[2144]);
    assign layer3_outputs[862] = ~(layer2_outputs[837]) | (layer2_outputs[955]);
    assign layer3_outputs[863] = ~((layer2_outputs[2140]) & (layer2_outputs[237]));
    assign layer3_outputs[864] = ~((layer2_outputs[1115]) & (layer2_outputs[45]));
    assign layer3_outputs[865] = layer2_outputs[688];
    assign layer3_outputs[866] = layer2_outputs[2067];
    assign layer3_outputs[867] = ~(layer2_outputs[1072]);
    assign layer3_outputs[868] = ~((layer2_outputs[685]) | (layer2_outputs[978]));
    assign layer3_outputs[869] = ~(layer2_outputs[1195]) | (layer2_outputs[2222]);
    assign layer3_outputs[870] = layer2_outputs[600];
    assign layer3_outputs[871] = layer2_outputs[755];
    assign layer3_outputs[872] = (layer2_outputs[1575]) & ~(layer2_outputs[1101]);
    assign layer3_outputs[873] = ~((layer2_outputs[342]) ^ (layer2_outputs[76]));
    assign layer3_outputs[874] = (layer2_outputs[994]) & ~(layer2_outputs[1322]);
    assign layer3_outputs[875] = (layer2_outputs[1009]) & ~(layer2_outputs[1131]);
    assign layer3_outputs[876] = ~(layer2_outputs[2187]) | (layer2_outputs[384]);
    assign layer3_outputs[877] = 1'b0;
    assign layer3_outputs[878] = layer2_outputs[1037];
    assign layer3_outputs[879] = (layer2_outputs[992]) & (layer2_outputs[2083]);
    assign layer3_outputs[880] = ~(layer2_outputs[729]);
    assign layer3_outputs[881] = ~(layer2_outputs[1491]) | (layer2_outputs[116]);
    assign layer3_outputs[882] = ~((layer2_outputs[932]) & (layer2_outputs[1481]));
    assign layer3_outputs[883] = 1'b1;
    assign layer3_outputs[884] = (layer2_outputs[1625]) & ~(layer2_outputs[1639]);
    assign layer3_outputs[885] = ~((layer2_outputs[19]) & (layer2_outputs[1675]));
    assign layer3_outputs[886] = ~(layer2_outputs[2236]);
    assign layer3_outputs[887] = (layer2_outputs[2099]) & ~(layer2_outputs[1936]);
    assign layer3_outputs[888] = ~(layer2_outputs[281]);
    assign layer3_outputs[889] = ~(layer2_outputs[1516]);
    assign layer3_outputs[890] = layer2_outputs[1446];
    assign layer3_outputs[891] = (layer2_outputs[2103]) & (layer2_outputs[2420]);
    assign layer3_outputs[892] = (layer2_outputs[1437]) & ~(layer2_outputs[1312]);
    assign layer3_outputs[893] = (layer2_outputs[490]) & (layer2_outputs[1961]);
    assign layer3_outputs[894] = (layer2_outputs[519]) & ~(layer2_outputs[400]);
    assign layer3_outputs[895] = ~(layer2_outputs[1225]);
    assign layer3_outputs[896] = ~(layer2_outputs[1767]);
    assign layer3_outputs[897] = (layer2_outputs[690]) & ~(layer2_outputs[927]);
    assign layer3_outputs[898] = ~(layer2_outputs[2444]) | (layer2_outputs[1896]);
    assign layer3_outputs[899] = (layer2_outputs[161]) | (layer2_outputs[556]);
    assign layer3_outputs[900] = ~(layer2_outputs[93]);
    assign layer3_outputs[901] = layer2_outputs[2448];
    assign layer3_outputs[902] = ~(layer2_outputs[2036]);
    assign layer3_outputs[903] = ~(layer2_outputs[1167]) | (layer2_outputs[873]);
    assign layer3_outputs[904] = (layer2_outputs[325]) ^ (layer2_outputs[397]);
    assign layer3_outputs[905] = ~(layer2_outputs[2197]);
    assign layer3_outputs[906] = (layer2_outputs[1398]) | (layer2_outputs[2165]);
    assign layer3_outputs[907] = ~(layer2_outputs[2186]) | (layer2_outputs[299]);
    assign layer3_outputs[908] = (layer2_outputs[1946]) | (layer2_outputs[2469]);
    assign layer3_outputs[909] = ~(layer2_outputs[2017]) | (layer2_outputs[423]);
    assign layer3_outputs[910] = ~(layer2_outputs[2185]);
    assign layer3_outputs[911] = layer2_outputs[2070];
    assign layer3_outputs[912] = (layer2_outputs[2405]) & (layer2_outputs[1657]);
    assign layer3_outputs[913] = (layer2_outputs[1783]) ^ (layer2_outputs[2384]);
    assign layer3_outputs[914] = (layer2_outputs[396]) & ~(layer2_outputs[1016]);
    assign layer3_outputs[915] = ~(layer2_outputs[1772]);
    assign layer3_outputs[916] = ~(layer2_outputs[2333]) | (layer2_outputs[803]);
    assign layer3_outputs[917] = (layer2_outputs[152]) & ~(layer2_outputs[577]);
    assign layer3_outputs[918] = layer2_outputs[2408];
    assign layer3_outputs[919] = (layer2_outputs[1804]) & ~(layer2_outputs[250]);
    assign layer3_outputs[920] = ~(layer2_outputs[295]) | (layer2_outputs[214]);
    assign layer3_outputs[921] = (layer2_outputs[1971]) & ~(layer2_outputs[1274]);
    assign layer3_outputs[922] = ~((layer2_outputs[180]) ^ (layer2_outputs[2534]));
    assign layer3_outputs[923] = ~((layer2_outputs[457]) ^ (layer2_outputs[1215]));
    assign layer3_outputs[924] = ~((layer2_outputs[460]) ^ (layer2_outputs[209]));
    assign layer3_outputs[925] = ~((layer2_outputs[2113]) | (layer2_outputs[1751]));
    assign layer3_outputs[926] = ~(layer2_outputs[514]) | (layer2_outputs[2537]);
    assign layer3_outputs[927] = 1'b0;
    assign layer3_outputs[928] = ~(layer2_outputs[209]);
    assign layer3_outputs[929] = (layer2_outputs[1213]) & ~(layer2_outputs[2478]);
    assign layer3_outputs[930] = ~(layer2_outputs[2278]);
    assign layer3_outputs[931] = layer2_outputs[410];
    assign layer3_outputs[932] = 1'b0;
    assign layer3_outputs[933] = (layer2_outputs[1353]) | (layer2_outputs[1202]);
    assign layer3_outputs[934] = layer2_outputs[378];
    assign layer3_outputs[935] = ~(layer2_outputs[1402]);
    assign layer3_outputs[936] = 1'b1;
    assign layer3_outputs[937] = (layer2_outputs[2148]) & (layer2_outputs[1995]);
    assign layer3_outputs[938] = ~((layer2_outputs[314]) ^ (layer2_outputs[1154]));
    assign layer3_outputs[939] = (layer2_outputs[115]) & ~(layer2_outputs[522]);
    assign layer3_outputs[940] = ~((layer2_outputs[847]) | (layer2_outputs[1861]));
    assign layer3_outputs[941] = ~((layer2_outputs[2458]) & (layer2_outputs[1509]));
    assign layer3_outputs[942] = layer2_outputs[2369];
    assign layer3_outputs[943] = ~((layer2_outputs[2182]) & (layer2_outputs[1477]));
    assign layer3_outputs[944] = (layer2_outputs[1755]) & ~(layer2_outputs[244]);
    assign layer3_outputs[945] = ~(layer2_outputs[2414]) | (layer2_outputs[608]);
    assign layer3_outputs[946] = layer2_outputs[1928];
    assign layer3_outputs[947] = layer2_outputs[512];
    assign layer3_outputs[948] = (layer2_outputs[1778]) | (layer2_outputs[2482]);
    assign layer3_outputs[949] = ~((layer2_outputs[2175]) | (layer2_outputs[1564]));
    assign layer3_outputs[950] = ~(layer2_outputs[167]) | (layer2_outputs[1419]);
    assign layer3_outputs[951] = layer2_outputs[343];
    assign layer3_outputs[952] = layer2_outputs[2196];
    assign layer3_outputs[953] = (layer2_outputs[1706]) & ~(layer2_outputs[1120]);
    assign layer3_outputs[954] = layer2_outputs[2557];
    assign layer3_outputs[955] = ~(layer2_outputs[1892]);
    assign layer3_outputs[956] = ~(layer2_outputs[568]) | (layer2_outputs[421]);
    assign layer3_outputs[957] = ~((layer2_outputs[259]) | (layer2_outputs[1816]));
    assign layer3_outputs[958] = 1'b1;
    assign layer3_outputs[959] = ~((layer2_outputs[1979]) & (layer2_outputs[1573]));
    assign layer3_outputs[960] = ~((layer2_outputs[717]) | (layer2_outputs[1513]));
    assign layer3_outputs[961] = layer2_outputs[2358];
    assign layer3_outputs[962] = ~(layer2_outputs[2256]) | (layer2_outputs[1140]);
    assign layer3_outputs[963] = layer2_outputs[201];
    assign layer3_outputs[964] = layer2_outputs[1828];
    assign layer3_outputs[965] = ~((layer2_outputs[1107]) & (layer2_outputs[2157]));
    assign layer3_outputs[966] = ~((layer2_outputs[2394]) | (layer2_outputs[2320]));
    assign layer3_outputs[967] = layer2_outputs[1870];
    assign layer3_outputs[968] = ~(layer2_outputs[1811]);
    assign layer3_outputs[969] = ~(layer2_outputs[1208]);
    assign layer3_outputs[970] = ~((layer2_outputs[1910]) & (layer2_outputs[1041]));
    assign layer3_outputs[971] = (layer2_outputs[716]) & ~(layer2_outputs[2433]);
    assign layer3_outputs[972] = (layer2_outputs[221]) & ~(layer2_outputs[2290]);
    assign layer3_outputs[973] = layer2_outputs[405];
    assign layer3_outputs[974] = (layer2_outputs[217]) | (layer2_outputs[698]);
    assign layer3_outputs[975] = layer2_outputs[1855];
    assign layer3_outputs[976] = ~(layer2_outputs[1493]);
    assign layer3_outputs[977] = ~(layer2_outputs[1212]);
    assign layer3_outputs[978] = layer2_outputs[2351];
    assign layer3_outputs[979] = ~(layer2_outputs[1120]);
    assign layer3_outputs[980] = ~((layer2_outputs[128]) & (layer2_outputs[849]));
    assign layer3_outputs[981] = ~((layer2_outputs[1374]) | (layer2_outputs[2548]));
    assign layer3_outputs[982] = ~(layer2_outputs[1108]);
    assign layer3_outputs[983] = layer2_outputs[2536];
    assign layer3_outputs[984] = (layer2_outputs[356]) & ~(layer2_outputs[1845]);
    assign layer3_outputs[985] = 1'b1;
    assign layer3_outputs[986] = ~((layer2_outputs[647]) & (layer2_outputs[67]));
    assign layer3_outputs[987] = ~(layer2_outputs[2253]) | (layer2_outputs[1458]);
    assign layer3_outputs[988] = layer2_outputs[560];
    assign layer3_outputs[989] = (layer2_outputs[2146]) & (layer2_outputs[28]);
    assign layer3_outputs[990] = (layer2_outputs[1901]) & ~(layer2_outputs[1877]);
    assign layer3_outputs[991] = ~(layer2_outputs[2130]);
    assign layer3_outputs[992] = 1'b0;
    assign layer3_outputs[993] = ~(layer2_outputs[1765]);
    assign layer3_outputs[994] = (layer2_outputs[1518]) & ~(layer2_outputs[507]);
    assign layer3_outputs[995] = ~((layer2_outputs[24]) & (layer2_outputs[1537]));
    assign layer3_outputs[996] = (layer2_outputs[1221]) & ~(layer2_outputs[2537]);
    assign layer3_outputs[997] = ~(layer2_outputs[1702]);
    assign layer3_outputs[998] = (layer2_outputs[525]) | (layer2_outputs[1924]);
    assign layer3_outputs[999] = (layer2_outputs[928]) & (layer2_outputs[68]);
    assign layer3_outputs[1000] = ~(layer2_outputs[1360]);
    assign layer3_outputs[1001] = layer2_outputs[564];
    assign layer3_outputs[1002] = 1'b0;
    assign layer3_outputs[1003] = layer2_outputs[798];
    assign layer3_outputs[1004] = ~(layer2_outputs[721]);
    assign layer3_outputs[1005] = layer2_outputs[1084];
    assign layer3_outputs[1006] = layer2_outputs[2220];
    assign layer3_outputs[1007] = ~((layer2_outputs[2025]) & (layer2_outputs[1991]));
    assign layer3_outputs[1008] = layer2_outputs[1655];
    assign layer3_outputs[1009] = (layer2_outputs[273]) & ~(layer2_outputs[1638]);
    assign layer3_outputs[1010] = ~(layer2_outputs[2143]) | (layer2_outputs[1793]);
    assign layer3_outputs[1011] = layer2_outputs[177];
    assign layer3_outputs[1012] = layer2_outputs[2048];
    assign layer3_outputs[1013] = layer2_outputs[805];
    assign layer3_outputs[1014] = 1'b0;
    assign layer3_outputs[1015] = layer2_outputs[2055];
    assign layer3_outputs[1016] = layer2_outputs[2178];
    assign layer3_outputs[1017] = (layer2_outputs[330]) ^ (layer2_outputs[1124]);
    assign layer3_outputs[1018] = ~(layer2_outputs[2419]) | (layer2_outputs[1877]);
    assign layer3_outputs[1019] = ~(layer2_outputs[119]);
    assign layer3_outputs[1020] = layer2_outputs[1926];
    assign layer3_outputs[1021] = (layer2_outputs[21]) ^ (layer2_outputs[557]);
    assign layer3_outputs[1022] = (layer2_outputs[1324]) & ~(layer2_outputs[802]);
    assign layer3_outputs[1023] = (layer2_outputs[2508]) & ~(layer2_outputs[121]);
    assign layer3_outputs[1024] = layer2_outputs[1661];
    assign layer3_outputs[1025] = ~(layer2_outputs[1982]);
    assign layer3_outputs[1026] = ~(layer2_outputs[387]) | (layer2_outputs[940]);
    assign layer3_outputs[1027] = layer2_outputs[1244];
    assign layer3_outputs[1028] = (layer2_outputs[417]) & ~(layer2_outputs[2391]);
    assign layer3_outputs[1029] = ~((layer2_outputs[1975]) | (layer2_outputs[1542]));
    assign layer3_outputs[1030] = (layer2_outputs[898]) & ~(layer2_outputs[1964]);
    assign layer3_outputs[1031] = ~((layer2_outputs[1406]) ^ (layer2_outputs[497]));
    assign layer3_outputs[1032] = ~(layer2_outputs[618]);
    assign layer3_outputs[1033] = layer2_outputs[1267];
    assign layer3_outputs[1034] = ~((layer2_outputs[1630]) ^ (layer2_outputs[227]));
    assign layer3_outputs[1035] = ~((layer2_outputs[182]) & (layer2_outputs[1028]));
    assign layer3_outputs[1036] = (layer2_outputs[2404]) & ~(layer2_outputs[799]);
    assign layer3_outputs[1037] = ~((layer2_outputs[981]) | (layer2_outputs[2545]));
    assign layer3_outputs[1038] = ~(layer2_outputs[1258]);
    assign layer3_outputs[1039] = ~(layer2_outputs[453]);
    assign layer3_outputs[1040] = ~(layer2_outputs[2188]);
    assign layer3_outputs[1041] = (layer2_outputs[2540]) | (layer2_outputs[838]);
    assign layer3_outputs[1042] = layer2_outputs[1247];
    assign layer3_outputs[1043] = (layer2_outputs[7]) | (layer2_outputs[1183]);
    assign layer3_outputs[1044] = (layer2_outputs[1045]) & ~(layer2_outputs[602]);
    assign layer3_outputs[1045] = 1'b1;
    assign layer3_outputs[1046] = 1'b1;
    assign layer3_outputs[1047] = layer2_outputs[1292];
    assign layer3_outputs[1048] = ~(layer2_outputs[860]);
    assign layer3_outputs[1049] = 1'b0;
    assign layer3_outputs[1050] = (layer2_outputs[1153]) | (layer2_outputs[1135]);
    assign layer3_outputs[1051] = ~(layer2_outputs[262]);
    assign layer3_outputs[1052] = (layer2_outputs[2522]) & (layer2_outputs[559]);
    assign layer3_outputs[1053] = (layer2_outputs[1661]) ^ (layer2_outputs[1205]);
    assign layer3_outputs[1054] = ~(layer2_outputs[1957]);
    assign layer3_outputs[1055] = layer2_outputs[2377];
    assign layer3_outputs[1056] = 1'b1;
    assign layer3_outputs[1057] = ~(layer2_outputs[853]) | (layer2_outputs[998]);
    assign layer3_outputs[1058] = layer2_outputs[1965];
    assign layer3_outputs[1059] = layer2_outputs[293];
    assign layer3_outputs[1060] = (layer2_outputs[2503]) & (layer2_outputs[261]);
    assign layer3_outputs[1061] = layer2_outputs[1943];
    assign layer3_outputs[1062] = ~(layer2_outputs[335]) | (layer2_outputs[424]);
    assign layer3_outputs[1063] = ~((layer2_outputs[1872]) | (layer2_outputs[1221]));
    assign layer3_outputs[1064] = layer2_outputs[956];
    assign layer3_outputs[1065] = 1'b0;
    assign layer3_outputs[1066] = ~((layer2_outputs[951]) & (layer2_outputs[956]));
    assign layer3_outputs[1067] = layer2_outputs[2254];
    assign layer3_outputs[1068] = ~((layer2_outputs[2238]) & (layer2_outputs[468]));
    assign layer3_outputs[1069] = layer2_outputs[530];
    assign layer3_outputs[1070] = (layer2_outputs[2008]) & ~(layer2_outputs[2003]);
    assign layer3_outputs[1071] = layer2_outputs[54];
    assign layer3_outputs[1072] = ~((layer2_outputs[171]) & (layer2_outputs[2286]));
    assign layer3_outputs[1073] = (layer2_outputs[685]) | (layer2_outputs[2385]);
    assign layer3_outputs[1074] = ~(layer2_outputs[1664]);
    assign layer3_outputs[1075] = ~(layer2_outputs[377]);
    assign layer3_outputs[1076] = layer2_outputs[1764];
    assign layer3_outputs[1077] = (layer2_outputs[1679]) | (layer2_outputs[974]);
    assign layer3_outputs[1078] = ~(layer2_outputs[921]);
    assign layer3_outputs[1079] = 1'b0;
    assign layer3_outputs[1080] = layer2_outputs[843];
    assign layer3_outputs[1081] = (layer2_outputs[1294]) & ~(layer2_outputs[1909]);
    assign layer3_outputs[1082] = layer2_outputs[1157];
    assign layer3_outputs[1083] = (layer2_outputs[1847]) & ~(layer2_outputs[1560]);
    assign layer3_outputs[1084] = layer2_outputs[2301];
    assign layer3_outputs[1085] = layer2_outputs[1809];
    assign layer3_outputs[1086] = (layer2_outputs[1311]) & ~(layer2_outputs[406]);
    assign layer3_outputs[1087] = ~((layer2_outputs[1535]) ^ (layer2_outputs[1667]));
    assign layer3_outputs[1088] = ~(layer2_outputs[831]) | (layer2_outputs[834]);
    assign layer3_outputs[1089] = ~(layer2_outputs[2299]);
    assign layer3_outputs[1090] = 1'b0;
    assign layer3_outputs[1091] = (layer2_outputs[2209]) | (layer2_outputs[1672]);
    assign layer3_outputs[1092] = ~((layer2_outputs[1328]) | (layer2_outputs[648]));
    assign layer3_outputs[1093] = ~(layer2_outputs[2046]) | (layer2_outputs[1354]);
    assign layer3_outputs[1094] = (layer2_outputs[2419]) & (layer2_outputs[939]);
    assign layer3_outputs[1095] = (layer2_outputs[261]) & ~(layer2_outputs[1241]);
    assign layer3_outputs[1096] = ~(layer2_outputs[1781]) | (layer2_outputs[2108]);
    assign layer3_outputs[1097] = (layer2_outputs[1482]) | (layer2_outputs[825]);
    assign layer3_outputs[1098] = ~(layer2_outputs[1497]);
    assign layer3_outputs[1099] = ~((layer2_outputs[2293]) & (layer2_outputs[1975]));
    assign layer3_outputs[1100] = (layer2_outputs[2462]) & (layer2_outputs[1649]);
    assign layer3_outputs[1101] = ~(layer2_outputs[1202]) | (layer2_outputs[1525]);
    assign layer3_outputs[1102] = ~(layer2_outputs[403]);
    assign layer3_outputs[1103] = (layer2_outputs[447]) ^ (layer2_outputs[208]);
    assign layer3_outputs[1104] = ~((layer2_outputs[2307]) & (layer2_outputs[817]));
    assign layer3_outputs[1105] = ~((layer2_outputs[412]) | (layer2_outputs[232]));
    assign layer3_outputs[1106] = layer2_outputs[1143];
    assign layer3_outputs[1107] = (layer2_outputs[862]) & (layer2_outputs[1107]);
    assign layer3_outputs[1108] = layer2_outputs[2502];
    assign layer3_outputs[1109] = ~(layer2_outputs[947]);
    assign layer3_outputs[1110] = ~(layer2_outputs[505]);
    assign layer3_outputs[1111] = ~(layer2_outputs[1629]) | (layer2_outputs[962]);
    assign layer3_outputs[1112] = layer2_outputs[432];
    assign layer3_outputs[1113] = ~(layer2_outputs[86]) | (layer2_outputs[1820]);
    assign layer3_outputs[1114] = ~(layer2_outputs[327]) | (layer2_outputs[1731]);
    assign layer3_outputs[1115] = ~((layer2_outputs[309]) ^ (layer2_outputs[2009]));
    assign layer3_outputs[1116] = ~(layer2_outputs[366]) | (layer2_outputs[2235]);
    assign layer3_outputs[1117] = ~(layer2_outputs[1522]);
    assign layer3_outputs[1118] = 1'b1;
    assign layer3_outputs[1119] = ~(layer2_outputs[966]);
    assign layer3_outputs[1120] = ~(layer2_outputs[47]) | (layer2_outputs[2283]);
    assign layer3_outputs[1121] = ~((layer2_outputs[2416]) | (layer2_outputs[1768]));
    assign layer3_outputs[1122] = ~(layer2_outputs[2517]) | (layer2_outputs[1506]);
    assign layer3_outputs[1123] = ~((layer2_outputs[1500]) | (layer2_outputs[278]));
    assign layer3_outputs[1124] = (layer2_outputs[153]) & ~(layer2_outputs[1118]);
    assign layer3_outputs[1125] = ~(layer2_outputs[376]);
    assign layer3_outputs[1126] = (layer2_outputs[1273]) ^ (layer2_outputs[569]);
    assign layer3_outputs[1127] = (layer2_outputs[1390]) & (layer2_outputs[305]);
    assign layer3_outputs[1128] = ~(layer2_outputs[1264]) | (layer2_outputs[1254]);
    assign layer3_outputs[1129] = ~(layer2_outputs[141]) | (layer2_outputs[1932]);
    assign layer3_outputs[1130] = (layer2_outputs[526]) & ~(layer2_outputs[1828]);
    assign layer3_outputs[1131] = (layer2_outputs[2272]) & ~(layer2_outputs[1043]);
    assign layer3_outputs[1132] = layer2_outputs[291];
    assign layer3_outputs[1133] = ~(layer2_outputs[1265]);
    assign layer3_outputs[1134] = ~(layer2_outputs[2200]);
    assign layer3_outputs[1135] = (layer2_outputs[1046]) | (layer2_outputs[683]);
    assign layer3_outputs[1136] = ~((layer2_outputs[1039]) & (layer2_outputs[106]));
    assign layer3_outputs[1137] = ~((layer2_outputs[1570]) & (layer2_outputs[1968]));
    assign layer3_outputs[1138] = ~((layer2_outputs[187]) & (layer2_outputs[2036]));
    assign layer3_outputs[1139] = ~(layer2_outputs[346]);
    assign layer3_outputs[1140] = ~(layer2_outputs[2499]);
    assign layer3_outputs[1141] = ~(layer2_outputs[1559]);
    assign layer3_outputs[1142] = (layer2_outputs[1134]) & ~(layer2_outputs[972]);
    assign layer3_outputs[1143] = layer2_outputs[633];
    assign layer3_outputs[1144] = ~(layer2_outputs[1385]);
    assign layer3_outputs[1145] = (layer2_outputs[1304]) & ~(layer2_outputs[587]);
    assign layer3_outputs[1146] = layer2_outputs[1291];
    assign layer3_outputs[1147] = (layer2_outputs[1831]) & ~(layer2_outputs[1556]);
    assign layer3_outputs[1148] = (layer2_outputs[589]) & ~(layer2_outputs[1444]);
    assign layer3_outputs[1149] = 1'b1;
    assign layer3_outputs[1150] = (layer2_outputs[1808]) & (layer2_outputs[2113]);
    assign layer3_outputs[1151] = ~(layer2_outputs[581]) | (layer2_outputs[807]);
    assign layer3_outputs[1152] = ~((layer2_outputs[2132]) & (layer2_outputs[658]));
    assign layer3_outputs[1153] = layer2_outputs[345];
    assign layer3_outputs[1154] = ~(layer2_outputs[1832]) | (layer2_outputs[1316]);
    assign layer3_outputs[1155] = layer2_outputs[1170];
    assign layer3_outputs[1156] = ~((layer2_outputs[2498]) ^ (layer2_outputs[1692]));
    assign layer3_outputs[1157] = (layer2_outputs[1091]) ^ (layer2_outputs[1281]);
    assign layer3_outputs[1158] = (layer2_outputs[2151]) & ~(layer2_outputs[1533]);
    assign layer3_outputs[1159] = ~(layer2_outputs[524]);
    assign layer3_outputs[1160] = ~(layer2_outputs[431]);
    assign layer3_outputs[1161] = ~(layer2_outputs[1376]);
    assign layer3_outputs[1162] = ~((layer2_outputs[1390]) | (layer2_outputs[868]));
    assign layer3_outputs[1163] = (layer2_outputs[2375]) & ~(layer2_outputs[1607]);
    assign layer3_outputs[1164] = layer2_outputs[867];
    assign layer3_outputs[1165] = ~((layer2_outputs[1257]) & (layer2_outputs[801]));
    assign layer3_outputs[1166] = ~((layer2_outputs[121]) & (layer2_outputs[1117]));
    assign layer3_outputs[1167] = ~(layer2_outputs[1280]);
    assign layer3_outputs[1168] = ~(layer2_outputs[788]);
    assign layer3_outputs[1169] = ~((layer2_outputs[1155]) ^ (layer2_outputs[1749]));
    assign layer3_outputs[1170] = layer2_outputs[2194];
    assign layer3_outputs[1171] = layer2_outputs[968];
    assign layer3_outputs[1172] = ~((layer2_outputs[1211]) | (layer2_outputs[1890]));
    assign layer3_outputs[1173] = (layer2_outputs[582]) & ~(layer2_outputs[2166]);
    assign layer3_outputs[1174] = ~(layer2_outputs[1676]);
    assign layer3_outputs[1175] = layer2_outputs[1683];
    assign layer3_outputs[1176] = ~(layer2_outputs[873]) | (layer2_outputs[1902]);
    assign layer3_outputs[1177] = layer2_outputs[1606];
    assign layer3_outputs[1178] = (layer2_outputs[137]) & ~(layer2_outputs[805]);
    assign layer3_outputs[1179] = layer2_outputs[1307];
    assign layer3_outputs[1180] = (layer2_outputs[1863]) | (layer2_outputs[1929]);
    assign layer3_outputs[1181] = layer2_outputs[467];
    assign layer3_outputs[1182] = layer2_outputs[18];
    assign layer3_outputs[1183] = 1'b0;
    assign layer3_outputs[1184] = ~(layer2_outputs[1750]);
    assign layer3_outputs[1185] = ~((layer2_outputs[1454]) ^ (layer2_outputs[1537]));
    assign layer3_outputs[1186] = 1'b0;
    assign layer3_outputs[1187] = layer2_outputs[1420];
    assign layer3_outputs[1188] = (layer2_outputs[1426]) & ~(layer2_outputs[669]);
    assign layer3_outputs[1189] = 1'b0;
    assign layer3_outputs[1190] = ~(layer2_outputs[1319]);
    assign layer3_outputs[1191] = layer2_outputs[2440];
    assign layer3_outputs[1192] = ~(layer2_outputs[1188]);
    assign layer3_outputs[1193] = layer2_outputs[1461];
    assign layer3_outputs[1194] = ~(layer2_outputs[145]);
    assign layer3_outputs[1195] = (layer2_outputs[1693]) & (layer2_outputs[178]);
    assign layer3_outputs[1196] = (layer2_outputs[1972]) & ~(layer2_outputs[77]);
    assign layer3_outputs[1197] = ~(layer2_outputs[1332]) | (layer2_outputs[963]);
    assign layer3_outputs[1198] = 1'b1;
    assign layer3_outputs[1199] = ~(layer2_outputs[897]);
    assign layer3_outputs[1200] = ~(layer2_outputs[2114]);
    assign layer3_outputs[1201] = ~(layer2_outputs[2222]);
    assign layer3_outputs[1202] = layer2_outputs[2432];
    assign layer3_outputs[1203] = ~((layer2_outputs[1927]) & (layer2_outputs[364]));
    assign layer3_outputs[1204] = ~(layer2_outputs[332]) | (layer2_outputs[2480]);
    assign layer3_outputs[1205] = ~((layer2_outputs[1497]) | (layer2_outputs[292]));
    assign layer3_outputs[1206] = ~((layer2_outputs[2180]) & (layer2_outputs[1479]));
    assign layer3_outputs[1207] = ~(layer2_outputs[1200]);
    assign layer3_outputs[1208] = ~((layer2_outputs[1952]) & (layer2_outputs[321]));
    assign layer3_outputs[1209] = ~(layer2_outputs[1959]);
    assign layer3_outputs[1210] = layer2_outputs[1048];
    assign layer3_outputs[1211] = (layer2_outputs[1007]) & ~(layer2_outputs[2049]);
    assign layer3_outputs[1212] = layer2_outputs[655];
    assign layer3_outputs[1213] = ~((layer2_outputs[606]) | (layer2_outputs[2238]));
    assign layer3_outputs[1214] = (layer2_outputs[1406]) & ~(layer2_outputs[142]);
    assign layer3_outputs[1215] = (layer2_outputs[2434]) & ~(layer2_outputs[505]);
    assign layer3_outputs[1216] = (layer2_outputs[2090]) | (layer2_outputs[1700]);
    assign layer3_outputs[1217] = 1'b1;
    assign layer3_outputs[1218] = ~(layer2_outputs[1448]);
    assign layer3_outputs[1219] = 1'b0;
    assign layer3_outputs[1220] = ~(layer2_outputs[522]);
    assign layer3_outputs[1221] = (layer2_outputs[592]) | (layer2_outputs[541]);
    assign layer3_outputs[1222] = ~(layer2_outputs[2167]) | (layer2_outputs[1266]);
    assign layer3_outputs[1223] = ~(layer2_outputs[149]) | (layer2_outputs[2089]);
    assign layer3_outputs[1224] = (layer2_outputs[2424]) & (layer2_outputs[2507]);
    assign layer3_outputs[1225] = (layer2_outputs[1468]) & ~(layer2_outputs[700]);
    assign layer3_outputs[1226] = ~(layer2_outputs[536]);
    assign layer3_outputs[1227] = (layer2_outputs[2336]) & ~(layer2_outputs[1395]);
    assign layer3_outputs[1228] = (layer2_outputs[921]) ^ (layer2_outputs[1285]);
    assign layer3_outputs[1229] = ~(layer2_outputs[851]);
    assign layer3_outputs[1230] = ~(layer2_outputs[1177]);
    assign layer3_outputs[1231] = ~(layer2_outputs[1381]);
    assign layer3_outputs[1232] = ~(layer2_outputs[37]) | (layer2_outputs[1626]);
    assign layer3_outputs[1233] = ~(layer2_outputs[1914]);
    assign layer3_outputs[1234] = ~(layer2_outputs[1249]) | (layer2_outputs[1409]);
    assign layer3_outputs[1235] = layer2_outputs[298];
    assign layer3_outputs[1236] = ~(layer2_outputs[2002]);
    assign layer3_outputs[1237] = ~(layer2_outputs[997]);
    assign layer3_outputs[1238] = layer2_outputs[1263];
    assign layer3_outputs[1239] = layer2_outputs[1591];
    assign layer3_outputs[1240] = layer2_outputs[684];
    assign layer3_outputs[1241] = (layer2_outputs[491]) & ~(layer2_outputs[444]);
    assign layer3_outputs[1242] = layer2_outputs[464];
    assign layer3_outputs[1243] = (layer2_outputs[1842]) | (layer2_outputs[2043]);
    assign layer3_outputs[1244] = layer2_outputs[811];
    assign layer3_outputs[1245] = (layer2_outputs[107]) ^ (layer2_outputs[686]);
    assign layer3_outputs[1246] = ~(layer2_outputs[1653]);
    assign layer3_outputs[1247] = ~((layer2_outputs[2059]) | (layer2_outputs[1779]));
    assign layer3_outputs[1248] = layer2_outputs[1761];
    assign layer3_outputs[1249] = ~((layer2_outputs[434]) & (layer2_outputs[1104]));
    assign layer3_outputs[1250] = ~((layer2_outputs[1571]) ^ (layer2_outputs[1141]));
    assign layer3_outputs[1251] = layer2_outputs[623];
    assign layer3_outputs[1252] = ~((layer2_outputs[434]) | (layer2_outputs[1905]));
    assign layer3_outputs[1253] = ~(layer2_outputs[2110]);
    assign layer3_outputs[1254] = (layer2_outputs[1456]) & ~(layer2_outputs[2088]);
    assign layer3_outputs[1255] = layer2_outputs[1695];
    assign layer3_outputs[1256] = ~(layer2_outputs[2124]);
    assign layer3_outputs[1257] = ~(layer2_outputs[1604]) | (layer2_outputs[386]);
    assign layer3_outputs[1258] = ~(layer2_outputs[2235]);
    assign layer3_outputs[1259] = (layer2_outputs[2441]) & ~(layer2_outputs[2317]);
    assign layer3_outputs[1260] = (layer2_outputs[297]) & ~(layer2_outputs[1377]);
    assign layer3_outputs[1261] = 1'b1;
    assign layer3_outputs[1262] = layer2_outputs[1582];
    assign layer3_outputs[1263] = (layer2_outputs[1722]) | (layer2_outputs[1462]);
    assign layer3_outputs[1264] = ~(layer2_outputs[1021]) | (layer2_outputs[176]);
    assign layer3_outputs[1265] = ~(layer2_outputs[1455]);
    assign layer3_outputs[1266] = ~(layer2_outputs[196]);
    assign layer3_outputs[1267] = (layer2_outputs[1974]) & (layer2_outputs[1378]);
    assign layer3_outputs[1268] = 1'b1;
    assign layer3_outputs[1269] = 1'b0;
    assign layer3_outputs[1270] = 1'b1;
    assign layer3_outputs[1271] = ~((layer2_outputs[491]) & (layer2_outputs[1476]));
    assign layer3_outputs[1272] = ~(layer2_outputs[634]);
    assign layer3_outputs[1273] = ~((layer2_outputs[737]) ^ (layer2_outputs[1714]));
    assign layer3_outputs[1274] = layer2_outputs[1017];
    assign layer3_outputs[1275] = (layer2_outputs[2401]) & ~(layer2_outputs[1426]);
    assign layer3_outputs[1276] = ~(layer2_outputs[322]);
    assign layer3_outputs[1277] = ~(layer2_outputs[761]) | (layer2_outputs[1607]);
    assign layer3_outputs[1278] = (layer2_outputs[2453]) | (layer2_outputs[1702]);
    assign layer3_outputs[1279] = ~(layer2_outputs[1391]) | (layer2_outputs[2468]);
    assign layer3_outputs[1280] = (layer2_outputs[437]) & ~(layer2_outputs[2429]);
    assign layer3_outputs[1281] = layer2_outputs[917];
    assign layer3_outputs[1282] = (layer2_outputs[1049]) | (layer2_outputs[1109]);
    assign layer3_outputs[1283] = layer2_outputs[353];
    assign layer3_outputs[1284] = layer2_outputs[2447];
    assign layer3_outputs[1285] = ~((layer2_outputs[700]) ^ (layer2_outputs[670]));
    assign layer3_outputs[1286] = ~(layer2_outputs[272]);
    assign layer3_outputs[1287] = (layer2_outputs[710]) & (layer2_outputs[2357]);
    assign layer3_outputs[1288] = (layer2_outputs[2524]) | (layer2_outputs[1224]);
    assign layer3_outputs[1289] = ~(layer2_outputs[587]) | (layer2_outputs[1806]);
    assign layer3_outputs[1290] = ~(layer2_outputs[210]);
    assign layer3_outputs[1291] = ~(layer2_outputs[62]) | (layer2_outputs[2106]);
    assign layer3_outputs[1292] = ~(layer2_outputs[68]);
    assign layer3_outputs[1293] = layer2_outputs[1316];
    assign layer3_outputs[1294] = ~(layer2_outputs[96]) | (layer2_outputs[1608]);
    assign layer3_outputs[1295] = (layer2_outputs[269]) & ~(layer2_outputs[2392]);
    assign layer3_outputs[1296] = ~(layer2_outputs[1216]);
    assign layer3_outputs[1297] = ~(layer2_outputs[2512]);
    assign layer3_outputs[1298] = ~((layer2_outputs[2115]) | (layer2_outputs[2159]));
    assign layer3_outputs[1299] = ~((layer2_outputs[2320]) & (layer2_outputs[282]));
    assign layer3_outputs[1300] = layer2_outputs[939];
    assign layer3_outputs[1301] = ~(layer2_outputs[1196]);
    assign layer3_outputs[1302] = ~((layer2_outputs[2449]) & (layer2_outputs[1642]));
    assign layer3_outputs[1303] = ~((layer2_outputs[2233]) | (layer2_outputs[2421]));
    assign layer3_outputs[1304] = (layer2_outputs[499]) ^ (layer2_outputs[612]);
    assign layer3_outputs[1305] = layer2_outputs[960];
    assign layer3_outputs[1306] = (layer2_outputs[816]) & (layer2_outputs[2499]);
    assign layer3_outputs[1307] = ~(layer2_outputs[2265]) | (layer2_outputs[1305]);
    assign layer3_outputs[1308] = (layer2_outputs[1224]) & (layer2_outputs[1248]);
    assign layer3_outputs[1309] = (layer2_outputs[1303]) | (layer2_outputs[964]);
    assign layer3_outputs[1310] = ~(layer2_outputs[2308]);
    assign layer3_outputs[1311] = 1'b1;
    assign layer3_outputs[1312] = (layer2_outputs[1929]) & (layer2_outputs[168]);
    assign layer3_outputs[1313] = ~(layer2_outputs[2135]);
    assign layer3_outputs[1314] = (layer2_outputs[1802]) & (layer2_outputs[1997]);
    assign layer3_outputs[1315] = layer2_outputs[1491];
    assign layer3_outputs[1316] = (layer2_outputs[1052]) & (layer2_outputs[2331]);
    assign layer3_outputs[1317] = (layer2_outputs[1857]) & ~(layer2_outputs[543]);
    assign layer3_outputs[1318] = (layer2_outputs[2245]) & (layer2_outputs[1503]);
    assign layer3_outputs[1319] = ~(layer2_outputs[170]);
    assign layer3_outputs[1320] = (layer2_outputs[2507]) ^ (layer2_outputs[1724]);
    assign layer3_outputs[1321] = ~(layer2_outputs[1958]);
    assign layer3_outputs[1322] = ~((layer2_outputs[465]) & (layer2_outputs[1142]));
    assign layer3_outputs[1323] = (layer2_outputs[1715]) & ~(layer2_outputs[1833]);
    assign layer3_outputs[1324] = (layer2_outputs[2133]) | (layer2_outputs[603]);
    assign layer3_outputs[1325] = ~(layer2_outputs[368]) | (layer2_outputs[1268]);
    assign layer3_outputs[1326] = ~((layer2_outputs[157]) & (layer2_outputs[2198]));
    assign layer3_outputs[1327] = layer2_outputs[1030];
    assign layer3_outputs[1328] = ~(layer2_outputs[856]);
    assign layer3_outputs[1329] = ~(layer2_outputs[2375]) | (layer2_outputs[669]);
    assign layer3_outputs[1330] = ~(layer2_outputs[390]);
    assign layer3_outputs[1331] = 1'b0;
    assign layer3_outputs[1332] = ~(layer2_outputs[1340]);
    assign layer3_outputs[1333] = ~(layer2_outputs[1450]) | (layer2_outputs[1541]);
    assign layer3_outputs[1334] = layer2_outputs[1687];
    assign layer3_outputs[1335] = layer2_outputs[2383];
    assign layer3_outputs[1336] = (layer2_outputs[179]) | (layer2_outputs[2215]);
    assign layer3_outputs[1337] = ~(layer2_outputs[760]);
    assign layer3_outputs[1338] = layer2_outputs[985];
    assign layer3_outputs[1339] = layer2_outputs[2034];
    assign layer3_outputs[1340] = (layer2_outputs[936]) | (layer2_outputs[1286]);
    assign layer3_outputs[1341] = ~(layer2_outputs[524]);
    assign layer3_outputs[1342] = (layer2_outputs[1871]) ^ (layer2_outputs[2186]);
    assign layer3_outputs[1343] = layer2_outputs[2393];
    assign layer3_outputs[1344] = layer2_outputs[461];
    assign layer3_outputs[1345] = layer2_outputs[1015];
    assign layer3_outputs[1346] = ~((layer2_outputs[1373]) & (layer2_outputs[311]));
    assign layer3_outputs[1347] = (layer2_outputs[1530]) & ~(layer2_outputs[2381]);
    assign layer3_outputs[1348] = ~((layer2_outputs[601]) & (layer2_outputs[920]));
    assign layer3_outputs[1349] = ~(layer2_outputs[1736]) | (layer2_outputs[1675]);
    assign layer3_outputs[1350] = layer2_outputs[1521];
    assign layer3_outputs[1351] = (layer2_outputs[1524]) & (layer2_outputs[1578]);
    assign layer3_outputs[1352] = ~(layer2_outputs[1716]) | (layer2_outputs[257]);
    assign layer3_outputs[1353] = ~(layer2_outputs[1755]);
    assign layer3_outputs[1354] = layer2_outputs[1548];
    assign layer3_outputs[1355] = ~((layer2_outputs[2317]) ^ (layer2_outputs[370]));
    assign layer3_outputs[1356] = (layer2_outputs[1612]) | (layer2_outputs[2260]);
    assign layer3_outputs[1357] = 1'b1;
    assign layer3_outputs[1358] = layer2_outputs[1908];
    assign layer3_outputs[1359] = ~(layer2_outputs[1713]);
    assign layer3_outputs[1360] = ~((layer2_outputs[1797]) ^ (layer2_outputs[1931]));
    assign layer3_outputs[1361] = ~(layer2_outputs[958]) | (layer2_outputs[693]);
    assign layer3_outputs[1362] = 1'b0;
    assign layer3_outputs[1363] = (layer2_outputs[2491]) | (layer2_outputs[490]);
    assign layer3_outputs[1364] = (layer2_outputs[2509]) & ~(layer2_outputs[1418]);
    assign layer3_outputs[1365] = ~(layer2_outputs[1945]);
    assign layer3_outputs[1366] = layer2_outputs[2111];
    assign layer3_outputs[1367] = layer2_outputs[1076];
    assign layer3_outputs[1368] = layer2_outputs[140];
    assign layer3_outputs[1369] = layer2_outputs[1556];
    assign layer3_outputs[1370] = (layer2_outputs[1422]) & ~(layer2_outputs[2260]);
    assign layer3_outputs[1371] = ~(layer2_outputs[1470]);
    assign layer3_outputs[1372] = (layer2_outputs[2059]) ^ (layer2_outputs[676]);
    assign layer3_outputs[1373] = ~((layer2_outputs[520]) & (layer2_outputs[2377]));
    assign layer3_outputs[1374] = 1'b1;
    assign layer3_outputs[1375] = ~(layer2_outputs[449]) | (layer2_outputs[1976]);
    assign layer3_outputs[1376] = (layer2_outputs[2226]) & ~(layer2_outputs[188]);
    assign layer3_outputs[1377] = layer2_outputs[1700];
    assign layer3_outputs[1378] = (layer2_outputs[1088]) | (layer2_outputs[1001]);
    assign layer3_outputs[1379] = ~(layer2_outputs[1267]);
    assign layer3_outputs[1380] = ~(layer2_outputs[162]) | (layer2_outputs[1614]);
    assign layer3_outputs[1381] = 1'b0;
    assign layer3_outputs[1382] = ~(layer2_outputs[34]);
    assign layer3_outputs[1383] = ~((layer2_outputs[1636]) | (layer2_outputs[1095]));
    assign layer3_outputs[1384] = layer2_outputs[1752];
    assign layer3_outputs[1385] = (layer2_outputs[1600]) & ~(layer2_outputs[442]);
    assign layer3_outputs[1386] = (layer2_outputs[628]) & (layer2_outputs[1071]);
    assign layer3_outputs[1387] = (layer2_outputs[1416]) ^ (layer2_outputs[66]);
    assign layer3_outputs[1388] = (layer2_outputs[759]) & ~(layer2_outputs[1415]);
    assign layer3_outputs[1389] = (layer2_outputs[775]) & ~(layer2_outputs[338]);
    assign layer3_outputs[1390] = 1'b1;
    assign layer3_outputs[1391] = 1'b0;
    assign layer3_outputs[1392] = ~(layer2_outputs[729]) | (layer2_outputs[1673]);
    assign layer3_outputs[1393] = (layer2_outputs[1081]) | (layer2_outputs[1179]);
    assign layer3_outputs[1394] = 1'b0;
    assign layer3_outputs[1395] = ~(layer2_outputs[1099]);
    assign layer3_outputs[1396] = ~(layer2_outputs[135]) | (layer2_outputs[2193]);
    assign layer3_outputs[1397] = layer2_outputs[336];
    assign layer3_outputs[1398] = ~((layer2_outputs[254]) | (layer2_outputs[2035]));
    assign layer3_outputs[1399] = (layer2_outputs[349]) & (layer2_outputs[806]);
    assign layer3_outputs[1400] = layer2_outputs[2459];
    assign layer3_outputs[1401] = ~(layer2_outputs[143]);
    assign layer3_outputs[1402] = ~((layer2_outputs[810]) ^ (layer2_outputs[86]));
    assign layer3_outputs[1403] = (layer2_outputs[2019]) & ~(layer2_outputs[5]);
    assign layer3_outputs[1404] = ~(layer2_outputs[1918]) | (layer2_outputs[880]);
    assign layer3_outputs[1405] = ~((layer2_outputs[1976]) | (layer2_outputs[2335]));
    assign layer3_outputs[1406] = (layer2_outputs[2134]) & ~(layer2_outputs[1038]);
    assign layer3_outputs[1407] = ~(layer2_outputs[2215]);
    assign layer3_outputs[1408] = layer2_outputs[2095];
    assign layer3_outputs[1409] = ~((layer2_outputs[2552]) ^ (layer2_outputs[1112]));
    assign layer3_outputs[1410] = ~((layer2_outputs[308]) ^ (layer2_outputs[159]));
    assign layer3_outputs[1411] = layer2_outputs[780];
    assign layer3_outputs[1412] = (layer2_outputs[1714]) & ~(layer2_outputs[1171]);
    assign layer3_outputs[1413] = ~(layer2_outputs[1459]) | (layer2_outputs[2244]);
    assign layer3_outputs[1414] = ~((layer2_outputs[942]) | (layer2_outputs[2327]));
    assign layer3_outputs[1415] = ~(layer2_outputs[22]);
    assign layer3_outputs[1416] = layer2_outputs[1735];
    assign layer3_outputs[1417] = ~((layer2_outputs[1977]) ^ (layer2_outputs[2]));
    assign layer3_outputs[1418] = ~((layer2_outputs[1401]) & (layer2_outputs[154]));
    assign layer3_outputs[1419] = ~(layer2_outputs[632]) | (layer2_outputs[201]);
    assign layer3_outputs[1420] = (layer2_outputs[1194]) & ~(layer2_outputs[2197]);
    assign layer3_outputs[1421] = layer2_outputs[612];
    assign layer3_outputs[1422] = layer2_outputs[919];
    assign layer3_outputs[1423] = (layer2_outputs[2075]) ^ (layer2_outputs[2313]);
    assign layer3_outputs[1424] = ~(layer2_outputs[1825]);
    assign layer3_outputs[1425] = layer2_outputs[2400];
    assign layer3_outputs[1426] = ~(layer2_outputs[941]) | (layer2_outputs[1340]);
    assign layer3_outputs[1427] = ~(layer2_outputs[1183]);
    assign layer3_outputs[1428] = (layer2_outputs[1597]) | (layer2_outputs[888]);
    assign layer3_outputs[1429] = ~(layer2_outputs[1097]);
    assign layer3_outputs[1430] = ~(layer2_outputs[2094]);
    assign layer3_outputs[1431] = (layer2_outputs[112]) & ~(layer2_outputs[1696]);
    assign layer3_outputs[1432] = layer2_outputs[1987];
    assign layer3_outputs[1433] = (layer2_outputs[1608]) & (layer2_outputs[1655]);
    assign layer3_outputs[1434] = layer2_outputs[2050];
    assign layer3_outputs[1435] = ~(layer2_outputs[1600]);
    assign layer3_outputs[1436] = 1'b1;
    assign layer3_outputs[1437] = ~(layer2_outputs[1754]) | (layer2_outputs[2029]);
    assign layer3_outputs[1438] = ~(layer2_outputs[1591]) | (layer2_outputs[306]);
    assign layer3_outputs[1439] = ~(layer2_outputs[2502]) | (layer2_outputs[1206]);
    assign layer3_outputs[1440] = ~((layer2_outputs[764]) & (layer2_outputs[1021]));
    assign layer3_outputs[1441] = ~(layer2_outputs[476]);
    assign layer3_outputs[1442] = ~(layer2_outputs[947]);
    assign layer3_outputs[1443] = ~((layer2_outputs[1481]) | (layer2_outputs[713]));
    assign layer3_outputs[1444] = ~(layer2_outputs[1533]) | (layer2_outputs[2199]);
    assign layer3_outputs[1445] = 1'b1;
    assign layer3_outputs[1446] = ~((layer2_outputs[2223]) ^ (layer2_outputs[714]));
    assign layer3_outputs[1447] = (layer2_outputs[1449]) ^ (layer2_outputs[1486]);
    assign layer3_outputs[1448] = 1'b0;
    assign layer3_outputs[1449] = layer2_outputs[2089];
    assign layer3_outputs[1450] = ~((layer2_outputs[71]) | (layer2_outputs[568]));
    assign layer3_outputs[1451] = 1'b1;
    assign layer3_outputs[1452] = (layer2_outputs[294]) & (layer2_outputs[675]);
    assign layer3_outputs[1453] = layer2_outputs[2058];
    assign layer3_outputs[1454] = (layer2_outputs[10]) & ~(layer2_outputs[2027]);
    assign layer3_outputs[1455] = ~(layer2_outputs[359]);
    assign layer3_outputs[1456] = ~((layer2_outputs[1159]) & (layer2_outputs[2294]));
    assign layer3_outputs[1457] = (layer2_outputs[1474]) & ~(layer2_outputs[1659]);
    assign layer3_outputs[1458] = ~(layer2_outputs[304]);
    assign layer3_outputs[1459] = (layer2_outputs[654]) ^ (layer2_outputs[1535]);
    assign layer3_outputs[1460] = (layer2_outputs[1185]) & (layer2_outputs[361]);
    assign layer3_outputs[1461] = layer2_outputs[2395];
    assign layer3_outputs[1462] = (layer2_outputs[126]) & ~(layer2_outputs[624]);
    assign layer3_outputs[1463] = layer2_outputs[1290];
    assign layer3_outputs[1464] = ~(layer2_outputs[2130]);
    assign layer3_outputs[1465] = layer2_outputs[578];
    assign layer3_outputs[1466] = layer2_outputs[385];
    assign layer3_outputs[1467] = ~(layer2_outputs[523]);
    assign layer3_outputs[1468] = ~(layer2_outputs[109]);
    assign layer3_outputs[1469] = ~((layer2_outputs[1992]) & (layer2_outputs[919]));
    assign layer3_outputs[1470] = ~(layer2_outputs[2296]);
    assign layer3_outputs[1471] = (layer2_outputs[1697]) & (layer2_outputs[1559]);
    assign layer3_outputs[1472] = 1'b1;
    assign layer3_outputs[1473] = layer2_outputs[1951];
    assign layer3_outputs[1474] = ~(layer2_outputs[473]);
    assign layer3_outputs[1475] = layer2_outputs[1750];
    assign layer3_outputs[1476] = ~(layer2_outputs[1584]);
    assign layer3_outputs[1477] = ~(layer2_outputs[236]);
    assign layer3_outputs[1478] = (layer2_outputs[1641]) & ~(layer2_outputs[347]);
    assign layer3_outputs[1479] = (layer2_outputs[1668]) ^ (layer2_outputs[1731]);
    assign layer3_outputs[1480] = ~(layer2_outputs[1246]);
    assign layer3_outputs[1481] = layer2_outputs[2447];
    assign layer3_outputs[1482] = 1'b0;
    assign layer3_outputs[1483] = (layer2_outputs[1130]) & (layer2_outputs[617]);
    assign layer3_outputs[1484] = (layer2_outputs[2227]) & ~(layer2_outputs[252]);
    assign layer3_outputs[1485] = ~(layer2_outputs[26]);
    assign layer3_outputs[1486] = layer2_outputs[696];
    assign layer3_outputs[1487] = (layer2_outputs[1944]) & ~(layer2_outputs[959]);
    assign layer3_outputs[1488] = ~((layer2_outputs[1577]) & (layer2_outputs[2368]));
    assign layer3_outputs[1489] = ~(layer2_outputs[1086]) | (layer2_outputs[243]);
    assign layer3_outputs[1490] = (layer2_outputs[2021]) | (layer2_outputs[264]);
    assign layer3_outputs[1491] = layer2_outputs[1164];
    assign layer3_outputs[1492] = ~((layer2_outputs[508]) ^ (layer2_outputs[2443]));
    assign layer3_outputs[1493] = ~(layer2_outputs[398]) | (layer2_outputs[1875]);
    assign layer3_outputs[1494] = (layer2_outputs[238]) ^ (layer2_outputs[1331]);
    assign layer3_outputs[1495] = layer2_outputs[1469];
    assign layer3_outputs[1496] = ~(layer2_outputs[114]);
    assign layer3_outputs[1497] = ~(layer2_outputs[757]);
    assign layer3_outputs[1498] = ~(layer2_outputs[1404]) | (layer2_outputs[1271]);
    assign layer3_outputs[1499] = 1'b1;
    assign layer3_outputs[1500] = ~(layer2_outputs[533]) | (layer2_outputs[2270]);
    assign layer3_outputs[1501] = ~(layer2_outputs[2141]) | (layer2_outputs[772]);
    assign layer3_outputs[1502] = layer2_outputs[739];
    assign layer3_outputs[1503] = layer2_outputs[1663];
    assign layer3_outputs[1504] = (layer2_outputs[2062]) & (layer2_outputs[207]);
    assign layer3_outputs[1505] = ~(layer2_outputs[2107]);
    assign layer3_outputs[1506] = ~(layer2_outputs[1907]) | (layer2_outputs[833]);
    assign layer3_outputs[1507] = ~(layer2_outputs[255]);
    assign layer3_outputs[1508] = ~((layer2_outputs[1174]) & (layer2_outputs[173]));
    assign layer3_outputs[1509] = ~(layer2_outputs[1108]);
    assign layer3_outputs[1510] = layer2_outputs[532];
    assign layer3_outputs[1511] = (layer2_outputs[1894]) & (layer2_outputs[2219]);
    assign layer3_outputs[1512] = 1'b1;
    assign layer3_outputs[1513] = (layer2_outputs[1040]) & ~(layer2_outputs[1072]);
    assign layer3_outputs[1514] = layer2_outputs[735];
    assign layer3_outputs[1515] = ~((layer2_outputs[72]) | (layer2_outputs[1883]));
    assign layer3_outputs[1516] = ~(layer2_outputs[116]);
    assign layer3_outputs[1517] = layer2_outputs[59];
    assign layer3_outputs[1518] = ~(layer2_outputs[1427]);
    assign layer3_outputs[1519] = ~(layer2_outputs[1810]) | (layer2_outputs[1482]);
    assign layer3_outputs[1520] = ~(layer2_outputs[1163]) | (layer2_outputs[1233]);
    assign layer3_outputs[1521] = layer2_outputs[1822];
    assign layer3_outputs[1522] = ~(layer2_outputs[547]) | (layer2_outputs[770]);
    assign layer3_outputs[1523] = (layer2_outputs[2263]) & (layer2_outputs[2119]);
    assign layer3_outputs[1524] = layer2_outputs[2174];
    assign layer3_outputs[1525] = layer2_outputs[655];
    assign layer3_outputs[1526] = ~(layer2_outputs[894]) | (layer2_outputs[2109]);
    assign layer3_outputs[1527] = layer2_outputs[1129];
    assign layer3_outputs[1528] = ~(layer2_outputs[2242]);
    assign layer3_outputs[1529] = (layer2_outputs[2258]) ^ (layer2_outputs[245]);
    assign layer3_outputs[1530] = (layer2_outputs[288]) & (layer2_outputs[1066]);
    assign layer3_outputs[1531] = layer2_outputs[583];
    assign layer3_outputs[1532] = ~((layer2_outputs[1939]) ^ (layer2_outputs[1860]));
    assign layer3_outputs[1533] = layer2_outputs[85];
    assign layer3_outputs[1534] = ~(layer2_outputs[1484]);
    assign layer3_outputs[1535] = layer2_outputs[49];
    assign layer3_outputs[1536] = layer2_outputs[868];
    assign layer3_outputs[1537] = layer2_outputs[800];
    assign layer3_outputs[1538] = ~(layer2_outputs[1298]) | (layer2_outputs[1351]);
    assign layer3_outputs[1539] = (layer2_outputs[2385]) & ~(layer2_outputs[1252]);
    assign layer3_outputs[1540] = (layer2_outputs[746]) | (layer2_outputs[948]);
    assign layer3_outputs[1541] = ~(layer2_outputs[1739]) | (layer2_outputs[1476]);
    assign layer3_outputs[1542] = ~(layer2_outputs[80]);
    assign layer3_outputs[1543] = (layer2_outputs[297]) & ~(layer2_outputs[1038]);
    assign layer3_outputs[1544] = (layer2_outputs[1251]) & ~(layer2_outputs[2319]);
    assign layer3_outputs[1545] = ~(layer2_outputs[1989]) | (layer2_outputs[1147]);
    assign layer3_outputs[1546] = ~(layer2_outputs[1431]) | (layer2_outputs[2047]);
    assign layer3_outputs[1547] = layer2_outputs[550];
    assign layer3_outputs[1548] = ~(layer2_outputs[87]) | (layer2_outputs[264]);
    assign layer3_outputs[1549] = layer2_outputs[216];
    assign layer3_outputs[1550] = (layer2_outputs[1396]) & ~(layer2_outputs[2268]);
    assign layer3_outputs[1551] = ~(layer2_outputs[1819]);
    assign layer3_outputs[1552] = (layer2_outputs[120]) | (layer2_outputs[89]);
    assign layer3_outputs[1553] = layer2_outputs[1470];
    assign layer3_outputs[1554] = ~((layer2_outputs[982]) ^ (layer2_outputs[1288]));
    assign layer3_outputs[1555] = ~((layer2_outputs[1904]) | (layer2_outputs[1019]));
    assign layer3_outputs[1556] = ~(layer2_outputs[306]);
    assign layer3_outputs[1557] = layer2_outputs[2203];
    assign layer3_outputs[1558] = layer2_outputs[566];
    assign layer3_outputs[1559] = ~((layer2_outputs[1455]) ^ (layer2_outputs[61]));
    assign layer3_outputs[1560] = ~(layer2_outputs[1555]) | (layer2_outputs[1719]);
    assign layer3_outputs[1561] = 1'b1;
    assign layer3_outputs[1562] = layer2_outputs[1889];
    assign layer3_outputs[1563] = ~(layer2_outputs[10]);
    assign layer3_outputs[1564] = (layer2_outputs[514]) & ~(layer2_outputs[590]);
    assign layer3_outputs[1565] = layer2_outputs[278];
    assign layer3_outputs[1566] = layer2_outputs[635];
    assign layer3_outputs[1567] = layer2_outputs[1621];
    assign layer3_outputs[1568] = (layer2_outputs[2154]) & ~(layer2_outputs[766]);
    assign layer3_outputs[1569] = (layer2_outputs[645]) & (layer2_outputs[453]);
    assign layer3_outputs[1570] = ~(layer2_outputs[1637]);
    assign layer3_outputs[1571] = ~(layer2_outputs[1498]) | (layer2_outputs[2544]);
    assign layer3_outputs[1572] = ~((layer2_outputs[1544]) & (layer2_outputs[788]));
    assign layer3_outputs[1573] = layer2_outputs[1883];
    assign layer3_outputs[1574] = layer2_outputs[995];
    assign layer3_outputs[1575] = ~(layer2_outputs[2263]);
    assign layer3_outputs[1576] = ~((layer2_outputs[2497]) | (layer2_outputs[242]));
    assign layer3_outputs[1577] = layer2_outputs[782];
    assign layer3_outputs[1578] = (layer2_outputs[2363]) & ~(layer2_outputs[2384]);
    assign layer3_outputs[1579] = 1'b1;
    assign layer3_outputs[1580] = (layer2_outputs[1369]) | (layer2_outputs[773]);
    assign layer3_outputs[1581] = layer2_outputs[1027];
    assign layer3_outputs[1582] = layer2_outputs[660];
    assign layer3_outputs[1583] = ~((layer2_outputs[2018]) & (layer2_outputs[2353]));
    assign layer3_outputs[1584] = ~((layer2_outputs[65]) | (layer2_outputs[276]));
    assign layer3_outputs[1585] = layer2_outputs[1562];
    assign layer3_outputs[1586] = (layer2_outputs[2038]) & ~(layer2_outputs[944]);
    assign layer3_outputs[1587] = (layer2_outputs[1414]) & ~(layer2_outputs[374]);
    assign layer3_outputs[1588] = (layer2_outputs[713]) | (layer2_outputs[495]);
    assign layer3_outputs[1589] = ~((layer2_outputs[2475]) | (layer2_outputs[1020]));
    assign layer3_outputs[1590] = 1'b0;
    assign layer3_outputs[1591] = ~(layer2_outputs[2363]);
    assign layer3_outputs[1592] = 1'b1;
    assign layer3_outputs[1593] = ~(layer2_outputs[1320]);
    assign layer3_outputs[1594] = ~(layer2_outputs[331]);
    assign layer3_outputs[1595] = (layer2_outputs[2514]) & ~(layer2_outputs[1631]);
    assign layer3_outputs[1596] = layer2_outputs[2171];
    assign layer3_outputs[1597] = layer2_outputs[2293];
    assign layer3_outputs[1598] = ~(layer2_outputs[1540]);
    assign layer3_outputs[1599] = layer2_outputs[1895];
    assign layer3_outputs[1600] = layer2_outputs[986];
    assign layer3_outputs[1601] = ~((layer2_outputs[1209]) | (layer2_outputs[808]));
    assign layer3_outputs[1602] = (layer2_outputs[1644]) | (layer2_outputs[52]);
    assign layer3_outputs[1603] = 1'b0;
    assign layer3_outputs[1604] = layer2_outputs[1699];
    assign layer3_outputs[1605] = ~(layer2_outputs[1498]);
    assign layer3_outputs[1606] = layer2_outputs[1382];
    assign layer3_outputs[1607] = ~(layer2_outputs[1500]);
    assign layer3_outputs[1608] = ~(layer2_outputs[995]);
    assign layer3_outputs[1609] = ~(layer2_outputs[2208]);
    assign layer3_outputs[1610] = (layer2_outputs[1443]) | (layer2_outputs[1574]);
    assign layer3_outputs[1611] = ~(layer2_outputs[2528]);
    assign layer3_outputs[1612] = ~(layer2_outputs[456]) | (layer2_outputs[1327]);
    assign layer3_outputs[1613] = layer2_outputs[4];
    assign layer3_outputs[1614] = (layer2_outputs[2557]) ^ (layer2_outputs[137]);
    assign layer3_outputs[1615] = (layer2_outputs[658]) & (layer2_outputs[1939]);
    assign layer3_outputs[1616] = (layer2_outputs[1475]) ^ (layer2_outputs[989]);
    assign layer3_outputs[1617] = ~(layer2_outputs[1033]);
    assign layer3_outputs[1618] = ~((layer2_outputs[2543]) | (layer2_outputs[732]));
    assign layer3_outputs[1619] = ~(layer2_outputs[2264]);
    assign layer3_outputs[1620] = ~(layer2_outputs[1155]) | (layer2_outputs[1248]);
    assign layer3_outputs[1621] = ~(layer2_outputs[2193]) | (layer2_outputs[631]);
    assign layer3_outputs[1622] = ~(layer2_outputs[1358]);
    assign layer3_outputs[1623] = (layer2_outputs[472]) & ~(layer2_outputs[1302]);
    assign layer3_outputs[1624] = ~(layer2_outputs[656]) | (layer2_outputs[478]);
    assign layer3_outputs[1625] = 1'b0;
    assign layer3_outputs[1626] = ~(layer2_outputs[1265]);
    assign layer3_outputs[1627] = ~(layer2_outputs[1756]);
    assign layer3_outputs[1628] = layer2_outputs[2389];
    assign layer3_outputs[1629] = ~(layer2_outputs[1253]);
    assign layer3_outputs[1630] = layer2_outputs[1298];
    assign layer3_outputs[1631] = ~(layer2_outputs[502]);
    assign layer3_outputs[1632] = layer2_outputs[1829];
    assign layer3_outputs[1633] = layer2_outputs[215];
    assign layer3_outputs[1634] = layer2_outputs[707];
    assign layer3_outputs[1635] = ~((layer2_outputs[320]) | (layer2_outputs[1450]));
    assign layer3_outputs[1636] = 1'b1;
    assign layer3_outputs[1637] = layer2_outputs[1452];
    assign layer3_outputs[1638] = layer2_outputs[2144];
    assign layer3_outputs[1639] = (layer2_outputs[45]) & ~(layer2_outputs[1320]);
    assign layer3_outputs[1640] = 1'b1;
    assign layer3_outputs[1641] = ~((layer2_outputs[1282]) ^ (layer2_outputs[1969]));
    assign layer3_outputs[1642] = (layer2_outputs[973]) & ~(layer2_outputs[1584]);
    assign layer3_outputs[1643] = ~(layer2_outputs[629]);
    assign layer3_outputs[1644] = (layer2_outputs[1192]) | (layer2_outputs[1422]);
    assign layer3_outputs[1645] = ~(layer2_outputs[2126]);
    assign layer3_outputs[1646] = ~(layer2_outputs[1730]);
    assign layer3_outputs[1647] = ~((layer2_outputs[2373]) | (layer2_outputs[2176]));
    assign layer3_outputs[1648] = (layer2_outputs[2288]) & ~(layer2_outputs[575]);
    assign layer3_outputs[1649] = ~(layer2_outputs[565]);
    assign layer3_outputs[1650] = 1'b0;
    assign layer3_outputs[1651] = ~((layer2_outputs[1669]) ^ (layer2_outputs[671]));
    assign layer3_outputs[1652] = (layer2_outputs[2400]) & (layer2_outputs[483]);
    assign layer3_outputs[1653] = ~((layer2_outputs[663]) ^ (layer2_outputs[1839]));
    assign layer3_outputs[1654] = (layer2_outputs[2086]) & (layer2_outputs[828]);
    assign layer3_outputs[1655] = ~(layer2_outputs[386]);
    assign layer3_outputs[1656] = (layer2_outputs[1656]) ^ (layer2_outputs[1874]);
    assign layer3_outputs[1657] = ~(layer2_outputs[2522]);
    assign layer3_outputs[1658] = ~((layer2_outputs[2552]) & (layer2_outputs[1541]));
    assign layer3_outputs[1659] = layer2_outputs[895];
    assign layer3_outputs[1660] = ~(layer2_outputs[1836]);
    assign layer3_outputs[1661] = 1'b1;
    assign layer3_outputs[1662] = ~(layer2_outputs[2007]);
    assign layer3_outputs[1663] = ~((layer2_outputs[547]) & (layer2_outputs[784]));
    assign layer3_outputs[1664] = 1'b1;
    assign layer3_outputs[1665] = ~(layer2_outputs[1879]);
    assign layer3_outputs[1666] = ~(layer2_outputs[1567]) | (layer2_outputs[2252]);
    assign layer3_outputs[1667] = ~(layer2_outputs[1011]);
    assign layer3_outputs[1668] = layer2_outputs[1090];
    assign layer3_outputs[1669] = (layer2_outputs[636]) & (layer2_outputs[2554]);
    assign layer3_outputs[1670] = ~((layer2_outputs[1034]) | (layer2_outputs[1734]));
    assign layer3_outputs[1671] = layer2_outputs[917];
    assign layer3_outputs[1672] = layer2_outputs[1984];
    assign layer3_outputs[1673] = ~(layer2_outputs[2324]) | (layer2_outputs[1432]);
    assign layer3_outputs[1674] = ~((layer2_outputs[2482]) & (layer2_outputs[1089]));
    assign layer3_outputs[1675] = ~(layer2_outputs[878]) | (layer2_outputs[1228]);
    assign layer3_outputs[1676] = ~(layer2_outputs[1005]);
    assign layer3_outputs[1677] = ~(layer2_outputs[215]) | (layer2_outputs[303]);
    assign layer3_outputs[1678] = (layer2_outputs[1349]) ^ (layer2_outputs[675]);
    assign layer3_outputs[1679] = ~((layer2_outputs[745]) ^ (layer2_outputs[1895]));
    assign layer3_outputs[1680] = (layer2_outputs[2304]) & (layer2_outputs[2367]);
    assign layer3_outputs[1681] = (layer2_outputs[836]) | (layer2_outputs[2515]);
    assign layer3_outputs[1682] = ~(layer2_outputs[918]) | (layer2_outputs[474]);
    assign layer3_outputs[1683] = layer2_outputs[999];
    assign layer3_outputs[1684] = ~(layer2_outputs[2163]);
    assign layer3_outputs[1685] = 1'b1;
    assign layer3_outputs[1686] = (layer2_outputs[2212]) | (layer2_outputs[2277]);
    assign layer3_outputs[1687] = layer2_outputs[2491];
    assign layer3_outputs[1688] = ~(layer2_outputs[724]);
    assign layer3_outputs[1689] = layer2_outputs[1326];
    assign layer3_outputs[1690] = (layer2_outputs[908]) & ~(layer2_outputs[2529]);
    assign layer3_outputs[1691] = ~((layer2_outputs[2431]) & (layer2_outputs[1246]));
    assign layer3_outputs[1692] = ~(layer2_outputs[1259]);
    assign layer3_outputs[1693] = layer2_outputs[2350];
    assign layer3_outputs[1694] = (layer2_outputs[2139]) ^ (layer2_outputs[1444]);
    assign layer3_outputs[1695] = (layer2_outputs[1841]) & (layer2_outputs[364]);
    assign layer3_outputs[1696] = layer2_outputs[2050];
    assign layer3_outputs[1697] = ~(layer2_outputs[1203]);
    assign layer3_outputs[1698] = layer2_outputs[1876];
    assign layer3_outputs[1699] = (layer2_outputs[225]) & (layer2_outputs[412]);
    assign layer3_outputs[1700] = ~(layer2_outputs[1277]);
    assign layer3_outputs[1701] = ~(layer2_outputs[2112]);
    assign layer3_outputs[1702] = (layer2_outputs[1504]) & ~(layer2_outputs[1430]);
    assign layer3_outputs[1703] = ~(layer2_outputs[928]);
    assign layer3_outputs[1704] = ~((layer2_outputs[2149]) ^ (layer2_outputs[731]));
    assign layer3_outputs[1705] = (layer2_outputs[425]) ^ (layer2_outputs[1957]);
    assign layer3_outputs[1706] = ~((layer2_outputs[332]) & (layer2_outputs[573]));
    assign layer3_outputs[1707] = (layer2_outputs[2199]) & ~(layer2_outputs[1123]);
    assign layer3_outputs[1708] = layer2_outputs[1558];
    assign layer3_outputs[1709] = ~(layer2_outputs[1903]);
    assign layer3_outputs[1710] = layer2_outputs[1835];
    assign layer3_outputs[1711] = layer2_outputs[565];
    assign layer3_outputs[1712] = ~((layer2_outputs[1285]) ^ (layer2_outputs[860]));
    assign layer3_outputs[1713] = (layer2_outputs[289]) ^ (layer2_outputs[667]);
    assign layer3_outputs[1714] = (layer2_outputs[446]) ^ (layer2_outputs[2503]);
    assign layer3_outputs[1715] = (layer2_outputs[1289]) & ~(layer2_outputs[2249]);
    assign layer3_outputs[1716] = layer2_outputs[1463];
    assign layer3_outputs[1717] = 1'b0;
    assign layer3_outputs[1718] = (layer2_outputs[1800]) & ~(layer2_outputs[661]);
    assign layer3_outputs[1719] = ~((layer2_outputs[1838]) ^ (layer2_outputs[1355]));
    assign layer3_outputs[1720] = (layer2_outputs[1736]) & ~(layer2_outputs[1794]);
    assign layer3_outputs[1721] = (layer2_outputs[678]) & ~(layer2_outputs[1916]);
    assign layer3_outputs[1722] = ~(layer2_outputs[2084]);
    assign layer3_outputs[1723] = ~((layer2_outputs[2261]) ^ (layer2_outputs[2042]));
    assign layer3_outputs[1724] = (layer2_outputs[696]) ^ (layer2_outputs[616]);
    assign layer3_outputs[1725] = ~((layer2_outputs[822]) ^ (layer2_outputs[1478]));
    assign layer3_outputs[1726] = (layer2_outputs[1036]) & ~(layer2_outputs[1254]);
    assign layer3_outputs[1727] = ~((layer2_outputs[2322]) ^ (layer2_outputs[858]));
    assign layer3_outputs[1728] = layer2_outputs[1878];
    assign layer3_outputs[1729] = ~(layer2_outputs[585]);
    assign layer3_outputs[1730] = (layer2_outputs[1151]) & ~(layer2_outputs[976]);
    assign layer3_outputs[1731] = (layer2_outputs[604]) | (layer2_outputs[918]);
    assign layer3_outputs[1732] = (layer2_outputs[1146]) | (layer2_outputs[227]);
    assign layer3_outputs[1733] = (layer2_outputs[2314]) & ~(layer2_outputs[2136]);
    assign layer3_outputs[1734] = ~(layer2_outputs[362]);
    assign layer3_outputs[1735] = layer2_outputs[409];
    assign layer3_outputs[1736] = (layer2_outputs[1865]) & ~(layer2_outputs[1241]);
    assign layer3_outputs[1737] = (layer2_outputs[1096]) & ~(layer2_outputs[1492]);
    assign layer3_outputs[1738] = layer2_outputs[2274];
    assign layer3_outputs[1739] = layer2_outputs[447];
    assign layer3_outputs[1740] = ~(layer2_outputs[1311]);
    assign layer3_outputs[1741] = ~(layer2_outputs[2046]) | (layer2_outputs[1866]);
    assign layer3_outputs[1742] = layer2_outputs[2104];
    assign layer3_outputs[1743] = ~(layer2_outputs[749]) | (layer2_outputs[1852]);
    assign layer3_outputs[1744] = ~((layer2_outputs[1146]) & (layer2_outputs[77]));
    assign layer3_outputs[1745] = layer2_outputs[2131];
    assign layer3_outputs[1746] = ~(layer2_outputs[1739]);
    assign layer3_outputs[1747] = ~(layer2_outputs[1557]) | (layer2_outputs[2492]);
    assign layer3_outputs[1748] = ~((layer2_outputs[1602]) & (layer2_outputs[1806]));
    assign layer3_outputs[1749] = ~(layer2_outputs[1428]) | (layer2_outputs[1595]);
    assign layer3_outputs[1750] = ~(layer2_outputs[2525]);
    assign layer3_outputs[1751] = ~(layer2_outputs[1647]);
    assign layer3_outputs[1752] = ~(layer2_outputs[923]);
    assign layer3_outputs[1753] = (layer2_outputs[1780]) & (layer2_outputs[2155]);
    assign layer3_outputs[1754] = layer2_outputs[1839];
    assign layer3_outputs[1755] = ~(layer2_outputs[2474]);
    assign layer3_outputs[1756] = (layer2_outputs[82]) & ~(layer2_outputs[1777]);
    assign layer3_outputs[1757] = 1'b0;
    assign layer3_outputs[1758] = 1'b1;
    assign layer3_outputs[1759] = ~(layer2_outputs[163]) | (layer2_outputs[470]);
    assign layer3_outputs[1760] = ~(layer2_outputs[1279]) | (layer2_outputs[301]);
    assign layer3_outputs[1761] = layer2_outputs[2230];
    assign layer3_outputs[1762] = ~((layer2_outputs[709]) & (layer2_outputs[1902]));
    assign layer3_outputs[1763] = ~(layer2_outputs[2163]);
    assign layer3_outputs[1764] = ~((layer2_outputs[1407]) & (layer2_outputs[629]));
    assign layer3_outputs[1765] = (layer2_outputs[2025]) ^ (layer2_outputs[2054]);
    assign layer3_outputs[1766] = ~((layer2_outputs[646]) & (layer2_outputs[732]));
    assign layer3_outputs[1767] = (layer2_outputs[720]) | (layer2_outputs[2395]);
    assign layer3_outputs[1768] = (layer2_outputs[1297]) & ~(layer2_outputs[1356]);
    assign layer3_outputs[1769] = ~(layer2_outputs[1759]);
    assign layer3_outputs[1770] = layer2_outputs[1922];
    assign layer3_outputs[1771] = ~(layer2_outputs[2002]);
    assign layer3_outputs[1772] = ~((layer2_outputs[31]) & (layer2_outputs[597]));
    assign layer3_outputs[1773] = ~(layer2_outputs[886]);
    assign layer3_outputs[1774] = (layer2_outputs[1638]) & ~(layer2_outputs[110]);
    assign layer3_outputs[1775] = (layer2_outputs[1670]) | (layer2_outputs[2346]);
    assign layer3_outputs[1776] = layer2_outputs[385];
    assign layer3_outputs[1777] = layer2_outputs[1186];
    assign layer3_outputs[1778] = layer2_outputs[493];
    assign layer3_outputs[1779] = ~((layer2_outputs[2311]) & (layer2_outputs[292]));
    assign layer3_outputs[1780] = ~((layer2_outputs[372]) | (layer2_outputs[199]));
    assign layer3_outputs[1781] = ~(layer2_outputs[2345]);
    assign layer3_outputs[1782] = (layer2_outputs[1852]) ^ (layer2_outputs[73]);
    assign layer3_outputs[1783] = ~((layer2_outputs[251]) & (layer2_outputs[1461]));
    assign layer3_outputs[1784] = ~(layer2_outputs[1496]);
    assign layer3_outputs[1785] = ~(layer2_outputs[1090]) | (layer2_outputs[1330]);
    assign layer3_outputs[1786] = (layer2_outputs[980]) & ~(layer2_outputs[390]);
    assign layer3_outputs[1787] = layer2_outputs[1341];
    assign layer3_outputs[1788] = layer2_outputs[2388];
    assign layer3_outputs[1789] = ~(layer2_outputs[590]);
    assign layer3_outputs[1790] = ~(layer2_outputs[1085]);
    assign layer3_outputs[1791] = (layer2_outputs[1933]) & ~(layer2_outputs[222]);
    assign layer3_outputs[1792] = (layer2_outputs[912]) ^ (layer2_outputs[1592]);
    assign layer3_outputs[1793] = (layer2_outputs[170]) | (layer2_outputs[394]);
    assign layer3_outputs[1794] = layer2_outputs[2480];
    assign layer3_outputs[1795] = (layer2_outputs[1490]) | (layer2_outputs[2268]);
    assign layer3_outputs[1796] = ~(layer2_outputs[2382]);
    assign layer3_outputs[1797] = (layer2_outputs[1032]) & (layer2_outputs[2082]);
    assign layer3_outputs[1798] = ~(layer2_outputs[2162]);
    assign layer3_outputs[1799] = layer2_outputs[241];
    assign layer3_outputs[1800] = (layer2_outputs[1176]) & ~(layer2_outputs[846]);
    assign layer3_outputs[1801] = ~((layer2_outputs[1969]) & (layer2_outputs[2181]));
    assign layer3_outputs[1802] = (layer2_outputs[72]) | (layer2_outputs[2531]);
    assign layer3_outputs[1803] = (layer2_outputs[1327]) & ~(layer2_outputs[2047]);
    assign layer3_outputs[1804] = ~((layer2_outputs[1583]) & (layer2_outputs[81]));
    assign layer3_outputs[1805] = ~(layer2_outputs[1849]);
    assign layer3_outputs[1806] = (layer2_outputs[2014]) & ~(layer2_outputs[1893]);
    assign layer3_outputs[1807] = (layer2_outputs[1433]) | (layer2_outputs[357]);
    assign layer3_outputs[1808] = layer2_outputs[1342];
    assign layer3_outputs[1809] = 1'b1;
    assign layer3_outputs[1810] = (layer2_outputs[657]) ^ (layer2_outputs[662]);
    assign layer3_outputs[1811] = (layer2_outputs[1947]) & ~(layer2_outputs[2302]);
    assign layer3_outputs[1812] = 1'b0;
    assign layer3_outputs[1813] = ~(layer2_outputs[223]);
    assign layer3_outputs[1814] = (layer2_outputs[1063]) & (layer2_outputs[42]);
    assign layer3_outputs[1815] = layer2_outputs[652];
    assign layer3_outputs[1816] = layer2_outputs[810];
    assign layer3_outputs[1817] = (layer2_outputs[1440]) & ~(layer2_outputs[139]);
    assign layer3_outputs[1818] = layer2_outputs[743];
    assign layer3_outputs[1819] = (layer2_outputs[1215]) & ~(layer2_outputs[604]);
    assign layer3_outputs[1820] = ~(layer2_outputs[1681]) | (layer2_outputs[1626]);
    assign layer3_outputs[1821] = ~(layer2_outputs[2420]) | (layer2_outputs[1593]);
    assign layer3_outputs[1822] = 1'b0;
    assign layer3_outputs[1823] = (layer2_outputs[585]) & ~(layer2_outputs[1240]);
    assign layer3_outputs[1824] = (layer2_outputs[913]) & (layer2_outputs[742]);
    assign layer3_outputs[1825] = ~(layer2_outputs[1227]);
    assign layer3_outputs[1826] = layer2_outputs[1694];
    assign layer3_outputs[1827] = ~((layer2_outputs[1833]) & (layer2_outputs[1199]));
    assign layer3_outputs[1828] = 1'b1;
    assign layer3_outputs[1829] = (layer2_outputs[2472]) & ~(layer2_outputs[2542]);
    assign layer3_outputs[1830] = (layer2_outputs[1633]) | (layer2_outputs[2170]);
    assign layer3_outputs[1831] = ~(layer2_outputs[235]);
    assign layer3_outputs[1832] = ~((layer2_outputs[1486]) & (layer2_outputs[1322]));
    assign layer3_outputs[1833] = (layer2_outputs[451]) & (layer2_outputs[2424]);
    assign layer3_outputs[1834] = ~(layer2_outputs[383]) | (layer2_outputs[818]);
    assign layer3_outputs[1835] = (layer2_outputs[19]) ^ (layer2_outputs[872]);
    assign layer3_outputs[1836] = ~(layer2_outputs[891]);
    assign layer3_outputs[1837] = layer2_outputs[136];
    assign layer3_outputs[1838] = (layer2_outputs[663]) ^ (layer2_outputs[1495]);
    assign layer3_outputs[1839] = ~(layer2_outputs[1905]);
    assign layer3_outputs[1840] = ~(layer2_outputs[2438]) | (layer2_outputs[875]);
    assign layer3_outputs[1841] = ~(layer2_outputs[668]) | (layer2_outputs[469]);
    assign layer3_outputs[1842] = ~((layer2_outputs[1125]) & (layer2_outputs[1742]));
    assign layer3_outputs[1843] = 1'b0;
    assign layer3_outputs[1844] = ~(layer2_outputs[1505]);
    assign layer3_outputs[1845] = (layer2_outputs[1712]) & ~(layer2_outputs[2373]);
    assign layer3_outputs[1846] = ~(layer2_outputs[2237]);
    assign layer3_outputs[1847] = layer2_outputs[2309];
    assign layer3_outputs[1848] = ~(layer2_outputs[146]);
    assign layer3_outputs[1849] = ~((layer2_outputs[1244]) | (layer2_outputs[151]));
    assign layer3_outputs[1850] = ~(layer2_outputs[961]);
    assign layer3_outputs[1851] = ~((layer2_outputs[738]) | (layer2_outputs[726]));
    assign layer3_outputs[1852] = (layer2_outputs[1718]) & (layer2_outputs[1448]);
    assign layer3_outputs[1853] = layer2_outputs[1920];
    assign layer3_outputs[1854] = 1'b0;
    assign layer3_outputs[1855] = layer2_outputs[1525];
    assign layer3_outputs[1856] = ~(layer2_outputs[299]);
    assign layer3_outputs[1857] = ~((layer2_outputs[1169]) & (layer2_outputs[876]));
    assign layer3_outputs[1858] = ~((layer2_outputs[2425]) | (layer2_outputs[641]));
    assign layer3_outputs[1859] = (layer2_outputs[1165]) & ~(layer2_outputs[1684]);
    assign layer3_outputs[1860] = ~(layer2_outputs[1938]);
    assign layer3_outputs[1861] = (layer2_outputs[1018]) & ~(layer2_outputs[1399]);
    assign layer3_outputs[1862] = 1'b0;
    assign layer3_outputs[1863] = 1'b1;
    assign layer3_outputs[1864] = (layer2_outputs[1154]) & ~(layer2_outputs[2539]);
    assign layer3_outputs[1865] = ~(layer2_outputs[229]) | (layer2_outputs[1546]);
    assign layer3_outputs[1866] = (layer2_outputs[821]) | (layer2_outputs[848]);
    assign layer3_outputs[1867] = ~((layer2_outputs[486]) & (layer2_outputs[2284]));
    assign layer3_outputs[1868] = layer2_outputs[2547];
    assign layer3_outputs[1869] = layer2_outputs[455];
    assign layer3_outputs[1870] = (layer2_outputs[736]) & (layer2_outputs[1752]);
    assign layer3_outputs[1871] = ~(layer2_outputs[855]) | (layer2_outputs[1521]);
    assign layer3_outputs[1872] = ~(layer2_outputs[212]);
    assign layer3_outputs[1873] = ~(layer2_outputs[832]);
    assign layer3_outputs[1874] = layer2_outputs[221];
    assign layer3_outputs[1875] = layer2_outputs[2352];
    assign layer3_outputs[1876] = (layer2_outputs[189]) & ~(layer2_outputs[1024]);
    assign layer3_outputs[1877] = ~(layer2_outputs[719]);
    assign layer3_outputs[1878] = (layer2_outputs[1058]) ^ (layer2_outputs[656]);
    assign layer3_outputs[1879] = layer2_outputs[1145];
    assign layer3_outputs[1880] = (layer2_outputs[394]) & (layer2_outputs[1204]);
    assign layer3_outputs[1881] = ~((layer2_outputs[722]) | (layer2_outputs[723]));
    assign layer3_outputs[1882] = ~(layer2_outputs[199]);
    assign layer3_outputs[1883] = layer2_outputs[1872];
    assign layer3_outputs[1884] = layer2_outputs[131];
    assign layer3_outputs[1885] = 1'b1;
    assign layer3_outputs[1886] = ~(layer2_outputs[2007]);
    assign layer3_outputs[1887] = ~(layer2_outputs[607]) | (layer2_outputs[1114]);
    assign layer3_outputs[1888] = ~(layer2_outputs[721]);
    assign layer3_outputs[1889] = ~(layer2_outputs[1610]);
    assign layer3_outputs[1890] = (layer2_outputs[1275]) & (layer2_outputs[1723]);
    assign layer3_outputs[1891] = layer2_outputs[1449];
    assign layer3_outputs[1892] = layer2_outputs[1868];
    assign layer3_outputs[1893] = layer2_outputs[1466];
    assign layer3_outputs[1894] = layer2_outputs[1286];
    assign layer3_outputs[1895] = ~((layer2_outputs[1669]) | (layer2_outputs[23]));
    assign layer3_outputs[1896] = ~(layer2_outputs[265]);
    assign layer3_outputs[1897] = layer2_outputs[2518];
    assign layer3_outputs[1898] = ~((layer2_outputs[1062]) | (layer2_outputs[1053]));
    assign layer3_outputs[1899] = ~((layer2_outputs[481]) & (layer2_outputs[1938]));
    assign layer3_outputs[1900] = ~((layer2_outputs[458]) ^ (layer2_outputs[1133]));
    assign layer3_outputs[1901] = ~(layer2_outputs[1027]) | (layer2_outputs[2389]);
    assign layer3_outputs[1902] = ~((layer2_outputs[1648]) & (layer2_outputs[2030]));
    assign layer3_outputs[1903] = ~(layer2_outputs[1467]);
    assign layer3_outputs[1904] = ~(layer2_outputs[2153]) | (layer2_outputs[819]);
    assign layer3_outputs[1905] = ~(layer2_outputs[27]);
    assign layer3_outputs[1906] = (layer2_outputs[744]) & (layer2_outputs[1571]);
    assign layer3_outputs[1907] = ~((layer2_outputs[328]) & (layer2_outputs[2294]));
    assign layer3_outputs[1908] = layer2_outputs[999];
    assign layer3_outputs[1909] = ~(layer2_outputs[1698]) | (layer2_outputs[1590]);
    assign layer3_outputs[1910] = (layer2_outputs[1651]) & ~(layer2_outputs[1580]);
    assign layer3_outputs[1911] = (layer2_outputs[1082]) | (layer2_outputs[2517]);
    assign layer3_outputs[1912] = layer2_outputs[2057];
    assign layer3_outputs[1913] = ~((layer2_outputs[760]) & (layer2_outputs[1020]));
    assign layer3_outputs[1914] = (layer2_outputs[1952]) & ~(layer2_outputs[687]);
    assign layer3_outputs[1915] = (layer2_outputs[145]) | (layer2_outputs[1727]);
    assign layer3_outputs[1916] = layer2_outputs[2224];
    assign layer3_outputs[1917] = layer2_outputs[1671];
    assign layer3_outputs[1918] = ~(layer2_outputs[2234]) | (layer2_outputs[1017]);
    assign layer3_outputs[1919] = (layer2_outputs[573]) & ~(layer2_outputs[443]);
    assign layer3_outputs[1920] = ~((layer2_outputs[770]) & (layer2_outputs[352]));
    assign layer3_outputs[1921] = (layer2_outputs[92]) | (layer2_outputs[1835]);
    assign layer3_outputs[1922] = layer2_outputs[1517];
    assign layer3_outputs[1923] = ~(layer2_outputs[515]);
    assign layer3_outputs[1924] = ~((layer2_outputs[850]) & (layer2_outputs[929]));
    assign layer3_outputs[1925] = ~((layer2_outputs[380]) | (layer2_outputs[2079]));
    assign layer3_outputs[1926] = (layer2_outputs[1989]) & ~(layer2_outputs[639]);
    assign layer3_outputs[1927] = (layer2_outputs[1181]) | (layer2_outputs[1832]);
    assign layer3_outputs[1928] = ~((layer2_outputs[454]) | (layer2_outputs[18]));
    assign layer3_outputs[1929] = (layer2_outputs[2207]) ^ (layer2_outputs[1310]);
    assign layer3_outputs[1930] = layer2_outputs[895];
    assign layer3_outputs[1931] = (layer2_outputs[1745]) & ~(layer2_outputs[1105]);
    assign layer3_outputs[1932] = ~(layer2_outputs[723]) | (layer2_outputs[1026]);
    assign layer3_outputs[1933] = layer2_outputs[330];
    assign layer3_outputs[1934] = ~((layer2_outputs[408]) & (layer2_outputs[811]));
    assign layer3_outputs[1935] = ~(layer2_outputs[1934]) | (layer2_outputs[1475]);
    assign layer3_outputs[1936] = layer2_outputs[2506];
    assign layer3_outputs[1937] = layer2_outputs[2284];
    assign layer3_outputs[1938] = ~((layer2_outputs[924]) ^ (layer2_outputs[594]));
    assign layer3_outputs[1939] = ~(layer2_outputs[697]) | (layer2_outputs[1741]);
    assign layer3_outputs[1940] = layer2_outputs[2020];
    assign layer3_outputs[1941] = ~(layer2_outputs[2465]);
    assign layer3_outputs[1942] = layer2_outputs[2473];
    assign layer3_outputs[1943] = ~(layer2_outputs[1250]) | (layer2_outputs[1983]);
    assign layer3_outputs[1944] = ~((layer2_outputs[367]) ^ (layer2_outputs[1866]));
    assign layer3_outputs[1945] = (layer2_outputs[1648]) & ~(layer2_outputs[1349]);
    assign layer3_outputs[1946] = ~(layer2_outputs[450]);
    assign layer3_outputs[1947] = layer2_outputs[2254];
    assign layer3_outputs[1948] = ~(layer2_outputs[2236]);
    assign layer3_outputs[1949] = ~((layer2_outputs[50]) | (layer2_outputs[1660]));
    assign layer3_outputs[1950] = (layer2_outputs[2044]) | (layer2_outputs[2328]);
    assign layer3_outputs[1951] = ~((layer2_outputs[2108]) | (layer2_outputs[1968]));
    assign layer3_outputs[1952] = (layer2_outputs[1848]) | (layer2_outputs[1070]);
    assign layer3_outputs[1953] = layer2_outputs[926];
    assign layer3_outputs[1954] = ~(layer2_outputs[181]);
    assign layer3_outputs[1955] = layer2_outputs[112];
    assign layer3_outputs[1956] = 1'b0;
    assign layer3_outputs[1957] = layer2_outputs[508];
    assign layer3_outputs[1958] = (layer2_outputs[180]) | (layer2_outputs[452]);
    assign layer3_outputs[1959] = ~(layer2_outputs[1765]);
    assign layer3_outputs[1960] = (layer2_outputs[1964]) & ~(layer2_outputs[1827]);
    assign layer3_outputs[1961] = (layer2_outputs[1830]) ^ (layer2_outputs[1620]);
    assign layer3_outputs[1962] = ~(layer2_outputs[800]);
    assign layer3_outputs[1963] = layer2_outputs[1508];
    assign layer3_outputs[1964] = layer2_outputs[1888];
    assign layer3_outputs[1965] = (layer2_outputs[582]) | (layer2_outputs[529]);
    assign layer3_outputs[1966] = ~((layer2_outputs[882]) | (layer2_outputs[882]));
    assign layer3_outputs[1967] = layer2_outputs[248];
    assign layer3_outputs[1968] = ~(layer2_outputs[382]);
    assign layer3_outputs[1969] = ~((layer2_outputs[1434]) & (layer2_outputs[907]));
    assign layer3_outputs[1970] = layer2_outputs[1503];
    assign layer3_outputs[1971] = ~((layer2_outputs[841]) | (layer2_outputs[1168]));
    assign layer3_outputs[1972] = ~(layer2_outputs[1057]);
    assign layer3_outputs[1973] = (layer2_outputs[337]) & ~(layer2_outputs[621]);
    assign layer3_outputs[1974] = ~(layer2_outputs[2135]);
    assign layer3_outputs[1975] = (layer2_outputs[2510]) | (layer2_outputs[1022]);
    assign layer3_outputs[1976] = (layer2_outputs[887]) & (layer2_outputs[284]);
    assign layer3_outputs[1977] = (layer2_outputs[272]) | (layer2_outputs[890]);
    assign layer3_outputs[1978] = layer2_outputs[1209];
    assign layer3_outputs[1979] = (layer2_outputs[1198]) & (layer2_outputs[1207]);
    assign layer3_outputs[1980] = ~(layer2_outputs[925]);
    assign layer3_outputs[1981] = layer2_outputs[1686];
    assign layer3_outputs[1982] = layer2_outputs[2354];
    assign layer3_outputs[1983] = (layer2_outputs[2008]) ^ (layer2_outputs[1640]);
    assign layer3_outputs[1984] = ~(layer2_outputs[2505]) | (layer2_outputs[747]);
    assign layer3_outputs[1985] = layer2_outputs[778];
    assign layer3_outputs[1986] = ~(layer2_outputs[2340]);
    assign layer3_outputs[1987] = 1'b1;
    assign layer3_outputs[1988] = ~(layer2_outputs[1953]);
    assign layer3_outputs[1989] = ~(layer2_outputs[2196]);
    assign layer3_outputs[1990] = (layer2_outputs[157]) ^ (layer2_outputs[625]);
    assign layer3_outputs[1991] = ~(layer2_outputs[2251]) | (layer2_outputs[407]);
    assign layer3_outputs[1992] = 1'b1;
    assign layer3_outputs[1993] = ~(layer2_outputs[2325]);
    assign layer3_outputs[1994] = (layer2_outputs[2380]) & ~(layer2_outputs[1603]);
    assign layer3_outputs[1995] = (layer2_outputs[694]) & ~(layer2_outputs[2559]);
    assign layer3_outputs[1996] = (layer2_outputs[1779]) & (layer2_outputs[2316]);
    assign layer3_outputs[1997] = (layer2_outputs[1945]) | (layer2_outputs[553]);
    assign layer3_outputs[1998] = layer2_outputs[2330];
    assign layer3_outputs[1999] = ~((layer2_outputs[1408]) | (layer2_outputs[55]));
    assign layer3_outputs[2000] = (layer2_outputs[826]) | (layer2_outputs[1314]);
    assign layer3_outputs[2001] = ~(layer2_outputs[432]);
    assign layer3_outputs[2002] = 1'b1;
    assign layer3_outputs[2003] = ~(layer2_outputs[224]) | (layer2_outputs[41]);
    assign layer3_outputs[2004] = (layer2_outputs[1915]) & ~(layer2_outputs[1639]);
    assign layer3_outputs[2005] = ~(layer2_outputs[354]);
    assign layer3_outputs[2006] = ~(layer2_outputs[699]);
    assign layer3_outputs[2007] = layer2_outputs[1313];
    assign layer3_outputs[2008] = layer2_outputs[2064];
    assign layer3_outputs[2009] = layer2_outputs[1126];
    assign layer3_outputs[2010] = ~(layer2_outputs[127]) | (layer2_outputs[652]);
    assign layer3_outputs[2011] = layer2_outputs[1561];
    assign layer3_outputs[2012] = ~((layer2_outputs[1993]) | (layer2_outputs[2487]));
    assign layer3_outputs[2013] = ~((layer2_outputs[835]) & (layer2_outputs[2368]));
    assign layer3_outputs[2014] = 1'b0;
    assign layer3_outputs[2015] = ~((layer2_outputs[1560]) ^ (layer2_outputs[100]));
    assign layer3_outputs[2016] = (layer2_outputs[776]) & ~(layer2_outputs[146]);
    assign layer3_outputs[2017] = layer2_outputs[898];
    assign layer3_outputs[2018] = layer2_outputs[2295];
    assign layer3_outputs[2019] = 1'b0;
    assign layer3_outputs[2020] = ~(layer2_outputs[1397]);
    assign layer3_outputs[2021] = layer2_outputs[1998];
    assign layer3_outputs[2022] = ~((layer2_outputs[1948]) | (layer2_outputs[511]));
    assign layer3_outputs[2023] = layer2_outputs[523];
    assign layer3_outputs[2024] = (layer2_outputs[2241]) & ~(layer2_outputs[1619]);
    assign layer3_outputs[2025] = layer2_outputs[414];
    assign layer3_outputs[2026] = ~((layer2_outputs[1814]) & (layer2_outputs[1913]));
    assign layer3_outputs[2027] = ~(layer2_outputs[2559]) | (layer2_outputs[2396]);
    assign layer3_outputs[2028] = (layer2_outputs[826]) & ~(layer2_outputs[561]);
    assign layer3_outputs[2029] = (layer2_outputs[1552]) ^ (layer2_outputs[1430]);
    assign layer3_outputs[2030] = ~((layer2_outputs[316]) ^ (layer2_outputs[973]));
    assign layer3_outputs[2031] = (layer2_outputs[637]) & (layer2_outputs[824]);
    assign layer3_outputs[2032] = ~((layer2_outputs[2164]) | (layer2_outputs[1653]));
    assign layer3_outputs[2033] = ~((layer2_outputs[1013]) ^ (layer2_outputs[2471]));
    assign layer3_outputs[2034] = ~(layer2_outputs[273]);
    assign layer3_outputs[2035] = ~((layer2_outputs[150]) & (layer2_outputs[913]));
    assign layer3_outputs[2036] = layer2_outputs[1288];
    assign layer3_outputs[2037] = ~((layer2_outputs[438]) | (layer2_outputs[2283]));
    assign layer3_outputs[2038] = ~((layer2_outputs[1308]) ^ (layer2_outputs[1177]));
    assign layer3_outputs[2039] = layer2_outputs[1894];
    assign layer3_outputs[2040] = layer2_outputs[436];
    assign layer3_outputs[2041] = layer2_outputs[515];
    assign layer3_outputs[2042] = ~(layer2_outputs[2151]) | (layer2_outputs[2077]);
    assign layer3_outputs[2043] = ~(layer2_outputs[88]) | (layer2_outputs[107]);
    assign layer3_outputs[2044] = (layer2_outputs[2154]) | (layer2_outputs[2105]);
    assign layer3_outputs[2045] = ~(layer2_outputs[563]) | (layer2_outputs[47]);
    assign layer3_outputs[2046] = (layer2_outputs[1359]) | (layer2_outputs[975]);
    assign layer3_outputs[2047] = ~(layer2_outputs[926]);
    assign layer3_outputs[2048] = ~(layer2_outputs[1370]);
    assign layer3_outputs[2049] = (layer2_outputs[1740]) | (layer2_outputs[270]);
    assign layer3_outputs[2050] = ~(layer2_outputs[1012]);
    assign layer3_outputs[2051] = ~(layer2_outputs[1954]);
    assign layer3_outputs[2052] = layer2_outputs[218];
    assign layer3_outputs[2053] = ~(layer2_outputs[521]);
    assign layer3_outputs[2054] = layer2_outputs[1646];
    assign layer3_outputs[2055] = ~(layer2_outputs[512]);
    assign layer3_outputs[2056] = layer2_outputs[1400];
    assign layer3_outputs[2057] = (layer2_outputs[2099]) & (layer2_outputs[2546]);
    assign layer3_outputs[2058] = ~(layer2_outputs[1605]);
    assign layer3_outputs[2059] = ~(layer2_outputs[233]);
    assign layer3_outputs[2060] = 1'b1;
    assign layer3_outputs[2061] = layer2_outputs[133];
    assign layer3_outputs[2062] = (layer2_outputs[1009]) ^ (layer2_outputs[2555]);
    assign layer3_outputs[2063] = ~((layer2_outputs[300]) | (layer2_outputs[2551]));
    assign layer3_outputs[2064] = (layer2_outputs[1392]) & ~(layer2_outputs[1792]);
    assign layer3_outputs[2065] = ~(layer2_outputs[1791]);
    assign layer3_outputs[2066] = (layer2_outputs[128]) | (layer2_outputs[2087]);
    assign layer3_outputs[2067] = layer2_outputs[1910];
    assign layer3_outputs[2068] = (layer2_outputs[789]) & ~(layer2_outputs[1139]);
    assign layer3_outputs[2069] = ~(layer2_outputs[680]) | (layer2_outputs[1613]);
    assign layer3_outputs[2070] = layer2_outputs[2074];
    assign layer3_outputs[2071] = (layer2_outputs[2489]) ^ (layer2_outputs[1425]);
    assign layer3_outputs[2072] = layer2_outputs[1415];
    assign layer3_outputs[2073] = (layer2_outputs[0]) & ~(layer2_outputs[1501]);
    assign layer3_outputs[2074] = (layer2_outputs[245]) & ~(layer2_outputs[1864]);
    assign layer3_outputs[2075] = layer2_outputs[1512];
    assign layer3_outputs[2076] = ~(layer2_outputs[360]);
    assign layer3_outputs[2077] = ~((layer2_outputs[613]) ^ (layer2_outputs[2043]));
    assign layer3_outputs[2078] = ~((layer2_outputs[1685]) ^ (layer2_outputs[1029]));
    assign layer3_outputs[2079] = ~(layer2_outputs[2456]) | (layer2_outputs[2225]);
    assign layer3_outputs[2080] = ~(layer2_outputs[2174]);
    assign layer3_outputs[2081] = (layer2_outputs[1375]) & (layer2_outputs[2327]);
    assign layer3_outputs[2082] = (layer2_outputs[2106]) ^ (layer2_outputs[1331]);
    assign layer3_outputs[2083] = ~((layer2_outputs[1628]) ^ (layer2_outputs[1909]));
    assign layer3_outputs[2084] = ~(layer2_outputs[2169]);
    assign layer3_outputs[2085] = ~(layer2_outputs[342]);
    assign layer3_outputs[2086] = layer2_outputs[34];
    assign layer3_outputs[2087] = ~(layer2_outputs[702]);
    assign layer3_outputs[2088] = (layer2_outputs[1205]) ^ (layer2_outputs[2530]);
    assign layer3_outputs[2089] = (layer2_outputs[1966]) | (layer2_outputs[2035]);
    assign layer3_outputs[2090] = ~((layer2_outputs[743]) | (layer2_outputs[1301]));
    assign layer3_outputs[2091] = 1'b0;
    assign layer3_outputs[2092] = ~((layer2_outputs[1635]) | (layer2_outputs[172]));
    assign layer3_outputs[2093] = (layer2_outputs[2051]) & (layer2_outputs[1869]);
    assign layer3_outputs[2094] = ~(layer2_outputs[78]) | (layer2_outputs[1352]);
    assign layer3_outputs[2095] = (layer2_outputs[2124]) & (layer2_outputs[1624]);
    assign layer3_outputs[2096] = (layer2_outputs[341]) & ~(layer2_outputs[2488]);
    assign layer3_outputs[2097] = layer2_outputs[1447];
    assign layer3_outputs[2098] = (layer2_outputs[1273]) ^ (layer2_outputs[1048]);
    assign layer3_outputs[2099] = layer2_outputs[1958];
    assign layer3_outputs[2100] = layer2_outputs[1243];
    assign layer3_outputs[2101] = ~((layer2_outputs[1403]) ^ (layer2_outputs[2084]));
    assign layer3_outputs[2102] = ~(layer2_outputs[1234]) | (layer2_outputs[1382]);
    assign layer3_outputs[2103] = ~(layer2_outputs[1182]);
    assign layer3_outputs[2104] = ~(layer2_outputs[1456]);
    assign layer3_outputs[2105] = ~(layer2_outputs[799]) | (layer2_outputs[1551]);
    assign layer3_outputs[2106] = (layer2_outputs[631]) | (layer2_outputs[2276]);
    assign layer3_outputs[2107] = ~(layer2_outputs[1262]) | (layer2_outputs[2281]);
    assign layer3_outputs[2108] = layer2_outputs[2053];
    assign layer3_outputs[2109] = layer2_outputs[449];
    assign layer3_outputs[2110] = layer2_outputs[2402];
    assign layer3_outputs[2111] = (layer2_outputs[957]) & (layer2_outputs[2102]);
    assign layer3_outputs[2112] = ~(layer2_outputs[758]) | (layer2_outputs[1149]);
    assign layer3_outputs[2113] = ~(layer2_outputs[1131]);
    assign layer3_outputs[2114] = layer2_outputs[1332];
    assign layer3_outputs[2115] = ~(layer2_outputs[1921]) | (layer2_outputs[1435]);
    assign layer3_outputs[2116] = ~(layer2_outputs[30]) | (layer2_outputs[1707]);
    assign layer3_outputs[2117] = layer2_outputs[2266];
    assign layer3_outputs[2118] = ~(layer2_outputs[1930]) | (layer2_outputs[777]);
    assign layer3_outputs[2119] = layer2_outputs[1437];
    assign layer3_outputs[2120] = (layer2_outputs[2056]) ^ (layer2_outputs[228]);
    assign layer3_outputs[2121] = ~(layer2_outputs[2276]);
    assign layer3_outputs[2122] = layer2_outputs[2458];
    assign layer3_outputs[2123] = (layer2_outputs[1100]) & ~(layer2_outputs[46]);
    assign layer3_outputs[2124] = ~(layer2_outputs[1843]) | (layer2_outputs[277]);
    assign layer3_outputs[2125] = ~(layer2_outputs[1816]);
    assign layer3_outputs[2126] = ~(layer2_outputs[2026]);
    assign layer3_outputs[2127] = ~(layer2_outputs[193]);
    assign layer3_outputs[2128] = (layer2_outputs[1876]) & ~(layer2_outputs[1687]);
    assign layer3_outputs[2129] = ~(layer2_outputs[1195]);
    assign layer3_outputs[2130] = layer2_outputs[1882];
    assign layer3_outputs[2131] = (layer2_outputs[2468]) ^ (layer2_outputs[1260]);
    assign layer3_outputs[2132] = 1'b0;
    assign layer3_outputs[2133] = ~(layer2_outputs[1239]);
    assign layer3_outputs[2134] = (layer2_outputs[1453]) ^ (layer2_outputs[1370]);
    assign layer3_outputs[2135] = ~(layer2_outputs[958]) | (layer2_outputs[2501]);
    assign layer3_outputs[2136] = layer2_outputs[773];
    assign layer3_outputs[2137] = ~((layer2_outputs[2156]) | (layer2_outputs[863]));
    assign layer3_outputs[2138] = (layer2_outputs[1098]) & ~(layer2_outputs[1574]);
    assign layer3_outputs[2139] = ~((layer2_outputs[969]) | (layer2_outputs[311]));
    assign layer3_outputs[2140] = ~(layer2_outputs[1044]);
    assign layer3_outputs[2141] = 1'b0;
    assign layer3_outputs[2142] = ~(layer2_outputs[419]) | (layer2_outputs[2349]);
    assign layer3_outputs[2143] = ~(layer2_outputs[1160]) | (layer2_outputs[413]);
    assign layer3_outputs[2144] = layer2_outputs[1473];
    assign layer3_outputs[2145] = (layer2_outputs[1514]) & ~(layer2_outputs[174]);
    assign layer3_outputs[2146] = (layer2_outputs[817]) & ~(layer2_outputs[28]);
    assign layer3_outputs[2147] = ~((layer2_outputs[768]) & (layer2_outputs[108]));
    assign layer3_outputs[2148] = 1'b0;
    assign layer3_outputs[2149] = (layer2_outputs[2286]) & (layer2_outputs[1873]);
    assign layer3_outputs[2150] = (layer2_outputs[2239]) & (layer2_outputs[2493]);
    assign layer3_outputs[2151] = 1'b1;
    assign layer3_outputs[2152] = (layer2_outputs[752]) | (layer2_outputs[70]);
    assign layer3_outputs[2153] = (layer2_outputs[1454]) & ~(layer2_outputs[83]);
    assign layer3_outputs[2154] = ~((layer2_outputs[833]) | (layer2_outputs[2422]));
    assign layer3_outputs[2155] = ~(layer2_outputs[579]);
    assign layer3_outputs[2156] = (layer2_outputs[948]) | (layer2_outputs[1484]);
    assign layer3_outputs[2157] = layer2_outputs[872];
    assign layer3_outputs[2158] = (layer2_outputs[351]) & (layer2_outputs[520]);
    assign layer3_outputs[2159] = ~(layer2_outputs[2358]);
    assign layer3_outputs[2160] = layer2_outputs[1023];
    assign layer3_outputs[2161] = (layer2_outputs[975]) & (layer2_outputs[9]);
    assign layer3_outputs[2162] = ~(layer2_outputs[1337]) | (layer2_outputs[1211]);
    assign layer3_outputs[2163] = (layer2_outputs[1594]) | (layer2_outputs[231]);
    assign layer3_outputs[2164] = (layer2_outputs[97]) ^ (layer2_outputs[436]);
    assign layer3_outputs[2165] = ~(layer2_outputs[1214]);
    assign layer3_outputs[2166] = (layer2_outputs[611]) & ~(layer2_outputs[662]);
    assign layer3_outputs[2167] = ~((layer2_outputs[2210]) ^ (layer2_outputs[73]));
    assign layer3_outputs[2168] = ~((layer2_outputs[694]) & (layer2_outputs[1928]));
    assign layer3_outputs[2169] = 1'b0;
    assign layer3_outputs[2170] = ~(layer2_outputs[1366]) | (layer2_outputs[1672]);
    assign layer3_outputs[2171] = ~(layer2_outputs[1704]) | (layer2_outputs[691]);
    assign layer3_outputs[2172] = ~(layer2_outputs[877]);
    assign layer3_outputs[2173] = (layer2_outputs[957]) & ~(layer2_outputs[2253]);
    assign layer3_outputs[2174] = ~((layer2_outputs[2486]) ^ (layer2_outputs[1355]));
    assign layer3_outputs[2175] = ~(layer2_outputs[1900]) | (layer2_outputs[1401]);
    assign layer3_outputs[2176] = ~((layer2_outputs[640]) ^ (layer2_outputs[1543]));
    assign layer3_outputs[2177] = ~(layer2_outputs[2262]);
    assign layer3_outputs[2178] = (layer2_outputs[561]) & (layer2_outputs[702]);
    assign layer3_outputs[2179] = ~(layer2_outputs[1650]) | (layer2_outputs[570]);
    assign layer3_outputs[2180] = ~(layer2_outputs[1142]);
    assign layer3_outputs[2181] = (layer2_outputs[340]) ^ (layer2_outputs[1662]);
    assign layer3_outputs[2182] = ~(layer2_outputs[1175]);
    assign layer3_outputs[2183] = (layer2_outputs[877]) ^ (layer2_outputs[2098]);
    assign layer3_outputs[2184] = ~((layer2_outputs[177]) | (layer2_outputs[2451]));
    assign layer3_outputs[2185] = 1'b1;
    assign layer3_outputs[2186] = layer2_outputs[2525];
    assign layer3_outputs[2187] = (layer2_outputs[341]) & ~(layer2_outputs[1993]);
    assign layer3_outputs[2188] = (layer2_outputs[1434]) & ~(layer2_outputs[85]);
    assign layer3_outputs[2189] = (layer2_outputs[1906]) | (layer2_outputs[2148]);
    assign layer3_outputs[2190] = layer2_outputs[363];
    assign layer3_outputs[2191] = ~((layer2_outputs[871]) | (layer2_outputs[914]));
    assign layer3_outputs[2192] = ~(layer2_outputs[881]) | (layer2_outputs[536]);
    assign layer3_outputs[2193] = ~((layer2_outputs[1378]) & (layer2_outputs[1986]));
    assign layer3_outputs[2194] = ~(layer2_outputs[674]);
    assign layer3_outputs[2195] = (layer2_outputs[517]) ^ (layer2_outputs[2129]);
    assign layer3_outputs[2196] = ~(layer2_outputs[494]) | (layer2_outputs[748]);
    assign layer3_outputs[2197] = ~(layer2_outputs[214]);
    assign layer3_outputs[2198] = ~(layer2_outputs[1918]) | (layer2_outputs[879]);
    assign layer3_outputs[2199] = layer2_outputs[983];
    assign layer3_outputs[2200] = layer2_outputs[783];
    assign layer3_outputs[2201] = (layer2_outputs[2152]) & ~(layer2_outputs[1682]);
    assign layer3_outputs[2202] = ~(layer2_outputs[1790]);
    assign layer3_outputs[2203] = ~((layer2_outputs[1585]) & (layer2_outputs[294]));
    assign layer3_outputs[2204] = ~((layer2_outputs[1067]) & (layer2_outputs[1869]));
    assign layer3_outputs[2205] = layer2_outputs[686];
    assign layer3_outputs[2206] = 1'b1;
    assign layer3_outputs[2207] = layer2_outputs[1302];
    assign layer3_outputs[2208] = ~((layer2_outputs[376]) | (layer2_outputs[1445]));
    assign layer3_outputs[2209] = ~(layer2_outputs[1911]);
    assign layer3_outputs[2210] = 1'b0;
    assign layer3_outputs[2211] = (layer2_outputs[389]) & ~(layer2_outputs[1862]);
    assign layer3_outputs[2212] = ~(layer2_outputs[104]);
    assign layer3_outputs[2213] = layer2_outputs[969];
    assign layer3_outputs[2214] = (layer2_outputs[383]) ^ (layer2_outputs[2257]);
    assign layer3_outputs[2215] = ~(layer2_outputs[1689]) | (layer2_outputs[1122]);
    assign layer3_outputs[2216] = layer2_outputs[1751];
    assign layer3_outputs[2217] = ~(layer2_outputs[2224]);
    assign layer3_outputs[2218] = ~((layer2_outputs[25]) ^ (layer2_outputs[715]));
    assign layer3_outputs[2219] = 1'b1;
    assign layer3_outputs[2220] = (layer2_outputs[1581]) & (layer2_outputs[1494]);
    assign layer3_outputs[2221] = ~(layer2_outputs[419]);
    assign layer3_outputs[2222] = layer2_outputs[1579];
    assign layer3_outputs[2223] = (layer2_outputs[1803]) | (layer2_outputs[267]);
    assign layer3_outputs[2224] = (layer2_outputs[1231]) ^ (layer2_outputs[1566]);
    assign layer3_outputs[2225] = layer2_outputs[1458];
    assign layer3_outputs[2226] = layer2_outputs[139];
    assign layer3_outputs[2227] = ~((layer2_outputs[2248]) ^ (layer2_outputs[1534]));
    assign layer3_outputs[2228] = ~(layer2_outputs[277]) | (layer2_outputs[785]);
    assign layer3_outputs[2229] = ~(layer2_outputs[1167]);
    assign layer3_outputs[2230] = ~(layer2_outputs[1424]);
    assign layer3_outputs[2231] = ~(layer2_outputs[2410]);
    assign layer3_outputs[2232] = ~(layer2_outputs[797]);
    assign layer3_outputs[2233] = layer2_outputs[677];
    assign layer3_outputs[2234] = ~((layer2_outputs[962]) | (layer2_outputs[775]));
    assign layer3_outputs[2235] = (layer2_outputs[1238]) & (layer2_outputs[843]);
    assign layer3_outputs[2236] = layer2_outputs[1407];
    assign layer3_outputs[2237] = layer2_outputs[2315];
    assign layer3_outputs[2238] = ~((layer2_outputs[2362]) | (layer2_outputs[1588]));
    assign layer3_outputs[2239] = (layer2_outputs[1269]) & ~(layer2_outputs[325]);
    assign layer3_outputs[2240] = layer2_outputs[1148];
    assign layer3_outputs[2241] = layer2_outputs[528];
    assign layer3_outputs[2242] = layer2_outputs[39];
    assign layer3_outputs[2243] = layer2_outputs[1796];
    assign layer3_outputs[2244] = ~((layer2_outputs[2255]) ^ (layer2_outputs[2053]));
    assign layer3_outputs[2245] = ~(layer2_outputs[124]);
    assign layer3_outputs[2246] = (layer2_outputs[260]) & ~(layer2_outputs[1152]);
    assign layer3_outputs[2247] = layer2_outputs[1026];
    assign layer3_outputs[2248] = layer2_outputs[598];
    assign layer3_outputs[2249] = ~(layer2_outputs[539]);
    assign layer3_outputs[2250] = ~(layer2_outputs[1688]) | (layer2_outputs[477]);
    assign layer3_outputs[2251] = ~(layer2_outputs[1076]);
    assign layer3_outputs[2252] = ~(layer2_outputs[1022]);
    assign layer3_outputs[2253] = (layer2_outputs[284]) & ~(layer2_outputs[17]);
    assign layer3_outputs[2254] = layer2_outputs[46];
    assign layer3_outputs[2255] = layer2_outputs[1222];
    assign layer3_outputs[2256] = layer2_outputs[793];
    assign layer3_outputs[2257] = layer2_outputs[1385];
    assign layer3_outputs[2258] = ~(layer2_outputs[1787]);
    assign layer3_outputs[2259] = (layer2_outputs[1594]) & (layer2_outputs[437]);
    assign layer3_outputs[2260] = layer2_outputs[1280];
    assign layer3_outputs[2261] = ~((layer2_outputs[102]) | (layer2_outputs[883]));
    assign layer3_outputs[2262] = layer2_outputs[530];
    assign layer3_outputs[2263] = layer2_outputs[594];
    assign layer3_outputs[2264] = layer2_outputs[1862];
    assign layer3_outputs[2265] = layer2_outputs[366];
    assign layer3_outputs[2266] = ~(layer2_outputs[60]) | (layer2_outputs[1008]);
    assign layer3_outputs[2267] = ~(layer2_outputs[2475]);
    assign layer3_outputs[2268] = (layer2_outputs[1255]) & (layer2_outputs[1103]);
    assign layer3_outputs[2269] = 1'b0;
    assign layer3_outputs[2270] = layer2_outputs[2336];
    assign layer3_outputs[2271] = (layer2_outputs[518]) & (layer2_outputs[1423]);
    assign layer3_outputs[2272] = ~((layer2_outputs[2073]) & (layer2_outputs[205]));
    assign layer3_outputs[2273] = (layer2_outputs[1451]) & ~(layer2_outputs[11]);
    assign layer3_outputs[2274] = ~((layer2_outputs[2231]) & (layer2_outputs[2463]));
    assign layer3_outputs[2275] = layer2_outputs[763];
    assign layer3_outputs[2276] = ~(layer2_outputs[427]) | (layer2_outputs[2476]);
    assign layer3_outputs[2277] = layer2_outputs[2039];
    assign layer3_outputs[2278] = ~(layer2_outputs[2515]);
    assign layer3_outputs[2279] = ~(layer2_outputs[509]);
    assign layer3_outputs[2280] = ~(layer2_outputs[2030]);
    assign layer3_outputs[2281] = ~(layer2_outputs[2514]);
    assign layer3_outputs[2282] = (layer2_outputs[1412]) & ~(layer2_outputs[1036]);
    assign layer3_outputs[2283] = (layer2_outputs[503]) & (layer2_outputs[1553]);
    assign layer3_outputs[2284] = (layer2_outputs[2142]) | (layer2_outputs[1483]);
    assign layer3_outputs[2285] = ~(layer2_outputs[1358]);
    assign layer3_outputs[2286] = ~((layer2_outputs[2279]) & (layer2_outputs[58]));
    assign layer3_outputs[2287] = (layer2_outputs[615]) & ~(layer2_outputs[2511]);
    assign layer3_outputs[2288] = layer2_outputs[1463];
    assign layer3_outputs[2289] = ~((layer2_outputs[175]) ^ (layer2_outputs[84]));
    assign layer3_outputs[2290] = layer2_outputs[1917];
    assign layer3_outputs[2291] = ~(layer2_outputs[1711]);
    assign layer3_outputs[2292] = layer2_outputs[2305];
    assign layer3_outputs[2293] = ~(layer2_outputs[993]);
    assign layer3_outputs[2294] = ~(layer2_outputs[1776]) | (layer2_outputs[1512]);
    assign layer3_outputs[2295] = layer2_outputs[1047];
    assign layer3_outputs[2296] = ~((layer2_outputs[793]) | (layer2_outputs[42]));
    assign layer3_outputs[2297] = ~((layer2_outputs[70]) | (layer2_outputs[334]));
    assign layer3_outputs[2298] = layer2_outputs[892];
    assign layer3_outputs[2299] = ~(layer2_outputs[2538]);
    assign layer3_outputs[2300] = ~((layer2_outputs[1487]) | (layer2_outputs[2534]));
    assign layer3_outputs[2301] = ~((layer2_outputs[2523]) & (layer2_outputs[318]));
    assign layer3_outputs[2302] = layer2_outputs[2364];
    assign layer3_outputs[2303] = layer2_outputs[527];
    assign layer3_outputs[2304] = ~(layer2_outputs[676]);
    assign layer3_outputs[2305] = ~(layer2_outputs[529]) | (layer2_outputs[1191]);
    assign layer3_outputs[2306] = ~(layer2_outputs[2427]);
    assign layer3_outputs[2307] = layer2_outputs[1867];
    assign layer3_outputs[2308] = ~(layer2_outputs[1429]);
    assign layer3_outputs[2309] = (layer2_outputs[2316]) | (layer2_outputs[1057]);
    assign layer3_outputs[2310] = layer2_outputs[191];
    assign layer3_outputs[2311] = ~(layer2_outputs[160]) | (layer2_outputs[1650]);
    assign layer3_outputs[2312] = ~(layer2_outputs[1917]);
    assign layer3_outputs[2313] = (layer2_outputs[2001]) & ~(layer2_outputs[2155]);
    assign layer3_outputs[2314] = (layer2_outputs[1554]) & ~(layer2_outputs[1083]);
    assign layer3_outputs[2315] = ~(layer2_outputs[1529]);
    assign layer3_outputs[2316] = layer2_outputs[33];
    assign layer3_outputs[2317] = ~((layer2_outputs[1935]) ^ (layer2_outputs[510]));
    assign layer3_outputs[2318] = (layer2_outputs[1228]) | (layer2_outputs[891]);
    assign layer3_outputs[2319] = (layer2_outputs[276]) ^ (layer2_outputs[1460]);
    assign layer3_outputs[2320] = layer2_outputs[226];
    assign layer3_outputs[2321] = layer2_outputs[2078];
    assign layer3_outputs[2322] = ~(layer2_outputs[1627]) | (layer2_outputs[69]);
    assign layer3_outputs[2323] = ~(layer2_outputs[2446]);
    assign layer3_outputs[2324] = ~(layer2_outputs[2003]) | (layer2_outputs[586]);
    assign layer3_outputs[2325] = ~(layer2_outputs[977]) | (layer2_outputs[786]);
    assign layer3_outputs[2326] = ~(layer2_outputs[1505]);
    assign layer3_outputs[2327] = ~(layer2_outputs[909]);
    assign layer3_outputs[2328] = layer2_outputs[1774];
    assign layer3_outputs[2329] = ~((layer2_outputs[53]) & (layer2_outputs[1329]));
    assign layer3_outputs[2330] = ~(layer2_outputs[355]);
    assign layer3_outputs[2331] = 1'b0;
    assign layer3_outputs[2332] = 1'b0;
    assign layer3_outputs[2333] = ~(layer2_outputs[952]);
    assign layer3_outputs[2334] = ~(layer2_outputs[1518]);
    assign layer3_outputs[2335] = layer2_outputs[809];
    assign layer3_outputs[2336] = ~(layer2_outputs[293]);
    assign layer3_outputs[2337] = ~(layer2_outputs[759]);
    assign layer3_outputs[2338] = (layer2_outputs[647]) | (layer2_outputs[1113]);
    assign layer3_outputs[2339] = ~(layer2_outputs[450]);
    assign layer3_outputs[2340] = (layer2_outputs[29]) & ~(layer2_outputs[2023]);
    assign layer3_outputs[2341] = 1'b0;
    assign layer3_outputs[2342] = ~(layer2_outputs[482]) | (layer2_outputs[1960]);
    assign layer3_outputs[2343] = ~(layer2_outputs[2300]);
    assign layer3_outputs[2344] = (layer2_outputs[62]) | (layer2_outputs[2335]);
    assign layer3_outputs[2345] = ~((layer2_outputs[312]) & (layer2_outputs[2431]));
    assign layer3_outputs[2346] = layer2_outputs[1116];
    assign layer3_outputs[2347] = 1'b0;
    assign layer3_outputs[2348] = ~((layer2_outputs[2146]) ^ (layer2_outputs[2125]));
    assign layer3_outputs[2349] = layer2_outputs[186];
    assign layer3_outputs[2350] = ~(layer2_outputs[1369]);
    assign layer3_outputs[2351] = ~((layer2_outputs[987]) & (layer2_outputs[674]));
    assign layer3_outputs[2352] = 1'b1;
    assign layer3_outputs[2353] = layer2_outputs[1616];
    assign layer3_outputs[2354] = ~(layer2_outputs[404]);
    assign layer3_outputs[2355] = ~((layer2_outputs[1408]) | (layer2_outputs[1801]));
    assign layer3_outputs[2356] = ~(layer2_outputs[967]);
    assign layer3_outputs[2357] = ~(layer2_outputs[75]);
    assign layer3_outputs[2358] = ~(layer2_outputs[2487]) | (layer2_outputs[2213]);
    assign layer3_outputs[2359] = (layer2_outputs[2301]) & ~(layer2_outputs[551]);
    assign layer3_outputs[2360] = (layer2_outputs[525]) | (layer2_outputs[781]);
    assign layer3_outputs[2361] = 1'b1;
    assign layer3_outputs[2362] = ~(layer2_outputs[728]);
    assign layer3_outputs[2363] = ~(layer2_outputs[94]);
    assign layer3_outputs[2364] = ~(layer2_outputs[946]);
    assign layer3_outputs[2365] = ~((layer2_outputs[2190]) | (layer2_outputs[1016]));
    assign layer3_outputs[2366] = ~(layer2_outputs[1554]) | (layer2_outputs[888]);
    assign layer3_outputs[2367] = ~(layer2_outputs[904]);
    assign layer3_outputs[2368] = (layer2_outputs[584]) & ~(layer2_outputs[1887]);
    assign layer3_outputs[2369] = (layer2_outputs[1171]) | (layer2_outputs[1885]);
    assign layer3_outputs[2370] = (layer2_outputs[2279]) & ~(layer2_outputs[763]);
    assign layer3_outputs[2371] = ~(layer2_outputs[2353]) | (layer2_outputs[1034]);
    assign layer3_outputs[2372] = 1'b1;
    assign layer3_outputs[2373] = layer2_outputs[422];
    assign layer3_outputs[2374] = layer2_outputs[1857];
    assign layer3_outputs[2375] = ~(layer2_outputs[965]);
    assign layer3_outputs[2376] = ~((layer2_outputs[570]) ^ (layer2_outputs[2453]));
    assign layer3_outputs[2377] = ~((layer2_outputs[2138]) & (layer2_outputs[1488]));
    assign layer3_outputs[2378] = (layer2_outputs[859]) & (layer2_outputs[1410]);
    assign layer3_outputs[2379] = 1'b1;
    assign layer3_outputs[2380] = ~(layer2_outputs[111]);
    assign layer3_outputs[2381] = ~((layer2_outputs[1634]) ^ (layer2_outputs[546]));
    assign layer3_outputs[2382] = layer2_outputs[679];
    assign layer3_outputs[2383] = ~((layer2_outputs[1959]) ^ (layer2_outputs[1539]));
    assign layer3_outputs[2384] = 1'b1;
    assign layer3_outputs[2385] = ~((layer2_outputs[326]) | (layer2_outputs[393]));
    assign layer3_outputs[2386] = ~(layer2_outputs[1515]) | (layer2_outputs[166]);
    assign layer3_outputs[2387] = ~((layer2_outputs[1616]) ^ (layer2_outputs[433]));
    assign layer3_outputs[2388] = 1'b0;
    assign layer3_outputs[2389] = ~((layer2_outputs[2206]) & (layer2_outputs[576]));
    assign layer3_outputs[2390] = ~(layer2_outputs[395]);
    assign layer3_outputs[2391] = ~((layer2_outputs[2469]) & (layer2_outputs[1660]));
    assign layer3_outputs[2392] = ~((layer2_outputs[1748]) & (layer2_outputs[1780]));
    assign layer3_outputs[2393] = (layer2_outputs[2319]) & (layer2_outputs[1421]);
    assign layer3_outputs[2394] = ~(layer2_outputs[1904]);
    assign layer3_outputs[2395] = ~((layer2_outputs[249]) & (layer2_outputs[684]));
    assign layer3_outputs[2396] = ~((layer2_outputs[795]) & (layer2_outputs[1078]));
    assign layer3_outputs[2397] = ~(layer2_outputs[1783]);
    assign layer3_outputs[2398] = (layer2_outputs[401]) & (layer2_outputs[2425]);
    assign layer3_outputs[2399] = ~(layer2_outputs[1313]) | (layer2_outputs[2204]);
    assign layer3_outputs[2400] = layer2_outputs[196];
    assign layer3_outputs[2401] = (layer2_outputs[2550]) ^ (layer2_outputs[1239]);
    assign layer3_outputs[2402] = 1'b0;
    assign layer3_outputs[2403] = ~(layer2_outputs[1465]);
    assign layer3_outputs[2404] = (layer2_outputs[1127]) ^ (layer2_outputs[1281]);
    assign layer3_outputs[2405] = ~(layer2_outputs[1982]);
    assign layer3_outputs[2406] = layer2_outputs[1066];
    assign layer3_outputs[2407] = layer2_outputs[1723];
    assign layer3_outputs[2408] = ~(layer2_outputs[1343]);
    assign layer3_outputs[2409] = 1'b0;
    assign layer3_outputs[2410] = layer2_outputs[780];
    assign layer3_outputs[2411] = ~(layer2_outputs[459]) | (layer2_outputs[2063]);
    assign layer3_outputs[2412] = (layer2_outputs[666]) & ~(layer2_outputs[118]);
    assign layer3_outputs[2413] = ~(layer2_outputs[1932]);
    assign layer3_outputs[2414] = ~(layer2_outputs[1092]);
    assign layer3_outputs[2415] = ~(layer2_outputs[922]);
    assign layer3_outputs[2416] = ~(layer2_outputs[1283]);
    assign layer3_outputs[2417] = ~(layer2_outputs[681]);
    assign layer3_outputs[2418] = (layer2_outputs[1442]) & ~(layer2_outputs[2121]);
    assign layer3_outputs[2419] = ~(layer2_outputs[580]) | (layer2_outputs[1268]);
    assign layer3_outputs[2420] = layer2_outputs[417];
    assign layer3_outputs[2421] = layer2_outputs[1054];
    assign layer3_outputs[2422] = ~(layer2_outputs[283]);
    assign layer3_outputs[2423] = (layer2_outputs[1803]) ^ (layer2_outputs[779]);
    assign layer3_outputs[2424] = layer2_outputs[621];
    assign layer3_outputs[2425] = ~((layer2_outputs[33]) & (layer2_outputs[1681]));
    assign layer3_outputs[2426] = ~(layer2_outputs[1738]);
    assign layer3_outputs[2427] = ~(layer2_outputs[931]);
    assign layer3_outputs[2428] = ~(layer2_outputs[801]);
    assign layer3_outputs[2429] = (layer2_outputs[279]) & ~(layer2_outputs[551]);
    assign layer3_outputs[2430] = ~(layer2_outputs[2032]);
    assign layer3_outputs[2431] = ~((layer2_outputs[1073]) | (layer2_outputs[103]));
    assign layer3_outputs[2432] = ~(layer2_outputs[1802]) | (layer2_outputs[2399]);
    assign layer3_outputs[2433] = (layer2_outputs[218]) & (layer2_outputs[2348]);
    assign layer3_outputs[2434] = ~(layer2_outputs[1808]) | (layer2_outputs[202]);
    assign layer3_outputs[2435] = (layer2_outputs[25]) & ~(layer2_outputs[933]);
    assign layer3_outputs[2436] = layer2_outputs[814];
    assign layer3_outputs[2437] = (layer2_outputs[2245]) & (layer2_outputs[2183]);
    assign layer3_outputs[2438] = ~(layer2_outputs[463]);
    assign layer3_outputs[2439] = ~(layer2_outputs[1589]);
    assign layer3_outputs[2440] = ~(layer2_outputs[1306]);
    assign layer3_outputs[2441] = ~((layer2_outputs[2180]) | (layer2_outputs[749]));
    assign layer3_outputs[2442] = layer2_outputs[858];
    assign layer3_outputs[2443] = layer2_outputs[35];
    assign layer3_outputs[2444] = (layer2_outputs[946]) | (layer2_outputs[126]);
    assign layer3_outputs[2445] = (layer2_outputs[1992]) ^ (layer2_outputs[1238]);
    assign layer3_outputs[2446] = ~(layer2_outputs[2071]);
    assign layer3_outputs[2447] = ~(layer2_outputs[2428]);
    assign layer3_outputs[2448] = ~(layer2_outputs[2167]);
    assign layer3_outputs[2449] = ~(layer2_outputs[2192]);
    assign layer3_outputs[2450] = 1'b0;
    assign layer3_outputs[2451] = ~(layer2_outputs[1666]) | (layer2_outputs[654]);
    assign layer3_outputs[2452] = ~((layer2_outputs[2273]) | (layer2_outputs[1583]));
    assign layer3_outputs[2453] = (layer2_outputs[1701]) & ~(layer2_outputs[2107]);
    assign layer3_outputs[2454] = ~(layer2_outputs[1570]);
    assign layer3_outputs[2455] = 1'b0;
    assign layer3_outputs[2456] = ~(layer2_outputs[2014]);
    assign layer3_outputs[2457] = (layer2_outputs[1438]) & ~(layer2_outputs[550]);
    assign layer3_outputs[2458] = (layer2_outputs[1807]) & (layer2_outputs[954]);
    assign layer3_outputs[2459] = (layer2_outputs[462]) & ~(layer2_outputs[2506]);
    assign layer3_outputs[2460] = ~(layer2_outputs[691]) | (layer2_outputs[1865]);
    assign layer3_outputs[2461] = layer2_outputs[1657];
    assign layer3_outputs[2462] = ~((layer2_outputs[1092]) ^ (layer2_outputs[1794]));
    assign layer3_outputs[2463] = layer2_outputs[2340];
    assign layer3_outputs[2464] = (layer2_outputs[2374]) ^ (layer2_outputs[1339]);
    assign layer3_outputs[2465] = ~(layer2_outputs[1879]) | (layer2_outputs[1152]);
    assign layer3_outputs[2466] = layer2_outputs[1346];
    assign layer3_outputs[2467] = ~((layer2_outputs[2093]) | (layer2_outputs[2190]));
    assign layer3_outputs[2468] = ~(layer2_outputs[1065]);
    assign layer3_outputs[2469] = (layer2_outputs[1858]) | (layer2_outputs[1460]);
    assign layer3_outputs[2470] = ~(layer2_outputs[1843]);
    assign layer3_outputs[2471] = ~(layer2_outputs[802]);
    assign layer3_outputs[2472] = ~(layer2_outputs[1304]) | (layer2_outputs[1079]);
    assign layer3_outputs[2473] = ~(layer2_outputs[1453]) | (layer2_outputs[2513]);
    assign layer3_outputs[2474] = ~(layer2_outputs[319]);
    assign layer3_outputs[2475] = (layer2_outputs[1760]) & (layer2_outputs[1093]);
    assign layer3_outputs[2476] = (layer2_outputs[574]) & ~(layer2_outputs[1567]);
    assign layer3_outputs[2477] = (layer2_outputs[846]) & ~(layer2_outputs[148]);
    assign layer3_outputs[2478] = 1'b0;
    assign layer3_outputs[2479] = ~(layer2_outputs[1787]);
    assign layer3_outputs[2480] = layer2_outputs[2015];
    assign layer3_outputs[2481] = ~(layer2_outputs[1654]);
    assign layer3_outputs[2482] = ~((layer2_outputs[1988]) | (layer2_outputs[1538]));
    assign layer3_outputs[2483] = (layer2_outputs[2173]) & ~(layer2_outputs[438]);
    assign layer3_outputs[2484] = ~(layer2_outputs[697]);
    assign layer3_outputs[2485] = (layer2_outputs[2227]) & ~(layer2_outputs[2140]);
    assign layer3_outputs[2486] = ~((layer2_outputs[1321]) ^ (layer2_outputs[1840]));
    assign layer3_outputs[2487] = ~(layer2_outputs[2020]);
    assign layer3_outputs[2488] = ~((layer2_outputs[195]) & (layer2_outputs[1405]));
    assign layer3_outputs[2489] = ~(layer2_outputs[532]);
    assign layer3_outputs[2490] = 1'b1;
    assign layer3_outputs[2491] = ~(layer2_outputs[1633]);
    assign layer3_outputs[2492] = ~(layer2_outputs[1698]);
    assign layer3_outputs[2493] = (layer2_outputs[1746]) & ~(layer2_outputs[730]);
    assign layer3_outputs[2494] = (layer2_outputs[2397]) & ~(layer2_outputs[572]);
    assign layer3_outputs[2495] = layer2_outputs[712];
    assign layer3_outputs[2496] = layer2_outputs[1781];
    assign layer3_outputs[2497] = 1'b0;
    assign layer3_outputs[2498] = ~(layer2_outputs[375]) | (layer2_outputs[526]);
    assign layer3_outputs[2499] = ~(layer2_outputs[1325]) | (layer2_outputs[659]);
    assign layer3_outputs[2500] = ~(layer2_outputs[1786]);
    assign layer3_outputs[2501] = ~((layer2_outputs[1819]) | (layer2_outputs[466]));
    assign layer3_outputs[2502] = layer2_outputs[246];
    assign layer3_outputs[2503] = ~(layer2_outputs[725]);
    assign layer3_outputs[2504] = (layer2_outputs[1499]) & (layer2_outputs[2134]);
    assign layer3_outputs[2505] = (layer2_outputs[1485]) & ~(layer2_outputs[2332]);
    assign layer3_outputs[2506] = ~(layer2_outputs[1381]);
    assign layer3_outputs[2507] = (layer2_outputs[894]) & ~(layer2_outputs[1595]);
    assign layer3_outputs[2508] = ~((layer2_outputs[1689]) ^ (layer2_outputs[564]));
    assign layer3_outputs[2509] = (layer2_outputs[746]) & ~(layer2_outputs[1812]);
    assign layer3_outputs[2510] = ~(layer2_outputs[418]);
    assign layer3_outputs[2511] = ~(layer2_outputs[2185]);
    assign layer3_outputs[2512] = ~(layer2_outputs[2028]);
    assign layer3_outputs[2513] = ~((layer2_outputs[954]) & (layer2_outputs[1523]));
    assign layer3_outputs[2514] = layer2_outputs[1301];
    assign layer3_outputs[2515] = layer2_outputs[535];
    assign layer3_outputs[2516] = layer2_outputs[5];
    assign layer3_outputs[2517] = ~(layer2_outputs[252]);
    assign layer3_outputs[2518] = layer2_outputs[1069];
    assign layer3_outputs[2519] = (layer2_outputs[2505]) & ~(layer2_outputs[420]);
    assign layer3_outputs[2520] = layer2_outputs[1225];
    assign layer3_outputs[2521] = ~(layer2_outputs[1614]);
    assign layer3_outputs[2522] = ~(layer2_outputs[2264]);
    assign layer3_outputs[2523] = layer2_outputs[2463];
    assign layer3_outputs[2524] = ~(layer2_outputs[2001]);
    assign layer3_outputs[2525] = ~(layer2_outputs[889]);
    assign layer3_outputs[2526] = ~((layer2_outputs[2555]) ^ (layer2_outputs[1335]));
    assign layer3_outputs[2527] = layer2_outputs[1937];
    assign layer3_outputs[2528] = layer2_outputs[2160];
    assign layer3_outputs[2529] = ~((layer2_outputs[2094]) & (layer2_outputs[1782]));
    assign layer3_outputs[2530] = (layer2_outputs[548]) & ~(layer2_outputs[2398]);
    assign layer3_outputs[2531] = ~(layer2_outputs[1830]);
    assign layer3_outputs[2532] = layer2_outputs[2504];
    assign layer3_outputs[2533] = 1'b0;
    assign layer3_outputs[2534] = ~((layer2_outputs[1379]) ^ (layer2_outputs[1576]));
    assign layer3_outputs[2535] = (layer2_outputs[298]) | (layer2_outputs[2247]);
    assign layer3_outputs[2536] = layer2_outputs[1587];
    assign layer3_outputs[2537] = ~((layer2_outputs[1028]) ^ (layer2_outputs[402]));
    assign layer3_outputs[2538] = ~((layer2_outputs[2261]) | (layer2_outputs[1981]));
    assign layer3_outputs[2539] = (layer2_outputs[1489]) & ~(layer2_outputs[321]);
    assign layer3_outputs[2540] = ~(layer2_outputs[994]);
    assign layer3_outputs[2541] = ~((layer2_outputs[153]) ^ (layer2_outputs[111]));
    assign layer3_outputs[2542] = layer2_outputs[1014];
    assign layer3_outputs[2543] = layer2_outputs[1599];
    assign layer3_outputs[2544] = (layer2_outputs[1291]) | (layer2_outputs[829]);
    assign layer3_outputs[2545] = ~(layer2_outputs[2455]);
    assign layer3_outputs[2546] = (layer2_outputs[2164]) | (layer2_outputs[1363]);
    assign layer3_outputs[2547] = layer2_outputs[1344];
    assign layer3_outputs[2548] = (layer2_outputs[2062]) & ~(layer2_outputs[821]);
    assign layer3_outputs[2549] = ~(layer2_outputs[117]);
    assign layer3_outputs[2550] = layer2_outputs[603];
    assign layer3_outputs[2551] = layer2_outputs[2206];
    assign layer3_outputs[2552] = ~(layer2_outputs[1740]);
    assign layer3_outputs[2553] = (layer2_outputs[441]) | (layer2_outputs[1536]);
    assign layer3_outputs[2554] = ~(layer2_outputs[392]);
    assign layer3_outputs[2555] = (layer2_outputs[1141]) & ~(layer2_outputs[1168]);
    assign layer3_outputs[2556] = ~(layer2_outputs[427]);
    assign layer3_outputs[2557] = ~(layer2_outputs[1411]) | (layer2_outputs[818]);
    assign layer3_outputs[2558] = (layer2_outputs[1854]) & ~(layer2_outputs[351]);
    assign layer3_outputs[2559] = ~(layer2_outputs[859]) | (layer2_outputs[812]);
    assign layer4_outputs[0] = layer3_outputs[130];
    assign layer4_outputs[1] = ~((layer3_outputs[313]) ^ (layer3_outputs[44]));
    assign layer4_outputs[2] = layer3_outputs[1536];
    assign layer4_outputs[3] = (layer3_outputs[1764]) ^ (layer3_outputs[1787]);
    assign layer4_outputs[4] = layer3_outputs[1076];
    assign layer4_outputs[5] = (layer3_outputs[2258]) & (layer3_outputs[2506]);
    assign layer4_outputs[6] = (layer3_outputs[2426]) & ~(layer3_outputs[1071]);
    assign layer4_outputs[7] = ~((layer3_outputs[138]) | (layer3_outputs[495]));
    assign layer4_outputs[8] = ~((layer3_outputs[2453]) & (layer3_outputs[680]));
    assign layer4_outputs[9] = (layer3_outputs[2508]) & (layer3_outputs[2240]);
    assign layer4_outputs[10] = layer3_outputs[1312];
    assign layer4_outputs[11] = ~(layer3_outputs[2035]);
    assign layer4_outputs[12] = ~((layer3_outputs[241]) ^ (layer3_outputs[2111]));
    assign layer4_outputs[13] = ~(layer3_outputs[635]);
    assign layer4_outputs[14] = layer3_outputs[72];
    assign layer4_outputs[15] = ~(layer3_outputs[2235]);
    assign layer4_outputs[16] = ~(layer3_outputs[2466]);
    assign layer4_outputs[17] = 1'b1;
    assign layer4_outputs[18] = ~(layer3_outputs[1770]);
    assign layer4_outputs[19] = ~(layer3_outputs[1396]) | (layer3_outputs[1455]);
    assign layer4_outputs[20] = ~(layer3_outputs[2173]);
    assign layer4_outputs[21] = (layer3_outputs[1144]) & (layer3_outputs[1935]);
    assign layer4_outputs[22] = (layer3_outputs[494]) & (layer3_outputs[809]);
    assign layer4_outputs[23] = ~(layer3_outputs[1181]) | (layer3_outputs[1092]);
    assign layer4_outputs[24] = ~(layer3_outputs[799]);
    assign layer4_outputs[25] = ~((layer3_outputs[143]) | (layer3_outputs[1020]));
    assign layer4_outputs[26] = ~((layer3_outputs[2458]) & (layer3_outputs[42]));
    assign layer4_outputs[27] = ~(layer3_outputs[1680]) | (layer3_outputs[1361]);
    assign layer4_outputs[28] = ~(layer3_outputs[584]) | (layer3_outputs[161]);
    assign layer4_outputs[29] = layer3_outputs[804];
    assign layer4_outputs[30] = 1'b0;
    assign layer4_outputs[31] = (layer3_outputs[357]) & (layer3_outputs[882]);
    assign layer4_outputs[32] = layer3_outputs[2337];
    assign layer4_outputs[33] = ~(layer3_outputs[664]);
    assign layer4_outputs[34] = ~((layer3_outputs[1678]) | (layer3_outputs[2083]));
    assign layer4_outputs[35] = ~(layer3_outputs[253]) | (layer3_outputs[339]);
    assign layer4_outputs[36] = ~(layer3_outputs[758]);
    assign layer4_outputs[37] = ~(layer3_outputs[417]) | (layer3_outputs[2471]);
    assign layer4_outputs[38] = 1'b1;
    assign layer4_outputs[39] = layer3_outputs[2167];
    assign layer4_outputs[40] = ~(layer3_outputs[775]);
    assign layer4_outputs[41] = ~((layer3_outputs[2167]) & (layer3_outputs[1270]));
    assign layer4_outputs[42] = 1'b1;
    assign layer4_outputs[43] = ~(layer3_outputs[46]);
    assign layer4_outputs[44] = ~(layer3_outputs[153]);
    assign layer4_outputs[45] = ~(layer3_outputs[945]) | (layer3_outputs[2327]);
    assign layer4_outputs[46] = (layer3_outputs[1752]) & ~(layer3_outputs[724]);
    assign layer4_outputs[47] = ~(layer3_outputs[307]);
    assign layer4_outputs[48] = ~((layer3_outputs[248]) | (layer3_outputs[2431]));
    assign layer4_outputs[49] = (layer3_outputs[470]) & (layer3_outputs[900]);
    assign layer4_outputs[50] = layer3_outputs[2503];
    assign layer4_outputs[51] = ~((layer3_outputs[536]) & (layer3_outputs[952]));
    assign layer4_outputs[52] = ~(layer3_outputs[1188]);
    assign layer4_outputs[53] = ~(layer3_outputs[1939]);
    assign layer4_outputs[54] = ~((layer3_outputs[549]) ^ (layer3_outputs[1844]));
    assign layer4_outputs[55] = layer3_outputs[419];
    assign layer4_outputs[56] = 1'b0;
    assign layer4_outputs[57] = ~((layer3_outputs[1635]) ^ (layer3_outputs[382]));
    assign layer4_outputs[58] = ~(layer3_outputs[906]) | (layer3_outputs[2172]);
    assign layer4_outputs[59] = layer3_outputs[1802];
    assign layer4_outputs[60] = ~((layer3_outputs[1099]) & (layer3_outputs[1311]));
    assign layer4_outputs[61] = ~(layer3_outputs[2136]);
    assign layer4_outputs[62] = (layer3_outputs[183]) | (layer3_outputs[609]);
    assign layer4_outputs[63] = ~(layer3_outputs[217]);
    assign layer4_outputs[64] = ~(layer3_outputs[552]);
    assign layer4_outputs[65] = ~(layer3_outputs[1344]);
    assign layer4_outputs[66] = ~(layer3_outputs[2371]);
    assign layer4_outputs[67] = ~((layer3_outputs[757]) & (layer3_outputs[553]));
    assign layer4_outputs[68] = (layer3_outputs[1207]) ^ (layer3_outputs[668]);
    assign layer4_outputs[69] = ~((layer3_outputs[788]) | (layer3_outputs[2267]));
    assign layer4_outputs[70] = (layer3_outputs[220]) & ~(layer3_outputs[2456]);
    assign layer4_outputs[71] = ~(layer3_outputs[2502]);
    assign layer4_outputs[72] = ~((layer3_outputs[408]) | (layer3_outputs[2144]));
    assign layer4_outputs[73] = ~((layer3_outputs[64]) & (layer3_outputs[296]));
    assign layer4_outputs[74] = ~(layer3_outputs[2299]);
    assign layer4_outputs[75] = (layer3_outputs[737]) & ~(layer3_outputs[2531]);
    assign layer4_outputs[76] = ~(layer3_outputs[1210]);
    assign layer4_outputs[77] = (layer3_outputs[2138]) ^ (layer3_outputs[628]);
    assign layer4_outputs[78] = ~((layer3_outputs[990]) | (layer3_outputs[900]));
    assign layer4_outputs[79] = (layer3_outputs[975]) ^ (layer3_outputs[499]);
    assign layer4_outputs[80] = ~(layer3_outputs[1485]);
    assign layer4_outputs[81] = (layer3_outputs[2083]) & ~(layer3_outputs[1757]);
    assign layer4_outputs[82] = layer3_outputs[1370];
    assign layer4_outputs[83] = (layer3_outputs[788]) & ~(layer3_outputs[1287]);
    assign layer4_outputs[84] = layer3_outputs[574];
    assign layer4_outputs[85] = ~(layer3_outputs[762]) | (layer3_outputs[2467]);
    assign layer4_outputs[86] = ~(layer3_outputs[92]);
    assign layer4_outputs[87] = layer3_outputs[1791];
    assign layer4_outputs[88] = 1'b0;
    assign layer4_outputs[89] = ~((layer3_outputs[915]) ^ (layer3_outputs[380]));
    assign layer4_outputs[90] = ~((layer3_outputs[2448]) ^ (layer3_outputs[937]));
    assign layer4_outputs[91] = ~(layer3_outputs[189]);
    assign layer4_outputs[92] = ~((layer3_outputs[2073]) ^ (layer3_outputs[1912]));
    assign layer4_outputs[93] = ~(layer3_outputs[1562]);
    assign layer4_outputs[94] = ~(layer3_outputs[2055]);
    assign layer4_outputs[95] = ~(layer3_outputs[571]);
    assign layer4_outputs[96] = ~((layer3_outputs[1624]) & (layer3_outputs[2428]));
    assign layer4_outputs[97] = ~((layer3_outputs[2401]) | (layer3_outputs[732]));
    assign layer4_outputs[98] = layer3_outputs[297];
    assign layer4_outputs[99] = (layer3_outputs[246]) & (layer3_outputs[831]);
    assign layer4_outputs[100] = ~(layer3_outputs[1882]) | (layer3_outputs[83]);
    assign layer4_outputs[101] = layer3_outputs[293];
    assign layer4_outputs[102] = ~(layer3_outputs[1317]);
    assign layer4_outputs[103] = ~((layer3_outputs[2078]) ^ (layer3_outputs[28]));
    assign layer4_outputs[104] = (layer3_outputs[2344]) | (layer3_outputs[872]);
    assign layer4_outputs[105] = layer3_outputs[2370];
    assign layer4_outputs[106] = ~((layer3_outputs[2266]) & (layer3_outputs[2548]));
    assign layer4_outputs[107] = layer3_outputs[633];
    assign layer4_outputs[108] = 1'b0;
    assign layer4_outputs[109] = ~(layer3_outputs[827]) | (layer3_outputs[324]);
    assign layer4_outputs[110] = ~(layer3_outputs[1397]);
    assign layer4_outputs[111] = ~((layer3_outputs[109]) & (layer3_outputs[1328]));
    assign layer4_outputs[112] = ~((layer3_outputs[2490]) | (layer3_outputs[1566]));
    assign layer4_outputs[113] = (layer3_outputs[2259]) | (layer3_outputs[1639]);
    assign layer4_outputs[114] = ~(layer3_outputs[633]);
    assign layer4_outputs[115] = ~(layer3_outputs[1518]);
    assign layer4_outputs[116] = ~(layer3_outputs[1771]);
    assign layer4_outputs[117] = ~(layer3_outputs[2175]);
    assign layer4_outputs[118] = ~((layer3_outputs[25]) ^ (layer3_outputs[1818]));
    assign layer4_outputs[119] = (layer3_outputs[1542]) | (layer3_outputs[110]);
    assign layer4_outputs[120] = ~(layer3_outputs[700]);
    assign layer4_outputs[121] = layer3_outputs[1112];
    assign layer4_outputs[122] = layer3_outputs[222];
    assign layer4_outputs[123] = ~(layer3_outputs[1277]);
    assign layer4_outputs[124] = ~(layer3_outputs[185]);
    assign layer4_outputs[125] = ~(layer3_outputs[237]);
    assign layer4_outputs[126] = ~(layer3_outputs[623]);
    assign layer4_outputs[127] = layer3_outputs[1568];
    assign layer4_outputs[128] = ~(layer3_outputs[1182]);
    assign layer4_outputs[129] = ~(layer3_outputs[664]) | (layer3_outputs[2057]);
    assign layer4_outputs[130] = ~(layer3_outputs[2419]);
    assign layer4_outputs[131] = ~(layer3_outputs[1307]) | (layer3_outputs[2351]);
    assign layer4_outputs[132] = layer3_outputs[364];
    assign layer4_outputs[133] = layer3_outputs[1739];
    assign layer4_outputs[134] = ~(layer3_outputs[13]);
    assign layer4_outputs[135] = ~(layer3_outputs[987]);
    assign layer4_outputs[136] = ~((layer3_outputs[1924]) | (layer3_outputs[1127]));
    assign layer4_outputs[137] = ~((layer3_outputs[1959]) ^ (layer3_outputs[745]));
    assign layer4_outputs[138] = ~(layer3_outputs[1657]);
    assign layer4_outputs[139] = ~(layer3_outputs[1593]);
    assign layer4_outputs[140] = ~((layer3_outputs[1337]) ^ (layer3_outputs[1012]));
    assign layer4_outputs[141] = ~((layer3_outputs[2357]) & (layer3_outputs[585]));
    assign layer4_outputs[142] = (layer3_outputs[2336]) ^ (layer3_outputs[485]);
    assign layer4_outputs[143] = ~(layer3_outputs[422]);
    assign layer4_outputs[144] = ~((layer3_outputs[421]) & (layer3_outputs[2555]));
    assign layer4_outputs[145] = layer3_outputs[1543];
    assign layer4_outputs[146] = (layer3_outputs[1755]) & ~(layer3_outputs[910]);
    assign layer4_outputs[147] = ~(layer3_outputs[635]);
    assign layer4_outputs[148] = layer3_outputs[1105];
    assign layer4_outputs[149] = ~((layer3_outputs[1582]) ^ (layer3_outputs[445]));
    assign layer4_outputs[150] = 1'b0;
    assign layer4_outputs[151] = ~(layer3_outputs[2027]);
    assign layer4_outputs[152] = layer3_outputs[1301];
    assign layer4_outputs[153] = layer3_outputs[874];
    assign layer4_outputs[154] = (layer3_outputs[1381]) ^ (layer3_outputs[1666]);
    assign layer4_outputs[155] = layer3_outputs[2253];
    assign layer4_outputs[156] = ~(layer3_outputs[698]);
    assign layer4_outputs[157] = ~(layer3_outputs[1646]);
    assign layer4_outputs[158] = (layer3_outputs[2298]) | (layer3_outputs[1340]);
    assign layer4_outputs[159] = ~((layer3_outputs[926]) & (layer3_outputs[939]));
    assign layer4_outputs[160] = (layer3_outputs[2471]) & ~(layer3_outputs[1332]);
    assign layer4_outputs[161] = layer3_outputs[1454];
    assign layer4_outputs[162] = ~(layer3_outputs[1919]);
    assign layer4_outputs[163] = (layer3_outputs[2129]) | (layer3_outputs[535]);
    assign layer4_outputs[164] = 1'b0;
    assign layer4_outputs[165] = ~(layer3_outputs[389]);
    assign layer4_outputs[166] = ~((layer3_outputs[455]) | (layer3_outputs[1371]));
    assign layer4_outputs[167] = layer3_outputs[121];
    assign layer4_outputs[168] = (layer3_outputs[398]) | (layer3_outputs[1472]);
    assign layer4_outputs[169] = (layer3_outputs[1118]) | (layer3_outputs[285]);
    assign layer4_outputs[170] = layer3_outputs[634];
    assign layer4_outputs[171] = (layer3_outputs[1679]) & ~(layer3_outputs[1484]);
    assign layer4_outputs[172] = layer3_outputs[320];
    assign layer4_outputs[173] = layer3_outputs[2255];
    assign layer4_outputs[174] = ~(layer3_outputs[311]);
    assign layer4_outputs[175] = ~(layer3_outputs[1815]);
    assign layer4_outputs[176] = ~(layer3_outputs[2127]);
    assign layer4_outputs[177] = ~((layer3_outputs[1693]) | (layer3_outputs[2460]));
    assign layer4_outputs[178] = (layer3_outputs[2221]) & ~(layer3_outputs[895]);
    assign layer4_outputs[179] = ~(layer3_outputs[2040]) | (layer3_outputs[2380]);
    assign layer4_outputs[180] = (layer3_outputs[838]) ^ (layer3_outputs[485]);
    assign layer4_outputs[181] = 1'b1;
    assign layer4_outputs[182] = ~((layer3_outputs[740]) | (layer3_outputs[2479]));
    assign layer4_outputs[183] = ~(layer3_outputs[1799]);
    assign layer4_outputs[184] = ~((layer3_outputs[491]) & (layer3_outputs[1736]));
    assign layer4_outputs[185] = layer3_outputs[1473];
    assign layer4_outputs[186] = ~(layer3_outputs[2201]);
    assign layer4_outputs[187] = ~((layer3_outputs[1812]) ^ (layer3_outputs[724]));
    assign layer4_outputs[188] = ~(layer3_outputs[162]);
    assign layer4_outputs[189] = (layer3_outputs[1027]) ^ (layer3_outputs[625]);
    assign layer4_outputs[190] = ~(layer3_outputs[1813]);
    assign layer4_outputs[191] = layer3_outputs[866];
    assign layer4_outputs[192] = (layer3_outputs[1481]) ^ (layer3_outputs[802]);
    assign layer4_outputs[193] = ~((layer3_outputs[1930]) & (layer3_outputs[1712]));
    assign layer4_outputs[194] = ~(layer3_outputs[1203]);
    assign layer4_outputs[195] = ~(layer3_outputs[2037]);
    assign layer4_outputs[196] = ~(layer3_outputs[165]);
    assign layer4_outputs[197] = ~(layer3_outputs[851]);
    assign layer4_outputs[198] = ~(layer3_outputs[123]) | (layer3_outputs[1776]);
    assign layer4_outputs[199] = (layer3_outputs[2336]) & ~(layer3_outputs[255]);
    assign layer4_outputs[200] = layer3_outputs[2126];
    assign layer4_outputs[201] = ~((layer3_outputs[1466]) | (layer3_outputs[2409]));
    assign layer4_outputs[202] = (layer3_outputs[179]) & ~(layer3_outputs[404]);
    assign layer4_outputs[203] = ~((layer3_outputs[959]) | (layer3_outputs[1639]));
    assign layer4_outputs[204] = ~(layer3_outputs[2539]);
    assign layer4_outputs[205] = layer3_outputs[1597];
    assign layer4_outputs[206] = ~((layer3_outputs[728]) | (layer3_outputs[657]));
    assign layer4_outputs[207] = ~(layer3_outputs[1289]) | (layer3_outputs[1530]);
    assign layer4_outputs[208] = ~((layer3_outputs[1933]) | (layer3_outputs[1415]));
    assign layer4_outputs[209] = (layer3_outputs[379]) & (layer3_outputs[1918]);
    assign layer4_outputs[210] = layer3_outputs[2348];
    assign layer4_outputs[211] = (layer3_outputs[1797]) | (layer3_outputs[8]);
    assign layer4_outputs[212] = ~(layer3_outputs[886]) | (layer3_outputs[1439]);
    assign layer4_outputs[213] = ~(layer3_outputs[2086]) | (layer3_outputs[1170]);
    assign layer4_outputs[214] = (layer3_outputs[979]) & (layer3_outputs[377]);
    assign layer4_outputs[215] = ~((layer3_outputs[1934]) & (layer3_outputs[2484]));
    assign layer4_outputs[216] = ~((layer3_outputs[1860]) & (layer3_outputs[160]));
    assign layer4_outputs[217] = (layer3_outputs[2463]) ^ (layer3_outputs[202]);
    assign layer4_outputs[218] = ~(layer3_outputs[1443]) | (layer3_outputs[2346]);
    assign layer4_outputs[219] = (layer3_outputs[1065]) & ~(layer3_outputs[52]);
    assign layer4_outputs[220] = ~((layer3_outputs[670]) ^ (layer3_outputs[2154]));
    assign layer4_outputs[221] = ~(layer3_outputs[736]) | (layer3_outputs[1754]);
    assign layer4_outputs[222] = ~(layer3_outputs[1610]) | (layer3_outputs[332]);
    assign layer4_outputs[223] = layer3_outputs[1167];
    assign layer4_outputs[224] = layer3_outputs[521];
    assign layer4_outputs[225] = ~((layer3_outputs[2321]) ^ (layer3_outputs[2327]));
    assign layer4_outputs[226] = ~(layer3_outputs[68]);
    assign layer4_outputs[227] = ~(layer3_outputs[336]);
    assign layer4_outputs[228] = layer3_outputs[2020];
    assign layer4_outputs[229] = ~(layer3_outputs[345]);
    assign layer4_outputs[230] = ~(layer3_outputs[852]);
    assign layer4_outputs[231] = ~(layer3_outputs[1769]) | (layer3_outputs[996]);
    assign layer4_outputs[232] = ~(layer3_outputs[2250]) | (layer3_outputs[1271]);
    assign layer4_outputs[233] = layer3_outputs[270];
    assign layer4_outputs[234] = (layer3_outputs[1317]) & ~(layer3_outputs[816]);
    assign layer4_outputs[235] = ~(layer3_outputs[2403]);
    assign layer4_outputs[236] = ~(layer3_outputs[914]);
    assign layer4_outputs[237] = ~(layer3_outputs[412]);
    assign layer4_outputs[238] = layer3_outputs[1154];
    assign layer4_outputs[239] = (layer3_outputs[251]) & ~(layer3_outputs[2118]);
    assign layer4_outputs[240] = ~(layer3_outputs[2143]);
    assign layer4_outputs[241] = ~((layer3_outputs[388]) ^ (layer3_outputs[932]));
    assign layer4_outputs[242] = layer3_outputs[879];
    assign layer4_outputs[243] = ~(layer3_outputs[441]);
    assign layer4_outputs[244] = ~(layer3_outputs[824]);
    assign layer4_outputs[245] = ~(layer3_outputs[518]) | (layer3_outputs[1147]);
    assign layer4_outputs[246] = ~(layer3_outputs[510]);
    assign layer4_outputs[247] = (layer3_outputs[631]) & ~(layer3_outputs[1798]);
    assign layer4_outputs[248] = layer3_outputs[2338];
    assign layer4_outputs[249] = ~(layer3_outputs[41]);
    assign layer4_outputs[250] = layer3_outputs[1738];
    assign layer4_outputs[251] = ~((layer3_outputs[2047]) | (layer3_outputs[360]));
    assign layer4_outputs[252] = layer3_outputs[145];
    assign layer4_outputs[253] = (layer3_outputs[1521]) ^ (layer3_outputs[1886]);
    assign layer4_outputs[254] = ~((layer3_outputs[316]) ^ (layer3_outputs[1748]));
    assign layer4_outputs[255] = ~(layer3_outputs[958]);
    assign layer4_outputs[256] = ~(layer3_outputs[2504]);
    assign layer4_outputs[257] = 1'b1;
    assign layer4_outputs[258] = ~(layer3_outputs[1064]);
    assign layer4_outputs[259] = (layer3_outputs[951]) & ~(layer3_outputs[118]);
    assign layer4_outputs[260] = layer3_outputs[1213];
    assign layer4_outputs[261] = (layer3_outputs[822]) & ~(layer3_outputs[418]);
    assign layer4_outputs[262] = layer3_outputs[1657];
    assign layer4_outputs[263] = (layer3_outputs[2461]) ^ (layer3_outputs[920]);
    assign layer4_outputs[264] = (layer3_outputs[2055]) & (layer3_outputs[468]);
    assign layer4_outputs[265] = layer3_outputs[1063];
    assign layer4_outputs[266] = ~((layer3_outputs[1117]) & (layer3_outputs[586]));
    assign layer4_outputs[267] = ~(layer3_outputs[1322]) | (layer3_outputs[451]);
    assign layer4_outputs[268] = ~((layer3_outputs[2520]) ^ (layer3_outputs[86]));
    assign layer4_outputs[269] = (layer3_outputs[2555]) & ~(layer3_outputs[1498]);
    assign layer4_outputs[270] = ~((layer3_outputs[321]) | (layer3_outputs[1184]));
    assign layer4_outputs[271] = ~((layer3_outputs[997]) ^ (layer3_outputs[2291]));
    assign layer4_outputs[272] = (layer3_outputs[2290]) | (layer3_outputs[406]);
    assign layer4_outputs[273] = ~(layer3_outputs[22]) | (layer3_outputs[564]);
    assign layer4_outputs[274] = layer3_outputs[1735];
    assign layer4_outputs[275] = ~((layer3_outputs[1765]) | (layer3_outputs[2195]));
    assign layer4_outputs[276] = layer3_outputs[1605];
    assign layer4_outputs[277] = (layer3_outputs[1011]) ^ (layer3_outputs[537]);
    assign layer4_outputs[278] = layer3_outputs[152];
    assign layer4_outputs[279] = (layer3_outputs[1023]) | (layer3_outputs[1609]);
    assign layer4_outputs[280] = layer3_outputs[420];
    assign layer4_outputs[281] = ~(layer3_outputs[1059]);
    assign layer4_outputs[282] = layer3_outputs[744];
    assign layer4_outputs[283] = ~((layer3_outputs[2274]) ^ (layer3_outputs[985]));
    assign layer4_outputs[284] = ~(layer3_outputs[18]);
    assign layer4_outputs[285] = (layer3_outputs[905]) & ~(layer3_outputs[1669]);
    assign layer4_outputs[286] = ~((layer3_outputs[1215]) ^ (layer3_outputs[1519]));
    assign layer4_outputs[287] = layer3_outputs[1710];
    assign layer4_outputs[288] = (layer3_outputs[46]) & ~(layer3_outputs[714]);
    assign layer4_outputs[289] = (layer3_outputs[216]) & ~(layer3_outputs[581]);
    assign layer4_outputs[290] = ~(layer3_outputs[1444]) | (layer3_outputs[2473]);
    assign layer4_outputs[291] = 1'b1;
    assign layer4_outputs[292] = layer3_outputs[167];
    assign layer4_outputs[293] = (layer3_outputs[903]) & ~(layer3_outputs[678]);
    assign layer4_outputs[294] = ~(layer3_outputs[566]) | (layer3_outputs[1375]);
    assign layer4_outputs[295] = layer3_outputs[60];
    assign layer4_outputs[296] = ~(layer3_outputs[1897]) | (layer3_outputs[993]);
    assign layer4_outputs[297] = layer3_outputs[54];
    assign layer4_outputs[298] = ~(layer3_outputs[224]);
    assign layer4_outputs[299] = ~(layer3_outputs[269]) | (layer3_outputs[258]);
    assign layer4_outputs[300] = layer3_outputs[1016];
    assign layer4_outputs[301] = ~(layer3_outputs[791]);
    assign layer4_outputs[302] = ~(layer3_outputs[493]);
    assign layer4_outputs[303] = layer3_outputs[1680];
    assign layer4_outputs[304] = (layer3_outputs[1400]) ^ (layer3_outputs[1093]);
    assign layer4_outputs[305] = ~(layer3_outputs[318]) | (layer3_outputs[971]);
    assign layer4_outputs[306] = ~(layer3_outputs[607]);
    assign layer4_outputs[307] = ~((layer3_outputs[2448]) & (layer3_outputs[329]));
    assign layer4_outputs[308] = layer3_outputs[493];
    assign layer4_outputs[309] = ~(layer3_outputs[1017]);
    assign layer4_outputs[310] = (layer3_outputs[1918]) & (layer3_outputs[2505]);
    assign layer4_outputs[311] = ~(layer3_outputs[1938]);
    assign layer4_outputs[312] = (layer3_outputs[2456]) | (layer3_outputs[1494]);
    assign layer4_outputs[313] = ~(layer3_outputs[2400]);
    assign layer4_outputs[314] = ~(layer3_outputs[90]);
    assign layer4_outputs[315] = ~((layer3_outputs[943]) | (layer3_outputs[1629]));
    assign layer4_outputs[316] = 1'b1;
    assign layer4_outputs[317] = ~(layer3_outputs[2247]);
    assign layer4_outputs[318] = ~(layer3_outputs[587]);
    assign layer4_outputs[319] = ~(layer3_outputs[1966]);
    assign layer4_outputs[320] = (layer3_outputs[85]) & ~(layer3_outputs[2475]);
    assign layer4_outputs[321] = layer3_outputs[1437];
    assign layer4_outputs[322] = ~(layer3_outputs[150]) | (layer3_outputs[2110]);
    assign layer4_outputs[323] = ~((layer3_outputs[1418]) & (layer3_outputs[1158]));
    assign layer4_outputs[324] = ~(layer3_outputs[1992]);
    assign layer4_outputs[325] = ~(layer3_outputs[1281]);
    assign layer4_outputs[326] = ~(layer3_outputs[2092]);
    assign layer4_outputs[327] = layer3_outputs[1607];
    assign layer4_outputs[328] = ~(layer3_outputs[70]);
    assign layer4_outputs[329] = layer3_outputs[2335];
    assign layer4_outputs[330] = ~(layer3_outputs[1755]);
    assign layer4_outputs[331] = layer3_outputs[107];
    assign layer4_outputs[332] = 1'b0;
    assign layer4_outputs[333] = ~((layer3_outputs[1926]) | (layer3_outputs[2178]));
    assign layer4_outputs[334] = ~(layer3_outputs[110]);
    assign layer4_outputs[335] = ~(layer3_outputs[1392]);
    assign layer4_outputs[336] = ~(layer3_outputs[2463]);
    assign layer4_outputs[337] = ~(layer3_outputs[837]);
    assign layer4_outputs[338] = ~(layer3_outputs[292]) | (layer3_outputs[1382]);
    assign layer4_outputs[339] = ~(layer3_outputs[15]);
    assign layer4_outputs[340] = ~((layer3_outputs[2349]) | (layer3_outputs[2018]));
    assign layer4_outputs[341] = ~(layer3_outputs[1973]);
    assign layer4_outputs[342] = ~((layer3_outputs[500]) & (layer3_outputs[1723]));
    assign layer4_outputs[343] = ~((layer3_outputs[1462]) | (layer3_outputs[1696]));
    assign layer4_outputs[344] = ~((layer3_outputs[2346]) | (layer3_outputs[2029]));
    assign layer4_outputs[345] = ~(layer3_outputs[545]);
    assign layer4_outputs[346] = (layer3_outputs[1007]) & ~(layer3_outputs[659]);
    assign layer4_outputs[347] = ~((layer3_outputs[91]) & (layer3_outputs[1539]));
    assign layer4_outputs[348] = ~(layer3_outputs[167]);
    assign layer4_outputs[349] = layer3_outputs[2330];
    assign layer4_outputs[350] = (layer3_outputs[898]) ^ (layer3_outputs[1522]);
    assign layer4_outputs[351] = layer3_outputs[1482];
    assign layer4_outputs[352] = ~(layer3_outputs[1147]);
    assign layer4_outputs[353] = ~(layer3_outputs[907]);
    assign layer4_outputs[354] = layer3_outputs[649];
    assign layer4_outputs[355] = ~((layer3_outputs[603]) ^ (layer3_outputs[965]));
    assign layer4_outputs[356] = ~(layer3_outputs[2080]) | (layer3_outputs[2476]);
    assign layer4_outputs[357] = ~((layer3_outputs[1656]) | (layer3_outputs[10]));
    assign layer4_outputs[358] = (layer3_outputs[97]) | (layer3_outputs[1060]);
    assign layer4_outputs[359] = ~(layer3_outputs[1115]);
    assign layer4_outputs[360] = ~(layer3_outputs[1655]);
    assign layer4_outputs[361] = ~(layer3_outputs[2299]);
    assign layer4_outputs[362] = layer3_outputs[1448];
    assign layer4_outputs[363] = ~(layer3_outputs[1963]) | (layer3_outputs[934]);
    assign layer4_outputs[364] = (layer3_outputs[241]) ^ (layer3_outputs[420]);
    assign layer4_outputs[365] = (layer3_outputs[50]) | (layer3_outputs[1960]);
    assign layer4_outputs[366] = (layer3_outputs[869]) & ~(layer3_outputs[1328]);
    assign layer4_outputs[367] = 1'b1;
    assign layer4_outputs[368] = ~(layer3_outputs[1531]) | (layer3_outputs[529]);
    assign layer4_outputs[369] = ~((layer3_outputs[1604]) ^ (layer3_outputs[2450]));
    assign layer4_outputs[370] = ~(layer3_outputs[2440]);
    assign layer4_outputs[371] = ~(layer3_outputs[2326]);
    assign layer4_outputs[372] = ~(layer3_outputs[1354]);
    assign layer4_outputs[373] = ~(layer3_outputs[1548]);
    assign layer4_outputs[374] = layer3_outputs[135];
    assign layer4_outputs[375] = (layer3_outputs[322]) & ~(layer3_outputs[1824]);
    assign layer4_outputs[376] = (layer3_outputs[614]) | (layer3_outputs[1489]);
    assign layer4_outputs[377] = ~((layer3_outputs[2295]) ^ (layer3_outputs[234]));
    assign layer4_outputs[378] = ~(layer3_outputs[2187]);
    assign layer4_outputs[379] = ~(layer3_outputs[26]);
    assign layer4_outputs[380] = ~(layer3_outputs[2119]) | (layer3_outputs[428]);
    assign layer4_outputs[381] = ~(layer3_outputs[1784]);
    assign layer4_outputs[382] = ~(layer3_outputs[2498]);
    assign layer4_outputs[383] = ~((layer3_outputs[1861]) & (layer3_outputs[54]));
    assign layer4_outputs[384] = (layer3_outputs[2477]) & (layer3_outputs[235]);
    assign layer4_outputs[385] = (layer3_outputs[1488]) | (layer3_outputs[2539]);
    assign layer4_outputs[386] = ~((layer3_outputs[1957]) & (layer3_outputs[579]));
    assign layer4_outputs[387] = (layer3_outputs[1958]) ^ (layer3_outputs[172]);
    assign layer4_outputs[388] = layer3_outputs[364];
    assign layer4_outputs[389] = layer3_outputs[182];
    assign layer4_outputs[390] = (layer3_outputs[314]) & ~(layer3_outputs[402]);
    assign layer4_outputs[391] = layer3_outputs[1591];
    assign layer4_outputs[392] = ~(layer3_outputs[1276]);
    assign layer4_outputs[393] = ~(layer3_outputs[1879]) | (layer3_outputs[2097]);
    assign layer4_outputs[394] = ~(layer3_outputs[2049]);
    assign layer4_outputs[395] = (layer3_outputs[1429]) | (layer3_outputs[1476]);
    assign layer4_outputs[396] = ~(layer3_outputs[1605]);
    assign layer4_outputs[397] = (layer3_outputs[619]) & (layer3_outputs[1761]);
    assign layer4_outputs[398] = ~((layer3_outputs[339]) ^ (layer3_outputs[881]));
    assign layer4_outputs[399] = ~((layer3_outputs[168]) & (layer3_outputs[1004]));
    assign layer4_outputs[400] = ~(layer3_outputs[1461]);
    assign layer4_outputs[401] = layer3_outputs[967];
    assign layer4_outputs[402] = (layer3_outputs[568]) & ~(layer3_outputs[1162]);
    assign layer4_outputs[403] = ~(layer3_outputs[2251]);
    assign layer4_outputs[404] = ~((layer3_outputs[2072]) | (layer3_outputs[279]));
    assign layer4_outputs[405] = layer3_outputs[78];
    assign layer4_outputs[406] = ~((layer3_outputs[1369]) | (layer3_outputs[260]));
    assign layer4_outputs[407] = layer3_outputs[1454];
    assign layer4_outputs[408] = layer3_outputs[2302];
    assign layer4_outputs[409] = ~(layer3_outputs[1869]) | (layer3_outputs[1623]);
    assign layer4_outputs[410] = (layer3_outputs[178]) | (layer3_outputs[1227]);
    assign layer4_outputs[411] = (layer3_outputs[2423]) & (layer3_outputs[1036]);
    assign layer4_outputs[412] = layer3_outputs[261];
    assign layer4_outputs[413] = ~(layer3_outputs[951]);
    assign layer4_outputs[414] = (layer3_outputs[1570]) & ~(layer3_outputs[293]);
    assign layer4_outputs[415] = ~((layer3_outputs[859]) & (layer3_outputs[1619]));
    assign layer4_outputs[416] = layer3_outputs[1402];
    assign layer4_outputs[417] = ~(layer3_outputs[2311]) | (layer3_outputs[543]);
    assign layer4_outputs[418] = ~(layer3_outputs[438]);
    assign layer4_outputs[419] = 1'b0;
    assign layer4_outputs[420] = ~(layer3_outputs[2324]);
    assign layer4_outputs[421] = ~((layer3_outputs[1771]) ^ (layer3_outputs[2328]));
    assign layer4_outputs[422] = ~(layer3_outputs[2147]) | (layer3_outputs[34]);
    assign layer4_outputs[423] = ~((layer3_outputs[367]) & (layer3_outputs[1998]));
    assign layer4_outputs[424] = ~(layer3_outputs[486]);
    assign layer4_outputs[425] = layer3_outputs[1733];
    assign layer4_outputs[426] = layer3_outputs[475];
    assign layer4_outputs[427] = ~(layer3_outputs[2378]) | (layer3_outputs[961]);
    assign layer4_outputs[428] = ~(layer3_outputs[1487]);
    assign layer4_outputs[429] = layer3_outputs[43];
    assign layer4_outputs[430] = ~((layer3_outputs[471]) & (layer3_outputs[1913]));
    assign layer4_outputs[431] = ~((layer3_outputs[1132]) & (layer3_outputs[1988]));
    assign layer4_outputs[432] = ~(layer3_outputs[1082]);
    assign layer4_outputs[433] = ~(layer3_outputs[2559]);
    assign layer4_outputs[434] = layer3_outputs[1698];
    assign layer4_outputs[435] = ~(layer3_outputs[2524]);
    assign layer4_outputs[436] = ~((layer3_outputs[1009]) | (layer3_outputs[1876]));
    assign layer4_outputs[437] = (layer3_outputs[467]) ^ (layer3_outputs[1388]);
    assign layer4_outputs[438] = (layer3_outputs[2191]) & (layer3_outputs[296]);
    assign layer4_outputs[439] = ~((layer3_outputs[806]) ^ (layer3_outputs[992]));
    assign layer4_outputs[440] = ~(layer3_outputs[1157]);
    assign layer4_outputs[441] = ~(layer3_outputs[860]);
    assign layer4_outputs[442] = ~((layer3_outputs[1526]) ^ (layer3_outputs[2120]));
    assign layer4_outputs[443] = ~((layer3_outputs[2118]) & (layer3_outputs[856]));
    assign layer4_outputs[444] = layer3_outputs[2260];
    assign layer4_outputs[445] = ~(layer3_outputs[1508]);
    assign layer4_outputs[446] = (layer3_outputs[1097]) ^ (layer3_outputs[828]);
    assign layer4_outputs[447] = (layer3_outputs[1812]) ^ (layer3_outputs[166]);
    assign layer4_outputs[448] = layer3_outputs[242];
    assign layer4_outputs[449] = ~(layer3_outputs[1177]) | (layer3_outputs[1969]);
    assign layer4_outputs[450] = 1'b0;
    assign layer4_outputs[451] = (layer3_outputs[2043]) & ~(layer3_outputs[826]);
    assign layer4_outputs[452] = ~(layer3_outputs[986]);
    assign layer4_outputs[453] = (layer3_outputs[738]) ^ (layer3_outputs[1928]);
    assign layer4_outputs[454] = ~(layer3_outputs[1894]);
    assign layer4_outputs[455] = ~(layer3_outputs[2425]);
    assign layer4_outputs[456] = (layer3_outputs[1524]) ^ (layer3_outputs[131]);
    assign layer4_outputs[457] = ~(layer3_outputs[1179]);
    assign layer4_outputs[458] = (layer3_outputs[1017]) & ~(layer3_outputs[726]);
    assign layer4_outputs[459] = ~(layer3_outputs[1087]);
    assign layer4_outputs[460] = ~((layer3_outputs[960]) | (layer3_outputs[1890]));
    assign layer4_outputs[461] = layer3_outputs[832];
    assign layer4_outputs[462] = (layer3_outputs[229]) ^ (layer3_outputs[294]);
    assign layer4_outputs[463] = ~(layer3_outputs[277]) | (layer3_outputs[2166]);
    assign layer4_outputs[464] = ~(layer3_outputs[798]);
    assign layer4_outputs[465] = (layer3_outputs[628]) ^ (layer3_outputs[1543]);
    assign layer4_outputs[466] = (layer3_outputs[576]) ^ (layer3_outputs[76]);
    assign layer4_outputs[467] = ~(layer3_outputs[1851]);
    assign layer4_outputs[468] = ~(layer3_outputs[2247]) | (layer3_outputs[2521]);
    assign layer4_outputs[469] = layer3_outputs[1806];
    assign layer4_outputs[470] = layer3_outputs[659];
    assign layer4_outputs[471] = (layer3_outputs[1256]) | (layer3_outputs[512]);
    assign layer4_outputs[472] = ~(layer3_outputs[554]);
    assign layer4_outputs[473] = (layer3_outputs[344]) ^ (layer3_outputs[891]);
    assign layer4_outputs[474] = layer3_outputs[1383];
    assign layer4_outputs[475] = layer3_outputs[1363];
    assign layer4_outputs[476] = ~((layer3_outputs[1215]) ^ (layer3_outputs[321]));
    assign layer4_outputs[477] = ~(layer3_outputs[2051]) | (layer3_outputs[1760]);
    assign layer4_outputs[478] = (layer3_outputs[1808]) & (layer3_outputs[723]);
    assign layer4_outputs[479] = (layer3_outputs[1467]) & ~(layer3_outputs[2342]);
    assign layer4_outputs[480] = ~(layer3_outputs[558]);
    assign layer4_outputs[481] = ~(layer3_outputs[1126]);
    assign layer4_outputs[482] = (layer3_outputs[1581]) & (layer3_outputs[101]);
    assign layer4_outputs[483] = ~(layer3_outputs[718]);
    assign layer4_outputs[484] = ~(layer3_outputs[2482]);
    assign layer4_outputs[485] = (layer3_outputs[1191]) & ~(layer3_outputs[1730]);
    assign layer4_outputs[486] = (layer3_outputs[1261]) | (layer3_outputs[1572]);
    assign layer4_outputs[487] = ~(layer3_outputs[1129]);
    assign layer4_outputs[488] = layer3_outputs[1342];
    assign layer4_outputs[489] = ~(layer3_outputs[1333]);
    assign layer4_outputs[490] = ~(layer3_outputs[2040]);
    assign layer4_outputs[491] = ~(layer3_outputs[1852]);
    assign layer4_outputs[492] = ~(layer3_outputs[102]);
    assign layer4_outputs[493] = ~(layer3_outputs[1075]);
    assign layer4_outputs[494] = layer3_outputs[2177];
    assign layer4_outputs[495] = ~(layer3_outputs[690]) | (layer3_outputs[36]);
    assign layer4_outputs[496] = (layer3_outputs[994]) & ~(layer3_outputs[787]);
    assign layer4_outputs[497] = (layer3_outputs[247]) | (layer3_outputs[1504]);
    assign layer4_outputs[498] = layer3_outputs[383];
    assign layer4_outputs[499] = layer3_outputs[1666];
    assign layer4_outputs[500] = layer3_outputs[2281];
    assign layer4_outputs[501] = layer3_outputs[924];
    assign layer4_outputs[502] = layer3_outputs[1497];
    assign layer4_outputs[503] = ~(layer3_outputs[1384]);
    assign layer4_outputs[504] = 1'b1;
    assign layer4_outputs[505] = layer3_outputs[271];
    assign layer4_outputs[506] = ~(layer3_outputs[1540]);
    assign layer4_outputs[507] = ~((layer3_outputs[2200]) ^ (layer3_outputs[1003]));
    assign layer4_outputs[508] = ~((layer3_outputs[2367]) | (layer3_outputs[2429]));
    assign layer4_outputs[509] = ~(layer3_outputs[1358]);
    assign layer4_outputs[510] = ~(layer3_outputs[2162]);
    assign layer4_outputs[511] = layer3_outputs[254];
    assign layer4_outputs[512] = layer3_outputs[284];
    assign layer4_outputs[513] = ~(layer3_outputs[259]);
    assign layer4_outputs[514] = ~(layer3_outputs[2500]);
    assign layer4_outputs[515] = layer3_outputs[264];
    assign layer4_outputs[516] = (layer3_outputs[2198]) ^ (layer3_outputs[760]);
    assign layer4_outputs[517] = ~((layer3_outputs[547]) | (layer3_outputs[1457]));
    assign layer4_outputs[518] = layer3_outputs[725];
    assign layer4_outputs[519] = layer3_outputs[2435];
    assign layer4_outputs[520] = ~(layer3_outputs[1874]) | (layer3_outputs[1836]);
    assign layer4_outputs[521] = layer3_outputs[2410];
    assign layer4_outputs[522] = (layer3_outputs[1800]) & ~(layer3_outputs[1648]);
    assign layer4_outputs[523] = layer3_outputs[1108];
    assign layer4_outputs[524] = ~(layer3_outputs[164]);
    assign layer4_outputs[525] = (layer3_outputs[511]) | (layer3_outputs[578]);
    assign layer4_outputs[526] = 1'b0;
    assign layer4_outputs[527] = (layer3_outputs[1782]) & (layer3_outputs[751]);
    assign layer4_outputs[528] = ~(layer3_outputs[756]);
    assign layer4_outputs[529] = ~(layer3_outputs[1912]);
    assign layer4_outputs[530] = layer3_outputs[1783];
    assign layer4_outputs[531] = ~(layer3_outputs[1875]);
    assign layer4_outputs[532] = ~(layer3_outputs[1128]);
    assign layer4_outputs[533] = ~(layer3_outputs[2096]);
    assign layer4_outputs[534] = ~(layer3_outputs[615]) | (layer3_outputs[898]);
    assign layer4_outputs[535] = ~(layer3_outputs[2545]);
    assign layer4_outputs[536] = ~((layer3_outputs[47]) | (layer3_outputs[1734]));
    assign layer4_outputs[537] = (layer3_outputs[127]) & ~(layer3_outputs[1611]);
    assign layer4_outputs[538] = (layer3_outputs[676]) & ~(layer3_outputs[851]);
    assign layer4_outputs[539] = ~(layer3_outputs[2466]);
    assign layer4_outputs[540] = layer3_outputs[927];
    assign layer4_outputs[541] = layer3_outputs[1220];
    assign layer4_outputs[542] = ~(layer3_outputs[1902]);
    assign layer4_outputs[543] = layer3_outputs[1529];
    assign layer4_outputs[544] = ~((layer3_outputs[1032]) & (layer3_outputs[2074]));
    assign layer4_outputs[545] = ~((layer3_outputs[1057]) | (layer3_outputs[1552]));
    assign layer4_outputs[546] = layer3_outputs[1209];
    assign layer4_outputs[547] = ~(layer3_outputs[256]);
    assign layer4_outputs[548] = ~((layer3_outputs[589]) & (layer3_outputs[245]));
    assign layer4_outputs[549] = ~(layer3_outputs[1534]);
    assign layer4_outputs[550] = layer3_outputs[140];
    assign layer4_outputs[551] = (layer3_outputs[1411]) & (layer3_outputs[1234]);
    assign layer4_outputs[552] = ~((layer3_outputs[1982]) & (layer3_outputs[282]));
    assign layer4_outputs[553] = ~(layer3_outputs[376]) | (layer3_outputs[1319]);
    assign layer4_outputs[554] = (layer3_outputs[1814]) & ~(layer3_outputs[1036]);
    assign layer4_outputs[555] = ~((layer3_outputs[538]) | (layer3_outputs[1707]));
    assign layer4_outputs[556] = ~(layer3_outputs[2297]);
    assign layer4_outputs[557] = layer3_outputs[1971];
    assign layer4_outputs[558] = ~(layer3_outputs[716]);
    assign layer4_outputs[559] = (layer3_outputs[1221]) & ~(layer3_outputs[1356]);
    assign layer4_outputs[560] = (layer3_outputs[2374]) & ~(layer3_outputs[891]);
    assign layer4_outputs[561] = layer3_outputs[1846];
    assign layer4_outputs[562] = ~(layer3_outputs[719]);
    assign layer4_outputs[563] = (layer3_outputs[231]) | (layer3_outputs[2433]);
    assign layer4_outputs[564] = ~((layer3_outputs[416]) | (layer3_outputs[2304]));
    assign layer4_outputs[565] = ~(layer3_outputs[964]);
    assign layer4_outputs[566] = layer3_outputs[1176];
    assign layer4_outputs[567] = ~(layer3_outputs[210]);
    assign layer4_outputs[568] = ~((layer3_outputs[2219]) ^ (layer3_outputs[1983]));
    assign layer4_outputs[569] = 1'b0;
    assign layer4_outputs[570] = (layer3_outputs[129]) ^ (layer3_outputs[221]);
    assign layer4_outputs[571] = layer3_outputs[1173];
    assign layer4_outputs[572] = (layer3_outputs[2418]) | (layer3_outputs[222]);
    assign layer4_outputs[573] = ~(layer3_outputs[1594]);
    assign layer4_outputs[574] = ~((layer3_outputs[596]) | (layer3_outputs[1474]));
    assign layer4_outputs[575] = layer3_outputs[400];
    assign layer4_outputs[576] = ~(layer3_outputs[2395]);
    assign layer4_outputs[577] = ~(layer3_outputs[1426]) | (layer3_outputs[1305]);
    assign layer4_outputs[578] = layer3_outputs[2214];
    assign layer4_outputs[579] = ~(layer3_outputs[1364]) | (layer3_outputs[1186]);
    assign layer4_outputs[580] = ~(layer3_outputs[439]);
    assign layer4_outputs[581] = layer3_outputs[2314];
    assign layer4_outputs[582] = ~(layer3_outputs[204]);
    assign layer4_outputs[583] = ~(layer3_outputs[1722]) | (layer3_outputs[2179]);
    assign layer4_outputs[584] = ~(layer3_outputs[2303]);
    assign layer4_outputs[585] = ~(layer3_outputs[2443]);
    assign layer4_outputs[586] = (layer3_outputs[1872]) & ~(layer3_outputs[854]);
    assign layer4_outputs[587] = ~(layer3_outputs[667]);
    assign layer4_outputs[588] = layer3_outputs[2188];
    assign layer4_outputs[589] = (layer3_outputs[2545]) & (layer3_outputs[98]);
    assign layer4_outputs[590] = ~((layer3_outputs[1156]) | (layer3_outputs[1049]));
    assign layer4_outputs[591] = layer3_outputs[394];
    assign layer4_outputs[592] = (layer3_outputs[1726]) & (layer3_outputs[1737]);
    assign layer4_outputs[593] = ~(layer3_outputs[1432]);
    assign layer4_outputs[594] = ~(layer3_outputs[1652]);
    assign layer4_outputs[595] = ~(layer3_outputs[2398]) | (layer3_outputs[158]);
    assign layer4_outputs[596] = ~((layer3_outputs[540]) ^ (layer3_outputs[572]));
    assign layer4_outputs[597] = ~(layer3_outputs[1674]) | (layer3_outputs[2093]);
    assign layer4_outputs[598] = (layer3_outputs[1715]) | (layer3_outputs[733]);
    assign layer4_outputs[599] = layer3_outputs[705];
    assign layer4_outputs[600] = ~(layer3_outputs[2279]);
    assign layer4_outputs[601] = ~((layer3_outputs[1925]) | (layer3_outputs[1790]));
    assign layer4_outputs[602] = (layer3_outputs[1373]) & (layer3_outputs[2186]);
    assign layer4_outputs[603] = layer3_outputs[1294];
    assign layer4_outputs[604] = layer3_outputs[463];
    assign layer4_outputs[605] = ~(layer3_outputs[1354]);
    assign layer4_outputs[606] = (layer3_outputs[701]) ^ (layer3_outputs[440]);
    assign layer4_outputs[607] = (layer3_outputs[1815]) ^ (layer3_outputs[2476]);
    assign layer4_outputs[608] = layer3_outputs[2308];
    assign layer4_outputs[609] = layer3_outputs[1783];
    assign layer4_outputs[610] = (layer3_outputs[1985]) | (layer3_outputs[37]);
    assign layer4_outputs[611] = layer3_outputs[1284];
    assign layer4_outputs[612] = (layer3_outputs[2417]) & (layer3_outputs[1306]);
    assign layer4_outputs[613] = ~((layer3_outputs[441]) ^ (layer3_outputs[2089]));
    assign layer4_outputs[614] = layer3_outputs[731];
    assign layer4_outputs[615] = ~(layer3_outputs[1850]) | (layer3_outputs[2509]);
    assign layer4_outputs[616] = layer3_outputs[2076];
    assign layer4_outputs[617] = layer3_outputs[2503];
    assign layer4_outputs[618] = ~(layer3_outputs[553]);
    assign layer4_outputs[619] = ~(layer3_outputs[921]);
    assign layer4_outputs[620] = layer3_outputs[1954];
    assign layer4_outputs[621] = ~((layer3_outputs[304]) & (layer3_outputs[1050]));
    assign layer4_outputs[622] = (layer3_outputs[375]) & (layer3_outputs[251]);
    assign layer4_outputs[623] = ~((layer3_outputs[1267]) & (layer3_outputs[1637]));
    assign layer4_outputs[624] = layer3_outputs[1637];
    assign layer4_outputs[625] = layer3_outputs[504];
    assign layer4_outputs[626] = ~((layer3_outputs[2523]) & (layer3_outputs[354]));
    assign layer4_outputs[627] = ~((layer3_outputs[108]) | (layer3_outputs[1229]));
    assign layer4_outputs[628] = layer3_outputs[1146];
    assign layer4_outputs[629] = layer3_outputs[1185];
    assign layer4_outputs[630] = layer3_outputs[651];
    assign layer4_outputs[631] = ~(layer3_outputs[1119]);
    assign layer4_outputs[632] = layer3_outputs[1141];
    assign layer4_outputs[633] = layer3_outputs[1073];
    assign layer4_outputs[634] = ~((layer3_outputs[1855]) ^ (layer3_outputs[1436]));
    assign layer4_outputs[635] = layer3_outputs[365];
    assign layer4_outputs[636] = ~(layer3_outputs[1642]);
    assign layer4_outputs[637] = (layer3_outputs[1645]) ^ (layer3_outputs[1596]);
    assign layer4_outputs[638] = ~(layer3_outputs[529]);
    assign layer4_outputs[639] = ~((layer3_outputs[2030]) & (layer3_outputs[1788]));
    assign layer4_outputs[640] = layer3_outputs[2124];
    assign layer4_outputs[641] = layer3_outputs[1716];
    assign layer4_outputs[642] = ~((layer3_outputs[850]) & (layer3_outputs[934]));
    assign layer4_outputs[643] = (layer3_outputs[148]) & ~(layer3_outputs[1423]);
    assign layer4_outputs[644] = ~((layer3_outputs[2381]) ^ (layer3_outputs[2041]));
    assign layer4_outputs[645] = layer3_outputs[661];
    assign layer4_outputs[646] = (layer3_outputs[1436]) & (layer3_outputs[207]);
    assign layer4_outputs[647] = layer3_outputs[2462];
    assign layer4_outputs[648] = layer3_outputs[1667];
    assign layer4_outputs[649] = (layer3_outputs[910]) ^ (layer3_outputs[1942]);
    assign layer4_outputs[650] = ~((layer3_outputs[880]) | (layer3_outputs[2275]));
    assign layer4_outputs[651] = ~(layer3_outputs[2005]) | (layer3_outputs[717]);
    assign layer4_outputs[652] = (layer3_outputs[796]) ^ (layer3_outputs[243]);
    assign layer4_outputs[653] = layer3_outputs[2103];
    assign layer4_outputs[654] = (layer3_outputs[1422]) & ~(layer3_outputs[1786]);
    assign layer4_outputs[655] = (layer3_outputs[1810]) & ~(layer3_outputs[1501]);
    assign layer4_outputs[656] = ~((layer3_outputs[2415]) & (layer3_outputs[1352]));
    assign layer4_outputs[657] = (layer3_outputs[1880]) & ~(layer3_outputs[2094]);
    assign layer4_outputs[658] = 1'b1;
    assign layer4_outputs[659] = (layer3_outputs[183]) ^ (layer3_outputs[719]);
    assign layer4_outputs[660] = ~((layer3_outputs[2245]) | (layer3_outputs[1908]));
    assign layer4_outputs[661] = ~(layer3_outputs[1352]);
    assign layer4_outputs[662] = ~(layer3_outputs[1349]);
    assign layer4_outputs[663] = ~(layer3_outputs[1506]);
    assign layer4_outputs[664] = layer3_outputs[941];
    assign layer4_outputs[665] = ~((layer3_outputs[2082]) | (layer3_outputs[3]));
    assign layer4_outputs[666] = ~((layer3_outputs[1069]) | (layer3_outputs[2512]));
    assign layer4_outputs[667] = (layer3_outputs[957]) ^ (layer3_outputs[1072]);
    assign layer4_outputs[668] = ~(layer3_outputs[863]) | (layer3_outputs[2318]);
    assign layer4_outputs[669] = layer3_outputs[905];
    assign layer4_outputs[670] = ~(layer3_outputs[2416]);
    assign layer4_outputs[671] = (layer3_outputs[2217]) & ~(layer3_outputs[1532]);
    assign layer4_outputs[672] = ~(layer3_outputs[16]);
    assign layer4_outputs[673] = 1'b0;
    assign layer4_outputs[674] = ~(layer3_outputs[1726]);
    assign layer4_outputs[675] = layer3_outputs[507];
    assign layer4_outputs[676] = ~(layer3_outputs[2549]);
    assign layer4_outputs[677] = (layer3_outputs[2226]) & (layer3_outputs[249]);
    assign layer4_outputs[678] = ~(layer3_outputs[981]);
    assign layer4_outputs[679] = ~(layer3_outputs[954]) | (layer3_outputs[1507]);
    assign layer4_outputs[680] = ~(layer3_outputs[2477]);
    assign layer4_outputs[681] = (layer3_outputs[593]) & ~(layer3_outputs[2205]);
    assign layer4_outputs[682] = (layer3_outputs[2514]) & (layer3_outputs[2292]);
    assign layer4_outputs[683] = (layer3_outputs[2035]) ^ (layer3_outputs[2491]);
    assign layer4_outputs[684] = layer3_outputs[370];
    assign layer4_outputs[685] = ~((layer3_outputs[882]) | (layer3_outputs[885]));
    assign layer4_outputs[686] = ~(layer3_outputs[1609]) | (layer3_outputs[58]);
    assign layer4_outputs[687] = layer3_outputs[2276];
    assign layer4_outputs[688] = ~(layer3_outputs[1923]);
    assign layer4_outputs[689] = layer3_outputs[806];
    assign layer4_outputs[690] = (layer3_outputs[772]) & (layer3_outputs[51]);
    assign layer4_outputs[691] = (layer3_outputs[1991]) & ~(layer3_outputs[332]);
    assign layer4_outputs[692] = (layer3_outputs[1676]) ^ (layer3_outputs[2161]);
    assign layer4_outputs[693] = ~(layer3_outputs[938]);
    assign layer4_outputs[694] = (layer3_outputs[1492]) & ~(layer3_outputs[1554]);
    assign layer4_outputs[695] = (layer3_outputs[1963]) | (layer3_outputs[2067]);
    assign layer4_outputs[696] = layer3_outputs[1000];
    assign layer4_outputs[697] = (layer3_outputs[75]) & ~(layer3_outputs[1488]);
    assign layer4_outputs[698] = ~(layer3_outputs[225]);
    assign layer4_outputs[699] = layer3_outputs[2488];
    assign layer4_outputs[700] = ~((layer3_outputs[1256]) ^ (layer3_outputs[1885]));
    assign layer4_outputs[701] = layer3_outputs[1441];
    assign layer4_outputs[702] = layer3_outputs[210];
    assign layer4_outputs[703] = layer3_outputs[1172];
    assign layer4_outputs[704] = layer3_outputs[1393];
    assign layer4_outputs[705] = ~(layer3_outputs[2192]);
    assign layer4_outputs[706] = layer3_outputs[43];
    assign layer4_outputs[707] = ~(layer3_outputs[930]);
    assign layer4_outputs[708] = layer3_outputs[1883];
    assign layer4_outputs[709] = layer3_outputs[1707];
    assign layer4_outputs[710] = layer3_outputs[1413];
    assign layer4_outputs[711] = (layer3_outputs[410]) & (layer3_outputs[2465]);
    assign layer4_outputs[712] = ~(layer3_outputs[2424]);
    assign layer4_outputs[713] = layer3_outputs[258];
    assign layer4_outputs[714] = layer3_outputs[756];
    assign layer4_outputs[715] = layer3_outputs[1456];
    assign layer4_outputs[716] = ~(layer3_outputs[778]);
    assign layer4_outputs[717] = layer3_outputs[1476];
    assign layer4_outputs[718] = ~((layer3_outputs[282]) ^ (layer3_outputs[1500]));
    assign layer4_outputs[719] = layer3_outputs[2069];
    assign layer4_outputs[720] = layer3_outputs[783];
    assign layer4_outputs[721] = (layer3_outputs[904]) & ~(layer3_outputs[1010]);
    assign layer4_outputs[722] = ~(layer3_outputs[1374]);
    assign layer4_outputs[723] = ~(layer3_outputs[2176]) | (layer3_outputs[2351]);
    assign layer4_outputs[724] = ~(layer3_outputs[59]);
    assign layer4_outputs[725] = ~(layer3_outputs[1040]);
    assign layer4_outputs[726] = (layer3_outputs[598]) | (layer3_outputs[281]);
    assign layer4_outputs[727] = ~((layer3_outputs[1198]) & (layer3_outputs[1925]));
    assign layer4_outputs[728] = (layer3_outputs[1667]) & (layer3_outputs[76]);
    assign layer4_outputs[729] = ~((layer3_outputs[297]) & (layer3_outputs[1636]));
    assign layer4_outputs[730] = ~(layer3_outputs[221]);
    assign layer4_outputs[731] = (layer3_outputs[1843]) & (layer3_outputs[964]);
    assign layer4_outputs[732] = ~(layer3_outputs[1415]) | (layer3_outputs[1008]);
    assign layer4_outputs[733] = ~(layer3_outputs[1616]);
    assign layer4_outputs[734] = layer3_outputs[691];
    assign layer4_outputs[735] = (layer3_outputs[1899]) & (layer3_outputs[87]);
    assign layer4_outputs[736] = layer3_outputs[1849];
    assign layer4_outputs[737] = layer3_outputs[2494];
    assign layer4_outputs[738] = ~((layer3_outputs[439]) | (layer3_outputs[1778]));
    assign layer4_outputs[739] = ~(layer3_outputs[399]);
    assign layer4_outputs[740] = ~(layer3_outputs[1464]);
    assign layer4_outputs[741] = layer3_outputs[1690];
    assign layer4_outputs[742] = ~(layer3_outputs[988]);
    assign layer4_outputs[743] = layer3_outputs[545];
    assign layer4_outputs[744] = ~((layer3_outputs[593]) | (layer3_outputs[242]));
    assign layer4_outputs[745] = ~(layer3_outputs[784]);
    assign layer4_outputs[746] = layer3_outputs[1533];
    assign layer4_outputs[747] = (layer3_outputs[2100]) & (layer3_outputs[230]);
    assign layer4_outputs[748] = ~(layer3_outputs[1954]) | (layer3_outputs[1979]);
    assign layer4_outputs[749] = ~(layer3_outputs[1900]);
    assign layer4_outputs[750] = ~(layer3_outputs[1613]);
    assign layer4_outputs[751] = ~((layer3_outputs[279]) | (layer3_outputs[1743]));
    assign layer4_outputs[752] = layer3_outputs[550];
    assign layer4_outputs[753] = ~(layer3_outputs[1893]);
    assign layer4_outputs[754] = ~(layer3_outputs[1670]);
    assign layer4_outputs[755] = layer3_outputs[2317];
    assign layer4_outputs[756] = (layer3_outputs[1274]) | (layer3_outputs[639]);
    assign layer4_outputs[757] = layer3_outputs[1509];
    assign layer4_outputs[758] = ~(layer3_outputs[1717]);
    assign layer4_outputs[759] = layer3_outputs[318];
    assign layer4_outputs[760] = ~((layer3_outputs[17]) ^ (layer3_outputs[2001]));
    assign layer4_outputs[761] = ~(layer3_outputs[367]) | (layer3_outputs[1151]);
    assign layer4_outputs[762] = ~(layer3_outputs[903]);
    assign layer4_outputs[763] = ~((layer3_outputs[1948]) | (layer3_outputs[1334]));
    assign layer4_outputs[764] = layer3_outputs[74];
    assign layer4_outputs[765] = ~(layer3_outputs[2419]) | (layer3_outputs[1641]);
    assign layer4_outputs[766] = ~((layer3_outputs[2128]) ^ (layer3_outputs[1999]));
    assign layer4_outputs[767] = (layer3_outputs[574]) & (layer3_outputs[1905]);
    assign layer4_outputs[768] = ~(layer3_outputs[558]);
    assign layer4_outputs[769] = ~(layer3_outputs[1922]) | (layer3_outputs[1163]);
    assign layer4_outputs[770] = ~(layer3_outputs[1692]);
    assign layer4_outputs[771] = ~((layer3_outputs[813]) ^ (layer3_outputs[1866]));
    assign layer4_outputs[772] = layer3_outputs[870];
    assign layer4_outputs[773] = ~((layer3_outputs[84]) ^ (layer3_outputs[2497]));
    assign layer4_outputs[774] = layer3_outputs[1383];
    assign layer4_outputs[775] = ~(layer3_outputs[681]);
    assign layer4_outputs[776] = ~(layer3_outputs[2128]);
    assign layer4_outputs[777] = layer3_outputs[2084];
    assign layer4_outputs[778] = ~(layer3_outputs[1545]) | (layer3_outputs[1132]);
    assign layer4_outputs[779] = layer3_outputs[495];
    assign layer4_outputs[780] = layer3_outputs[685];
    assign layer4_outputs[781] = ~((layer3_outputs[1620]) ^ (layer3_outputs[2017]));
    assign layer4_outputs[782] = layer3_outputs[2278];
    assign layer4_outputs[783] = ~(layer3_outputs[2]);
    assign layer4_outputs[784] = layer3_outputs[2367];
    assign layer4_outputs[785] = ~((layer3_outputs[2345]) ^ (layer3_outputs[1917]));
    assign layer4_outputs[786] = layer3_outputs[870];
    assign layer4_outputs[787] = ~(layer3_outputs[114]) | (layer3_outputs[146]);
    assign layer4_outputs[788] = (layer3_outputs[547]) ^ (layer3_outputs[281]);
    assign layer4_outputs[789] = ~(layer3_outputs[1980]) | (layer3_outputs[1308]);
    assign layer4_outputs[790] = ~(layer3_outputs[413]);
    assign layer4_outputs[791] = layer3_outputs[2386];
    assign layer4_outputs[792] = (layer3_outputs[191]) & ~(layer3_outputs[98]);
    assign layer4_outputs[793] = ~(layer3_outputs[2416]);
    assign layer4_outputs[794] = (layer3_outputs[995]) & ~(layer3_outputs[1013]);
    assign layer4_outputs[795] = ~(layer3_outputs[94]);
    assign layer4_outputs[796] = (layer3_outputs[268]) | (layer3_outputs[1381]);
    assign layer4_outputs[797] = ~((layer3_outputs[286]) & (layer3_outputs[1167]));
    assign layer4_outputs[798] = layer3_outputs[1615];
    assign layer4_outputs[799] = (layer3_outputs[754]) & ~(layer3_outputs[2026]);
    assign layer4_outputs[800] = ~(layer3_outputs[1964]);
    assign layer4_outputs[801] = (layer3_outputs[413]) & (layer3_outputs[344]);
    assign layer4_outputs[802] = ~(layer3_outputs[1555]);
    assign layer4_outputs[803] = ~(layer3_outputs[625]);
    assign layer4_outputs[804] = ~(layer3_outputs[502]) | (layer3_outputs[1258]);
    assign layer4_outputs[805] = ~((layer3_outputs[1144]) & (layer3_outputs[1176]));
    assign layer4_outputs[806] = ~(layer3_outputs[250]) | (layer3_outputs[568]);
    assign layer4_outputs[807] = ~(layer3_outputs[518]);
    assign layer4_outputs[808] = ~(layer3_outputs[1860]);
    assign layer4_outputs[809] = (layer3_outputs[1318]) & ~(layer3_outputs[1153]);
    assign layer4_outputs[810] = ~(layer3_outputs[2312]);
    assign layer4_outputs[811] = layer3_outputs[814];
    assign layer4_outputs[812] = ~(layer3_outputs[2418]);
    assign layer4_outputs[813] = ~(layer3_outputs[181]);
    assign layer4_outputs[814] = ~(layer3_outputs[2199]) | (layer3_outputs[1628]);
    assign layer4_outputs[815] = layer3_outputs[252];
    assign layer4_outputs[816] = (layer3_outputs[482]) ^ (layer3_outputs[1313]);
    assign layer4_outputs[817] = (layer3_outputs[100]) | (layer3_outputs[1749]);
    assign layer4_outputs[818] = ~(layer3_outputs[1200]);
    assign layer4_outputs[819] = ~((layer3_outputs[2461]) ^ (layer3_outputs[2301]));
    assign layer4_outputs[820] = layer3_outputs[2039];
    assign layer4_outputs[821] = layer3_outputs[1005];
    assign layer4_outputs[822] = layer3_outputs[1119];
    assign layer4_outputs[823] = (layer3_outputs[1660]) | (layer3_outputs[2253]);
    assign layer4_outputs[824] = ~((layer3_outputs[199]) ^ (layer3_outputs[1011]));
    assign layer4_outputs[825] = (layer3_outputs[1592]) & (layer3_outputs[1271]);
    assign layer4_outputs[826] = layer3_outputs[1804];
    assign layer4_outputs[827] = (layer3_outputs[1149]) & ~(layer3_outputs[2006]);
    assign layer4_outputs[828] = ~(layer3_outputs[1254]);
    assign layer4_outputs[829] = ~(layer3_outputs[309]);
    assign layer4_outputs[830] = (layer3_outputs[1165]) & (layer3_outputs[1220]);
    assign layer4_outputs[831] = 1'b0;
    assign layer4_outputs[832] = layer3_outputs[1461];
    assign layer4_outputs[833] = layer3_outputs[920];
    assign layer4_outputs[834] = ~(layer3_outputs[966]);
    assign layer4_outputs[835] = (layer3_outputs[570]) & ~(layer3_outputs[986]);
    assign layer4_outputs[836] = (layer3_outputs[637]) | (layer3_outputs[2354]);
    assign layer4_outputs[837] = ~(layer3_outputs[1131]) | (layer3_outputs[1208]);
    assign layer4_outputs[838] = (layer3_outputs[1611]) & ~(layer3_outputs[39]);
    assign layer4_outputs[839] = ~(layer3_outputs[148]);
    assign layer4_outputs[840] = layer3_outputs[1972];
    assign layer4_outputs[841] = ~(layer3_outputs[492]);
    assign layer4_outputs[842] = ~((layer3_outputs[682]) & (layer3_outputs[1717]));
    assign layer4_outputs[843] = ~(layer3_outputs[2071]);
    assign layer4_outputs[844] = (layer3_outputs[653]) & (layer3_outputs[676]);
    assign layer4_outputs[845] = ~(layer3_outputs[2059]);
    assign layer4_outputs[846] = ~(layer3_outputs[1701]);
    assign layer4_outputs[847] = ~(layer3_outputs[147]);
    assign layer4_outputs[848] = (layer3_outputs[1260]) & ~(layer3_outputs[531]);
    assign layer4_outputs[849] = ~(layer3_outputs[1949]) | (layer3_outputs[2041]);
    assign layer4_outputs[850] = 1'b0;
    assign layer4_outputs[851] = ~((layer3_outputs[515]) | (layer3_outputs[315]));
    assign layer4_outputs[852] = ~((layer3_outputs[2092]) | (layer3_outputs[1395]));
    assign layer4_outputs[853] = (layer3_outputs[1597]) & ~(layer3_outputs[1752]);
    assign layer4_outputs[854] = ~((layer3_outputs[519]) & (layer3_outputs[1366]));
    assign layer4_outputs[855] = (layer3_outputs[749]) & (layer3_outputs[507]);
    assign layer4_outputs[856] = ~(layer3_outputs[1060]);
    assign layer4_outputs[857] = layer3_outputs[1089];
    assign layer4_outputs[858] = layer3_outputs[2312];
    assign layer4_outputs[859] = layer3_outputs[1403];
    assign layer4_outputs[860] = (layer3_outputs[1357]) & ~(layer3_outputs[1725]);
    assign layer4_outputs[861] = (layer3_outputs[2241]) & (layer3_outputs[1424]);
    assign layer4_outputs[862] = (layer3_outputs[734]) & (layer3_outputs[1034]);
    assign layer4_outputs[863] = 1'b1;
    assign layer4_outputs[864] = (layer3_outputs[680]) ^ (layer3_outputs[1621]);
    assign layer4_outputs[865] = ~(layer3_outputs[468]);
    assign layer4_outputs[866] = ~(layer3_outputs[469]);
    assign layer4_outputs[867] = ~((layer3_outputs[2485]) & (layer3_outputs[2375]));
    assign layer4_outputs[868] = (layer3_outputs[2308]) ^ (layer3_outputs[1223]);
    assign layer4_outputs[869] = (layer3_outputs[1051]) | (layer3_outputs[2387]);
    assign layer4_outputs[870] = ~(layer3_outputs[1048]) | (layer3_outputs[570]);
    assign layer4_outputs[871] = layer3_outputs[1742];
    assign layer4_outputs[872] = (layer3_outputs[428]) | (layer3_outputs[834]);
    assign layer4_outputs[873] = ~((layer3_outputs[2206]) ^ (layer3_outputs[801]));
    assign layer4_outputs[874] = ~(layer3_outputs[2522]) | (layer3_outputs[48]);
    assign layer4_outputs[875] = layer3_outputs[415];
    assign layer4_outputs[876] = layer3_outputs[1031];
    assign layer4_outputs[877] = layer3_outputs[901];
    assign layer4_outputs[878] = (layer3_outputs[2478]) & ~(layer3_outputs[650]);
    assign layer4_outputs[879] = ~(layer3_outputs[1184]);
    assign layer4_outputs[880] = layer3_outputs[2249];
    assign layer4_outputs[881] = layer3_outputs[38];
    assign layer4_outputs[882] = ~(layer3_outputs[2426]);
    assign layer4_outputs[883] = ~(layer3_outputs[2139]) | (layer3_outputs[1613]);
    assign layer4_outputs[884] = 1'b1;
    assign layer4_outputs[885] = (layer3_outputs[1456]) & ~(layer3_outputs[1490]);
    assign layer4_outputs[886] = layer3_outputs[1022];
    assign layer4_outputs[887] = ~((layer3_outputs[1504]) | (layer3_outputs[901]));
    assign layer4_outputs[888] = (layer3_outputs[670]) ^ (layer3_outputs[1127]);
    assign layer4_outputs[889] = ~(layer3_outputs[1920]) | (layer3_outputs[2431]);
    assign layer4_outputs[890] = (layer3_outputs[1029]) & (layer3_outputs[2156]);
    assign layer4_outputs[891] = layer3_outputs[1361];
    assign layer4_outputs[892] = (layer3_outputs[2437]) ^ (layer3_outputs[1422]);
    assign layer4_outputs[893] = ~((layer3_outputs[1447]) | (layer3_outputs[842]));
    assign layer4_outputs[894] = ~((layer3_outputs[971]) | (layer3_outputs[1101]));
    assign layer4_outputs[895] = (layer3_outputs[2470]) & ~(layer3_outputs[1031]);
    assign layer4_outputs[896] = ~((layer3_outputs[168]) | (layer3_outputs[41]));
    assign layer4_outputs[897] = ~(layer3_outputs[1402]) | (layer3_outputs[1736]);
    assign layer4_outputs[898] = ~((layer3_outputs[169]) & (layer3_outputs[2323]));
    assign layer4_outputs[899] = (layer3_outputs[2383]) & (layer3_outputs[2507]);
    assign layer4_outputs[900] = ~(layer3_outputs[350]);
    assign layer4_outputs[901] = layer3_outputs[1146];
    assign layer4_outputs[902] = (layer3_outputs[2289]) | (layer3_outputs[2087]);
    assign layer4_outputs[903] = (layer3_outputs[1069]) ^ (layer3_outputs[1270]);
    assign layer4_outputs[904] = ~((layer3_outputs[72]) | (layer3_outputs[1073]));
    assign layer4_outputs[905] = ~(layer3_outputs[1549]);
    assign layer4_outputs[906] = layer3_outputs[879];
    assign layer4_outputs[907] = ~(layer3_outputs[1041]) | (layer3_outputs[1896]);
    assign layer4_outputs[908] = layer3_outputs[33];
    assign layer4_outputs[909] = ~(layer3_outputs[455]);
    assign layer4_outputs[910] = ~(layer3_outputs[324]) | (layer3_outputs[2201]);
    assign layer4_outputs[911] = ~((layer3_outputs[50]) | (layer3_outputs[2190]));
    assign layer4_outputs[912] = layer3_outputs[1206];
    assign layer4_outputs[913] = layer3_outputs[2364];
    assign layer4_outputs[914] = ~((layer3_outputs[2220]) ^ (layer3_outputs[1433]));
    assign layer4_outputs[915] = ~(layer3_outputs[2089]);
    assign layer4_outputs[916] = layer3_outputs[1760];
    assign layer4_outputs[917] = (layer3_outputs[35]) | (layer3_outputs[1793]);
    assign layer4_outputs[918] = ~(layer3_outputs[918]) | (layer3_outputs[2420]);
    assign layer4_outputs[919] = ~(layer3_outputs[1449]) | (layer3_outputs[2148]);
    assign layer4_outputs[920] = ~(layer3_outputs[1655]);
    assign layer4_outputs[921] = (layer3_outputs[2013]) & ~(layer3_outputs[12]);
    assign layer4_outputs[922] = (layer3_outputs[91]) & ~(layer3_outputs[153]);
    assign layer4_outputs[923] = (layer3_outputs[1038]) & (layer3_outputs[1405]);
    assign layer4_outputs[924] = ~((layer3_outputs[695]) ^ (layer3_outputs[973]));
    assign layer4_outputs[925] = (layer3_outputs[2170]) & ~(layer3_outputs[1384]);
    assign layer4_outputs[926] = layer3_outputs[440];
    assign layer4_outputs[927] = layer3_outputs[861];
    assign layer4_outputs[928] = layer3_outputs[1867];
    assign layer4_outputs[929] = ~((layer3_outputs[1523]) ^ (layer3_outputs[2280]));
    assign layer4_outputs[930] = layer3_outputs[1106];
    assign layer4_outputs[931] = (layer3_outputs[1246]) & ~(layer3_outputs[2069]);
    assign layer4_outputs[932] = ~((layer3_outputs[1692]) ^ (layer3_outputs[706]));
    assign layer4_outputs[933] = (layer3_outputs[1405]) & ~(layer3_outputs[1298]);
    assign layer4_outputs[934] = (layer3_outputs[2274]) ^ (layer3_outputs[970]);
    assign layer4_outputs[935] = layer3_outputs[883];
    assign layer4_outputs[936] = (layer3_outputs[754]) & ~(layer3_outputs[478]);
    assign layer4_outputs[937] = ~(layer3_outputs[397]);
    assign layer4_outputs[938] = 1'b1;
    assign layer4_outputs[939] = ~((layer3_outputs[1445]) ^ (layer3_outputs[2469]));
    assign layer4_outputs[940] = layer3_outputs[1721];
    assign layer4_outputs[941] = layer3_outputs[1864];
    assign layer4_outputs[942] = layer3_outputs[2114];
    assign layer4_outputs[943] = ~(layer3_outputs[2411]) | (layer3_outputs[696]);
    assign layer4_outputs[944] = (layer3_outputs[1024]) & (layer3_outputs[1161]);
    assign layer4_outputs[945] = (layer3_outputs[508]) | (layer3_outputs[1745]);
    assign layer4_outputs[946] = layer3_outputs[124];
    assign layer4_outputs[947] = ~(layer3_outputs[818]) | (layer3_outputs[963]);
    assign layer4_outputs[948] = (layer3_outputs[342]) & (layer3_outputs[1620]);
    assign layer4_outputs[949] = ~(layer3_outputs[697]);
    assign layer4_outputs[950] = ~((layer3_outputs[1398]) ^ (layer3_outputs[471]));
    assign layer4_outputs[951] = (layer3_outputs[45]) ^ (layer3_outputs[884]);
    assign layer4_outputs[952] = (layer3_outputs[949]) ^ (layer3_outputs[2481]);
    assign layer4_outputs[953] = layer3_outputs[442];
    assign layer4_outputs[954] = ~(layer3_outputs[735]);
    assign layer4_outputs[955] = ~(layer3_outputs[1057]) | (layer3_outputs[1539]);
    assign layer4_outputs[956] = 1'b0;
    assign layer4_outputs[957] = layer3_outputs[1104];
    assign layer4_outputs[958] = ~(layer3_outputs[942]);
    assign layer4_outputs[959] = ~(layer3_outputs[391]);
    assign layer4_outputs[960] = (layer3_outputs[70]) | (layer3_outputs[1082]);
    assign layer4_outputs[961] = ~((layer3_outputs[2023]) ^ (layer3_outputs[353]));
    assign layer4_outputs[962] = ~(layer3_outputs[540]);
    assign layer4_outputs[963] = ~((layer3_outputs[1894]) ^ (layer3_outputs[1749]));
    assign layer4_outputs[964] = ~(layer3_outputs[1187]);
    assign layer4_outputs[965] = ~(layer3_outputs[763]) | (layer3_outputs[2257]);
    assign layer4_outputs[966] = layer3_outputs[838];
    assign layer4_outputs[967] = ~(layer3_outputs[577]);
    assign layer4_outputs[968] = ~(layer3_outputs[443]);
    assign layer4_outputs[969] = ~(layer3_outputs[2102]) | (layer3_outputs[620]);
    assign layer4_outputs[970] = layer3_outputs[1340];
    assign layer4_outputs[971] = (layer3_outputs[2425]) ^ (layer3_outputs[2066]);
    assign layer4_outputs[972] = ~(layer3_outputs[2049]);
    assign layer4_outputs[973] = ~(layer3_outputs[1790]);
    assign layer4_outputs[974] = layer3_outputs[860];
    assign layer4_outputs[975] = (layer3_outputs[1716]) & ~(layer3_outputs[1314]);
    assign layer4_outputs[976] = layer3_outputs[2054];
    assign layer4_outputs[977] = layer3_outputs[1569];
    assign layer4_outputs[978] = ~(layer3_outputs[381]);
    assign layer4_outputs[979] = (layer3_outputs[1825]) | (layer3_outputs[2468]);
    assign layer4_outputs[980] = layer3_outputs[634];
    assign layer4_outputs[981] = layer3_outputs[1932];
    assign layer4_outputs[982] = (layer3_outputs[170]) & (layer3_outputs[2296]);
    assign layer4_outputs[983] = ~(layer3_outputs[1411]);
    assign layer4_outputs[984] = layer3_outputs[1373];
    assign layer4_outputs[985] = ~(layer3_outputs[1553]) | (layer3_outputs[2123]);
    assign layer4_outputs[986] = layer3_outputs[1191];
    assign layer4_outputs[987] = layer3_outputs[1739];
    assign layer4_outputs[988] = (layer3_outputs[1852]) ^ (layer3_outputs[1225]);
    assign layer4_outputs[989] = layer3_outputs[1647];
    assign layer4_outputs[990] = (layer3_outputs[2474]) | (layer3_outputs[1410]);
    assign layer4_outputs[991] = ~((layer3_outputs[1070]) | (layer3_outputs[1066]));
    assign layer4_outputs[992] = (layer3_outputs[2048]) & ~(layer3_outputs[311]);
    assign layer4_outputs[993] = layer3_outputs[2517];
    assign layer4_outputs[994] = ~((layer3_outputs[1479]) | (layer3_outputs[772]));
    assign layer4_outputs[995] = (layer3_outputs[1109]) | (layer3_outputs[2433]);
    assign layer4_outputs[996] = (layer3_outputs[1175]) & ~(layer3_outputs[159]);
    assign layer4_outputs[997] = layer3_outputs[450];
    assign layer4_outputs[998] = layer3_outputs[2363];
    assign layer4_outputs[999] = ~(layer3_outputs[1071]);
    assign layer4_outputs[1000] = ~(layer3_outputs[2527]) | (layer3_outputs[889]);
    assign layer4_outputs[1001] = ~(layer3_outputs[1940]) | (layer3_outputs[363]);
    assign layer4_outputs[1002] = layer3_outputs[69];
    assign layer4_outputs[1003] = (layer3_outputs[1277]) ^ (layer3_outputs[1997]);
    assign layer4_outputs[1004] = layer3_outputs[770];
    assign layer4_outputs[1005] = (layer3_outputs[808]) & ~(layer3_outputs[1824]);
    assign layer4_outputs[1006] = ~(layer3_outputs[32]) | (layer3_outputs[2214]);
    assign layer4_outputs[1007] = layer3_outputs[1901];
    assign layer4_outputs[1008] = ~(layer3_outputs[459]);
    assign layer4_outputs[1009] = layer3_outputs[287];
    assign layer4_outputs[1010] = ~(layer3_outputs[1826]);
    assign layer4_outputs[1011] = layer3_outputs[1723];
    assign layer4_outputs[1012] = ~(layer3_outputs[113]);
    assign layer4_outputs[1013] = ~(layer3_outputs[1856]) | (layer3_outputs[2054]);
    assign layer4_outputs[1014] = ~((layer3_outputs[679]) & (layer3_outputs[820]));
    assign layer4_outputs[1015] = layer3_outputs[1844];
    assign layer4_outputs[1016] = (layer3_outputs[2065]) & ~(layer3_outputs[684]);
    assign layer4_outputs[1017] = layer3_outputs[1495];
    assign layer4_outputs[1018] = ~((layer3_outputs[66]) ^ (layer3_outputs[1733]));
    assign layer4_outputs[1019] = layer3_outputs[2263];
    assign layer4_outputs[1020] = layer3_outputs[807];
    assign layer4_outputs[1021] = (layer3_outputs[983]) & (layer3_outputs[430]);
    assign layer4_outputs[1022] = ~(layer3_outputs[1985]);
    assign layer4_outputs[1023] = (layer3_outputs[1727]) & ~(layer3_outputs[748]);
    assign layer4_outputs[1024] = ~((layer3_outputs[2372]) & (layer3_outputs[520]));
    assign layer4_outputs[1025] = layer3_outputs[1699];
    assign layer4_outputs[1026] = layer3_outputs[268];
    assign layer4_outputs[1027] = (layer3_outputs[1160]) ^ (layer3_outputs[1737]);
    assign layer4_outputs[1028] = (layer3_outputs[1839]) & ~(layer3_outputs[833]);
    assign layer4_outputs[1029] = (layer3_outputs[2533]) & ~(layer3_outputs[319]);
    assign layer4_outputs[1030] = layer3_outputs[2015];
    assign layer4_outputs[1031] = 1'b0;
    assign layer4_outputs[1032] = ~(layer3_outputs[1506]) | (layer3_outputs[280]);
    assign layer4_outputs[1033] = ~(layer3_outputs[789]) | (layer3_outputs[2380]);
    assign layer4_outputs[1034] = (layer3_outputs[935]) & ~(layer3_outputs[2217]);
    assign layer4_outputs[1035] = ~((layer3_outputs[791]) | (layer3_outputs[203]));
    assign layer4_outputs[1036] = ~(layer3_outputs[58]);
    assign layer4_outputs[1037] = ~(layer3_outputs[1103]);
    assign layer4_outputs[1038] = ~(layer3_outputs[1989]);
    assign layer4_outputs[1039] = ~((layer3_outputs[2064]) ^ (layer3_outputs[1278]));
    assign layer4_outputs[1040] = ~(layer3_outputs[575]) | (layer3_outputs[924]);
    assign layer4_outputs[1041] = ~(layer3_outputs[2438]);
    assign layer4_outputs[1042] = ~(layer3_outputs[2099]);
    assign layer4_outputs[1043] = (layer3_outputs[1970]) & ~(layer3_outputs[589]);
    assign layer4_outputs[1044] = (layer3_outputs[1106]) & ~(layer3_outputs[774]);
    assign layer4_outputs[1045] = layer3_outputs[1896];
    assign layer4_outputs[1046] = ~((layer3_outputs[1218]) ^ (layer3_outputs[2094]));
    assign layer4_outputs[1047] = (layer3_outputs[1598]) & ~(layer3_outputs[1406]);
    assign layer4_outputs[1048] = ~(layer3_outputs[976]);
    assign layer4_outputs[1049] = ~(layer3_outputs[2314]);
    assign layer4_outputs[1050] = ~(layer3_outputs[740]);
    assign layer4_outputs[1051] = ~(layer3_outputs[2184]);
    assign layer4_outputs[1052] = ~(layer3_outputs[1350]);
    assign layer4_outputs[1053] = layer3_outputs[136];
    assign layer4_outputs[1054] = layer3_outputs[2180];
    assign layer4_outputs[1055] = ~((layer3_outputs[1283]) ^ (layer3_outputs[2306]));
    assign layer4_outputs[1056] = ~(layer3_outputs[2173]);
    assign layer4_outputs[1057] = layer3_outputs[1431];
    assign layer4_outputs[1058] = layer3_outputs[2042];
    assign layer4_outputs[1059] = ~(layer3_outputs[66]) | (layer3_outputs[115]);
    assign layer4_outputs[1060] = (layer3_outputs[1510]) | (layer3_outputs[1471]);
    assign layer4_outputs[1061] = layer3_outputs[1098];
    assign layer4_outputs[1062] = ~(layer3_outputs[2043]) | (layer3_outputs[2090]);
    assign layer4_outputs[1063] = ~(layer3_outputs[2552]) | (layer3_outputs[447]);
    assign layer4_outputs[1064] = (layer3_outputs[2427]) | (layer3_outputs[2518]);
    assign layer4_outputs[1065] = (layer3_outputs[2429]) ^ (layer3_outputs[1560]);
    assign layer4_outputs[1066] = (layer3_outputs[2398]) & ~(layer3_outputs[1348]);
    assign layer4_outputs[1067] = (layer3_outputs[341]) & ~(layer3_outputs[425]);
    assign layer4_outputs[1068] = ~(layer3_outputs[1001]) | (layer3_outputs[953]);
    assign layer4_outputs[1069] = (layer3_outputs[1030]) | (layer3_outputs[1517]);
    assign layer4_outputs[1070] = ~(layer3_outputs[1345]) | (layer3_outputs[1635]);
    assign layer4_outputs[1071] = (layer3_outputs[713]) & ~(layer3_outputs[1786]);
    assign layer4_outputs[1072] = layer3_outputs[2437];
    assign layer4_outputs[1073] = layer3_outputs[235];
    assign layer4_outputs[1074] = ~(layer3_outputs[1900]);
    assign layer4_outputs[1075] = layer3_outputs[350];
    assign layer4_outputs[1076] = ~(layer3_outputs[804]);
    assign layer4_outputs[1077] = ~(layer3_outputs[1845]) | (layer3_outputs[289]);
    assign layer4_outputs[1078] = ~(layer3_outputs[839]);
    assign layer4_outputs[1079] = layer3_outputs[1526];
    assign layer4_outputs[1080] = (layer3_outputs[395]) & ~(layer3_outputs[1503]);
    assign layer4_outputs[1081] = (layer3_outputs[945]) | (layer3_outputs[1641]);
    assign layer4_outputs[1082] = 1'b1;
    assign layer4_outputs[1083] = ~((layer3_outputs[193]) | (layer3_outputs[640]));
    assign layer4_outputs[1084] = (layer3_outputs[595]) | (layer3_outputs[854]);
    assign layer4_outputs[1085] = layer3_outputs[2220];
    assign layer4_outputs[1086] = ~(layer3_outputs[1263]);
    assign layer4_outputs[1087] = layer3_outputs[1377];
    assign layer4_outputs[1088] = (layer3_outputs[612]) & (layer3_outputs[917]);
    assign layer4_outputs[1089] = ~((layer3_outputs[2305]) | (layer3_outputs[90]));
    assign layer4_outputs[1090] = ~((layer3_outputs[601]) | (layer3_outputs[239]));
    assign layer4_outputs[1091] = (layer3_outputs[2276]) ^ (layer3_outputs[2003]);
    assign layer4_outputs[1092] = layer3_outputs[287];
    assign layer4_outputs[1093] = 1'b1;
    assign layer4_outputs[1094] = layer3_outputs[1216];
    assign layer4_outputs[1095] = 1'b1;
    assign layer4_outputs[1096] = (layer3_outputs[2288]) & (layer3_outputs[1135]);
    assign layer4_outputs[1097] = ~(layer3_outputs[828]);
    assign layer4_outputs[1098] = layer3_outputs[1133];
    assign layer4_outputs[1099] = ~(layer3_outputs[2036]);
    assign layer4_outputs[1100] = ~((layer3_outputs[1241]) ^ (layer3_outputs[317]));
    assign layer4_outputs[1101] = ~((layer3_outputs[1302]) & (layer3_outputs[985]));
    assign layer4_outputs[1102] = ~((layer3_outputs[257]) ^ (layer3_outputs[1780]));
    assign layer4_outputs[1103] = (layer3_outputs[1647]) ^ (layer3_outputs[79]);
    assign layer4_outputs[1104] = (layer3_outputs[474]) & (layer3_outputs[2441]);
    assign layer4_outputs[1105] = ~(layer3_outputs[1486]);
    assign layer4_outputs[1106] = (layer3_outputs[2528]) & (layer3_outputs[2558]);
    assign layer4_outputs[1107] = ~(layer3_outputs[2397]);
    assign layer4_outputs[1108] = ~((layer3_outputs[703]) & (layer3_outputs[1320]));
    assign layer4_outputs[1109] = ~(layer3_outputs[858]) | (layer3_outputs[1847]);
    assign layer4_outputs[1110] = (layer3_outputs[1738]) ^ (layer3_outputs[2031]);
    assign layer4_outputs[1111] = (layer3_outputs[57]) & ~(layer3_outputs[2487]);
    assign layer4_outputs[1112] = ~(layer3_outputs[1990]);
    assign layer4_outputs[1113] = (layer3_outputs[1083]) & (layer3_outputs[1380]);
    assign layer4_outputs[1114] = ~(layer3_outputs[2042]);
    assign layer4_outputs[1115] = (layer3_outputs[2166]) & ~(layer3_outputs[1731]);
    assign layer4_outputs[1116] = ~((layer3_outputs[1364]) & (layer3_outputs[973]));
    assign layer4_outputs[1117] = ~(layer3_outputs[2352]);
    assign layer4_outputs[1118] = (layer3_outputs[1711]) & (layer3_outputs[2119]);
    assign layer4_outputs[1119] = ~(layer3_outputs[1997]);
    assign layer4_outputs[1120] = ~(layer3_outputs[744]) | (layer3_outputs[21]);
    assign layer4_outputs[1121] = ~((layer3_outputs[1314]) & (layer3_outputs[1173]));
    assign layer4_outputs[1122] = ~(layer3_outputs[1531]);
    assign layer4_outputs[1123] = ~(layer3_outputs[830]);
    assign layer4_outputs[1124] = layer3_outputs[1025];
    assign layer4_outputs[1125] = layer3_outputs[1120];
    assign layer4_outputs[1126] = ~(layer3_outputs[1721]);
    assign layer4_outputs[1127] = ~(layer3_outputs[775]);
    assign layer4_outputs[1128] = layer3_outputs[1700];
    assign layer4_outputs[1129] = ~(layer3_outputs[1214]);
    assign layer4_outputs[1130] = layer3_outputs[944];
    assign layer4_outputs[1131] = ~((layer3_outputs[1921]) & (layer3_outputs[349]));
    assign layer4_outputs[1132] = ~(layer3_outputs[2383]) | (layer3_outputs[1888]);
    assign layer4_outputs[1133] = layer3_outputs[1484];
    assign layer4_outputs[1134] = layer3_outputs[1793];
    assign layer4_outputs[1135] = layer3_outputs[2359];
    assign layer4_outputs[1136] = (layer3_outputs[560]) | (layer3_outputs[2538]);
    assign layer4_outputs[1137] = ~(layer3_outputs[2171]);
    assign layer4_outputs[1138] = 1'b1;
    assign layer4_outputs[1139] = ~((layer3_outputs[1045]) | (layer3_outputs[884]));
    assign layer4_outputs[1140] = (layer3_outputs[2249]) & ~(layer3_outputs[929]);
    assign layer4_outputs[1141] = ~((layer3_outputs[864]) | (layer3_outputs[595]));
    assign layer4_outputs[1142] = ~(layer3_outputs[1243]);
    assign layer4_outputs[1143] = ~(layer3_outputs[2348]);
    assign layer4_outputs[1144] = (layer3_outputs[19]) ^ (layer3_outputs[23]);
    assign layer4_outputs[1145] = (layer3_outputs[1214]) & ~(layer3_outputs[2218]);
    assign layer4_outputs[1146] = ~(layer3_outputs[698]);
    assign layer4_outputs[1147] = (layer3_outputs[2081]) ^ (layer3_outputs[1054]);
    assign layer4_outputs[1148] = layer3_outputs[84];
    assign layer4_outputs[1149] = layer3_outputs[776];
    assign layer4_outputs[1150] = ~(layer3_outputs[822]) | (layer3_outputs[677]);
    assign layer4_outputs[1151] = ~(layer3_outputs[53]);
    assign layer4_outputs[1152] = ~(layer3_outputs[1266]);
    assign layer4_outputs[1153] = ~(layer3_outputs[1264]);
    assign layer4_outputs[1154] = layer3_outputs[617];
    assign layer4_outputs[1155] = ~(layer3_outputs[2289]) | (layer3_outputs[2550]);
    assign layer4_outputs[1156] = layer3_outputs[1976];
    assign layer4_outputs[1157] = (layer3_outputs[2340]) | (layer3_outputs[911]);
    assign layer4_outputs[1158] = ~(layer3_outputs[1112]);
    assign layer4_outputs[1159] = ~((layer3_outputs[2061]) ^ (layer3_outputs[166]));
    assign layer4_outputs[1160] = (layer3_outputs[379]) & ~(layer3_outputs[2271]);
    assign layer4_outputs[1161] = (layer3_outputs[640]) ^ (layer3_outputs[1809]);
    assign layer4_outputs[1162] = ~(layer3_outputs[832]) | (layer3_outputs[1168]);
    assign layer4_outputs[1163] = layer3_outputs[2388];
    assign layer4_outputs[1164] = (layer3_outputs[2374]) & (layer3_outputs[693]);
    assign layer4_outputs[1165] = ~(layer3_outputs[830]);
    assign layer4_outputs[1166] = (layer3_outputs[1831]) | (layer3_outputs[1534]);
    assign layer4_outputs[1167] = ~((layer3_outputs[1881]) ^ (layer3_outputs[214]));
    assign layer4_outputs[1168] = ~(layer3_outputs[1865]);
    assign layer4_outputs[1169] = 1'b1;
    assign layer4_outputs[1170] = ~(layer3_outputs[223]) | (layer3_outputs[283]);
    assign layer4_outputs[1171] = ~((layer3_outputs[1316]) ^ (layer3_outputs[61]));
    assign layer4_outputs[1172] = ~(layer3_outputs[498]) | (layer3_outputs[2464]);
    assign layer4_outputs[1173] = layer3_outputs[997];
    assign layer4_outputs[1174] = ~(layer3_outputs[65]);
    assign layer4_outputs[1175] = ~(layer3_outputs[65]) | (layer3_outputs[32]);
    assign layer4_outputs[1176] = ~(layer3_outputs[1205]);
    assign layer4_outputs[1177] = (layer3_outputs[338]) & ~(layer3_outputs[2378]);
    assign layer4_outputs[1178] = ~(layer3_outputs[192]);
    assign layer4_outputs[1179] = ~((layer3_outputs[2342]) ^ (layer3_outputs[496]));
    assign layer4_outputs[1180] = ~(layer3_outputs[2213]);
    assign layer4_outputs[1181] = layer3_outputs[611];
    assign layer4_outputs[1182] = (layer3_outputs[486]) & ~(layer3_outputs[2033]);
    assign layer4_outputs[1183] = layer3_outputs[1547];
    assign layer4_outputs[1184] = ~(layer3_outputs[2097]);
    assign layer4_outputs[1185] = (layer3_outputs[519]) & ~(layer3_outputs[1139]);
    assign layer4_outputs[1186] = (layer3_outputs[1110]) & ~(layer3_outputs[1841]);
    assign layer4_outputs[1187] = (layer3_outputs[1273]) & ~(layer3_outputs[2498]);
    assign layer4_outputs[1188] = ~(layer3_outputs[1742]) | (layer3_outputs[1563]);
    assign layer4_outputs[1189] = (layer3_outputs[1688]) & (layer3_outputs[1003]);
    assign layer4_outputs[1190] = ~(layer3_outputs[1781]);
    assign layer4_outputs[1191] = 1'b0;
    assign layer4_outputs[1192] = ~(layer3_outputs[972]);
    assign layer4_outputs[1193] = layer3_outputs[2447];
    assign layer4_outputs[1194] = layer3_outputs[661];
    assign layer4_outputs[1195] = ~(layer3_outputs[2265]);
    assign layer4_outputs[1196] = (layer3_outputs[1502]) & ~(layer3_outputs[1125]);
    assign layer4_outputs[1197] = layer3_outputs[1179];
    assign layer4_outputs[1198] = (layer3_outputs[1329]) & (layer3_outputs[768]);
    assign layer4_outputs[1199] = ~(layer3_outputs[1043]);
    assign layer4_outputs[1200] = ~(layer3_outputs[1190]);
    assign layer4_outputs[1201] = layer3_outputs[1282];
    assign layer4_outputs[1202] = ~(layer3_outputs[81]);
    assign layer4_outputs[1203] = (layer3_outputs[966]) & (layer3_outputs[2204]);
    assign layer4_outputs[1204] = ~(layer3_outputs[887]);
    assign layer4_outputs[1205] = layer3_outputs[2138];
    assign layer4_outputs[1206] = layer3_outputs[2369];
    assign layer4_outputs[1207] = ~(layer3_outputs[206]) | (layer3_outputs[2386]);
    assign layer4_outputs[1208] = (layer3_outputs[2488]) & ~(layer3_outputs[432]);
    assign layer4_outputs[1209] = ~(layer3_outputs[1741]);
    assign layer4_outputs[1210] = ~((layer3_outputs[1324]) ^ (layer3_outputs[1032]));
    assign layer4_outputs[1211] = ~(layer3_outputs[836]);
    assign layer4_outputs[1212] = (layer3_outputs[944]) ^ (layer3_outputs[96]);
    assign layer4_outputs[1213] = layer3_outputs[2522];
    assign layer4_outputs[1214] = layer3_outputs[233];
    assign layer4_outputs[1215] = layer3_outputs[2462];
    assign layer4_outputs[1216] = ~(layer3_outputs[1948]);
    assign layer4_outputs[1217] = (layer3_outputs[198]) | (layer3_outputs[2333]);
    assign layer4_outputs[1218] = ~(layer3_outputs[177]);
    assign layer4_outputs[1219] = ~(layer3_outputs[1358]) | (layer3_outputs[2132]);
    assign layer4_outputs[1220] = layer3_outputs[2246];
    assign layer4_outputs[1221] = (layer3_outputs[1964]) & (layer3_outputs[2406]);
    assign layer4_outputs[1222] = layer3_outputs[1413];
    assign layer4_outputs[1223] = ~(layer3_outputs[583]);
    assign layer4_outputs[1224] = ~((layer3_outputs[184]) | (layer3_outputs[2459]));
    assign layer4_outputs[1225] = ~(layer3_outputs[2239]);
    assign layer4_outputs[1226] = ~(layer3_outputs[2202]) | (layer3_outputs[1293]);
    assign layer4_outputs[1227] = layer3_outputs[337];
    assign layer4_outputs[1228] = (layer3_outputs[1193]) & ~(layer3_outputs[1386]);
    assign layer4_outputs[1229] = layer3_outputs[2307];
    assign layer4_outputs[1230] = (layer3_outputs[564]) | (layer3_outputs[1409]);
    assign layer4_outputs[1231] = (layer3_outputs[702]) & ~(layer3_outputs[1653]);
    assign layer4_outputs[1232] = layer3_outputs[1563];
    assign layer4_outputs[1233] = ~(layer3_outputs[2382]);
    assign layer4_outputs[1234] = (layer3_outputs[273]) & ~(layer3_outputs[22]);
    assign layer4_outputs[1235] = ~((layer3_outputs[1138]) | (layer3_outputs[1310]));
    assign layer4_outputs[1236] = layer3_outputs[1148];
    assign layer4_outputs[1237] = layer3_outputs[85];
    assign layer4_outputs[1238] = ~(layer3_outputs[1077]);
    assign layer4_outputs[1239] = ~(layer3_outputs[1728]);
    assign layer4_outputs[1240] = layer3_outputs[1868];
    assign layer4_outputs[1241] = ~((layer3_outputs[1514]) | (layer3_outputs[2125]));
    assign layer4_outputs[1242] = ~(layer3_outputs[1818]) | (layer3_outputs[1006]);
    assign layer4_outputs[1243] = (layer3_outputs[211]) & ~(layer3_outputs[1475]);
    assign layer4_outputs[1244] = layer3_outputs[859];
    assign layer4_outputs[1245] = layer3_outputs[1114];
    assign layer4_outputs[1246] = ~(layer3_outputs[1367]);
    assign layer4_outputs[1247] = layer3_outputs[310];
    assign layer4_outputs[1248] = layer3_outputs[270];
    assign layer4_outputs[1249] = ~(layer3_outputs[2207]);
    assign layer4_outputs[1250] = (layer3_outputs[360]) | (layer3_outputs[2127]);
    assign layer4_outputs[1251] = (layer3_outputs[1039]) | (layer3_outputs[1240]);
    assign layer4_outputs[1252] = layer3_outputs[1204];
    assign layer4_outputs[1253] = (layer3_outputs[894]) & ~(layer3_outputs[641]);
    assign layer4_outputs[1254] = (layer3_outputs[1312]) | (layer3_outputs[1428]);
    assign layer4_outputs[1255] = (layer3_outputs[2321]) ^ (layer3_outputs[675]);
    assign layer4_outputs[1256] = ~(layer3_outputs[1096]);
    assign layer4_outputs[1257] = (layer3_outputs[1107]) ^ (layer3_outputs[808]);
    assign layer4_outputs[1258] = ~((layer3_outputs[490]) & (layer3_outputs[968]));
    assign layer4_outputs[1259] = ~((layer3_outputs[785]) | (layer3_outputs[810]));
    assign layer4_outputs[1260] = layer3_outputs[1800];
    assign layer4_outputs[1261] = ~(layer3_outputs[1445]) | (layer3_outputs[1541]);
    assign layer4_outputs[1262] = (layer3_outputs[1505]) ^ (layer3_outputs[371]);
    assign layer4_outputs[1263] = layer3_outputs[626];
    assign layer4_outputs[1264] = layer3_outputs[1109];
    assign layer4_outputs[1265] = ~(layer3_outputs[1569]);
    assign layer4_outputs[1266] = layer3_outputs[1251];
    assign layer4_outputs[1267] = 1'b0;
    assign layer4_outputs[1268] = ~(layer3_outputs[2095]);
    assign layer4_outputs[1269] = layer3_outputs[352];
    assign layer4_outputs[1270] = ~(layer3_outputs[2052]);
    assign layer4_outputs[1271] = (layer3_outputs[346]) & ~(layer3_outputs[1623]);
    assign layer4_outputs[1272] = (layer3_outputs[1718]) ^ (layer3_outputs[299]);
    assign layer4_outputs[1273] = ~(layer3_outputs[513]);
    assign layer4_outputs[1274] = ~(layer3_outputs[423]);
    assign layer4_outputs[1275] = ~((layer3_outputs[656]) & (layer3_outputs[779]));
    assign layer4_outputs[1276] = layer3_outputs[780];
    assign layer4_outputs[1277] = (layer3_outputs[226]) ^ (layer3_outputs[1614]);
    assign layer4_outputs[1278] = ~((layer3_outputs[1325]) & (layer3_outputs[687]));
    assign layer4_outputs[1279] = (layer3_outputs[2331]) & ~(layer3_outputs[137]);
    assign layer4_outputs[1280] = (layer3_outputs[2459]) & (layer3_outputs[1735]);
    assign layer4_outputs[1281] = layer3_outputs[1385];
    assign layer4_outputs[1282] = layer3_outputs[2215];
    assign layer4_outputs[1283] = layer3_outputs[1424];
    assign layer4_outputs[1284] = layer3_outputs[487];
    assign layer4_outputs[1285] = (layer3_outputs[2219]) & ~(layer3_outputs[2339]);
    assign layer4_outputs[1286] = (layer3_outputs[190]) & ~(layer3_outputs[500]);
    assign layer4_outputs[1287] = layer3_outputs[1518];
    assign layer4_outputs[1288] = ~(layer3_outputs[516]);
    assign layer4_outputs[1289] = (layer3_outputs[2248]) & ~(layer3_outputs[692]);
    assign layer4_outputs[1290] = layer3_outputs[1245];
    assign layer4_outputs[1291] = ~(layer3_outputs[97]);
    assign layer4_outputs[1292] = ~(layer3_outputs[528]);
    assign layer4_outputs[1293] = ~((layer3_outputs[1795]) & (layer3_outputs[1094]));
    assign layer4_outputs[1294] = (layer3_outputs[747]) & ~(layer3_outputs[608]);
    assign layer4_outputs[1295] = layer3_outputs[1855];
    assign layer4_outputs[1296] = ~(layer3_outputs[1779]);
    assign layer4_outputs[1297] = layer3_outputs[2053];
    assign layer4_outputs[1298] = layer3_outputs[913];
    assign layer4_outputs[1299] = layer3_outputs[1128];
    assign layer4_outputs[1300] = 1'b1;
    assign layer4_outputs[1301] = layer3_outputs[611];
    assign layer4_outputs[1302] = (layer3_outputs[1395]) & ~(layer3_outputs[520]);
    assign layer4_outputs[1303] = (layer3_outputs[1907]) ^ (layer3_outputs[2088]);
    assign layer4_outputs[1304] = (layer3_outputs[2098]) & ~(layer3_outputs[365]);
    assign layer4_outputs[1305] = ~(layer3_outputs[1100]) | (layer3_outputs[989]);
    assign layer4_outputs[1306] = ~(layer3_outputs[406]);
    assign layer4_outputs[1307] = ~(layer3_outputs[1375]);
    assign layer4_outputs[1308] = layer3_outputs[2553];
    assign layer4_outputs[1309] = 1'b0;
    assign layer4_outputs[1310] = ~(layer3_outputs[29]) | (layer3_outputs[138]);
    assign layer4_outputs[1311] = layer3_outputs[1659];
    assign layer4_outputs[1312] = ~((layer3_outputs[2149]) ^ (layer3_outputs[1033]));
    assign layer4_outputs[1313] = ~(layer3_outputs[27]);
    assign layer4_outputs[1314] = layer3_outputs[652];
    assign layer4_outputs[1315] = (layer3_outputs[1775]) & (layer3_outputs[2172]);
    assign layer4_outputs[1316] = ~(layer3_outputs[1633]);
    assign layer4_outputs[1317] = ~(layer3_outputs[78]) | (layer3_outputs[1427]);
    assign layer4_outputs[1318] = (layer3_outputs[403]) & ~(layer3_outputs[1452]);
    assign layer4_outputs[1319] = (layer3_outputs[157]) ^ (layer3_outputs[1615]);
    assign layer4_outputs[1320] = (layer3_outputs[1745]) & ~(layer3_outputs[1584]);
    assign layer4_outputs[1321] = ~((layer3_outputs[1053]) & (layer3_outputs[432]));
    assign layer4_outputs[1322] = layer3_outputs[2211];
    assign layer4_outputs[1323] = layer3_outputs[2046];
    assign layer4_outputs[1324] = ~(layer3_outputs[1110]);
    assign layer4_outputs[1325] = ~(layer3_outputs[697]);
    assign layer4_outputs[1326] = ~(layer3_outputs[1614]) | (layer3_outputs[765]);
    assign layer4_outputs[1327] = layer3_outputs[2427];
    assign layer4_outputs[1328] = layer3_outputs[342];
    assign layer4_outputs[1329] = layer3_outputs[1407];
    assign layer4_outputs[1330] = ~(layer3_outputs[2079]);
    assign layer4_outputs[1331] = (layer3_outputs[1472]) ^ (layer3_outputs[26]);
    assign layer4_outputs[1332] = ~(layer3_outputs[1584]);
    assign layer4_outputs[1333] = ~(layer3_outputs[1360]);
    assign layer4_outputs[1334] = ~(layer3_outputs[106]);
    assign layer4_outputs[1335] = ~((layer3_outputs[386]) | (layer3_outputs[916]));
    assign layer4_outputs[1336] = ~(layer3_outputs[289]);
    assign layer4_outputs[1337] = (layer3_outputs[1676]) & (layer3_outputs[275]);
    assign layer4_outputs[1338] = ~(layer3_outputs[2036]) | (layer3_outputs[1018]);
    assign layer4_outputs[1339] = ~((layer3_outputs[1748]) & (layer3_outputs[2421]));
    assign layer4_outputs[1340] = (layer3_outputs[1280]) | (layer3_outputs[2082]);
    assign layer4_outputs[1341] = ~((layer3_outputs[2073]) | (layer3_outputs[588]));
    assign layer4_outputs[1342] = layer3_outputs[605];
    assign layer4_outputs[1343] = (layer3_outputs[2087]) & (layer3_outputs[1479]);
    assign layer4_outputs[1344] = (layer3_outputs[875]) & ~(layer3_outputs[2058]);
    assign layer4_outputs[1345] = ~(layer3_outputs[2387]);
    assign layer4_outputs[1346] = layer3_outputs[1943];
    assign layer4_outputs[1347] = ~(layer3_outputs[1778]) | (layer3_outputs[1588]);
    assign layer4_outputs[1348] = layer3_outputs[476];
    assign layer4_outputs[1349] = layer3_outputs[2521];
    assign layer4_outputs[1350] = ~((layer3_outputs[2528]) & (layer3_outputs[2157]));
    assign layer4_outputs[1351] = layer3_outputs[844];
    assign layer4_outputs[1352] = (layer3_outputs[2358]) ^ (layer3_outputs[690]);
    assign layer4_outputs[1353] = ~(layer3_outputs[415]);
    assign layer4_outputs[1354] = (layer3_outputs[1810]) & ~(layer3_outputs[2420]);
    assign layer4_outputs[1355] = ~((layer3_outputs[1537]) & (layer3_outputs[2228]));
    assign layer4_outputs[1356] = (layer3_outputs[1965]) ^ (layer3_outputs[1217]);
    assign layer4_outputs[1357] = ~(layer3_outputs[2294]);
    assign layer4_outputs[1358] = ~((layer3_outputs[781]) ^ (layer3_outputs[1906]));
    assign layer4_outputs[1359] = layer3_outputs[1718];
    assign layer4_outputs[1360] = ~(layer3_outputs[525]) | (layer3_outputs[2210]);
    assign layer4_outputs[1361] = ~(layer3_outputs[646]);
    assign layer4_outputs[1362] = ~(layer3_outputs[2458]);
    assign layer4_outputs[1363] = 1'b0;
    assign layer4_outputs[1364] = layer3_outputs[580];
    assign layer4_outputs[1365] = layer3_outputs[1257];
    assign layer4_outputs[1366] = ~(layer3_outputs[1898]);
    assign layer4_outputs[1367] = (layer3_outputs[336]) ^ (layer3_outputs[1792]);
    assign layer4_outputs[1368] = ~(layer3_outputs[2318]) | (layer3_outputs[865]);
    assign layer4_outputs[1369] = layer3_outputs[2184];
    assign layer4_outputs[1370] = ~(layer3_outputs[136]) | (layer3_outputs[62]);
    assign layer4_outputs[1371] = ~((layer3_outputs[1834]) | (layer3_outputs[2075]));
    assign layer4_outputs[1372] = layer3_outputs[479];
    assign layer4_outputs[1373] = 1'b0;
    assign layer4_outputs[1374] = layer3_outputs[1198];
    assign layer4_outputs[1375] = ~(layer3_outputs[526]);
    assign layer4_outputs[1376] = 1'b0;
    assign layer4_outputs[1377] = (layer3_outputs[111]) ^ (layer3_outputs[1244]);
    assign layer4_outputs[1378] = ~((layer3_outputs[2174]) ^ (layer3_outputs[1877]));
    assign layer4_outputs[1379] = (layer3_outputs[483]) & (layer3_outputs[1390]);
    assign layer4_outputs[1380] = layer3_outputs[621];
    assign layer4_outputs[1381] = (layer3_outputs[2223]) ^ (layer3_outputs[984]);
    assign layer4_outputs[1382] = (layer3_outputs[363]) ^ (layer3_outputs[1123]);
    assign layer4_outputs[1383] = layer3_outputs[4];
    assign layer4_outputs[1384] = layer3_outputs[906];
    assign layer4_outputs[1385] = (layer3_outputs[1565]) & ~(layer3_outputs[506]);
    assign layer4_outputs[1386] = layer3_outputs[288];
    assign layer4_outputs[1387] = (layer3_outputs[2487]) & ~(layer3_outputs[605]);
    assign layer4_outputs[1388] = layer3_outputs[2194];
    assign layer4_outputs[1389] = (layer3_outputs[999]) ^ (layer3_outputs[215]);
    assign layer4_outputs[1390] = ~(layer3_outputs[2320]);
    assign layer4_outputs[1391] = (layer3_outputs[2382]) ^ (layer3_outputs[1185]);
    assign layer4_outputs[1392] = layer3_outputs[2553];
    assign layer4_outputs[1393] = ~(layer3_outputs[1335]);
    assign layer4_outputs[1394] = ~((layer3_outputs[2526]) & (layer3_outputs[2191]));
    assign layer4_outputs[1395] = ~((layer3_outputs[845]) & (layer3_outputs[73]));
    assign layer4_outputs[1396] = (layer3_outputs[290]) & ~(layer3_outputs[23]);
    assign layer4_outputs[1397] = ~((layer3_outputs[2517]) | (layer3_outputs[1816]));
    assign layer4_outputs[1398] = ~(layer3_outputs[328]);
    assign layer4_outputs[1399] = ~((layer3_outputs[1394]) | (layer3_outputs[1121]));
    assign layer4_outputs[1400] = layer3_outputs[213];
    assign layer4_outputs[1401] = ~(layer3_outputs[2133]);
    assign layer4_outputs[1402] = layer3_outputs[1728];
    assign layer4_outputs[1403] = ~(layer3_outputs[2164]);
    assign layer4_outputs[1404] = ~(layer3_outputs[1371]);
    assign layer4_outputs[1405] = (layer3_outputs[654]) ^ (layer3_outputs[893]);
    assign layer4_outputs[1406] = layer3_outputs[1195];
    assign layer4_outputs[1407] = ~(layer3_outputs[1768]) | (layer3_outputs[1612]);
    assign layer4_outputs[1408] = (layer3_outputs[2024]) ^ (layer3_outputs[1311]);
    assign layer4_outputs[1409] = ~(layer3_outputs[886]);
    assign layer4_outputs[1410] = ~((layer3_outputs[837]) & (layer3_outputs[590]));
    assign layer4_outputs[1411] = layer3_outputs[1586];
    assign layer4_outputs[1412] = layer3_outputs[362];
    assign layer4_outputs[1413] = layer3_outputs[1414];
    assign layer4_outputs[1414] = 1'b0;
    assign layer4_outputs[1415] = ~(layer3_outputs[542]);
    assign layer4_outputs[1416] = ~(layer3_outputs[1801]);
    assign layer4_outputs[1417] = (layer3_outputs[1310]) & ~(layer3_outputs[1143]);
    assign layer4_outputs[1418] = ~(layer3_outputs[800]) | (layer3_outputs[2113]);
    assign layer4_outputs[1419] = ~(layer3_outputs[613]);
    assign layer4_outputs[1420] = ~(layer3_outputs[285]);
    assign layer4_outputs[1421] = layer3_outputs[2234];
    assign layer4_outputs[1422] = layer3_outputs[675];
    assign layer4_outputs[1423] = ~((layer3_outputs[205]) & (layer3_outputs[1520]));
    assign layer4_outputs[1424] = layer3_outputs[2257];
    assign layer4_outputs[1425] = ~((layer3_outputs[2379]) | (layer3_outputs[2391]));
    assign layer4_outputs[1426] = layer3_outputs[1212];
    assign layer4_outputs[1427] = layer3_outputs[1473];
    assign layer4_outputs[1428] = (layer3_outputs[2474]) & (layer3_outputs[189]);
    assign layer4_outputs[1429] = ~(layer3_outputs[1763]);
    assign layer4_outputs[1430] = ~(layer3_outputs[618]) | (layer3_outputs[1854]);
    assign layer4_outputs[1431] = ~((layer3_outputs[1257]) & (layer3_outputs[1662]));
    assign layer4_outputs[1432] = layer3_outputs[1346];
    assign layer4_outputs[1433] = layer3_outputs[1899];
    assign layer4_outputs[1434] = (layer3_outputs[330]) & ~(layer3_outputs[610]);
    assign layer4_outputs[1435] = ~((layer3_outputs[1971]) ^ (layer3_outputs[2388]));
    assign layer4_outputs[1436] = ~(layer3_outputs[716]) | (layer3_outputs[1490]);
    assign layer4_outputs[1437] = (layer3_outputs[1762]) & (layer3_outputs[831]);
    assign layer4_outputs[1438] = (layer3_outputs[2032]) & ~(layer3_outputs[566]);
    assign layer4_outputs[1439] = ~(layer3_outputs[1999]);
    assign layer4_outputs[1440] = (layer3_outputs[876]) & (layer3_outputs[105]);
    assign layer4_outputs[1441] = ~((layer3_outputs[2353]) ^ (layer3_outputs[1512]));
    assign layer4_outputs[1442] = ~(layer3_outputs[1142]) | (layer3_outputs[451]);
    assign layer4_outputs[1443] = ~(layer3_outputs[1882]);
    assign layer4_outputs[1444] = layer3_outputs[1080];
    assign layer4_outputs[1445] = (layer3_outputs[1095]) | (layer3_outputs[1244]);
    assign layer4_outputs[1446] = ~((layer3_outputs[2105]) & (layer3_outputs[1612]));
    assign layer4_outputs[1447] = layer3_outputs[745];
    assign layer4_outputs[1448] = layer3_outputs[372];
    assign layer4_outputs[1449] = layer3_outputs[510];
    assign layer4_outputs[1450] = ~((layer3_outputs[2366]) & (layer3_outputs[1989]));
    assign layer4_outputs[1451] = (layer3_outputs[880]) | (layer3_outputs[1333]);
    assign layer4_outputs[1452] = ~(layer3_outputs[857]);
    assign layer4_outputs[1453] = (layer3_outputs[764]) & (layer3_outputs[1345]);
    assign layer4_outputs[1454] = ~((layer3_outputs[1174]) | (layer3_outputs[1816]));
    assign layer4_outputs[1455] = ~(layer3_outputs[587]);
    assign layer4_outputs[1456] = ~((layer3_outputs[479]) | (layer3_outputs[620]));
    assign layer4_outputs[1457] = (layer3_outputs[2215]) & ~(layer3_outputs[684]);
    assign layer4_outputs[1458] = ~(layer3_outputs[2350]);
    assign layer4_outputs[1459] = ~((layer3_outputs[2467]) | (layer3_outputs[67]));
    assign layer4_outputs[1460] = ~(layer3_outputs[711]);
    assign layer4_outputs[1461] = ~(layer3_outputs[454]);
    assign layer4_outputs[1462] = layer3_outputs[848];
    assign layer4_outputs[1463] = ~(layer3_outputs[38]) | (layer3_outputs[1309]);
    assign layer4_outputs[1464] = (layer3_outputs[341]) | (layer3_outputs[2542]);
    assign layer4_outputs[1465] = ~(layer3_outputs[2278]);
    assign layer4_outputs[1466] = ~((layer3_outputs[803]) & (layer3_outputs[1064]));
    assign layer4_outputs[1467] = ~(layer3_outputs[861]);
    assign layer4_outputs[1468] = (layer3_outputs[2365]) | (layer3_outputs[2406]);
    assign layer4_outputs[1469] = ~(layer3_outputs[2335]);
    assign layer4_outputs[1470] = (layer3_outputs[2130]) & ~(layer3_outputs[1589]);
    assign layer4_outputs[1471] = ~(layer3_outputs[1570]);
    assign layer4_outputs[1472] = (layer3_outputs[368]) ^ (layer3_outputs[1640]);
    assign layer4_outputs[1473] = (layer3_outputs[123]) & (layer3_outputs[24]);
    assign layer4_outputs[1474] = ~(layer3_outputs[556]);
    assign layer4_outputs[1475] = (layer3_outputs[916]) & (layer3_outputs[2360]);
    assign layer4_outputs[1476] = (layer3_outputs[1532]) ^ (layer3_outputs[2062]);
    assign layer4_outputs[1477] = (layer3_outputs[1137]) & ~(layer3_outputs[1825]);
    assign layer4_outputs[1478] = ~(layer3_outputs[2031]) | (layer3_outputs[2264]);
    assign layer4_outputs[1479] = (layer3_outputs[117]) | (layer3_outputs[2446]);
    assign layer4_outputs[1480] = ~(layer3_outputs[421]);
    assign layer4_outputs[1481] = layer3_outputs[692];
    assign layer4_outputs[1482] = ~((layer3_outputs[1746]) | (layer3_outputs[2015]));
    assign layer4_outputs[1483] = 1'b0;
    assign layer4_outputs[1484] = ~(layer3_outputs[1356]);
    assign layer4_outputs[1485] = ~((layer3_outputs[624]) | (layer3_outputs[1804]));
    assign layer4_outputs[1486] = ~(layer3_outputs[272]);
    assign layer4_outputs[1487] = layer3_outputs[523];
    assign layer4_outputs[1488] = 1'b0;
    assign layer4_outputs[1489] = (layer3_outputs[1325]) ^ (layer3_outputs[1097]);
    assign layer4_outputs[1490] = ~((layer3_outputs[1561]) ^ (layer3_outputs[1192]));
    assign layer4_outputs[1491] = layer3_outputs[2272];
    assign layer4_outputs[1492] = ~(layer3_outputs[2182]);
    assign layer4_outputs[1493] = ~(layer3_outputs[1150]);
    assign layer4_outputs[1494] = ~((layer3_outputs[433]) ^ (layer3_outputs[248]));
    assign layer4_outputs[1495] = ~(layer3_outputs[876]) | (layer3_outputs[846]);
    assign layer4_outputs[1496] = ~(layer3_outputs[2254]);
    assign layer4_outputs[1497] = layer3_outputs[2104];
    assign layer4_outputs[1498] = ~((layer3_outputs[2145]) & (layer3_outputs[461]));
    assign layer4_outputs[1499] = ~((layer3_outputs[157]) ^ (layer3_outputs[1062]));
    assign layer4_outputs[1500] = ~((layer3_outputs[1580]) & (layer3_outputs[93]));
    assign layer4_outputs[1501] = layer3_outputs[912];
    assign layer4_outputs[1502] = layer3_outputs[1329];
    assign layer4_outputs[1503] = layer3_outputs[2294];
    assign layer4_outputs[1504] = layer3_outputs[871];
    assign layer4_outputs[1505] = (layer3_outputs[824]) & ~(layer3_outputs[1426]);
    assign layer4_outputs[1506] = ~(layer3_outputs[2298]) | (layer3_outputs[120]);
    assign layer4_outputs[1507] = ~(layer3_outputs[1512]);
    assign layer4_outputs[1508] = ~((layer3_outputs[950]) & (layer3_outputs[1024]));
    assign layer4_outputs[1509] = layer3_outputs[2016];
    assign layer4_outputs[1510] = layer3_outputs[541];
    assign layer4_outputs[1511] = (layer3_outputs[1431]) ^ (layer3_outputs[2224]);
    assign layer4_outputs[1512] = ~((layer3_outputs[1823]) ^ (layer3_outputs[2044]));
    assign layer4_outputs[1513] = layer3_outputs[1859];
    assign layer4_outputs[1514] = (layer3_outputs[2359]) & ~(layer3_outputs[1706]);
    assign layer4_outputs[1515] = layer3_outputs[2291];
    assign layer4_outputs[1516] = (layer3_outputs[2281]) ^ (layer3_outputs[313]);
    assign layer4_outputs[1517] = 1'b1;
    assign layer4_outputs[1518] = (layer3_outputs[358]) & ~(layer3_outputs[343]);
    assign layer4_outputs[1519] = layer3_outputs[783];
    assign layer4_outputs[1520] = (layer3_outputs[1307]) & ~(layer3_outputs[1001]);
    assign layer4_outputs[1521] = ~(layer3_outputs[562]);
    assign layer4_outputs[1522] = ~((layer3_outputs[1600]) & (layer3_outputs[487]));
    assign layer4_outputs[1523] = (layer3_outputs[1019]) & ~(layer3_outputs[523]);
    assign layer4_outputs[1524] = ~((layer3_outputs[1111]) | (layer3_outputs[1336]));
    assign layer4_outputs[1525] = ~((layer3_outputs[1266]) | (layer3_outputs[216]));
    assign layer4_outputs[1526] = ~(layer3_outputs[1291]) | (layer3_outputs[1873]);
    assign layer4_outputs[1527] = layer3_outputs[1840];
    assign layer4_outputs[1528] = ~(layer3_outputs[2204]);
    assign layer4_outputs[1529] = ~(layer3_outputs[1915]);
    assign layer4_outputs[1530] = ~(layer3_outputs[576]);
    assign layer4_outputs[1531] = layer3_outputs[667];
    assign layer4_outputs[1532] = ~(layer3_outputs[1047]);
    assign layer4_outputs[1533] = layer3_outputs[149];
    assign layer4_outputs[1534] = ~(layer3_outputs[2393]) | (layer3_outputs[750]);
    assign layer4_outputs[1535] = ~((layer3_outputs[218]) | (layer3_outputs[1272]));
    assign layer4_outputs[1536] = (layer3_outputs[2168]) | (layer3_outputs[260]);
    assign layer4_outputs[1537] = layer3_outputs[1457];
    assign layer4_outputs[1538] = (layer3_outputs[1419]) & ~(layer3_outputs[1616]);
    assign layer4_outputs[1539] = (layer3_outputs[1697]) ^ (layer3_outputs[1058]);
    assign layer4_outputs[1540] = layer3_outputs[2229];
    assign layer4_outputs[1541] = (layer3_outputs[1018]) | (layer3_outputs[1067]);
    assign layer4_outputs[1542] = ~(layer3_outputs[1]);
    assign layer4_outputs[1543] = ~(layer3_outputs[627]);
    assign layer4_outputs[1544] = (layer3_outputs[1363]) ^ (layer3_outputs[2050]);
    assign layer4_outputs[1545] = ~((layer3_outputs[1055]) & (layer3_outputs[2107]));
    assign layer4_outputs[1546] = ~(layer3_outputs[330]);
    assign layer4_outputs[1547] = (layer3_outputs[1904]) & ~(layer3_outputs[1451]);
    assign layer4_outputs[1548] = ~(layer3_outputs[2480]);
    assign layer4_outputs[1549] = ~(layer3_outputs[1116]);
    assign layer4_outputs[1550] = ~(layer3_outputs[741]);
    assign layer4_outputs[1551] = ~(layer3_outputs[1973]);
    assign layer4_outputs[1552] = ~(layer3_outputs[1148]) | (layer3_outputs[199]);
    assign layer4_outputs[1553] = layer3_outputs[27];
    assign layer4_outputs[1554] = (layer3_outputs[146]) & ~(layer3_outputs[52]);
    assign layer4_outputs[1555] = layer3_outputs[244];
    assign layer4_outputs[1556] = ~(layer3_outputs[814]) | (layer3_outputs[2032]);
    assign layer4_outputs[1557] = (layer3_outputs[190]) ^ (layer3_outputs[1890]);
    assign layer4_outputs[1558] = ~((layer3_outputs[2323]) & (layer3_outputs[2493]));
    assign layer4_outputs[1559] = ~(layer3_outputs[443]);
    assign layer4_outputs[1560] = (layer3_outputs[1688]) | (layer3_outputs[1362]);
    assign layer4_outputs[1561] = layer3_outputs[329];
    assign layer4_outputs[1562] = layer3_outputs[2525];
    assign layer4_outputs[1563] = ~(layer3_outputs[498]) | (layer3_outputs[2169]);
    assign layer4_outputs[1564] = ~(layer3_outputs[347]);
    assign layer4_outputs[1565] = layer3_outputs[134];
    assign layer4_outputs[1566] = ~((layer3_outputs[1993]) | (layer3_outputs[878]));
    assign layer4_outputs[1567] = ~(layer3_outputs[111]);
    assign layer4_outputs[1568] = ~(layer3_outputs[1440]) | (layer3_outputs[2010]);
    assign layer4_outputs[1569] = ~(layer3_outputs[424]);
    assign layer4_outputs[1570] = ~(layer3_outputs[630]);
    assign layer4_outputs[1571] = layer3_outputs[1981];
    assign layer4_outputs[1572] = layer3_outputs[996];
    assign layer4_outputs[1573] = (layer3_outputs[1747]) & ~(layer3_outputs[396]);
    assign layer4_outputs[1574] = ~(layer3_outputs[1135]) | (layer3_outputs[1309]);
    assign layer4_outputs[1575] = (layer3_outputs[1720]) | (layer3_outputs[686]);
    assign layer4_outputs[1576] = ~(layer3_outputs[1315]);
    assign layer4_outputs[1577] = layer3_outputs[669];
    assign layer4_outputs[1578] = layer3_outputs[1496];
    assign layer4_outputs[1579] = ~((layer3_outputs[1224]) ^ (layer3_outputs[703]));
    assign layer4_outputs[1580] = ~(layer3_outputs[2445]);
    assign layer4_outputs[1581] = ~(layer3_outputs[573]);
    assign layer4_outputs[1582] = (layer3_outputs[1722]) ^ (layer3_outputs[1228]);
    assign layer4_outputs[1583] = layer3_outputs[1944];
    assign layer4_outputs[1584] = (layer3_outputs[2315]) & ~(layer3_outputs[2234]);
    assign layer4_outputs[1585] = ~((layer3_outputs[1566]) & (layer3_outputs[1703]));
    assign layer4_outputs[1586] = layer3_outputs[1873];
    assign layer4_outputs[1587] = 1'b0;
    assign layer4_outputs[1588] = ~(layer3_outputs[79]) | (layer3_outputs[873]);
    assign layer4_outputs[1589] = layer3_outputs[1832];
    assign layer4_outputs[1590] = ~(layer3_outputs[669]) | (layer3_outputs[825]);
    assign layer4_outputs[1591] = (layer3_outputs[1346]) & (layer3_outputs[1165]);
    assign layer4_outputs[1592] = ~((layer3_outputs[835]) & (layer3_outputs[2293]));
    assign layer4_outputs[1593] = ~(layer3_outputs[2106]);
    assign layer4_outputs[1594] = ~(layer3_outputs[2175]);
    assign layer4_outputs[1595] = ~(layer3_outputs[2152]);
    assign layer4_outputs[1596] = ~(layer3_outputs[1260]) | (layer3_outputs[122]);
    assign layer4_outputs[1597] = layer3_outputs[1048];
    assign layer4_outputs[1598] = ~(layer3_outputs[894]);
    assign layer4_outputs[1599] = (layer3_outputs[265]) | (layer3_outputs[2443]);
    assign layer4_outputs[1600] = ~(layer3_outputs[1105]);
    assign layer4_outputs[1601] = layer3_outputs[1380];
    assign layer4_outputs[1602] = layer3_outputs[1967];
    assign layer4_outputs[1603] = ~(layer3_outputs[2309]);
    assign layer4_outputs[1604] = layer3_outputs[968];
    assign layer4_outputs[1605] = (layer3_outputs[736]) | (layer3_outputs[488]);
    assign layer4_outputs[1606] = ~((layer3_outputs[803]) & (layer3_outputs[442]));
    assign layer4_outputs[1607] = ~((layer3_outputs[1466]) | (layer3_outputs[209]));
    assign layer4_outputs[1608] = ~(layer3_outputs[708]);
    assign layer4_outputs[1609] = layer3_outputs[908];
    assign layer4_outputs[1610] = ~((layer3_outputs[2343]) ^ (layer3_outputs[673]));
    assign layer4_outputs[1611] = ~((layer3_outputs[1323]) ^ (layer3_outputs[2187]));
    assign layer4_outputs[1612] = ~(layer3_outputs[705]);
    assign layer4_outputs[1613] = ~(layer3_outputs[1322]);
    assign layer4_outputs[1614] = ~(layer3_outputs[2449]);
    assign layer4_outputs[1615] = layer3_outputs[228];
    assign layer4_outputs[1616] = layer3_outputs[142];
    assign layer4_outputs[1617] = ~(layer3_outputs[1095]);
    assign layer4_outputs[1618] = ~(layer3_outputs[2142]) | (layer3_outputs[256]);
    assign layer4_outputs[1619] = layer3_outputs[1416];
    assign layer4_outputs[1620] = layer3_outputs[1895];
    assign layer4_outputs[1621] = layer3_outputs[71];
    assign layer4_outputs[1622] = layer3_outputs[424];
    assign layer4_outputs[1623] = ~(layer3_outputs[177]);
    assign layer4_outputs[1624] = ~(layer3_outputs[1914]);
    assign layer4_outputs[1625] = layer3_outputs[1974];
    assign layer4_outputs[1626] = (layer3_outputs[2493]) | (layer3_outputs[1789]);
    assign layer4_outputs[1627] = (layer3_outputs[1911]) & (layer3_outputs[606]);
    assign layer4_outputs[1628] = ~(layer3_outputs[1145]) | (layer3_outputs[1606]);
    assign layer4_outputs[1629] = ~((layer3_outputs[786]) ^ (layer3_outputs[2170]));
    assign layer4_outputs[1630] = ~(layer3_outputs[2550]) | (layer3_outputs[2453]);
    assign layer4_outputs[1631] = ~(layer3_outputs[1510]);
    assign layer4_outputs[1632] = ~((layer3_outputs[2358]) & (layer3_outputs[2164]));
    assign layer4_outputs[1633] = layer3_outputs[2159];
    assign layer4_outputs[1634] = ~((layer3_outputs[2347]) & (layer3_outputs[2547]));
    assign layer4_outputs[1635] = layer3_outputs[263];
    assign layer4_outputs[1636] = layer3_outputs[1801];
    assign layer4_outputs[1637] = ~(layer3_outputs[671]);
    assign layer4_outputs[1638] = (layer3_outputs[1642]) & ~(layer3_outputs[2556]);
    assign layer4_outputs[1639] = (layer3_outputs[543]) | (layer3_outputs[1969]);
    assign layer4_outputs[1640] = layer3_outputs[1835];
    assign layer4_outputs[1641] = layer3_outputs[1368];
    assign layer4_outputs[1642] = ~(layer3_outputs[1646]);
    assign layer4_outputs[1643] = ~(layer3_outputs[290]) | (layer3_outputs[1883]);
    assign layer4_outputs[1644] = (layer3_outputs[1556]) | (layer3_outputs[1142]);
    assign layer4_outputs[1645] = ~(layer3_outputs[149]);
    assign layer4_outputs[1646] = (layer3_outputs[2364]) & ~(layer3_outputs[522]);
    assign layer4_outputs[1647] = ~(layer3_outputs[1608]);
    assign layer4_outputs[1648] = ~(layer3_outputs[630]);
    assign layer4_outputs[1649] = (layer3_outputs[1796]) ^ (layer3_outputs[77]);
    assign layer4_outputs[1650] = ~(layer3_outputs[2326]);
    assign layer4_outputs[1651] = ~(layer3_outputs[1817]);
    assign layer4_outputs[1652] = (layer3_outputs[897]) & (layer3_outputs[2122]);
    assign layer4_outputs[1653] = (layer3_outputs[368]) & (layer3_outputs[913]);
    assign layer4_outputs[1654] = (layer3_outputs[1591]) & (layer3_outputs[2034]);
    assign layer4_outputs[1655] = ~(layer3_outputs[9]);
    assign layer4_outputs[1656] = 1'b1;
    assign layer4_outputs[1657] = ~(layer3_outputs[562]) | (layer3_outputs[2357]);
    assign layer4_outputs[1658] = (layer3_outputs[5]) & ~(layer3_outputs[82]);
    assign layer4_outputs[1659] = (layer3_outputs[466]) & ~(layer3_outputs[1111]);
    assign layer4_outputs[1660] = ~((layer3_outputs[802]) ^ (layer3_outputs[1130]));
    assign layer4_outputs[1661] = ~(layer3_outputs[1996]);
    assign layer4_outputs[1662] = ~(layer3_outputs[489]);
    assign layer4_outputs[1663] = layer3_outputs[2246];
    assign layer4_outputs[1664] = (layer3_outputs[1564]) & ~(layer3_outputs[734]);
    assign layer4_outputs[1665] = (layer3_outputs[653]) & ~(layer3_outputs[1556]);
    assign layer4_outputs[1666] = (layer3_outputs[1947]) ^ (layer3_outputs[1155]);
    assign layer4_outputs[1667] = ~(layer3_outputs[308]);
    assign layer4_outputs[1668] = layer3_outputs[1689];
    assign layer4_outputs[1669] = layer3_outputs[2504];
    assign layer4_outputs[1670] = ~(layer3_outputs[163]) | (layer3_outputs[1935]);
    assign layer4_outputs[1671] = ~(layer3_outputs[1903]);
    assign layer4_outputs[1672] = (layer3_outputs[836]) | (layer3_outputs[795]);
    assign layer4_outputs[1673] = layer3_outputs[1544];
    assign layer4_outputs[1674] = ~(layer3_outputs[2244]) | (layer3_outputs[2150]);
    assign layer4_outputs[1675] = ~((layer3_outputs[841]) & (layer3_outputs[2068]));
    assign layer4_outputs[1676] = ~(layer3_outputs[2012]) | (layer3_outputs[980]);
    assign layer4_outputs[1677] = ~((layer3_outputs[1630]) | (layer3_outputs[1608]));
    assign layer4_outputs[1678] = ~(layer3_outputs[764]);
    assign layer4_outputs[1679] = ~(layer3_outputs[771]);
    assign layer4_outputs[1680] = 1'b1;
    assign layer4_outputs[1681] = ~((layer3_outputs[946]) & (layer3_outputs[1365]));
    assign layer4_outputs[1682] = layer3_outputs[1199];
    assign layer4_outputs[1683] = ~((layer3_outputs[224]) ^ (layer3_outputs[2500]));
    assign layer4_outputs[1684] = layer3_outputs[48];
    assign layer4_outputs[1685] = (layer3_outputs[918]) & ~(layer3_outputs[1661]);
    assign layer4_outputs[1686] = (layer3_outputs[2375]) & (layer3_outputs[2245]);
    assign layer4_outputs[1687] = layer3_outputs[941];
    assign layer4_outputs[1688] = 1'b0;
    assign layer4_outputs[1689] = ~(layer3_outputs[2519]);
    assign layer4_outputs[1690] = ~(layer3_outputs[2142]);
    assign layer4_outputs[1691] = layer3_outputs[410];
    assign layer4_outputs[1692] = ~((layer3_outputs[1947]) ^ (layer3_outputs[391]));
    assign layer4_outputs[1693] = ~(layer3_outputs[2231]);
    assign layer4_outputs[1694] = layer3_outputs[2183];
    assign layer4_outputs[1695] = (layer3_outputs[1864]) & ~(layer3_outputs[750]);
    assign layer4_outputs[1696] = ~(layer3_outputs[542]);
    assign layer4_outputs[1697] = ~((layer3_outputs[1222]) & (layer3_outputs[340]));
    assign layer4_outputs[1698] = layer3_outputs[650];
    assign layer4_outputs[1699] = ~((layer3_outputs[1065]) ^ (layer3_outputs[1009]));
    assign layer4_outputs[1700] = layer3_outputs[1227];
    assign layer4_outputs[1701] = layer3_outputs[1981];
    assign layer4_outputs[1702] = (layer3_outputs[195]) & ~(layer3_outputs[665]);
    assign layer4_outputs[1703] = ~(layer3_outputs[1908]);
    assign layer4_outputs[1704] = (layer3_outputs[1576]) & ~(layer3_outputs[1878]);
    assign layer4_outputs[1705] = (layer3_outputs[94]) & (layer3_outputs[2350]);
    assign layer4_outputs[1706] = layer3_outputs[62];
    assign layer4_outputs[1707] = layer3_outputs[1104];
    assign layer4_outputs[1708] = ~(layer3_outputs[1525]);
    assign layer4_outputs[1709] = (layer3_outputs[206]) ^ (layer3_outputs[569]);
    assign layer4_outputs[1710] = ~((layer3_outputs[1249]) ^ (layer3_outputs[2019]));
    assign layer4_outputs[1711] = layer3_outputs[757];
    assign layer4_outputs[1712] = ~((layer3_outputs[1535]) & (layer3_outputs[1744]));
    assign layer4_outputs[1713] = ~((layer3_outputs[1067]) & (layer3_outputs[1697]));
    assign layer4_outputs[1714] = ~((layer3_outputs[359]) | (layer3_outputs[92]));
    assign layer4_outputs[1715] = ~((layer3_outputs[1203]) & (layer3_outputs[396]));
    assign layer4_outputs[1716] = ~((layer3_outputs[456]) ^ (layer3_outputs[1416]));
    assign layer4_outputs[1717] = layer3_outputs[1337];
    assign layer4_outputs[1718] = ~(layer3_outputs[865]);
    assign layer4_outputs[1719] = (layer3_outputs[1589]) & (layer3_outputs[1833]);
    assign layer4_outputs[1720] = ~((layer3_outputs[1367]) & (layer3_outputs[1491]));
    assign layer4_outputs[1721] = layer3_outputs[939];
    assign layer4_outputs[1722] = ~(layer3_outputs[323]);
    assign layer4_outputs[1723] = ~((layer3_outputs[722]) | (layer3_outputs[2538]));
    assign layer4_outputs[1724] = layer3_outputs[526];
    assign layer4_outputs[1725] = ~(layer3_outputs[2085]);
    assign layer4_outputs[1726] = ~(layer3_outputs[1175]);
    assign layer4_outputs[1727] = ~(layer3_outputs[33]);
    assign layer4_outputs[1728] = (layer3_outputs[1631]) ^ (layer3_outputs[1513]);
    assign layer4_outputs[1729] = layer3_outputs[2340];
    assign layer4_outputs[1730] = ~((layer3_outputs[252]) ^ (layer3_outputs[721]));
    assign layer4_outputs[1731] = (layer3_outputs[15]) & ~(layer3_outputs[2021]);
    assign layer4_outputs[1732] = layer3_outputs[178];
    assign layer4_outputs[1733] = layer3_outputs[395];
    assign layer4_outputs[1734] = layer3_outputs[581];
    assign layer4_outputs[1735] = layer3_outputs[1207];
    assign layer4_outputs[1736] = ~(layer3_outputs[2319]);
    assign layer4_outputs[1737] = (layer3_outputs[2515]) | (layer3_outputs[521]);
    assign layer4_outputs[1738] = (layer3_outputs[1156]) & ~(layer3_outputs[1710]);
    assign layer4_outputs[1739] = ~(layer3_outputs[95]);
    assign layer4_outputs[1740] = ~((layer3_outputs[2133]) ^ (layer3_outputs[928]));
    assign layer4_outputs[1741] = ~(layer3_outputs[1773]);
    assign layer4_outputs[1742] = ~((layer3_outputs[1630]) | (layer3_outputs[2145]));
    assign layer4_outputs[1743] = (layer3_outputs[1453]) ^ (layer3_outputs[325]);
    assign layer4_outputs[1744] = (layer3_outputs[820]) & ~(layer3_outputs[615]);
    assign layer4_outputs[1745] = (layer3_outputs[1513]) ^ (layer3_outputs[1686]);
    assign layer4_outputs[1746] = ~(layer3_outputs[1166]);
    assign layer4_outputs[1747] = (layer3_outputs[1193]) & ~(layer3_outputs[790]);
    assign layer4_outputs[1748] = ~((layer3_outputs[1471]) & (layer3_outputs[436]));
    assign layer4_outputs[1749] = ~(layer3_outputs[1884]) | (layer3_outputs[1241]);
    assign layer4_outputs[1750] = (layer3_outputs[133]) & ~(layer3_outputs[947]);
    assign layer4_outputs[1751] = ~(layer3_outputs[1096]) | (layer3_outputs[1028]);
    assign layer4_outputs[1752] = ~(layer3_outputs[2190]) | (layer3_outputs[1197]);
    assign layer4_outputs[1753] = ~(layer3_outputs[1681]);
    assign layer4_outputs[1754] = ~((layer3_outputs[579]) ^ (layer3_outputs[1134]));
    assign layer4_outputs[1755] = (layer3_outputs[2158]) ^ (layer3_outputs[11]);
    assign layer4_outputs[1756] = ~(layer3_outputs[1194]) | (layer3_outputs[1953]);
    assign layer4_outputs[1757] = (layer3_outputs[2558]) & ~(layer3_outputs[2457]);
    assign layer4_outputs[1758] = (layer3_outputs[1984]) & (layer3_outputs[1959]);
    assign layer4_outputs[1759] = (layer3_outputs[2320]) & (layer3_outputs[1551]);
    assign layer4_outputs[1760] = (layer3_outputs[1714]) & ~(layer3_outputs[1055]);
    assign layer4_outputs[1761] = ~(layer3_outputs[2296]);
    assign layer4_outputs[1762] = (layer3_outputs[1050]) | (layer3_outputs[2005]);
    assign layer4_outputs[1763] = ~(layer3_outputs[1509]);
    assign layer4_outputs[1764] = layer3_outputs[642];
    assign layer4_outputs[1765] = (layer3_outputs[619]) & ~(layer3_outputs[2155]);
    assign layer4_outputs[1766] = ~(layer3_outputs[2404]);
    assign layer4_outputs[1767] = layer3_outputs[1285];
    assign layer4_outputs[1768] = layer3_outputs[1181];
    assign layer4_outputs[1769] = ~((layer3_outputs[554]) ^ (layer3_outputs[2325]));
    assign layer4_outputs[1770] = ~((layer3_outputs[2486]) | (layer3_outputs[2237]));
    assign layer4_outputs[1771] = ~(layer3_outputs[1649]) | (layer3_outputs[1820]);
    assign layer4_outputs[1772] = layer3_outputs[377];
    assign layer4_outputs[1773] = layer3_outputs[2390];
    assign layer4_outputs[1774] = ~((layer3_outputs[317]) & (layer3_outputs[1840]));
    assign layer4_outputs[1775] = ~((layer3_outputs[171]) | (layer3_outputs[1480]));
    assign layer4_outputs[1776] = ~(layer3_outputs[1263]);
    assign layer4_outputs[1777] = ~(layer3_outputs[1462]);
    assign layer4_outputs[1778] = ~(layer3_outputs[1684]);
    assign layer4_outputs[1779] = layer3_outputs[1075];
    assign layer4_outputs[1780] = ~(layer3_outputs[30]);
    assign layer4_outputs[1781] = (layer3_outputs[2356]) & (layer3_outputs[262]);
    assign layer4_outputs[1782] = layer3_outputs[980];
    assign layer4_outputs[1783] = 1'b0;
    assign layer4_outputs[1784] = ~((layer3_outputs[952]) ^ (layer3_outputs[969]));
    assign layer4_outputs[1785] = layer3_outputs[63];
    assign layer4_outputs[1786] = ~((layer3_outputs[1830]) | (layer3_outputs[1695]));
    assign layer4_outputs[1787] = ~((layer3_outputs[203]) | (layer3_outputs[853]));
    assign layer4_outputs[1788] = ~(layer3_outputs[366]) | (layer3_outputs[600]);
    assign layer4_outputs[1789] = ~(layer3_outputs[427]);
    assign layer4_outputs[1790] = (layer3_outputs[1886]) ^ (layer3_outputs[1691]);
    assign layer4_outputs[1791] = ~(layer3_outputs[1389]) | (layer3_outputs[2136]);
    assign layer4_outputs[1792] = ~(layer3_outputs[2288]) | (layer3_outputs[2180]);
    assign layer4_outputs[1793] = (layer3_outputs[2163]) & ~(layer3_outputs[2252]);
    assign layer4_outputs[1794] = layer3_outputs[243];
    assign layer4_outputs[1795] = ~((layer3_outputs[1715]) | (layer3_outputs[1129]));
    assign layer4_outputs[1796] = ~(layer3_outputs[2541]) | (layer3_outputs[569]);
    assign layer4_outputs[1797] = ~(layer3_outputs[1631]);
    assign layer4_outputs[1798] = ~((layer3_outputs[970]) & (layer3_outputs[1879]));
    assign layer4_outputs[1799] = layer3_outputs[1010];
    assign layer4_outputs[1800] = (layer3_outputs[2238]) & (layer3_outputs[93]);
    assign layer4_outputs[1801] = (layer3_outputs[2422]) & ~(layer3_outputs[401]);
    assign layer4_outputs[1802] = ~(layer3_outputs[621]);
    assign layer4_outputs[1803] = layer3_outputs[1026];
    assign layer4_outputs[1804] = layer3_outputs[2030];
    assign layer4_outputs[1805] = (layer3_outputs[135]) | (layer3_outputs[1362]);
    assign layer4_outputs[1806] = (layer3_outputs[1780]) & ~(layer3_outputs[1022]);
    assign layer4_outputs[1807] = (layer3_outputs[666]) & (layer3_outputs[681]);
    assign layer4_outputs[1808] = ~(layer3_outputs[1951]);
    assign layer4_outputs[1809] = ~((layer3_outputs[1833]) ^ (layer3_outputs[431]));
    assign layer4_outputs[1810] = ~(layer3_outputs[1475]);
    assign layer4_outputs[1811] = ~((layer3_outputs[237]) | (layer3_outputs[2051]));
    assign layer4_outputs[1812] = (layer3_outputs[509]) & ~(layer3_outputs[331]);
    assign layer4_outputs[1813] = ~(layer3_outputs[662]);
    assign layer4_outputs[1814] = ~(layer3_outputs[334]) | (layer3_outputs[810]);
    assign layer4_outputs[1815] = ~(layer3_outputs[2229]) | (layer3_outputs[295]);
    assign layer4_outputs[1816] = layer3_outputs[1888];
    assign layer4_outputs[1817] = ~(layer3_outputs[1698]);
    assign layer4_outputs[1818] = layer3_outputs[1686];
    assign layer4_outputs[1819] = layer3_outputs[141];
    assign layer4_outputs[1820] = ~(layer3_outputs[987]) | (layer3_outputs[1967]);
    assign layer4_outputs[1821] = (layer3_outputs[175]) ^ (layer3_outputs[805]);
    assign layer4_outputs[1822] = ~(layer3_outputs[2202]);
    assign layer4_outputs[1823] = ~(layer3_outputs[674]);
    assign layer4_outputs[1824] = 1'b0;
    assign layer4_outputs[1825] = (layer3_outputs[2192]) ^ (layer3_outputs[821]);
    assign layer4_outputs[1826] = layer3_outputs[1600];
    assign layer4_outputs[1827] = ~((layer3_outputs[2232]) & (layer3_outputs[1268]));
    assign layer4_outputs[1828] = ~(layer3_outputs[2440]);
    assign layer4_outputs[1829] = ~(layer3_outputs[1719]);
    assign layer4_outputs[1830] = ~(layer3_outputs[2213]) | (layer3_outputs[276]);
    assign layer4_outputs[1831] = ~(layer3_outputs[1477]) | (layer3_outputs[2328]);
    assign layer4_outputs[1832] = layer3_outputs[2492];
    assign layer4_outputs[1833] = layer3_outputs[414];
    assign layer4_outputs[1834] = ~(layer3_outputs[75]);
    assign layer4_outputs[1835] = 1'b0;
    assign layer4_outputs[1836] = ~((layer3_outputs[796]) ^ (layer3_outputs[494]));
    assign layer4_outputs[1837] = layer3_outputs[333];
    assign layer4_outputs[1838] = ~(layer3_outputs[2496]);
    assign layer4_outputs[1839] = ~((layer3_outputs[812]) ^ (layer3_outputs[1113]));
    assign layer4_outputs[1840] = ~((layer3_outputs[2373]) ^ (layer3_outputs[74]));
    assign layer4_outputs[1841] = (layer3_outputs[116]) | (layer3_outputs[2258]);
    assign layer4_outputs[1842] = ~((layer3_outputs[172]) ^ (layer3_outputs[1928]));
    assign layer4_outputs[1843] = ~(layer3_outputs[1338]);
    assign layer4_outputs[1844] = ~(layer3_outputs[1571]) | (layer3_outputs[2171]);
    assign layer4_outputs[1845] = (layer3_outputs[1727]) & ~(layer3_outputs[1811]);
    assign layer4_outputs[1846] = ~(layer3_outputs[868]) | (layer3_outputs[129]);
    assign layer4_outputs[1847] = ~(layer3_outputs[603]);
    assign layer4_outputs[1848] = ~(layer3_outputs[1025]) | (layer3_outputs[1225]);
    assign layer4_outputs[1849] = (layer3_outputs[1481]) | (layer3_outputs[1259]);
    assign layer4_outputs[1850] = ~(layer3_outputs[127]);
    assign layer4_outputs[1851] = ~(layer3_outputs[1962]);
    assign layer4_outputs[1852] = ~(layer3_outputs[1459]) | (layer3_outputs[2179]);
    assign layer4_outputs[1853] = ~(layer3_outputs[2060]) | (layer3_outputs[2153]);
    assign layer4_outputs[1854] = (layer3_outputs[49]) & (layer3_outputs[445]);
    assign layer4_outputs[1855] = (layer3_outputs[114]) & ~(layer3_outputs[1433]);
    assign layer4_outputs[1856] = ~(layer3_outputs[457]) | (layer3_outputs[732]);
    assign layer4_outputs[1857] = (layer3_outputs[47]) & ~(layer3_outputs[1171]);
    assign layer4_outputs[1858] = ~(layer3_outputs[1892]);
    assign layer4_outputs[1859] = ~(layer3_outputs[460]);
    assign layer4_outputs[1860] = (layer3_outputs[1949]) & (layer3_outputs[1560]);
    assign layer4_outputs[1861] = ~(layer3_outputs[577]);
    assign layer4_outputs[1862] = ~(layer3_outputs[207]);
    assign layer4_outputs[1863] = ~(layer3_outputs[156]) | (layer3_outputs[663]);
    assign layer4_outputs[1864] = ~((layer3_outputs[1379]) & (layer3_outputs[1034]));
    assign layer4_outputs[1865] = layer3_outputs[34];
    assign layer4_outputs[1866] = ~(layer3_outputs[1126]);
    assign layer4_outputs[1867] = ~(layer3_outputs[1921]);
    assign layer4_outputs[1868] = layer3_outputs[1758];
    assign layer4_outputs[1869] = ~(layer3_outputs[1903]);
    assign layer4_outputs[1870] = ~(layer3_outputs[2452]) | (layer3_outputs[1202]);
    assign layer4_outputs[1871] = ~(layer3_outputs[192]);
    assign layer4_outputs[1872] = ~(layer3_outputs[777]);
    assign layer4_outputs[1873] = 1'b0;
    assign layer4_outputs[1874] = ~((layer3_outputs[1696]) & (layer3_outputs[1643]));
    assign layer4_outputs[1875] = (layer3_outputs[1799]) & (layer3_outputs[1579]);
    assign layer4_outputs[1876] = ~((layer3_outputs[2025]) ^ (layer3_outputs[1831]));
    assign layer4_outputs[1877] = ~((layer3_outputs[160]) ^ (layer3_outputs[1592]));
    assign layer4_outputs[1878] = (layer3_outputs[2101]) & ~(layer3_outputs[1138]);
    assign layer4_outputs[1879] = (layer3_outputs[588]) | (layer3_outputs[2554]);
    assign layer4_outputs[1880] = ~(layer3_outputs[2106]) | (layer3_outputs[688]);
    assign layer4_outputs[1881] = layer3_outputs[2009];
    assign layer4_outputs[1882] = ~((layer3_outputs[2121]) ^ (layer3_outputs[1074]));
    assign layer4_outputs[1883] = ~((layer3_outputs[877]) ^ (layer3_outputs[1758]));
    assign layer4_outputs[1884] = (layer3_outputs[2519]) & ~(layer3_outputs[919]);
    assign layer4_outputs[1885] = (layer3_outputs[2046]) | (layer3_outputs[1575]);
    assign layer4_outputs[1886] = ~(layer3_outputs[768]);
    assign layer4_outputs[1887] = ~(layer3_outputs[1419]);
    assign layer4_outputs[1888] = ~((layer3_outputs[1068]) ^ (layer3_outputs[2547]));
    assign layer4_outputs[1889] = 1'b0;
    assign layer4_outputs[1890] = ~((layer3_outputs[2279]) | (layer3_outputs[539]));
    assign layer4_outputs[1891] = ~(layer3_outputs[2265]) | (layer3_outputs[895]);
    assign layer4_outputs[1892] = layer3_outputs[1574];
    assign layer4_outputs[1893] = layer3_outputs[534];
    assign layer4_outputs[1894] = (layer3_outputs[1740]) & ~(layer3_outputs[1308]);
    assign layer4_outputs[1895] = (layer3_outputs[349]) & ~(layer3_outputs[875]);
    assign layer4_outputs[1896] = ~((layer3_outputs[2514]) | (layer3_outputs[356]));
    assign layer4_outputs[1897] = ~(layer3_outputs[2300]) | (layer3_outputs[1607]);
    assign layer4_outputs[1898] = ~(layer3_outputs[1626]);
    assign layer4_outputs[1899] = layer3_outputs[1862];
    assign layer4_outputs[1900] = layer3_outputs[333];
    assign layer4_outputs[1901] = ~(layer3_outputs[1468]) | (layer3_outputs[1553]);
    assign layer4_outputs[1902] = (layer3_outputs[1157]) & (layer3_outputs[1625]);
    assign layer4_outputs[1903] = ~(layer3_outputs[2108]) | (layer3_outputs[522]);
    assign layer4_outputs[1904] = ~(layer3_outputs[1684]);
    assign layer4_outputs[1905] = ~(layer3_outputs[2251]) | (layer3_outputs[2216]);
    assign layer4_outputs[1906] = layer3_outputs[516];
    assign layer4_outputs[1907] = (layer3_outputs[1099]) ^ (layer3_outputs[928]);
    assign layer4_outputs[1908] = ~(layer3_outputs[1580]);
    assign layer4_outputs[1909] = ~((layer3_outputs[2099]) ^ (layer3_outputs[1196]));
    assign layer4_outputs[1910] = (layer3_outputs[378]) ^ (layer3_outputs[877]);
    assign layer4_outputs[1911] = ~((layer3_outputs[919]) ^ (layer3_outputs[2196]));
    assign layer4_outputs[1912] = (layer3_outputs[912]) ^ (layer3_outputs[815]);
    assign layer4_outputs[1913] = ~(layer3_outputs[925]);
    assign layer4_outputs[1914] = layer3_outputs[176];
    assign layer4_outputs[1915] = layer3_outputs[1290];
    assign layer4_outputs[1916] = layer3_outputs[1573];
    assign layer4_outputs[1917] = ~(layer3_outputs[1756]);
    assign layer4_outputs[1918] = ~(layer3_outputs[40]);
    assign layer4_outputs[1919] = 1'b1;
    assign layer4_outputs[1920] = ~(layer3_outputs[472]);
    assign layer4_outputs[1921] = ~((layer3_outputs[1672]) | (layer3_outputs[2233]));
    assign layer4_outputs[1922] = (layer3_outputs[567]) | (layer3_outputs[1702]);
    assign layer4_outputs[1923] = ~(layer3_outputs[215]) | (layer3_outputs[1288]);
    assign layer4_outputs[1924] = ~(layer3_outputs[1527]) | (layer3_outputs[933]);
    assign layer4_outputs[1925] = layer3_outputs[39];
    assign layer4_outputs[1926] = ~(layer3_outputs[578]);
    assign layer4_outputs[1927] = ~((layer3_outputs[528]) ^ (layer3_outputs[974]));
    assign layer4_outputs[1928] = 1'b1;
    assign layer4_outputs[1929] = ~(layer3_outputs[1276]);
    assign layer4_outputs[1930] = layer3_outputs[2322];
    assign layer4_outputs[1931] = layer3_outputs[2131];
    assign layer4_outputs[1932] = (layer3_outputs[1538]) & ~(layer3_outputs[1533]);
    assign layer4_outputs[1933] = (layer3_outputs[1281]) | (layer3_outputs[1839]);
    assign layer4_outputs[1934] = ~(layer3_outputs[908]);
    assign layer4_outputs[1935] = layer3_outputs[871];
    assign layer4_outputs[1936] = layer3_outputs[538];
    assign layer4_outputs[1937] = (layer3_outputs[1059]) & (layer3_outputs[1568]);
    assign layer4_outputs[1938] = (layer3_outputs[255]) | (layer3_outputs[2077]);
    assign layer4_outputs[1939] = (layer3_outputs[1540]) ^ (layer3_outputs[1813]);
    assign layer4_outputs[1940] = layer3_outputs[718];
    assign layer4_outputs[1941] = ~(layer3_outputs[185]);
    assign layer4_outputs[1942] = ~((layer3_outputs[613]) & (layer3_outputs[1699]));
    assign layer4_outputs[1943] = (layer3_outputs[532]) & ~(layer3_outputs[1619]);
    assign layer4_outputs[1944] = (layer3_outputs[402]) | (layer3_outputs[1785]);
    assign layer4_outputs[1945] = ~(layer3_outputs[1581]) | (layer3_outputs[1243]);
    assign layer4_outputs[1946] = layer3_outputs[1741];
    assign layer4_outputs[1947] = (layer3_outputs[1446]) & ~(layer3_outputs[1323]);
    assign layer4_outputs[1948] = layer3_outputs[1299];
    assign layer4_outputs[1949] = 1'b1;
    assign layer4_outputs[1950] = ~(layer3_outputs[531]) | (layer3_outputs[915]);
    assign layer4_outputs[1951] = layer3_outputs[2381];
    assign layer4_outputs[1952] = ~(layer3_outputs[1331]) | (layer3_outputs[1677]);
    assign layer4_outputs[1953] = layer3_outputs[1634];
    assign layer4_outputs[1954] = (layer3_outputs[89]) ^ (layer3_outputs[761]);
    assign layer4_outputs[1955] = ~((layer3_outputs[1644]) ^ (layer3_outputs[2248]));
    assign layer4_outputs[1956] = layer3_outputs[1549];
    assign layer4_outputs[1957] = ~((layer3_outputs[2059]) | (layer3_outputs[196]));
    assign layer4_outputs[1958] = ~(layer3_outputs[357]) | (layer3_outputs[777]);
    assign layer4_outputs[1959] = layer3_outputs[715];
    assign layer4_outputs[1960] = (layer3_outputs[308]) | (layer3_outputs[2081]);
    assign layer4_outputs[1961] = 1'b0;
    assign layer4_outputs[1962] = ~((layer3_outputs[867]) ^ (layer3_outputs[1545]));
    assign layer4_outputs[1963] = ~((layer3_outputs[1103]) | (layer3_outputs[1937]));
    assign layer4_outputs[1964] = ~((layer3_outputs[2495]) & (layer3_outputs[626]));
    assign layer4_outputs[1965] = (layer3_outputs[283]) ^ (layer3_outputs[1124]);
    assign layer4_outputs[1966] = (layer3_outputs[1366]) & ~(layer3_outputs[2365]);
    assign layer4_outputs[1967] = layer3_outputs[263];
    assign layer4_outputs[1968] = ~(layer3_outputs[982]);
    assign layer4_outputs[1969] = ~(layer3_outputs[1880]);
    assign layer4_outputs[1970] = ~(layer3_outputs[453]) | (layer3_outputs[480]);
    assign layer4_outputs[1971] = ~(layer3_outputs[2112]);
    assign layer4_outputs[1972] = ~(layer3_outputs[1823]);
    assign layer4_outputs[1973] = ~(layer3_outputs[1877]);
    assign layer4_outputs[1974] = ~(layer3_outputs[103]);
    assign layer4_outputs[1975] = (layer3_outputs[204]) ^ (layer3_outputs[1732]);
    assign layer4_outputs[1976] = layer3_outputs[1685];
    assign layer4_outputs[1977] = layer3_outputs[1114];
    assign layer4_outputs[1978] = (layer3_outputs[73]) | (layer3_outputs[1360]);
    assign layer4_outputs[1979] = (layer3_outputs[2520]) & ~(layer3_outputs[2491]);
    assign layer4_outputs[1980] = layer3_outputs[751];
    assign layer4_outputs[1981] = ~(layer3_outputs[286]);
    assign layer4_outputs[1982] = layer3_outputs[101];
    assign layer4_outputs[1983] = ~(layer3_outputs[2525]) | (layer3_outputs[1936]);
    assign layer4_outputs[1984] = (layer3_outputs[638]) ^ (layer3_outputs[598]);
    assign layer4_outputs[1985] = ~(layer3_outputs[956]) | (layer3_outputs[2371]);
    assign layer4_outputs[1986] = ~(layer3_outputs[1898]);
    assign layer4_outputs[1987] = layer3_outputs[2026];
    assign layer4_outputs[1988] = ~(layer3_outputs[599]);
    assign layer4_outputs[1989] = ~(layer3_outputs[2422]);
    assign layer4_outputs[1990] = layer3_outputs[1204];
    assign layer4_outputs[1991] = ~(layer3_outputs[855]);
    assign layer4_outputs[1992] = ~(layer3_outputs[2212]);
    assign layer4_outputs[1993] = ~(layer3_outputs[699]);
    assign layer4_outputs[1994] = ~((layer3_outputs[2091]) ^ (layer3_outputs[187]));
    assign layer4_outputs[1995] = ~((layer3_outputs[2405]) | (layer3_outputs[1261]));
    assign layer4_outputs[1996] = layer3_outputs[155];
    assign layer4_outputs[1997] = ~(layer3_outputs[1962]);
    assign layer4_outputs[1998] = ~(layer3_outputs[1133]);
    assign layer4_outputs[1999] = ~((layer3_outputs[761]) ^ (layer3_outputs[677]));
    assign layer4_outputs[2000] = (layer3_outputs[151]) ^ (layer3_outputs[602]);
    assign layer4_outputs[2001] = ~(layer3_outputs[2022]);
    assign layer4_outputs[2002] = ~(layer3_outputs[606]);
    assign layer4_outputs[2003] = ~(layer3_outputs[2338]);
    assign layer4_outputs[2004] = ~((layer3_outputs[13]) | (layer3_outputs[1093]));
    assign layer4_outputs[2005] = ~(layer3_outputs[1529]);
    assign layer4_outputs[2006] = layer3_outputs[1986];
    assign layer4_outputs[2007] = ~((layer3_outputs[946]) ^ (layer3_outputs[1046]));
    assign layer4_outputs[2008] = (layer3_outputs[1552]) & ~(layer3_outputs[194]);
    assign layer4_outputs[2009] = (layer3_outputs[1805]) & ~(layer3_outputs[2150]);
    assign layer4_outputs[2010] = ~(layer3_outputs[2495]);
    assign layer4_outputs[2011] = layer3_outputs[762];
    assign layer4_outputs[2012] = ~(layer3_outputs[1766]) | (layer3_outputs[1398]);
    assign layer4_outputs[2013] = ~(layer3_outputs[16]);
    assign layer4_outputs[2014] = layer3_outputs[715];
    assign layer4_outputs[2015] = ~(layer3_outputs[488]) | (layer3_outputs[1924]);
    assign layer4_outputs[2016] = layer3_outputs[2039];
    assign layer4_outputs[2017] = ~(layer3_outputs[2077]);
    assign layer4_outputs[2018] = ~(layer3_outputs[1134]);
    assign layer4_outputs[2019] = ~(layer3_outputs[2108]);
    assign layer4_outputs[2020] = ~((layer3_outputs[1535]) & (layer3_outputs[2061]));
    assign layer4_outputs[2021] = (layer3_outputs[1601]) & ~(layer3_outputs[1180]);
    assign layer4_outputs[2022] = layer3_outputs[1199];
    assign layer4_outputs[2023] = ~((layer3_outputs[326]) | (layer3_outputs[28]));
    assign layer4_outputs[2024] = 1'b1;
    assign layer4_outputs[2025] = layer3_outputs[829];
    assign layer4_outputs[2026] = layer3_outputs[816];
    assign layer4_outputs[2027] = ~((layer3_outputs[278]) ^ (layer3_outputs[1604]));
    assign layer4_outputs[2028] = (layer3_outputs[2115]) ^ (layer3_outputs[2341]);
    assign layer4_outputs[2029] = 1'b1;
    assign layer4_outputs[2030] = layer3_outputs[1910];
    assign layer4_outputs[2031] = ~(layer3_outputs[685]);
    assign layer4_outputs[2032] = (layer3_outputs[2062]) ^ (layer3_outputs[96]);
    assign layer4_outputs[2033] = (layer3_outputs[1290]) & (layer3_outputs[2072]);
    assign layer4_outputs[2034] = ~(layer3_outputs[688]);
    assign layer4_outputs[2035] = ~((layer3_outputs[86]) ^ (layer3_outputs[1593]));
    assign layer4_outputs[2036] = layer3_outputs[2113];
    assign layer4_outputs[2037] = ~(layer3_outputs[447]);
    assign layer4_outputs[2038] = ~((layer3_outputs[228]) | (layer3_outputs[721]));
    assign layer4_outputs[2039] = ~(layer3_outputs[18]);
    assign layer4_outputs[2040] = layer3_outputs[1202];
    assign layer4_outputs[2041] = ~(layer3_outputs[476]) | (layer3_outputs[1301]);
    assign layer4_outputs[2042] = ~(layer3_outputs[1180]);
    assign layer4_outputs[2043] = ~(layer3_outputs[473]) | (layer3_outputs[1249]);
    assign layer4_outputs[2044] = (layer3_outputs[1237]) & ~(layer3_outputs[1694]);
    assign layer4_outputs[2045] = (layer3_outputs[864]) ^ (layer3_outputs[2309]);
    assign layer4_outputs[2046] = layer3_outputs[291];
    assign layer4_outputs[2047] = layer3_outputs[1102];
    assign layer4_outputs[2048] = layer3_outputs[4];
    assign layer4_outputs[2049] = ~(layer3_outputs[472]);
    assign layer4_outputs[2050] = ~(layer3_outputs[535]);
    assign layer4_outputs[2051] = (layer3_outputs[57]) ^ (layer3_outputs[655]);
    assign layer4_outputs[2052] = ~((layer3_outputs[729]) ^ (layer3_outputs[878]));
    assign layer4_outputs[2053] = ~(layer3_outputs[1711]);
    assign layer4_outputs[2054] = ~(layer3_outputs[2317]);
    assign layer4_outputs[2055] = ~((layer3_outputs[1603]) ^ (layer3_outputs[107]));
    assign layer4_outputs[2056] = ~(layer3_outputs[2324]) | (layer3_outputs[957]);
    assign layer4_outputs[2057] = layer3_outputs[461];
    assign layer4_outputs[2058] = (layer3_outputs[1761]) & ~(layer3_outputs[2292]);
    assign layer4_outputs[2059] = ~(layer3_outputs[2428]);
    assign layer4_outputs[2060] = ~(layer3_outputs[644]);
    assign layer4_outputs[2061] = ~((layer3_outputs[1847]) | (layer3_outputs[1719]));
    assign layer4_outputs[2062] = ~((layer3_outputs[512]) ^ (layer3_outputs[2221]));
    assign layer4_outputs[2063] = layer3_outputs[301];
    assign layer4_outputs[2064] = ~(layer3_outputs[793]);
    assign layer4_outputs[2065] = layer3_outputs[1562];
    assign layer4_outputs[2066] = ~((layer3_outputs[847]) | (layer3_outputs[1668]));
    assign layer4_outputs[2067] = ~((layer3_outputs[327]) & (layer3_outputs[583]));
    assign layer4_outputs[2068] = ~(layer3_outputs[695]);
    assign layer4_outputs[2069] = (layer3_outputs[1789]) ^ (layer3_outputs[1248]);
    assign layer4_outputs[2070] = (layer3_outputs[142]) | (layer3_outputs[627]);
    assign layer4_outputs[2071] = ~(layer3_outputs[2044]) | (layer3_outputs[1991]);
    assign layer4_outputs[2072] = ~((layer3_outputs[1287]) ^ (layer3_outputs[306]));
    assign layer4_outputs[2073] = ~(layer3_outputs[303]);
    assign layer4_outputs[2074] = layer3_outputs[533];
    assign layer4_outputs[2075] = ~(layer3_outputs[658]);
    assign layer4_outputs[2076] = ~((layer3_outputs[1234]) & (layer3_outputs[373]));
    assign layer4_outputs[2077] = ~(layer3_outputs[0]) | (layer3_outputs[1656]);
    assign layer4_outputs[2078] = ~(layer3_outputs[1982]);
    assign layer4_outputs[2079] = ~(layer3_outputs[2496]) | (layer3_outputs[429]);
    assign layer4_outputs[2080] = ~(layer3_outputs[2479]);
    assign layer4_outputs[2081] = layer3_outputs[1724];
    assign layer4_outputs[2082] = layer3_outputs[2302];
    assign layer4_outputs[2083] = (layer3_outputs[88]) & ~(layer3_outputs[503]);
    assign layer4_outputs[2084] = ~(layer3_outputs[2088]);
    assign layer4_outputs[2085] = (layer3_outputs[1027]) ^ (layer3_outputs[1929]);
    assign layer4_outputs[2086] = ~(layer3_outputs[1762]);
    assign layer4_outputs[2087] = (layer3_outputs[1720]) & (layer3_outputs[2468]);
    assign layer4_outputs[2088] = ~((layer3_outputs[505]) | (layer3_outputs[618]));
    assign layer4_outputs[2089] = (layer3_outputs[2261]) & ~(layer3_outputs[1232]);
    assign layer4_outputs[2090] = ~(layer3_outputs[1849]) | (layer3_outputs[209]);
    assign layer4_outputs[2091] = ~(layer3_outputs[1391]);
    assign layer4_outputs[2092] = (layer3_outputs[1627]) & ~(layer3_outputs[1442]);
    assign layer4_outputs[2093] = ~(layer3_outputs[459]);
    assign layer4_outputs[2094] = (layer3_outputs[154]) & ~(layer3_outputs[1451]);
    assign layer4_outputs[2095] = ~(layer3_outputs[1170]);
    assign layer4_outputs[2096] = layer3_outputs[1286];
    assign layer4_outputs[2097] = (layer3_outputs[359]) & ~(layer3_outputs[1265]);
    assign layer4_outputs[2098] = layer3_outputs[1197];
    assign layer4_outputs[2099] = ~(layer3_outputs[1159]);
    assign layer4_outputs[2100] = ~((layer3_outputs[2353]) ^ (layer3_outputs[2141]));
    assign layer4_outputs[2101] = (layer3_outputs[380]) ^ (layer3_outputs[2414]);
    assign layer4_outputs[2102] = layer3_outputs[1238];
    assign layer4_outputs[2103] = 1'b0;
    assign layer4_outputs[2104] = 1'b0;
    assign layer4_outputs[2105] = ~(layer3_outputs[2559]);
    assign layer4_outputs[2106] = (layer3_outputs[1700]) ^ (layer3_outputs[1499]);
    assign layer4_outputs[2107] = ~(layer3_outputs[253]);
    assign layer4_outputs[2108] = ~(layer3_outputs[1578]);
    assign layer4_outputs[2109] = ~(layer3_outputs[991]) | (layer3_outputs[1674]);
    assign layer4_outputs[2110] = ~(layer3_outputs[2272]);
    assign layer4_outputs[2111] = ~((layer3_outputs[1811]) | (layer3_outputs[1351]));
    assign layer4_outputs[2112] = (layer3_outputs[561]) & (layer3_outputs[517]);
    assign layer4_outputs[2113] = layer3_outputs[1941];
    assign layer4_outputs[2114] = layer3_outputs[1968];
    assign layer4_outputs[2115] = (layer3_outputs[2086]) & ~(layer3_outputs[1574]);
    assign layer4_outputs[2116] = (layer3_outputs[219]) | (layer3_outputs[259]);
    assign layer4_outputs[2117] = ~(layer3_outputs[1772]) | (layer3_outputs[817]);
    assign layer4_outputs[2118] = layer3_outputs[534];
    assign layer4_outputs[2119] = (layer3_outputs[2252]) | (layer3_outputs[1764]);
    assign layer4_outputs[2120] = ~((layer3_outputs[2237]) | (layer3_outputs[1945]));
    assign layer4_outputs[2121] = layer3_outputs[2033];
    assign layer4_outputs[2122] = layer3_outputs[2080];
    assign layer4_outputs[2123] = ~(layer3_outputs[141]);
    assign layer4_outputs[2124] = layer3_outputs[1895];
    assign layer4_outputs[2125] = layer3_outputs[2243];
    assign layer4_outputs[2126] = (layer3_outputs[152]) & ~(layer3_outputs[2268]);
    assign layer4_outputs[2127] = ~((layer3_outputs[1327]) | (layer3_outputs[1960]));
    assign layer4_outputs[2128] = ~((layer3_outputs[2016]) & (layer3_outputs[37]));
    assign layer4_outputs[2129] = ~(layer3_outputs[1428]) | (layer3_outputs[1339]);
    assign layer4_outputs[2130] = ~((layer3_outputs[1887]) ^ (layer3_outputs[119]));
    assign layer4_outputs[2131] = layer3_outputs[2444];
    assign layer4_outputs[2132] = ~((layer3_outputs[2384]) ^ (layer3_outputs[477]));
    assign layer4_outputs[2133] = layer3_outputs[1355];
    assign layer4_outputs[2134] = layer3_outputs[1565];
    assign layer4_outputs[2135] = layer3_outputs[1136];
    assign layer4_outputs[2136] = (layer3_outputs[1348]) & ~(layer3_outputs[1998]);
    assign layer4_outputs[2137] = ~(layer3_outputs[465]);
    assign layer4_outputs[2138] = (layer3_outputs[191]) | (layer3_outputs[2285]);
    assign layer4_outputs[2139] = ~(layer3_outputs[1174]) | (layer3_outputs[1595]);
    assign layer4_outputs[2140] = layer3_outputs[469];
    assign layer4_outputs[2141] = layer3_outputs[2438];
    assign layer4_outputs[2142] = ~(layer3_outputs[1516]);
    assign layer4_outputs[2143] = ~(layer3_outputs[1122]);
    assign layer4_outputs[2144] = (layer3_outputs[1326]) & ~(layer3_outputs[983]);
    assign layer4_outputs[2145] = layer3_outputs[1634];
    assign layer4_outputs[2146] = ~(layer3_outputs[629]);
    assign layer4_outputs[2147] = layer3_outputs[497];
    assign layer4_outputs[2148] = ~(layer3_outputs[1101]);
    assign layer4_outputs[2149] = ~(layer3_outputs[1638]);
    assign layer4_outputs[2150] = ~(layer3_outputs[857]);
    assign layer4_outputs[2151] = ~(layer3_outputs[1302]);
    assign layer4_outputs[2152] = ~(layer3_outputs[2063]);
    assign layer4_outputs[2153] = ~(layer3_outputs[2485]);
    assign layer4_outputs[2154] = ~(layer3_outputs[1278]) | (layer3_outputs[338]);
    assign layer4_outputs[2155] = ~((layer3_outputs[1300]) ^ (layer3_outputs[2546]));
    assign layer4_outputs[2156] = ~(layer3_outputs[1961]) | (layer3_outputs[2018]);
    assign layer4_outputs[2157] = ~((layer3_outputs[218]) ^ (layer3_outputs[1206]));
    assign layer4_outputs[2158] = (layer3_outputs[1246]) & (layer3_outputs[2489]);
    assign layer4_outputs[2159] = ~(layer3_outputs[1767]) | (layer3_outputs[347]);
    assign layer4_outputs[2160] = (layer3_outputs[467]) ^ (layer3_outputs[1286]);
    assign layer4_outputs[2161] = ~(layer3_outputs[1231]);
    assign layer4_outputs[2162] = ~((layer3_outputs[2465]) & (layer3_outputs[335]));
    assign layer4_outputs[2163] = ~(layer3_outputs[2502]) | (layer3_outputs[2195]);
    assign layer4_outputs[2164] = layer3_outputs[992];
    assign layer4_outputs[2165] = ~(layer3_outputs[1182]);
    assign layer4_outputs[2166] = layer3_outputs[2037];
    assign layer4_outputs[2167] = (layer3_outputs[1336]) ^ (layer3_outputs[1042]);
    assign layer4_outputs[2168] = layer3_outputs[2227];
    assign layer4_outputs[2169] = (layer3_outputs[335]) ^ (layer3_outputs[431]);
    assign layer4_outputs[2170] = ~(layer3_outputs[1231]);
    assign layer4_outputs[2171] = layer3_outputs[1026];
    assign layer4_outputs[2172] = (layer3_outputs[922]) & ~(layer3_outputs[834]);
    assign layer4_outputs[2173] = ~(layer3_outputs[2109]);
    assign layer4_outputs[2174] = ~(layer3_outputs[176]);
    assign layer4_outputs[2175] = layer3_outputs[1683];
    assign layer4_outputs[2176] = (layer3_outputs[2085]) & ~(layer3_outputs[1305]);
    assign layer4_outputs[2177] = ~(layer3_outputs[188]);
    assign layer4_outputs[2178] = ~(layer3_outputs[454]);
    assign layer4_outputs[2179] = layer3_outputs[1934];
    assign layer4_outputs[2180] = ~((layer3_outputs[5]) & (layer3_outputs[1006]));
    assign layer4_outputs[2181] = ~(layer3_outputs[1892]);
    assign layer4_outputs[2182] = ~((layer3_outputs[1275]) | (layer3_outputs[637]));
    assign layer4_outputs[2183] = ~(layer3_outputs[1485]);
    assign layer4_outputs[2184] = ~(layer3_outputs[1297]);
    assign layer4_outputs[2185] = (layer3_outputs[1136]) ^ (layer3_outputs[211]);
    assign layer4_outputs[2186] = ~(layer3_outputs[990]) | (layer3_outputs[767]);
    assign layer4_outputs[2187] = layer3_outputs[713];
    assign layer4_outputs[2188] = ~(layer3_outputs[1904]);
    assign layer4_outputs[2189] = ~(layer3_outputs[2510]) | (layer3_outputs[1235]);
    assign layer4_outputs[2190] = ~(layer3_outputs[2506]);
    assign layer4_outputs[2191] = ~(layer3_outputs[1120]);
    assign layer4_outputs[2192] = (layer3_outputs[656]) ^ (layer3_outputs[2070]);
    assign layer4_outputs[2193] = ~(layer3_outputs[2551]) | (layer3_outputs[1701]);
    assign layer4_outputs[2194] = ~((layer3_outputs[29]) & (layer3_outputs[1624]));
    assign layer4_outputs[2195] = layer3_outputs[1522];
    assign layer4_outputs[2196] = ~((layer3_outputs[1315]) | (layer3_outputs[1015]));
    assign layer4_outputs[2197] = ~((layer3_outputs[2409]) ^ (layer3_outputs[1052]));
    assign layer4_outputs[2198] = (layer3_outputs[1913]) & ~(layer3_outputs[1575]);
    assign layer4_outputs[2199] = ~((layer3_outputs[940]) & (layer3_outputs[265]));
    assign layer4_outputs[2200] = ~(layer3_outputs[1869]) | (layer3_outputs[636]);
    assign layer4_outputs[2201] = ~((layer3_outputs[2515]) | (layer3_outputs[393]));
    assign layer4_outputs[2202] = (layer3_outputs[385]) & (layer3_outputs[1083]);
    assign layer4_outputs[2203] = ~(layer3_outputs[112]);
    assign layer4_outputs[2204] = layer3_outputs[2263];
    assign layer4_outputs[2205] = ~((layer3_outputs[87]) & (layer3_outputs[1703]));
    assign layer4_outputs[2206] = ~((layer3_outputs[1819]) | (layer3_outputs[2011]));
    assign layer4_outputs[2207] = ~((layer3_outputs[780]) | (layer3_outputs[2554]));
    assign layer4_outputs[2208] = layer3_outputs[2401];
    assign layer4_outputs[2209] = ~(layer3_outputs[2543]);
    assign layer4_outputs[2210] = ~((layer3_outputs[2112]) | (layer3_outputs[1794]));
    assign layer4_outputs[2211] = layer3_outputs[1521];
    assign layer4_outputs[2212] = (layer3_outputs[1089]) & (layer3_outputs[1938]);
    assign layer4_outputs[2213] = (layer3_outputs[1567]) & ~(layer3_outputs[708]);
    assign layer4_outputs[2214] = layer3_outputs[2199];
    assign layer4_outputs[2215] = ~(layer3_outputs[1868]);
    assign layer4_outputs[2216] = ~(layer3_outputs[2436]);
    assign layer4_outputs[2217] = (layer3_outputs[1195]) & ~(layer3_outputs[2300]);
    assign layer4_outputs[2218] = ~((layer3_outputs[614]) ^ (layer3_outputs[1387]));
    assign layer4_outputs[2219] = ~(layer3_outputs[2530]) | (layer3_outputs[2027]);
    assign layer4_outputs[2220] = layer3_outputs[116];
    assign layer4_outputs[2221] = ~(layer3_outputs[1511]);
    assign layer4_outputs[2222] = ~(layer3_outputs[1427]);
    assign layer4_outputs[2223] = ~(layer3_outputs[1683]);
    assign layer4_outputs[2224] = ~((layer3_outputs[2004]) ^ (layer3_outputs[1561]));
    assign layer4_outputs[2225] = layer3_outputs[1159];
    assign layer4_outputs[2226] = ~(layer3_outputs[1275]);
    assign layer4_outputs[2227] = ~(layer3_outputs[352]);
    assign layer4_outputs[2228] = (layer3_outputs[1558]) & ~(layer3_outputs[1258]);
    assign layer4_outputs[2229] = layer3_outputs[1827];
    assign layer4_outputs[2230] = ~((layer3_outputs[1161]) & (layer3_outputs[21]));
    assign layer4_outputs[2231] = ~(layer3_outputs[1946]);
    assign layer4_outputs[2232] = ~(layer3_outputs[742]);
    assign layer4_outputs[2233] = layer3_outputs[1372];
    assign layer4_outputs[2234] = (layer3_outputs[1016]) | (layer3_outputs[399]);
    assign layer4_outputs[2235] = layer3_outputs[2];
    assign layer4_outputs[2236] = ~((layer3_outputs[709]) & (layer3_outputs[546]));
    assign layer4_outputs[2237] = (layer3_outputs[1648]) & ~(layer3_outputs[1546]);
    assign layer4_outputs[2238] = layer3_outputs[1221];
    assign layer4_outputs[2239] = layer3_outputs[1239];
    assign layer4_outputs[2240] = ~(layer3_outputs[2363]);
    assign layer4_outputs[2241] = ~(layer3_outputs[2343]);
    assign layer4_outputs[2242] = layer3_outputs[1140];
    assign layer4_outputs[2243] = ~(layer3_outputs[121]);
    assign layer4_outputs[2244] = ~((layer3_outputs[1807]) ^ (layer3_outputs[448]));
    assign layer4_outputs[2245] = ~(layer3_outputs[2454]) | (layer3_outputs[1285]);
    assign layer4_outputs[2246] = (layer3_outputs[819]) & ~(layer3_outputs[689]);
    assign layer4_outputs[2247] = ~(layer3_outputs[988]);
    assign layer4_outputs[2248] = ~(layer3_outputs[602]);
    assign layer4_outputs[2249] = ~(layer3_outputs[1524]);
    assign layer4_outputs[2250] = layer3_outputs[1417];
    assign layer4_outputs[2251] = ~(layer3_outputs[1537]) | (layer3_outputs[1791]);
    assign layer4_outputs[2252] = ~(layer3_outputs[437]) | (layer3_outputs[909]);
    assign layer4_outputs[2253] = ~(layer3_outputs[1585]);
    assign layer4_outputs[2254] = (layer3_outputs[2047]) & ~(layer3_outputs[845]);
    assign layer4_outputs[2255] = ~(layer3_outputs[770]);
    assign layer4_outputs[2256] = ~((layer3_outputs[1394]) | (layer3_outputs[1272]));
    assign layer4_outputs[2257] = layer3_outputs[1986];
    assign layer4_outputs[2258] = (layer3_outputs[604]) ^ (layer3_outputs[743]);
    assign layer4_outputs[2259] = ~(layer3_outputs[959]);
    assign layer4_outputs[2260] = ~(layer3_outputs[1004]);
    assign layer4_outputs[2261] = ~((layer3_outputs[2210]) ^ (layer3_outputs[2424]));
    assign layer4_outputs[2262] = ~(layer3_outputs[1706]);
    assign layer4_outputs[2263] = layer3_outputs[1598];
    assign layer4_outputs[2264] = ~((layer3_outputs[1876]) & (layer3_outputs[374]));
    assign layer4_outputs[2265] = layer3_outputs[2283];
    assign layer4_outputs[2266] = ~(layer3_outputs[2243]);
    assign layer4_outputs[2267] = layer3_outputs[159];
    assign layer4_outputs[2268] = ~(layer3_outputs[2451]);
    assign layer4_outputs[2269] = ~(layer3_outputs[1240]);
    assign layer4_outputs[2270] = layer3_outputs[2369];
    assign layer4_outputs[2271] = ~(layer3_outputs[1047]);
    assign layer4_outputs[2272] = (layer3_outputs[1013]) & ~(layer3_outputs[904]);
    assign layer4_outputs[2273] = ~(layer3_outputs[2176]);
    assign layer4_outputs[2274] = layer3_outputs[2389];
    assign layer4_outputs[2275] = layer3_outputs[1994];
    assign layer4_outputs[2276] = layer3_outputs[1675];
    assign layer4_outputs[2277] = 1'b0;
    assign layer4_outputs[2278] = layer3_outputs[1946];
    assign layer4_outputs[2279] = layer3_outputs[2235];
    assign layer4_outputs[2280] = ~(layer3_outputs[573]);
    assign layer4_outputs[2281] = ~(layer3_outputs[2060]) | (layer3_outputs[2146]);
    assign layer4_outputs[2282] = ~((layer3_outputs[1440]) ^ (layer3_outputs[2023]));
    assign layer4_outputs[2283] = layer3_outputs[645];
    assign layer4_outputs[2284] = layer3_outputs[2115];
    assign layer4_outputs[2285] = layer3_outputs[2435];
    assign layer4_outputs[2286] = ~(layer3_outputs[1299]);
    assign layer4_outputs[2287] = ~(layer3_outputs[2325]);
    assign layer4_outputs[2288] = ~((layer3_outputs[1658]) | (layer3_outputs[262]));
    assign layer4_outputs[2289] = layer3_outputs[1547];
    assign layer4_outputs[2290] = (layer3_outputs[501]) & ~(layer3_outputs[1320]);
    assign layer4_outputs[2291] = ~((layer3_outputs[1150]) ^ (layer3_outputs[2185]));
    assign layer4_outputs[2292] = ~(layer3_outputs[2222]);
    assign layer4_outputs[2293] = ~((layer3_outputs[1370]) ^ (layer3_outputs[1113]));
    assign layer4_outputs[2294] = ~(layer3_outputs[1412]);
    assign layer4_outputs[2295] = (layer3_outputs[2264]) & ~(layer3_outputs[1939]);
    assign layer4_outputs[2296] = ~(layer3_outputs[1343]);
    assign layer4_outputs[2297] = (layer3_outputs[867]) ^ (layer3_outputs[821]);
    assign layer4_outputs[2298] = (layer3_outputs[2100]) & ~(layer3_outputs[760]);
    assign layer4_outputs[2299] = ~((layer3_outputs[1618]) ^ (layer3_outputs[712]));
    assign layer4_outputs[2300] = ~(layer3_outputs[164]);
    assign layer4_outputs[2301] = 1'b0;
    assign layer4_outputs[2302] = layer3_outputs[1245];
    assign layer4_outputs[2303] = ~(layer3_outputs[250]);
    assign layer4_outputs[2304] = layer3_outputs[1335];
    assign layer4_outputs[2305] = ~((layer3_outputs[1577]) & (layer3_outputs[1835]));
    assign layer4_outputs[2306] = (layer3_outputs[2038]) & ~(layer3_outputs[1965]);
    assign layer4_outputs[2307] = ~((layer3_outputs[1673]) ^ (layer3_outputs[1478]));
    assign layer4_outputs[2308] = (layer3_outputs[1242]) | (layer3_outputs[1247]);
    assign layer4_outputs[2309] = layer3_outputs[2368];
    assign layer4_outputs[2310] = layer3_outputs[720];
    assign layer4_outputs[2311] = layer3_outputs[44];
    assign layer4_outputs[2312] = ~(layer3_outputs[68]);
    assign layer4_outputs[2313] = ~((layer3_outputs[1056]) | (layer3_outputs[2413]));
    assign layer4_outputs[2314] = (layer3_outputs[2510]) & (layer3_outputs[1914]);
    assign layer4_outputs[2315] = ~(layer3_outputs[1974]);
    assign layer4_outputs[2316] = layer3_outputs[1678];
    assign layer4_outputs[2317] = ~((layer3_outputs[1253]) | (layer3_outputs[397]));
    assign layer4_outputs[2318] = ~((layer3_outputs[1279]) ^ (layer3_outputs[1137]));
    assign layer4_outputs[2319] = layer3_outputs[2527];
    assign layer4_outputs[2320] = ~((layer3_outputs[753]) ^ (layer3_outputs[1633]));
    assign layer4_outputs[2321] = (layer3_outputs[437]) & ~(layer3_outputs[2355]);
    assign layer4_outputs[2322] = ~((layer3_outputs[853]) ^ (layer3_outputs[2169]));
    assign layer4_outputs[2323] = layer3_outputs[462];
    assign layer4_outputs[2324] = ~(layer3_outputs[622]);
    assign layer4_outputs[2325] = ~(layer3_outputs[1995]);
    assign layer4_outputs[2326] = (layer3_outputs[132]) & (layer3_outputs[173]);
    assign layer4_outputs[2327] = ~((layer3_outputs[1525]) & (layer3_outputs[887]));
    assign layer4_outputs[2328] = layer3_outputs[1805];
    assign layer4_outputs[2329] = layer3_outputs[462];
    assign layer4_outputs[2330] = ~(layer3_outputs[1374]);
    assign layer4_outputs[2331] = layer3_outputs[1250];
    assign layer4_outputs[2332] = layer3_outputs[2260];
    assign layer4_outputs[2333] = ~(layer3_outputs[1682]) | (layer3_outputs[2412]);
    assign layer4_outputs[2334] = layer3_outputs[1019];
    assign layer4_outputs[2335] = layer3_outputs[1768];
    assign layer4_outputs[2336] = (layer3_outputs[319]) ^ (layer3_outputs[2254]);
    assign layer4_outputs[2337] = (layer3_outputs[1916]) & (layer3_outputs[2240]);
    assign layer4_outputs[2338] = (layer3_outputs[1045]) & ~(layer3_outputs[1293]);
    assign layer4_outputs[2339] = ~(layer3_outputs[2469]);
    assign layer4_outputs[2340] = ~(layer3_outputs[1339]);
    assign layer4_outputs[2341] = (layer3_outputs[2501]) | (layer3_outputs[1081]);
    assign layer4_outputs[2342] = ~(layer3_outputs[1640]);
    assign layer4_outputs[2343] = (layer3_outputs[1255]) ^ (layer3_outputs[2415]);
    assign layer4_outputs[2344] = (layer3_outputs[651]) ^ (layer3_outputs[1809]);
    assign layer4_outputs[2345] = ~(layer3_outputs[601]);
    assign layer4_outputs[2346] = ~(layer3_outputs[427]);
    assign layer4_outputs[2347] = ~(layer3_outputs[956]);
    assign layer4_outputs[2348] = ~(layer3_outputs[2188]);
    assign layer4_outputs[2349] = ~(layer3_outputs[1848]) | (layer3_outputs[1042]);
    assign layer4_outputs[2350] = ~(layer3_outputs[1353]);
    assign layer4_outputs[2351] = layer3_outputs[2322];
    assign layer4_outputs[2352] = (layer3_outputs[1377]) | (layer3_outputs[1453]);
    assign layer4_outputs[2353] = ~((layer3_outputs[2011]) ^ (layer3_outputs[1390]));
    assign layer4_outputs[2354] = ~((layer3_outputs[205]) ^ (layer3_outputs[1832]));
    assign layer4_outputs[2355] = layer3_outputs[246];
    assign layer4_outputs[2356] = ~((layer3_outputs[1465]) | (layer3_outputs[310]));
    assign layer4_outputs[2357] = ~(layer3_outputs[2137]) | (layer3_outputs[1303]);
    assign layer4_outputs[2358] = ~((layer3_outputs[137]) & (layer3_outputs[1359]));
    assign layer4_outputs[2359] = ~(layer3_outputs[1496]);
    assign layer4_outputs[2360] = ~(layer3_outputs[1838]);
    assign layer4_outputs[2361] = ~((layer3_outputs[1483]) & (layer3_outputs[309]));
    assign layer4_outputs[2362] = (layer3_outputs[2129]) & ~(layer3_outputs[2268]);
    assign layer4_outputs[2363] = ~((layer3_outputs[2002]) ^ (layer3_outputs[555]));
    assign layer4_outputs[2364] = ~(layer3_outputs[738]);
    assign layer4_outputs[2365] = layer3_outputs[1229];
    assign layer4_outputs[2366] = ~((layer3_outputs[1164]) & (layer3_outputs[419]));
    assign layer4_outputs[2367] = ~(layer3_outputs[1626]);
    assign layer4_outputs[2368] = layer3_outputs[930];
    assign layer4_outputs[2369] = layer3_outputs[2130];
    assign layer4_outputs[2370] = ~((layer3_outputs[1188]) | (layer3_outputs[264]));
    assign layer4_outputs[2371] = layer3_outputs[2532];
    assign layer4_outputs[2372] = (layer3_outputs[2228]) & ~(layer3_outputs[266]);
    assign layer4_outputs[2373] = ~(layer3_outputs[361]);
    assign layer4_outputs[2374] = ~(layer3_outputs[2139]);
    assign layer4_outputs[2375] = ~(layer3_outputs[2484]) | (layer3_outputs[873]);
    assign layer4_outputs[2376] = (layer3_outputs[1443]) & ~(layer3_outputs[1108]);
    assign layer4_outputs[2377] = ~(layer3_outputs[2122]);
    assign layer4_outputs[2378] = ~(layer3_outputs[1838]);
    assign layer4_outputs[2379] = ~(layer3_outputs[852]);
    assign layer4_outputs[2380] = ~(layer3_outputs[2189]);
    assign layer4_outputs[2381] = (layer3_outputs[1183]) ^ (layer3_outputs[2535]);
    assign layer4_outputs[2382] = ~(layer3_outputs[2377]) | (layer3_outputs[1196]);
    assign layer4_outputs[2383] = (layer3_outputs[426]) & ~(layer3_outputs[723]);
    assign layer4_outputs[2384] = (layer3_outputs[2181]) & ~(layer3_outputs[2226]);
    assign layer4_outputs[2385] = ~(layer3_outputs[64]) | (layer3_outputs[817]);
    assign layer4_outputs[2386] = layer3_outputs[704];
    assign layer4_outputs[2387] = ~(layer3_outputs[687]) | (layer3_outputs[2516]);
    assign layer4_outputs[2388] = ~(layer3_outputs[312]);
    assign layer4_outputs[2389] = layer3_outputs[885];
    assign layer4_outputs[2390] = layer3_outputs[345];
    assign layer4_outputs[2391] = ~((layer3_outputs[2132]) ^ (layer3_outputs[1088]));
    assign layer4_outputs[2392] = ~(layer3_outputs[2377]);
    assign layer4_outputs[2393] = layer3_outputs[1658];
    assign layer4_outputs[2394] = ~(layer3_outputs[623]);
    assign layer4_outputs[2395] = ~(layer3_outputs[1945]);
    assign layer4_outputs[2396] = layer3_outputs[1393];
    assign layer4_outputs[2397] = ~((layer3_outputs[2439]) & (layer3_outputs[1463]));
    assign layer4_outputs[2398] = ~((layer3_outputs[1163]) ^ (layer3_outputs[763]));
    assign layer4_outputs[2399] = (layer3_outputs[1712]) | (layer3_outputs[1192]);
    assign layer4_outputs[2400] = (layer3_outputs[1403]) & ~(layer3_outputs[422]);
    assign layer4_outputs[2401] = ~((layer3_outputs[2052]) | (layer3_outputs[2352]));
    assign layer4_outputs[2402] = ~(layer3_outputs[1536]);
    assign layer4_outputs[2403] = ~(layer3_outputs[1300]) | (layer3_outputs[1901]);
    assign layer4_outputs[2404] = layer3_outputs[1957];
    assign layer4_outputs[2405] = ~(layer3_outputs[1766]);
    assign layer4_outputs[2406] = ~((layer3_outputs[1713]) & (layer3_outputs[1250]));
    assign layer4_outputs[2407] = ~(layer3_outputs[1130]) | (layer3_outputs[1211]);
    assign layer4_outputs[2408] = ~(layer3_outputs[1750]);
    assign layer4_outputs[2409] = ~(layer3_outputs[1452]) | (layer3_outputs[2293]);
    assign layer4_outputs[2410] = layer3_outputs[2430];
    assign layer4_outputs[2411] = ~(layer3_outputs[1995]);
    assign layer4_outputs[2412] = ~(layer3_outputs[155]) | (layer3_outputs[563]);
    assign layer4_outputs[2413] = ~((layer3_outputs[2540]) ^ (layer3_outputs[105]));
    assign layer4_outputs[2414] = ~(layer3_outputs[1750]);
    assign layer4_outputs[2415] = layer3_outputs[759];
    assign layer4_outputs[2416] = ~((layer3_outputs[2516]) & (layer3_outputs[403]));
    assign layer4_outputs[2417] = ~(layer3_outputs[1351]);
    assign layer4_outputs[2418] = layer3_outputs[1212];
    assign layer4_outputs[2419] = layer3_outputs[2012];
    assign layer4_outputs[2420] = ~(layer3_outputs[771]);
    assign layer4_outputs[2421] = ~((layer3_outputs[1627]) ^ (layer3_outputs[434]));
    assign layer4_outputs[2422] = (layer3_outputs[755]) & ~(layer3_outputs[2194]);
    assign layer4_outputs[2423] = ~(layer3_outputs[2283]);
    assign layer4_outputs[2424] = (layer3_outputs[1343]) & ~(layer3_outputs[9]);
    assign layer4_outputs[2425] = ~(layer3_outputs[2544]);
    assign layer4_outputs[2426] = ~(layer3_outputs[537]);
    assign layer4_outputs[2427] = ~((layer3_outputs[947]) | (layer3_outputs[657]));
    assign layer4_outputs[2428] = ~(layer3_outputs[2123]);
    assign layer4_outputs[2429] = (layer3_outputs[497]) ^ (layer3_outputs[2232]);
    assign layer4_outputs[2430] = layer3_outputs[1052];
    assign layer4_outputs[2431] = layer3_outputs[1498];
    assign layer4_outputs[2432] = (layer3_outputs[273]) & (layer3_outputs[709]);
    assign layer4_outputs[2433] = ~(layer3_outputs[325]);
    assign layer4_outputs[2434] = (layer3_outputs[823]) ^ (layer3_outputs[868]);
    assign layer4_outputs[2435] = ~((layer3_outputs[113]) ^ (layer3_outputs[446]));
    assign layer4_outputs[2436] = ~((layer3_outputs[2200]) & (layer3_outputs[1434]));
    assign layer4_outputs[2437] = (layer3_outputs[559]) ^ (layer3_outputs[128]);
    assign layer4_outputs[2438] = ~(layer3_outputs[1689]) | (layer3_outputs[162]);
    assign layer4_outputs[2439] = layer3_outputs[1429];
    assign layer4_outputs[2440] = ~(layer3_outputs[1121]) | (layer3_outputs[1503]);
    assign layer4_outputs[2441] = ~(layer3_outputs[1432]) | (layer3_outputs[1100]);
    assign layer4_outputs[2442] = ~(layer3_outputs[174]) | (layer3_outputs[2354]);
    assign layer4_outputs[2443] = (layer3_outputs[1079]) ^ (layer3_outputs[383]);
    assign layer4_outputs[2444] = layer3_outputs[2186];
    assign layer4_outputs[2445] = ~((layer3_outputs[1458]) | (layer3_outputs[188]));
    assign layer4_outputs[2446] = ~((layer3_outputs[1951]) & (layer3_outputs[1085]));
    assign layer4_outputs[2447] = ~(layer3_outputs[316]);
    assign layer4_outputs[2448] = (layer3_outputs[797]) & (layer3_outputs[2434]);
    assign layer4_outputs[2449] = ~(layer3_outputs[2394]) | (layer3_outputs[230]);
    assign layer4_outputs[2450] = ~((layer3_outputs[2256]) ^ (layer3_outputs[278]));
    assign layer4_outputs[2451] = ~(layer3_outputs[1881]);
    assign layer4_outputs[2452] = ~(layer3_outputs[850]);
    assign layer4_outputs[2453] = (layer3_outputs[1145]) & ~(layer3_outputs[2277]);
    assign layer4_outputs[2454] = ~(layer3_outputs[567]);
    assign layer4_outputs[2455] = ~(layer3_outputs[1306]) | (layer3_outputs[1870]);
    assign layer4_outputs[2456] = layer3_outputs[546];
    assign layer4_outputs[2457] = (layer3_outputs[1557]) & ~(layer3_outputs[730]);
    assign layer4_outputs[2458] = ~(layer3_outputs[1298]);
    assign layer4_outputs[2459] = layer3_outputs[1669];
    assign layer4_outputs[2460] = layer3_outputs[1644];
    assign layer4_outputs[2461] = ~(layer3_outputs[118]);
    assign layer4_outputs[2462] = ~((layer3_outputs[1399]) | (layer3_outputs[2444]));
    assign layer4_outputs[2463] = ~((layer3_outputs[706]) | (layer3_outputs[1740]));
    assign layer4_outputs[2464] = ~(layer3_outputs[1734]);
    assign layer4_outputs[2465] = ~((layer3_outputs[2376]) ^ (layer3_outputs[1507]));
    assign layer4_outputs[2466] = ~((layer3_outputs[1751]) & (layer3_outputs[2405]));
    assign layer4_outputs[2467] = (layer3_outputs[752]) | (layer3_outputs[272]);
    assign layer4_outputs[2468] = 1'b1;
    assign layer4_outputs[2469] = layer3_outputs[1021];
    assign layer4_outputs[2470] = ~(layer3_outputs[2212]);
    assign layer4_outputs[2471] = ~(layer3_outputs[1224]);
    assign layer4_outputs[2472] = ~(layer3_outputs[1916]);
    assign layer4_outputs[2473] = ~(layer3_outputs[2203]);
    assign layer4_outputs[2474] = (layer3_outputs[503]) & ~(layer3_outputs[1217]);
    assign layer4_outputs[2475] = layer3_outputs[1237];
    assign layer4_outputs[2476] = ~(layer3_outputs[343]) | (layer3_outputs[1629]);
    assign layer4_outputs[2477] = ~(layer3_outputs[1757]);
    assign layer4_outputs[2478] = layer3_outputs[180];
    assign layer4_outputs[2479] = (layer3_outputs[355]) | (layer3_outputs[1210]);
    assign layer4_outputs[2480] = layer3_outputs[2182];
    assign layer4_outputs[2481] = 1'b0;
    assign layer4_outputs[2482] = layer3_outputs[1837];
    assign layer4_outputs[2483] = ~(layer3_outputs[799]);
    assign layer4_outputs[2484] = ~(layer3_outputs[1053]) | (layer3_outputs[893]);
    assign layer4_outputs[2485] = ~(layer3_outputs[717]);
    assign layer4_outputs[2486] = layer3_outputs[2111];
    assign layer4_outputs[2487] = layer3_outputs[238];
    assign layer4_outputs[2488] = ~(layer3_outputs[610]) | (layer3_outputs[888]);
    assign layer4_outputs[2489] = layer3_outputs[508];
    assign layer4_outputs[2490] = ~(layer3_outputs[2508]);
    assign layer4_outputs[2491] = ~(layer3_outputs[2395]);
    assign layer4_outputs[2492] = ~(layer3_outputs[914]);
    assign layer4_outputs[2493] = ~((layer3_outputs[212]) ^ (layer3_outputs[511]));
    assign layer4_outputs[2494] = ~(layer3_outputs[102]) | (layer3_outputs[1505]);
    assign layer4_outputs[2495] = (layer3_outputs[645]) ^ (layer3_outputs[1140]);
    assign layer4_outputs[2496] = ~(layer3_outputs[1841]);
    assign layer4_outputs[2497] = layer3_outputs[1341];
    assign layer4_outputs[2498] = layer3_outputs[1567];
    assign layer4_outputs[2499] = (layer3_outputs[1653]) & ~(layer3_outputs[2349]);
    assign layer4_outputs[2500] = ~(layer3_outputs[1468]) | (layer3_outputs[381]);
    assign layer4_outputs[2501] = ~((layer3_outputs[712]) | (layer3_outputs[2222]));
    assign layer4_outputs[2502] = layer3_outputs[1084];
    assign layer4_outputs[2503] = layer3_outputs[1929];
    assign layer4_outputs[2504] = ~(layer3_outputs[2549]) | (layer3_outputs[390]);
    assign layer4_outputs[2505] = ~(layer3_outputs[67]);
    assign layer4_outputs[2506] = layer3_outputs[95];
    assign layer4_outputs[2507] = ~(layer3_outputs[1932]);
    assign layer4_outputs[2508] = 1'b1;
    assign layer4_outputs[2509] = ~((layer3_outputs[227]) & (layer3_outputs[2091]));
    assign layer4_outputs[2510] = ~(layer3_outputs[369]) | (layer3_outputs[1037]);
    assign layer4_outputs[2511] = ~(layer3_outputs[337]);
    assign layer4_outputs[2512] = (layer3_outputs[644]) & ~(layer3_outputs[921]);
    assign layer4_outputs[2513] = ~(layer3_outputs[1379]);
    assign layer4_outputs[2514] = layer3_outputs[1638];
    assign layer4_outputs[2515] = ~(layer3_outputs[1663]);
    assign layer4_outputs[2516] = (layer3_outputs[984]) ^ (layer3_outputs[1889]);
    assign layer4_outputs[2517] = ~(layer3_outputs[1061]);
    assign layer4_outputs[2518] = (layer3_outputs[1401]) ^ (layer3_outputs[1950]);
    assign layer4_outputs[2519] = ~(layer3_outputs[532]);
    assign layer4_outputs[2520] = ~((layer3_outputs[388]) | (layer3_outputs[2152]));
    assign layer4_outputs[2521] = ~(layer3_outputs[2535]);
    assign layer4_outputs[2522] = layer3_outputs[2104];
    assign layer4_outputs[2523] = layer3_outputs[266];
    assign layer4_outputs[2524] = ~(layer3_outputs[782]);
    assign layer4_outputs[2525] = layer3_outputs[2064];
    assign layer4_outputs[2526] = (layer3_outputs[1599]) ^ (layer3_outputs[240]);
    assign layer4_outputs[2527] = layer3_outputs[2120];
    assign layer4_outputs[2528] = (layer3_outputs[1469]) & ~(layer3_outputs[1704]);
    assign layer4_outputs[2529] = (layer3_outputs[2445]) & ~(layer3_outputs[106]);
    assign layer4_outputs[2530] = 1'b1;
    assign layer4_outputs[2531] = (layer3_outputs[490]) & ~(layer3_outputs[1483]);
    assign layer4_outputs[2532] = (layer3_outputs[2524]) & ~(layer3_outputs[800]);
    assign layer4_outputs[2533] = ~(layer3_outputs[907]);
    assign layer4_outputs[2534] = ~(layer3_outputs[315]);
    assign layer4_outputs[2535] = (layer3_outputs[416]) & ~(layer3_outputs[1458]);
    assign layer4_outputs[2536] = ~(layer3_outputs[809]);
    assign layer4_outputs[2537] = layer3_outputs[217];
    assign layer4_outputs[2538] = ~(layer3_outputs[575]);
    assign layer4_outputs[2539] = layer3_outputs[103];
    assign layer4_outputs[2540] = ~(layer3_outputs[8]);
    assign layer4_outputs[2541] = ~(layer3_outputs[2116]);
    assign layer4_outputs[2542] = 1'b0;
    assign layer4_outputs[2543] = (layer3_outputs[1514]) ^ (layer3_outputs[1677]);
    assign layer4_outputs[2544] = ~(layer3_outputs[2536]);
    assign layer4_outputs[2545] = ~(layer3_outputs[849]);
    assign layer4_outputs[2546] = ~(layer3_outputs[1846]);
    assign layer4_outputs[2547] = layer3_outputs[2284];
    assign layer4_outputs[2548] = ~((layer3_outputs[1955]) & (layer3_outputs[1850]));
    assign layer4_outputs[2549] = 1'b0;
    assign layer4_outputs[2550] = (layer3_outputs[131]) ^ (layer3_outputs[658]);
    assign layer4_outputs[2551] = (layer3_outputs[1606]) & ~(layer3_outputs[622]);
    assign layer4_outputs[2552] = (layer3_outputs[132]) ^ (layer3_outputs[1420]);
    assign layer4_outputs[2553] = ~(layer3_outputs[1594]);
    assign layer4_outputs[2554] = ~(layer3_outputs[2287]);
    assign layer4_outputs[2555] = ~(layer3_outputs[2117]);
    assign layer4_outputs[2556] = ~((layer3_outputs[2000]) | (layer3_outputs[818]));
    assign layer4_outputs[2557] = ~(layer3_outputs[109]);
    assign layer4_outputs[2558] = layer3_outputs[2208];
    assign layer4_outputs[2559] = ~((layer3_outputs[599]) & (layer3_outputs[2095]));
    assign outputs[0] = ~(layer4_outputs[2425]);
    assign outputs[1] = ~(layer4_outputs[1789]);
    assign outputs[2] = ~(layer4_outputs[2262]);
    assign outputs[3] = layer4_outputs[1411];
    assign outputs[4] = ~(layer4_outputs[2272]);
    assign outputs[5] = ~(layer4_outputs[623]);
    assign outputs[6] = (layer4_outputs[1139]) ^ (layer4_outputs[1025]);
    assign outputs[7] = layer4_outputs[488];
    assign outputs[8] = (layer4_outputs[652]) & (layer4_outputs[504]);
    assign outputs[9] = ~(layer4_outputs[600]);
    assign outputs[10] = ~(layer4_outputs[2093]);
    assign outputs[11] = ~(layer4_outputs[1307]);
    assign outputs[12] = ~(layer4_outputs[1568]);
    assign outputs[13] = ~(layer4_outputs[1545]);
    assign outputs[14] = ~(layer4_outputs[819]);
    assign outputs[15] = ~(layer4_outputs[1142]);
    assign outputs[16] = (layer4_outputs[2104]) ^ (layer4_outputs[1481]);
    assign outputs[17] = layer4_outputs[1328];
    assign outputs[18] = (layer4_outputs[2423]) & ~(layer4_outputs[600]);
    assign outputs[19] = layer4_outputs[963];
    assign outputs[20] = ~(layer4_outputs[859]);
    assign outputs[21] = layer4_outputs[125];
    assign outputs[22] = layer4_outputs[2537];
    assign outputs[23] = ~(layer4_outputs[1378]);
    assign outputs[24] = (layer4_outputs[761]) & ~(layer4_outputs[2060]);
    assign outputs[25] = (layer4_outputs[1992]) & ~(layer4_outputs[2388]);
    assign outputs[26] = (layer4_outputs[2490]) & (layer4_outputs[1699]);
    assign outputs[27] = ~(layer4_outputs[2139]);
    assign outputs[28] = layer4_outputs[2358];
    assign outputs[29] = (layer4_outputs[122]) & ~(layer4_outputs[2500]);
    assign outputs[30] = ~(layer4_outputs[2416]);
    assign outputs[31] = layer4_outputs[1515];
    assign outputs[32] = layer4_outputs[24];
    assign outputs[33] = ~(layer4_outputs[846]);
    assign outputs[34] = ~(layer4_outputs[1098]);
    assign outputs[35] = ~(layer4_outputs[2336]);
    assign outputs[36] = ~(layer4_outputs[1718]);
    assign outputs[37] = ~(layer4_outputs[1950]);
    assign outputs[38] = layer4_outputs[1129];
    assign outputs[39] = ~(layer4_outputs[631]);
    assign outputs[40] = layer4_outputs[1109];
    assign outputs[41] = (layer4_outputs[2144]) | (layer4_outputs[519]);
    assign outputs[42] = ~((layer4_outputs[1019]) | (layer4_outputs[2185]));
    assign outputs[43] = ~(layer4_outputs[1942]);
    assign outputs[44] = layer4_outputs[1067];
    assign outputs[45] = layer4_outputs[1459];
    assign outputs[46] = layer4_outputs[2452];
    assign outputs[47] = ~(layer4_outputs[2480]);
    assign outputs[48] = ~(layer4_outputs[2260]);
    assign outputs[49] = ~(layer4_outputs[134]);
    assign outputs[50] = (layer4_outputs[302]) & ~(layer4_outputs[223]);
    assign outputs[51] = layer4_outputs[2298];
    assign outputs[52] = (layer4_outputs[282]) & ~(layer4_outputs[462]);
    assign outputs[53] = ~(layer4_outputs[2244]);
    assign outputs[54] = layer4_outputs[1330];
    assign outputs[55] = ~(layer4_outputs[2328]);
    assign outputs[56] = (layer4_outputs[2287]) & ~(layer4_outputs[720]);
    assign outputs[57] = ~(layer4_outputs[1150]);
    assign outputs[58] = ~(layer4_outputs[2484]);
    assign outputs[59] = ~(layer4_outputs[857]);
    assign outputs[60] = layer4_outputs[1816];
    assign outputs[61] = (layer4_outputs[841]) & ~(layer4_outputs[2324]);
    assign outputs[62] = ~(layer4_outputs[431]);
    assign outputs[63] = ~(layer4_outputs[1739]);
    assign outputs[64] = (layer4_outputs[57]) & ~(layer4_outputs[1068]);
    assign outputs[65] = layer4_outputs[1914];
    assign outputs[66] = layer4_outputs[787];
    assign outputs[67] = ~(layer4_outputs[2477]) | (layer4_outputs[1827]);
    assign outputs[68] = layer4_outputs[254];
    assign outputs[69] = ~(layer4_outputs[2395]);
    assign outputs[70] = ~(layer4_outputs[2063]);
    assign outputs[71] = ~(layer4_outputs[1765]);
    assign outputs[72] = (layer4_outputs[521]) & (layer4_outputs[2250]);
    assign outputs[73] = ~((layer4_outputs[347]) ^ (layer4_outputs[852]));
    assign outputs[74] = ~(layer4_outputs[1032]);
    assign outputs[75] = (layer4_outputs[115]) & (layer4_outputs[1092]);
    assign outputs[76] = ~(layer4_outputs[2369]);
    assign outputs[77] = (layer4_outputs[214]) ^ (layer4_outputs[372]);
    assign outputs[78] = (layer4_outputs[617]) & (layer4_outputs[1559]);
    assign outputs[79] = ~(layer4_outputs[49]);
    assign outputs[80] = ~(layer4_outputs[1316]);
    assign outputs[81] = ~(layer4_outputs[651]);
    assign outputs[82] = ~(layer4_outputs[1218]);
    assign outputs[83] = ~(layer4_outputs[1101]);
    assign outputs[84] = layer4_outputs[2271];
    assign outputs[85] = (layer4_outputs[1870]) & (layer4_outputs[2097]);
    assign outputs[86] = ~((layer4_outputs[590]) | (layer4_outputs[1426]));
    assign outputs[87] = (layer4_outputs[551]) ^ (layer4_outputs[1995]);
    assign outputs[88] = ~(layer4_outputs[390]);
    assign outputs[89] = (layer4_outputs[1644]) & (layer4_outputs[2090]);
    assign outputs[90] = (layer4_outputs[1532]) & ~(layer4_outputs[1289]);
    assign outputs[91] = ~(layer4_outputs[2038]);
    assign outputs[92] = layer4_outputs[1472];
    assign outputs[93] = ~(layer4_outputs[90]);
    assign outputs[94] = layer4_outputs[866];
    assign outputs[95] = (layer4_outputs[2456]) & (layer4_outputs[1402]);
    assign outputs[96] = ~((layer4_outputs[823]) ^ (layer4_outputs[1899]));
    assign outputs[97] = ~(layer4_outputs[818]);
    assign outputs[98] = ~(layer4_outputs[359]) | (layer4_outputs[975]);
    assign outputs[99] = layer4_outputs[2261];
    assign outputs[100] = ~(layer4_outputs[1000]);
    assign outputs[101] = ~(layer4_outputs[1729]);
    assign outputs[102] = layer4_outputs[1026];
    assign outputs[103] = layer4_outputs[1600];
    assign outputs[104] = (layer4_outputs[2138]) & (layer4_outputs[240]);
    assign outputs[105] = ~(layer4_outputs[1555]);
    assign outputs[106] = ~((layer4_outputs[2244]) ^ (layer4_outputs[1688]));
    assign outputs[107] = ~(layer4_outputs[311]);
    assign outputs[108] = ~(layer4_outputs[2032]);
    assign outputs[109] = ~(layer4_outputs[1978]);
    assign outputs[110] = (layer4_outputs[1026]) & ~(layer4_outputs[1627]);
    assign outputs[111] = ~(layer4_outputs[1772]);
    assign outputs[112] = layer4_outputs[521];
    assign outputs[113] = ~((layer4_outputs[2447]) | (layer4_outputs[2551]));
    assign outputs[114] = (layer4_outputs[1418]) ^ (layer4_outputs[379]);
    assign outputs[115] = ~((layer4_outputs[953]) ^ (layer4_outputs[103]));
    assign outputs[116] = ~(layer4_outputs[1592]);
    assign outputs[117] = layer4_outputs[665];
    assign outputs[118] = ~(layer4_outputs[2434]);
    assign outputs[119] = ~(layer4_outputs[556]);
    assign outputs[120] = layer4_outputs[1182];
    assign outputs[121] = layer4_outputs[480];
    assign outputs[122] = ~(layer4_outputs[51]) | (layer4_outputs[872]);
    assign outputs[123] = layer4_outputs[225];
    assign outputs[124] = (layer4_outputs[145]) | (layer4_outputs[1510]);
    assign outputs[125] = layer4_outputs[1212];
    assign outputs[126] = layer4_outputs[1118];
    assign outputs[127] = layer4_outputs[211];
    assign outputs[128] = (layer4_outputs[1989]) ^ (layer4_outputs[2292]);
    assign outputs[129] = (layer4_outputs[2200]) & ~(layer4_outputs[1761]);
    assign outputs[130] = layer4_outputs[766];
    assign outputs[131] = ~((layer4_outputs[1784]) | (layer4_outputs[1289]));
    assign outputs[132] = ~(layer4_outputs[811]);
    assign outputs[133] = (layer4_outputs[1293]) & ~(layer4_outputs[1458]);
    assign outputs[134] = layer4_outputs[1096];
    assign outputs[135] = layer4_outputs[773];
    assign outputs[136] = ~(layer4_outputs[2165]);
    assign outputs[137] = layer4_outputs[653];
    assign outputs[138] = (layer4_outputs[57]) ^ (layer4_outputs[450]);
    assign outputs[139] = layer4_outputs[1854];
    assign outputs[140] = layer4_outputs[1655];
    assign outputs[141] = ~(layer4_outputs[1958]);
    assign outputs[142] = ~((layer4_outputs[1735]) | (layer4_outputs[2535]));
    assign outputs[143] = (layer4_outputs[1944]) & ~(layer4_outputs[880]);
    assign outputs[144] = ~((layer4_outputs[1128]) ^ (layer4_outputs[2404]));
    assign outputs[145] = layer4_outputs[2011];
    assign outputs[146] = layer4_outputs[821];
    assign outputs[147] = layer4_outputs[711];
    assign outputs[148] = ~(layer4_outputs[2266]);
    assign outputs[149] = ~(layer4_outputs[2053]);
    assign outputs[150] = (layer4_outputs[1389]) ^ (layer4_outputs[2259]);
    assign outputs[151] = ~(layer4_outputs[1623]);
    assign outputs[152] = ~(layer4_outputs[1845]);
    assign outputs[153] = (layer4_outputs[853]) | (layer4_outputs[1425]);
    assign outputs[154] = (layer4_outputs[2498]) ^ (layer4_outputs[42]);
    assign outputs[155] = layer4_outputs[457];
    assign outputs[156] = ~(layer4_outputs[2165]);
    assign outputs[157] = ~((layer4_outputs[1683]) & (layer4_outputs[163]));
    assign outputs[158] = ~(layer4_outputs[262]);
    assign outputs[159] = layer4_outputs[2097];
    assign outputs[160] = layer4_outputs[1083];
    assign outputs[161] = layer4_outputs[2112];
    assign outputs[162] = (layer4_outputs[27]) & (layer4_outputs[679]);
    assign outputs[163] = ~((layer4_outputs[1635]) ^ (layer4_outputs[456]));
    assign outputs[164] = ~(layer4_outputs[1543]) | (layer4_outputs[2443]);
    assign outputs[165] = ~((layer4_outputs[1693]) ^ (layer4_outputs[832]));
    assign outputs[166] = (layer4_outputs[635]) & ~(layer4_outputs[6]);
    assign outputs[167] = (layer4_outputs[1136]) & ~(layer4_outputs[793]);
    assign outputs[168] = layer4_outputs[2456];
    assign outputs[169] = layer4_outputs[1492];
    assign outputs[170] = ~((layer4_outputs[327]) ^ (layer4_outputs[2541]));
    assign outputs[171] = layer4_outputs[783];
    assign outputs[172] = ~((layer4_outputs[1894]) | (layer4_outputs[2459]));
    assign outputs[173] = ~(layer4_outputs[1470]);
    assign outputs[174] = ~((layer4_outputs[2317]) | (layer4_outputs[1524]));
    assign outputs[175] = layer4_outputs[301];
    assign outputs[176] = ~(layer4_outputs[793]);
    assign outputs[177] = (layer4_outputs[520]) & ~(layer4_outputs[541]);
    assign outputs[178] = ~(layer4_outputs[2157]);
    assign outputs[179] = layer4_outputs[2220];
    assign outputs[180] = ~(layer4_outputs[2322]);
    assign outputs[181] = layer4_outputs[1925];
    assign outputs[182] = layer4_outputs[1660];
    assign outputs[183] = ~(layer4_outputs[1563]);
    assign outputs[184] = (layer4_outputs[903]) & (layer4_outputs[389]);
    assign outputs[185] = (layer4_outputs[496]) ^ (layer4_outputs[1333]);
    assign outputs[186] = (layer4_outputs[1076]) ^ (layer4_outputs[1280]);
    assign outputs[187] = layer4_outputs[872];
    assign outputs[188] = layer4_outputs[550];
    assign outputs[189] = ~(layer4_outputs[1555]);
    assign outputs[190] = ~(layer4_outputs[129]);
    assign outputs[191] = (layer4_outputs[2094]) | (layer4_outputs[2289]);
    assign outputs[192] = layer4_outputs[2523];
    assign outputs[193] = ~(layer4_outputs[1447]);
    assign outputs[194] = ~((layer4_outputs[767]) ^ (layer4_outputs[2399]));
    assign outputs[195] = (layer4_outputs[1277]) & ~(layer4_outputs[1018]);
    assign outputs[196] = layer4_outputs[113];
    assign outputs[197] = ~(layer4_outputs[1589]);
    assign outputs[198] = ~((layer4_outputs[905]) ^ (layer4_outputs[383]));
    assign outputs[199] = layer4_outputs[1109];
    assign outputs[200] = layer4_outputs[772];
    assign outputs[201] = ~(layer4_outputs[1891]);
    assign outputs[202] = ~(layer4_outputs[2003]);
    assign outputs[203] = ~((layer4_outputs[471]) | (layer4_outputs[289]));
    assign outputs[204] = ~((layer4_outputs[1419]) | (layer4_outputs[2302]));
    assign outputs[205] = layer4_outputs[1888];
    assign outputs[206] = ~(layer4_outputs[1145]);
    assign outputs[207] = layer4_outputs[2379];
    assign outputs[208] = layer4_outputs[2449];
    assign outputs[209] = ~(layer4_outputs[2472]);
    assign outputs[210] = ~(layer4_outputs[1320]);
    assign outputs[211] = layer4_outputs[2483];
    assign outputs[212] = ~(layer4_outputs[993]) | (layer4_outputs[571]);
    assign outputs[213] = ~(layer4_outputs[977]);
    assign outputs[214] = layer4_outputs[2478];
    assign outputs[215] = layer4_outputs[913];
    assign outputs[216] = layer4_outputs[43];
    assign outputs[217] = (layer4_outputs[1798]) & ~(layer4_outputs[1567]);
    assign outputs[218] = ~(layer4_outputs[1792]) | (layer4_outputs[2158]);
    assign outputs[219] = layer4_outputs[1042];
    assign outputs[220] = layer4_outputs[1548];
    assign outputs[221] = layer4_outputs[325];
    assign outputs[222] = ~(layer4_outputs[2354]);
    assign outputs[223] = ~(layer4_outputs[1956]);
    assign outputs[224] = ~((layer4_outputs[1769]) ^ (layer4_outputs[648]));
    assign outputs[225] = layer4_outputs[1438];
    assign outputs[226] = layer4_outputs[910];
    assign outputs[227] = layer4_outputs[699];
    assign outputs[228] = ~(layer4_outputs[1098]);
    assign outputs[229] = ~(layer4_outputs[1965]);
    assign outputs[230] = ~(layer4_outputs[687]);
    assign outputs[231] = ~(layer4_outputs[236]);
    assign outputs[232] = ~(layer4_outputs[2492]);
    assign outputs[233] = layer4_outputs[1927];
    assign outputs[234] = layer4_outputs[60];
    assign outputs[235] = ~(layer4_outputs[2555]) | (layer4_outputs[2552]);
    assign outputs[236] = layer4_outputs[447];
    assign outputs[237] = layer4_outputs[821];
    assign outputs[238] = layer4_outputs[50];
    assign outputs[239] = ~(layer4_outputs[153]);
    assign outputs[240] = (layer4_outputs[1213]) & (layer4_outputs[2101]);
    assign outputs[241] = ~((layer4_outputs[1838]) ^ (layer4_outputs[2477]));
    assign outputs[242] = layer4_outputs[2000];
    assign outputs[243] = ~(layer4_outputs[26]) | (layer4_outputs[529]);
    assign outputs[244] = ~(layer4_outputs[927]);
    assign outputs[245] = ~((layer4_outputs[2065]) | (layer4_outputs[1781]));
    assign outputs[246] = layer4_outputs[2359];
    assign outputs[247] = ~(layer4_outputs[1084]);
    assign outputs[248] = layer4_outputs[2386];
    assign outputs[249] = (layer4_outputs[2483]) & (layer4_outputs[444]);
    assign outputs[250] = ~(layer4_outputs[1698]);
    assign outputs[251] = (layer4_outputs[910]) & ~(layer4_outputs[1080]);
    assign outputs[252] = (layer4_outputs[138]) & ~(layer4_outputs[1263]);
    assign outputs[253] = layer4_outputs[1904];
    assign outputs[254] = (layer4_outputs[1770]) & ~(layer4_outputs[2275]);
    assign outputs[255] = ~(layer4_outputs[14]);
    assign outputs[256] = layer4_outputs[1280];
    assign outputs[257] = ~(layer4_outputs[1759]);
    assign outputs[258] = (layer4_outputs[528]) & (layer4_outputs[2141]);
    assign outputs[259] = (layer4_outputs[68]) & ~(layer4_outputs[1822]);
    assign outputs[260] = (layer4_outputs[1950]) & ~(layer4_outputs[348]);
    assign outputs[261] = (layer4_outputs[1436]) & ~(layer4_outputs[2417]);
    assign outputs[262] = layer4_outputs[1528];
    assign outputs[263] = (layer4_outputs[120]) & ~(layer4_outputs[478]);
    assign outputs[264] = (layer4_outputs[1663]) & ~(layer4_outputs[1794]);
    assign outputs[265] = (layer4_outputs[1806]) & ~(layer4_outputs[2327]);
    assign outputs[266] = (layer4_outputs[814]) & ~(layer4_outputs[1559]);
    assign outputs[267] = ~(layer4_outputs[1017]);
    assign outputs[268] = (layer4_outputs[267]) & ~(layer4_outputs[2516]);
    assign outputs[269] = (layer4_outputs[919]) & ~(layer4_outputs[1075]);
    assign outputs[270] = layer4_outputs[1917];
    assign outputs[271] = ~(layer4_outputs[2028]);
    assign outputs[272] = ~((layer4_outputs[2156]) | (layer4_outputs[901]));
    assign outputs[273] = layer4_outputs[124];
    assign outputs[274] = ~(layer4_outputs[1212]);
    assign outputs[275] = ~(layer4_outputs[1368]);
    assign outputs[276] = ~((layer4_outputs[2411]) ^ (layer4_outputs[1657]));
    assign outputs[277] = (layer4_outputs[655]) & (layer4_outputs[1304]);
    assign outputs[278] = (layer4_outputs[780]) | (layer4_outputs[1163]);
    assign outputs[279] = ~((layer4_outputs[1352]) ^ (layer4_outputs[7]));
    assign outputs[280] = ~((layer4_outputs[12]) | (layer4_outputs[1882]));
    assign outputs[281] = (layer4_outputs[1382]) ^ (layer4_outputs[1217]);
    assign outputs[282] = (layer4_outputs[16]) & ~(layer4_outputs[499]);
    assign outputs[283] = (layer4_outputs[1614]) & ~(layer4_outputs[1177]);
    assign outputs[284] = (layer4_outputs[1752]) & (layer4_outputs[141]);
    assign outputs[285] = layer4_outputs[807];
    assign outputs[286] = (layer4_outputs[536]) & (layer4_outputs[317]);
    assign outputs[287] = ~(layer4_outputs[1278]);
    assign outputs[288] = ~((layer4_outputs[544]) & (layer4_outputs[188]));
    assign outputs[289] = ~(layer4_outputs[756]) | (layer4_outputs[1695]);
    assign outputs[290] = ~(layer4_outputs[1366]);
    assign outputs[291] = layer4_outputs[2030];
    assign outputs[292] = (layer4_outputs[2471]) ^ (layer4_outputs[35]);
    assign outputs[293] = ~((layer4_outputs[1102]) | (layer4_outputs[170]));
    assign outputs[294] = ~(layer4_outputs[1864]);
    assign outputs[295] = (layer4_outputs[2442]) & ~(layer4_outputs[1094]);
    assign outputs[296] = (layer4_outputs[1024]) & ~(layer4_outputs[852]);
    assign outputs[297] = layer4_outputs[236];
    assign outputs[298] = (layer4_outputs[549]) & ~(layer4_outputs[2485]);
    assign outputs[299] = ~(layer4_outputs[1841]);
    assign outputs[300] = (layer4_outputs[576]) & (layer4_outputs[310]);
    assign outputs[301] = ~(layer4_outputs[2284]);
    assign outputs[302] = ~(layer4_outputs[1923]);
    assign outputs[303] = (layer4_outputs[2145]) & (layer4_outputs[6]);
    assign outputs[304] = (layer4_outputs[631]) ^ (layer4_outputs[649]);
    assign outputs[305] = ~(layer4_outputs[1924]);
    assign outputs[306] = layer4_outputs[1492];
    assign outputs[307] = ~((layer4_outputs[212]) | (layer4_outputs[1925]));
    assign outputs[308] = ~((layer4_outputs[1593]) | (layer4_outputs[466]));
    assign outputs[309] = layer4_outputs[1603];
    assign outputs[310] = ~(layer4_outputs[2024]) | (layer4_outputs[1322]);
    assign outputs[311] = ~((layer4_outputs[2070]) | (layer4_outputs[2454]));
    assign outputs[312] = ~(layer4_outputs[59]);
    assign outputs[313] = layer4_outputs[2445];
    assign outputs[314] = (layer4_outputs[892]) & ~(layer4_outputs[493]);
    assign outputs[315] = layer4_outputs[1302];
    assign outputs[316] = ~((layer4_outputs[855]) | (layer4_outputs[1417]));
    assign outputs[317] = ~((layer4_outputs[2286]) ^ (layer4_outputs[193]));
    assign outputs[318] = (layer4_outputs[477]) ^ (layer4_outputs[2191]);
    assign outputs[319] = (layer4_outputs[1535]) & ~(layer4_outputs[460]);
    assign outputs[320] = layer4_outputs[2052];
    assign outputs[321] = (layer4_outputs[408]) & ~(layer4_outputs[988]);
    assign outputs[322] = layer4_outputs[2453];
    assign outputs[323] = layer4_outputs[1781];
    assign outputs[324] = ~(layer4_outputs[1972]);
    assign outputs[325] = (layer4_outputs[2293]) ^ (layer4_outputs[2094]);
    assign outputs[326] = ~(layer4_outputs[463]) | (layer4_outputs[771]);
    assign outputs[327] = ~((layer4_outputs[1224]) | (layer4_outputs[595]));
    assign outputs[328] = ~(layer4_outputs[380]) | (layer4_outputs[203]);
    assign outputs[329] = layer4_outputs[1127];
    assign outputs[330] = ~(layer4_outputs[1903]);
    assign outputs[331] = (layer4_outputs[382]) & (layer4_outputs[8]);
    assign outputs[332] = layer4_outputs[604];
    assign outputs[333] = layer4_outputs[2554];
    assign outputs[334] = (layer4_outputs[601]) & ~(layer4_outputs[2085]);
    assign outputs[335] = (layer4_outputs[1538]) & ~(layer4_outputs[1679]);
    assign outputs[336] = layer4_outputs[1509];
    assign outputs[337] = (layer4_outputs[705]) ^ (layer4_outputs[2368]);
    assign outputs[338] = (layer4_outputs[937]) & ~(layer4_outputs[865]);
    assign outputs[339] = ~(layer4_outputs[1478]);
    assign outputs[340] = (layer4_outputs[1175]) ^ (layer4_outputs[1952]);
    assign outputs[341] = ~(layer4_outputs[1305]);
    assign outputs[342] = ~(layer4_outputs[843]);
    assign outputs[343] = layer4_outputs[1523];
    assign outputs[344] = (layer4_outputs[859]) & (layer4_outputs[1900]);
    assign outputs[345] = ~((layer4_outputs[2326]) ^ (layer4_outputs[1536]));
    assign outputs[346] = layer4_outputs[1358];
    assign outputs[347] = (layer4_outputs[2145]) & ~(layer4_outputs[232]);
    assign outputs[348] = (layer4_outputs[2382]) & ~(layer4_outputs[826]);
    assign outputs[349] = (layer4_outputs[2491]) & ~(layer4_outputs[1642]);
    assign outputs[350] = layer4_outputs[2267];
    assign outputs[351] = (layer4_outputs[1236]) & (layer4_outputs[2161]);
    assign outputs[352] = (layer4_outputs[1161]) & ~(layer4_outputs[1033]);
    assign outputs[353] = layer4_outputs[990];
    assign outputs[354] = (layer4_outputs[917]) & ~(layer4_outputs[1643]);
    assign outputs[355] = (layer4_outputs[379]) & ~(layer4_outputs[2168]);
    assign outputs[356] = ~(layer4_outputs[2134]);
    assign outputs[357] = ~(layer4_outputs[1207]);
    assign outputs[358] = (layer4_outputs[433]) ^ (layer4_outputs[411]);
    assign outputs[359] = ~(layer4_outputs[154]) | (layer4_outputs[2313]);
    assign outputs[360] = (layer4_outputs[373]) ^ (layer4_outputs[1989]);
    assign outputs[361] = (layer4_outputs[2492]) ^ (layer4_outputs[772]);
    assign outputs[362] = ~(layer4_outputs[744]);
    assign outputs[363] = layer4_outputs[2290];
    assign outputs[364] = ~((layer4_outputs[1739]) | (layer4_outputs[976]));
    assign outputs[365] = ~(layer4_outputs[1875]);
    assign outputs[366] = layer4_outputs[1595];
    assign outputs[367] = (layer4_outputs[2243]) & (layer4_outputs[1646]);
    assign outputs[368] = ~((layer4_outputs[796]) | (layer4_outputs[2156]));
    assign outputs[369] = layer4_outputs[1396];
    assign outputs[370] = ~(layer4_outputs[2420]);
    assign outputs[371] = ~(layer4_outputs[2186]);
    assign outputs[372] = ~(layer4_outputs[1893]);
    assign outputs[373] = ~(layer4_outputs[945]) | (layer4_outputs[1633]);
    assign outputs[374] = (layer4_outputs[579]) & (layer4_outputs[1743]);
    assign outputs[375] = ~(layer4_outputs[2502]);
    assign outputs[376] = ~(layer4_outputs[1935]);
    assign outputs[377] = (layer4_outputs[2246]) ^ (layer4_outputs[2474]);
    assign outputs[378] = (layer4_outputs[2264]) ^ (layer4_outputs[291]);
    assign outputs[379] = ~((layer4_outputs[1631]) | (layer4_outputs[1175]));
    assign outputs[380] = ~(layer4_outputs[395]);
    assign outputs[381] = ~(layer4_outputs[2349]);
    assign outputs[382] = (layer4_outputs[1957]) & (layer4_outputs[940]);
    assign outputs[383] = ~(layer4_outputs[1970]);
    assign outputs[384] = (layer4_outputs[899]) & (layer4_outputs[627]);
    assign outputs[385] = ~(layer4_outputs[2332]);
    assign outputs[386] = (layer4_outputs[2146]) & ~(layer4_outputs[1465]);
    assign outputs[387] = ~(layer4_outputs[1745]);
    assign outputs[388] = (layer4_outputs[1620]) ^ (layer4_outputs[419]);
    assign outputs[389] = layer4_outputs[1006];
    assign outputs[390] = (layer4_outputs[86]) & ~(layer4_outputs[1416]);
    assign outputs[391] = (layer4_outputs[1627]) & (layer4_outputs[99]);
    assign outputs[392] = (layer4_outputs[1156]) & ~(layer4_outputs[192]);
    assign outputs[393] = (layer4_outputs[2345]) & (layer4_outputs[296]);
    assign outputs[394] = layer4_outputs[1529];
    assign outputs[395] = layer4_outputs[1066];
    assign outputs[396] = layer4_outputs[861];
    assign outputs[397] = ~(layer4_outputs[1816]);
    assign outputs[398] = ~(layer4_outputs[64]);
    assign outputs[399] = ~((layer4_outputs[2286]) | (layer4_outputs[1305]));
    assign outputs[400] = (layer4_outputs[97]) & ~(layer4_outputs[2017]);
    assign outputs[401] = (layer4_outputs[914]) ^ (layer4_outputs[2305]);
    assign outputs[402] = ~((layer4_outputs[836]) ^ (layer4_outputs[2401]));
    assign outputs[403] = layer4_outputs[1005];
    assign outputs[404] = ~(layer4_outputs[175]);
    assign outputs[405] = layer4_outputs[308];
    assign outputs[406] = (layer4_outputs[1137]) ^ (layer4_outputs[2147]);
    assign outputs[407] = ~((layer4_outputs[1221]) | (layer4_outputs[83]));
    assign outputs[408] = (layer4_outputs[1302]) & ~(layer4_outputs[1915]);
    assign outputs[409] = (layer4_outputs[1606]) ^ (layer4_outputs[501]);
    assign outputs[410] = layer4_outputs[2004];
    assign outputs[411] = ~((layer4_outputs[2066]) | (layer4_outputs[119]));
    assign outputs[412] = (layer4_outputs[362]) & ~(layer4_outputs[1244]);
    assign outputs[413] = layer4_outputs[2105];
    assign outputs[414] = ~(layer4_outputs[1676]);
    assign outputs[415] = (layer4_outputs[2075]) & (layer4_outputs[1122]);
    assign outputs[416] = layer4_outputs[1501];
    assign outputs[417] = ~((layer4_outputs[849]) | (layer4_outputs[1118]));
    assign outputs[418] = (layer4_outputs[1462]) & (layer4_outputs[1463]);
    assign outputs[419] = layer4_outputs[722];
    assign outputs[420] = ~(layer4_outputs[546]);
    assign outputs[421] = (layer4_outputs[1229]) & (layer4_outputs[1091]);
    assign outputs[422] = ~(layer4_outputs[207]);
    assign outputs[423] = (layer4_outputs[1803]) & ~(layer4_outputs[238]);
    assign outputs[424] = (layer4_outputs[1209]) & ~(layer4_outputs[50]);
    assign outputs[425] = (layer4_outputs[919]) & (layer4_outputs[1456]);
    assign outputs[426] = (layer4_outputs[2448]) & (layer4_outputs[1322]);
    assign outputs[427] = ~((layer4_outputs[2238]) ^ (layer4_outputs[934]));
    assign outputs[428] = ~(layer4_outputs[1771]);
    assign outputs[429] = (layer4_outputs[448]) ^ (layer4_outputs[206]);
    assign outputs[430] = layer4_outputs[985];
    assign outputs[431] = (layer4_outputs[1987]) & ~(layer4_outputs[10]);
    assign outputs[432] = ~((layer4_outputs[2432]) ^ (layer4_outputs[1876]));
    assign outputs[433] = (layer4_outputs[2263]) & ~(layer4_outputs[175]);
    assign outputs[434] = layer4_outputs[1047];
    assign outputs[435] = layer4_outputs[1341];
    assign outputs[436] = (layer4_outputs[1450]) & (layer4_outputs[532]);
    assign outputs[437] = (layer4_outputs[190]) & (layer4_outputs[275]);
    assign outputs[438] = layer4_outputs[1787];
    assign outputs[439] = (layer4_outputs[999]) & (layer4_outputs[1717]);
    assign outputs[440] = (layer4_outputs[806]) & (layer4_outputs[655]);
    assign outputs[441] = (layer4_outputs[1613]) & ~(layer4_outputs[410]);
    assign outputs[442] = ~(layer4_outputs[1179]);
    assign outputs[443] = ~(layer4_outputs[385]);
    assign outputs[444] = (layer4_outputs[1523]) & ~(layer4_outputs[734]);
    assign outputs[445] = ~(layer4_outputs[1254]);
    assign outputs[446] = ~(layer4_outputs[1788]);
    assign outputs[447] = (layer4_outputs[2239]) & ~(layer4_outputs[2393]);
    assign outputs[448] = (layer4_outputs[1157]) & ~(layer4_outputs[1035]);
    assign outputs[449] = ~(layer4_outputs[507]);
    assign outputs[450] = layer4_outputs[47];
    assign outputs[451] = (layer4_outputs[1512]) & ~(layer4_outputs[248]);
    assign outputs[452] = (layer4_outputs[346]) & ~(layer4_outputs[2220]);
    assign outputs[453] = layer4_outputs[320];
    assign outputs[454] = layer4_outputs[182];
    assign outputs[455] = ~(layer4_outputs[1132]);
    assign outputs[456] = ~(layer4_outputs[1814]);
    assign outputs[457] = ~((layer4_outputs[435]) | (layer4_outputs[1700]));
    assign outputs[458] = layer4_outputs[2507];
    assign outputs[459] = (layer4_outputs[2297]) ^ (layer4_outputs[674]);
    assign outputs[460] = (layer4_outputs[189]) & (layer4_outputs[1580]);
    assign outputs[461] = (layer4_outputs[1663]) & ~(layer4_outputs[1670]);
    assign outputs[462] = ~((layer4_outputs[1179]) | (layer4_outputs[2085]));
    assign outputs[463] = layer4_outputs[2309];
    assign outputs[464] = ~(layer4_outputs[1264]);
    assign outputs[465] = ~(layer4_outputs[1058]);
    assign outputs[466] = ~(layer4_outputs[1306]);
    assign outputs[467] = ~(layer4_outputs[1578]);
    assign outputs[468] = ~((layer4_outputs[7]) ^ (layer4_outputs[1441]));
    assign outputs[469] = ~(layer4_outputs[2211]);
    assign outputs[470] = (layer4_outputs[665]) ^ (layer4_outputs[696]);
    assign outputs[471] = (layer4_outputs[2462]) & (layer4_outputs[2497]);
    assign outputs[472] = layer4_outputs[1314];
    assign outputs[473] = ~((layer4_outputs[1843]) | (layer4_outputs[715]));
    assign outputs[474] = (layer4_outputs[1055]) & ~(layer4_outputs[404]);
    assign outputs[475] = (layer4_outputs[2453]) | (layer4_outputs[1513]);
    assign outputs[476] = (layer4_outputs[1612]) & (layer4_outputs[1859]);
    assign outputs[477] = layer4_outputs[2556];
    assign outputs[478] = ~((layer4_outputs[2219]) | (layer4_outputs[1364]));
    assign outputs[479] = (layer4_outputs[560]) & (layer4_outputs[2363]);
    assign outputs[480] = ~((layer4_outputs[817]) | (layer4_outputs[1226]));
    assign outputs[481] = (layer4_outputs[353]) & (layer4_outputs[297]);
    assign outputs[482] = (layer4_outputs[2486]) & (layer4_outputs[834]);
    assign outputs[483] = ~(layer4_outputs[2409]);
    assign outputs[484] = ~(layer4_outputs[323]);
    assign outputs[485] = (layer4_outputs[1859]) & ~(layer4_outputs[2128]);
    assign outputs[486] = (layer4_outputs[2366]) & (layer4_outputs[2142]);
    assign outputs[487] = (layer4_outputs[651]) & ~(layer4_outputs[1398]);
    assign outputs[488] = (layer4_outputs[2057]) & (layer4_outputs[2064]);
    assign outputs[489] = layer4_outputs[685];
    assign outputs[490] = ~(layer4_outputs[2230]);
    assign outputs[491] = (layer4_outputs[1476]) ^ (layer4_outputs[756]);
    assign outputs[492] = layer4_outputs[991];
    assign outputs[493] = ~(layer4_outputs[1823]);
    assign outputs[494] = layer4_outputs[1470];
    assign outputs[495] = (layer4_outputs[1440]) & (layer4_outputs[1860]);
    assign outputs[496] = layer4_outputs[1878];
    assign outputs[497] = ~(layer4_outputs[1756]);
    assign outputs[498] = (layer4_outputs[2557]) & ~(layer4_outputs[1338]);
    assign outputs[499] = layer4_outputs[2336];
    assign outputs[500] = ~((layer4_outputs[2022]) | (layer4_outputs[2361]));
    assign outputs[501] = ~((layer4_outputs[440]) | (layer4_outputs[1342]));
    assign outputs[502] = ~((layer4_outputs[178]) | (layer4_outputs[2067]));
    assign outputs[503] = layer4_outputs[1065];
    assign outputs[504] = (layer4_outputs[473]) & ~(layer4_outputs[754]);
    assign outputs[505] = layer4_outputs[142];
    assign outputs[506] = (layer4_outputs[2092]) & ~(layer4_outputs[555]);
    assign outputs[507] = ~(layer4_outputs[2302]);
    assign outputs[508] = ~((layer4_outputs[1552]) ^ (layer4_outputs[670]));
    assign outputs[509] = ~((layer4_outputs[2020]) ^ (layer4_outputs[84]));
    assign outputs[510] = layer4_outputs[1786];
    assign outputs[511] = (layer4_outputs[533]) & ~(layer4_outputs[1797]);
    assign outputs[512] = layer4_outputs[1858];
    assign outputs[513] = ~(layer4_outputs[1655]);
    assign outputs[514] = ~((layer4_outputs[167]) | (layer4_outputs[1843]));
    assign outputs[515] = layer4_outputs[504];
    assign outputs[516] = (layer4_outputs[858]) & (layer4_outputs[2402]);
    assign outputs[517] = layer4_outputs[74];
    assign outputs[518] = layer4_outputs[1101];
    assign outputs[519] = ~(layer4_outputs[555]);
    assign outputs[520] = ~(layer4_outputs[167]) | (layer4_outputs[2002]);
    assign outputs[521] = layer4_outputs[1203];
    assign outputs[522] = ~((layer4_outputs[2367]) | (layer4_outputs[264]));
    assign outputs[523] = ~(layer4_outputs[1789]);
    assign outputs[524] = (layer4_outputs[604]) ^ (layer4_outputs[614]);
    assign outputs[525] = ~(layer4_outputs[1933]);
    assign outputs[526] = ~(layer4_outputs[368]);
    assign outputs[527] = layer4_outputs[1126];
    assign outputs[528] = layer4_outputs[1602];
    assign outputs[529] = layer4_outputs[1517];
    assign outputs[530] = (layer4_outputs[2247]) & (layer4_outputs[1915]);
    assign outputs[531] = layer4_outputs[89];
    assign outputs[532] = ~(layer4_outputs[1817]);
    assign outputs[533] = ~(layer4_outputs[1712]);
    assign outputs[534] = ~(layer4_outputs[155]);
    assign outputs[535] = ~(layer4_outputs[639]) | (layer4_outputs[2438]);
    assign outputs[536] = ~(layer4_outputs[1877]);
    assign outputs[537] = ~(layer4_outputs[945]);
    assign outputs[538] = (layer4_outputs[847]) & ~(layer4_outputs[1736]);
    assign outputs[539] = ~(layer4_outputs[2042]) | (layer4_outputs[1532]);
    assign outputs[540] = layer4_outputs[2403];
    assign outputs[541] = layer4_outputs[1943];
    assign outputs[542] = ~(layer4_outputs[243]);
    assign outputs[543] = ~(layer4_outputs[575]);
    assign outputs[544] = ~(layer4_outputs[2254]) | (layer4_outputs[2294]);
    assign outputs[545] = ~(layer4_outputs[1199]);
    assign outputs[546] = ~((layer4_outputs[2497]) ^ (layer4_outputs[1752]));
    assign outputs[547] = ~(layer4_outputs[14]);
    assign outputs[548] = ~(layer4_outputs[1451]);
    assign outputs[549] = ~(layer4_outputs[1276]);
    assign outputs[550] = (layer4_outputs[998]) & ~(layer4_outputs[1011]);
    assign outputs[551] = ~((layer4_outputs[1567]) | (layer4_outputs[1982]));
    assign outputs[552] = ~(layer4_outputs[1722]);
    assign outputs[553] = (layer4_outputs[2481]) ^ (layer4_outputs[1315]);
    assign outputs[554] = layer4_outputs[511];
    assign outputs[555] = layer4_outputs[2491];
    assign outputs[556] = layer4_outputs[2444];
    assign outputs[557] = layer4_outputs[58];
    assign outputs[558] = ~(layer4_outputs[269]);
    assign outputs[559] = layer4_outputs[525];
    assign outputs[560] = ~(layer4_outputs[952]);
    assign outputs[561] = layer4_outputs[1953];
    assign outputs[562] = layer4_outputs[543];
    assign outputs[563] = (layer4_outputs[136]) | (layer4_outputs[1131]);
    assign outputs[564] = ~(layer4_outputs[2269]);
    assign outputs[565] = ~(layer4_outputs[299]);
    assign outputs[566] = (layer4_outputs[675]) ^ (layer4_outputs[569]);
    assign outputs[567] = layer4_outputs[1399];
    assign outputs[568] = (layer4_outputs[996]) & ~(layer4_outputs[268]);
    assign outputs[569] = layer4_outputs[32];
    assign outputs[570] = ~(layer4_outputs[416]);
    assign outputs[571] = ~(layer4_outputs[2013]);
    assign outputs[572] = ~(layer4_outputs[107]);
    assign outputs[573] = layer4_outputs[2523];
    assign outputs[574] = layer4_outputs[91];
    assign outputs[575] = ~(layer4_outputs[1935]);
    assign outputs[576] = (layer4_outputs[1759]) ^ (layer4_outputs[1868]);
    assign outputs[577] = ~(layer4_outputs[133]);
    assign outputs[578] = layer4_outputs[1495];
    assign outputs[579] = ~(layer4_outputs[947]);
    assign outputs[580] = layer4_outputs[306];
    assign outputs[581] = layer4_outputs[648];
    assign outputs[582] = layer4_outputs[535];
    assign outputs[583] = layer4_outputs[718];
    assign outputs[584] = ~(layer4_outputs[769]);
    assign outputs[585] = ~(layer4_outputs[1847]);
    assign outputs[586] = layer4_outputs[2231];
    assign outputs[587] = ~(layer4_outputs[788]);
    assign outputs[588] = ~((layer4_outputs[943]) & (layer4_outputs[1490]));
    assign outputs[589] = ~(layer4_outputs[554]);
    assign outputs[590] = ~(layer4_outputs[1974]) | (layer4_outputs[1688]);
    assign outputs[591] = ~(layer4_outputs[457]);
    assign outputs[592] = ~(layer4_outputs[2031]);
    assign outputs[593] = (layer4_outputs[331]) & ~(layer4_outputs[1346]);
    assign outputs[594] = layer4_outputs[2182];
    assign outputs[595] = (layer4_outputs[1325]) & ~(layer4_outputs[1926]);
    assign outputs[596] = ~(layer4_outputs[1357]);
    assign outputs[597] = ~(layer4_outputs[1334]);
    assign outputs[598] = ~(layer4_outputs[1981]);
    assign outputs[599] = ~(layer4_outputs[1960]);
    assign outputs[600] = (layer4_outputs[1574]) & (layer4_outputs[1074]);
    assign outputs[601] = layer4_outputs[1579];
    assign outputs[602] = ~((layer4_outputs[758]) ^ (layer4_outputs[1204]));
    assign outputs[603] = layer4_outputs[1348];
    assign outputs[604] = layer4_outputs[768];
    assign outputs[605] = layer4_outputs[2035];
    assign outputs[606] = (layer4_outputs[953]) ^ (layer4_outputs[1991]);
    assign outputs[607] = layer4_outputs[2512];
    assign outputs[608] = ~((layer4_outputs[1961]) ^ (layer4_outputs[628]));
    assign outputs[609] = (layer4_outputs[2525]) | (layer4_outputs[2501]);
    assign outputs[610] = (layer4_outputs[67]) | (layer4_outputs[1373]);
    assign outputs[611] = (layer4_outputs[2355]) ^ (layer4_outputs[2481]);
    assign outputs[612] = ~(layer4_outputs[820]);
    assign outputs[613] = ~(layer4_outputs[2068]);
    assign outputs[614] = layer4_outputs[2057];
    assign outputs[615] = ~(layer4_outputs[2426]);
    assign outputs[616] = layer4_outputs[511];
    assign outputs[617] = (layer4_outputs[307]) ^ (layer4_outputs[789]);
    assign outputs[618] = (layer4_outputs[1216]) & (layer4_outputs[1246]);
    assign outputs[619] = ~(layer4_outputs[1847]);
    assign outputs[620] = (layer4_outputs[2357]) & ~(layer4_outputs[1373]);
    assign outputs[621] = ~(layer4_outputs[2110]);
    assign outputs[622] = ~((layer4_outputs[211]) | (layer4_outputs[2086]));
    assign outputs[623] = ~(layer4_outputs[2391]) | (layer4_outputs[1196]);
    assign outputs[624] = ~(layer4_outputs[933]);
    assign outputs[625] = ~(layer4_outputs[1509]);
    assign outputs[626] = ~(layer4_outputs[1585]);
    assign outputs[627] = (layer4_outputs[298]) ^ (layer4_outputs[108]);
    assign outputs[628] = layer4_outputs[2440];
    assign outputs[629] = (layer4_outputs[441]) ^ (layer4_outputs[2458]);
    assign outputs[630] = (layer4_outputs[1846]) & ~(layer4_outputs[599]);
    assign outputs[631] = ~(layer4_outputs[1429]);
    assign outputs[632] = (layer4_outputs[1964]) & ~(layer4_outputs[1346]);
    assign outputs[633] = ~(layer4_outputs[2299]);
    assign outputs[634] = ~(layer4_outputs[1477]);
    assign outputs[635] = ~(layer4_outputs[2055]);
    assign outputs[636] = (layer4_outputs[2118]) & ~(layer4_outputs[775]);
    assign outputs[637] = ~((layer4_outputs[946]) & (layer4_outputs[2169]));
    assign outputs[638] = ~(layer4_outputs[813]);
    assign outputs[639] = (layer4_outputs[2160]) ^ (layer4_outputs[44]);
    assign outputs[640] = (layer4_outputs[205]) & ~(layer4_outputs[423]);
    assign outputs[641] = ~((layer4_outputs[102]) ^ (layer4_outputs[1748]));
    assign outputs[642] = (layer4_outputs[876]) ^ (layer4_outputs[1650]);
    assign outputs[643] = layer4_outputs[1460];
    assign outputs[644] = layer4_outputs[1997];
    assign outputs[645] = ~(layer4_outputs[2339]);
    assign outputs[646] = ~(layer4_outputs[2460]);
    assign outputs[647] = ~(layer4_outputs[2380]);
    assign outputs[648] = layer4_outputs[622];
    assign outputs[649] = ~(layer4_outputs[796]);
    assign outputs[650] = ~(layer4_outputs[73]);
    assign outputs[651] = layer4_outputs[1485];
    assign outputs[652] = ~(layer4_outputs[522]);
    assign outputs[653] = layer4_outputs[1068];
    assign outputs[654] = ~(layer4_outputs[1931]) | (layer4_outputs[1215]);
    assign outputs[655] = ~(layer4_outputs[2162]) | (layer4_outputs[746]);
    assign outputs[656] = ~((layer4_outputs[295]) ^ (layer4_outputs[1762]));
    assign outputs[657] = ~(layer4_outputs[1355]);
    assign outputs[658] = (layer4_outputs[294]) & (layer4_outputs[98]);
    assign outputs[659] = ~(layer4_outputs[566]);
    assign outputs[660] = (layer4_outputs[640]) ^ (layer4_outputs[1420]);
    assign outputs[661] = ~(layer4_outputs[429]);
    assign outputs[662] = layer4_outputs[578];
    assign outputs[663] = (layer4_outputs[1810]) & ~(layer4_outputs[1371]);
    assign outputs[664] = layer4_outputs[1677];
    assign outputs[665] = (layer4_outputs[2266]) & ~(layer4_outputs[740]);
    assign outputs[666] = (layer4_outputs[1622]) & (layer4_outputs[1671]);
    assign outputs[667] = (layer4_outputs[1745]) ^ (layer4_outputs[2108]);
    assign outputs[668] = (layer4_outputs[1669]) ^ (layer4_outputs[468]);
    assign outputs[669] = ~(layer4_outputs[1713]) | (layer4_outputs[2408]);
    assign outputs[670] = (layer4_outputs[2375]) & ~(layer4_outputs[1842]);
    assign outputs[671] = ~(layer4_outputs[729]);
    assign outputs[672] = (layer4_outputs[1044]) & ~(layer4_outputs[1250]);
    assign outputs[673] = ~(layer4_outputs[2235]);
    assign outputs[674] = ~(layer4_outputs[739]);
    assign outputs[675] = (layer4_outputs[1135]) & ~(layer4_outputs[1211]);
    assign outputs[676] = layer4_outputs[1437];
    assign outputs[677] = layer4_outputs[364];
    assign outputs[678] = ~(layer4_outputs[1317]);
    assign outputs[679] = layer4_outputs[609];
    assign outputs[680] = layer4_outputs[1708];
    assign outputs[681] = layer4_outputs[1195];
    assign outputs[682] = ~(layer4_outputs[248]);
    assign outputs[683] = ~((layer4_outputs[1320]) & (layer4_outputs[1121]));
    assign outputs[684] = layer4_outputs[497];
    assign outputs[685] = layer4_outputs[1232];
    assign outputs[686] = (layer4_outputs[356]) & (layer4_outputs[1720]);
    assign outputs[687] = layer4_outputs[361];
    assign outputs[688] = ~(layer4_outputs[1823]);
    assign outputs[689] = ~(layer4_outputs[1723]);
    assign outputs[690] = layer4_outputs[179];
    assign outputs[691] = (layer4_outputs[495]) & (layer4_outputs[1308]);
    assign outputs[692] = layer4_outputs[384];
    assign outputs[693] = (layer4_outputs[1006]) & ~(layer4_outputs[2113]);
    assign outputs[694] = layer4_outputs[398];
    assign outputs[695] = ~(layer4_outputs[2460]);
    assign outputs[696] = (layer4_outputs[2074]) | (layer4_outputs[1505]);
    assign outputs[697] = ~(layer4_outputs[2475]);
    assign outputs[698] = (layer4_outputs[2509]) ^ (layer4_outputs[315]);
    assign outputs[699] = ~(layer4_outputs[776]) | (layer4_outputs[637]);
    assign outputs[700] = ~((layer4_outputs[1020]) ^ (layer4_outputs[1149]));
    assign outputs[701] = ~(layer4_outputs[408]) | (layer4_outputs[1746]);
    assign outputs[702] = ~(layer4_outputs[258]);
    assign outputs[703] = ~((layer4_outputs[2511]) | (layer4_outputs[1906]));
    assign outputs[704] = layer4_outputs[1506];
    assign outputs[705] = layer4_outputs[2413];
    assign outputs[706] = ~(layer4_outputs[1564]);
    assign outputs[707] = layer4_outputs[1424];
    assign outputs[708] = ~((layer4_outputs[292]) & (layer4_outputs[1792]));
    assign outputs[709] = ~(layer4_outputs[2318]);
    assign outputs[710] = layer4_outputs[1471];
    assign outputs[711] = layer4_outputs[1459];
    assign outputs[712] = ~(layer4_outputs[964]);
    assign outputs[713] = layer4_outputs[2045];
    assign outputs[714] = layer4_outputs[1740];
    assign outputs[715] = ~((layer4_outputs[1223]) ^ (layer4_outputs[1979]));
    assign outputs[716] = ~((layer4_outputs[611]) | (layer4_outputs[1825]));
    assign outputs[717] = ~((layer4_outputs[2273]) ^ (layer4_outputs[582]));
    assign outputs[718] = ~(layer4_outputs[2346]);
    assign outputs[719] = layer4_outputs[1622];
    assign outputs[720] = ~((layer4_outputs[828]) ^ (layer4_outputs[762]));
    assign outputs[721] = layer4_outputs[1237];
    assign outputs[722] = layer4_outputs[18];
    assign outputs[723] = layer4_outputs[861];
    assign outputs[724] = layer4_outputs[660];
    assign outputs[725] = layer4_outputs[32];
    assign outputs[726] = layer4_outputs[1733];
    assign outputs[727] = ~(layer4_outputs[126]);
    assign outputs[728] = ~(layer4_outputs[470]);
    assign outputs[729] = layer4_outputs[2464];
    assign outputs[730] = ~((layer4_outputs[742]) ^ (layer4_outputs[1464]));
    assign outputs[731] = layer4_outputs[428];
    assign outputs[732] = ~(layer4_outputs[107]);
    assign outputs[733] = layer4_outputs[146];
    assign outputs[734] = layer4_outputs[1325];
    assign outputs[735] = ~(layer4_outputs[1960]);
    assign outputs[736] = ~((layer4_outputs[2530]) ^ (layer4_outputs[862]));
    assign outputs[737] = layer4_outputs[1431];
    assign outputs[738] = (layer4_outputs[2350]) & ~(layer4_outputs[1249]);
    assign outputs[739] = ~(layer4_outputs[1749]);
    assign outputs[740] = ~(layer4_outputs[1711]) | (layer4_outputs[1205]);
    assign outputs[741] = layer4_outputs[1434];
    assign outputs[742] = ~((layer4_outputs[2396]) & (layer4_outputs[1301]));
    assign outputs[743] = ~(layer4_outputs[2299]);
    assign outputs[744] = ~(layer4_outputs[797]);
    assign outputs[745] = (layer4_outputs[154]) & (layer4_outputs[513]);
    assign outputs[746] = ~(layer4_outputs[712]);
    assign outputs[747] = ~(layer4_outputs[931]) | (layer4_outputs[1271]);
    assign outputs[748] = ~(layer4_outputs[1782]);
    assign outputs[749] = layer4_outputs[1419];
    assign outputs[750] = (layer4_outputs[221]) ^ (layer4_outputs[2034]);
    assign outputs[751] = ~(layer4_outputs[96]);
    assign outputs[752] = ~(layer4_outputs[1133]);
    assign outputs[753] = ~(layer4_outputs[640]);
    assign outputs[754] = layer4_outputs[23];
    assign outputs[755] = layer4_outputs[703];
    assign outputs[756] = ~((layer4_outputs[1563]) ^ (layer4_outputs[1187]));
    assign outputs[757] = layer4_outputs[1572];
    assign outputs[758] = ~((layer4_outputs[2385]) | (layer4_outputs[1802]));
    assign outputs[759] = layer4_outputs[1164];
    assign outputs[760] = layer4_outputs[213];
    assign outputs[761] = ~(layer4_outputs[1753]);
    assign outputs[762] = ~(layer4_outputs[2380]);
    assign outputs[763] = ~(layer4_outputs[826]);
    assign outputs[764] = (layer4_outputs[963]) & ~(layer4_outputs[2447]);
    assign outputs[765] = ~(layer4_outputs[1829]);
    assign outputs[766] = (layer4_outputs[1936]) ^ (layer4_outputs[1731]);
    assign outputs[767] = layer4_outputs[377];
    assign outputs[768] = layer4_outputs[284];
    assign outputs[769] = layer4_outputs[1803];
    assign outputs[770] = layer4_outputs[709];
    assign outputs[771] = ~(layer4_outputs[143]);
    assign outputs[772] = layer4_outputs[854];
    assign outputs[773] = ~(layer4_outputs[2005]);
    assign outputs[774] = ~(layer4_outputs[2018]);
    assign outputs[775] = layer4_outputs[1078];
    assign outputs[776] = layer4_outputs[2228];
    assign outputs[777] = (layer4_outputs[1240]) | (layer4_outputs[2540]);
    assign outputs[778] = ~((layer4_outputs[1445]) ^ (layer4_outputs[1628]));
    assign outputs[779] = ~(layer4_outputs[1581]);
    assign outputs[780] = (layer4_outputs[816]) & ~(layer4_outputs[1851]);
    assign outputs[781] = (layer4_outputs[322]) & ~(layer4_outputs[400]);
    assign outputs[782] = ~(layer4_outputs[1866]);
    assign outputs[783] = ~(layer4_outputs[224]);
    assign outputs[784] = (layer4_outputs[617]) & ~(layer4_outputs[388]);
    assign outputs[785] = layer4_outputs[2061];
    assign outputs[786] = ~((layer4_outputs[605]) | (layer4_outputs[401]));
    assign outputs[787] = ~(layer4_outputs[1866]) | (layer4_outputs[108]);
    assign outputs[788] = layer4_outputs[39];
    assign outputs[789] = layer4_outputs[2048];
    assign outputs[790] = ~(layer4_outputs[525]);
    assign outputs[791] = layer4_outputs[235];
    assign outputs[792] = ~(layer4_outputs[1394]);
    assign outputs[793] = ~(layer4_outputs[92]);
    assign outputs[794] = ~(layer4_outputs[1637]);
    assign outputs[795] = layer4_outputs[1319];
    assign outputs[796] = (layer4_outputs[1200]) ^ (layer4_outputs[2256]);
    assign outputs[797] = ~(layer4_outputs[710]) | (layer4_outputs[1946]);
    assign outputs[798] = (layer4_outputs[2405]) & ~(layer4_outputs[924]);
    assign outputs[799] = ~((layer4_outputs[1908]) ^ (layer4_outputs[321]));
    assign outputs[800] = (layer4_outputs[1180]) ^ (layer4_outputs[421]);
    assign outputs[801] = (layer4_outputs[432]) | (layer4_outputs[285]);
    assign outputs[802] = layer4_outputs[1076];
    assign outputs[803] = ~(layer4_outputs[1787]);
    assign outputs[804] = (layer4_outputs[838]) & ~(layer4_outputs[625]);
    assign outputs[805] = (layer4_outputs[396]) & (layer4_outputs[195]);
    assign outputs[806] = layer4_outputs[472];
    assign outputs[807] = ~(layer4_outputs[1999]);
    assign outputs[808] = ~(layer4_outputs[2163]);
    assign outputs[809] = ~(layer4_outputs[358]);
    assign outputs[810] = (layer4_outputs[2520]) ^ (layer4_outputs[1253]);
    assign outputs[811] = ~(layer4_outputs[2082]);
    assign outputs[812] = layer4_outputs[927];
    assign outputs[813] = ~(layer4_outputs[1406]);
    assign outputs[814] = ~(layer4_outputs[37]);
    assign outputs[815] = ~((layer4_outputs[1416]) | (layer4_outputs[702]));
    assign outputs[816] = ~(layer4_outputs[1630]);
    assign outputs[817] = layer4_outputs[571];
    assign outputs[818] = layer4_outputs[2181];
    assign outputs[819] = ~((layer4_outputs[488]) | (layer4_outputs[1940]));
    assign outputs[820] = (layer4_outputs[1639]) & ~(layer4_outputs[1798]);
    assign outputs[821] = ~(layer4_outputs[1574]);
    assign outputs[822] = ~(layer4_outputs[1886]);
    assign outputs[823] = layer4_outputs[1198];
    assign outputs[824] = layer4_outputs[2193];
    assign outputs[825] = ~((layer4_outputs[1274]) ^ (layer4_outputs[708]));
    assign outputs[826] = ~(layer4_outputs[262]);
    assign outputs[827] = ~((layer4_outputs[314]) | (layer4_outputs[2444]));
    assign outputs[828] = layer4_outputs[1785];
    assign outputs[829] = layer4_outputs[2076];
    assign outputs[830] = ~(layer4_outputs[2256]);
    assign outputs[831] = layer4_outputs[1388];
    assign outputs[832] = layer4_outputs[2137];
    assign outputs[833] = ~(layer4_outputs[470]);
    assign outputs[834] = ~(layer4_outputs[491]) | (layer4_outputs[2326]);
    assign outputs[835] = layer4_outputs[453];
    assign outputs[836] = (layer4_outputs[420]) & ~(layer4_outputs[1658]);
    assign outputs[837] = layer4_outputs[2532];
    assign outputs[838] = layer4_outputs[1291];
    assign outputs[839] = ~(layer4_outputs[2050]);
    assign outputs[840] = ~((layer4_outputs[1596]) & (layer4_outputs[250]));
    assign outputs[841] = (layer4_outputs[907]) | (layer4_outputs[419]);
    assign outputs[842] = ~(layer4_outputs[1273]);
    assign outputs[843] = layer4_outputs[980];
    assign outputs[844] = layer4_outputs[618];
    assign outputs[845] = ~(layer4_outputs[49]);
    assign outputs[846] = ~(layer4_outputs[868]);
    assign outputs[847] = layer4_outputs[2117];
    assign outputs[848] = (layer4_outputs[2486]) & ~(layer4_outputs[2348]);
    assign outputs[849] = ~(layer4_outputs[231]);
    assign outputs[850] = ~(layer4_outputs[2246]);
    assign outputs[851] = ~(layer4_outputs[1105]);
    assign outputs[852] = ~(layer4_outputs[613]);
    assign outputs[853] = ~((layer4_outputs[2026]) ^ (layer4_outputs[2455]));
    assign outputs[854] = ~(layer4_outputs[233]);
    assign outputs[855] = ~((layer4_outputs[1397]) ^ (layer4_outputs[2320]));
    assign outputs[856] = layer4_outputs[2376];
    assign outputs[857] = ~(layer4_outputs[1353]);
    assign outputs[858] = ~(layer4_outputs[393]);
    assign outputs[859] = ~((layer4_outputs[310]) | (layer4_outputs[535]));
    assign outputs[860] = layer4_outputs[923];
    assign outputs[861] = ~(layer4_outputs[1152]);
    assign outputs[862] = ~((layer4_outputs[1602]) | (layer4_outputs[1630]));
    assign outputs[863] = layer4_outputs[434];
    assign outputs[864] = ~(layer4_outputs[1503]);
    assign outputs[865] = ~(layer4_outputs[874]);
    assign outputs[866] = ~(layer4_outputs[800]);
    assign outputs[867] = ~(layer4_outputs[491]);
    assign outputs[868] = layer4_outputs[109];
    assign outputs[869] = ~(layer4_outputs[1508]);
    assign outputs[870] = ~(layer4_outputs[1941]) | (layer4_outputs[515]);
    assign outputs[871] = ~(layer4_outputs[2536]);
    assign outputs[872] = ~((layer4_outputs[260]) | (layer4_outputs[2264]));
    assign outputs[873] = layer4_outputs[72];
    assign outputs[874] = ~(layer4_outputs[1293]);
    assign outputs[875] = ~(layer4_outputs[476]);
    assign outputs[876] = ~(layer4_outputs[520]);
    assign outputs[877] = layer4_outputs[473];
    assign outputs[878] = ~((layer4_outputs[1091]) ^ (layer4_outputs[2347]));
    assign outputs[879] = ~((layer4_outputs[1255]) ^ (layer4_outputs[365]));
    assign outputs[880] = ~(layer4_outputs[1084]);
    assign outputs[881] = ~((layer4_outputs[1598]) & (layer4_outputs[1161]));
    assign outputs[882] = layer4_outputs[1036];
    assign outputs[883] = layer4_outputs[1762];
    assign outputs[884] = (layer4_outputs[1312]) & (layer4_outputs[1042]);
    assign outputs[885] = ~(layer4_outputs[1386]);
    assign outputs[886] = layer4_outputs[359];
    assign outputs[887] = ~(layer4_outputs[1321]);
    assign outputs[888] = layer4_outputs[567];
    assign outputs[889] = ~(layer4_outputs[1813]);
    assign outputs[890] = ~(layer4_outputs[2369]);
    assign outputs[891] = (layer4_outputs[2411]) & (layer4_outputs[1041]);
    assign outputs[892] = layer4_outputs[1252];
    assign outputs[893] = layer4_outputs[661];
    assign outputs[894] = layer4_outputs[406];
    assign outputs[895] = ~(layer4_outputs[1465]);
    assign outputs[896] = ~(layer4_outputs[2485]);
    assign outputs[897] = ~((layer4_outputs[1726]) & (layer4_outputs[1072]));
    assign outputs[898] = ~(layer4_outputs[387]);
    assign outputs[899] = (layer4_outputs[1703]) & ~(layer4_outputs[1754]);
    assign outputs[900] = (layer4_outputs[1756]) ^ (layer4_outputs[952]);
    assign outputs[901] = ~(layer4_outputs[997]);
    assign outputs[902] = layer4_outputs[2372];
    assign outputs[903] = ~((layer4_outputs[1667]) | (layer4_outputs[801]));
    assign outputs[904] = ~(layer4_outputs[719]);
    assign outputs[905] = ~(layer4_outputs[2217]);
    assign outputs[906] = ~(layer4_outputs[1111]);
    assign outputs[907] = ~(layer4_outputs[1300]) | (layer4_outputs[2149]);
    assign outputs[908] = layer4_outputs[1473];
    assign outputs[909] = ~(layer4_outputs[1194]);
    assign outputs[910] = (layer4_outputs[2223]) & ~(layer4_outputs[1697]);
    assign outputs[911] = ~(layer4_outputs[410]);
    assign outputs[912] = (layer4_outputs[2184]) & ~(layer4_outputs[330]);
    assign outputs[913] = layer4_outputs[1500];
    assign outputs[914] = ~(layer4_outputs[218]);
    assign outputs[915] = (layer4_outputs[222]) & ~(layer4_outputs[1472]);
    assign outputs[916] = layer4_outputs[1481];
    assign outputs[917] = layer4_outputs[2171];
    assign outputs[918] = ~(layer4_outputs[635]);
    assign outputs[919] = ~(layer4_outputs[2518]);
    assign outputs[920] = (layer4_outputs[1143]) & (layer4_outputs[1059]);
    assign outputs[921] = ~(layer4_outputs[1206]);
    assign outputs[922] = ~(layer4_outputs[1991]);
    assign outputs[923] = layer4_outputs[730];
    assign outputs[924] = ~((layer4_outputs[1028]) ^ (layer4_outputs[1273]));
    assign outputs[925] = ~(layer4_outputs[1120]) | (layer4_outputs[559]);
    assign outputs[926] = ~((layer4_outputs[1162]) & (layer4_outputs[368]));
    assign outputs[927] = layer4_outputs[374];
    assign outputs[928] = ~(layer4_outputs[2270]);
    assign outputs[929] = (layer4_outputs[87]) ^ (layer4_outputs[1123]);
    assign outputs[930] = layer4_outputs[15];
    assign outputs[931] = ~(layer4_outputs[882]);
    assign outputs[932] = layer4_outputs[1825];
    assign outputs[933] = layer4_outputs[1599];
    assign outputs[934] = layer4_outputs[2020];
    assign outputs[935] = layer4_outputs[714];
    assign outputs[936] = layer4_outputs[1641];
    assign outputs[937] = (layer4_outputs[1428]) ^ (layer4_outputs[1717]);
    assign outputs[938] = layer4_outputs[2430];
    assign outputs[939] = layer4_outputs[151];
    assign outputs[940] = ~(layer4_outputs[2107]);
    assign outputs[941] = layer4_outputs[364];
    assign outputs[942] = (layer4_outputs[1498]) & ~(layer4_outputs[1432]);
    assign outputs[943] = (layer4_outputs[2332]) & (layer4_outputs[2435]);
    assign outputs[944] = layer4_outputs[889];
    assign outputs[945] = ~(layer4_outputs[1777]);
    assign outputs[946] = ~((layer4_outputs[898]) ^ (layer4_outputs[972]));
    assign outputs[947] = layer4_outputs[1281];
    assign outputs[948] = ~(layer4_outputs[1467]);
    assign outputs[949] = (layer4_outputs[1550]) | (layer4_outputs[988]);
    assign outputs[950] = ~(layer4_outputs[1171]);
    assign outputs[951] = (layer4_outputs[1898]) & ~(layer4_outputs[2294]);
    assign outputs[952] = layer4_outputs[561];
    assign outputs[953] = ~(layer4_outputs[89]);
    assign outputs[954] = layer4_outputs[2019];
    assign outputs[955] = ~(layer4_outputs[1134]);
    assign outputs[956] = ~(layer4_outputs[2054]);
    assign outputs[957] = (layer4_outputs[2027]) | (layer4_outputs[285]);
    assign outputs[958] = layer4_outputs[345];
    assign outputs[959] = ~(layer4_outputs[706]);
    assign outputs[960] = ~(layer4_outputs[968]);
    assign outputs[961] = (layer4_outputs[673]) | (layer4_outputs[479]);
    assign outputs[962] = ~(layer4_outputs[1687]);
    assign outputs[963] = layer4_outputs[2044];
    assign outputs[964] = layer4_outputs[923];
    assign outputs[965] = ~(layer4_outputs[229]);
    assign outputs[966] = (layer4_outputs[2012]) & ~(layer4_outputs[152]);
    assign outputs[967] = ~(layer4_outputs[372]);
    assign outputs[968] = ~(layer4_outputs[1106]);
    assign outputs[969] = ~(layer4_outputs[2551]);
    assign outputs[970] = layer4_outputs[1985];
    assign outputs[971] = layer4_outputs[63];
    assign outputs[972] = (layer4_outputs[1360]) & ~(layer4_outputs[941]);
    assign outputs[973] = layer4_outputs[2325];
    assign outputs[974] = layer4_outputs[2181];
    assign outputs[975] = ~(layer4_outputs[330]) | (layer4_outputs[803]);
    assign outputs[976] = layer4_outputs[884];
    assign outputs[977] = ~(layer4_outputs[768]);
    assign outputs[978] = ~(layer4_outputs[528]);
    assign outputs[979] = layer4_outputs[1123];
    assign outputs[980] = (layer4_outputs[596]) & (layer4_outputs[838]);
    assign outputs[981] = ~((layer4_outputs[917]) ^ (layer4_outputs[2021]));
    assign outputs[982] = layer4_outputs[779];
    assign outputs[983] = (layer4_outputs[2559]) & (layer4_outputs[2340]);
    assign outputs[984] = layer4_outputs[598];
    assign outputs[985] = ~(layer4_outputs[1099]);
    assign outputs[986] = ~(layer4_outputs[263]);
    assign outputs[987] = (layer4_outputs[1410]) & ~(layer4_outputs[776]);
    assign outputs[988] = (layer4_outputs[420]) & ~(layer4_outputs[1083]);
    assign outputs[989] = layer4_outputs[950];
    assign outputs[990] = layer4_outputs[2124];
    assign outputs[991] = ~(layer4_outputs[1111]);
    assign outputs[992] = ~(layer4_outputs[1588]);
    assign outputs[993] = (layer4_outputs[1727]) & (layer4_outputs[422]);
    assign outputs[994] = ~(layer4_outputs[2524]);
    assign outputs[995] = (layer4_outputs[707]) & (layer4_outputs[764]);
    assign outputs[996] = (layer4_outputs[1918]) & ~(layer4_outputs[1107]);
    assign outputs[997] = ~(layer4_outputs[1671]);
    assign outputs[998] = (layer4_outputs[2237]) ^ (layer4_outputs[803]);
    assign outputs[999] = layer4_outputs[1779];
    assign outputs[1000] = layer4_outputs[22];
    assign outputs[1001] = layer4_outputs[816];
    assign outputs[1002] = layer4_outputs[157];
    assign outputs[1003] = layer4_outputs[1652];
    assign outputs[1004] = ~(layer4_outputs[523]);
    assign outputs[1005] = ~(layer4_outputs[143]);
    assign outputs[1006] = ~(layer4_outputs[1901]);
    assign outputs[1007] = ~(layer4_outputs[2308]);
    assign outputs[1008] = ~(layer4_outputs[203]);
    assign outputs[1009] = ~(layer4_outputs[234]);
    assign outputs[1010] = layer4_outputs[779];
    assign outputs[1011] = ~(layer4_outputs[909]);
    assign outputs[1012] = layer4_outputs[959];
    assign outputs[1013] = layer4_outputs[2499];
    assign outputs[1014] = (layer4_outputs[438]) & ~(layer4_outputs[2189]);
    assign outputs[1015] = layer4_outputs[2128];
    assign outputs[1016] = ~(layer4_outputs[2002]);
    assign outputs[1017] = ~((layer4_outputs[2179]) ^ (layer4_outputs[671]));
    assign outputs[1018] = layer4_outputs[561];
    assign outputs[1019] = (layer4_outputs[243]) ^ (layer4_outputs[1801]);
    assign outputs[1020] = ~(layer4_outputs[2353]);
    assign outputs[1021] = ~((layer4_outputs[601]) | (layer4_outputs[1962]));
    assign outputs[1022] = ~((layer4_outputs[2356]) ^ (layer4_outputs[59]));
    assign outputs[1023] = ~(layer4_outputs[805]);
    assign outputs[1024] = ~(layer4_outputs[464]);
    assign outputs[1025] = ~(layer4_outputs[142]);
    assign outputs[1026] = layer4_outputs[2133];
    assign outputs[1027] = ~(layer4_outputs[2304]);
    assign outputs[1028] = ~((layer4_outputs[2342]) ^ (layer4_outputs[2274]));
    assign outputs[1029] = (layer4_outputs[1631]) ^ (layer4_outputs[2542]);
    assign outputs[1030] = (layer4_outputs[422]) & ~(layer4_outputs[1702]);
    assign outputs[1031] = ~(layer4_outputs[2254]);
    assign outputs[1032] = ~(layer4_outputs[2100]);
    assign outputs[1033] = layer4_outputs[734];
    assign outputs[1034] = layer4_outputs[1417];
    assign outputs[1035] = layer4_outputs[117];
    assign outputs[1036] = (layer4_outputs[1908]) & ~(layer4_outputs[974]);
    assign outputs[1037] = ~((layer4_outputs[1495]) ^ (layer4_outputs[1656]));
    assign outputs[1038] = ~(layer4_outputs[544]) | (layer4_outputs[994]);
    assign outputs[1039] = layer4_outputs[1485];
    assign outputs[1040] = ~(layer4_outputs[1863]);
    assign outputs[1041] = (layer4_outputs[1421]) & (layer4_outputs[1239]);
    assign outputs[1042] = layer4_outputs[1910];
    assign outputs[1043] = ~(layer4_outputs[17]) | (layer4_outputs[2191]);
    assign outputs[1044] = layer4_outputs[2307];
    assign outputs[1045] = ~(layer4_outputs[480]);
    assign outputs[1046] = layer4_outputs[350];
    assign outputs[1047] = ~((layer4_outputs[265]) ^ (layer4_outputs[1518]));
    assign outputs[1048] = (layer4_outputs[1073]) & ~(layer4_outputs[1480]);
    assign outputs[1049] = ~((layer4_outputs[94]) | (layer4_outputs[873]));
    assign outputs[1050] = (layer4_outputs[667]) & (layer4_outputs[1890]);
    assign outputs[1051] = layer4_outputs[879];
    assign outputs[1052] = ~((layer4_outputs[547]) | (layer4_outputs[939]));
    assign outputs[1053] = layer4_outputs[1996];
    assign outputs[1054] = ~(layer4_outputs[761]);
    assign outputs[1055] = ~(layer4_outputs[1056]);
    assign outputs[1056] = ~(layer4_outputs[1754]);
    assign outputs[1057] = layer4_outputs[482];
    assign outputs[1058] = (layer4_outputs[2183]) & (layer4_outputs[1455]);
    assign outputs[1059] = (layer4_outputs[2330]) & (layer4_outputs[1734]);
    assign outputs[1060] = (layer4_outputs[58]) & ~(layer4_outputs[1746]);
    assign outputs[1061] = layer4_outputs[215];
    assign outputs[1062] = (layer4_outputs[1254]) & ~(layer4_outputs[1033]);
    assign outputs[1063] = ~(layer4_outputs[1451]);
    assign outputs[1064] = (layer4_outputs[573]) & ~(layer4_outputs[2109]);
    assign outputs[1065] = (layer4_outputs[748]) & ~(layer4_outputs[344]);
    assign outputs[1066] = layer4_outputs[264];
    assign outputs[1067] = layer4_outputs[2406];
    assign outputs[1068] = layer4_outputs[650];
    assign outputs[1069] = layer4_outputs[220];
    assign outputs[1070] = layer4_outputs[1884];
    assign outputs[1071] = layer4_outputs[53];
    assign outputs[1072] = layer4_outputs[246];
    assign outputs[1073] = layer4_outputs[751];
    assign outputs[1074] = ~(layer4_outputs[2135]);
    assign outputs[1075] = layer4_outputs[2185];
    assign outputs[1076] = ~(layer4_outputs[216]) | (layer4_outputs[890]);
    assign outputs[1077] = ~(layer4_outputs[891]);
    assign outputs[1078] = ~(layer4_outputs[1527]);
    assign outputs[1079] = ~((layer4_outputs[411]) | (layer4_outputs[2376]));
    assign outputs[1080] = layer4_outputs[2102];
    assign outputs[1081] = ~(layer4_outputs[1296]);
    assign outputs[1082] = ~(layer4_outputs[1341]);
    assign outputs[1083] = layer4_outputs[942];
    assign outputs[1084] = (layer4_outputs[1966]) | (layer4_outputs[88]);
    assign outputs[1085] = layer4_outputs[1648];
    assign outputs[1086] = layer4_outputs[886];
    assign outputs[1087] = layer4_outputs[1659];
    assign outputs[1088] = layer4_outputs[1665];
    assign outputs[1089] = layer4_outputs[149];
    assign outputs[1090] = layer4_outputs[105];
    assign outputs[1091] = layer4_outputs[1679];
    assign outputs[1092] = ~(layer4_outputs[806]) | (layer4_outputs[1884]);
    assign outputs[1093] = layer4_outputs[886];
    assign outputs[1094] = (layer4_outputs[1561]) & (layer4_outputs[124]);
    assign outputs[1095] = layer4_outputs[1531];
    assign outputs[1096] = layer4_outputs[1560];
    assign outputs[1097] = layer4_outputs[973];
    assign outputs[1098] = layer4_outputs[2126];
    assign outputs[1099] = layer4_outputs[482];
    assign outputs[1100] = ~(layer4_outputs[682]);
    assign outputs[1101] = layer4_outputs[896];
    assign outputs[1102] = ~(layer4_outputs[2395]);
    assign outputs[1103] = ~(layer4_outputs[1706]) | (layer4_outputs[2176]);
    assign outputs[1104] = layer4_outputs[703];
    assign outputs[1105] = ~((layer4_outputs[2043]) ^ (layer4_outputs[1113]));
    assign outputs[1106] = ~(layer4_outputs[1808]);
    assign outputs[1107] = (layer4_outputs[2534]) & ~(layer4_outputs[1354]);
    assign outputs[1108] = ~(layer4_outputs[1553]);
    assign outputs[1109] = ~((layer4_outputs[1230]) | (layer4_outputs[370]));
    assign outputs[1110] = layer4_outputs[775];
    assign outputs[1111] = (layer4_outputs[1533]) ^ (layer4_outputs[626]);
    assign outputs[1112] = (layer4_outputs[123]) & (layer4_outputs[901]);
    assign outputs[1113] = ~((layer4_outputs[81]) ^ (layer4_outputs[1088]));
    assign outputs[1114] = layer4_outputs[664];
    assign outputs[1115] = ~(layer4_outputs[2226]);
    assign outputs[1116] = ~((layer4_outputs[531]) ^ (layer4_outputs[1193]));
    assign outputs[1117] = ~(layer4_outputs[390]);
    assign outputs[1118] = (layer4_outputs[502]) ^ (layer4_outputs[2281]);
    assign outputs[1119] = layer4_outputs[1466];
    assign outputs[1120] = ~((layer4_outputs[1647]) | (layer4_outputs[2292]));
    assign outputs[1121] = layer4_outputs[228];
    assign outputs[1122] = (layer4_outputs[2058]) & ~(layer4_outputs[1719]);
    assign outputs[1123] = (layer4_outputs[2047]) & (layer4_outputs[1009]);
    assign outputs[1124] = layer4_outputs[541];
    assign outputs[1125] = (layer4_outputs[1535]) & ~(layer4_outputs[2334]);
    assign outputs[1126] = ~(layer4_outputs[2334]);
    assign outputs[1127] = layer4_outputs[701];
    assign outputs[1128] = layer4_outputs[1687];
    assign outputs[1129] = ~(layer4_outputs[1060]);
    assign outputs[1130] = ~((layer4_outputs[220]) ^ (layer4_outputs[1976]));
    assign outputs[1131] = layer4_outputs[139];
    assign outputs[1132] = ~((layer4_outputs[539]) | (layer4_outputs[678]));
    assign outputs[1133] = (layer4_outputs[1689]) ^ (layer4_outputs[198]);
    assign outputs[1134] = (layer4_outputs[2558]) & ~(layer4_outputs[164]);
    assign outputs[1135] = layer4_outputs[366];
    assign outputs[1136] = ~((layer4_outputs[2132]) ^ (layer4_outputs[104]));
    assign outputs[1137] = ~(layer4_outputs[2487]);
    assign outputs[1138] = layer4_outputs[1054];
    assign outputs[1139] = ~(layer4_outputs[1612]);
    assign outputs[1140] = ~(layer4_outputs[999]);
    assign outputs[1141] = layer4_outputs[928];
    assign outputs[1142] = ~((layer4_outputs[1047]) | (layer4_outputs[2552]));
    assign outputs[1143] = ~(layer4_outputs[1556]);
    assign outputs[1144] = ~(layer4_outputs[1998]);
    assign outputs[1145] = layer4_outputs[1669];
    assign outputs[1146] = (layer4_outputs[1641]) ^ (layer4_outputs[477]);
    assign outputs[1147] = ~(layer4_outputs[1992]);
    assign outputs[1148] = layer4_outputs[442];
    assign outputs[1149] = layer4_outputs[753];
    assign outputs[1150] = layer4_outputs[1202];
    assign outputs[1151] = ~((layer4_outputs[1799]) & (layer4_outputs[2446]));
    assign outputs[1152] = ~(layer4_outputs[579]) | (layer4_outputs[1309]);
    assign outputs[1153] = (layer4_outputs[2215]) & ~(layer4_outputs[1909]);
    assign outputs[1154] = ~(layer4_outputs[458]);
    assign outputs[1155] = layer4_outputs[672];
    assign outputs[1156] = layer4_outputs[1406];
    assign outputs[1157] = (layer4_outputs[2389]) & ~(layer4_outputs[2549]);
    assign outputs[1158] = ~(layer4_outputs[245]);
    assign outputs[1159] = (layer4_outputs[278]) ^ (layer4_outputs[2519]);
    assign outputs[1160] = layer4_outputs[2281];
    assign outputs[1161] = layer4_outputs[5];
    assign outputs[1162] = ~(layer4_outputs[1892]);
    assign outputs[1163] = ~(layer4_outputs[2129]);
    assign outputs[1164] = layer4_outputs[634];
    assign outputs[1165] = (layer4_outputs[2337]) ^ (layer4_outputs[1208]);
    assign outputs[1166] = layer4_outputs[75];
    assign outputs[1167] = ~((layer4_outputs[181]) ^ (layer4_outputs[249]));
    assign outputs[1168] = ~((layer4_outputs[1064]) ^ (layer4_outputs[2496]));
    assign outputs[1169] = ~(layer4_outputs[1258]);
    assign outputs[1170] = ~(layer4_outputs[2108]);
    assign outputs[1171] = ~((layer4_outputs[2109]) & (layer4_outputs[1558]));
    assign outputs[1172] = layer4_outputs[674];
    assign outputs[1173] = (layer4_outputs[2530]) & ~(layer4_outputs[195]);
    assign outputs[1174] = layer4_outputs[1645];
    assign outputs[1175] = (layer4_outputs[2114]) & ~(layer4_outputs[2425]);
    assign outputs[1176] = layer4_outputs[752];
    assign outputs[1177] = ~(layer4_outputs[113]);
    assign outputs[1178] = ~(layer4_outputs[1834]);
    assign outputs[1179] = (layer4_outputs[1486]) & (layer4_outputs[1489]);
    assign outputs[1180] = (layer4_outputs[1566]) & ~(layer4_outputs[1810]);
    assign outputs[1181] = ~((layer4_outputs[1129]) | (layer4_outputs[1227]));
    assign outputs[1182] = ~(layer4_outputs[1881]);
    assign outputs[1183] = layer4_outputs[932];
    assign outputs[1184] = layer4_outputs[2515];
    assign outputs[1185] = ~(layer4_outputs[1258]);
    assign outputs[1186] = ~(layer4_outputs[1538]);
    assign outputs[1187] = ~(layer4_outputs[1282]);
    assign outputs[1188] = ~((layer4_outputs[2218]) ^ (layer4_outputs[369]));
    assign outputs[1189] = (layer4_outputs[1133]) ^ (layer4_outputs[235]);
    assign outputs[1190] = layer4_outputs[1521];
    assign outputs[1191] = ~((layer4_outputs[2245]) ^ (layer4_outputs[332]));
    assign outputs[1192] = ~(layer4_outputs[1449]);
    assign outputs[1193] = ~(layer4_outputs[1172]);
    assign outputs[1194] = ~(layer4_outputs[1913]);
    assign outputs[1195] = (layer4_outputs[2368]) ^ (layer4_outputs[1968]);
    assign outputs[1196] = (layer4_outputs[984]) ^ (layer4_outputs[2051]);
    assign outputs[1197] = ~(layer4_outputs[1401]);
    assign outputs[1198] = layer4_outputs[21];
    assign outputs[1199] = (layer4_outputs[258]) ^ (layer4_outputs[876]);
    assign outputs[1200] = (layer4_outputs[1526]) & (layer4_outputs[1392]);
    assign outputs[1201] = ~(layer4_outputs[1522]);
    assign outputs[1202] = ~(layer4_outputs[1820]);
    assign outputs[1203] = layer4_outputs[2420];
    assign outputs[1204] = (layer4_outputs[415]) & ~(layer4_outputs[1188]);
    assign outputs[1205] = ~(layer4_outputs[930]);
    assign outputs[1206] = layer4_outputs[1962];
    assign outputs[1207] = ~(layer4_outputs[2506]);
    assign outputs[1208] = ~((layer4_outputs[34]) | (layer4_outputs[1062]));
    assign outputs[1209] = (layer4_outputs[2544]) & ~(layer4_outputs[1345]);
    assign outputs[1210] = ~(layer4_outputs[370]);
    assign outputs[1211] = layer4_outputs[2329];
    assign outputs[1212] = (layer4_outputs[1287]) & ~(layer4_outputs[162]);
    assign outputs[1213] = (layer4_outputs[481]) ^ (layer4_outputs[1824]);
    assign outputs[1214] = layer4_outputs[615];
    assign outputs[1215] = layer4_outputs[469];
    assign outputs[1216] = layer4_outputs[2528];
    assign outputs[1217] = (layer4_outputs[2008]) & ~(layer4_outputs[159]);
    assign outputs[1218] = layer4_outputs[735];
    assign outputs[1219] = ~(layer4_outputs[2163]) | (layer4_outputs[2210]);
    assign outputs[1220] = layer4_outputs[1295];
    assign outputs[1221] = ~(layer4_outputs[2231]);
    assign outputs[1222] = (layer4_outputs[585]) & ~(layer4_outputs[2285]);
    assign outputs[1223] = layer4_outputs[1514];
    assign outputs[1224] = ~(layer4_outputs[941]) | (layer4_outputs[1435]);
    assign outputs[1225] = ~(layer4_outputs[1158]);
    assign outputs[1226] = layer4_outputs[1105];
    assign outputs[1227] = layer4_outputs[1478];
    assign outputs[1228] = layer4_outputs[2428];
    assign outputs[1229] = layer4_outputs[192];
    assign outputs[1230] = ~(layer4_outputs[1323]);
    assign outputs[1231] = (layer4_outputs[750]) & ~(layer4_outputs[602]);
    assign outputs[1232] = (layer4_outputs[311]) & (layer4_outputs[2240]);
    assign outputs[1233] = ~((layer4_outputs[2207]) | (layer4_outputs[1468]));
    assign outputs[1234] = ~(layer4_outputs[2123]);
    assign outputs[1235] = layer4_outputs[1784];
    assign outputs[1236] = ~((layer4_outputs[1170]) ^ (layer4_outputs[1879]));
    assign outputs[1237] = layer4_outputs[318];
    assign outputs[1238] = ~(layer4_outputs[1832]);
    assign outputs[1239] = ~((layer4_outputs[2451]) ^ (layer4_outputs[1193]));
    assign outputs[1240] = ~(layer4_outputs[1370]);
    assign outputs[1241] = ~(layer4_outputs[1609]);
    assign outputs[1242] = ~(layer4_outputs[1616]);
    assign outputs[1243] = layer4_outputs[2295];
    assign outputs[1244] = (layer4_outputs[743]) & ~(layer4_outputs[2536]);
    assign outputs[1245] = ~(layer4_outputs[666]);
    assign outputs[1246] = ~(layer4_outputs[279]);
    assign outputs[1247] = (layer4_outputs[719]) & ~(layer4_outputs[2070]);
    assign outputs[1248] = layer4_outputs[105];
    assign outputs[1249] = ~(layer4_outputs[2077]);
    assign outputs[1250] = layer4_outputs[634];
    assign outputs[1251] = ~((layer4_outputs[81]) | (layer4_outputs[977]));
    assign outputs[1252] = layer4_outputs[1653];
    assign outputs[1253] = layer4_outputs[1301];
    assign outputs[1254] = ~(layer4_outputs[531]);
    assign outputs[1255] = ~(layer4_outputs[1512]);
    assign outputs[1256] = layer4_outputs[1819];
    assign outputs[1257] = ~(layer4_outputs[562]);
    assign outputs[1258] = ~((layer4_outputs[1082]) ^ (layer4_outputs[312]));
    assign outputs[1259] = ~(layer4_outputs[532]);
    assign outputs[1260] = ~((layer4_outputs[1336]) | (layer4_outputs[2467]));
    assign outputs[1261] = (layer4_outputs[2427]) & ~(layer4_outputs[274]);
    assign outputs[1262] = ~(layer4_outputs[1624]);
    assign outputs[1263] = ~(layer4_outputs[1829]);
    assign outputs[1264] = (layer4_outputs[19]) & (layer4_outputs[54]);
    assign outputs[1265] = ~(layer4_outputs[1262]);
    assign outputs[1266] = ~(layer4_outputs[712]);
    assign outputs[1267] = (layer4_outputs[992]) & ~(layer4_outputs[2233]);
    assign outputs[1268] = layer4_outputs[736];
    assign outputs[1269] = (layer4_outputs[2016]) & ~(layer4_outputs[436]);
    assign outputs[1270] = ~((layer4_outputs[2397]) ^ (layer4_outputs[350]));
    assign outputs[1271] = layer4_outputs[1566];
    assign outputs[1272] = layer4_outputs[1368];
    assign outputs[1273] = ~(layer4_outputs[2303]);
    assign outputs[1274] = ~(layer4_outputs[1977]);
    assign outputs[1275] = (layer4_outputs[638]) & ~(layer4_outputs[338]);
    assign outputs[1276] = (layer4_outputs[1009]) & (layer4_outputs[2058]);
    assign outputs[1277] = ~(layer4_outputs[2412]);
    assign outputs[1278] = (layer4_outputs[339]) ^ (layer4_outputs[397]);
    assign outputs[1279] = layer4_outputs[61];
    assign outputs[1280] = layer4_outputs[1516];
    assign outputs[1281] = ~((layer4_outputs[1312]) | (layer4_outputs[1940]));
    assign outputs[1282] = layer4_outputs[371];
    assign outputs[1283] = layer4_outputs[1732];
    assign outputs[1284] = (layer4_outputs[729]) & (layer4_outputs[871]);
    assign outputs[1285] = ~(layer4_outputs[1601]);
    assign outputs[1286] = ~(layer4_outputs[1534]) | (layer4_outputs[650]);
    assign outputs[1287] = ~((layer4_outputs[140]) ^ (layer4_outputs[396]));
    assign outputs[1288] = layer4_outputs[570];
    assign outputs[1289] = layer4_outputs[381];
    assign outputs[1290] = ~(layer4_outputs[1626]);
    assign outputs[1291] = (layer4_outputs[1053]) & (layer4_outputs[1]);
    assign outputs[1292] = (layer4_outputs[1646]) & ~(layer4_outputs[2431]);
    assign outputs[1293] = (layer4_outputs[2449]) & (layer4_outputs[580]);
    assign outputs[1294] = ~(layer4_outputs[2290]);
    assign outputs[1295] = ~(layer4_outputs[1045]);
    assign outputs[1296] = layer4_outputs[1608];
    assign outputs[1297] = layer4_outputs[877];
    assign outputs[1298] = ~(layer4_outputs[558]);
    assign outputs[1299] = layer4_outputs[1467];
    assign outputs[1300] = ~(layer4_outputs[497]);
    assign outputs[1301] = ~(layer4_outputs[2270]);
    assign outputs[1302] = ~(layer4_outputs[1019]);
    assign outputs[1303] = layer4_outputs[182];
    assign outputs[1304] = layer4_outputs[552];
    assign outputs[1305] = (layer4_outputs[1330]) ^ (layer4_outputs[822]);
    assign outputs[1306] = layer4_outputs[1981];
    assign outputs[1307] = (layer4_outputs[1381]) & ~(layer4_outputs[349]);
    assign outputs[1308] = ~((layer4_outputs[1113]) | (layer4_outputs[908]));
    assign outputs[1309] = (layer4_outputs[2060]) & ~(layer4_outputs[942]);
    assign outputs[1310] = ~(layer4_outputs[256]);
    assign outputs[1311] = layer4_outputs[1704];
    assign outputs[1312] = ~(layer4_outputs[209]);
    assign outputs[1313] = ~(layer4_outputs[490]);
    assign outputs[1314] = (layer4_outputs[2101]) & (layer4_outputs[1550]);
    assign outputs[1315] = ~(layer4_outputs[1266]);
    assign outputs[1316] = ~(layer4_outputs[1769]);
    assign outputs[1317] = ~((layer4_outputs[72]) | (layer4_outputs[781]));
    assign outputs[1318] = layer4_outputs[649];
    assign outputs[1319] = (layer4_outputs[118]) & ~(layer4_outputs[1067]);
    assign outputs[1320] = ~((layer4_outputs[1857]) | (layer4_outputs[400]));
    assign outputs[1321] = ~(layer4_outputs[1879]);
    assign outputs[1322] = (layer4_outputs[1388]) ^ (layer4_outputs[2040]);
    assign outputs[1323] = (layer4_outputs[2450]) | (layer4_outputs[1007]);
    assign outputs[1324] = ~(layer4_outputs[500]);
    assign outputs[1325] = layer4_outputs[2418];
    assign outputs[1326] = (layer4_outputs[588]) & (layer4_outputs[1131]);
    assign outputs[1327] = ~(layer4_outputs[1210]);
    assign outputs[1328] = layer4_outputs[681];
    assign outputs[1329] = layer4_outputs[412];
    assign outputs[1330] = ~(layer4_outputs[1480]);
    assign outputs[1331] = layer4_outputs[505];
    assign outputs[1332] = ~(layer4_outputs[99]);
    assign outputs[1333] = layer4_outputs[1003];
    assign outputs[1334] = ~((layer4_outputs[1537]) ^ (layer4_outputs[928]));
    assign outputs[1335] = ~(layer4_outputs[144]);
    assign outputs[1336] = ~(layer4_outputs[1804]);
    assign outputs[1337] = layer4_outputs[810];
    assign outputs[1338] = layer4_outputs[1760];
    assign outputs[1339] = ~(layer4_outputs[1152]);
    assign outputs[1340] = layer4_outputs[586];
    assign outputs[1341] = ~(layer4_outputs[451]);
    assign outputs[1342] = ~(layer4_outputs[2265]);
    assign outputs[1343] = (layer4_outputs[2271]) | (layer4_outputs[1861]);
    assign outputs[1344] = ~((layer4_outputs[2306]) | (layer4_outputs[1081]));
    assign outputs[1345] = ~((layer4_outputs[208]) ^ (layer4_outputs[1242]));
    assign outputs[1346] = ~(layer4_outputs[174]) | (layer4_outputs[895]);
    assign outputs[1347] = layer4_outputs[2452];
    assign outputs[1348] = ~(layer4_outputs[1765]);
    assign outputs[1349] = ~(layer4_outputs[724]);
    assign outputs[1350] = ~((layer4_outputs[1114]) | (layer4_outputs[2196]));
    assign outputs[1351] = layer4_outputs[31];
    assign outputs[1352] = layer4_outputs[925];
    assign outputs[1353] = (layer4_outputs[2543]) | (layer4_outputs[1153]);
    assign outputs[1354] = ~(layer4_outputs[1670]);
    assign outputs[1355] = ~(layer4_outputs[2171]);
    assign outputs[1356] = ~(layer4_outputs[949]);
    assign outputs[1357] = (layer4_outputs[955]) ^ (layer4_outputs[2173]);
    assign outputs[1358] = ~((layer4_outputs[1654]) ^ (layer4_outputs[1013]));
    assign outputs[1359] = layer4_outputs[2206];
    assign outputs[1360] = layer4_outputs[1855];
    assign outputs[1361] = layer4_outputs[66];
    assign outputs[1362] = layer4_outputs[1531];
    assign outputs[1363] = (layer4_outputs[2482]) & ~(layer4_outputs[301]);
    assign outputs[1364] = ~(layer4_outputs[37]);
    assign outputs[1365] = ~(layer4_outputs[918]);
    assign outputs[1366] = layer4_outputs[557];
    assign outputs[1367] = layer4_outputs[1148];
    assign outputs[1368] = ~((layer4_outputs[581]) | (layer4_outputs[392]));
    assign outputs[1369] = layer4_outputs[340];
    assign outputs[1370] = ~(layer4_outputs[188]) | (layer4_outputs[2499]);
    assign outputs[1371] = ~((layer4_outputs[691]) ^ (layer4_outputs[455]));
    assign outputs[1372] = layer4_outputs[1484];
    assign outputs[1373] = ~(layer4_outputs[1137]);
    assign outputs[1374] = layer4_outputs[2372];
    assign outputs[1375] = ~((layer4_outputs[1313]) & (layer4_outputs[1401]));
    assign outputs[1376] = layer4_outputs[1794];
    assign outputs[1377] = ~(layer4_outputs[1733]);
    assign outputs[1378] = ~(layer4_outputs[1079]);
    assign outputs[1379] = (layer4_outputs[229]) & (layer4_outputs[230]);
    assign outputs[1380] = (layer4_outputs[1730]) & (layer4_outputs[2152]);
    assign outputs[1381] = (layer4_outputs[2249]) & (layer4_outputs[279]);
    assign outputs[1382] = (layer4_outputs[2]) & (layer4_outputs[689]);
    assign outputs[1383] = (layer4_outputs[1297]) & ~(layer4_outputs[352]);
    assign outputs[1384] = (layer4_outputs[777]) & (layer4_outputs[2543]);
    assign outputs[1385] = layer4_outputs[2083];
    assign outputs[1386] = (layer4_outputs[2122]) & ~(layer4_outputs[757]);
    assign outputs[1387] = ~(layer4_outputs[2010]);
    assign outputs[1388] = layer4_outputs[1993];
    assign outputs[1389] = layer4_outputs[666];
    assign outputs[1390] = ~(layer4_outputs[659]);
    assign outputs[1391] = ~(layer4_outputs[2195]);
    assign outputs[1392] = layer4_outputs[96];
    assign outputs[1393] = ~((layer4_outputs[1049]) ^ (layer4_outputs[1675]));
    assign outputs[1394] = layer4_outputs[2039];
    assign outputs[1395] = ~(layer4_outputs[690]);
    assign outputs[1396] = ~(layer4_outputs[533]);
    assign outputs[1397] = layer4_outputs[2039];
    assign outputs[1398] = ~(layer4_outputs[1720]);
    assign outputs[1399] = layer4_outputs[790];
    assign outputs[1400] = (layer4_outputs[351]) ^ (layer4_outputs[508]);
    assign outputs[1401] = (layer4_outputs[1824]) ^ (layer4_outputs[1475]);
    assign outputs[1402] = (layer4_outputs[875]) ^ (layer4_outputs[373]);
    assign outputs[1403] = ~(layer4_outputs[1246]);
    assign outputs[1404] = ~(layer4_outputs[361]);
    assign outputs[1405] = layer4_outputs[1575];
    assign outputs[1406] = (layer4_outputs[508]) & (layer4_outputs[1148]);
    assign outputs[1407] = layer4_outputs[524];
    assign outputs[1408] = ~(layer4_outputs[725]);
    assign outputs[1409] = ~(layer4_outputs[1015]) | (layer4_outputs[274]);
    assign outputs[1410] = layer4_outputs[1393];
    assign outputs[1411] = ~((layer4_outputs[489]) | (layer4_outputs[714]));
    assign outputs[1412] = (layer4_outputs[2174]) & ~(layer4_outputs[971]);
    assign outputs[1413] = ~(layer4_outputs[744]);
    assign outputs[1414] = layer4_outputs[1848];
    assign outputs[1415] = (layer4_outputs[1324]) & ~(layer4_outputs[439]);
    assign outputs[1416] = ~((layer4_outputs[1917]) ^ (layer4_outputs[856]));
    assign outputs[1417] = layer4_outputs[1931];
    assign outputs[1418] = layer4_outputs[2187];
    assign outputs[1419] = ~(layer4_outputs[238]);
    assign outputs[1420] = ~(layer4_outputs[620]);
    assign outputs[1421] = (layer4_outputs[750]) & (layer4_outputs[567]);
    assign outputs[1422] = layer4_outputs[1504];
    assign outputs[1423] = layer4_outputs[102];
    assign outputs[1424] = (layer4_outputs[1546]) & ~(layer4_outputs[1299]);
    assign outputs[1425] = layer4_outputs[2090];
    assign outputs[1426] = layer4_outputs[269];
    assign outputs[1427] = ~(layer4_outputs[1601]);
    assign outputs[1428] = layer4_outputs[1038];
    assign outputs[1429] = ~(layer4_outputs[1043]);
    assign outputs[1430] = (layer4_outputs[938]) ^ (layer4_outputs[1222]);
    assign outputs[1431] = ~(layer4_outputs[12]);
    assign outputs[1432] = layer4_outputs[733];
    assign outputs[1433] = ~(layer4_outputs[1757]);
    assign outputs[1434] = layer4_outputs[402];
    assign outputs[1435] = (layer4_outputs[48]) & ~(layer4_outputs[1557]);
    assign outputs[1436] = layer4_outputs[967];
    assign outputs[1437] = (layer4_outputs[1458]) ^ (layer4_outputs[813]);
    assign outputs[1438] = (layer4_outputs[608]) & ~(layer4_outputs[2017]);
    assign outputs[1439] = ~((layer4_outputs[251]) | (layer4_outputs[241]));
    assign outputs[1440] = ~((layer4_outputs[1871]) | (layer4_outputs[1967]));
    assign outputs[1441] = ~(layer4_outputs[2505]);
    assign outputs[1442] = ~(layer4_outputs[357]);
    assign outputs[1443] = layer4_outputs[799];
    assign outputs[1444] = ~((layer4_outputs[417]) ^ (layer4_outputs[2433]));
    assign outputs[1445] = ~((layer4_outputs[2067]) ^ (layer4_outputs[833]));
    assign outputs[1446] = (layer4_outputs[1354]) & ~(layer4_outputs[137]);
    assign outputs[1447] = ~(layer4_outputs[1329]);
    assign outputs[1448] = ~((layer4_outputs[116]) ^ (layer4_outputs[1809]));
    assign outputs[1449] = ~(layer4_outputs[352]);
    assign outputs[1450] = (layer4_outputs[870]) & (layer4_outputs[680]);
    assign outputs[1451] = ~(layer4_outputs[1050]) | (layer4_outputs[272]);
    assign outputs[1452] = (layer4_outputs[53]) & ~(layer4_outputs[1901]);
    assign outputs[1453] = ~((layer4_outputs[2133]) ^ (layer4_outputs[2391]));
    assign outputs[1454] = ~(layer4_outputs[1182]);
    assign outputs[1455] = (layer4_outputs[1741]) & ~(layer4_outputs[186]);
    assign outputs[1456] = ~(layer4_outputs[465]) | (layer4_outputs[1518]);
    assign outputs[1457] = (layer4_outputs[2187]) & ~(layer4_outputs[660]);
    assign outputs[1458] = (layer4_outputs[970]) ^ (layer4_outputs[1097]);
    assign outputs[1459] = ~(layer4_outputs[1836]);
    assign outputs[1460] = (layer4_outputs[1454]) ^ (layer4_outputs[2558]);
    assign outputs[1461] = (layer4_outputs[717]) | (layer4_outputs[1615]);
    assign outputs[1462] = ~(layer4_outputs[2353]);
    assign outputs[1463] = (layer4_outputs[668]) ^ (layer4_outputs[239]);
    assign outputs[1464] = ~((layer4_outputs[2053]) ^ (layer4_outputs[1466]));
    assign outputs[1465] = ~(layer4_outputs[75]);
    assign outputs[1466] = ~(layer4_outputs[2118]) | (layer4_outputs[951]);
    assign outputs[1467] = ~((layer4_outputs[590]) ^ (layer4_outputs[2291]));
    assign outputs[1468] = layer4_outputs[2494];
    assign outputs[1469] = layer4_outputs[2031];
    assign outputs[1470] = ~((layer4_outputs[2188]) & (layer4_outputs[358]));
    assign outputs[1471] = ~(layer4_outputs[1955]);
    assign outputs[1472] = (layer4_outputs[2119]) ^ (layer4_outputs[1251]);
    assign outputs[1473] = (layer4_outputs[1778]) & ~(layer4_outputs[1916]);
    assign outputs[1474] = layer4_outputs[764];
    assign outputs[1475] = ~(layer4_outputs[1219]);
    assign outputs[1476] = ~((layer4_outputs[1954]) ^ (layer4_outputs[177]));
    assign outputs[1477] = layer4_outputs[1904];
    assign outputs[1478] = ~((layer4_outputs[173]) ^ (layer4_outputs[435]));
    assign outputs[1479] = ~((layer4_outputs[104]) ^ (layer4_outputs[1921]));
    assign outputs[1480] = ~(layer4_outputs[1742]);
    assign outputs[1481] = ~(layer4_outputs[866]);
    assign outputs[1482] = layer4_outputs[1449];
    assign outputs[1483] = ~(layer4_outputs[1639]);
    assign outputs[1484] = ~(layer4_outputs[2431]);
    assign outputs[1485] = ~(layer4_outputs[1144]);
    assign outputs[1486] = ~(layer4_outputs[2378]);
    assign outputs[1487] = ~(layer4_outputs[1284]);
    assign outputs[1488] = layer4_outputs[483];
    assign outputs[1489] = ~(layer4_outputs[1164]) | (layer4_outputs[958]);
    assign outputs[1490] = (layer4_outputs[1023]) ^ (layer4_outputs[1528]);
    assign outputs[1491] = ~(layer4_outputs[2328]);
    assign outputs[1492] = layer4_outputs[1291];
    assign outputs[1493] = (layer4_outputs[842]) ^ (layer4_outputs[189]);
    assign outputs[1494] = (layer4_outputs[1592]) ^ (layer4_outputs[1795]);
    assign outputs[1495] = layer4_outputs[461];
    assign outputs[1496] = ~(layer4_outputs[636]);
    assign outputs[1497] = layer4_outputs[2080];
    assign outputs[1498] = ~((layer4_outputs[2134]) | (layer4_outputs[2393]));
    assign outputs[1499] = layer4_outputs[681];
    assign outputs[1500] = ~(layer4_outputs[183]);
    assign outputs[1501] = ~(layer4_outputs[1684]);
    assign outputs[1502] = layer4_outputs[957];
    assign outputs[1503] = ~(layer4_outputs[407]);
    assign outputs[1504] = layer4_outputs[522];
    assign outputs[1505] = layer4_outputs[881];
    assign outputs[1506] = (layer4_outputs[2178]) & (layer4_outputs[2155]);
    assign outputs[1507] = (layer4_outputs[1297]) & ~(layer4_outputs[77]);
    assign outputs[1508] = layer4_outputs[1640];
    assign outputs[1509] = ~(layer4_outputs[1290]);
    assign outputs[1510] = (layer4_outputs[323]) & ~(layer4_outputs[890]);
    assign outputs[1511] = (layer4_outputs[1349]) & ~(layer4_outputs[1387]);
    assign outputs[1512] = layer4_outputs[1314];
    assign outputs[1513] = ~(layer4_outputs[176]);
    assign outputs[1514] = ~((layer4_outputs[1224]) ^ (layer4_outputs[1232]));
    assign outputs[1515] = ~(layer4_outputs[1625]) | (layer4_outputs[926]);
    assign outputs[1516] = (layer4_outputs[2054]) & ~(layer4_outputs[1839]);
    assign outputs[1517] = ~((layer4_outputs[244]) ^ (layer4_outputs[1830]));
    assign outputs[1518] = (layer4_outputs[2416]) & (layer4_outputs[606]);
    assign outputs[1519] = ~(layer4_outputs[2317]);
    assign outputs[1520] = layer4_outputs[2213];
    assign outputs[1521] = ~((layer4_outputs[602]) | (layer4_outputs[1667]));
    assign outputs[1522] = layer4_outputs[2272];
    assign outputs[1523] = ~(layer4_outputs[1124]);
    assign outputs[1524] = layer4_outputs[925];
    assign outputs[1525] = (layer4_outputs[244]) & ~(layer4_outputs[1184]);
    assign outputs[1526] = ~(layer4_outputs[1415]);
    assign outputs[1527] = ~(layer4_outputs[2204]);
    assign outputs[1528] = ~(layer4_outputs[1146]);
    assign outputs[1529] = ~((layer4_outputs[2374]) & (layer4_outputs[700]));
    assign outputs[1530] = (layer4_outputs[1856]) ^ (layer4_outputs[2199]);
    assign outputs[1531] = layer4_outputs[1059];
    assign outputs[1532] = layer4_outputs[2073];
    assign outputs[1533] = ~((layer4_outputs[1108]) & (layer4_outputs[1890]));
    assign outputs[1534] = layer4_outputs[1726];
    assign outputs[1535] = (layer4_outputs[1203]) | (layer4_outputs[948]);
    assign outputs[1536] = ~(layer4_outputs[2441]);
    assign outputs[1537] = (layer4_outputs[995]) & ~(layer4_outputs[1125]);
    assign outputs[1538] = layer4_outputs[1264];
    assign outputs[1539] = ~((layer4_outputs[284]) ^ (layer4_outputs[1835]));
    assign outputs[1540] = layer4_outputs[305];
    assign outputs[1541] = layer4_outputs[2306];
    assign outputs[1542] = layer4_outputs[1775];
    assign outputs[1543] = layer4_outputs[172];
    assign outputs[1544] = ~(layer4_outputs[33]);
    assign outputs[1545] = ~(layer4_outputs[2150]) | (layer4_outputs[1240]);
    assign outputs[1546] = (layer4_outputs[309]) & ~(layer4_outputs[920]);
    assign outputs[1547] = ~(layer4_outputs[287]);
    assign outputs[1548] = (layer4_outputs[1822]) | (layer4_outputs[2099]);
    assign outputs[1549] = layer4_outputs[1619];
    assign outputs[1550] = ~(layer4_outputs[1426]);
    assign outputs[1551] = (layer4_outputs[2079]) & (layer4_outputs[2194]);
    assign outputs[1552] = (layer4_outputs[308]) & ~(layer4_outputs[1403]);
    assign outputs[1553] = (layer4_outputs[1584]) | (layer4_outputs[612]);
    assign outputs[1554] = ~((layer4_outputs[2282]) ^ (layer4_outputs[2493]));
    assign outputs[1555] = ~(layer4_outputs[2077]);
    assign outputs[1556] = ~(layer4_outputs[653]);
    assign outputs[1557] = ~(layer4_outputs[2333]);
    assign outputs[1558] = layer4_outputs[46];
    assign outputs[1559] = ~(layer4_outputs[849]);
    assign outputs[1560] = (layer4_outputs[1476]) & ~(layer4_outputs[1438]);
    assign outputs[1561] = (layer4_outputs[995]) & (layer4_outputs[281]);
    assign outputs[1562] = ~(layer4_outputs[2439]);
    assign outputs[1563] = ~(layer4_outputs[427]);
    assign outputs[1564] = ~(layer4_outputs[669]);
    assign outputs[1565] = layer4_outputs[992];
    assign outputs[1566] = ~(layer4_outputs[2098]);
    assign outputs[1567] = layer4_outputs[1356];
    assign outputs[1568] = layer4_outputs[328];
    assign outputs[1569] = ~((layer4_outputs[106]) & (layer4_outputs[2505]));
    assign outputs[1570] = layer4_outputs[481];
    assign outputs[1571] = ~(layer4_outputs[2315]) | (layer4_outputs[2312]);
    assign outputs[1572] = (layer4_outputs[2516]) & (layer4_outputs[2548]);
    assign outputs[1573] = layer4_outputs[430];
    assign outputs[1574] = layer4_outputs[2414];
    assign outputs[1575] = ~((layer4_outputs[2164]) ^ (layer4_outputs[1331]));
    assign outputs[1576] = ~(layer4_outputs[292]);
    assign outputs[1577] = ~((layer4_outputs[349]) | (layer4_outputs[2207]));
    assign outputs[1578] = layer4_outputs[172];
    assign outputs[1579] = layer4_outputs[1424];
    assign outputs[1580] = ~(layer4_outputs[1990]);
    assign outputs[1581] = layer4_outputs[845];
    assign outputs[1582] = (layer4_outputs[2011]) & ~(layer4_outputs[645]);
    assign outputs[1583] = (layer4_outputs[111]) & (layer4_outputs[1275]);
    assign outputs[1584] = ~((layer4_outputs[1651]) | (layer4_outputs[889]));
    assign outputs[1585] = ~((layer4_outputs[1500]) ^ (layer4_outputs[906]));
    assign outputs[1586] = (layer4_outputs[1583]) & ~(layer4_outputs[710]);
    assign outputs[1587] = ~(layer4_outputs[168]) | (layer4_outputs[1272]);
    assign outputs[1588] = (layer4_outputs[791]) | (layer4_outputs[895]);
    assign outputs[1589] = ~((layer4_outputs[2212]) ^ (layer4_outputs[2276]));
    assign outputs[1590] = ~(layer4_outputs[1872]) | (layer4_outputs[251]);
    assign outputs[1591] = ~(layer4_outputs[1922]);
    assign outputs[1592] = layer4_outputs[739];
    assign outputs[1593] = ~(layer4_outputs[2197]);
    assign outputs[1594] = layer4_outputs[335];
    assign outputs[1595] = ~(layer4_outputs[2197]);
    assign outputs[1596] = ~((layer4_outputs[2047]) | (layer4_outputs[1855]));
    assign outputs[1597] = ~(layer4_outputs[1805]);
    assign outputs[1598] = layer4_outputs[2180];
    assign outputs[1599] = (layer4_outputs[2414]) & (layer4_outputs[2073]);
    assign outputs[1600] = (layer4_outputs[1919]) ^ (layer4_outputs[1181]);
    assign outputs[1601] = layer4_outputs[1850];
    assign outputs[1602] = ~(layer4_outputs[1678]);
    assign outputs[1603] = (layer4_outputs[1031]) | (layer4_outputs[2224]);
    assign outputs[1604] = ~((layer4_outputs[1172]) ^ (layer4_outputs[954]));
    assign outputs[1605] = ~((layer4_outputs[2072]) ^ (layer4_outputs[267]));
    assign outputs[1606] = ~(layer4_outputs[2161]);
    assign outputs[1607] = layer4_outputs[2473];
    assign outputs[1608] = ~(layer4_outputs[1821]) | (layer4_outputs[2147]);
    assign outputs[1609] = ~(layer4_outputs[278]);
    assign outputs[1610] = layer4_outputs[2394];
    assign outputs[1611] = layer4_outputs[1506];
    assign outputs[1612] = ~((layer4_outputs[2476]) | (layer4_outputs[93]));
    assign outputs[1613] = (layer4_outputs[1385]) | (layer4_outputs[166]);
    assign outputs[1614] = layer4_outputs[336];
    assign outputs[1615] = ~(layer4_outputs[459]);
    assign outputs[1616] = ~((layer4_outputs[2547]) & (layer4_outputs[1632]));
    assign outputs[1617] = ~(layer4_outputs[1252]);
    assign outputs[1618] = ~(layer4_outputs[2116]);
    assign outputs[1619] = layer4_outputs[2210];
    assign outputs[1620] = ~(layer4_outputs[2236]) | (layer4_outputs[1188]);
    assign outputs[1621] = layer4_outputs[2111];
    assign outputs[1622] = layer4_outputs[877];
    assign outputs[1623] = layer4_outputs[1072];
    assign outputs[1624] = layer4_outputs[1151];
    assign outputs[1625] = layer4_outputs[2394];
    assign outputs[1626] = ~(layer4_outputs[1369]);
    assign outputs[1627] = ~(layer4_outputs[1527]) | (layer4_outputs[1719]);
    assign outputs[1628] = layer4_outputs[1234];
    assign outputs[1629] = ~(layer4_outputs[1367]);
    assign outputs[1630] = (layer4_outputs[2510]) ^ (layer4_outputs[1064]);
    assign outputs[1631] = ~(layer4_outputs[307]);
    assign outputs[1632] = layer4_outputs[2265];
    assign outputs[1633] = ~(layer4_outputs[354]);
    assign outputs[1634] = (layer4_outputs[1582]) ^ (layer4_outputs[498]);
    assign outputs[1635] = ~(layer4_outputs[85]);
    assign outputs[1636] = ~((layer4_outputs[671]) ^ (layer4_outputs[2169]));
    assign outputs[1637] = ~(layer4_outputs[881]);
    assign outputs[1638] = ~(layer4_outputs[728]);
    assign outputs[1639] = ~(layer4_outputs[784]);
    assign outputs[1640] = layer4_outputs[1241];
    assign outputs[1641] = ~((layer4_outputs[2026]) | (layer4_outputs[1768]));
    assign outputs[1642] = layer4_outputs[2312];
    assign outputs[1643] = ~((layer4_outputs[735]) | (layer4_outputs[2190]));
    assign outputs[1644] = layer4_outputs[1696];
    assign outputs[1645] = ~(layer4_outputs[2428]);
    assign outputs[1646] = ~(layer4_outputs[161]);
    assign outputs[1647] = ~(layer4_outputs[1741]);
    assign outputs[1648] = layer4_outputs[809];
    assign outputs[1649] = ~(layer4_outputs[1695]);
    assign outputs[1650] = ~(layer4_outputs[378]);
    assign outputs[1651] = ~((layer4_outputs[1764]) ^ (layer4_outputs[506]));
    assign outputs[1652] = (layer4_outputs[1619]) & (layer4_outputs[385]);
    assign outputs[1653] = layer4_outputs[1285];
    assign outputs[1654] = (layer4_outputs[128]) & ~(layer4_outputs[914]);
    assign outputs[1655] = layer4_outputs[1645];
    assign outputs[1656] = (layer4_outputs[460]) & ~(layer4_outputs[1087]);
    assign outputs[1657] = layer4_outputs[1266];
    assign outputs[1658] = layer4_outputs[767];
    assign outputs[1659] = (layer4_outputs[2517]) ^ (layer4_outputs[534]);
    assign outputs[1660] = (layer4_outputs[553]) & (layer4_outputs[1278]);
    assign outputs[1661] = layer4_outputs[1496];
    assign outputs[1662] = ~(layer4_outputs[1150]);
    assign outputs[1663] = ~(layer4_outputs[41]);
    assign outputs[1664] = ~(layer4_outputs[1534]);
    assign outputs[1665] = layer4_outputs[695];
    assign outputs[1666] = (layer4_outputs[191]) ^ (layer4_outputs[1993]);
    assign outputs[1667] = ~(layer4_outputs[1490]);
    assign outputs[1668] = ~((layer4_outputs[1094]) | (layer4_outputs[1484]));
    assign outputs[1669] = layer4_outputs[830];
    assign outputs[1670] = ~(layer4_outputs[704]);
    assign outputs[1671] = (layer4_outputs[1051]) & (layer4_outputs[1971]);
    assign outputs[1672] = layer4_outputs[908];
    assign outputs[1673] = (layer4_outputs[2188]) & ~(layer4_outputs[2055]);
    assign outputs[1674] = ~(layer4_outputs[782]);
    assign outputs[1675] = layer4_outputs[1496];
    assign outputs[1676] = ~(layer4_outputs[1448]);
    assign outputs[1677] = layer4_outputs[495];
    assign outputs[1678] = (layer4_outputs[427]) ^ (layer4_outputs[486]);
    assign outputs[1679] = layer4_outputs[1966];
    assign outputs[1680] = (layer4_outputs[1579]) & ~(layer4_outputs[1691]);
    assign outputs[1681] = ~(layer4_outputs[2295]) | (layer4_outputs[1267]);
    assign outputs[1682] = (layer4_outputs[1276]) & (layer4_outputs[902]);
    assign outputs[1683] = layer4_outputs[384];
    assign outputs[1684] = (layer4_outputs[848]) ^ (layer4_outputs[2006]);
    assign outputs[1685] = ~(layer4_outputs[974]);
    assign outputs[1686] = layer4_outputs[1674];
    assign outputs[1687] = layer4_outputs[1820];
    assign outputs[1688] = ~(layer4_outputs[2015]);
    assign outputs[1689] = ~(layer4_outputs[883]);
    assign outputs[1690] = ~(layer4_outputs[709]);
    assign outputs[1691] = ~(layer4_outputs[817]);
    assign outputs[1692] = (layer4_outputs[1146]) & (layer4_outputs[2300]);
    assign outputs[1693] = (layer4_outputs[2436]) & ~(layer4_outputs[1616]);
    assign outputs[1694] = layer4_outputs[547];
    assign outputs[1695] = (layer4_outputs[383]) ^ (layer4_outputs[484]);
    assign outputs[1696] = ~(layer4_outputs[2048]);
    assign outputs[1697] = ~(layer4_outputs[1250]);
    assign outputs[1698] = ~(layer4_outputs[275]);
    assign outputs[1699] = layer4_outputs[1285];
    assign outputs[1700] = ~((layer4_outputs[2540]) & (layer4_outputs[646]));
    assign outputs[1701] = ~(layer4_outputs[409]);
    assign outputs[1702] = (layer4_outputs[839]) & (layer4_outputs[54]);
    assign outputs[1703] = ~(layer4_outputs[854]);
    assign outputs[1704] = (layer4_outputs[1895]) & (layer4_outputs[2259]);
    assign outputs[1705] = (layer4_outputs[553]) ^ (layer4_outputs[1835]);
    assign outputs[1706] = ~((layer4_outputs[2042]) | (layer4_outputs[159]));
    assign outputs[1707] = layer4_outputs[864];
    assign outputs[1708] = (layer4_outputs[1071]) ^ (layer4_outputs[1139]);
    assign outputs[1709] = layer4_outputs[1875];
    assign outputs[1710] = layer4_outputs[732];
    assign outputs[1711] = layer4_outputs[1867];
    assign outputs[1712] = layer4_outputs[2429];
    assign outputs[1713] = layer4_outputs[830];
    assign outputs[1714] = ~(layer4_outputs[1168]);
    assign outputs[1715] = layer4_outputs[899];
    assign outputs[1716] = ~((layer4_outputs[1428]) ^ (layer4_outputs[811]));
    assign outputs[1717] = layer4_outputs[1840];
    assign outputs[1718] = (layer4_outputs[664]) & (layer4_outputs[1696]);
    assign outputs[1719] = ~(layer4_outputs[669]);
    assign outputs[1720] = ~(layer4_outputs[2321]);
    assign outputs[1721] = ~(layer4_outputs[443]);
    assign outputs[1722] = (layer4_outputs[2151]) & ~(layer4_outputs[2095]);
    assign outputs[1723] = ~(layer4_outputs[2016]);
    assign outputs[1724] = ~(layer4_outputs[1392]);
    assign outputs[1725] = ~(layer4_outputs[500]);
    assign outputs[1726] = ~(layer4_outputs[52]);
    assign outputs[1727] = (layer4_outputs[1885]) & ~(layer4_outputs[1844]);
    assign outputs[1728] = layer4_outputs[778];
    assign outputs[1729] = layer4_outputs[2100];
    assign outputs[1730] = layer4_outputs[2151];
    assign outputs[1731] = layer4_outputs[1079];
    assign outputs[1732] = ~(layer4_outputs[1014]);
    assign outputs[1733] = ~(layer4_outputs[1265]);
    assign outputs[1734] = ~(layer4_outputs[587]);
    assign outputs[1735] = layer4_outputs[971];
    assign outputs[1736] = ~(layer4_outputs[2418]) | (layer4_outputs[2432]);
    assign outputs[1737] = layer4_outputs[173];
    assign outputs[1738] = ~((layer4_outputs[29]) ^ (layer4_outputs[168]));
    assign outputs[1739] = ~(layer4_outputs[2373]);
    assign outputs[1740] = ~(layer4_outputs[1620]);
    assign outputs[1741] = ~((layer4_outputs[2446]) ^ (layer4_outputs[1997]));
    assign outputs[1742] = ~(layer4_outputs[78]);
    assign outputs[1743] = ~((layer4_outputs[494]) | (layer4_outputs[1483]));
    assign outputs[1744] = (layer4_outputs[878]) ^ (layer4_outputs[2454]);
    assign outputs[1745] = (layer4_outputs[2537]) ^ (layer4_outputs[745]);
    assign outputs[1746] = ~(layer4_outputs[0]);
    assign outputs[1747] = ~((layer4_outputs[935]) & (layer4_outputs[1452]));
    assign outputs[1748] = layer4_outputs[2025];
    assign outputs[1749] = ~(layer4_outputs[1160]);
    assign outputs[1750] = ~(layer4_outputs[517]);
    assign outputs[1751] = ~(layer4_outputs[93]) | (layer4_outputs[1549]);
    assign outputs[1752] = ~(layer4_outputs[1828]);
    assign outputs[1753] = ~(layer4_outputs[2385]);
    assign outputs[1754] = ~((layer4_outputs[1540]) & (layer4_outputs[633]));
    assign outputs[1755] = ~(layer4_outputs[2423]);
    assign outputs[1756] = ~(layer4_outputs[1348]);
    assign outputs[1757] = ~(layer4_outputs[1263]);
    assign outputs[1758] = ~(layer4_outputs[2482]);
    assign outputs[1759] = layer4_outputs[1342];
    assign outputs[1760] = layer4_outputs[513];
    assign outputs[1761] = ~(layer4_outputs[129]);
    assign outputs[1762] = ~(layer4_outputs[2208]);
    assign outputs[1763] = layer4_outputs[493];
    assign outputs[1764] = layer4_outputs[1048];
    assign outputs[1765] = layer4_outputs[4];
    assign outputs[1766] = layer4_outputs[1423];
    assign outputs[1767] = (layer4_outputs[1408]) ^ (layer4_outputs[1119]);
    assign outputs[1768] = ~(layer4_outputs[2371]);
    assign outputs[1769] = layer4_outputs[234];
    assign outputs[1770] = ~(layer4_outputs[759]);
    assign outputs[1771] = ~((layer4_outputs[745]) ^ (layer4_outputs[1087]));
    assign outputs[1772] = (layer4_outputs[564]) ^ (layer4_outputs[1456]);
    assign outputs[1773] = ~((layer4_outputs[1048]) ^ (layer4_outputs[1095]));
    assign outputs[1774] = ~(layer4_outputs[538]);
    assign outputs[1775] = ~(layer4_outputs[1514]);
    assign outputs[1776] = layer4_outputs[1259];
    assign outputs[1777] = (layer4_outputs[446]) ^ (layer4_outputs[831]);
    assign outputs[1778] = layer4_outputs[1504];
    assign outputs[1779] = ~(layer4_outputs[707]);
    assign outputs[1780] = ~(layer4_outputs[933]);
    assign outputs[1781] = (layer4_outputs[2282]) | (layer4_outputs[478]);
    assign outputs[1782] = layer4_outputs[2255];
    assign outputs[1783] = (layer4_outputs[1422]) | (layer4_outputs[1356]);
    assign outputs[1784] = layer4_outputs[126];
    assign outputs[1785] = layer4_outputs[2226];
    assign outputs[1786] = ~(layer4_outputs[442]);
    assign outputs[1787] = (layer4_outputs[42]) & (layer4_outputs[2034]);
    assign outputs[1788] = ~(layer4_outputs[827]);
    assign outputs[1789] = ~((layer4_outputs[1367]) ^ (layer4_outputs[2110]));
    assign outputs[1790] = ~(layer4_outputs[1691]);
    assign outputs[1791] = ~(layer4_outputs[1658]);
    assign outputs[1792] = ~(layer4_outputs[1561]) | (layer4_outputs[661]);
    assign outputs[1793] = layer4_outputs[2202];
    assign outputs[1794] = ~((layer4_outputs[1397]) | (layer4_outputs[676]));
    assign outputs[1795] = ~(layer4_outputs[1415]);
    assign outputs[1796] = ~((layer4_outputs[1916]) | (layer4_outputs[1140]));
    assign outputs[1797] = ~(layer4_outputs[1501]);
    assign outputs[1798] = ~((layer4_outputs[1173]) | (layer4_outputs[1221]));
    assign outputs[1799] = ~(layer4_outputs[802]);
    assign outputs[1800] = ~(layer4_outputs[1347]);
    assign outputs[1801] = ~(layer4_outputs[979]);
    assign outputs[1802] = ~((layer4_outputs[55]) | (layer4_outputs[2252]));
    assign outputs[1803] = ~(layer4_outputs[281]);
    assign outputs[1804] = (layer4_outputs[1827]) & (layer4_outputs[1089]);
    assign outputs[1805] = layer4_outputs[893];
    assign outputs[1806] = ~(layer4_outputs[1112]);
    assign outputs[1807] = layer4_outputs[527];
    assign outputs[1808] = ~((layer4_outputs[1598]) ^ (layer4_outputs[1149]));
    assign outputs[1809] = ~(layer4_outputs[1826]);
    assign outputs[1810] = ~(layer4_outputs[230]);
    assign outputs[1811] = ~(layer4_outputs[2504]);
    assign outputs[1812] = ~((layer4_outputs[625]) | (layer4_outputs[60]));
    assign outputs[1813] = ~(layer4_outputs[1551]);
    assign outputs[1814] = ~(layer4_outputs[837]);
    assign outputs[1815] = ~(layer4_outputs[2442]);
    assign outputs[1816] = layer4_outputs[2314];
    assign outputs[1817] = ~((layer4_outputs[936]) ^ (layer4_outputs[387]));
    assign outputs[1818] = layer4_outputs[2149];
    assign outputs[1819] = layer4_outputs[964];
    assign outputs[1820] = layer4_outputs[912];
    assign outputs[1821] = (layer4_outputs[2279]) & ~(layer4_outputs[2496]);
    assign outputs[1822] = (layer4_outputs[1303]) & (layer4_outputs[2014]);
    assign outputs[1823] = ~((layer4_outputs[170]) | (layer4_outputs[1028]));
    assign outputs[1824] = layer4_outputs[1871];
    assign outputs[1825] = layer4_outputs[1386];
    assign outputs[1826] = ~((layer4_outputs[2010]) | (layer4_outputs[1198]));
    assign outputs[1827] = layer4_outputs[1673];
    assign outputs[1828] = ~(layer4_outputs[466]) | (layer4_outputs[2319]);
    assign outputs[1829] = ~(layer4_outputs[405]);
    assign outputs[1830] = layer4_outputs[589];
    assign outputs[1831] = layer4_outputs[2069];
    assign outputs[1832] = layer4_outputs[1747];
    assign outputs[1833] = (layer4_outputs[976]) & ~(layer4_outputs[1196]);
    assign outputs[1834] = (layer4_outputs[1996]) & ~(layer4_outputs[628]);
    assign outputs[1835] = (layer4_outputs[485]) & (layer4_outputs[1122]);
    assign outputs[1836] = ~(layer4_outputs[1590]);
    assign outputs[1837] = (layer4_outputs[1805]) & ~(layer4_outputs[607]);
    assign outputs[1838] = ~(layer4_outputs[298]);
    assign outputs[1839] = ~(layer4_outputs[880]);
    assign outputs[1840] = (layer4_outputs[780]) & ~(layer4_outputs[894]);
    assign outputs[1841] = (layer4_outputs[2261]) & ~(layer4_outputs[1230]);
    assign outputs[1842] = layer4_outputs[679];
    assign outputs[1843] = ~(layer4_outputs[2080]);
    assign outputs[1844] = ~(layer4_outputs[1571]);
    assign outputs[1845] = (layer4_outputs[1766]) & ~(layer4_outputs[2384]);
    assign outputs[1846] = ~((layer4_outputs[305]) | (layer4_outputs[2180]));
    assign outputs[1847] = ~((layer4_outputs[913]) & (layer4_outputs[1086]));
    assign outputs[1848] = (layer4_outputs[369]) ^ (layer4_outputs[1069]);
    assign outputs[1849] = (layer4_outputs[1597]) & ~(layer4_outputs[905]);
    assign outputs[1850] = layer4_outputs[2529];
    assign outputs[1851] = (layer4_outputs[1225]) & ~(layer4_outputs[1744]);
    assign outputs[1852] = ~(layer4_outputs[1183]);
    assign outputs[1853] = layer4_outputs[774];
    assign outputs[1854] = ~(layer4_outputs[1796]);
    assign outputs[1855] = layer4_outputs[386];
    assign outputs[1856] = ~((layer4_outputs[402]) | (layer4_outputs[242]));
    assign outputs[1857] = ~(layer4_outputs[1311]);
    assign outputs[1858] = (layer4_outputs[130]) & (layer4_outputs[2315]);
    assign outputs[1859] = (layer4_outputs[77]) & ~(layer4_outputs[1243]);
    assign outputs[1860] = (layer4_outputs[1405]) ^ (layer4_outputs[1565]);
    assign outputs[1861] = ~(layer4_outputs[1350]);
    assign outputs[1862] = ~((layer4_outputs[2021]) ^ (layer4_outputs[2467]));
    assign outputs[1863] = layer4_outputs[1260];
    assign outputs[1864] = (layer4_outputs[2419]) & (layer4_outputs[716]);
    assign outputs[1865] = ~((layer4_outputs[1103]) | (layer4_outputs[819]));
    assign outputs[1866] = (layer4_outputs[1586]) & ~(layer4_outputs[10]);
    assign outputs[1867] = (layer4_outputs[1853]) & ~(layer4_outputs[2354]);
    assign outputs[1868] = ~(layer4_outputs[1445]);
    assign outputs[1869] = ~((layer4_outputs[226]) | (layer4_outputs[1308]));
    assign outputs[1870] = ~(layer4_outputs[543]);
    assign outputs[1871] = (layer4_outputs[82]) & (layer4_outputs[1235]);
    assign outputs[1872] = ~(layer4_outputs[1615]);
    assign outputs[1873] = ~((layer4_outputs[1027]) | (layer4_outputs[260]));
    assign outputs[1874] = layer4_outputs[1651];
    assign outputs[1875] = (layer4_outputs[266]) & ~(layer4_outputs[615]);
    assign outputs[1876] = ~(layer4_outputs[299]);
    assign outputs[1877] = ~(layer4_outputs[1227]);
    assign outputs[1878] = layer4_outputs[2545];
    assign outputs[1879] = (layer4_outputs[1959]) & ~(layer4_outputs[277]);
    assign outputs[1880] = ~((layer4_outputs[23]) | (layer4_outputs[2141]));
    assign outputs[1881] = (layer4_outputs[1178]) & (layer4_outputs[1441]);
    assign outputs[1882] = layer4_outputs[2361];
    assign outputs[1883] = (layer4_outputs[2284]) & ~(layer4_outputs[1638]);
    assign outputs[1884] = ~(layer4_outputs[2135]);
    assign outputs[1885] = layer4_outputs[937];
    assign outputs[1886] = (layer4_outputs[1130]) & (layer4_outputs[2304]);
    assign outputs[1887] = layer4_outputs[70];
    assign outputs[1888] = (layer4_outputs[1905]) ^ (layer4_outputs[831]);
    assign outputs[1889] = ~(layer4_outputs[1945]);
    assign outputs[1890] = ~(layer4_outputs[322]);
    assign outputs[1891] = (layer4_outputs[2190]) & ~(layer4_outputs[1016]);
    assign outputs[1892] = ~((layer4_outputs[1086]) ^ (layer4_outputs[1961]));
    assign outputs[1893] = ~(layer4_outputs[2203]);
    assign outputs[1894] = ~(layer4_outputs[382]);
    assign outputs[1895] = layer4_outputs[559];
    assign outputs[1896] = layer4_outputs[1758];
    assign outputs[1897] = ~(layer4_outputs[1807]);
    assign outputs[1898] = layer4_outputs[1790];
    assign outputs[1899] = layer4_outputs[1937];
    assign outputs[1900] = (layer4_outputs[180]) & ~(layer4_outputs[786]);
    assign outputs[1901] = ~((layer4_outputs[1808]) ^ (layer4_outputs[462]));
    assign outputs[1902] = layer4_outputs[320];
    assign outputs[1903] = ~((layer4_outputs[1934]) | (layer4_outputs[331]));
    assign outputs[1904] = (layer4_outputs[1958]) ^ (layer4_outputs[1298]);
    assign outputs[1905] = ~(layer4_outputs[641]);
    assign outputs[1906] = layer4_outputs[161];
    assign outputs[1907] = layer4_outputs[2202];
    assign outputs[1908] = ~((layer4_outputs[1636]) ^ (layer4_outputs[1833]));
    assign outputs[1909] = ~(layer4_outputs[1624]);
    assign outputs[1910] = layer4_outputs[727];
    assign outputs[1911] = ~(layer4_outputs[723]);
    assign outputs[1912] = (layer4_outputs[374]) & (layer4_outputs[1984]);
    assign outputs[1913] = layer4_outputs[763];
    assign outputs[1914] = ~((layer4_outputs[1714]) | (layer4_outputs[1155]));
    assign outputs[1915] = (layer4_outputs[407]) & ~(layer4_outputs[825]);
    assign outputs[1916] = ~((layer4_outputs[2132]) ^ (layer4_outputs[2217]));
    assign outputs[1917] = layer4_outputs[327];
    assign outputs[1918] = ~(layer4_outputs[1948]);
    assign outputs[1919] = ~(layer4_outputs[1201]);
    assign outputs[1920] = layer4_outputs[1106];
    assign outputs[1921] = (layer4_outputs[2170]) & (layer4_outputs[1570]);
    assign outputs[1922] = ~(layer4_outputs[456]);
    assign outputs[1923] = ~((layer4_outputs[970]) | (layer4_outputs[1724]));
    assign outputs[1924] = (layer4_outputs[978]) ^ (layer4_outputs[2063]);
    assign outputs[1925] = ~(layer4_outputs[1233]);
    assign outputs[1926] = (layer4_outputs[1017]) & ~(layer4_outputs[80]);
    assign outputs[1927] = (layer4_outputs[1022]) & ~(layer4_outputs[1793]);
    assign outputs[1928] = layer4_outputs[1572];
    assign outputs[1929] = ~((layer4_outputs[1763]) | (layer4_outputs[333]));
    assign outputs[1930] = layer4_outputs[1318];
    assign outputs[1931] = layer4_outputs[2422];
    assign outputs[1932] = ~(layer4_outputs[2500]);
    assign outputs[1933] = ~(layer4_outputs[501]);
    assign outputs[1934] = ~((layer4_outputs[911]) | (layer4_outputs[1165]));
    assign outputs[1935] = ~(layer4_outputs[1707]);
    assign outputs[1936] = (layer4_outputs[1115]) ^ (layer4_outputs[1573]);
    assign outputs[1937] = layer4_outputs[1050];
    assign outputs[1938] = ~(layer4_outputs[2407]);
    assign outputs[1939] = ~(layer4_outputs[2387]);
    assign outputs[1940] = ~((layer4_outputs[121]) | (layer4_outputs[2487]));
    assign outputs[1941] = layer4_outputs[2136];
    assign outputs[1942] = (layer4_outputs[475]) & ~(layer4_outputs[1608]);
    assign outputs[1943] = ~(layer4_outputs[1012]);
    assign outputs[1944] = (layer4_outputs[2443]) & ~(layer4_outputs[2260]);
    assign outputs[1945] = (layer4_outputs[2347]) | (layer4_outputs[1021]);
    assign outputs[1946] = ~(layer4_outputs[2514]);
    assign outputs[1947] = layer4_outputs[2170];
    assign outputs[1948] = ~(layer4_outputs[207]);
    assign outputs[1949] = ~(layer4_outputs[1590]);
    assign outputs[1950] = ~(layer4_outputs[1125]);
    assign outputs[1951] = (layer4_outputs[1600]) & ~(layer4_outputs[1403]);
    assign outputs[1952] = (layer4_outputs[2421]) & (layer4_outputs[2338]);
    assign outputs[1953] = (layer4_outputs[798]) & (layer4_outputs[2280]);
    assign outputs[1954] = layer4_outputs[759];
    assign outputs[1955] = ~(layer4_outputs[67]);
    assign outputs[1956] = (layer4_outputs[2008]) & ~(layer4_outputs[975]);
    assign outputs[1957] = ~(layer4_outputs[1233]);
    assign outputs[1958] = layer4_outputs[76];
    assign outputs[1959] = ~(layer4_outputs[1929]);
    assign outputs[1960] = layer4_outputs[1819];
    assign outputs[1961] = (layer4_outputs[2511]) & (layer4_outputs[704]);
    assign outputs[1962] = layer4_outputs[354];
    assign outputs[1963] = (layer4_outputs[2424]) ^ (layer4_outputs[851]);
    assign outputs[1964] = ~(layer4_outputs[1323]);
    assign outputs[1965] = (layer4_outputs[303]) ^ (layer4_outputs[1887]);
    assign outputs[1966] = ~(layer4_outputs[1831]);
    assign outputs[1967] = layer4_outputs[1621];
    assign outputs[1968] = layer4_outputs[47];
    assign outputs[1969] = layer4_outputs[940];
    assign outputs[1970] = (layer4_outputs[1715]) & ~(layer4_outputs[2268]);
    assign outputs[1971] = layer4_outputs[252];
    assign outputs[1972] = ~(layer4_outputs[965]);
    assign outputs[1973] = ~(layer4_outputs[684]);
    assign outputs[1974] = ~(layer4_outputs[2183]);
    assign outputs[1975] = (layer4_outputs[1044]) & ~(layer4_outputs[100]);
    assign outputs[1976] = ~(layer4_outputs[1728]);
    assign outputs[1977] = layer4_outputs[498];
    assign outputs[1978] = ~(layer4_outputs[149]);
    assign outputs[1979] = layer4_outputs[1057];
    assign outputs[1980] = ~((layer4_outputs[534]) ^ (layer4_outputs[672]));
    assign outputs[1981] = layer4_outputs[2472];
    assign outputs[1982] = ~(layer4_outputs[1508]);
    assign outputs[1983] = ~(layer4_outputs[715]);
    assign outputs[1984] = ~(layer4_outputs[259]);
    assign outputs[1985] = ~((layer4_outputs[829]) ^ (layer4_outputs[1755]));
    assign outputs[1986] = ~((layer4_outputs[2364]) ^ (layer4_outputs[966]));
    assign outputs[1987] = ~(layer4_outputs[394]);
    assign outputs[1988] = (layer4_outputs[2198]) ^ (layer4_outputs[1943]);
    assign outputs[1989] = (layer4_outputs[1873]) ^ (layer4_outputs[1898]);
    assign outputs[1990] = layer4_outputs[63];
    assign outputs[1991] = layer4_outputs[1758];
    assign outputs[1992] = ~((layer4_outputs[1524]) ^ (layer4_outputs[884]));
    assign outputs[1993] = (layer4_outputs[2545]) & ~(layer4_outputs[733]);
    assign outputs[1994] = layer4_outputs[944];
    assign outputs[1995] = ~(layer4_outputs[1892]);
    assign outputs[1996] = (layer4_outputs[474]) & (layer4_outputs[578]);
    assign outputs[1997] = ~((layer4_outputs[808]) & (layer4_outputs[2389]));
    assign outputs[1998] = ~(layer4_outputs[539]);
    assign outputs[1999] = layer4_outputs[2291];
    assign outputs[2000] = layer4_outputs[1189];
    assign outputs[2001] = ~(layer4_outputs[2129]);
    assign outputs[2002] = ~(layer4_outputs[1971]);
    assign outputs[2003] = (layer4_outputs[1575]) & ~(layer4_outputs[1214]);
    assign outputs[2004] = layer4_outputs[903];
    assign outputs[2005] = ~(layer4_outputs[1487]);
    assign outputs[2006] = ~(layer4_outputs[100]);
    assign outputs[2007] = (layer4_outputs[1235]) & (layer4_outputs[632]);
    assign outputs[2008] = ~(layer4_outputs[3]);
    assign outputs[2009] = ~(layer4_outputs[2489]);
    assign outputs[2010] = ~(layer4_outputs[1493]);
    assign outputs[2011] = ~(layer4_outputs[2276]);
    assign outputs[2012] = layer4_outputs[1433];
    assign outputs[2013] = (layer4_outputs[340]) & ~(layer4_outputs[1862]);
    assign outputs[2014] = ~(layer4_outputs[2548]);
    assign outputs[2015] = layer4_outputs[130];
    assign outputs[2016] = (layer4_outputs[1036]) & (layer4_outputs[413]);
    assign outputs[2017] = (layer4_outputs[158]) & (layer4_outputs[2007]);
    assign outputs[2018] = layer4_outputs[1711];
    assign outputs[2019] = ~(layer4_outputs[1103]);
    assign outputs[2020] = layer4_outputs[1184];
    assign outputs[2021] = (layer4_outputs[2382]) ^ (layer4_outputs[286]);
    assign outputs[2022] = layer4_outputs[1398];
    assign outputs[2023] = (layer4_outputs[1370]) ^ (layer4_outputs[237]);
    assign outputs[2024] = ~(layer4_outputs[1243]);
    assign outputs[2025] = layer4_outputs[1];
    assign outputs[2026] = layer4_outputs[2538];
    assign outputs[2027] = layer4_outputs[1413];
    assign outputs[2028] = ~(layer4_outputs[897]);
    assign outputs[2029] = ~(layer4_outputs[363]) | (layer4_outputs[1244]);
    assign outputs[2030] = (layer4_outputs[566]) & ~(layer4_outputs[1315]);
    assign outputs[2031] = (layer4_outputs[458]) & (layer4_outputs[401]);
    assign outputs[2032] = ~(layer4_outputs[668]);
    assign outputs[2033] = (layer4_outputs[1460]) & ~(layer4_outputs[1520]);
    assign outputs[2034] = (layer4_outputs[197]) & ~(layer4_outputs[2203]);
    assign outputs[2035] = layer4_outputs[1841];
    assign outputs[2036] = ~(layer4_outputs[1964]);
    assign outputs[2037] = (layer4_outputs[1482]) & (layer4_outputs[2075]);
    assign outputs[2038] = (layer4_outputs[1444]) & ~(layer4_outputs[870]);
    assign outputs[2039] = ~(layer4_outputs[1447]);
    assign outputs[2040] = ~(layer4_outputs[1394]);
    assign outputs[2041] = layer4_outputs[160];
    assign outputs[2042] = (layer4_outputs[163]) & ~(layer4_outputs[64]);
    assign outputs[2043] = ~(layer4_outputs[2037]);
    assign outputs[2044] = ~(layer4_outputs[837]);
    assign outputs[2045] = ~(layer4_outputs[2248]);
    assign outputs[2046] = ~(layer4_outputs[2251]);
    assign outputs[2047] = layer4_outputs[1089];
    assign outputs[2048] = layer4_outputs[431];
    assign outputs[2049] = (layer4_outputs[1536]) | (layer4_outputs[2137]);
    assign outputs[2050] = (layer4_outputs[1491]) & ~(layer4_outputs[1100]);
    assign outputs[2051] = ~(layer4_outputs[162]);
    assign outputs[2052] = layer4_outputs[1080];
    assign outputs[2053] = ~((layer4_outputs[1222]) ^ (layer4_outputs[2083]));
    assign outputs[2054] = (layer4_outputs[313]) & (layer4_outputs[347]);
    assign outputs[2055] = layer4_outputs[1261];
    assign outputs[2056] = ~(layer4_outputs[1666]);
    assign outputs[2057] = layer4_outputs[1491];
    assign outputs[2058] = ~(layer4_outputs[43]);
    assign outputs[2059] = (layer4_outputs[45]) & (layer4_outputs[2352]);
    assign outputs[2060] = ~(layer4_outputs[1644]);
    assign outputs[2061] = layer4_outputs[770];
    assign outputs[2062] = ~(layer4_outputs[1686]) | (layer4_outputs[1554]);
    assign outputs[2063] = ~(layer4_outputs[1593]);
    assign outputs[2064] = ~(layer4_outputs[84]);
    assign outputs[2065] = ~(layer4_outputs[241]);
    assign outputs[2066] = ~(layer4_outputs[2176]);
    assign outputs[2067] = ~(layer4_outputs[1849]);
    assign outputs[2068] = layer4_outputs[2507];
    assign outputs[2069] = ~(layer4_outputs[2093]);
    assign outputs[2070] = layer4_outputs[766];
    assign outputs[2071] = ~(layer4_outputs[2553]) | (layer4_outputs[1678]);
    assign outputs[2072] = (layer4_outputs[1347]) & ~(layer4_outputs[145]);
    assign outputs[2073] = ~(layer4_outputs[2365]);
    assign outputs[2074] = layer4_outputs[713];
    assign outputs[2075] = ~(layer4_outputs[2168]);
    assign outputs[2076] = layer4_outputs[1499];
    assign outputs[2077] = ~(layer4_outputs[1668]);
    assign outputs[2078] = layer4_outputs[1724];
    assign outputs[2079] = (layer4_outputs[737]) & (layer4_outputs[2475]);
    assign outputs[2080] = ~(layer4_outputs[290]);
    assign outputs[2081] = layer4_outputs[810];
    assign outputs[2082] = layer4_outputs[309];
    assign outputs[2083] = ~(layer4_outputs[2088]) | (layer4_outputs[741]);
    assign outputs[2084] = ~(layer4_outputs[2517]);
    assign outputs[2085] = ~(layer4_outputs[2457]) | (layer4_outputs[1660]);
    assign outputs[2086] = ~(layer4_outputs[2338]);
    assign outputs[2087] = ~((layer4_outputs[343]) | (layer4_outputs[2257]));
    assign outputs[2088] = (layer4_outputs[760]) & (layer4_outputs[1283]);
    assign outputs[2089] = ~(layer4_outputs[2396]);
    assign outputs[2090] = layer4_outputs[194];
    assign outputs[2091] = layer4_outputs[738];
    assign outputs[2092] = (layer4_outputs[921]) & ~(layer4_outputs[71]);
    assign outputs[2093] = layer4_outputs[843];
    assign outputs[2094] = ~(layer4_outputs[22]);
    assign outputs[2095] = (layer4_outputs[121]) ^ (layer4_outputs[1294]);
    assign outputs[2096] = ~(layer4_outputs[282]);
    assign outputs[2097] = ~(layer4_outputs[1548]);
    assign outputs[2098] = ~(layer4_outputs[1990]) | (layer4_outputs[2076]);
    assign outputs[2099] = (layer4_outputs[2392]) ^ (layer4_outputs[494]);
    assign outputs[2100] = ~(layer4_outputs[2321]);
    assign outputs[2101] = (layer4_outputs[1980]) ^ (layer4_outputs[1138]);
    assign outputs[2102] = ~(layer4_outputs[1849]);
    assign outputs[2103] = ~(layer4_outputs[1051]);
    assign outputs[2104] = layer4_outputs[1292];
    assign outputs[2105] = layer4_outputs[1738];
    assign outputs[2106] = ~(layer4_outputs[749]);
    assign outputs[2107] = (layer4_outputs[1767]) ^ (layer4_outputs[2490]);
    assign outputs[2108] = (layer4_outputs[1893]) & ~(layer4_outputs[62]);
    assign outputs[2109] = layer4_outputs[1625];
    assign outputs[2110] = ~(layer4_outputs[176]);
    assign outputs[2111] = ~(layer4_outputs[749]);
    assign outputs[2112] = layer4_outputs[738];
    assign outputs[2113] = (layer4_outputs[403]) ^ (layer4_outputs[1001]);
    assign outputs[2114] = layer4_outputs[2249];
    assign outputs[2115] = ~(layer4_outputs[684]);
    assign outputs[2116] = ~((layer4_outputs[155]) ^ (layer4_outputs[1412]));
    assign outputs[2117] = (layer4_outputs[2363]) ^ (layer4_outputs[677]);
    assign outputs[2118] = (layer4_outputs[1269]) & (layer4_outputs[471]);
    assign outputs[2119] = ~(layer4_outputs[1171]);
    assign outputs[2120] = ~(layer4_outputs[444]);
    assign outputs[2121] = (layer4_outputs[1983]) & (layer4_outputs[1228]);
    assign outputs[2122] = ~(layer4_outputs[1708]);
    assign outputs[2123] = ~(layer4_outputs[217]);
    assign outputs[2124] = ~(layer4_outputs[127]);
    assign outputs[2125] = ~(layer4_outputs[304]);
    assign outputs[2126] = ~(layer4_outputs[1763]);
    assign outputs[2127] = ~(layer4_outputs[1431]);
    assign outputs[2128] = ~(layer4_outputs[2316]) | (layer4_outputs[2469]);
    assign outputs[2129] = ~((layer4_outputs[2470]) | (layer4_outputs[530]));
    assign outputs[2130] = layer4_outputs[2522];
    assign outputs[2131] = (layer4_outputs[503]) & (layer4_outputs[1577]);
    assign outputs[2132] = ~(layer4_outputs[800]);
    assign outputs[2133] = ~((layer4_outputs[1967]) ^ (layer4_outputs[2269]));
    assign outputs[2134] = (layer4_outputs[156]) ^ (layer4_outputs[2205]);
    assign outputs[2135] = ~(layer4_outputs[2105]);
    assign outputs[2136] = layer4_outputs[5];
    assign outputs[2137] = layer4_outputs[1120];
    assign outputs[2138] = ~((layer4_outputs[969]) & (layer4_outputs[687]));
    assign outputs[2139] = layer4_outputs[1039];
    assign outputs[2140] = layer4_outputs[1268];
    assign outputs[2141] = ~(layer4_outputs[2238]);
    assign outputs[2142] = ~((layer4_outputs[2521]) ^ (layer4_outputs[56]));
    assign outputs[2143] = ~(layer4_outputs[2082]);
    assign outputs[2144] = layer4_outputs[1062];
    assign outputs[2145] = ~((layer4_outputs[1200]) ^ (layer4_outputs[65]));
    assign outputs[2146] = layer4_outputs[1831];
    assign outputs[2147] = layer4_outputs[701];
    assign outputs[2148] = (layer4_outputs[1907]) & (layer4_outputs[1650]);
    assign outputs[2149] = layer4_outputs[1145];
    assign outputs[2150] = ~(layer4_outputs[2166]);
    assign outputs[2151] = ~(layer4_outputs[1378]);
    assign outputs[2152] = ~(layer4_outputs[2033]);
    assign outputs[2153] = layer4_outputs[1112];
    assign outputs[2154] = (layer4_outputs[239]) ^ (layer4_outputs[1181]);
    assign outputs[2155] = ~((layer4_outputs[377]) ^ (layer4_outputs[1444]));
    assign outputs[2156] = layer4_outputs[1610];
    assign outputs[2157] = ~(layer4_outputs[1166]);
    assign outputs[2158] = ~(layer4_outputs[1384]);
    assign outputs[2159] = ~(layer4_outputs[1618]);
    assign outputs[2160] = ~((layer4_outputs[598]) ^ (layer4_outputs[1657]));
    assign outputs[2161] = ~(layer4_outputs[1040]) | (layer4_outputs[39]);
    assign outputs[2162] = (layer4_outputs[35]) | (layer4_outputs[1099]);
    assign outputs[2163] = ~(layer4_outputs[214]);
    assign outputs[2164] = layer4_outputs[223];
    assign outputs[2165] = layer4_outputs[1462];
    assign outputs[2166] = ~(layer4_outputs[31]) | (layer4_outputs[1437]);
    assign outputs[2167] = layer4_outputs[1011];
    assign outputs[2168] = layer4_outputs[2099];
    assign outputs[2169] = ~(layer4_outputs[295]);
    assign outputs[2170] = ~(layer4_outputs[1063]);
    assign outputs[2171] = ~((layer4_outputs[510]) ^ (layer4_outputs[1015]));
    assign outputs[2172] = ~((layer4_outputs[720]) | (layer4_outputs[926]));
    assign outputs[2173] = layer4_outputs[66];
    assign outputs[2174] = ~(layer4_outputs[132]);
    assign outputs[2175] = ~(layer4_outputs[1551]) | (layer4_outputs[2503]);
    assign outputs[2176] = layer4_outputs[865];
    assign outputs[2177] = ~(layer4_outputs[846]) | (layer4_outputs[1238]);
    assign outputs[2178] = ~(layer4_outputs[864]);
    assign outputs[2179] = ~((layer4_outputs[1779]) ^ (layer4_outputs[1052]));
    assign outputs[2180] = ~((layer4_outputs[1988]) | (layer4_outputs[139]));
    assign outputs[2181] = ~(layer4_outputs[2159]);
    assign outputs[2182] = layer4_outputs[165];
    assign outputs[2183] = layer4_outputs[2175];
    assign outputs[2184] = ~(layer4_outputs[2547]) | (layer4_outputs[1206]);
    assign outputs[2185] = (layer4_outputs[848]) ^ (layer4_outputs[272]);
    assign outputs[2186] = layer4_outputs[15];
    assign outputs[2187] = layer4_outputs[1761];
    assign outputs[2188] = layer4_outputs[562];
    assign outputs[2189] = ~(layer4_outputs[2225]) | (layer4_outputs[2112]);
    assign outputs[2190] = layer4_outputs[897];
    assign outputs[2191] = (layer4_outputs[2078]) & ~(layer4_outputs[690]);
    assign outputs[2192] = ~(layer4_outputs[667]) | (layer4_outputs[920]);
    assign outputs[2193] = layer4_outputs[1497];
    assign outputs[2194] = ~((layer4_outputs[1407]) ^ (layer4_outputs[2439]));
    assign outputs[2195] = (layer4_outputs[823]) & (layer4_outputs[51]);
    assign outputs[2196] = ~(layer4_outputs[1013]);
    assign outputs[2197] = layer4_outputs[647];
    assign outputs[2198] = ~((layer4_outputs[1918]) ^ (layer4_outputs[2330]));
    assign outputs[2199] = ~(layer4_outputs[888]);
    assign outputs[2200] = layer4_outputs[1457];
    assign outputs[2201] = ~(layer4_outputs[1903]);
    assign outputs[2202] = (layer4_outputs[181]) ^ (layer4_outputs[1703]);
    assign outputs[2203] = ~(layer4_outputs[1768]);
    assign outputs[2204] = ~(layer4_outputs[179]) | (layer4_outputs[94]);
    assign outputs[2205] = (layer4_outputs[1889]) ^ (layer4_outputs[2009]);
    assign outputs[2206] = ~((layer4_outputs[1409]) | (layer4_outputs[536]));
    assign outputs[2207] = ~(layer4_outputs[1968]);
    assign outputs[2208] = layer4_outputs[2120];
    assign outputs[2209] = ~(layer4_outputs[137]);
    assign outputs[2210] = ~(layer4_outputs[2378]);
    assign outputs[2211] = layer4_outputs[1839];
    assign outputs[2212] = layer4_outputs[2066];
    assign outputs[2213] = (layer4_outputs[38]) & ~(layer4_outputs[1519]);
    assign outputs[2214] = ~(layer4_outputs[1853]);
    assign outputs[2215] = ~(layer4_outputs[271]);
    assign outputs[2216] = layer4_outputs[708];
    assign outputs[2217] = ~(layer4_outputs[512]);
    assign outputs[2218] = ~(layer4_outputs[433]);
    assign outputs[2219] = ~(layer4_outputs[1216]);
    assign outputs[2220] = (layer4_outputs[2350]) ^ (layer4_outputs[879]);
    assign outputs[2221] = (layer4_outputs[1585]) & ~(layer4_outputs[2206]);
    assign outputs[2222] = ~((layer4_outputs[228]) ^ (layer4_outputs[362]));
    assign outputs[2223] = ~(layer4_outputs[1672]);
    assign outputs[2224] = ~((layer4_outputs[572]) | (layer4_outputs[233]));
    assign outputs[2225] = layer4_outputs[392];
    assign outputs[2226] = layer4_outputs[2522];
    assign outputs[2227] = ~(layer4_outputs[1721]);
    assign outputs[2228] = layer4_outputs[755];
    assign outputs[2229] = ~(layer4_outputs[981]);
    assign outputs[2230] = layer4_outputs[1269];
    assign outputs[2231] = ~(layer4_outputs[912]);
    assign outputs[2232] = layer4_outputs[2480];
    assign outputs[2233] = (layer4_outputs[1727]) & ~(layer4_outputs[1328]);
    assign outputs[2234] = ~(layer4_outputs[2102]);
    assign outputs[2235] = ~(layer4_outputs[2357]);
    assign outputs[2236] = layer4_outputs[647];
    assign outputs[2237] = (layer4_outputs[1371]) & ~(layer4_outputs[451]);
    assign outputs[2238] = ~(layer4_outputs[2538]);
    assign outputs[2239] = layer4_outputs[732];
    assign outputs[2240] = ~((layer4_outputs[517]) | (layer4_outputs[128]));
    assign outputs[2241] = ~(layer4_outputs[1190]) | (layer4_outputs[2113]);
    assign outputs[2242] = layer4_outputs[2285];
    assign outputs[2243] = ~(layer4_outputs[180]);
    assign outputs[2244] = ~(layer4_outputs[115]);
    assign outputs[2245] = ~((layer4_outputs[55]) | (layer4_outputs[765]));
    assign outputs[2246] = (layer4_outputs[112]) ^ (layer4_outputs[1265]);
    assign outputs[2247] = ~(layer4_outputs[1130]);
    assign outputs[2248] = layer4_outputs[847];
    assign outputs[2249] = ~(layer4_outputs[2367]);
    assign outputs[2250] = (layer4_outputs[2146]) & ~(layer4_outputs[1750]);
    assign outputs[2251] = ~(layer4_outputs[426]);
    assign outputs[2252] = layer4_outputs[2550];
    assign outputs[2253] = (layer4_outputs[551]) & (layer4_outputs[338]);
    assign outputs[2254] = layer4_outputs[1813];
    assign outputs[2255] = ~(layer4_outputs[530]);
    assign outputs[2256] = ~(layer4_outputs[1780]);
    assign outputs[2257] = (layer4_outputs[860]) ^ (layer4_outputs[1255]);
    assign outputs[2258] = (layer4_outputs[2209]) ^ (layer4_outputs[1706]);
    assign outputs[2259] = ~(layer4_outputs[1005]);
    assign outputs[2260] = ~(layer4_outputs[1716]);
    assign outputs[2261] = ~((layer4_outputs[2225]) ^ (layer4_outputs[1279]));
    assign outputs[2262] = layer4_outputs[131];
    assign outputs[2263] = ~(layer4_outputs[778]);
    assign outputs[2264] = (layer4_outputs[2116]) & ~(layer4_outputs[2018]);
    assign outputs[2265] = ~((layer4_outputs[245]) ^ (layer4_outputs[202]));
    assign outputs[2266] = ~((layer4_outputs[196]) ^ (layer4_outputs[197]));
    assign outputs[2267] = ~(layer4_outputs[1571]);
    assign outputs[2268] = layer4_outputs[642];
    assign outputs[2269] = ~(layer4_outputs[342]);
    assign outputs[2270] = layer4_outputs[2241];
    assign outputs[2271] = ~(layer4_outputs[1025]);
    assign outputs[2272] = layer4_outputs[317];
    assign outputs[2273] = ~(layer4_outputs[1728]);
    assign outputs[2274] = (layer4_outputs[2143]) | (layer4_outputs[1364]);
    assign outputs[2275] = (layer4_outputs[325]) ^ (layer4_outputs[2437]);
    assign outputs[2276] = layer4_outputs[2121];
    assign outputs[2277] = (layer4_outputs[1147]) ^ (layer4_outputs[109]);
    assign outputs[2278] = ~(layer4_outputs[1737]) | (layer4_outputs[2143]);
    assign outputs[2279] = (layer4_outputs[1932]) ^ (layer4_outputs[2131]);
    assign outputs[2280] = ~((layer4_outputs[1767]) ^ (layer4_outputs[52]));
    assign outputs[2281] = (layer4_outputs[11]) ^ (layer4_outputs[148]);
    assign outputs[2282] = ~(layer4_outputs[300]);
    assign outputs[2283] = layer4_outputs[1704];
    assign outputs[2284] = layer4_outputs[2065];
    assign outputs[2285] = ~(layer4_outputs[1327]);
    assign outputs[2286] = (layer4_outputs[1885]) ^ (layer4_outputs[1586]);
    assign outputs[2287] = ~(layer4_outputs[2179]);
    assign outputs[2288] = (layer4_outputs[80]) & ~(layer4_outputs[485]);
    assign outputs[2289] = layer4_outputs[2311];
    assign outputs[2290] = (layer4_outputs[1395]) & ~(layer4_outputs[259]);
    assign outputs[2291] = layer4_outputs[2122];
    assign outputs[2292] = layer4_outputs[645];
    assign outputs[2293] = ~(layer4_outputs[986]);
    assign outputs[2294] = layer4_outputs[1876];
    assign outputs[2295] = (layer4_outputs[2177]) & ~(layer4_outputs[1187]);
    assign outputs[2296] = (layer4_outputs[2253]) ^ (layer4_outputs[2465]);
    assign outputs[2297] = ~((layer4_outputs[1065]) | (layer4_outputs[900]));
    assign outputs[2298] = (layer4_outputs[2237]) ^ (layer4_outputs[1782]);
    assign outputs[2299] = layer4_outputs[98];
    assign outputs[2300] = ~((layer4_outputs[1780]) | (layer4_outputs[152]));
    assign outputs[2301] = ~((layer4_outputs[1402]) | (layer4_outputs[318]));
    assign outputs[2302] = ~((layer4_outputs[1533]) ^ (layer4_outputs[2221]));
    assign outputs[2303] = ~(layer4_outputs[2003]);
    assign outputs[2304] = ~((layer4_outputs[591]) ^ (layer4_outputs[1493]));
    assign outputs[2305] = layer4_outputs[2115];
    assign outputs[2306] = ~(layer4_outputs[2218]);
    assign outputs[2307] = (layer4_outputs[1063]) & (layer4_outputs[268]);
    assign outputs[2308] = layer4_outputs[2278];
    assign outputs[2309] = layer4_outputs[2526];
    assign outputs[2310] = layer4_outputs[593];
    assign outputs[2311] = (layer4_outputs[204]) & ~(layer4_outputs[2040]);
    assign outputs[2312] = (layer4_outputs[1796]) & ~(layer4_outputs[304]);
    assign outputs[2313] = layer4_outputs[1223];
    assign outputs[2314] = layer4_outputs[966];
    assign outputs[2315] = ~((layer4_outputs[1021]) | (layer4_outputs[939]));
    assign outputs[2316] = ~((layer4_outputs[1817]) ^ (layer4_outputs[2404]));
    assign outputs[2317] = ~(layer4_outputs[1874]);
    assign outputs[2318] = ~(layer4_outputs[900]);
    assign outputs[2319] = (layer4_outputs[871]) ^ (layer4_outputs[2313]);
    assign outputs[2320] = (layer4_outputs[2095]) & (layer4_outputs[1189]);
    assign outputs[2321] = layer4_outputs[1649];
    assign outputs[2322] = ~(layer4_outputs[2316]);
    assign outputs[2323] = (layer4_outputs[1353]) & ~(layer4_outputs[1510]);
    assign outputs[2324] = layer4_outputs[1569];
    assign outputs[2325] = layer4_outputs[1560];
    assign outputs[2326] = ~((layer4_outputs[1948]) ^ (layer4_outputs[954]));
    assign outputs[2327] = ~((layer4_outputs[443]) ^ (layer4_outputs[1081]));
    assign outputs[2328] = ~(layer4_outputs[1939]);
    assign outputs[2329] = ~((layer4_outputs[1552]) ^ (layer4_outputs[1446]));
    assign outputs[2330] = layer4_outputs[9];
    assign outputs[2331] = ~(layer4_outputs[1637]);
    assign outputs[2332] = ~(layer4_outputs[2355]);
    assign outputs[2333] = ~((layer4_outputs[171]) | (layer4_outputs[2412]));
    assign outputs[2334] = ~(layer4_outputs[1440]);
    assign outputs[2335] = ~(layer4_outputs[297]);
    assign outputs[2336] = ~(layer4_outputs[2390]);
    assign outputs[2337] = ~(layer4_outputs[2071]);
    assign outputs[2338] = ~(layer4_outputs[1987]);
    assign outputs[2339] = layer4_outputs[487];
    assign outputs[2340] = (layer4_outputs[2240]) & (layer4_outputs[1282]);
    assign outputs[2341] = layer4_outputs[2459];
    assign outputs[2342] = (layer4_outputs[1292]) | (layer4_outputs[2158]);
    assign outputs[2343] = (layer4_outputs[2199]) & ~(layer4_outputs[957]);
    assign outputs[2344] = layer4_outputs[2410];
    assign outputs[2345] = ~(layer4_outputs[948]);
    assign outputs[2346] = layer4_outputs[2406];
    assign outputs[2347] = layer4_outputs[2370];
    assign outputs[2348] = ~(layer4_outputs[2331]);
    assign outputs[2349] = ~((layer4_outputs[1423]) & (layer4_outputs[144]));
    assign outputs[2350] = layer4_outputs[2013];
    assign outputs[2351] = (layer4_outputs[2535]) & ~(layer4_outputs[2193]);
    assign outputs[2352] = ~((layer4_outputs[199]) | (layer4_outputs[2059]));
    assign outputs[2353] = layer4_outputs[2400];
    assign outputs[2354] = ~((layer4_outputs[584]) ^ (layer4_outputs[2531]));
    assign outputs[2355] = ~((layer4_outputs[1863]) ^ (layer4_outputs[1664]));
    assign outputs[2356] = ~(layer4_outputs[805]);
    assign outputs[2357] = ~(layer4_outputs[1004]);
    assign outputs[2358] = ~(layer4_outputs[1412]);
    assign outputs[2359] = (layer4_outputs[36]) & ~(layer4_outputs[839]);
    assign outputs[2360] = ~((layer4_outputs[1379]) ^ (layer4_outputs[2012]));
    assign outputs[2361] = (layer4_outputs[969]) & (layer4_outputs[1228]);
    assign outputs[2362] = ~((layer4_outputs[1405]) & (layer4_outputs[2268]));
    assign outputs[2363] = (layer4_outputs[418]) ^ (layer4_outputs[2275]);
    assign outputs[2364] = (layer4_outputs[1141]) ^ (layer4_outputs[1391]);
    assign outputs[2365] = layer4_outputs[2398];
    assign outputs[2366] = ~(layer4_outputs[2539]);
    assign outputs[2367] = layer4_outputs[1471];
    assign outputs[2368] = ~((layer4_outputs[449]) ^ (layer4_outputs[1692]));
    assign outputs[2369] = (layer4_outputs[1525]) & ~(layer4_outputs[199]);
    assign outputs[2370] = ~((layer4_outputs[326]) | (layer4_outputs[510]));
    assign outputs[2371] = layer4_outputs[736];
    assign outputs[2372] = ~(layer4_outputs[2071]);
    assign outputs[2373] = (layer4_outputs[1914]) & ~(layer4_outputs[1511]);
    assign outputs[2374] = (layer4_outputs[1436]) ^ (layer4_outputs[2519]);
    assign outputs[2375] = ~((layer4_outputs[753]) ^ (layer4_outputs[1208]));
    assign outputs[2376] = layer4_outputs[575];
    assign outputs[2377] = layer4_outputs[1578];
    assign outputs[2378] = (layer4_outputs[328]) & ~(layer4_outputs[670]);
    assign outputs[2379] = ~(layer4_outputs[1116]);
    assign outputs[2380] = layer4_outputs[1337];
    assign outputs[2381] = layer4_outputs[2311];
    assign outputs[2382] = (layer4_outputs[2340]) ^ (layer4_outputs[1117]);
    assign outputs[2383] = ~((layer4_outputs[2525]) | (layer4_outputs[546]));
    assign outputs[2384] = ~(layer4_outputs[985]);
    assign outputs[2385] = layer4_outputs[724];
    assign outputs[2386] = (layer4_outputs[1897]) ^ (layer4_outputs[1432]);
    assign outputs[2387] = layer4_outputs[452];
    assign outputs[2388] = layer4_outputs[677];
    assign outputs[2389] = (layer4_outputs[1156]) & ~(layer4_outputs[1826]);
    assign outputs[2390] = layer4_outputs[1957];
    assign outputs[2391] = ~(layer4_outputs[841]);
    assign outputs[2392] = ~(layer4_outputs[630]);
    assign outputs[2393] = layer4_outputs[1686];
    assign outputs[2394] = (layer4_outputs[663]) ^ (layer4_outputs[1010]);
    assign outputs[2395] = (layer4_outputs[9]) & ~(layer4_outputs[1896]);
    assign outputs[2396] = ~(layer4_outputs[2051]);
    assign outputs[2397] = ~(layer4_outputs[610]);
    assign outputs[2398] = ~(layer4_outputs[1959]);
    assign outputs[2399] = ~((layer4_outputs[1662]) ^ (layer4_outputs[1095]));
    assign outputs[2400] = ~((layer4_outputs[1737]) ^ (layer4_outputs[2035]));
    assign outputs[2401] = (layer4_outputs[844]) & ~(layer4_outputs[225]);
    assign outputs[2402] = ~((layer4_outputs[1389]) ^ (layer4_outputs[2410]));
    assign outputs[2403] = layer4_outputs[2381];
    assign outputs[2404] = layer4_outputs[1604];
    assign outputs[2405] = (layer4_outputs[1818]) & ~(layer4_outputs[1753]);
    assign outputs[2406] = ~((layer4_outputs[1054]) ^ (layer4_outputs[117]));
    assign outputs[2407] = ~(layer4_outputs[1069]) | (layer4_outputs[1454]);
    assign outputs[2408] = (layer4_outputs[127]) & ~(layer4_outputs[770]);
    assign outputs[2409] = (layer4_outputs[426]) ^ (layer4_outputs[673]);
    assign outputs[2410] = ~(layer4_outputs[713]);
    assign outputs[2411] = (layer4_outputs[1804]) & ~(layer4_outputs[1681]);
    assign outputs[2412] = layer4_outputs[2127];
    assign outputs[2413] = (layer4_outputs[2341]) & ~(layer4_outputs[1463]);
    assign outputs[2414] = ~((layer4_outputs[2331]) | (layer4_outputs[13]));
    assign outputs[2415] = ~(layer4_outputs[909]);
    assign outputs[2416] = (layer4_outputs[465]) & ~(layer4_outputs[792]);
    assign outputs[2417] = ~((layer4_outputs[2059]) | (layer4_outputs[2390]));
    assign outputs[2418] = ~((layer4_outputs[376]) | (layer4_outputs[1473]));
    assign outputs[2419] = ~(layer4_outputs[1116]);
    assign outputs[2420] = (layer4_outputs[1143]) & (layer4_outputs[2344]);
    assign outputs[2421] = ~(layer4_outputs[1912]);
    assign outputs[2422] = ~(layer4_outputs[609]);
    assign outputs[2423] = (layer4_outputs[716]) ^ (layer4_outputs[1409]);
    assign outputs[2424] = ~(layer4_outputs[1939]);
    assign outputs[2425] = ~(layer4_outputs[1772]);
    assign outputs[2426] = (layer4_outputs[961]) ^ (layer4_outputs[1085]);
    assign outputs[2427] = ~((layer4_outputs[1975]) | (layer4_outputs[659]));
    assign outputs[2428] = layer4_outputs[1290];
    assign outputs[2429] = (layer4_outputs[2417]) & (layer4_outputs[1751]);
    assign outputs[2430] = layer4_outputs[1387];
    assign outputs[2431] = ~(layer4_outputs[135]);
    assign outputs[2432] = ~(layer4_outputs[1060]);
    assign outputs[2433] = ~((layer4_outputs[1895]) ^ (layer4_outputs[454]));
    assign outputs[2434] = ~(layer4_outputs[678]);
    assign outputs[2435] = (layer4_outputs[514]) ^ (layer4_outputs[1809]);
    assign outputs[2436] = ~(layer4_outputs[2189]);
    assign outputs[2437] = ~(layer4_outputs[341]);
    assign outputs[2438] = layer4_outputs[1453];
    assign outputs[2439] = ~((layer4_outputs[2153]) ^ (layer4_outputs[878]));
    assign outputs[2440] = layer4_outputs[73];
    assign outputs[2441] = ~(layer4_outputs[1295]);
    assign outputs[2442] = (layer4_outputs[1675]) & (layer4_outputs[2216]);
    assign outputs[2443] = layer4_outputs[1570];
    assign outputs[2444] = ~((layer4_outputs[376]) | (layer4_outputs[0]));
    assign outputs[2445] = ~(layer4_outputs[213]);
    assign outputs[2446] = ~(layer4_outputs[2250]);
    assign outputs[2447] = ~((layer4_outputs[1110]) ^ (layer4_outputs[1430]));
    assign outputs[2448] = ~(layer4_outputs[1433]);
    assign outputs[2449] = ~((layer4_outputs[1380]) & (layer4_outputs[428]));
    assign outputs[2450] = ~((layer4_outputs[1930]) | (layer4_outputs[1840]));
    assign outputs[2451] = (layer4_outputs[1383]) & ~(layer4_outputs[205]);
    assign outputs[2452] = ~((layer4_outputs[1487]) ^ (layer4_outputs[416]));
    assign outputs[2453] = ~(layer4_outputs[787]);
    assign outputs[2454] = ~(layer4_outputs[312]);
    assign outputs[2455] = layer4_outputs[1023];
    assign outputs[2456] = layer4_outputs[1214];
    assign outputs[2457] = ~(layer4_outputs[1842]);
    assign outputs[2458] = layer4_outputs[1557];
    assign outputs[2459] = layer4_outputs[818];
    assign outputs[2460] = ~(layer4_outputs[1975]);
    assign outputs[2461] = ~(layer4_outputs[1004]);
    assign outputs[2462] = ~(layer4_outputs[1776]);
    assign outputs[2463] = layer4_outputs[393];
    assign outputs[2464] = layer4_outputs[1231];
    assign outputs[2465] = ~(layer4_outputs[801]);
    assign outputs[2466] = ~((layer4_outputs[1003]) | (layer4_outputs[1677]));
    assign outputs[2467] = ~(layer4_outputs[1262]);
    assign outputs[2468] = layer4_outputs[1795];
    assign outputs[2469] = (layer4_outputs[1705]) ^ (layer4_outputs[1710]);
    assign outputs[2470] = layer4_outputs[476];
    assign outputs[2471] = ~(layer4_outputs[1070]);
    assign outputs[2472] = layer4_outputs[1963];
    assign outputs[2473] = layer4_outputs[1697];
    assign outputs[2474] = ~(layer4_outputs[1154]);
    assign outputs[2475] = ~((layer4_outputs[484]) | (layer4_outputs[1599]));
    assign outputs[2476] = ~(layer4_outputs[1611]);
    assign outputs[2477] = ~(layer4_outputs[187]);
    assign outputs[2478] = layer4_outputs[1404];
    assign outputs[2479] = (layer4_outputs[1562]) & ~(layer4_outputs[958]);
    assign outputs[2480] = layer4_outputs[1268];
    assign outputs[2481] = layer4_outputs[1034];
    assign outputs[2482] = ~(layer4_outputs[2387]);
    assign outputs[2483] = layer4_outputs[270];
    assign outputs[2484] = (layer4_outputs[397]) & ~(layer4_outputs[436]);
    assign outputs[2485] = (layer4_outputs[116]) & (layer4_outputs[589]);
    assign outputs[2486] = layer4_outputs[357];
    assign outputs[2487] = (layer4_outputs[987]) & (layer4_outputs[597]);
    assign outputs[2488] = ~(layer4_outputs[16]);
    assign outputs[2489] = layer4_outputs[763];
    assign outputs[2490] = ~(layer4_outputs[341]);
    assign outputs[2491] = layer4_outputs[2023];
    assign outputs[2492] = ~((layer4_outputs[1257]) ^ (layer4_outputs[280]));
    assign outputs[2493] = ~(layer4_outputs[2064]);
    assign outputs[2494] = layer4_outputs[2204];
    assign outputs[2495] = layer4_outputs[574];
    assign outputs[2496] = (layer4_outputs[874]) & ~(layer4_outputs[1192]);
    assign outputs[2497] = ~(layer4_outputs[638]);
    assign outputs[2498] = ~(layer4_outputs[1310]);
    assign outputs[2499] = layer4_outputs[663];
    assign outputs[2500] = (layer4_outputs[1502]) ^ (layer4_outputs[682]);
    assign outputs[2501] = (layer4_outputs[1365]) & (layer4_outputs[1270]);
    assign outputs[2502] = layer4_outputs[1865];
    assign outputs[2503] = layer4_outputs[360];
    assign outputs[2504] = ~(layer4_outputs[20]);
    assign outputs[2505] = (layer4_outputs[2513]) ^ (layer4_outputs[2216]);
    assign outputs[2506] = (layer4_outputs[657]) ^ (layer4_outputs[403]);
    assign outputs[2507] = layer4_outputs[1515];
    assign outputs[2508] = ~(layer4_outputs[990]);
    assign outputs[2509] = (layer4_outputs[1489]) & ~(layer4_outputs[1640]);
    assign outputs[2510] = layer4_outputs[440];
    assign outputs[2511] = layer4_outputs[979];
    assign outputs[2512] = ~(layer4_outputs[2273]);
    assign outputs[2513] = layer4_outputs[469];
    assign outputs[2514] = ~((layer4_outputs[717]) ^ (layer4_outputs[1945]));
    assign outputs[2515] = (layer4_outputs[459]) & ~(layer4_outputs[343]);
    assign outputs[2516] = layer4_outputs[160];
    assign outputs[2517] = ~(layer4_outputs[986]);
    assign outputs[2518] = ~((layer4_outputs[641]) | (layer4_outputs[240]));
    assign outputs[2519] = ~((layer4_outputs[1539]) | (layer4_outputs[2098]));
    assign outputs[2520] = layer4_outputs[1864];
    assign outputs[2521] = (layer4_outputs[1351]) ^ (layer4_outputs[133]);
    assign outputs[2522] = ~((layer4_outputs[565]) ^ (layer4_outputs[1751]));
    assign outputs[2523] = layer4_outputs[2148];
    assign outputs[2524] = (layer4_outputs[812]) ^ (layer4_outputs[2351]);
    assign outputs[2525] = (layer4_outputs[1486]) ^ (layer4_outputs[87]);
    assign outputs[2526] = layer4_outputs[437];
    assign outputs[2527] = ~((layer4_outputs[2104]) ^ (layer4_outputs[2167]));
    assign outputs[2528] = ~(layer4_outputs[867]);
    assign outputs[2529] = ~((layer4_outputs[1030]) | (layer4_outputs[2201]));
    assign outputs[2530] = layer4_outputs[632];
    assign outputs[2531] = layer4_outputs[70];
    assign outputs[2532] = layer4_outputs[1856];
    assign outputs[2533] = layer4_outputs[799];
    assign outputs[2534] = (layer4_outputs[1581]) & ~(layer4_outputs[1340]);
    assign outputs[2535] = (layer4_outputs[399]) & ~(layer4_outputs[570]);
    assign outputs[2536] = ~((layer4_outputs[147]) | (layer4_outputs[563]));
    assign outputs[2537] = ~(layer4_outputs[1553]);
    assign outputs[2538] = (layer4_outputs[573]) ^ (layer4_outputs[1701]);
    assign outputs[2539] = (layer4_outputs[191]) ^ (layer4_outputs[1905]);
    assign outputs[2540] = ~(layer4_outputs[138]);
    assign outputs[2541] = layer4_outputs[2553];
    assign outputs[2542] = (layer4_outputs[1676]) & ~(layer4_outputs[1167]);
    assign outputs[2543] = ~(layer4_outputs[610]);
    assign outputs[2544] = layer4_outputs[79];
    assign outputs[2545] = (layer4_outputs[2457]) ^ (layer4_outputs[982]);
    assign outputs[2546] = (layer4_outputs[1665]) | (layer4_outputs[1267]);
    assign outputs[2547] = layer4_outputs[538];
    assign outputs[2548] = ~(layer4_outputs[355]);
    assign outputs[2549] = ~(layer4_outputs[334]);
    assign outputs[2550] = layer4_outputs[2413];
    assign outputs[2551] = (layer4_outputs[1226]) & (layer4_outputs[832]);
    assign outputs[2552] = layer4_outputs[1034];
    assign outputs[2553] = (layer4_outputs[907]) & (layer4_outputs[1155]);
    assign outputs[2554] = layer4_outputs[946];
    assign outputs[2555] = layer4_outputs[2278];
    assign outputs[2556] = layer4_outputs[1562];
    assign outputs[2557] = layer4_outputs[1248];
    assign outputs[2558] = ~(layer4_outputs[2234]) | (layer4_outputs[894]);
    assign outputs[2559] = (layer4_outputs[389]) ^ (layer4_outputs[577]);
endmodule
