library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs : in std_logic_vector(255 downto 0);
        outputs : out std_logic_vector(9 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs : std_logic_vector(10239 downto 0);

begin

    layer0_outputs(0) <= (inputs(184)) and not (inputs(213));
    layer0_outputs(1) <= not((inputs(75)) xor (inputs(165)));
    layer0_outputs(2) <= (inputs(254)) and not (inputs(49));
    layer0_outputs(3) <= (inputs(185)) or (inputs(155));
    layer0_outputs(4) <= (inputs(83)) xor (inputs(211));
    layer0_outputs(5) <= not((inputs(109)) or (inputs(255)));
    layer0_outputs(6) <= inputs(221);
    layer0_outputs(7) <= (inputs(111)) or (inputs(115));
    layer0_outputs(8) <= not((inputs(158)) xor (inputs(202)));
    layer0_outputs(9) <= not((inputs(239)) and (inputs(113)));
    layer0_outputs(10) <= (inputs(37)) or (inputs(51));
    layer0_outputs(11) <= not(inputs(37)) or (inputs(140));
    layer0_outputs(12) <= (inputs(107)) or (inputs(234));
    layer0_outputs(13) <= (inputs(232)) and not (inputs(52));
    layer0_outputs(14) <= (inputs(223)) and not (inputs(10));
    layer0_outputs(15) <= not(inputs(164)) or (inputs(210));
    layer0_outputs(16) <= not((inputs(234)) xor (inputs(137)));
    layer0_outputs(17) <= inputs(229);
    layer0_outputs(18) <= inputs(118);
    layer0_outputs(19) <= not(inputs(217)) or (inputs(59));
    layer0_outputs(20) <= not((inputs(96)) xor (inputs(180)));
    layer0_outputs(21) <= inputs(194);
    layer0_outputs(22) <= (inputs(169)) xor (inputs(19));
    layer0_outputs(23) <= (inputs(212)) and not (inputs(44));
    layer0_outputs(24) <= not((inputs(141)) xor (inputs(62)));
    layer0_outputs(25) <= '0';
    layer0_outputs(26) <= not((inputs(164)) or (inputs(167)));
    layer0_outputs(27) <= (inputs(39)) or (inputs(0));
    layer0_outputs(28) <= (inputs(129)) xor (inputs(236));
    layer0_outputs(29) <= (inputs(53)) and not (inputs(95));
    layer0_outputs(30) <= not((inputs(170)) xor (inputs(83)));
    layer0_outputs(31) <= inputs(164);
    layer0_outputs(32) <= not(inputs(118));
    layer0_outputs(33) <= inputs(80);
    layer0_outputs(34) <= not((inputs(135)) or (inputs(129)));
    layer0_outputs(35) <= not((inputs(245)) xor (inputs(141)));
    layer0_outputs(36) <= (inputs(113)) and not (inputs(19));
    layer0_outputs(37) <= (inputs(151)) and not (inputs(112));
    layer0_outputs(38) <= (inputs(155)) or (inputs(253));
    layer0_outputs(39) <= not(inputs(104));
    layer0_outputs(40) <= (inputs(56)) and not (inputs(109));
    layer0_outputs(41) <= not((inputs(59)) xor (inputs(144)));
    layer0_outputs(42) <= not((inputs(182)) or (inputs(142)));
    layer0_outputs(43) <= (inputs(192)) and not (inputs(245));
    layer0_outputs(44) <= (inputs(71)) and (inputs(54));
    layer0_outputs(45) <= (inputs(27)) or (inputs(132));
    layer0_outputs(46) <= (inputs(251)) and (inputs(30));
    layer0_outputs(47) <= '0';
    layer0_outputs(48) <= (inputs(198)) or (inputs(250));
    layer0_outputs(49) <= inputs(55);
    layer0_outputs(50) <= (inputs(124)) and not (inputs(2));
    layer0_outputs(51) <= '1';
    layer0_outputs(52) <= (inputs(93)) and not (inputs(79));
    layer0_outputs(53) <= (inputs(165)) or (inputs(85));
    layer0_outputs(54) <= (inputs(187)) xor (inputs(161));
    layer0_outputs(55) <= not(inputs(95)) or (inputs(237));
    layer0_outputs(56) <= inputs(137);
    layer0_outputs(57) <= not((inputs(240)) and (inputs(245)));
    layer0_outputs(58) <= (inputs(135)) or (inputs(151));
    layer0_outputs(59) <= not((inputs(221)) and (inputs(16)));
    layer0_outputs(60) <= not((inputs(135)) and (inputs(21)));
    layer0_outputs(61) <= (inputs(117)) and not (inputs(83));
    layer0_outputs(62) <= (inputs(9)) xor (inputs(47));
    layer0_outputs(63) <= (inputs(241)) or (inputs(200));
    layer0_outputs(64) <= not(inputs(139)) or (inputs(18));
    layer0_outputs(65) <= not((inputs(120)) or (inputs(195)));
    layer0_outputs(66) <= not((inputs(13)) xor (inputs(74)));
    layer0_outputs(67) <= (inputs(178)) or (inputs(79));
    layer0_outputs(68) <= not((inputs(38)) or (inputs(243)));
    layer0_outputs(69) <= (inputs(87)) and not (inputs(242));
    layer0_outputs(70) <= not(inputs(183));
    layer0_outputs(71) <= not((inputs(52)) xor (inputs(193)));
    layer0_outputs(72) <= not(inputs(189)) or (inputs(167));
    layer0_outputs(73) <= (inputs(179)) xor (inputs(197));
    layer0_outputs(74) <= (inputs(206)) and not (inputs(249));
    layer0_outputs(75) <= not((inputs(200)) xor (inputs(14)));
    layer0_outputs(76) <= not(inputs(232));
    layer0_outputs(77) <= inputs(156);
    layer0_outputs(78) <= inputs(7);
    layer0_outputs(79) <= not((inputs(67)) or (inputs(156)));
    layer0_outputs(80) <= inputs(56);
    layer0_outputs(81) <= (inputs(249)) and not (inputs(193));
    layer0_outputs(82) <= not(inputs(181));
    layer0_outputs(83) <= inputs(122);
    layer0_outputs(84) <= (inputs(223)) and not (inputs(40));
    layer0_outputs(85) <= (inputs(217)) or (inputs(127));
    layer0_outputs(86) <= inputs(207);
    layer0_outputs(87) <= not(inputs(175)) or (inputs(208));
    layer0_outputs(88) <= (inputs(253)) xor (inputs(198));
    layer0_outputs(89) <= not(inputs(119));
    layer0_outputs(90) <= (inputs(113)) or (inputs(138));
    layer0_outputs(91) <= not((inputs(140)) and (inputs(9)));
    layer0_outputs(92) <= inputs(201);
    layer0_outputs(93) <= (inputs(179)) xor (inputs(38));
    layer0_outputs(94) <= inputs(75);
    layer0_outputs(95) <= (inputs(201)) and not (inputs(123));
    layer0_outputs(96) <= not(inputs(46)) or (inputs(5));
    layer0_outputs(97) <= not(inputs(189)) or (inputs(129));
    layer0_outputs(98) <= (inputs(154)) xor (inputs(79));
    layer0_outputs(99) <= not(inputs(188));
    layer0_outputs(100) <= not(inputs(183)) or (inputs(76));
    layer0_outputs(101) <= (inputs(102)) or (inputs(223));
    layer0_outputs(102) <= not((inputs(56)) xor (inputs(25)));
    layer0_outputs(103) <= not((inputs(194)) xor (inputs(239)));
    layer0_outputs(104) <= not((inputs(77)) and (inputs(217)));
    layer0_outputs(105) <= (inputs(185)) or (inputs(21));
    layer0_outputs(106) <= inputs(215);
    layer0_outputs(107) <= '0';
    layer0_outputs(108) <= (inputs(32)) and (inputs(184));
    layer0_outputs(109) <= (inputs(37)) or (inputs(178));
    layer0_outputs(110) <= inputs(34);
    layer0_outputs(111) <= inputs(158);
    layer0_outputs(112) <= (inputs(243)) and (inputs(1));
    layer0_outputs(113) <= not((inputs(77)) or (inputs(103)));
    layer0_outputs(114) <= (inputs(169)) or (inputs(134));
    layer0_outputs(115) <= (inputs(38)) or (inputs(64));
    layer0_outputs(116) <= inputs(166);
    layer0_outputs(117) <= (inputs(211)) or (inputs(138));
    layer0_outputs(118) <= '1';
    layer0_outputs(119) <= inputs(220);
    layer0_outputs(120) <= inputs(7);
    layer0_outputs(121) <= (inputs(248)) or (inputs(107));
    layer0_outputs(122) <= not(inputs(198));
    layer0_outputs(123) <= not(inputs(112)) or (inputs(246));
    layer0_outputs(124) <= not(inputs(244));
    layer0_outputs(125) <= (inputs(236)) and (inputs(144));
    layer0_outputs(126) <= (inputs(183)) or (inputs(242));
    layer0_outputs(127) <= not(inputs(22));
    layer0_outputs(128) <= not((inputs(115)) or (inputs(125)));
    layer0_outputs(129) <= not((inputs(102)) or (inputs(149)));
    layer0_outputs(130) <= '1';
    layer0_outputs(131) <= '0';
    layer0_outputs(132) <= (inputs(132)) and not (inputs(245));
    layer0_outputs(133) <= not(inputs(139)) or (inputs(4));
    layer0_outputs(134) <= inputs(139);
    layer0_outputs(135) <= not(inputs(132)) or (inputs(1));
    layer0_outputs(136) <= (inputs(239)) and not (inputs(2));
    layer0_outputs(137) <= not((inputs(205)) xor (inputs(119)));
    layer0_outputs(138) <= inputs(203);
    layer0_outputs(139) <= (inputs(91)) xor (inputs(69));
    layer0_outputs(140) <= not((inputs(114)) or (inputs(2)));
    layer0_outputs(141) <= (inputs(0)) or (inputs(140));
    layer0_outputs(142) <= not((inputs(205)) xor (inputs(138)));
    layer0_outputs(143) <= (inputs(35)) xor (inputs(123));
    layer0_outputs(144) <= not(inputs(196)) or (inputs(5));
    layer0_outputs(145) <= (inputs(230)) and not (inputs(62));
    layer0_outputs(146) <= not(inputs(74)) or (inputs(99));
    layer0_outputs(147) <= (inputs(62)) and (inputs(125));
    layer0_outputs(148) <= inputs(250);
    layer0_outputs(149) <= (inputs(190)) xor (inputs(30));
    layer0_outputs(150) <= (inputs(214)) and not (inputs(48));
    layer0_outputs(151) <= (inputs(245)) and (inputs(200));
    layer0_outputs(152) <= (inputs(108)) and not (inputs(159));
    layer0_outputs(153) <= (inputs(238)) or (inputs(90));
    layer0_outputs(154) <= (inputs(16)) or (inputs(78));
    layer0_outputs(155) <= not(inputs(180)) or (inputs(40));
    layer0_outputs(156) <= (inputs(245)) xor (inputs(69));
    layer0_outputs(157) <= not(inputs(62));
    layer0_outputs(158) <= (inputs(93)) and not (inputs(124));
    layer0_outputs(159) <= inputs(51);
    layer0_outputs(160) <= inputs(138);
    layer0_outputs(161) <= not((inputs(158)) or (inputs(172)));
    layer0_outputs(162) <= not((inputs(64)) or (inputs(233)));
    layer0_outputs(163) <= not((inputs(18)) xor (inputs(106)));
    layer0_outputs(164) <= not(inputs(136)) or (inputs(27));
    layer0_outputs(165) <= '1';
    layer0_outputs(166) <= inputs(152);
    layer0_outputs(167) <= (inputs(128)) and not (inputs(237));
    layer0_outputs(168) <= (inputs(118)) and not (inputs(14));
    layer0_outputs(169) <= not((inputs(237)) or (inputs(49)));
    layer0_outputs(170) <= not((inputs(130)) or (inputs(153)));
    layer0_outputs(171) <= inputs(34);
    layer0_outputs(172) <= (inputs(73)) xor (inputs(29));
    layer0_outputs(173) <= (inputs(47)) or (inputs(107));
    layer0_outputs(174) <= not(inputs(195));
    layer0_outputs(175) <= not((inputs(201)) or (inputs(78)));
    layer0_outputs(176) <= not(inputs(72)) or (inputs(179));
    layer0_outputs(177) <= '1';
    layer0_outputs(178) <= (inputs(159)) and not (inputs(14));
    layer0_outputs(179) <= inputs(51);
    layer0_outputs(180) <= not((inputs(241)) or (inputs(108)));
    layer0_outputs(181) <= (inputs(64)) or (inputs(205));
    layer0_outputs(182) <= not(inputs(135));
    layer0_outputs(183) <= not((inputs(31)) xor (inputs(38)));
    layer0_outputs(184) <= '0';
    layer0_outputs(185) <= inputs(68);
    layer0_outputs(186) <= (inputs(14)) and not (inputs(11));
    layer0_outputs(187) <= inputs(246);
    layer0_outputs(188) <= (inputs(107)) and not (inputs(233));
    layer0_outputs(189) <= not(inputs(39)) or (inputs(62));
    layer0_outputs(190) <= inputs(151);
    layer0_outputs(191) <= not(inputs(19));
    layer0_outputs(192) <= not((inputs(193)) and (inputs(111)));
    layer0_outputs(193) <= not((inputs(137)) or (inputs(67)));
    layer0_outputs(194) <= not(inputs(215)) or (inputs(195));
    layer0_outputs(195) <= not((inputs(105)) or (inputs(237)));
    layer0_outputs(196) <= not((inputs(177)) xor (inputs(19)));
    layer0_outputs(197) <= not(inputs(109));
    layer0_outputs(198) <= inputs(117);
    layer0_outputs(199) <= (inputs(138)) or (inputs(229));
    layer0_outputs(200) <= not((inputs(125)) and (inputs(112)));
    layer0_outputs(201) <= (inputs(250)) and (inputs(128));
    layer0_outputs(202) <= not(inputs(231)) or (inputs(191));
    layer0_outputs(203) <= not((inputs(177)) or (inputs(12)));
    layer0_outputs(204) <= (inputs(114)) and (inputs(249));
    layer0_outputs(205) <= '1';
    layer0_outputs(206) <= not(inputs(166)) or (inputs(75));
    layer0_outputs(207) <= '0';
    layer0_outputs(208) <= inputs(211);
    layer0_outputs(209) <= not(inputs(33)) or (inputs(127));
    layer0_outputs(210) <= (inputs(222)) xor (inputs(249));
    layer0_outputs(211) <= (inputs(23)) and not (inputs(252));
    layer0_outputs(212) <= (inputs(223)) and (inputs(238));
    layer0_outputs(213) <= not(inputs(42));
    layer0_outputs(214) <= (inputs(120)) and not (inputs(172));
    layer0_outputs(215) <= (inputs(10)) and not (inputs(44));
    layer0_outputs(216) <= not(inputs(232));
    layer0_outputs(217) <= (inputs(194)) and not (inputs(252));
    layer0_outputs(218) <= not(inputs(186)) or (inputs(100));
    layer0_outputs(219) <= not((inputs(126)) or (inputs(20)));
    layer0_outputs(220) <= not((inputs(125)) xor (inputs(11)));
    layer0_outputs(221) <= not((inputs(107)) or (inputs(128)));
    layer0_outputs(222) <= not((inputs(202)) xor (inputs(139)));
    layer0_outputs(223) <= not((inputs(41)) or (inputs(123)));
    layer0_outputs(224) <= inputs(187);
    layer0_outputs(225) <= (inputs(49)) or (inputs(0));
    layer0_outputs(226) <= inputs(107);
    layer0_outputs(227) <= not(inputs(182));
    layer0_outputs(228) <= (inputs(179)) and not (inputs(29));
    layer0_outputs(229) <= not((inputs(39)) xor (inputs(136)));
    layer0_outputs(230) <= (inputs(25)) and not (inputs(247));
    layer0_outputs(231) <= (inputs(20)) and not (inputs(237));
    layer0_outputs(232) <= not(inputs(106));
    layer0_outputs(233) <= not(inputs(145)) or (inputs(109));
    layer0_outputs(234) <= not((inputs(171)) xor (inputs(254)));
    layer0_outputs(235) <= (inputs(181)) and not (inputs(140));
    layer0_outputs(236) <= not((inputs(78)) xor (inputs(52)));
    layer0_outputs(237) <= not((inputs(121)) or (inputs(130)));
    layer0_outputs(238) <= not(inputs(248));
    layer0_outputs(239) <= inputs(252);
    layer0_outputs(240) <= inputs(116);
    layer0_outputs(241) <= (inputs(25)) or (inputs(69));
    layer0_outputs(242) <= (inputs(169)) and not (inputs(190));
    layer0_outputs(243) <= (inputs(85)) or (inputs(34));
    layer0_outputs(244) <= not(inputs(70)) or (inputs(158));
    layer0_outputs(245) <= not(inputs(145));
    layer0_outputs(246) <= not((inputs(14)) xor (inputs(188)));
    layer0_outputs(247) <= inputs(89);
    layer0_outputs(248) <= inputs(132);
    layer0_outputs(249) <= not(inputs(94)) or (inputs(14));
    layer0_outputs(250) <= not(inputs(40));
    layer0_outputs(251) <= (inputs(2)) xor (inputs(211));
    layer0_outputs(252) <= not((inputs(14)) xor (inputs(165)));
    layer0_outputs(253) <= not(inputs(228)) or (inputs(63));
    layer0_outputs(254) <= not((inputs(217)) xor (inputs(1)));
    layer0_outputs(255) <= not((inputs(48)) or (inputs(108)));
    layer0_outputs(256) <= not(inputs(120)) or (inputs(204));
    layer0_outputs(257) <= (inputs(188)) xor (inputs(233));
    layer0_outputs(258) <= not(inputs(131));
    layer0_outputs(259) <= not(inputs(157)) or (inputs(240));
    layer0_outputs(260) <= (inputs(140)) or (inputs(96));
    layer0_outputs(261) <= not(inputs(253));
    layer0_outputs(262) <= not(inputs(41));
    layer0_outputs(263) <= not((inputs(251)) or (inputs(0)));
    layer0_outputs(264) <= inputs(117);
    layer0_outputs(265) <= '0';
    layer0_outputs(266) <= inputs(204);
    layer0_outputs(267) <= (inputs(209)) and not (inputs(69));
    layer0_outputs(268) <= not(inputs(115)) or (inputs(178));
    layer0_outputs(269) <= (inputs(63)) and not (inputs(43));
    layer0_outputs(270) <= (inputs(202)) and not (inputs(247));
    layer0_outputs(271) <= (inputs(60)) or (inputs(110));
    layer0_outputs(272) <= not((inputs(122)) or (inputs(229)));
    layer0_outputs(273) <= (inputs(236)) or (inputs(4));
    layer0_outputs(274) <= not((inputs(186)) and (inputs(104)));
    layer0_outputs(275) <= (inputs(205)) or (inputs(61));
    layer0_outputs(276) <= not(inputs(85));
    layer0_outputs(277) <= inputs(134);
    layer0_outputs(278) <= inputs(54);
    layer0_outputs(279) <= not((inputs(255)) or (inputs(59)));
    layer0_outputs(280) <= (inputs(149)) or (inputs(246));
    layer0_outputs(281) <= '0';
    layer0_outputs(282) <= (inputs(75)) or (inputs(206));
    layer0_outputs(283) <= inputs(223);
    layer0_outputs(284) <= (inputs(17)) or (inputs(199));
    layer0_outputs(285) <= not((inputs(254)) or (inputs(92)));
    layer0_outputs(286) <= not(inputs(104));
    layer0_outputs(287) <= (inputs(141)) xor (inputs(90));
    layer0_outputs(288) <= inputs(166);
    layer0_outputs(289) <= (inputs(242)) or (inputs(136));
    layer0_outputs(290) <= (inputs(64)) or (inputs(191));
    layer0_outputs(291) <= not((inputs(87)) xor (inputs(169)));
    layer0_outputs(292) <= (inputs(87)) and not (inputs(245));
    layer0_outputs(293) <= inputs(120);
    layer0_outputs(294) <= not((inputs(142)) and (inputs(163)));
    layer0_outputs(295) <= (inputs(249)) and (inputs(148));
    layer0_outputs(296) <= inputs(198);
    layer0_outputs(297) <= inputs(180);
    layer0_outputs(298) <= inputs(239);
    layer0_outputs(299) <= (inputs(237)) xor (inputs(61));
    layer0_outputs(300) <= not((inputs(87)) or (inputs(136)));
    layer0_outputs(301) <= (inputs(212)) or (inputs(57));
    layer0_outputs(302) <= not((inputs(211)) and (inputs(33)));
    layer0_outputs(303) <= (inputs(90)) and not (inputs(43));
    layer0_outputs(304) <= not(inputs(154)) or (inputs(32));
    layer0_outputs(305) <= (inputs(235)) and not (inputs(240));
    layer0_outputs(306) <= (inputs(167)) and not (inputs(76));
    layer0_outputs(307) <= (inputs(196)) and not (inputs(17));
    layer0_outputs(308) <= not((inputs(50)) or (inputs(152)));
    layer0_outputs(309) <= (inputs(44)) xor (inputs(12));
    layer0_outputs(310) <= (inputs(94)) or (inputs(11));
    layer0_outputs(311) <= (inputs(203)) and not (inputs(224));
    layer0_outputs(312) <= (inputs(91)) or (inputs(149));
    layer0_outputs(313) <= (inputs(40)) or (inputs(137));
    layer0_outputs(314) <= (inputs(236)) or (inputs(19));
    layer0_outputs(315) <= not((inputs(244)) or (inputs(164)));
    layer0_outputs(316) <= (inputs(123)) and not (inputs(81));
    layer0_outputs(317) <= (inputs(22)) and not (inputs(46));
    layer0_outputs(318) <= (inputs(120)) and not (inputs(93));
    layer0_outputs(319) <= (inputs(133)) and not (inputs(187));
    layer0_outputs(320) <= (inputs(85)) and not (inputs(12));
    layer0_outputs(321) <= inputs(115);
    layer0_outputs(322) <= inputs(204);
    layer0_outputs(323) <= '0';
    layer0_outputs(324) <= inputs(49);
    layer0_outputs(325) <= (inputs(28)) or (inputs(42));
    layer0_outputs(326) <= not(inputs(79));
    layer0_outputs(327) <= not(inputs(70)) or (inputs(220));
    layer0_outputs(328) <= (inputs(125)) and (inputs(157));
    layer0_outputs(329) <= (inputs(11)) xor (inputs(38));
    layer0_outputs(330) <= inputs(140);
    layer0_outputs(331) <= (inputs(29)) or (inputs(152));
    layer0_outputs(332) <= not(inputs(218));
    layer0_outputs(333) <= inputs(175);
    layer0_outputs(334) <= not((inputs(26)) or (inputs(134)));
    layer0_outputs(335) <= inputs(151);
    layer0_outputs(336) <= '0';
    layer0_outputs(337) <= not(inputs(182)) or (inputs(65));
    layer0_outputs(338) <= (inputs(213)) or (inputs(82));
    layer0_outputs(339) <= not(inputs(88));
    layer0_outputs(340) <= '1';
    layer0_outputs(341) <= (inputs(23)) and not (inputs(110));
    layer0_outputs(342) <= not((inputs(4)) or (inputs(76)));
    layer0_outputs(343) <= not(inputs(158));
    layer0_outputs(344) <= (inputs(215)) and not (inputs(195));
    layer0_outputs(345) <= (inputs(159)) or (inputs(191));
    layer0_outputs(346) <= not((inputs(174)) xor (inputs(97)));
    layer0_outputs(347) <= not(inputs(114));
    layer0_outputs(348) <= (inputs(211)) and not (inputs(111));
    layer0_outputs(349) <= (inputs(118)) or (inputs(4));
    layer0_outputs(350) <= '1';
    layer0_outputs(351) <= (inputs(94)) and (inputs(4));
    layer0_outputs(352) <= not((inputs(170)) or (inputs(116)));
    layer0_outputs(353) <= not((inputs(193)) and (inputs(14)));
    layer0_outputs(354) <= not((inputs(58)) xor (inputs(63)));
    layer0_outputs(355) <= not(inputs(63));
    layer0_outputs(356) <= not((inputs(10)) or (inputs(97)));
    layer0_outputs(357) <= not((inputs(54)) or (inputs(99)));
    layer0_outputs(358) <= not(inputs(167)) or (inputs(178));
    layer0_outputs(359) <= inputs(52);
    layer0_outputs(360) <= (inputs(211)) or (inputs(7));
    layer0_outputs(361) <= (inputs(151)) or (inputs(125));
    layer0_outputs(362) <= inputs(115);
    layer0_outputs(363) <= (inputs(107)) or (inputs(140));
    layer0_outputs(364) <= not((inputs(79)) or (inputs(54)));
    layer0_outputs(365) <= inputs(136);
    layer0_outputs(366) <= not(inputs(20)) or (inputs(21));
    layer0_outputs(367) <= not((inputs(198)) xor (inputs(162)));
    layer0_outputs(368) <= not(inputs(13));
    layer0_outputs(369) <= (inputs(186)) and not (inputs(110));
    layer0_outputs(370) <= not(inputs(167));
    layer0_outputs(371) <= not(inputs(203));
    layer0_outputs(372) <= (inputs(165)) or (inputs(196));
    layer0_outputs(373) <= (inputs(155)) and not (inputs(20));
    layer0_outputs(374) <= not((inputs(230)) or (inputs(62)));
    layer0_outputs(375) <= not(inputs(104));
    layer0_outputs(376) <= (inputs(168)) xor (inputs(81));
    layer0_outputs(377) <= inputs(76);
    layer0_outputs(378) <= not(inputs(133));
    layer0_outputs(379) <= (inputs(246)) or (inputs(180));
    layer0_outputs(380) <= (inputs(160)) xor (inputs(247));
    layer0_outputs(381) <= (inputs(73)) and not (inputs(16));
    layer0_outputs(382) <= '0';
    layer0_outputs(383) <= not(inputs(61));
    layer0_outputs(384) <= not(inputs(120));
    layer0_outputs(385) <= not((inputs(188)) xor (inputs(139)));
    layer0_outputs(386) <= not((inputs(42)) or (inputs(15)));
    layer0_outputs(387) <= (inputs(159)) and not (inputs(53));
    layer0_outputs(388) <= not((inputs(79)) xor (inputs(100)));
    layer0_outputs(389) <= not((inputs(31)) xor (inputs(152)));
    layer0_outputs(390) <= not((inputs(144)) or (inputs(197)));
    layer0_outputs(391) <= not(inputs(76));
    layer0_outputs(392) <= not((inputs(232)) or (inputs(231)));
    layer0_outputs(393) <= not((inputs(249)) xor (inputs(177)));
    layer0_outputs(394) <= (inputs(67)) xor (inputs(29));
    layer0_outputs(395) <= not((inputs(156)) or (inputs(250)));
    layer0_outputs(396) <= not((inputs(239)) and (inputs(221)));
    layer0_outputs(397) <= inputs(33);
    layer0_outputs(398) <= not(inputs(116));
    layer0_outputs(399) <= (inputs(68)) and not (inputs(142));
    layer0_outputs(400) <= (inputs(85)) or (inputs(97));
    layer0_outputs(401) <= inputs(169);
    layer0_outputs(402) <= not((inputs(227)) and (inputs(113)));
    layer0_outputs(403) <= not((inputs(29)) or (inputs(166)));
    layer0_outputs(404) <= (inputs(216)) or (inputs(206));
    layer0_outputs(405) <= not((inputs(31)) xor (inputs(167)));
    layer0_outputs(406) <= not((inputs(121)) or (inputs(81)));
    layer0_outputs(407) <= (inputs(39)) xor (inputs(2));
    layer0_outputs(408) <= (inputs(229)) and not (inputs(79));
    layer0_outputs(409) <= not(inputs(214));
    layer0_outputs(410) <= not(inputs(165));
    layer0_outputs(411) <= not((inputs(160)) or (inputs(162)));
    layer0_outputs(412) <= (inputs(98)) and not (inputs(189));
    layer0_outputs(413) <= not(inputs(60)) or (inputs(255));
    layer0_outputs(414) <= not(inputs(10));
    layer0_outputs(415) <= inputs(13);
    layer0_outputs(416) <= not(inputs(55)) or (inputs(114));
    layer0_outputs(417) <= not((inputs(35)) xor (inputs(126)));
    layer0_outputs(418) <= not(inputs(144)) or (inputs(217));
    layer0_outputs(419) <= not((inputs(140)) or (inputs(186)));
    layer0_outputs(420) <= not(inputs(185));
    layer0_outputs(421) <= '0';
    layer0_outputs(422) <= not(inputs(84)) or (inputs(94));
    layer0_outputs(423) <= (inputs(93)) and not (inputs(206));
    layer0_outputs(424) <= inputs(47);
    layer0_outputs(425) <= not(inputs(106)) or (inputs(30));
    layer0_outputs(426) <= (inputs(196)) xor (inputs(6));
    layer0_outputs(427) <= (inputs(251)) and (inputs(157));
    layer0_outputs(428) <= inputs(111);
    layer0_outputs(429) <= (inputs(251)) xor (inputs(175));
    layer0_outputs(430) <= inputs(141);
    layer0_outputs(431) <= inputs(138);
    layer0_outputs(432) <= (inputs(106)) and not (inputs(163));
    layer0_outputs(433) <= inputs(119);
    layer0_outputs(434) <= not((inputs(57)) or (inputs(205)));
    layer0_outputs(435) <= (inputs(76)) and not (inputs(10));
    layer0_outputs(436) <= not(inputs(163)) or (inputs(11));
    layer0_outputs(437) <= not(inputs(59));
    layer0_outputs(438) <= not((inputs(4)) xor (inputs(116)));
    layer0_outputs(439) <= inputs(116);
    layer0_outputs(440) <= not(inputs(27)) or (inputs(112));
    layer0_outputs(441) <= (inputs(209)) and (inputs(65));
    layer0_outputs(442) <= (inputs(86)) and not (inputs(111));
    layer0_outputs(443) <= not(inputs(142)) or (inputs(112));
    layer0_outputs(444) <= (inputs(187)) or (inputs(43));
    layer0_outputs(445) <= not((inputs(227)) or (inputs(212)));
    layer0_outputs(446) <= (inputs(145)) and (inputs(113));
    layer0_outputs(447) <= (inputs(152)) or (inputs(244));
    layer0_outputs(448) <= inputs(27);
    layer0_outputs(449) <= (inputs(208)) or (inputs(203));
    layer0_outputs(450) <= not((inputs(22)) xor (inputs(212)));
    layer0_outputs(451) <= not((inputs(228)) or (inputs(156)));
    layer0_outputs(452) <= not(inputs(181));
    layer0_outputs(453) <= inputs(181);
    layer0_outputs(454) <= not((inputs(7)) or (inputs(86)));
    layer0_outputs(455) <= not((inputs(255)) xor (inputs(131)));
    layer0_outputs(456) <= (inputs(165)) xor (inputs(81));
    layer0_outputs(457) <= (inputs(211)) or (inputs(133));
    layer0_outputs(458) <= not((inputs(3)) and (inputs(128)));
    layer0_outputs(459) <= (inputs(148)) and not (inputs(244));
    layer0_outputs(460) <= not(inputs(179)) or (inputs(118));
    layer0_outputs(461) <= (inputs(104)) or (inputs(196));
    layer0_outputs(462) <= not((inputs(165)) or (inputs(106)));
    layer0_outputs(463) <= inputs(120);
    layer0_outputs(464) <= not((inputs(19)) or (inputs(101)));
    layer0_outputs(465) <= inputs(94);
    layer0_outputs(466) <= (inputs(54)) or (inputs(79));
    layer0_outputs(467) <= (inputs(149)) and not (inputs(1));
    layer0_outputs(468) <= not((inputs(12)) xor (inputs(142)));
    layer0_outputs(469) <= not((inputs(110)) xor (inputs(104)));
    layer0_outputs(470) <= (inputs(104)) and not (inputs(238));
    layer0_outputs(471) <= (inputs(174)) xor (inputs(250));
    layer0_outputs(472) <= not(inputs(54));
    layer0_outputs(473) <= not(inputs(46)) or (inputs(6));
    layer0_outputs(474) <= not(inputs(67)) or (inputs(236));
    layer0_outputs(475) <= inputs(200);
    layer0_outputs(476) <= (inputs(86)) xor (inputs(160));
    layer0_outputs(477) <= not((inputs(110)) or (inputs(113)));
    layer0_outputs(478) <= not(inputs(227)) or (inputs(146));
    layer0_outputs(479) <= (inputs(179)) xor (inputs(198));
    layer0_outputs(480) <= not(inputs(99)) or (inputs(249));
    layer0_outputs(481) <= inputs(19);
    layer0_outputs(482) <= inputs(109);
    layer0_outputs(483) <= not((inputs(160)) and (inputs(145)));
    layer0_outputs(484) <= not((inputs(10)) xor (inputs(100)));
    layer0_outputs(485) <= not(inputs(241));
    layer0_outputs(486) <= (inputs(96)) or (inputs(167));
    layer0_outputs(487) <= not(inputs(22)) or (inputs(254));
    layer0_outputs(488) <= not(inputs(112));
    layer0_outputs(489) <= not(inputs(63));
    layer0_outputs(490) <= (inputs(27)) or (inputs(166));
    layer0_outputs(491) <= inputs(126);
    layer0_outputs(492) <= not(inputs(119)) or (inputs(144));
    layer0_outputs(493) <= not(inputs(93)) or (inputs(35));
    layer0_outputs(494) <= not(inputs(50)) or (inputs(147));
    layer0_outputs(495) <= (inputs(163)) xor (inputs(136));
    layer0_outputs(496) <= not(inputs(252));
    layer0_outputs(497) <= not((inputs(130)) and (inputs(112)));
    layer0_outputs(498) <= '1';
    layer0_outputs(499) <= inputs(108);
    layer0_outputs(500) <= not((inputs(114)) or (inputs(220)));
    layer0_outputs(501) <= not(inputs(22));
    layer0_outputs(502) <= not(inputs(214)) or (inputs(44));
    layer0_outputs(503) <= inputs(163);
    layer0_outputs(504) <= not((inputs(211)) or (inputs(106)));
    layer0_outputs(505) <= not((inputs(212)) or (inputs(160)));
    layer0_outputs(506) <= not((inputs(229)) xor (inputs(211)));
    layer0_outputs(507) <= not((inputs(146)) or (inputs(230)));
    layer0_outputs(508) <= not(inputs(152)) or (inputs(121));
    layer0_outputs(509) <= not((inputs(218)) or (inputs(40)));
    layer0_outputs(510) <= (inputs(161)) xor (inputs(231));
    layer0_outputs(511) <= not(inputs(165));
    layer0_outputs(512) <= not(inputs(40));
    layer0_outputs(513) <= not(inputs(253)) or (inputs(163));
    layer0_outputs(514) <= (inputs(167)) and not (inputs(81));
    layer0_outputs(515) <= (inputs(179)) or (inputs(7));
    layer0_outputs(516) <= (inputs(47)) or (inputs(117));
    layer0_outputs(517) <= not((inputs(149)) or (inputs(65)));
    layer0_outputs(518) <= inputs(152);
    layer0_outputs(519) <= inputs(59);
    layer0_outputs(520) <= not((inputs(116)) xor (inputs(117)));
    layer0_outputs(521) <= not(inputs(10)) or (inputs(176));
    layer0_outputs(522) <= inputs(21);
    layer0_outputs(523) <= (inputs(114)) or (inputs(127));
    layer0_outputs(524) <= not((inputs(22)) or (inputs(121)));
    layer0_outputs(525) <= inputs(180);
    layer0_outputs(526) <= (inputs(200)) and not (inputs(182));
    layer0_outputs(527) <= not(inputs(19));
    layer0_outputs(528) <= (inputs(71)) xor (inputs(65));
    layer0_outputs(529) <= not((inputs(180)) or (inputs(93)));
    layer0_outputs(530) <= not((inputs(98)) or (inputs(198)));
    layer0_outputs(531) <= (inputs(61)) xor (inputs(65));
    layer0_outputs(532) <= not(inputs(126)) or (inputs(206));
    layer0_outputs(533) <= (inputs(164)) or (inputs(35));
    layer0_outputs(534) <= not((inputs(242)) xor (inputs(115)));
    layer0_outputs(535) <= not((inputs(46)) xor (inputs(86)));
    layer0_outputs(536) <= not(inputs(130)) or (inputs(115));
    layer0_outputs(537) <= (inputs(155)) xor (inputs(171));
    layer0_outputs(538) <= not((inputs(122)) or (inputs(133)));
    layer0_outputs(539) <= not((inputs(176)) xor (inputs(234)));
    layer0_outputs(540) <= not(inputs(184)) or (inputs(9));
    layer0_outputs(541) <= not(inputs(119));
    layer0_outputs(542) <= inputs(229);
    layer0_outputs(543) <= not(inputs(117)) or (inputs(155));
    layer0_outputs(544) <= not(inputs(88));
    layer0_outputs(545) <= (inputs(201)) and (inputs(85));
    layer0_outputs(546) <= not((inputs(196)) or (inputs(17)));
    layer0_outputs(547) <= (inputs(108)) xor (inputs(142));
    layer0_outputs(548) <= (inputs(214)) or (inputs(52));
    layer0_outputs(549) <= (inputs(183)) and (inputs(83));
    layer0_outputs(550) <= not(inputs(0)) or (inputs(226));
    layer0_outputs(551) <= not(inputs(150));
    layer0_outputs(552) <= not((inputs(141)) and (inputs(141)));
    layer0_outputs(553) <= (inputs(11)) xor (inputs(105));
    layer0_outputs(554) <= not(inputs(125));
    layer0_outputs(555) <= (inputs(182)) or (inputs(149));
    layer0_outputs(556) <= not(inputs(80)) or (inputs(227));
    layer0_outputs(557) <= not((inputs(227)) and (inputs(245)));
    layer0_outputs(558) <= not(inputs(132));
    layer0_outputs(559) <= not((inputs(69)) xor (inputs(160)));
    layer0_outputs(560) <= '1';
    layer0_outputs(561) <= (inputs(119)) and not (inputs(147));
    layer0_outputs(562) <= not((inputs(106)) or (inputs(219)));
    layer0_outputs(563) <= not(inputs(62));
    layer0_outputs(564) <= (inputs(150)) and not (inputs(144));
    layer0_outputs(565) <= not(inputs(97));
    layer0_outputs(566) <= not(inputs(189));
    layer0_outputs(567) <= not((inputs(148)) or (inputs(91)));
    layer0_outputs(568) <= inputs(53);
    layer0_outputs(569) <= (inputs(57)) or (inputs(188));
    layer0_outputs(570) <= not((inputs(206)) or (inputs(35)));
    layer0_outputs(571) <= not((inputs(254)) and (inputs(126)));
    layer0_outputs(572) <= (inputs(21)) or (inputs(72));
    layer0_outputs(573) <= not(inputs(124)) or (inputs(40));
    layer0_outputs(574) <= not((inputs(232)) xor (inputs(174)));
    layer0_outputs(575) <= (inputs(130)) or (inputs(89));
    layer0_outputs(576) <= not((inputs(226)) or (inputs(227)));
    layer0_outputs(577) <= (inputs(194)) and (inputs(111));
    layer0_outputs(578) <= not((inputs(39)) xor (inputs(225)));
    layer0_outputs(579) <= (inputs(140)) and not (inputs(216));
    layer0_outputs(580) <= not(inputs(136)) or (inputs(234));
    layer0_outputs(581) <= (inputs(118)) and not (inputs(100));
    layer0_outputs(582) <= not((inputs(105)) xor (inputs(112)));
    layer0_outputs(583) <= not((inputs(224)) and (inputs(94)));
    layer0_outputs(584) <= not(inputs(148)) or (inputs(160));
    layer0_outputs(585) <= (inputs(121)) and not (inputs(119));
    layer0_outputs(586) <= (inputs(113)) xor (inputs(165));
    layer0_outputs(587) <= not(inputs(134)) or (inputs(246));
    layer0_outputs(588) <= not((inputs(250)) or (inputs(224)));
    layer0_outputs(589) <= not((inputs(84)) xor (inputs(99)));
    layer0_outputs(590) <= inputs(53);
    layer0_outputs(591) <= not((inputs(167)) xor (inputs(89)));
    layer0_outputs(592) <= not((inputs(149)) or (inputs(109)));
    layer0_outputs(593) <= not(inputs(102)) or (inputs(166));
    layer0_outputs(594) <= not(inputs(221));
    layer0_outputs(595) <= not(inputs(152));
    layer0_outputs(596) <= (inputs(224)) and not (inputs(57));
    layer0_outputs(597) <= inputs(107);
    layer0_outputs(598) <= (inputs(196)) xor (inputs(19));
    layer0_outputs(599) <= not((inputs(193)) xor (inputs(0)));
    layer0_outputs(600) <= inputs(95);
    layer0_outputs(601) <= (inputs(52)) and not (inputs(45));
    layer0_outputs(602) <= not((inputs(124)) or (inputs(109)));
    layer0_outputs(603) <= not((inputs(49)) xor (inputs(142)));
    layer0_outputs(604) <= not((inputs(22)) or (inputs(186)));
    layer0_outputs(605) <= inputs(212);
    layer0_outputs(606) <= not((inputs(208)) or (inputs(60)));
    layer0_outputs(607) <= not((inputs(74)) or (inputs(41)));
    layer0_outputs(608) <= (inputs(184)) and not (inputs(92));
    layer0_outputs(609) <= (inputs(173)) and not (inputs(17));
    layer0_outputs(610) <= not(inputs(118));
    layer0_outputs(611) <= not(inputs(68)) or (inputs(45));
    layer0_outputs(612) <= (inputs(253)) and (inputs(86));
    layer0_outputs(613) <= not(inputs(250)) or (inputs(161));
    layer0_outputs(614) <= not((inputs(10)) xor (inputs(247)));
    layer0_outputs(615) <= (inputs(71)) xor (inputs(59));
    layer0_outputs(616) <= not((inputs(67)) or (inputs(45)));
    layer0_outputs(617) <= not((inputs(81)) xor (inputs(47)));
    layer0_outputs(618) <= (inputs(168)) and not (inputs(112));
    layer0_outputs(619) <= inputs(175);
    layer0_outputs(620) <= not(inputs(175)) or (inputs(11));
    layer0_outputs(621) <= (inputs(40)) and not (inputs(229));
    layer0_outputs(622) <= (inputs(97)) and not (inputs(1));
    layer0_outputs(623) <= not(inputs(174)) or (inputs(31));
    layer0_outputs(624) <= not(inputs(75)) or (inputs(240));
    layer0_outputs(625) <= inputs(107);
    layer0_outputs(626) <= not((inputs(116)) or (inputs(16)));
    layer0_outputs(627) <= inputs(94);
    layer0_outputs(628) <= (inputs(158)) or (inputs(155));
    layer0_outputs(629) <= (inputs(110)) or (inputs(207));
    layer0_outputs(630) <= not(inputs(234)) or (inputs(161));
    layer0_outputs(631) <= (inputs(0)) and (inputs(170));
    layer0_outputs(632) <= (inputs(49)) or (inputs(247));
    layer0_outputs(633) <= (inputs(248)) and not (inputs(142));
    layer0_outputs(634) <= (inputs(94)) xor (inputs(232));
    layer0_outputs(635) <= (inputs(90)) and (inputs(250));
    layer0_outputs(636) <= inputs(121);
    layer0_outputs(637) <= (inputs(195)) and not (inputs(250));
    layer0_outputs(638) <= not(inputs(189));
    layer0_outputs(639) <= not((inputs(9)) or (inputs(226)));
    layer0_outputs(640) <= not((inputs(121)) xor (inputs(98)));
    layer0_outputs(641) <= not((inputs(194)) or (inputs(195)));
    layer0_outputs(642) <= not(inputs(106));
    layer0_outputs(643) <= not((inputs(68)) or (inputs(152)));
    layer0_outputs(644) <= (inputs(203)) xor (inputs(186));
    layer0_outputs(645) <= inputs(89);
    layer0_outputs(646) <= not(inputs(86));
    layer0_outputs(647) <= (inputs(34)) xor (inputs(182));
    layer0_outputs(648) <= not((inputs(224)) or (inputs(36)));
    layer0_outputs(649) <= inputs(233);
    layer0_outputs(650) <= (inputs(223)) and not (inputs(156));
    layer0_outputs(651) <= (inputs(116)) and not (inputs(192));
    layer0_outputs(652) <= (inputs(108)) and not (inputs(53));
    layer0_outputs(653) <= not(inputs(216)) or (inputs(144));
    layer0_outputs(654) <= not(inputs(58));
    layer0_outputs(655) <= not((inputs(153)) xor (inputs(240)));
    layer0_outputs(656) <= (inputs(193)) or (inputs(237));
    layer0_outputs(657) <= not(inputs(247)) or (inputs(193));
    layer0_outputs(658) <= (inputs(202)) xor (inputs(154));
    layer0_outputs(659) <= (inputs(150)) and not (inputs(156));
    layer0_outputs(660) <= not(inputs(52)) or (inputs(75));
    layer0_outputs(661) <= (inputs(45)) xor (inputs(205));
    layer0_outputs(662) <= (inputs(121)) and not (inputs(228));
    layer0_outputs(663) <= not((inputs(31)) and (inputs(190)));
    layer0_outputs(664) <= (inputs(71)) or (inputs(13));
    layer0_outputs(665) <= not(inputs(71)) or (inputs(121));
    layer0_outputs(666) <= (inputs(210)) and not (inputs(227));
    layer0_outputs(667) <= inputs(20);
    layer0_outputs(668) <= (inputs(137)) and not (inputs(62));
    layer0_outputs(669) <= inputs(38);
    layer0_outputs(670) <= (inputs(59)) or (inputs(120));
    layer0_outputs(671) <= not((inputs(230)) or (inputs(25)));
    layer0_outputs(672) <= not((inputs(162)) xor (inputs(9)));
    layer0_outputs(673) <= not(inputs(86)) or (inputs(228));
    layer0_outputs(674) <= (inputs(81)) or (inputs(96));
    layer0_outputs(675) <= inputs(137);
    layer0_outputs(676) <= not(inputs(143));
    layer0_outputs(677) <= not(inputs(248));
    layer0_outputs(678) <= (inputs(69)) or (inputs(98));
    layer0_outputs(679) <= not((inputs(243)) xor (inputs(122)));
    layer0_outputs(680) <= inputs(181);
    layer0_outputs(681) <= inputs(111);
    layer0_outputs(682) <= (inputs(253)) xor (inputs(92));
    layer0_outputs(683) <= not((inputs(175)) xor (inputs(248)));
    layer0_outputs(684) <= not(inputs(241));
    layer0_outputs(685) <= not(inputs(87)) or (inputs(15));
    layer0_outputs(686) <= (inputs(129)) and not (inputs(177));
    layer0_outputs(687) <= not((inputs(241)) or (inputs(126)));
    layer0_outputs(688) <= (inputs(45)) and (inputs(79));
    layer0_outputs(689) <= '0';
    layer0_outputs(690) <= not((inputs(44)) or (inputs(32)));
    layer0_outputs(691) <= (inputs(93)) xor (inputs(173));
    layer0_outputs(692) <= not(inputs(123)) or (inputs(226));
    layer0_outputs(693) <= (inputs(123)) and (inputs(15));
    layer0_outputs(694) <= (inputs(26)) xor (inputs(44));
    layer0_outputs(695) <= inputs(1);
    layer0_outputs(696) <= not((inputs(129)) or (inputs(99)));
    layer0_outputs(697) <= inputs(46);
    layer0_outputs(698) <= (inputs(2)) and (inputs(41));
    layer0_outputs(699) <= (inputs(127)) and (inputs(248));
    layer0_outputs(700) <= not(inputs(216));
    layer0_outputs(701) <= not(inputs(182));
    layer0_outputs(702) <= not((inputs(125)) or (inputs(39)));
    layer0_outputs(703) <= not(inputs(81));
    layer0_outputs(704) <= not(inputs(144));
    layer0_outputs(705) <= (inputs(219)) or (inputs(137));
    layer0_outputs(706) <= inputs(13);
    layer0_outputs(707) <= (inputs(52)) or (inputs(204));
    layer0_outputs(708) <= not((inputs(219)) or (inputs(236)));
    layer0_outputs(709) <= (inputs(126)) and not (inputs(190));
    layer0_outputs(710) <= inputs(172);
    layer0_outputs(711) <= not((inputs(12)) xor (inputs(106)));
    layer0_outputs(712) <= (inputs(188)) or (inputs(220));
    layer0_outputs(713) <= (inputs(210)) xor (inputs(171));
    layer0_outputs(714) <= not(inputs(195));
    layer0_outputs(715) <= (inputs(81)) and (inputs(68));
    layer0_outputs(716) <= not((inputs(97)) and (inputs(26)));
    layer0_outputs(717) <= (inputs(53)) and not (inputs(115));
    layer0_outputs(718) <= (inputs(177)) xor (inputs(83));
    layer0_outputs(719) <= not((inputs(102)) xor (inputs(70)));
    layer0_outputs(720) <= inputs(101);
    layer0_outputs(721) <= inputs(27);
    layer0_outputs(722) <= not((inputs(208)) or (inputs(133)));
    layer0_outputs(723) <= (inputs(123)) and not (inputs(204));
    layer0_outputs(724) <= not((inputs(24)) or (inputs(78)));
    layer0_outputs(725) <= (inputs(210)) and not (inputs(209));
    layer0_outputs(726) <= not((inputs(39)) xor (inputs(216)));
    layer0_outputs(727) <= (inputs(23)) xor (inputs(134));
    layer0_outputs(728) <= not((inputs(220)) or (inputs(241)));
    layer0_outputs(729) <= (inputs(176)) or (inputs(55));
    layer0_outputs(730) <= inputs(148);
    layer0_outputs(731) <= not((inputs(39)) and (inputs(29)));
    layer0_outputs(732) <= (inputs(197)) xor (inputs(67));
    layer0_outputs(733) <= not((inputs(44)) or (inputs(140)));
    layer0_outputs(734) <= (inputs(244)) or (inputs(100));
    layer0_outputs(735) <= (inputs(37)) and not (inputs(212));
    layer0_outputs(736) <= '0';
    layer0_outputs(737) <= inputs(102);
    layer0_outputs(738) <= (inputs(218)) xor (inputs(131));
    layer0_outputs(739) <= (inputs(174)) xor (inputs(179));
    layer0_outputs(740) <= not((inputs(210)) and (inputs(7)));
    layer0_outputs(741) <= not(inputs(129));
    layer0_outputs(742) <= (inputs(42)) xor (inputs(89));
    layer0_outputs(743) <= '1';
    layer0_outputs(744) <= not((inputs(164)) or (inputs(172)));
    layer0_outputs(745) <= not((inputs(219)) xor (inputs(149)));
    layer0_outputs(746) <= inputs(131);
    layer0_outputs(747) <= (inputs(47)) and not (inputs(161));
    layer0_outputs(748) <= not(inputs(135)) or (inputs(4));
    layer0_outputs(749) <= (inputs(17)) and not (inputs(74));
    layer0_outputs(750) <= '0';
    layer0_outputs(751) <= '0';
    layer0_outputs(752) <= not(inputs(198)) or (inputs(144));
    layer0_outputs(753) <= inputs(90);
    layer0_outputs(754) <= inputs(35);
    layer0_outputs(755) <= not(inputs(132)) or (inputs(23));
    layer0_outputs(756) <= inputs(157);
    layer0_outputs(757) <= not((inputs(55)) or (inputs(94)));
    layer0_outputs(758) <= not((inputs(125)) xor (inputs(172)));
    layer0_outputs(759) <= not((inputs(187)) or (inputs(7)));
    layer0_outputs(760) <= not((inputs(41)) or (inputs(195)));
    layer0_outputs(761) <= (inputs(154)) and not (inputs(198));
    layer0_outputs(762) <= not((inputs(172)) xor (inputs(227)));
    layer0_outputs(763) <= not((inputs(104)) xor (inputs(20)));
    layer0_outputs(764) <= not((inputs(211)) xor (inputs(155)));
    layer0_outputs(765) <= inputs(140);
    layer0_outputs(766) <= not(inputs(35));
    layer0_outputs(767) <= not((inputs(67)) xor (inputs(185)));
    layer0_outputs(768) <= inputs(208);
    layer0_outputs(769) <= not((inputs(171)) or (inputs(51)));
    layer0_outputs(770) <= not((inputs(34)) or (inputs(197)));
    layer0_outputs(771) <= inputs(162);
    layer0_outputs(772) <= (inputs(214)) and not (inputs(28));
    layer0_outputs(773) <= inputs(85);
    layer0_outputs(774) <= not(inputs(232)) or (inputs(110));
    layer0_outputs(775) <= (inputs(182)) and not (inputs(7));
    layer0_outputs(776) <= (inputs(234)) xor (inputs(104));
    layer0_outputs(777) <= (inputs(221)) and (inputs(139));
    layer0_outputs(778) <= (inputs(167)) and (inputs(187));
    layer0_outputs(779) <= (inputs(127)) xor (inputs(152));
    layer0_outputs(780) <= inputs(135);
    layer0_outputs(781) <= inputs(59);
    layer0_outputs(782) <= (inputs(200)) and not (inputs(224));
    layer0_outputs(783) <= not(inputs(219));
    layer0_outputs(784) <= not((inputs(209)) or (inputs(227)));
    layer0_outputs(785) <= inputs(2);
    layer0_outputs(786) <= (inputs(97)) or (inputs(103));
    layer0_outputs(787) <= (inputs(205)) and not (inputs(8));
    layer0_outputs(788) <= inputs(20);
    layer0_outputs(789) <= not(inputs(235));
    layer0_outputs(790) <= (inputs(155)) xor (inputs(193));
    layer0_outputs(791) <= not(inputs(123));
    layer0_outputs(792) <= not(inputs(88));
    layer0_outputs(793) <= (inputs(196)) or (inputs(84));
    layer0_outputs(794) <= (inputs(46)) or (inputs(180));
    layer0_outputs(795) <= (inputs(170)) and (inputs(136));
    layer0_outputs(796) <= not((inputs(22)) xor (inputs(82)));
    layer0_outputs(797) <= (inputs(179)) and not (inputs(233));
    layer0_outputs(798) <= not(inputs(247)) or (inputs(173));
    layer0_outputs(799) <= (inputs(135)) and not (inputs(34));
    layer0_outputs(800) <= (inputs(73)) or (inputs(180));
    layer0_outputs(801) <= not(inputs(249)) or (inputs(255));
    layer0_outputs(802) <= (inputs(90)) and not (inputs(254));
    layer0_outputs(803) <= not(inputs(234)) or (inputs(140));
    layer0_outputs(804) <= (inputs(95)) xor (inputs(29));
    layer0_outputs(805) <= not((inputs(159)) xor (inputs(7)));
    layer0_outputs(806) <= (inputs(13)) or (inputs(248));
    layer0_outputs(807) <= (inputs(129)) and not (inputs(201));
    layer0_outputs(808) <= inputs(61);
    layer0_outputs(809) <= (inputs(159)) and (inputs(64));
    layer0_outputs(810) <= not(inputs(55)) or (inputs(205));
    layer0_outputs(811) <= inputs(193);
    layer0_outputs(812) <= not(inputs(197)) or (inputs(28));
    layer0_outputs(813) <= not(inputs(107));
    layer0_outputs(814) <= not(inputs(132));
    layer0_outputs(815) <= not((inputs(196)) or (inputs(92)));
    layer0_outputs(816) <= not((inputs(137)) or (inputs(130)));
    layer0_outputs(817) <= not(inputs(246));
    layer0_outputs(818) <= '0';
    layer0_outputs(819) <= (inputs(166)) or (inputs(29));
    layer0_outputs(820) <= (inputs(177)) or (inputs(73));
    layer0_outputs(821) <= not(inputs(18)) or (inputs(163));
    layer0_outputs(822) <= (inputs(152)) or (inputs(98));
    layer0_outputs(823) <= (inputs(105)) and (inputs(4));
    layer0_outputs(824) <= not(inputs(116));
    layer0_outputs(825) <= not(inputs(188)) or (inputs(7));
    layer0_outputs(826) <= (inputs(204)) or (inputs(38));
    layer0_outputs(827) <= inputs(109);
    layer0_outputs(828) <= '0';
    layer0_outputs(829) <= not((inputs(60)) or (inputs(77)));
    layer0_outputs(830) <= not((inputs(54)) xor (inputs(196)));
    layer0_outputs(831) <= not((inputs(65)) or (inputs(53)));
    layer0_outputs(832) <= not(inputs(197)) or (inputs(130));
    layer0_outputs(833) <= (inputs(244)) and not (inputs(110));
    layer0_outputs(834) <= not((inputs(95)) xor (inputs(87)));
    layer0_outputs(835) <= (inputs(249)) and not (inputs(47));
    layer0_outputs(836) <= not((inputs(22)) and (inputs(14)));
    layer0_outputs(837) <= inputs(133);
    layer0_outputs(838) <= inputs(34);
    layer0_outputs(839) <= (inputs(201)) or (inputs(187));
    layer0_outputs(840) <= inputs(157);
    layer0_outputs(841) <= not(inputs(153)) or (inputs(68));
    layer0_outputs(842) <= not((inputs(86)) or (inputs(79)));
    layer0_outputs(843) <= (inputs(144)) xor (inputs(94));
    layer0_outputs(844) <= not((inputs(208)) xor (inputs(230)));
    layer0_outputs(845) <= not(inputs(119));
    layer0_outputs(846) <= not((inputs(99)) or (inputs(98)));
    layer0_outputs(847) <= '0';
    layer0_outputs(848) <= not(inputs(255));
    layer0_outputs(849) <= not((inputs(255)) xor (inputs(210)));
    layer0_outputs(850) <= not(inputs(60)) or (inputs(227));
    layer0_outputs(851) <= inputs(137);
    layer0_outputs(852) <= inputs(199);
    layer0_outputs(853) <= not(inputs(117));
    layer0_outputs(854) <= (inputs(121)) and (inputs(170));
    layer0_outputs(855) <= (inputs(187)) or (inputs(35));
    layer0_outputs(856) <= not(inputs(59));
    layer0_outputs(857) <= (inputs(123)) and not (inputs(207));
    layer0_outputs(858) <= not(inputs(185)) or (inputs(226));
    layer0_outputs(859) <= inputs(189);
    layer0_outputs(860) <= (inputs(242)) or (inputs(101));
    layer0_outputs(861) <= not((inputs(9)) xor (inputs(87)));
    layer0_outputs(862) <= not((inputs(178)) or (inputs(59)));
    layer0_outputs(863) <= not(inputs(88));
    layer0_outputs(864) <= not(inputs(168));
    layer0_outputs(865) <= (inputs(6)) or (inputs(116));
    layer0_outputs(866) <= (inputs(89)) and not (inputs(193));
    layer0_outputs(867) <= not(inputs(136)) or (inputs(166));
    layer0_outputs(868) <= (inputs(119)) or (inputs(107));
    layer0_outputs(869) <= not((inputs(208)) or (inputs(199)));
    layer0_outputs(870) <= not((inputs(10)) and (inputs(80)));
    layer0_outputs(871) <= (inputs(132)) and not (inputs(238));
    layer0_outputs(872) <= not(inputs(41));
    layer0_outputs(873) <= not(inputs(57));
    layer0_outputs(874) <= (inputs(213)) and not (inputs(156));
    layer0_outputs(875) <= not((inputs(143)) xor (inputs(236)));
    layer0_outputs(876) <= not((inputs(240)) and (inputs(61)));
    layer0_outputs(877) <= not(inputs(133)) or (inputs(189));
    layer0_outputs(878) <= (inputs(54)) xor (inputs(20));
    layer0_outputs(879) <= not((inputs(36)) or (inputs(57)));
    layer0_outputs(880) <= not((inputs(191)) and (inputs(254)));
    layer0_outputs(881) <= not((inputs(172)) xor (inputs(65)));
    layer0_outputs(882) <= not(inputs(144)) or (inputs(46));
    layer0_outputs(883) <= (inputs(235)) or (inputs(100));
    layer0_outputs(884) <= inputs(216);
    layer0_outputs(885) <= (inputs(50)) xor (inputs(203));
    layer0_outputs(886) <= (inputs(201)) and not (inputs(234));
    layer0_outputs(887) <= not((inputs(203)) or (inputs(125)));
    layer0_outputs(888) <= not(inputs(196)) or (inputs(248));
    layer0_outputs(889) <= (inputs(59)) xor (inputs(7));
    layer0_outputs(890) <= not(inputs(119)) or (inputs(167));
    layer0_outputs(891) <= not((inputs(157)) or (inputs(187)));
    layer0_outputs(892) <= '0';
    layer0_outputs(893) <= not((inputs(224)) xor (inputs(117)));
    layer0_outputs(894) <= '1';
    layer0_outputs(895) <= not((inputs(75)) or (inputs(84)));
    layer0_outputs(896) <= not(inputs(217)) or (inputs(23));
    layer0_outputs(897) <= (inputs(91)) and not (inputs(236));
    layer0_outputs(898) <= not(inputs(196));
    layer0_outputs(899) <= '1';
    layer0_outputs(900) <= not(inputs(3)) or (inputs(65));
    layer0_outputs(901) <= not((inputs(73)) or (inputs(220)));
    layer0_outputs(902) <= inputs(166);
    layer0_outputs(903) <= not(inputs(180)) or (inputs(235));
    layer0_outputs(904) <= not((inputs(235)) or (inputs(67)));
    layer0_outputs(905) <= not(inputs(51)) or (inputs(60));
    layer0_outputs(906) <= not((inputs(42)) xor (inputs(188)));
    layer0_outputs(907) <= (inputs(253)) and (inputs(79));
    layer0_outputs(908) <= not((inputs(51)) or (inputs(153)));
    layer0_outputs(909) <= not(inputs(24)) or (inputs(51));
    layer0_outputs(910) <= not(inputs(232)) or (inputs(72));
    layer0_outputs(911) <= not((inputs(223)) xor (inputs(82)));
    layer0_outputs(912) <= not((inputs(243)) or (inputs(208)));
    layer0_outputs(913) <= not((inputs(118)) xor (inputs(125)));
    layer0_outputs(914) <= not(inputs(186)) or (inputs(19));
    layer0_outputs(915) <= (inputs(70)) xor (inputs(174));
    layer0_outputs(916) <= not((inputs(220)) or (inputs(123)));
    layer0_outputs(917) <= not((inputs(19)) or (inputs(0)));
    layer0_outputs(918) <= not((inputs(18)) xor (inputs(231)));
    layer0_outputs(919) <= (inputs(11)) and not (inputs(94));
    layer0_outputs(920) <= (inputs(121)) or (inputs(242));
    layer0_outputs(921) <= not(inputs(54));
    layer0_outputs(922) <= '0';
    layer0_outputs(923) <= not((inputs(36)) xor (inputs(175)));
    layer0_outputs(924) <= (inputs(110)) or (inputs(100));
    layer0_outputs(925) <= (inputs(157)) xor (inputs(105));
    layer0_outputs(926) <= not((inputs(185)) xor (inputs(9)));
    layer0_outputs(927) <= (inputs(137)) or (inputs(25));
    layer0_outputs(928) <= inputs(53);
    layer0_outputs(929) <= not((inputs(91)) and (inputs(222)));
    layer0_outputs(930) <= (inputs(151)) xor (inputs(136));
    layer0_outputs(931) <= (inputs(67)) and not (inputs(19));
    layer0_outputs(932) <= (inputs(45)) and not (inputs(111));
    layer0_outputs(933) <= not((inputs(97)) or (inputs(8)));
    layer0_outputs(934) <= not(inputs(107));
    layer0_outputs(935) <= not(inputs(199));
    layer0_outputs(936) <= '1';
    layer0_outputs(937) <= inputs(230);
    layer0_outputs(938) <= (inputs(235)) and not (inputs(145));
    layer0_outputs(939) <= (inputs(42)) xor (inputs(169));
    layer0_outputs(940) <= inputs(76);
    layer0_outputs(941) <= not(inputs(14));
    layer0_outputs(942) <= (inputs(165)) xor (inputs(141));
    layer0_outputs(943) <= inputs(165);
    layer0_outputs(944) <= not((inputs(99)) or (inputs(121)));
    layer0_outputs(945) <= '1';
    layer0_outputs(946) <= not(inputs(41));
    layer0_outputs(947) <= (inputs(49)) xor (inputs(79));
    layer0_outputs(948) <= not(inputs(19)) or (inputs(28));
    layer0_outputs(949) <= (inputs(120)) and not (inputs(189));
    layer0_outputs(950) <= (inputs(86)) or (inputs(75));
    layer0_outputs(951) <= not(inputs(73));
    layer0_outputs(952) <= (inputs(197)) xor (inputs(30));
    layer0_outputs(953) <= not(inputs(170));
    layer0_outputs(954) <= not(inputs(212));
    layer0_outputs(955) <= (inputs(203)) or (inputs(198));
    layer0_outputs(956) <= inputs(150);
    layer0_outputs(957) <= not(inputs(220)) or (inputs(2));
    layer0_outputs(958) <= '1';
    layer0_outputs(959) <= not(inputs(91));
    layer0_outputs(960) <= '0';
    layer0_outputs(961) <= (inputs(207)) and not (inputs(235));
    layer0_outputs(962) <= inputs(1);
    layer0_outputs(963) <= not(inputs(91));
    layer0_outputs(964) <= '0';
    layer0_outputs(965) <= not(inputs(221)) or (inputs(173));
    layer0_outputs(966) <= (inputs(3)) and (inputs(34));
    layer0_outputs(967) <= inputs(127);
    layer0_outputs(968) <= not(inputs(153));
    layer0_outputs(969) <= inputs(107);
    layer0_outputs(970) <= (inputs(107)) or (inputs(221));
    layer0_outputs(971) <= not((inputs(191)) or (inputs(19)));
    layer0_outputs(972) <= (inputs(88)) and not (inputs(243));
    layer0_outputs(973) <= inputs(137);
    layer0_outputs(974) <= not(inputs(122));
    layer0_outputs(975) <= (inputs(203)) xor (inputs(135));
    layer0_outputs(976) <= not(inputs(107)) or (inputs(195));
    layer0_outputs(977) <= not(inputs(143)) or (inputs(3));
    layer0_outputs(978) <= (inputs(209)) xor (inputs(91));
    layer0_outputs(979) <= not((inputs(161)) or (inputs(238)));
    layer0_outputs(980) <= (inputs(220)) xor (inputs(79));
    layer0_outputs(981) <= '0';
    layer0_outputs(982) <= (inputs(69)) xor (inputs(235));
    layer0_outputs(983) <= not(inputs(124)) or (inputs(111));
    layer0_outputs(984) <= not((inputs(19)) and (inputs(176)));
    layer0_outputs(985) <= (inputs(57)) xor (inputs(219));
    layer0_outputs(986) <= not((inputs(98)) or (inputs(173)));
    layer0_outputs(987) <= (inputs(70)) and not (inputs(195));
    layer0_outputs(988) <= not(inputs(216)) or (inputs(96));
    layer0_outputs(989) <= (inputs(18)) or (inputs(221));
    layer0_outputs(990) <= not((inputs(34)) or (inputs(202)));
    layer0_outputs(991) <= inputs(132);
    layer0_outputs(992) <= '1';
    layer0_outputs(993) <= not(inputs(74));
    layer0_outputs(994) <= (inputs(40)) and (inputs(90));
    layer0_outputs(995) <= inputs(159);
    layer0_outputs(996) <= not(inputs(77));
    layer0_outputs(997) <= (inputs(95)) or (inputs(208));
    layer0_outputs(998) <= (inputs(50)) and not (inputs(208));
    layer0_outputs(999) <= not((inputs(182)) xor (inputs(74)));
    layer0_outputs(1000) <= not(inputs(136)) or (inputs(48));
    layer0_outputs(1001) <= (inputs(86)) xor (inputs(8));
    layer0_outputs(1002) <= (inputs(68)) or (inputs(50));
    layer0_outputs(1003) <= (inputs(75)) xor (inputs(120));
    layer0_outputs(1004) <= (inputs(48)) and not (inputs(1));
    layer0_outputs(1005) <= (inputs(234)) or (inputs(85));
    layer0_outputs(1006) <= not(inputs(122)) or (inputs(73));
    layer0_outputs(1007) <= not(inputs(79));
    layer0_outputs(1008) <= (inputs(83)) or (inputs(150));
    layer0_outputs(1009) <= (inputs(182)) or (inputs(166));
    layer0_outputs(1010) <= (inputs(171)) or (inputs(107));
    layer0_outputs(1011) <= not(inputs(36));
    layer0_outputs(1012) <= '1';
    layer0_outputs(1013) <= not(inputs(54)) or (inputs(26));
    layer0_outputs(1014) <= not(inputs(160)) or (inputs(27));
    layer0_outputs(1015) <= inputs(171);
    layer0_outputs(1016) <= inputs(162);
    layer0_outputs(1017) <= not((inputs(60)) xor (inputs(43)));
    layer0_outputs(1018) <= not(inputs(38)) or (inputs(32));
    layer0_outputs(1019) <= not((inputs(202)) or (inputs(211)));
    layer0_outputs(1020) <= (inputs(167)) and not (inputs(131));
    layer0_outputs(1021) <= not(inputs(117)) or (inputs(245));
    layer0_outputs(1022) <= not(inputs(216)) or (inputs(165));
    layer0_outputs(1023) <= inputs(231);
    layer0_outputs(1024) <= not(inputs(90)) or (inputs(246));
    layer0_outputs(1025) <= '0';
    layer0_outputs(1026) <= not((inputs(199)) and (inputs(89)));
    layer0_outputs(1027) <= not((inputs(97)) or (inputs(86)));
    layer0_outputs(1028) <= (inputs(153)) and not (inputs(200));
    layer0_outputs(1029) <= (inputs(197)) xor (inputs(0));
    layer0_outputs(1030) <= not((inputs(146)) or (inputs(212)));
    layer0_outputs(1031) <= not((inputs(55)) or (inputs(189)));
    layer0_outputs(1032) <= not((inputs(96)) xor (inputs(211)));
    layer0_outputs(1033) <= not((inputs(209)) or (inputs(231)));
    layer0_outputs(1034) <= not(inputs(211)) or (inputs(8));
    layer0_outputs(1035) <= inputs(104);
    layer0_outputs(1036) <= not(inputs(249)) or (inputs(107));
    layer0_outputs(1037) <= not((inputs(198)) or (inputs(109)));
    layer0_outputs(1038) <= not((inputs(129)) xor (inputs(44)));
    layer0_outputs(1039) <= not((inputs(103)) xor (inputs(116)));
    layer0_outputs(1040) <= (inputs(127)) or (inputs(167));
    layer0_outputs(1041) <= inputs(79);
    layer0_outputs(1042) <= not((inputs(120)) xor (inputs(180)));
    layer0_outputs(1043) <= inputs(216);
    layer0_outputs(1044) <= (inputs(174)) and (inputs(46));
    layer0_outputs(1045) <= not((inputs(69)) or (inputs(68)));
    layer0_outputs(1046) <= not(inputs(227));
    layer0_outputs(1047) <= not(inputs(182)) or (inputs(228));
    layer0_outputs(1048) <= inputs(168);
    layer0_outputs(1049) <= not((inputs(179)) or (inputs(69)));
    layer0_outputs(1050) <= not((inputs(168)) or (inputs(96)));
    layer0_outputs(1051) <= not((inputs(72)) or (inputs(23)));
    layer0_outputs(1052) <= not(inputs(64));
    layer0_outputs(1053) <= not((inputs(184)) or (inputs(96)));
    layer0_outputs(1054) <= inputs(6);
    layer0_outputs(1055) <= not(inputs(221)) or (inputs(32));
    layer0_outputs(1056) <= (inputs(64)) and (inputs(177));
    layer0_outputs(1057) <= inputs(110);
    layer0_outputs(1058) <= not(inputs(219)) or (inputs(47));
    layer0_outputs(1059) <= not((inputs(38)) xor (inputs(80)));
    layer0_outputs(1060) <= not((inputs(53)) or (inputs(13)));
    layer0_outputs(1061) <= inputs(46);
    layer0_outputs(1062) <= not(inputs(72)) or (inputs(236));
    layer0_outputs(1063) <= not((inputs(168)) xor (inputs(43)));
    layer0_outputs(1064) <= inputs(112);
    layer0_outputs(1065) <= (inputs(44)) or (inputs(193));
    layer0_outputs(1066) <= not((inputs(65)) or (inputs(241)));
    layer0_outputs(1067) <= '0';
    layer0_outputs(1068) <= (inputs(250)) or (inputs(121));
    layer0_outputs(1069) <= not(inputs(13));
    layer0_outputs(1070) <= not(inputs(191));
    layer0_outputs(1071) <= not(inputs(69)) or (inputs(250));
    layer0_outputs(1072) <= (inputs(62)) or (inputs(249));
    layer0_outputs(1073) <= (inputs(32)) and not (inputs(3));
    layer0_outputs(1074) <= (inputs(154)) or (inputs(127));
    layer0_outputs(1075) <= not((inputs(94)) or (inputs(218)));
    layer0_outputs(1076) <= not((inputs(157)) xor (inputs(242)));
    layer0_outputs(1077) <= not(inputs(93));
    layer0_outputs(1078) <= inputs(78);
    layer0_outputs(1079) <= not((inputs(212)) or (inputs(213)));
    layer0_outputs(1080) <= inputs(43);
    layer0_outputs(1081) <= not(inputs(204)) or (inputs(161));
    layer0_outputs(1082) <= not((inputs(207)) and (inputs(209)));
    layer0_outputs(1083) <= (inputs(239)) or (inputs(122));
    layer0_outputs(1084) <= not(inputs(200)) or (inputs(5));
    layer0_outputs(1085) <= inputs(119);
    layer0_outputs(1086) <= not(inputs(151));
    layer0_outputs(1087) <= inputs(3);
    layer0_outputs(1088) <= not((inputs(212)) xor (inputs(85)));
    layer0_outputs(1089) <= (inputs(230)) xor (inputs(5));
    layer0_outputs(1090) <= inputs(135);
    layer0_outputs(1091) <= not(inputs(51)) or (inputs(110));
    layer0_outputs(1092) <= inputs(205);
    layer0_outputs(1093) <= (inputs(74)) and not (inputs(64));
    layer0_outputs(1094) <= not(inputs(204)) or (inputs(224));
    layer0_outputs(1095) <= not(inputs(39)) or (inputs(255));
    layer0_outputs(1096) <= not(inputs(104));
    layer0_outputs(1097) <= not(inputs(214));
    layer0_outputs(1098) <= (inputs(217)) or (inputs(224));
    layer0_outputs(1099) <= not((inputs(192)) or (inputs(1)));
    layer0_outputs(1100) <= (inputs(128)) xor (inputs(48));
    layer0_outputs(1101) <= not((inputs(5)) xor (inputs(148)));
    layer0_outputs(1102) <= not((inputs(25)) xor (inputs(114)));
    layer0_outputs(1103) <= (inputs(170)) and not (inputs(211));
    layer0_outputs(1104) <= not((inputs(51)) and (inputs(51)));
    layer0_outputs(1105) <= (inputs(31)) and not (inputs(136));
    layer0_outputs(1106) <= not(inputs(15));
    layer0_outputs(1107) <= '1';
    layer0_outputs(1108) <= not(inputs(199));
    layer0_outputs(1109) <= (inputs(45)) or (inputs(247));
    layer0_outputs(1110) <= (inputs(73)) xor (inputs(251));
    layer0_outputs(1111) <= not((inputs(131)) and (inputs(127)));
    layer0_outputs(1112) <= (inputs(166)) or (inputs(229));
    layer0_outputs(1113) <= not(inputs(114));
    layer0_outputs(1114) <= '1';
    layer0_outputs(1115) <= not(inputs(88)) or (inputs(22));
    layer0_outputs(1116) <= not((inputs(72)) or (inputs(62)));
    layer0_outputs(1117) <= (inputs(37)) and not (inputs(250));
    layer0_outputs(1118) <= (inputs(67)) and (inputs(32));
    layer0_outputs(1119) <= not(inputs(202)) or (inputs(126));
    layer0_outputs(1120) <= not(inputs(138));
    layer0_outputs(1121) <= not(inputs(73)) or (inputs(241));
    layer0_outputs(1122) <= not(inputs(86)) or (inputs(160));
    layer0_outputs(1123) <= '0';
    layer0_outputs(1124) <= (inputs(37)) or (inputs(25));
    layer0_outputs(1125) <= not(inputs(111));
    layer0_outputs(1126) <= inputs(213);
    layer0_outputs(1127) <= (inputs(167)) xor (inputs(173));
    layer0_outputs(1128) <= '0';
    layer0_outputs(1129) <= not(inputs(119)) or (inputs(253));
    layer0_outputs(1130) <= not((inputs(73)) xor (inputs(111)));
    layer0_outputs(1131) <= (inputs(167)) or (inputs(77));
    layer0_outputs(1132) <= not(inputs(36));
    layer0_outputs(1133) <= inputs(220);
    layer0_outputs(1134) <= (inputs(192)) and not (inputs(163));
    layer0_outputs(1135) <= (inputs(202)) or (inputs(63));
    layer0_outputs(1136) <= not((inputs(145)) or (inputs(100)));
    layer0_outputs(1137) <= (inputs(83)) xor (inputs(113));
    layer0_outputs(1138) <= (inputs(165)) or (inputs(182));
    layer0_outputs(1139) <= (inputs(97)) xor (inputs(58));
    layer0_outputs(1140) <= inputs(55);
    layer0_outputs(1141) <= (inputs(179)) xor (inputs(30));
    layer0_outputs(1142) <= (inputs(156)) or (inputs(207));
    layer0_outputs(1143) <= '1';
    layer0_outputs(1144) <= (inputs(211)) or (inputs(196));
    layer0_outputs(1145) <= '0';
    layer0_outputs(1146) <= inputs(197);
    layer0_outputs(1147) <= (inputs(212)) xor (inputs(109));
    layer0_outputs(1148) <= not(inputs(16)) or (inputs(236));
    layer0_outputs(1149) <= inputs(111);
    layer0_outputs(1150) <= (inputs(36)) or (inputs(150));
    layer0_outputs(1151) <= not((inputs(33)) or (inputs(68)));
    layer0_outputs(1152) <= not((inputs(96)) or (inputs(75)));
    layer0_outputs(1153) <= (inputs(174)) or (inputs(165));
    layer0_outputs(1154) <= '1';
    layer0_outputs(1155) <= not(inputs(186));
    layer0_outputs(1156) <= not((inputs(52)) xor (inputs(132)));
    layer0_outputs(1157) <= (inputs(43)) and not (inputs(190));
    layer0_outputs(1158) <= not((inputs(10)) and (inputs(243)));
    layer0_outputs(1159) <= inputs(46);
    layer0_outputs(1160) <= (inputs(132)) xor (inputs(234));
    layer0_outputs(1161) <= inputs(242);
    layer0_outputs(1162) <= '1';
    layer0_outputs(1163) <= (inputs(117)) or (inputs(141));
    layer0_outputs(1164) <= inputs(117);
    layer0_outputs(1165) <= inputs(121);
    layer0_outputs(1166) <= not((inputs(43)) or (inputs(125)));
    layer0_outputs(1167) <= not(inputs(226)) or (inputs(116));
    layer0_outputs(1168) <= (inputs(123)) xor (inputs(116));
    layer0_outputs(1169) <= (inputs(218)) and (inputs(246));
    layer0_outputs(1170) <= not((inputs(231)) or (inputs(246)));
    layer0_outputs(1171) <= not(inputs(83)) or (inputs(178));
    layer0_outputs(1172) <= not(inputs(41)) or (inputs(145));
    layer0_outputs(1173) <= (inputs(164)) and not (inputs(27));
    layer0_outputs(1174) <= '1';
    layer0_outputs(1175) <= not((inputs(238)) and (inputs(36)));
    layer0_outputs(1176) <= not(inputs(117)) or (inputs(219));
    layer0_outputs(1177) <= not(inputs(53)) or (inputs(248));
    layer0_outputs(1178) <= not(inputs(46));
    layer0_outputs(1179) <= inputs(76);
    layer0_outputs(1180) <= '0';
    layer0_outputs(1181) <= (inputs(198)) and not (inputs(35));
    layer0_outputs(1182) <= inputs(183);
    layer0_outputs(1183) <= not(inputs(55));
    layer0_outputs(1184) <= (inputs(177)) and not (inputs(247));
    layer0_outputs(1185) <= (inputs(238)) or (inputs(200));
    layer0_outputs(1186) <= inputs(132);
    layer0_outputs(1187) <= (inputs(221)) or (inputs(72));
    layer0_outputs(1188) <= not(inputs(102)) or (inputs(39));
    layer0_outputs(1189) <= '0';
    layer0_outputs(1190) <= not((inputs(40)) or (inputs(134)));
    layer0_outputs(1191) <= '1';
    layer0_outputs(1192) <= (inputs(201)) and not (inputs(24));
    layer0_outputs(1193) <= (inputs(85)) xor (inputs(129));
    layer0_outputs(1194) <= '1';
    layer0_outputs(1195) <= not(inputs(59)) or (inputs(222));
    layer0_outputs(1196) <= (inputs(132)) or (inputs(188));
    layer0_outputs(1197) <= not(inputs(221)) or (inputs(99));
    layer0_outputs(1198) <= (inputs(204)) or (inputs(50));
    layer0_outputs(1199) <= (inputs(8)) xor (inputs(88));
    layer0_outputs(1200) <= not(inputs(182)) or (inputs(243));
    layer0_outputs(1201) <= not((inputs(73)) or (inputs(122)));
    layer0_outputs(1202) <= (inputs(161)) or (inputs(163));
    layer0_outputs(1203) <= '0';
    layer0_outputs(1204) <= not(inputs(151)) or (inputs(98));
    layer0_outputs(1205) <= (inputs(62)) xor (inputs(202));
    layer0_outputs(1206) <= not(inputs(11));
    layer0_outputs(1207) <= inputs(82);
    layer0_outputs(1208) <= (inputs(85)) and not (inputs(172));
    layer0_outputs(1209) <= (inputs(169)) and (inputs(53));
    layer0_outputs(1210) <= not((inputs(86)) xor (inputs(70)));
    layer0_outputs(1211) <= (inputs(66)) xor (inputs(5));
    layer0_outputs(1212) <= not(inputs(226)) or (inputs(239));
    layer0_outputs(1213) <= (inputs(75)) and not (inputs(147));
    layer0_outputs(1214) <= not(inputs(106));
    layer0_outputs(1215) <= not(inputs(76)) or (inputs(3));
    layer0_outputs(1216) <= (inputs(202)) and not (inputs(184));
    layer0_outputs(1217) <= (inputs(1)) and not (inputs(203));
    layer0_outputs(1218) <= (inputs(234)) or (inputs(249));
    layer0_outputs(1219) <= not((inputs(39)) and (inputs(200)));
    layer0_outputs(1220) <= not(inputs(150));
    layer0_outputs(1221) <= inputs(59);
    layer0_outputs(1222) <= (inputs(235)) and not (inputs(30));
    layer0_outputs(1223) <= not(inputs(119)) or (inputs(165));
    layer0_outputs(1224) <= inputs(10);
    layer0_outputs(1225) <= (inputs(249)) or (inputs(228));
    layer0_outputs(1226) <= not((inputs(235)) or (inputs(190)));
    layer0_outputs(1227) <= inputs(245);
    layer0_outputs(1228) <= (inputs(166)) and not (inputs(233));
    layer0_outputs(1229) <= not(inputs(60)) or (inputs(138));
    layer0_outputs(1230) <= not(inputs(166)) or (inputs(132));
    layer0_outputs(1231) <= not((inputs(244)) xor (inputs(60)));
    layer0_outputs(1232) <= not((inputs(23)) or (inputs(147)));
    layer0_outputs(1233) <= not(inputs(107));
    layer0_outputs(1234) <= inputs(158);
    layer0_outputs(1235) <= not(inputs(92)) or (inputs(19));
    layer0_outputs(1236) <= inputs(53);
    layer0_outputs(1237) <= not((inputs(32)) xor (inputs(65)));
    layer0_outputs(1238) <= not(inputs(1)) or (inputs(173));
    layer0_outputs(1239) <= (inputs(36)) and not (inputs(29));
    layer0_outputs(1240) <= not((inputs(59)) xor (inputs(2)));
    layer0_outputs(1241) <= not((inputs(152)) xor (inputs(128)));
    layer0_outputs(1242) <= (inputs(78)) and not (inputs(241));
    layer0_outputs(1243) <= (inputs(166)) or (inputs(32));
    layer0_outputs(1244) <= (inputs(82)) or (inputs(215));
    layer0_outputs(1245) <= not(inputs(204));
    layer0_outputs(1246) <= not((inputs(161)) xor (inputs(234)));
    layer0_outputs(1247) <= not(inputs(169));
    layer0_outputs(1248) <= (inputs(184)) and not (inputs(33));
    layer0_outputs(1249) <= not((inputs(109)) or (inputs(113)));
    layer0_outputs(1250) <= inputs(139);
    layer0_outputs(1251) <= not((inputs(51)) or (inputs(193)));
    layer0_outputs(1252) <= (inputs(219)) and not (inputs(232));
    layer0_outputs(1253) <= inputs(114);
    layer0_outputs(1254) <= not((inputs(119)) or (inputs(206)));
    layer0_outputs(1255) <= (inputs(115)) xor (inputs(255));
    layer0_outputs(1256) <= (inputs(91)) and not (inputs(23));
    layer0_outputs(1257) <= (inputs(145)) and not (inputs(236));
    layer0_outputs(1258) <= (inputs(116)) and not (inputs(83));
    layer0_outputs(1259) <= not(inputs(198));
    layer0_outputs(1260) <= not(inputs(154));
    layer0_outputs(1261) <= (inputs(48)) and (inputs(176));
    layer0_outputs(1262) <= (inputs(237)) or (inputs(40));
    layer0_outputs(1263) <= not((inputs(114)) xor (inputs(109)));
    layer0_outputs(1264) <= not(inputs(77)) or (inputs(24));
    layer0_outputs(1265) <= not(inputs(172)) or (inputs(251));
    layer0_outputs(1266) <= not((inputs(90)) xor (inputs(33)));
    layer0_outputs(1267) <= (inputs(138)) or (inputs(250));
    layer0_outputs(1268) <= not((inputs(78)) or (inputs(135)));
    layer0_outputs(1269) <= (inputs(118)) and not (inputs(8));
    layer0_outputs(1270) <= (inputs(158)) and not (inputs(188));
    layer0_outputs(1271) <= (inputs(112)) xor (inputs(89));
    layer0_outputs(1272) <= (inputs(193)) xor (inputs(87));
    layer0_outputs(1273) <= not(inputs(149));
    layer0_outputs(1274) <= not((inputs(60)) xor (inputs(183)));
    layer0_outputs(1275) <= (inputs(177)) xor (inputs(28));
    layer0_outputs(1276) <= (inputs(199)) or (inputs(177));
    layer0_outputs(1277) <= (inputs(59)) and not (inputs(237));
    layer0_outputs(1278) <= inputs(37);
    layer0_outputs(1279) <= '0';
    layer0_outputs(1280) <= (inputs(214)) or (inputs(124));
    layer0_outputs(1281) <= not(inputs(192));
    layer0_outputs(1282) <= (inputs(253)) xor (inputs(33));
    layer0_outputs(1283) <= inputs(10);
    layer0_outputs(1284) <= not((inputs(150)) xor (inputs(221)));
    layer0_outputs(1285) <= not(inputs(249)) or (inputs(4));
    layer0_outputs(1286) <= inputs(138);
    layer0_outputs(1287) <= (inputs(22)) xor (inputs(201));
    layer0_outputs(1288) <= (inputs(70)) and not (inputs(239));
    layer0_outputs(1289) <= not(inputs(167));
    layer0_outputs(1290) <= not(inputs(63));
    layer0_outputs(1291) <= not(inputs(198)) or (inputs(173));
    layer0_outputs(1292) <= not((inputs(108)) xor (inputs(225)));
    layer0_outputs(1293) <= not((inputs(235)) or (inputs(39)));
    layer0_outputs(1294) <= inputs(239);
    layer0_outputs(1295) <= not(inputs(87)) or (inputs(158));
    layer0_outputs(1296) <= not((inputs(199)) or (inputs(34)));
    layer0_outputs(1297) <= not(inputs(196));
    layer0_outputs(1298) <= (inputs(59)) and (inputs(39));
    layer0_outputs(1299) <= '1';
    layer0_outputs(1300) <= inputs(58);
    layer0_outputs(1301) <= not(inputs(168)) or (inputs(180));
    layer0_outputs(1302) <= not((inputs(37)) xor (inputs(8)));
    layer0_outputs(1303) <= (inputs(89)) xor (inputs(112));
    layer0_outputs(1304) <= not(inputs(116));
    layer0_outputs(1305) <= (inputs(111)) or (inputs(98));
    layer0_outputs(1306) <= not(inputs(67)) or (inputs(31));
    layer0_outputs(1307) <= not(inputs(155)) or (inputs(199));
    layer0_outputs(1308) <= '1';
    layer0_outputs(1309) <= (inputs(200)) or (inputs(244));
    layer0_outputs(1310) <= not(inputs(198)) or (inputs(81));
    layer0_outputs(1311) <= (inputs(148)) xor (inputs(248));
    layer0_outputs(1312) <= inputs(162);
    layer0_outputs(1313) <= (inputs(184)) and not (inputs(7));
    layer0_outputs(1314) <= not((inputs(204)) or (inputs(179)));
    layer0_outputs(1315) <= (inputs(133)) and not (inputs(180));
    layer0_outputs(1316) <= not(inputs(170)) or (inputs(130));
    layer0_outputs(1317) <= (inputs(90)) and not (inputs(53));
    layer0_outputs(1318) <= not(inputs(173)) or (inputs(27));
    layer0_outputs(1319) <= not(inputs(48));
    layer0_outputs(1320) <= not((inputs(181)) xor (inputs(238)));
    layer0_outputs(1321) <= (inputs(13)) or (inputs(191));
    layer0_outputs(1322) <= (inputs(204)) or (inputs(221));
    layer0_outputs(1323) <= not((inputs(118)) xor (inputs(218)));
    layer0_outputs(1324) <= not(inputs(166));
    layer0_outputs(1325) <= not(inputs(183)) or (inputs(217));
    layer0_outputs(1326) <= '0';
    layer0_outputs(1327) <= inputs(60);
    layer0_outputs(1328) <= (inputs(52)) xor (inputs(148));
    layer0_outputs(1329) <= (inputs(65)) or (inputs(243));
    layer0_outputs(1330) <= not((inputs(139)) or (inputs(85)));
    layer0_outputs(1331) <= (inputs(23)) or (inputs(182));
    layer0_outputs(1332) <= (inputs(184)) or (inputs(157));
    layer0_outputs(1333) <= not((inputs(57)) xor (inputs(44)));
    layer0_outputs(1334) <= not((inputs(26)) and (inputs(196)));
    layer0_outputs(1335) <= (inputs(71)) and not (inputs(142));
    layer0_outputs(1336) <= not(inputs(141));
    layer0_outputs(1337) <= (inputs(194)) or (inputs(78));
    layer0_outputs(1338) <= not(inputs(18));
    layer0_outputs(1339) <= (inputs(149)) and not (inputs(110));
    layer0_outputs(1340) <= inputs(231);
    layer0_outputs(1341) <= not(inputs(147));
    layer0_outputs(1342) <= not((inputs(87)) or (inputs(77)));
    layer0_outputs(1343) <= not(inputs(184));
    layer0_outputs(1344) <= (inputs(115)) and not (inputs(50));
    layer0_outputs(1345) <= not(inputs(158));
    layer0_outputs(1346) <= (inputs(155)) xor (inputs(124));
    layer0_outputs(1347) <= (inputs(228)) or (inputs(113));
    layer0_outputs(1348) <= not(inputs(152)) or (inputs(98));
    layer0_outputs(1349) <= not((inputs(131)) or (inputs(215)));
    layer0_outputs(1350) <= (inputs(88)) and not (inputs(9));
    layer0_outputs(1351) <= (inputs(86)) xor (inputs(6));
    layer0_outputs(1352) <= (inputs(221)) or (inputs(221));
    layer0_outputs(1353) <= not(inputs(47)) or (inputs(226));
    layer0_outputs(1354) <= inputs(203);
    layer0_outputs(1355) <= not((inputs(22)) xor (inputs(195)));
    layer0_outputs(1356) <= '1';
    layer0_outputs(1357) <= (inputs(158)) and not (inputs(110));
    layer0_outputs(1358) <= not(inputs(120)) or (inputs(143));
    layer0_outputs(1359) <= (inputs(59)) and (inputs(195));
    layer0_outputs(1360) <= inputs(117);
    layer0_outputs(1361) <= (inputs(102)) and not (inputs(108));
    layer0_outputs(1362) <= (inputs(163)) or (inputs(180));
    layer0_outputs(1363) <= not((inputs(253)) xor (inputs(151)));
    layer0_outputs(1364) <= not(inputs(88)) or (inputs(1));
    layer0_outputs(1365) <= not((inputs(174)) and (inputs(71)));
    layer0_outputs(1366) <= (inputs(191)) and not (inputs(174));
    layer0_outputs(1367) <= (inputs(8)) or (inputs(93));
    layer0_outputs(1368) <= not(inputs(57)) or (inputs(177));
    layer0_outputs(1369) <= not((inputs(226)) and (inputs(32)));
    layer0_outputs(1370) <= not(inputs(199));
    layer0_outputs(1371) <= not(inputs(67)) or (inputs(219));
    layer0_outputs(1372) <= (inputs(53)) and not (inputs(10));
    layer0_outputs(1373) <= not(inputs(117));
    layer0_outputs(1374) <= not(inputs(102));
    layer0_outputs(1375) <= inputs(220);
    layer0_outputs(1376) <= not((inputs(73)) or (inputs(215)));
    layer0_outputs(1377) <= (inputs(254)) and not (inputs(50));
    layer0_outputs(1378) <= inputs(246);
    layer0_outputs(1379) <= not(inputs(1)) or (inputs(241));
    layer0_outputs(1380) <= inputs(102);
    layer0_outputs(1381) <= inputs(117);
    layer0_outputs(1382) <= not((inputs(75)) xor (inputs(31)));
    layer0_outputs(1383) <= not(inputs(227)) or (inputs(190));
    layer0_outputs(1384) <= not(inputs(171)) or (inputs(61));
    layer0_outputs(1385) <= not((inputs(226)) and (inputs(17)));
    layer0_outputs(1386) <= not((inputs(88)) xor (inputs(194)));
    layer0_outputs(1387) <= not((inputs(252)) xor (inputs(188)));
    layer0_outputs(1388) <= not((inputs(114)) or (inputs(168)));
    layer0_outputs(1389) <= not(inputs(197));
    layer0_outputs(1390) <= not(inputs(152));
    layer0_outputs(1391) <= not(inputs(66));
    layer0_outputs(1392) <= not(inputs(108));
    layer0_outputs(1393) <= (inputs(245)) xor (inputs(101));
    layer0_outputs(1394) <= not((inputs(68)) and (inputs(177)));
    layer0_outputs(1395) <= not((inputs(246)) and (inputs(238)));
    layer0_outputs(1396) <= not((inputs(142)) xor (inputs(73)));
    layer0_outputs(1397) <= not(inputs(56)) or (inputs(1));
    layer0_outputs(1398) <= inputs(102);
    layer0_outputs(1399) <= (inputs(95)) or (inputs(140));
    layer0_outputs(1400) <= (inputs(249)) and not (inputs(9));
    layer0_outputs(1401) <= not(inputs(55));
    layer0_outputs(1402) <= not(inputs(186));
    layer0_outputs(1403) <= not((inputs(98)) xor (inputs(162)));
    layer0_outputs(1404) <= (inputs(40)) or (inputs(26));
    layer0_outputs(1405) <= (inputs(242)) and not (inputs(62));
    layer0_outputs(1406) <= not(inputs(92));
    layer0_outputs(1407) <= not(inputs(119));
    layer0_outputs(1408) <= '0';
    layer0_outputs(1409) <= not(inputs(32));
    layer0_outputs(1410) <= (inputs(179)) xor (inputs(11));
    layer0_outputs(1411) <= not((inputs(211)) or (inputs(247)));
    layer0_outputs(1412) <= inputs(42);
    layer0_outputs(1413) <= (inputs(114)) xor (inputs(242));
    layer0_outputs(1414) <= not(inputs(82)) or (inputs(38));
    layer0_outputs(1415) <= (inputs(128)) xor (inputs(107));
    layer0_outputs(1416) <= not((inputs(168)) or (inputs(34)));
    layer0_outputs(1417) <= (inputs(153)) xor (inputs(247));
    layer0_outputs(1418) <= (inputs(71)) and not (inputs(58));
    layer0_outputs(1419) <= inputs(113);
    layer0_outputs(1420) <= (inputs(162)) or (inputs(254));
    layer0_outputs(1421) <= (inputs(30)) xor (inputs(152));
    layer0_outputs(1422) <= (inputs(102)) and not (inputs(240));
    layer0_outputs(1423) <= not(inputs(125)) or (inputs(78));
    layer0_outputs(1424) <= inputs(60);
    layer0_outputs(1425) <= not(inputs(238)) or (inputs(5));
    layer0_outputs(1426) <= (inputs(65)) or (inputs(63));
    layer0_outputs(1427) <= not(inputs(190));
    layer0_outputs(1428) <= (inputs(247)) xor (inputs(251));
    layer0_outputs(1429) <= not((inputs(116)) or (inputs(45)));
    layer0_outputs(1430) <= (inputs(192)) and not (inputs(16));
    layer0_outputs(1431) <= inputs(185);
    layer0_outputs(1432) <= (inputs(238)) and (inputs(66));
    layer0_outputs(1433) <= not((inputs(219)) or (inputs(56)));
    layer0_outputs(1434) <= not(inputs(117));
    layer0_outputs(1435) <= (inputs(105)) and not (inputs(14));
    layer0_outputs(1436) <= (inputs(187)) or (inputs(43));
    layer0_outputs(1437) <= not(inputs(112));
    layer0_outputs(1438) <= (inputs(179)) xor (inputs(148));
    layer0_outputs(1439) <= not(inputs(121));
    layer0_outputs(1440) <= not(inputs(101));
    layer0_outputs(1441) <= not((inputs(245)) xor (inputs(235)));
    layer0_outputs(1442) <= (inputs(232)) and not (inputs(36));
    layer0_outputs(1443) <= not(inputs(215));
    layer0_outputs(1444) <= not((inputs(135)) xor (inputs(79)));
    layer0_outputs(1445) <= (inputs(124)) or (inputs(234));
    layer0_outputs(1446) <= inputs(34);
    layer0_outputs(1447) <= (inputs(204)) and not (inputs(99));
    layer0_outputs(1448) <= (inputs(142)) and not (inputs(113));
    layer0_outputs(1449) <= inputs(82);
    layer0_outputs(1450) <= not((inputs(54)) xor (inputs(56)));
    layer0_outputs(1451) <= not((inputs(218)) xor (inputs(234)));
    layer0_outputs(1452) <= (inputs(247)) or (inputs(1));
    layer0_outputs(1453) <= (inputs(11)) xor (inputs(172));
    layer0_outputs(1454) <= (inputs(254)) xor (inputs(191));
    layer0_outputs(1455) <= inputs(234);
    layer0_outputs(1456) <= (inputs(214)) and not (inputs(94));
    layer0_outputs(1457) <= '0';
    layer0_outputs(1458) <= not((inputs(152)) xor (inputs(59)));
    layer0_outputs(1459) <= (inputs(206)) or (inputs(155));
    layer0_outputs(1460) <= not((inputs(65)) or (inputs(88)));
    layer0_outputs(1461) <= inputs(155);
    layer0_outputs(1462) <= not((inputs(170)) xor (inputs(246)));
    layer0_outputs(1463) <= not((inputs(166)) or (inputs(123)));
    layer0_outputs(1464) <= inputs(81);
    layer0_outputs(1465) <= inputs(189);
    layer0_outputs(1466) <= not(inputs(60));
    layer0_outputs(1467) <= (inputs(235)) or (inputs(229));
    layer0_outputs(1468) <= (inputs(7)) or (inputs(152));
    layer0_outputs(1469) <= (inputs(190)) xor (inputs(132));
    layer0_outputs(1470) <= (inputs(44)) xor (inputs(9));
    layer0_outputs(1471) <= inputs(150);
    layer0_outputs(1472) <= '1';
    layer0_outputs(1473) <= not((inputs(5)) or (inputs(35)));
    layer0_outputs(1474) <= not(inputs(177));
    layer0_outputs(1475) <= not(inputs(184));
    layer0_outputs(1476) <= not(inputs(93));
    layer0_outputs(1477) <= (inputs(13)) xor (inputs(54));
    layer0_outputs(1478) <= (inputs(52)) xor (inputs(15));
    layer0_outputs(1479) <= not(inputs(54));
    layer0_outputs(1480) <= not(inputs(150));
    layer0_outputs(1481) <= not(inputs(107));
    layer0_outputs(1482) <= not((inputs(214)) or (inputs(115)));
    layer0_outputs(1483) <= inputs(71);
    layer0_outputs(1484) <= (inputs(165)) and not (inputs(44));
    layer0_outputs(1485) <= not((inputs(181)) or (inputs(71)));
    layer0_outputs(1486) <= (inputs(231)) or (inputs(66));
    layer0_outputs(1487) <= not((inputs(61)) xor (inputs(119)));
    layer0_outputs(1488) <= (inputs(45)) xor (inputs(135));
    layer0_outputs(1489) <= (inputs(240)) and not (inputs(177));
    layer0_outputs(1490) <= not((inputs(235)) or (inputs(155)));
    layer0_outputs(1491) <= not(inputs(72));
    layer0_outputs(1492) <= (inputs(56)) and (inputs(57));
    layer0_outputs(1493) <= inputs(192);
    layer0_outputs(1494) <= inputs(92);
    layer0_outputs(1495) <= not((inputs(82)) or (inputs(61)));
    layer0_outputs(1496) <= not((inputs(247)) or (inputs(199)));
    layer0_outputs(1497) <= not((inputs(213)) xor (inputs(181)));
    layer0_outputs(1498) <= (inputs(120)) or (inputs(156));
    layer0_outputs(1499) <= (inputs(136)) xor (inputs(180));
    layer0_outputs(1500) <= inputs(136);
    layer0_outputs(1501) <= (inputs(77)) xor (inputs(181));
    layer0_outputs(1502) <= not((inputs(201)) xor (inputs(3)));
    layer0_outputs(1503) <= not(inputs(192));
    layer0_outputs(1504) <= (inputs(177)) and (inputs(238));
    layer0_outputs(1505) <= inputs(80);
    layer0_outputs(1506) <= not((inputs(240)) or (inputs(188)));
    layer0_outputs(1507) <= not((inputs(54)) xor (inputs(21)));
    layer0_outputs(1508) <= (inputs(150)) or (inputs(187));
    layer0_outputs(1509) <= not((inputs(86)) xor (inputs(84)));
    layer0_outputs(1510) <= not(inputs(43)) or (inputs(63));
    layer0_outputs(1511) <= not(inputs(72)) or (inputs(142));
    layer0_outputs(1512) <= (inputs(42)) and not (inputs(16));
    layer0_outputs(1513) <= not((inputs(211)) xor (inputs(167)));
    layer0_outputs(1514) <= (inputs(111)) xor (inputs(166));
    layer0_outputs(1515) <= (inputs(194)) or (inputs(193));
    layer0_outputs(1516) <= not(inputs(232)) or (inputs(145));
    layer0_outputs(1517) <= (inputs(7)) xor (inputs(37));
    layer0_outputs(1518) <= not((inputs(84)) or (inputs(92)));
    layer0_outputs(1519) <= not(inputs(10));
    layer0_outputs(1520) <= not((inputs(121)) xor (inputs(177)));
    layer0_outputs(1521) <= not(inputs(95)) or (inputs(16));
    layer0_outputs(1522) <= not(inputs(233)) or (inputs(226));
    layer0_outputs(1523) <= (inputs(225)) and (inputs(251));
    layer0_outputs(1524) <= not(inputs(201)) or (inputs(220));
    layer0_outputs(1525) <= (inputs(26)) or (inputs(224));
    layer0_outputs(1526) <= not((inputs(105)) or (inputs(254)));
    layer0_outputs(1527) <= not((inputs(153)) xor (inputs(105)));
    layer0_outputs(1528) <= not(inputs(21)) or (inputs(198));
    layer0_outputs(1529) <= inputs(51);
    layer0_outputs(1530) <= not((inputs(64)) or (inputs(152)));
    layer0_outputs(1531) <= not((inputs(108)) xor (inputs(113)));
    layer0_outputs(1532) <= not(inputs(41));
    layer0_outputs(1533) <= (inputs(77)) or (inputs(213));
    layer0_outputs(1534) <= not((inputs(107)) or (inputs(89)));
    layer0_outputs(1535) <= inputs(196);
    layer0_outputs(1536) <= inputs(104);
    layer0_outputs(1537) <= (inputs(199)) xor (inputs(6));
    layer0_outputs(1538) <= not((inputs(104)) xor (inputs(177)));
    layer0_outputs(1539) <= (inputs(192)) xor (inputs(200));
    layer0_outputs(1540) <= (inputs(132)) xor (inputs(45));
    layer0_outputs(1541) <= (inputs(80)) and not (inputs(117));
    layer0_outputs(1542) <= (inputs(233)) xor (inputs(235));
    layer0_outputs(1543) <= (inputs(116)) and not (inputs(31));
    layer0_outputs(1544) <= (inputs(70)) and not (inputs(61));
    layer0_outputs(1545) <= inputs(199);
    layer0_outputs(1546) <= (inputs(94)) or (inputs(179));
    layer0_outputs(1547) <= (inputs(211)) and not (inputs(28));
    layer0_outputs(1548) <= (inputs(236)) or (inputs(55));
    layer0_outputs(1549) <= (inputs(240)) and not (inputs(177));
    layer0_outputs(1550) <= (inputs(78)) and not (inputs(228));
    layer0_outputs(1551) <= (inputs(112)) xor (inputs(138));
    layer0_outputs(1552) <= (inputs(245)) xor (inputs(67));
    layer0_outputs(1553) <= not(inputs(64));
    layer0_outputs(1554) <= not((inputs(32)) or (inputs(190)));
    layer0_outputs(1555) <= not((inputs(61)) xor (inputs(227)));
    layer0_outputs(1556) <= not((inputs(147)) or (inputs(117)));
    layer0_outputs(1557) <= (inputs(63)) and (inputs(224));
    layer0_outputs(1558) <= (inputs(71)) and not (inputs(174));
    layer0_outputs(1559) <= inputs(57);
    layer0_outputs(1560) <= (inputs(215)) xor (inputs(83));
    layer0_outputs(1561) <= not(inputs(198));
    layer0_outputs(1562) <= not((inputs(65)) or (inputs(147)));
    layer0_outputs(1563) <= (inputs(176)) and not (inputs(219));
    layer0_outputs(1564) <= (inputs(133)) and not (inputs(249));
    layer0_outputs(1565) <= not((inputs(33)) or (inputs(207)));
    layer0_outputs(1566) <= (inputs(229)) or (inputs(219));
    layer0_outputs(1567) <= not(inputs(189));
    layer0_outputs(1568) <= not((inputs(11)) or (inputs(120)));
    layer0_outputs(1569) <= not((inputs(104)) or (inputs(57)));
    layer0_outputs(1570) <= '0';
    layer0_outputs(1571) <= not((inputs(77)) or (inputs(26)));
    layer0_outputs(1572) <= not(inputs(93)) or (inputs(231));
    layer0_outputs(1573) <= not(inputs(230));
    layer0_outputs(1574) <= (inputs(148)) or (inputs(30));
    layer0_outputs(1575) <= not(inputs(115));
    layer0_outputs(1576) <= inputs(72);
    layer0_outputs(1577) <= (inputs(117)) and not (inputs(114));
    layer0_outputs(1578) <= inputs(166);
    layer0_outputs(1579) <= not(inputs(10)) or (inputs(236));
    layer0_outputs(1580) <= (inputs(43)) xor (inputs(66));
    layer0_outputs(1581) <= inputs(60);
    layer0_outputs(1582) <= (inputs(113)) or (inputs(20));
    layer0_outputs(1583) <= (inputs(243)) and (inputs(163));
    layer0_outputs(1584) <= not(inputs(55)) or (inputs(32));
    layer0_outputs(1585) <= (inputs(148)) and not (inputs(98));
    layer0_outputs(1586) <= (inputs(151)) xor (inputs(168));
    layer0_outputs(1587) <= (inputs(13)) or (inputs(226));
    layer0_outputs(1588) <= inputs(195);
    layer0_outputs(1589) <= (inputs(120)) xor (inputs(240));
    layer0_outputs(1590) <= (inputs(227)) and not (inputs(251));
    layer0_outputs(1591) <= not((inputs(239)) xor (inputs(133)));
    layer0_outputs(1592) <= inputs(183);
    layer0_outputs(1593) <= inputs(116);
    layer0_outputs(1594) <= not((inputs(148)) or (inputs(4)));
    layer0_outputs(1595) <= (inputs(143)) or (inputs(147));
    layer0_outputs(1596) <= inputs(51);
    layer0_outputs(1597) <= (inputs(173)) or (inputs(199));
    layer0_outputs(1598) <= (inputs(214)) or (inputs(104));
    layer0_outputs(1599) <= not(inputs(236));
    layer0_outputs(1600) <= not(inputs(245)) or (inputs(98));
    layer0_outputs(1601) <= inputs(201);
    layer0_outputs(1602) <= not(inputs(89));
    layer0_outputs(1603) <= (inputs(15)) or (inputs(157));
    layer0_outputs(1604) <= not((inputs(94)) xor (inputs(138)));
    layer0_outputs(1605) <= (inputs(151)) and not (inputs(127));
    layer0_outputs(1606) <= inputs(153);
    layer0_outputs(1607) <= not((inputs(14)) xor (inputs(201)));
    layer0_outputs(1608) <= not((inputs(93)) xor (inputs(232)));
    layer0_outputs(1609) <= not((inputs(36)) and (inputs(236)));
    layer0_outputs(1610) <= (inputs(205)) and not (inputs(115));
    layer0_outputs(1611) <= (inputs(52)) or (inputs(255));
    layer0_outputs(1612) <= not(inputs(205)) or (inputs(208));
    layer0_outputs(1613) <= not((inputs(72)) xor (inputs(167)));
    layer0_outputs(1614) <= (inputs(23)) and not (inputs(28));
    layer0_outputs(1615) <= not((inputs(88)) or (inputs(250)));
    layer0_outputs(1616) <= not(inputs(53)) or (inputs(159));
    layer0_outputs(1617) <= inputs(183);
    layer0_outputs(1618) <= not(inputs(27));
    layer0_outputs(1619) <= (inputs(38)) and not (inputs(208));
    layer0_outputs(1620) <= inputs(186);
    layer0_outputs(1621) <= (inputs(243)) and (inputs(221));
    layer0_outputs(1622) <= (inputs(68)) or (inputs(170));
    layer0_outputs(1623) <= not(inputs(132));
    layer0_outputs(1624) <= not((inputs(137)) or (inputs(232)));
    layer0_outputs(1625) <= not(inputs(183)) or (inputs(90));
    layer0_outputs(1626) <= not((inputs(247)) xor (inputs(2)));
    layer0_outputs(1627) <= (inputs(49)) and not (inputs(34));
    layer0_outputs(1628) <= inputs(201);
    layer0_outputs(1629) <= inputs(194);
    layer0_outputs(1630) <= (inputs(2)) and (inputs(12));
    layer0_outputs(1631) <= (inputs(172)) xor (inputs(70));
    layer0_outputs(1632) <= (inputs(106)) and not (inputs(101));
    layer0_outputs(1633) <= (inputs(93)) or (inputs(179));
    layer0_outputs(1634) <= not(inputs(250));
    layer0_outputs(1635) <= (inputs(58)) or (inputs(235));
    layer0_outputs(1636) <= not(inputs(104)) or (inputs(36));
    layer0_outputs(1637) <= (inputs(198)) and not (inputs(202));
    layer0_outputs(1638) <= not(inputs(141));
    layer0_outputs(1639) <= not((inputs(245)) xor (inputs(54)));
    layer0_outputs(1640) <= not((inputs(144)) or (inputs(92)));
    layer0_outputs(1641) <= (inputs(118)) and not (inputs(229));
    layer0_outputs(1642) <= not((inputs(64)) or (inputs(169)));
    layer0_outputs(1643) <= (inputs(231)) xor (inputs(146));
    layer0_outputs(1644) <= not(inputs(51)) or (inputs(47));
    layer0_outputs(1645) <= not(inputs(148));
    layer0_outputs(1646) <= not(inputs(79)) or (inputs(252));
    layer0_outputs(1647) <= not((inputs(122)) xor (inputs(22)));
    layer0_outputs(1648) <= inputs(154);
    layer0_outputs(1649) <= (inputs(45)) xor (inputs(204));
    layer0_outputs(1650) <= not(inputs(252)) or (inputs(128));
    layer0_outputs(1651) <= not((inputs(94)) xor (inputs(125)));
    layer0_outputs(1652) <= not(inputs(106)) or (inputs(29));
    layer0_outputs(1653) <= not((inputs(21)) xor (inputs(55)));
    layer0_outputs(1654) <= not(inputs(100)) or (inputs(248));
    layer0_outputs(1655) <= (inputs(243)) xor (inputs(68));
    layer0_outputs(1656) <= inputs(28);
    layer0_outputs(1657) <= (inputs(104)) or (inputs(181));
    layer0_outputs(1658) <= not((inputs(217)) or (inputs(41)));
    layer0_outputs(1659) <= not((inputs(70)) and (inputs(57)));
    layer0_outputs(1660) <= not((inputs(6)) xor (inputs(209)));
    layer0_outputs(1661) <= (inputs(127)) or (inputs(196));
    layer0_outputs(1662) <= not(inputs(196)) or (inputs(207));
    layer0_outputs(1663) <= not((inputs(226)) or (inputs(134)));
    layer0_outputs(1664) <= not((inputs(229)) and (inputs(8)));
    layer0_outputs(1665) <= (inputs(175)) or (inputs(58));
    layer0_outputs(1666) <= (inputs(121)) and not (inputs(114));
    layer0_outputs(1667) <= not(inputs(72)) or (inputs(234));
    layer0_outputs(1668) <= not(inputs(135)) or (inputs(246));
    layer0_outputs(1669) <= (inputs(36)) or (inputs(174));
    layer0_outputs(1670) <= (inputs(55)) xor (inputs(253));
    layer0_outputs(1671) <= not(inputs(32));
    layer0_outputs(1672) <= (inputs(101)) and not (inputs(240));
    layer0_outputs(1673) <= (inputs(165)) and not (inputs(116));
    layer0_outputs(1674) <= (inputs(110)) xor (inputs(104));
    layer0_outputs(1675) <= (inputs(209)) xor (inputs(4));
    layer0_outputs(1676) <= not(inputs(131));
    layer0_outputs(1677) <= (inputs(232)) and not (inputs(242));
    layer0_outputs(1678) <= (inputs(64)) and not (inputs(249));
    layer0_outputs(1679) <= not(inputs(78)) or (inputs(11));
    layer0_outputs(1680) <= not((inputs(4)) xor (inputs(56)));
    layer0_outputs(1681) <= not((inputs(253)) and (inputs(235)));
    layer0_outputs(1682) <= '1';
    layer0_outputs(1683) <= inputs(147);
    layer0_outputs(1684) <= (inputs(173)) xor (inputs(223));
    layer0_outputs(1685) <= not(inputs(64));
    layer0_outputs(1686) <= (inputs(158)) or (inputs(83));
    layer0_outputs(1687) <= (inputs(122)) and not (inputs(37));
    layer0_outputs(1688) <= not(inputs(254)) or (inputs(83));
    layer0_outputs(1689) <= (inputs(16)) xor (inputs(118));
    layer0_outputs(1690) <= not(inputs(71)) or (inputs(42));
    layer0_outputs(1691) <= not(inputs(114)) or (inputs(207));
    layer0_outputs(1692) <= inputs(25);
    layer0_outputs(1693) <= not((inputs(54)) or (inputs(150)));
    layer0_outputs(1694) <= (inputs(111)) and (inputs(59));
    layer0_outputs(1695) <= not(inputs(29)) or (inputs(134));
    layer0_outputs(1696) <= (inputs(149)) and not (inputs(251));
    layer0_outputs(1697) <= (inputs(231)) and (inputs(247));
    layer0_outputs(1698) <= not(inputs(255));
    layer0_outputs(1699) <= not((inputs(241)) xor (inputs(54)));
    layer0_outputs(1700) <= (inputs(84)) and not (inputs(142));
    layer0_outputs(1701) <= (inputs(70)) and not (inputs(49));
    layer0_outputs(1702) <= not((inputs(56)) xor (inputs(183)));
    layer0_outputs(1703) <= (inputs(33)) xor (inputs(68));
    layer0_outputs(1704) <= (inputs(244)) or (inputs(17));
    layer0_outputs(1705) <= (inputs(87)) and not (inputs(180));
    layer0_outputs(1706) <= not(inputs(135));
    layer0_outputs(1707) <= (inputs(66)) or (inputs(68));
    layer0_outputs(1708) <= not((inputs(76)) or (inputs(215)));
    layer0_outputs(1709) <= (inputs(7)) or (inputs(211));
    layer0_outputs(1710) <= inputs(247);
    layer0_outputs(1711) <= not(inputs(253));
    layer0_outputs(1712) <= inputs(38);
    layer0_outputs(1713) <= not(inputs(182));
    layer0_outputs(1714) <= inputs(254);
    layer0_outputs(1715) <= not(inputs(19));
    layer0_outputs(1716) <= (inputs(215)) and not (inputs(95));
    layer0_outputs(1717) <= not((inputs(156)) xor (inputs(105)));
    layer0_outputs(1718) <= (inputs(126)) xor (inputs(195));
    layer0_outputs(1719) <= inputs(189);
    layer0_outputs(1720) <= (inputs(235)) xor (inputs(11));
    layer0_outputs(1721) <= (inputs(186)) and not (inputs(154));
    layer0_outputs(1722) <= not(inputs(55)) or (inputs(234));
    layer0_outputs(1723) <= not(inputs(79)) or (inputs(48));
    layer0_outputs(1724) <= not((inputs(248)) xor (inputs(42)));
    layer0_outputs(1725) <= not((inputs(55)) or (inputs(247)));
    layer0_outputs(1726) <= not((inputs(144)) or (inputs(218)));
    layer0_outputs(1727) <= (inputs(64)) or (inputs(109));
    layer0_outputs(1728) <= (inputs(137)) and not (inputs(17));
    layer0_outputs(1729) <= not(inputs(245));
    layer0_outputs(1730) <= (inputs(64)) and not (inputs(228));
    layer0_outputs(1731) <= inputs(140);
    layer0_outputs(1732) <= inputs(84);
    layer0_outputs(1733) <= not((inputs(247)) xor (inputs(155)));
    layer0_outputs(1734) <= not(inputs(82)) or (inputs(111));
    layer0_outputs(1735) <= (inputs(69)) and not (inputs(204));
    layer0_outputs(1736) <= not((inputs(2)) xor (inputs(153)));
    layer0_outputs(1737) <= (inputs(53)) or (inputs(125));
    layer0_outputs(1738) <= not((inputs(194)) or (inputs(180)));
    layer0_outputs(1739) <= (inputs(214)) and not (inputs(187));
    layer0_outputs(1740) <= not((inputs(184)) or (inputs(45)));
    layer0_outputs(1741) <= not((inputs(68)) xor (inputs(193)));
    layer0_outputs(1742) <= inputs(202);
    layer0_outputs(1743) <= (inputs(43)) xor (inputs(201));
    layer0_outputs(1744) <= (inputs(255)) and (inputs(247));
    layer0_outputs(1745) <= (inputs(169)) or (inputs(28));
    layer0_outputs(1746) <= inputs(105);
    layer0_outputs(1747) <= '0';
    layer0_outputs(1748) <= not(inputs(240)) or (inputs(183));
    layer0_outputs(1749) <= not(inputs(152));
    layer0_outputs(1750) <= not((inputs(185)) xor (inputs(16)));
    layer0_outputs(1751) <= not((inputs(149)) or (inputs(54)));
    layer0_outputs(1752) <= not(inputs(148)) or (inputs(41));
    layer0_outputs(1753) <= (inputs(149)) and not (inputs(6));
    layer0_outputs(1754) <= not(inputs(155)) or (inputs(15));
    layer0_outputs(1755) <= (inputs(134)) and not (inputs(105));
    layer0_outputs(1756) <= not(inputs(119));
    layer0_outputs(1757) <= (inputs(187)) and not (inputs(31));
    layer0_outputs(1758) <= not((inputs(241)) xor (inputs(152)));
    layer0_outputs(1759) <= not(inputs(121));
    layer0_outputs(1760) <= (inputs(0)) or (inputs(72));
    layer0_outputs(1761) <= not((inputs(205)) xor (inputs(219)));
    layer0_outputs(1762) <= not((inputs(3)) or (inputs(118)));
    layer0_outputs(1763) <= not((inputs(150)) xor (inputs(7)));
    layer0_outputs(1764) <= not((inputs(241)) or (inputs(120)));
    layer0_outputs(1765) <= not((inputs(134)) xor (inputs(193)));
    layer0_outputs(1766) <= not(inputs(188));
    layer0_outputs(1767) <= not(inputs(122)) or (inputs(13));
    layer0_outputs(1768) <= not(inputs(135));
    layer0_outputs(1769) <= (inputs(75)) and not (inputs(245));
    layer0_outputs(1770) <= not((inputs(238)) or (inputs(94)));
    layer0_outputs(1771) <= (inputs(128)) xor (inputs(34));
    layer0_outputs(1772) <= not((inputs(67)) xor (inputs(147)));
    layer0_outputs(1773) <= not(inputs(200));
    layer0_outputs(1774) <= '1';
    layer0_outputs(1775) <= not((inputs(146)) xor (inputs(163)));
    layer0_outputs(1776) <= not(inputs(58)) or (inputs(144));
    layer0_outputs(1777) <= (inputs(36)) xor (inputs(44));
    layer0_outputs(1778) <= not(inputs(71)) or (inputs(66));
    layer0_outputs(1779) <= (inputs(145)) and not (inputs(176));
    layer0_outputs(1780) <= (inputs(215)) and not (inputs(190));
    layer0_outputs(1781) <= inputs(180);
    layer0_outputs(1782) <= (inputs(99)) and not (inputs(255));
    layer0_outputs(1783) <= not((inputs(45)) xor (inputs(235)));
    layer0_outputs(1784) <= not((inputs(86)) xor (inputs(224)));
    layer0_outputs(1785) <= (inputs(95)) xor (inputs(138));
    layer0_outputs(1786) <= inputs(184);
    layer0_outputs(1787) <= (inputs(144)) and not (inputs(251));
    layer0_outputs(1788) <= not((inputs(138)) xor (inputs(65)));
    layer0_outputs(1789) <= not((inputs(38)) or (inputs(79)));
    layer0_outputs(1790) <= '1';
    layer0_outputs(1791) <= not(inputs(98));
    layer0_outputs(1792) <= not(inputs(136)) or (inputs(165));
    layer0_outputs(1793) <= (inputs(236)) xor (inputs(92));
    layer0_outputs(1794) <= not((inputs(221)) xor (inputs(84)));
    layer0_outputs(1795) <= not((inputs(127)) or (inputs(170)));
    layer0_outputs(1796) <= not((inputs(1)) or (inputs(194)));
    layer0_outputs(1797) <= (inputs(171)) or (inputs(54));
    layer0_outputs(1798) <= inputs(92);
    layer0_outputs(1799) <= not(inputs(60)) or (inputs(214));
    layer0_outputs(1800) <= not((inputs(80)) or (inputs(156)));
    layer0_outputs(1801) <= not(inputs(100)) or (inputs(223));
    layer0_outputs(1802) <= not(inputs(66));
    layer0_outputs(1803) <= (inputs(126)) and not (inputs(221));
    layer0_outputs(1804) <= not((inputs(123)) or (inputs(4)));
    layer0_outputs(1805) <= inputs(10);
    layer0_outputs(1806) <= not(inputs(137));
    layer0_outputs(1807) <= (inputs(13)) xor (inputs(239));
    layer0_outputs(1808) <= (inputs(29)) and not (inputs(166));
    layer0_outputs(1809) <= not((inputs(253)) xor (inputs(138)));
    layer0_outputs(1810) <= not((inputs(216)) or (inputs(43)));
    layer0_outputs(1811) <= not((inputs(237)) or (inputs(195)));
    layer0_outputs(1812) <= (inputs(196)) and not (inputs(249));
    layer0_outputs(1813) <= (inputs(47)) and not (inputs(248));
    layer0_outputs(1814) <= not(inputs(143)) or (inputs(244));
    layer0_outputs(1815) <= (inputs(18)) and not (inputs(6));
    layer0_outputs(1816) <= inputs(51);
    layer0_outputs(1817) <= (inputs(194)) and not (inputs(18));
    layer0_outputs(1818) <= not((inputs(81)) or (inputs(85)));
    layer0_outputs(1819) <= inputs(36);
    layer0_outputs(1820) <= not(inputs(92));
    layer0_outputs(1821) <= not(inputs(121));
    layer0_outputs(1822) <= not(inputs(217)) or (inputs(23));
    layer0_outputs(1823) <= inputs(82);
    layer0_outputs(1824) <= not((inputs(104)) or (inputs(250)));
    layer0_outputs(1825) <= not(inputs(46)) or (inputs(254));
    layer0_outputs(1826) <= not(inputs(122)) or (inputs(64));
    layer0_outputs(1827) <= not(inputs(235)) or (inputs(93));
    layer0_outputs(1828) <= not(inputs(151));
    layer0_outputs(1829) <= (inputs(82)) and not (inputs(230));
    layer0_outputs(1830) <= not(inputs(64));
    layer0_outputs(1831) <= not((inputs(81)) xor (inputs(216)));
    layer0_outputs(1832) <= not((inputs(25)) or (inputs(90)));
    layer0_outputs(1833) <= not((inputs(38)) xor (inputs(13)));
    layer0_outputs(1834) <= (inputs(180)) and not (inputs(141));
    layer0_outputs(1835) <= inputs(133);
    layer0_outputs(1836) <= not(inputs(163));
    layer0_outputs(1837) <= (inputs(188)) and not (inputs(28));
    layer0_outputs(1838) <= not(inputs(6));
    layer0_outputs(1839) <= not((inputs(230)) or (inputs(117)));
    layer0_outputs(1840) <= (inputs(188)) or (inputs(74));
    layer0_outputs(1841) <= inputs(100);
    layer0_outputs(1842) <= inputs(84);
    layer0_outputs(1843) <= not(inputs(199));
    layer0_outputs(1844) <= not(inputs(135)) or (inputs(154));
    layer0_outputs(1845) <= not(inputs(121));
    layer0_outputs(1846) <= not(inputs(168)) or (inputs(0));
    layer0_outputs(1847) <= inputs(220);
    layer0_outputs(1848) <= inputs(117);
    layer0_outputs(1849) <= inputs(123);
    layer0_outputs(1850) <= not(inputs(250)) or (inputs(190));
    layer0_outputs(1851) <= not((inputs(194)) or (inputs(79)));
    layer0_outputs(1852) <= (inputs(158)) xor (inputs(193));
    layer0_outputs(1853) <= inputs(163);
    layer0_outputs(1854) <= not((inputs(115)) xor (inputs(176)));
    layer0_outputs(1855) <= not((inputs(65)) or (inputs(84)));
    layer0_outputs(1856) <= not((inputs(176)) or (inputs(181)));
    layer0_outputs(1857) <= inputs(118);
    layer0_outputs(1858) <= (inputs(148)) and not (inputs(230));
    layer0_outputs(1859) <= not((inputs(113)) and (inputs(114)));
    layer0_outputs(1860) <= not(inputs(136)) or (inputs(247));
    layer0_outputs(1861) <= inputs(109);
    layer0_outputs(1862) <= not(inputs(54)) or (inputs(176));
    layer0_outputs(1863) <= not((inputs(172)) or (inputs(184)));
    layer0_outputs(1864) <= (inputs(55)) or (inputs(193));
    layer0_outputs(1865) <= not(inputs(232));
    layer0_outputs(1866) <= inputs(89);
    layer0_outputs(1867) <= not((inputs(32)) xor (inputs(102)));
    layer0_outputs(1868) <= not((inputs(163)) or (inputs(86)));
    layer0_outputs(1869) <= not(inputs(17)) or (inputs(204));
    layer0_outputs(1870) <= (inputs(149)) and not (inputs(12));
    layer0_outputs(1871) <= not(inputs(100)) or (inputs(164));
    layer0_outputs(1872) <= (inputs(16)) xor (inputs(69));
    layer0_outputs(1873) <= (inputs(93)) or (inputs(205));
    layer0_outputs(1874) <= (inputs(149)) and not (inputs(219));
    layer0_outputs(1875) <= inputs(165);
    layer0_outputs(1876) <= not((inputs(211)) xor (inputs(1)));
    layer0_outputs(1877) <= (inputs(114)) or (inputs(93));
    layer0_outputs(1878) <= inputs(146);
    layer0_outputs(1879) <= not(inputs(179)) or (inputs(41));
    layer0_outputs(1880) <= not(inputs(177)) or (inputs(189));
    layer0_outputs(1881) <= (inputs(189)) and not (inputs(222));
    layer0_outputs(1882) <= not(inputs(166)) or (inputs(110));
    layer0_outputs(1883) <= not(inputs(95)) or (inputs(45));
    layer0_outputs(1884) <= not((inputs(60)) or (inputs(48)));
    layer0_outputs(1885) <= (inputs(117)) and not (inputs(175));
    layer0_outputs(1886) <= (inputs(5)) or (inputs(44));
    layer0_outputs(1887) <= (inputs(56)) and (inputs(106));
    layer0_outputs(1888) <= (inputs(112)) or (inputs(192));
    layer0_outputs(1889) <= not(inputs(139)) or (inputs(8));
    layer0_outputs(1890) <= (inputs(255)) or (inputs(228));
    layer0_outputs(1891) <= (inputs(33)) or (inputs(136));
    layer0_outputs(1892) <= inputs(75);
    layer0_outputs(1893) <= not(inputs(12));
    layer0_outputs(1894) <= (inputs(86)) and not (inputs(158));
    layer0_outputs(1895) <= not((inputs(42)) or (inputs(191)));
    layer0_outputs(1896) <= (inputs(38)) or (inputs(36));
    layer0_outputs(1897) <= (inputs(233)) or (inputs(87));
    layer0_outputs(1898) <= not(inputs(45));
    layer0_outputs(1899) <= not((inputs(54)) or (inputs(94)));
    layer0_outputs(1900) <= (inputs(182)) or (inputs(122));
    layer0_outputs(1901) <= inputs(45);
    layer0_outputs(1902) <= not((inputs(203)) xor (inputs(170)));
    layer0_outputs(1903) <= (inputs(222)) and not (inputs(244));
    layer0_outputs(1904) <= inputs(181);
    layer0_outputs(1905) <= not(inputs(11));
    layer0_outputs(1906) <= (inputs(185)) and not (inputs(111));
    layer0_outputs(1907) <= not(inputs(85));
    layer0_outputs(1908) <= not(inputs(19));
    layer0_outputs(1909) <= (inputs(158)) or (inputs(152));
    layer0_outputs(1910) <= inputs(74);
    layer0_outputs(1911) <= not(inputs(60)) or (inputs(210));
    layer0_outputs(1912) <= not((inputs(90)) or (inputs(108)));
    layer0_outputs(1913) <= (inputs(106)) and (inputs(149));
    layer0_outputs(1914) <= not(inputs(86)) or (inputs(172));
    layer0_outputs(1915) <= not(inputs(148));
    layer0_outputs(1916) <= (inputs(251)) and (inputs(206));
    layer0_outputs(1917) <= (inputs(186)) and not (inputs(113));
    layer0_outputs(1918) <= not((inputs(201)) or (inputs(247)));
    layer0_outputs(1919) <= not(inputs(57));
    layer0_outputs(1920) <= (inputs(106)) and not (inputs(118));
    layer0_outputs(1921) <= not((inputs(197)) or (inputs(74)));
    layer0_outputs(1922) <= not((inputs(89)) or (inputs(9)));
    layer0_outputs(1923) <= (inputs(27)) and not (inputs(47));
    layer0_outputs(1924) <= not(inputs(250)) or (inputs(36));
    layer0_outputs(1925) <= not(inputs(252)) or (inputs(110));
    layer0_outputs(1926) <= not((inputs(156)) xor (inputs(205)));
    layer0_outputs(1927) <= (inputs(209)) and not (inputs(49));
    layer0_outputs(1928) <= (inputs(155)) and not (inputs(237));
    layer0_outputs(1929) <= not((inputs(33)) xor (inputs(134)));
    layer0_outputs(1930) <= not(inputs(221)) or (inputs(83));
    layer0_outputs(1931) <= inputs(64);
    layer0_outputs(1932) <= not((inputs(63)) xor (inputs(100)));
    layer0_outputs(1933) <= inputs(153);
    layer0_outputs(1934) <= not((inputs(70)) or (inputs(23)));
    layer0_outputs(1935) <= (inputs(106)) and not (inputs(156));
    layer0_outputs(1936) <= not(inputs(230)) or (inputs(33));
    layer0_outputs(1937) <= not(inputs(52));
    layer0_outputs(1938) <= (inputs(27)) or (inputs(170));
    layer0_outputs(1939) <= not((inputs(32)) or (inputs(53)));
    layer0_outputs(1940) <= (inputs(183)) and not (inputs(42));
    layer0_outputs(1941) <= not((inputs(21)) or (inputs(53)));
    layer0_outputs(1942) <= not(inputs(84));
    layer0_outputs(1943) <= not((inputs(39)) or (inputs(242)));
    layer0_outputs(1944) <= inputs(225);
    layer0_outputs(1945) <= inputs(109);
    layer0_outputs(1946) <= inputs(197);
    layer0_outputs(1947) <= (inputs(199)) and not (inputs(67));
    layer0_outputs(1948) <= not(inputs(163));
    layer0_outputs(1949) <= (inputs(250)) xor (inputs(251));
    layer0_outputs(1950) <= inputs(180);
    layer0_outputs(1951) <= not((inputs(236)) xor (inputs(187)));
    layer0_outputs(1952) <= not(inputs(216)) or (inputs(42));
    layer0_outputs(1953) <= not((inputs(251)) and (inputs(143)));
    layer0_outputs(1954) <= not(inputs(96));
    layer0_outputs(1955) <= not(inputs(145));
    layer0_outputs(1956) <= not((inputs(25)) or (inputs(106)));
    layer0_outputs(1957) <= not(inputs(56));
    layer0_outputs(1958) <= (inputs(79)) xor (inputs(232));
    layer0_outputs(1959) <= inputs(109);
    layer0_outputs(1960) <= not(inputs(73));
    layer0_outputs(1961) <= (inputs(66)) and not (inputs(15));
    layer0_outputs(1962) <= inputs(70);
    layer0_outputs(1963) <= '1';
    layer0_outputs(1964) <= not((inputs(241)) xor (inputs(98)));
    layer0_outputs(1965) <= not(inputs(150)) or (inputs(62));
    layer0_outputs(1966) <= (inputs(149)) or (inputs(27));
    layer0_outputs(1967) <= not((inputs(117)) or (inputs(239)));
    layer0_outputs(1968) <= inputs(254);
    layer0_outputs(1969) <= (inputs(90)) and not (inputs(238));
    layer0_outputs(1970) <= not(inputs(230));
    layer0_outputs(1971) <= not((inputs(43)) or (inputs(49)));
    layer0_outputs(1972) <= (inputs(88)) or (inputs(227));
    layer0_outputs(1973) <= not((inputs(2)) xor (inputs(244)));
    layer0_outputs(1974) <= (inputs(218)) xor (inputs(185));
    layer0_outputs(1975) <= inputs(171);
    layer0_outputs(1976) <= (inputs(198)) or (inputs(178));
    layer0_outputs(1977) <= not(inputs(193)) or (inputs(9));
    layer0_outputs(1978) <= (inputs(220)) and (inputs(141));
    layer0_outputs(1979) <= (inputs(193)) and (inputs(127));
    layer0_outputs(1980) <= (inputs(188)) xor (inputs(56));
    layer0_outputs(1981) <= not((inputs(94)) or (inputs(76)));
    layer0_outputs(1982) <= '1';
    layer0_outputs(1983) <= inputs(103);
    layer0_outputs(1984) <= (inputs(130)) or (inputs(137));
    layer0_outputs(1985) <= not(inputs(71));
    layer0_outputs(1986) <= (inputs(192)) or (inputs(238));
    layer0_outputs(1987) <= not((inputs(148)) xor (inputs(119)));
    layer0_outputs(1988) <= (inputs(95)) xor (inputs(177));
    layer0_outputs(1989) <= not((inputs(186)) or (inputs(224)));
    layer0_outputs(1990) <= not(inputs(243));
    layer0_outputs(1991) <= inputs(236);
    layer0_outputs(1992) <= not(inputs(141));
    layer0_outputs(1993) <= (inputs(9)) and (inputs(46));
    layer0_outputs(1994) <= not(inputs(96)) or (inputs(0));
    layer0_outputs(1995) <= not((inputs(78)) xor (inputs(151)));
    layer0_outputs(1996) <= not(inputs(216));
    layer0_outputs(1997) <= (inputs(252)) or (inputs(45));
    layer0_outputs(1998) <= not((inputs(200)) or (inputs(147)));
    layer0_outputs(1999) <= not(inputs(123)) or (inputs(176));
    layer0_outputs(2000) <= (inputs(181)) and (inputs(207));
    layer0_outputs(2001) <= '1';
    layer0_outputs(2002) <= not(inputs(77)) or (inputs(222));
    layer0_outputs(2003) <= not(inputs(164)) or (inputs(178));
    layer0_outputs(2004) <= inputs(201);
    layer0_outputs(2005) <= not((inputs(220)) or (inputs(57)));
    layer0_outputs(2006) <= not((inputs(254)) and (inputs(111)));
    layer0_outputs(2007) <= (inputs(97)) or (inputs(107));
    layer0_outputs(2008) <= not(inputs(108)) or (inputs(42));
    layer0_outputs(2009) <= not(inputs(203));
    layer0_outputs(2010) <= (inputs(55)) xor (inputs(42));
    layer0_outputs(2011) <= not(inputs(195));
    layer0_outputs(2012) <= (inputs(73)) and not (inputs(109));
    layer0_outputs(2013) <= (inputs(96)) or (inputs(186));
    layer0_outputs(2014) <= (inputs(132)) or (inputs(133));
    layer0_outputs(2015) <= (inputs(179)) and (inputs(13));
    layer0_outputs(2016) <= inputs(125);
    layer0_outputs(2017) <= not(inputs(56));
    layer0_outputs(2018) <= not((inputs(131)) xor (inputs(51)));
    layer0_outputs(2019) <= not((inputs(82)) xor (inputs(29)));
    layer0_outputs(2020) <= not((inputs(100)) and (inputs(78)));
    layer0_outputs(2021) <= not((inputs(4)) or (inputs(118)));
    layer0_outputs(2022) <= not((inputs(100)) xor (inputs(176)));
    layer0_outputs(2023) <= not((inputs(171)) or (inputs(22)));
    layer0_outputs(2024) <= (inputs(243)) or (inputs(72));
    layer0_outputs(2025) <= '0';
    layer0_outputs(2026) <= not(inputs(222)) or (inputs(45));
    layer0_outputs(2027) <= inputs(137);
    layer0_outputs(2028) <= '0';
    layer0_outputs(2029) <= inputs(240);
    layer0_outputs(2030) <= not(inputs(109));
    layer0_outputs(2031) <= not(inputs(164));
    layer0_outputs(2032) <= inputs(191);
    layer0_outputs(2033) <= not(inputs(162)) or (inputs(218));
    layer0_outputs(2034) <= '0';
    layer0_outputs(2035) <= not(inputs(24)) or (inputs(0));
    layer0_outputs(2036) <= not(inputs(107));
    layer0_outputs(2037) <= not(inputs(254)) or (inputs(50));
    layer0_outputs(2038) <= (inputs(233)) or (inputs(47));
    layer0_outputs(2039) <= not((inputs(86)) or (inputs(4)));
    layer0_outputs(2040) <= (inputs(120)) and not (inputs(189));
    layer0_outputs(2041) <= not(inputs(119));
    layer0_outputs(2042) <= inputs(73);
    layer0_outputs(2043) <= not((inputs(58)) xor (inputs(123)));
    layer0_outputs(2044) <= (inputs(187)) or (inputs(34));
    layer0_outputs(2045) <= '0';
    layer0_outputs(2046) <= (inputs(95)) or (inputs(135));
    layer0_outputs(2047) <= not(inputs(234)) or (inputs(98));
    layer0_outputs(2048) <= (inputs(86)) and not (inputs(52));
    layer0_outputs(2049) <= (inputs(81)) xor (inputs(233));
    layer0_outputs(2050) <= not(inputs(229)) or (inputs(242));
    layer0_outputs(2051) <= inputs(85);
    layer0_outputs(2052) <= not(inputs(132)) or (inputs(22));
    layer0_outputs(2053) <= inputs(215);
    layer0_outputs(2054) <= not((inputs(220)) or (inputs(116)));
    layer0_outputs(2055) <= (inputs(131)) and not (inputs(18));
    layer0_outputs(2056) <= (inputs(147)) or (inputs(178));
    layer0_outputs(2057) <= not(inputs(93)) or (inputs(13));
    layer0_outputs(2058) <= not((inputs(56)) or (inputs(47)));
    layer0_outputs(2059) <= inputs(149);
    layer0_outputs(2060) <= not((inputs(203)) or (inputs(144)));
    layer0_outputs(2061) <= not((inputs(96)) or (inputs(132)));
    layer0_outputs(2062) <= (inputs(2)) xor (inputs(225));
    layer0_outputs(2063) <= (inputs(135)) and not (inputs(225));
    layer0_outputs(2064) <= not((inputs(154)) or (inputs(4)));
    layer0_outputs(2065) <= not((inputs(73)) or (inputs(180)));
    layer0_outputs(2066) <= (inputs(35)) or (inputs(172));
    layer0_outputs(2067) <= (inputs(86)) and not (inputs(4));
    layer0_outputs(2068) <= not(inputs(136)) or (inputs(187));
    layer0_outputs(2069) <= not((inputs(84)) or (inputs(144)));
    layer0_outputs(2070) <= '0';
    layer0_outputs(2071) <= (inputs(202)) or (inputs(240));
    layer0_outputs(2072) <= not((inputs(159)) or (inputs(163)));
    layer0_outputs(2073) <= not(inputs(120)) or (inputs(39));
    layer0_outputs(2074) <= not(inputs(161)) or (inputs(67));
    layer0_outputs(2075) <= (inputs(165)) or (inputs(157));
    layer0_outputs(2076) <= not(inputs(151)) or (inputs(95));
    layer0_outputs(2077) <= not(inputs(12));
    layer0_outputs(2078) <= (inputs(163)) xor (inputs(202));
    layer0_outputs(2079) <= not((inputs(30)) or (inputs(213)));
    layer0_outputs(2080) <= not((inputs(255)) or (inputs(210)));
    layer0_outputs(2081) <= not((inputs(100)) or (inputs(61)));
    layer0_outputs(2082) <= (inputs(195)) xor (inputs(169));
    layer0_outputs(2083) <= (inputs(4)) and not (inputs(66));
    layer0_outputs(2084) <= inputs(43);
    layer0_outputs(2085) <= not(inputs(131)) or (inputs(222));
    layer0_outputs(2086) <= (inputs(58)) and not (inputs(242));
    layer0_outputs(2087) <= not(inputs(185));
    layer0_outputs(2088) <= not((inputs(133)) xor (inputs(142)));
    layer0_outputs(2089) <= not(inputs(181));
    layer0_outputs(2090) <= (inputs(164)) xor (inputs(25));
    layer0_outputs(2091) <= not((inputs(245)) xor (inputs(72)));
    layer0_outputs(2092) <= inputs(38);
    layer0_outputs(2093) <= inputs(238);
    layer0_outputs(2094) <= not((inputs(92)) xor (inputs(18)));
    layer0_outputs(2095) <= not(inputs(123));
    layer0_outputs(2096) <= not(inputs(75)) or (inputs(223));
    layer0_outputs(2097) <= not(inputs(187));
    layer0_outputs(2098) <= not(inputs(134));
    layer0_outputs(2099) <= (inputs(41)) or (inputs(77));
    layer0_outputs(2100) <= inputs(161);
    layer0_outputs(2101) <= (inputs(157)) or (inputs(118));
    layer0_outputs(2102) <= (inputs(128)) xor (inputs(46));
    layer0_outputs(2103) <= (inputs(61)) or (inputs(183));
    layer0_outputs(2104) <= inputs(45);
    layer0_outputs(2105) <= (inputs(9)) xor (inputs(38));
    layer0_outputs(2106) <= inputs(139);
    layer0_outputs(2107) <= not(inputs(138));
    layer0_outputs(2108) <= not((inputs(141)) and (inputs(234)));
    layer0_outputs(2109) <= '0';
    layer0_outputs(2110) <= '0';
    layer0_outputs(2111) <= '0';
    layer0_outputs(2112) <= not((inputs(237)) xor (inputs(129)));
    layer0_outputs(2113) <= not(inputs(73));
    layer0_outputs(2114) <= '0';
    layer0_outputs(2115) <= not(inputs(92));
    layer0_outputs(2116) <= not((inputs(251)) xor (inputs(254)));
    layer0_outputs(2117) <= not(inputs(147)) or (inputs(39));
    layer0_outputs(2118) <= inputs(57);
    layer0_outputs(2119) <= (inputs(87)) and not (inputs(195));
    layer0_outputs(2120) <= (inputs(52)) or (inputs(12));
    layer0_outputs(2121) <= (inputs(40)) and not (inputs(112));
    layer0_outputs(2122) <= not(inputs(234)) or (inputs(189));
    layer0_outputs(2123) <= not(inputs(182));
    layer0_outputs(2124) <= (inputs(147)) and not (inputs(239));
    layer0_outputs(2125) <= (inputs(186)) xor (inputs(111));
    layer0_outputs(2126) <= '1';
    layer0_outputs(2127) <= (inputs(31)) and (inputs(72));
    layer0_outputs(2128) <= not(inputs(138)) or (inputs(22));
    layer0_outputs(2129) <= (inputs(229)) xor (inputs(6));
    layer0_outputs(2130) <= (inputs(97)) and not (inputs(179));
    layer0_outputs(2131) <= (inputs(102)) xor (inputs(223));
    layer0_outputs(2132) <= not((inputs(72)) or (inputs(163)));
    layer0_outputs(2133) <= (inputs(118)) or (inputs(173));
    layer0_outputs(2134) <= (inputs(201)) and not (inputs(105));
    layer0_outputs(2135) <= not((inputs(172)) xor (inputs(177)));
    layer0_outputs(2136) <= not((inputs(82)) or (inputs(99)));
    layer0_outputs(2137) <= '0';
    layer0_outputs(2138) <= not((inputs(204)) xor (inputs(63)));
    layer0_outputs(2139) <= (inputs(31)) and not (inputs(43));
    layer0_outputs(2140) <= (inputs(50)) and (inputs(65));
    layer0_outputs(2141) <= (inputs(26)) xor (inputs(50));
    layer0_outputs(2142) <= (inputs(87)) xor (inputs(218));
    layer0_outputs(2143) <= (inputs(189)) xor (inputs(123));
    layer0_outputs(2144) <= not((inputs(171)) or (inputs(74)));
    layer0_outputs(2145) <= not((inputs(90)) or (inputs(142)));
    layer0_outputs(2146) <= (inputs(78)) xor (inputs(155));
    layer0_outputs(2147) <= (inputs(101)) xor (inputs(221));
    layer0_outputs(2148) <= not(inputs(251)) or (inputs(255));
    layer0_outputs(2149) <= (inputs(249)) and (inputs(50));
    layer0_outputs(2150) <= (inputs(243)) xor (inputs(163));
    layer0_outputs(2151) <= inputs(61);
    layer0_outputs(2152) <= not(inputs(199)) or (inputs(241));
    layer0_outputs(2153) <= (inputs(24)) and (inputs(80));
    layer0_outputs(2154) <= not((inputs(158)) or (inputs(171)));
    layer0_outputs(2155) <= not(inputs(113)) or (inputs(143));
    layer0_outputs(2156) <= inputs(122);
    layer0_outputs(2157) <= inputs(152);
    layer0_outputs(2158) <= (inputs(246)) and not (inputs(1));
    layer0_outputs(2159) <= not((inputs(125)) or (inputs(50)));
    layer0_outputs(2160) <= (inputs(176)) xor (inputs(108));
    layer0_outputs(2161) <= (inputs(119)) xor (inputs(145));
    layer0_outputs(2162) <= (inputs(9)) and (inputs(121));
    layer0_outputs(2163) <= not(inputs(201));
    layer0_outputs(2164) <= (inputs(71)) or (inputs(94));
    layer0_outputs(2165) <= (inputs(218)) and not (inputs(248));
    layer0_outputs(2166) <= not(inputs(149));
    layer0_outputs(2167) <= not(inputs(55));
    layer0_outputs(2168) <= (inputs(72)) and (inputs(121));
    layer0_outputs(2169) <= (inputs(57)) xor (inputs(177));
    layer0_outputs(2170) <= '1';
    layer0_outputs(2171) <= '0';
    layer0_outputs(2172) <= (inputs(147)) or (inputs(167));
    layer0_outputs(2173) <= not(inputs(26)) or (inputs(2));
    layer0_outputs(2174) <= not(inputs(233)) or (inputs(189));
    layer0_outputs(2175) <= not(inputs(69));
    layer0_outputs(2176) <= inputs(255);
    layer0_outputs(2177) <= (inputs(179)) or (inputs(39));
    layer0_outputs(2178) <= not((inputs(16)) xor (inputs(101)));
    layer0_outputs(2179) <= inputs(253);
    layer0_outputs(2180) <= (inputs(181)) xor (inputs(241));
    layer0_outputs(2181) <= not(inputs(87)) or (inputs(125));
    layer0_outputs(2182) <= (inputs(112)) xor (inputs(172));
    layer0_outputs(2183) <= (inputs(251)) or (inputs(120));
    layer0_outputs(2184) <= inputs(164);
    layer0_outputs(2185) <= not((inputs(198)) or (inputs(39)));
    layer0_outputs(2186) <= (inputs(188)) xor (inputs(117));
    layer0_outputs(2187) <= not((inputs(208)) and (inputs(255)));
    layer0_outputs(2188) <= (inputs(183)) and not (inputs(229));
    layer0_outputs(2189) <= (inputs(48)) and not (inputs(127));
    layer0_outputs(2190) <= (inputs(121)) and not (inputs(120));
    layer0_outputs(2191) <= (inputs(247)) or (inputs(149));
    layer0_outputs(2192) <= not(inputs(167));
    layer0_outputs(2193) <= not((inputs(77)) xor (inputs(237)));
    layer0_outputs(2194) <= not(inputs(148));
    layer0_outputs(2195) <= '1';
    layer0_outputs(2196) <= (inputs(20)) and not (inputs(98));
    layer0_outputs(2197) <= inputs(152);
    layer0_outputs(2198) <= not((inputs(87)) and (inputs(201)));
    layer0_outputs(2199) <= not((inputs(36)) and (inputs(23)));
    layer0_outputs(2200) <= (inputs(209)) and not (inputs(14));
    layer0_outputs(2201) <= (inputs(95)) xor (inputs(215));
    layer0_outputs(2202) <= (inputs(27)) or (inputs(99));
    layer0_outputs(2203) <= not((inputs(231)) or (inputs(191)));
    layer0_outputs(2204) <= not(inputs(56));
    layer0_outputs(2205) <= not(inputs(43));
    layer0_outputs(2206) <= not((inputs(149)) or (inputs(168)));
    layer0_outputs(2207) <= not(inputs(102)) or (inputs(233));
    layer0_outputs(2208) <= not((inputs(213)) or (inputs(66)));
    layer0_outputs(2209) <= (inputs(114)) and (inputs(217));
    layer0_outputs(2210) <= (inputs(93)) and not (inputs(160));
    layer0_outputs(2211) <= (inputs(182)) xor (inputs(33));
    layer0_outputs(2212) <= (inputs(74)) and not (inputs(128));
    layer0_outputs(2213) <= (inputs(99)) or (inputs(220));
    layer0_outputs(2214) <= inputs(196);
    layer0_outputs(2215) <= (inputs(29)) and (inputs(204));
    layer0_outputs(2216) <= not(inputs(168)) or (inputs(207));
    layer0_outputs(2217) <= (inputs(146)) or (inputs(91));
    layer0_outputs(2218) <= (inputs(95)) and (inputs(46));
    layer0_outputs(2219) <= not(inputs(143));
    layer0_outputs(2220) <= (inputs(213)) or (inputs(93));
    layer0_outputs(2221) <= (inputs(255)) xor (inputs(32));
    layer0_outputs(2222) <= not((inputs(236)) xor (inputs(156)));
    layer0_outputs(2223) <= not(inputs(89));
    layer0_outputs(2224) <= (inputs(171)) xor (inputs(67));
    layer0_outputs(2225) <= not(inputs(233)) or (inputs(175));
    layer0_outputs(2226) <= inputs(153);
    layer0_outputs(2227) <= not(inputs(197));
    layer0_outputs(2228) <= not((inputs(119)) and (inputs(108)));
    layer0_outputs(2229) <= (inputs(101)) and not (inputs(160));
    layer0_outputs(2230) <= '1';
    layer0_outputs(2231) <= not((inputs(172)) xor (inputs(81)));
    layer0_outputs(2232) <= not((inputs(147)) or (inputs(191)));
    layer0_outputs(2233) <= not(inputs(164)) or (inputs(248));
    layer0_outputs(2234) <= not(inputs(55));
    layer0_outputs(2235) <= not(inputs(135));
    layer0_outputs(2236) <= not(inputs(154));
    layer0_outputs(2237) <= (inputs(163)) and not (inputs(20));
    layer0_outputs(2238) <= inputs(163);
    layer0_outputs(2239) <= (inputs(75)) or (inputs(73));
    layer0_outputs(2240) <= not((inputs(253)) or (inputs(121)));
    layer0_outputs(2241) <= (inputs(182)) and not (inputs(111));
    layer0_outputs(2242) <= (inputs(18)) and not (inputs(63));
    layer0_outputs(2243) <= '1';
    layer0_outputs(2244) <= not(inputs(106));
    layer0_outputs(2245) <= not(inputs(69)) or (inputs(224));
    layer0_outputs(2246) <= not((inputs(178)) xor (inputs(53)));
    layer0_outputs(2247) <= (inputs(140)) or (inputs(5));
    layer0_outputs(2248) <= (inputs(61)) xor (inputs(54));
    layer0_outputs(2249) <= (inputs(230)) and not (inputs(175));
    layer0_outputs(2250) <= not((inputs(196)) xor (inputs(126)));
    layer0_outputs(2251) <= not((inputs(6)) xor (inputs(21)));
    layer0_outputs(2252) <= (inputs(0)) and not (inputs(251));
    layer0_outputs(2253) <= not(inputs(164));
    layer0_outputs(2254) <= (inputs(254)) or (inputs(186));
    layer0_outputs(2255) <= not(inputs(114)) or (inputs(7));
    layer0_outputs(2256) <= not(inputs(89)) or (inputs(189));
    layer0_outputs(2257) <= not(inputs(173)) or (inputs(92));
    layer0_outputs(2258) <= inputs(3);
    layer0_outputs(2259) <= not((inputs(183)) xor (inputs(232)));
    layer0_outputs(2260) <= not((inputs(26)) or (inputs(214)));
    layer0_outputs(2261) <= (inputs(4)) and (inputs(101));
    layer0_outputs(2262) <= (inputs(33)) and not (inputs(33));
    layer0_outputs(2263) <= not((inputs(102)) xor (inputs(98)));
    layer0_outputs(2264) <= not((inputs(83)) xor (inputs(70)));
    layer0_outputs(2265) <= (inputs(135)) and not (inputs(78));
    layer0_outputs(2266) <= not(inputs(200)) or (inputs(205));
    layer0_outputs(2267) <= (inputs(185)) xor (inputs(158));
    layer0_outputs(2268) <= not(inputs(106));
    layer0_outputs(2269) <= (inputs(249)) or (inputs(29));
    layer0_outputs(2270) <= inputs(58);
    layer0_outputs(2271) <= (inputs(31)) or (inputs(63));
    layer0_outputs(2272) <= (inputs(136)) and not (inputs(28));
    layer0_outputs(2273) <= (inputs(232)) or (inputs(161));
    layer0_outputs(2274) <= not(inputs(196));
    layer0_outputs(2275) <= not(inputs(63));
    layer0_outputs(2276) <= not(inputs(120)) or (inputs(158));
    layer0_outputs(2277) <= not((inputs(122)) xor (inputs(224)));
    layer0_outputs(2278) <= (inputs(133)) and not (inputs(92));
    layer0_outputs(2279) <= (inputs(108)) and not (inputs(194));
    layer0_outputs(2280) <= (inputs(193)) or (inputs(175));
    layer0_outputs(2281) <= (inputs(171)) or (inputs(234));
    layer0_outputs(2282) <= (inputs(143)) xor (inputs(69));
    layer0_outputs(2283) <= not((inputs(196)) xor (inputs(220)));
    layer0_outputs(2284) <= not((inputs(110)) and (inputs(58)));
    layer0_outputs(2285) <= not(inputs(169));
    layer0_outputs(2286) <= (inputs(167)) and not (inputs(64));
    layer0_outputs(2287) <= not((inputs(225)) xor (inputs(197)));
    layer0_outputs(2288) <= (inputs(106)) and not (inputs(110));
    layer0_outputs(2289) <= (inputs(48)) and not (inputs(30));
    layer0_outputs(2290) <= (inputs(53)) and not (inputs(44));
    layer0_outputs(2291) <= not(inputs(70));
    layer0_outputs(2292) <= not((inputs(214)) or (inputs(76)));
    layer0_outputs(2293) <= (inputs(155)) xor (inputs(33));
    layer0_outputs(2294) <= (inputs(213)) and not (inputs(97));
    layer0_outputs(2295) <= (inputs(115)) and not (inputs(209));
    layer0_outputs(2296) <= not((inputs(15)) xor (inputs(226)));
    layer0_outputs(2297) <= not(inputs(58));
    layer0_outputs(2298) <= not(inputs(73)) or (inputs(175));
    layer0_outputs(2299) <= not((inputs(149)) and (inputs(171)));
    layer0_outputs(2300) <= inputs(69);
    layer0_outputs(2301) <= not((inputs(21)) xor (inputs(179)));
    layer0_outputs(2302) <= not((inputs(34)) or (inputs(229)));
    layer0_outputs(2303) <= (inputs(183)) and not (inputs(10));
    layer0_outputs(2304) <= (inputs(251)) or (inputs(58));
    layer0_outputs(2305) <= not((inputs(178)) xor (inputs(244)));
    layer0_outputs(2306) <= (inputs(103)) or (inputs(124));
    layer0_outputs(2307) <= not((inputs(187)) or (inputs(93)));
    layer0_outputs(2308) <= inputs(107);
    layer0_outputs(2309) <= not(inputs(121));
    layer0_outputs(2310) <= '1';
    layer0_outputs(2311) <= (inputs(137)) or (inputs(182));
    layer0_outputs(2312) <= (inputs(235)) and not (inputs(50));
    layer0_outputs(2313) <= inputs(43);
    layer0_outputs(2314) <= (inputs(65)) and (inputs(50));
    layer0_outputs(2315) <= not((inputs(224)) xor (inputs(232)));
    layer0_outputs(2316) <= '1';
    layer0_outputs(2317) <= inputs(181);
    layer0_outputs(2318) <= not(inputs(225));
    layer0_outputs(2319) <= (inputs(170)) and not (inputs(85));
    layer0_outputs(2320) <= not((inputs(34)) xor (inputs(255)));
    layer0_outputs(2321) <= '1';
    layer0_outputs(2322) <= not(inputs(152)) or (inputs(94));
    layer0_outputs(2323) <= inputs(52);
    layer0_outputs(2324) <= (inputs(3)) xor (inputs(14));
    layer0_outputs(2325) <= (inputs(153)) or (inputs(104));
    layer0_outputs(2326) <= not((inputs(174)) xor (inputs(88)));
    layer0_outputs(2327) <= (inputs(97)) or (inputs(84));
    layer0_outputs(2328) <= inputs(147);
    layer0_outputs(2329) <= inputs(151);
    layer0_outputs(2330) <= (inputs(110)) and (inputs(133));
    layer0_outputs(2331) <= (inputs(155)) and not (inputs(51));
    layer0_outputs(2332) <= inputs(100);
    layer0_outputs(2333) <= not(inputs(227)) or (inputs(15));
    layer0_outputs(2334) <= not((inputs(47)) or (inputs(182)));
    layer0_outputs(2335) <= not((inputs(5)) xor (inputs(172)));
    layer0_outputs(2336) <= inputs(136);
    layer0_outputs(2337) <= (inputs(36)) and not (inputs(82));
    layer0_outputs(2338) <= not(inputs(94));
    layer0_outputs(2339) <= not(inputs(0)) or (inputs(89));
    layer0_outputs(2340) <= not(inputs(109));
    layer0_outputs(2341) <= not(inputs(71)) or (inputs(60));
    layer0_outputs(2342) <= (inputs(101)) or (inputs(61));
    layer0_outputs(2343) <= not((inputs(22)) and (inputs(198)));
    layer0_outputs(2344) <= not((inputs(215)) or (inputs(175)));
    layer0_outputs(2345) <= (inputs(237)) xor (inputs(53));
    layer0_outputs(2346) <= (inputs(92)) or (inputs(49));
    layer0_outputs(2347) <= (inputs(120)) and not (inputs(187));
    layer0_outputs(2348) <= not(inputs(11)) or (inputs(47));
    layer0_outputs(2349) <= (inputs(179)) xor (inputs(216));
    layer0_outputs(2350) <= (inputs(231)) or (inputs(209));
    layer0_outputs(2351) <= (inputs(229)) or (inputs(184));
    layer0_outputs(2352) <= (inputs(17)) and (inputs(146));
    layer0_outputs(2353) <= not(inputs(45));
    layer0_outputs(2354) <= '0';
    layer0_outputs(2355) <= inputs(105);
    layer0_outputs(2356) <= not(inputs(142)) or (inputs(161));
    layer0_outputs(2357) <= (inputs(14)) or (inputs(202));
    layer0_outputs(2358) <= inputs(186);
    layer0_outputs(2359) <= '1';
    layer0_outputs(2360) <= not((inputs(35)) and (inputs(20)));
    layer0_outputs(2361) <= not((inputs(17)) or (inputs(24)));
    layer0_outputs(2362) <= not(inputs(58));
    layer0_outputs(2363) <= inputs(168);
    layer0_outputs(2364) <= inputs(132);
    layer0_outputs(2365) <= not((inputs(37)) xor (inputs(178)));
    layer0_outputs(2366) <= (inputs(43)) or (inputs(184));
    layer0_outputs(2367) <= inputs(125);
    layer0_outputs(2368) <= (inputs(2)) or (inputs(145));
    layer0_outputs(2369) <= not((inputs(92)) xor (inputs(168)));
    layer0_outputs(2370) <= inputs(13);
    layer0_outputs(2371) <= not(inputs(90));
    layer0_outputs(2372) <= not(inputs(134)) or (inputs(98));
    layer0_outputs(2373) <= (inputs(207)) or (inputs(166));
    layer0_outputs(2374) <= not(inputs(181));
    layer0_outputs(2375) <= (inputs(68)) or (inputs(107));
    layer0_outputs(2376) <= (inputs(98)) and not (inputs(110));
    layer0_outputs(2377) <= not(inputs(234)) or (inputs(83));
    layer0_outputs(2378) <= not(inputs(56));
    layer0_outputs(2379) <= not(inputs(114)) or (inputs(51));
    layer0_outputs(2380) <= '1';
    layer0_outputs(2381) <= not(inputs(218)) or (inputs(109));
    layer0_outputs(2382) <= (inputs(195)) or (inputs(74));
    layer0_outputs(2383) <= not(inputs(181));
    layer0_outputs(2384) <= not(inputs(54));
    layer0_outputs(2385) <= not((inputs(131)) xor (inputs(61)));
    layer0_outputs(2386) <= (inputs(29)) or (inputs(197));
    layer0_outputs(2387) <= inputs(73);
    layer0_outputs(2388) <= '1';
    layer0_outputs(2389) <= not(inputs(114));
    layer0_outputs(2390) <= not(inputs(119)) or (inputs(234));
    layer0_outputs(2391) <= not(inputs(251)) or (inputs(59));
    layer0_outputs(2392) <= not((inputs(228)) or (inputs(249)));
    layer0_outputs(2393) <= not((inputs(146)) or (inputs(143)));
    layer0_outputs(2394) <= (inputs(140)) or (inputs(103));
    layer0_outputs(2395) <= not(inputs(148));
    layer0_outputs(2396) <= inputs(157);
    layer0_outputs(2397) <= inputs(0);
    layer0_outputs(2398) <= not(inputs(197)) or (inputs(77));
    layer0_outputs(2399) <= not(inputs(185)) or (inputs(1));
    layer0_outputs(2400) <= (inputs(216)) xor (inputs(217));
    layer0_outputs(2401) <= not(inputs(161));
    layer0_outputs(2402) <= not(inputs(199));
    layer0_outputs(2403) <= inputs(53);
    layer0_outputs(2404) <= not((inputs(249)) or (inputs(1)));
    layer0_outputs(2405) <= not(inputs(155)) or (inputs(3));
    layer0_outputs(2406) <= not((inputs(167)) and (inputs(183)));
    layer0_outputs(2407) <= not(inputs(147));
    layer0_outputs(2408) <= (inputs(77)) or (inputs(120));
    layer0_outputs(2409) <= not(inputs(217));
    layer0_outputs(2410) <= (inputs(156)) or (inputs(191));
    layer0_outputs(2411) <= not((inputs(208)) and (inputs(210)));
    layer0_outputs(2412) <= inputs(22);
    layer0_outputs(2413) <= (inputs(90)) and not (inputs(221));
    layer0_outputs(2414) <= not(inputs(169)) or (inputs(58));
    layer0_outputs(2415) <= inputs(13);
    layer0_outputs(2416) <= not(inputs(238));
    layer0_outputs(2417) <= not(inputs(69));
    layer0_outputs(2418) <= (inputs(105)) and not (inputs(110));
    layer0_outputs(2419) <= inputs(165);
    layer0_outputs(2420) <= (inputs(10)) and not (inputs(219));
    layer0_outputs(2421) <= not((inputs(166)) xor (inputs(217)));
    layer0_outputs(2422) <= not((inputs(90)) and (inputs(151)));
    layer0_outputs(2423) <= '0';
    layer0_outputs(2424) <= not(inputs(57)) or (inputs(228));
    layer0_outputs(2425) <= not((inputs(53)) xor (inputs(189)));
    layer0_outputs(2426) <= (inputs(193)) or (inputs(69));
    layer0_outputs(2427) <= not((inputs(71)) xor (inputs(229)));
    layer0_outputs(2428) <= (inputs(20)) and not (inputs(127));
    layer0_outputs(2429) <= not((inputs(79)) xor (inputs(76)));
    layer0_outputs(2430) <= not(inputs(89)) or (inputs(112));
    layer0_outputs(2431) <= not((inputs(156)) or (inputs(163)));
    layer0_outputs(2432) <= (inputs(17)) and not (inputs(141));
    layer0_outputs(2433) <= not(inputs(165)) or (inputs(17));
    layer0_outputs(2434) <= (inputs(211)) xor (inputs(23));
    layer0_outputs(2435) <= (inputs(223)) or (inputs(74));
    layer0_outputs(2436) <= not((inputs(248)) xor (inputs(169)));
    layer0_outputs(2437) <= not((inputs(33)) xor (inputs(12)));
    layer0_outputs(2438) <= (inputs(92)) xor (inputs(61));
    layer0_outputs(2439) <= not((inputs(221)) or (inputs(158)));
    layer0_outputs(2440) <= (inputs(106)) and not (inputs(49));
    layer0_outputs(2441) <= not((inputs(148)) xor (inputs(138)));
    layer0_outputs(2442) <= not((inputs(136)) and (inputs(171)));
    layer0_outputs(2443) <= (inputs(115)) and not (inputs(225));
    layer0_outputs(2444) <= (inputs(124)) xor (inputs(88));
    layer0_outputs(2445) <= not((inputs(190)) xor (inputs(178)));
    layer0_outputs(2446) <= not(inputs(230));
    layer0_outputs(2447) <= not((inputs(122)) or (inputs(119)));
    layer0_outputs(2448) <= (inputs(40)) or (inputs(55));
    layer0_outputs(2449) <= (inputs(42)) or (inputs(133));
    layer0_outputs(2450) <= not(inputs(59));
    layer0_outputs(2451) <= not(inputs(201)) or (inputs(67));
    layer0_outputs(2452) <= not(inputs(92));
    layer0_outputs(2453) <= (inputs(54)) or (inputs(232));
    layer0_outputs(2454) <= not(inputs(158));
    layer0_outputs(2455) <= (inputs(105)) xor (inputs(97));
    layer0_outputs(2456) <= not(inputs(188));
    layer0_outputs(2457) <= not((inputs(80)) and (inputs(203)));
    layer0_outputs(2458) <= (inputs(99)) xor (inputs(188));
    layer0_outputs(2459) <= (inputs(227)) and not (inputs(13));
    layer0_outputs(2460) <= inputs(235);
    layer0_outputs(2461) <= inputs(200);
    layer0_outputs(2462) <= not(inputs(68)) or (inputs(161));
    layer0_outputs(2463) <= not((inputs(6)) xor (inputs(3)));
    layer0_outputs(2464) <= (inputs(8)) and (inputs(204));
    layer0_outputs(2465) <= not(inputs(150));
    layer0_outputs(2466) <= inputs(14);
    layer0_outputs(2467) <= not((inputs(173)) xor (inputs(27)));
    layer0_outputs(2468) <= not(inputs(152)) or (inputs(157));
    layer0_outputs(2469) <= not((inputs(70)) or (inputs(200)));
    layer0_outputs(2470) <= not((inputs(208)) or (inputs(152)));
    layer0_outputs(2471) <= not((inputs(54)) or (inputs(52)));
    layer0_outputs(2472) <= inputs(102);
    layer0_outputs(2473) <= inputs(71);
    layer0_outputs(2474) <= not(inputs(136)) or (inputs(60));
    layer0_outputs(2475) <= not(inputs(152)) or (inputs(249));
    layer0_outputs(2476) <= (inputs(244)) xor (inputs(27));
    layer0_outputs(2477) <= inputs(73);
    layer0_outputs(2478) <= not(inputs(49));
    layer0_outputs(2479) <= '1';
    layer0_outputs(2480) <= not((inputs(53)) xor (inputs(166)));
    layer0_outputs(2481) <= (inputs(41)) or (inputs(35));
    layer0_outputs(2482) <= not(inputs(3));
    layer0_outputs(2483) <= inputs(90);
    layer0_outputs(2484) <= not(inputs(96)) or (inputs(37));
    layer0_outputs(2485) <= not(inputs(76));
    layer0_outputs(2486) <= (inputs(73)) and (inputs(73));
    layer0_outputs(2487) <= not(inputs(171)) or (inputs(19));
    layer0_outputs(2488) <= not((inputs(31)) or (inputs(58)));
    layer0_outputs(2489) <= not(inputs(150));
    layer0_outputs(2490) <= (inputs(30)) or (inputs(86));
    layer0_outputs(2491) <= not((inputs(191)) xor (inputs(131)));
    layer0_outputs(2492) <= (inputs(105)) and not (inputs(183));
    layer0_outputs(2493) <= not((inputs(197)) or (inputs(37)));
    layer0_outputs(2494) <= not(inputs(16));
    layer0_outputs(2495) <= inputs(104);
    layer0_outputs(2496) <= inputs(80);
    layer0_outputs(2497) <= not((inputs(234)) xor (inputs(9)));
    layer0_outputs(2498) <= (inputs(179)) and not (inputs(78));
    layer0_outputs(2499) <= inputs(13);
    layer0_outputs(2500) <= (inputs(188)) or (inputs(97));
    layer0_outputs(2501) <= not(inputs(117));
    layer0_outputs(2502) <= (inputs(79)) or (inputs(23));
    layer0_outputs(2503) <= not((inputs(172)) and (inputs(66)));
    layer0_outputs(2504) <= not((inputs(40)) xor (inputs(4)));
    layer0_outputs(2505) <= not((inputs(41)) xor (inputs(23)));
    layer0_outputs(2506) <= inputs(98);
    layer0_outputs(2507) <= inputs(151);
    layer0_outputs(2508) <= (inputs(206)) xor (inputs(187));
    layer0_outputs(2509) <= '0';
    layer0_outputs(2510) <= inputs(243);
    layer0_outputs(2511) <= not((inputs(204)) or (inputs(133)));
    layer0_outputs(2512) <= (inputs(131)) and not (inputs(25));
    layer0_outputs(2513) <= (inputs(99)) xor (inputs(227));
    layer0_outputs(2514) <= not((inputs(151)) or (inputs(21)));
    layer0_outputs(2515) <= not(inputs(9)) or (inputs(173));
    layer0_outputs(2516) <= (inputs(120)) and not (inputs(190));
    layer0_outputs(2517) <= inputs(203);
    layer0_outputs(2518) <= not(inputs(187)) or (inputs(253));
    layer0_outputs(2519) <= not(inputs(132)) or (inputs(42));
    layer0_outputs(2520) <= (inputs(7)) xor (inputs(27));
    layer0_outputs(2521) <= not(inputs(124)) or (inputs(62));
    layer0_outputs(2522) <= (inputs(140)) or (inputs(215));
    layer0_outputs(2523) <= (inputs(106)) and not (inputs(40));
    layer0_outputs(2524) <= (inputs(21)) xor (inputs(119));
    layer0_outputs(2525) <= not(inputs(38)) or (inputs(5));
    layer0_outputs(2526) <= not(inputs(165));
    layer0_outputs(2527) <= not((inputs(128)) xor (inputs(60)));
    layer0_outputs(2528) <= (inputs(17)) and not (inputs(190));
    layer0_outputs(2529) <= inputs(148);
    layer0_outputs(2530) <= '1';
    layer0_outputs(2531) <= (inputs(76)) xor (inputs(90));
    layer0_outputs(2532) <= inputs(187);
    layer0_outputs(2533) <= not((inputs(62)) xor (inputs(215)));
    layer0_outputs(2534) <= '0';
    layer0_outputs(2535) <= (inputs(55)) and not (inputs(249));
    layer0_outputs(2536) <= not(inputs(245)) or (inputs(232));
    layer0_outputs(2537) <= (inputs(37)) xor (inputs(30));
    layer0_outputs(2538) <= inputs(140);
    layer0_outputs(2539) <= inputs(106);
    layer0_outputs(2540) <= (inputs(11)) and not (inputs(175));
    layer0_outputs(2541) <= (inputs(150)) and (inputs(10));
    layer0_outputs(2542) <= not((inputs(206)) and (inputs(13)));
    layer0_outputs(2543) <= not(inputs(164)) or (inputs(81));
    layer0_outputs(2544) <= (inputs(73)) and not (inputs(97));
    layer0_outputs(2545) <= not(inputs(228)) or (inputs(254));
    layer0_outputs(2546) <= not((inputs(20)) or (inputs(12)));
    layer0_outputs(2547) <= (inputs(169)) and not (inputs(164));
    layer0_outputs(2548) <= inputs(165);
    layer0_outputs(2549) <= inputs(135);
    layer0_outputs(2550) <= (inputs(85)) or (inputs(236));
    layer0_outputs(2551) <= not(inputs(29));
    layer0_outputs(2552) <= not(inputs(230));
    layer0_outputs(2553) <= not((inputs(90)) or (inputs(177)));
    layer0_outputs(2554) <= (inputs(163)) or (inputs(244));
    layer0_outputs(2555) <= (inputs(32)) or (inputs(18));
    layer0_outputs(2556) <= not(inputs(250));
    layer0_outputs(2557) <= not(inputs(75)) or (inputs(3));
    layer0_outputs(2558) <= inputs(127);
    layer0_outputs(2559) <= (inputs(139)) or (inputs(138));
    layer0_outputs(2560) <= not(inputs(86)) or (inputs(97));
    layer0_outputs(2561) <= inputs(175);
    layer0_outputs(2562) <= (inputs(61)) and not (inputs(228));
    layer0_outputs(2563) <= (inputs(171)) xor (inputs(204));
    layer0_outputs(2564) <= (inputs(194)) and not (inputs(203));
    layer0_outputs(2565) <= not(inputs(113)) or (inputs(247));
    layer0_outputs(2566) <= not((inputs(230)) or (inputs(90)));
    layer0_outputs(2567) <= (inputs(97)) and not (inputs(144));
    layer0_outputs(2568) <= '1';
    layer0_outputs(2569) <= (inputs(55)) and not (inputs(17));
    layer0_outputs(2570) <= (inputs(167)) xor (inputs(241));
    layer0_outputs(2571) <= (inputs(85)) and not (inputs(129));
    layer0_outputs(2572) <= (inputs(88)) and not (inputs(110));
    layer0_outputs(2573) <= not(inputs(198)) or (inputs(25));
    layer0_outputs(2574) <= not((inputs(112)) or (inputs(201)));
    layer0_outputs(2575) <= not((inputs(179)) or (inputs(128)));
    layer0_outputs(2576) <= not(inputs(245));
    layer0_outputs(2577) <= (inputs(36)) and not (inputs(29));
    layer0_outputs(2578) <= not(inputs(107)) or (inputs(141));
    layer0_outputs(2579) <= not(inputs(106));
    layer0_outputs(2580) <= not((inputs(239)) or (inputs(43)));
    layer0_outputs(2581) <= '1';
    layer0_outputs(2582) <= (inputs(85)) or (inputs(99));
    layer0_outputs(2583) <= inputs(236);
    layer0_outputs(2584) <= not((inputs(38)) xor (inputs(141)));
    layer0_outputs(2585) <= not(inputs(135)) or (inputs(180));
    layer0_outputs(2586) <= (inputs(240)) and not (inputs(245));
    layer0_outputs(2587) <= inputs(243);
    layer0_outputs(2588) <= (inputs(149)) or (inputs(152));
    layer0_outputs(2589) <= not(inputs(74)) or (inputs(181));
    layer0_outputs(2590) <= (inputs(42)) xor (inputs(72));
    layer0_outputs(2591) <= not(inputs(86)) or (inputs(60));
    layer0_outputs(2592) <= (inputs(37)) and (inputs(113));
    layer0_outputs(2593) <= not(inputs(94)) or (inputs(206));
    layer0_outputs(2594) <= not(inputs(232)) or (inputs(59));
    layer0_outputs(2595) <= not(inputs(153));
    layer0_outputs(2596) <= not(inputs(118)) or (inputs(146));
    layer0_outputs(2597) <= (inputs(239)) xor (inputs(191));
    layer0_outputs(2598) <= (inputs(17)) or (inputs(188));
    layer0_outputs(2599) <= not(inputs(217));
    layer0_outputs(2600) <= not((inputs(86)) xor (inputs(112)));
    layer0_outputs(2601) <= not((inputs(90)) xor (inputs(89)));
    layer0_outputs(2602) <= not((inputs(179)) xor (inputs(240)));
    layer0_outputs(2603) <= not((inputs(99)) xor (inputs(222)));
    layer0_outputs(2604) <= not((inputs(232)) and (inputs(223)));
    layer0_outputs(2605) <= not((inputs(97)) and (inputs(9)));
    layer0_outputs(2606) <= (inputs(59)) xor (inputs(147));
    layer0_outputs(2607) <= not((inputs(252)) or (inputs(122)));
    layer0_outputs(2608) <= not((inputs(74)) xor (inputs(76)));
    layer0_outputs(2609) <= not(inputs(211));
    layer0_outputs(2610) <= not(inputs(180)) or (inputs(17));
    layer0_outputs(2611) <= not(inputs(196));
    layer0_outputs(2612) <= not((inputs(20)) xor (inputs(141)));
    layer0_outputs(2613) <= inputs(118);
    layer0_outputs(2614) <= not((inputs(208)) and (inputs(192)));
    layer0_outputs(2615) <= (inputs(207)) and (inputs(117));
    layer0_outputs(2616) <= (inputs(138)) and not (inputs(180));
    layer0_outputs(2617) <= not(inputs(121)) or (inputs(243));
    layer0_outputs(2618) <= inputs(119);
    layer0_outputs(2619) <= not((inputs(84)) or (inputs(196)));
    layer0_outputs(2620) <= not((inputs(105)) or (inputs(6)));
    layer0_outputs(2621) <= not(inputs(169)) or (inputs(212));
    layer0_outputs(2622) <= (inputs(124)) xor (inputs(187));
    layer0_outputs(2623) <= not(inputs(77));
    layer0_outputs(2624) <= not(inputs(45));
    layer0_outputs(2625) <= (inputs(120)) xor (inputs(188));
    layer0_outputs(2626) <= not(inputs(54)) or (inputs(125));
    layer0_outputs(2627) <= not(inputs(207)) or (inputs(250));
    layer0_outputs(2628) <= not(inputs(218));
    layer0_outputs(2629) <= (inputs(78)) and (inputs(254));
    layer0_outputs(2630) <= (inputs(37)) and not (inputs(128));
    layer0_outputs(2631) <= inputs(91);
    layer0_outputs(2632) <= (inputs(155)) xor (inputs(112));
    layer0_outputs(2633) <= (inputs(198)) xor (inputs(209));
    layer0_outputs(2634) <= inputs(125);
    layer0_outputs(2635) <= (inputs(37)) and (inputs(239));
    layer0_outputs(2636) <= (inputs(150)) xor (inputs(64));
    layer0_outputs(2637) <= inputs(10);
    layer0_outputs(2638) <= (inputs(241)) xor (inputs(186));
    layer0_outputs(2639) <= not((inputs(121)) or (inputs(3)));
    layer0_outputs(2640) <= not(inputs(216)) or (inputs(81));
    layer0_outputs(2641) <= inputs(138);
    layer0_outputs(2642) <= (inputs(166)) and not (inputs(253));
    layer0_outputs(2643) <= not((inputs(140)) xor (inputs(204)));
    layer0_outputs(2644) <= not(inputs(137));
    layer0_outputs(2645) <= not(inputs(105)) or (inputs(0));
    layer0_outputs(2646) <= (inputs(21)) and (inputs(22));
    layer0_outputs(2647) <= '1';
    layer0_outputs(2648) <= not(inputs(172));
    layer0_outputs(2649) <= not(inputs(39)) or (inputs(108));
    layer0_outputs(2650) <= not((inputs(35)) xor (inputs(107)));
    layer0_outputs(2651) <= (inputs(248)) or (inputs(193));
    layer0_outputs(2652) <= not((inputs(190)) and (inputs(243)));
    layer0_outputs(2653) <= inputs(198);
    layer0_outputs(2654) <= not((inputs(37)) or (inputs(155)));
    layer0_outputs(2655) <= not(inputs(91)) or (inputs(45));
    layer0_outputs(2656) <= not((inputs(46)) xor (inputs(82)));
    layer0_outputs(2657) <= not(inputs(75));
    layer0_outputs(2658) <= not(inputs(227)) or (inputs(160));
    layer0_outputs(2659) <= (inputs(225)) or (inputs(239));
    layer0_outputs(2660) <= (inputs(24)) xor (inputs(221));
    layer0_outputs(2661) <= (inputs(134)) and not (inputs(223));
    layer0_outputs(2662) <= (inputs(103)) xor (inputs(255));
    layer0_outputs(2663) <= (inputs(252)) or (inputs(78));
    layer0_outputs(2664) <= not((inputs(72)) or (inputs(206)));
    layer0_outputs(2665) <= (inputs(188)) xor (inputs(172));
    layer0_outputs(2666) <= (inputs(197)) xor (inputs(128));
    layer0_outputs(2667) <= not((inputs(133)) or (inputs(77)));
    layer0_outputs(2668) <= (inputs(40)) xor (inputs(100));
    layer0_outputs(2669) <= (inputs(148)) or (inputs(225));
    layer0_outputs(2670) <= not((inputs(88)) xor (inputs(180)));
    layer0_outputs(2671) <= not(inputs(43)) or (inputs(249));
    layer0_outputs(2672) <= (inputs(202)) or (inputs(150));
    layer0_outputs(2673) <= not(inputs(24));
    layer0_outputs(2674) <= not(inputs(37));
    layer0_outputs(2675) <= (inputs(78)) and not (inputs(206));
    layer0_outputs(2676) <= inputs(111);
    layer0_outputs(2677) <= not(inputs(138));
    layer0_outputs(2678) <= (inputs(175)) and not (inputs(208));
    layer0_outputs(2679) <= (inputs(217)) and not (inputs(27));
    layer0_outputs(2680) <= not((inputs(247)) or (inputs(193)));
    layer0_outputs(2681) <= not(inputs(45));
    layer0_outputs(2682) <= inputs(241);
    layer0_outputs(2683) <= inputs(146);
    layer0_outputs(2684) <= not((inputs(38)) or (inputs(0)));
    layer0_outputs(2685) <= not((inputs(99)) or (inputs(233)));
    layer0_outputs(2686) <= not(inputs(91)) or (inputs(129));
    layer0_outputs(2687) <= not((inputs(154)) xor (inputs(98)));
    layer0_outputs(2688) <= (inputs(169)) and not (inputs(173));
    layer0_outputs(2689) <= inputs(120);
    layer0_outputs(2690) <= (inputs(219)) xor (inputs(243));
    layer0_outputs(2691) <= not((inputs(1)) xor (inputs(97)));
    layer0_outputs(2692) <= (inputs(147)) or (inputs(94));
    layer0_outputs(2693) <= inputs(102);
    layer0_outputs(2694) <= not(inputs(165));
    layer0_outputs(2695) <= not(inputs(235));
    layer0_outputs(2696) <= not(inputs(129)) or (inputs(9));
    layer0_outputs(2697) <= inputs(55);
    layer0_outputs(2698) <= '1';
    layer0_outputs(2699) <= not((inputs(156)) or (inputs(68)));
    layer0_outputs(2700) <= not(inputs(203)) or (inputs(18));
    layer0_outputs(2701) <= not((inputs(85)) or (inputs(83)));
    layer0_outputs(2702) <= not((inputs(226)) or (inputs(29)));
    layer0_outputs(2703) <= not(inputs(165));
    layer0_outputs(2704) <= (inputs(149)) and not (inputs(83));
    layer0_outputs(2705) <= not((inputs(145)) and (inputs(146)));
    layer0_outputs(2706) <= inputs(63);
    layer0_outputs(2707) <= (inputs(24)) or (inputs(164));
    layer0_outputs(2708) <= not(inputs(118)) or (inputs(236));
    layer0_outputs(2709) <= not((inputs(82)) or (inputs(5)));
    layer0_outputs(2710) <= (inputs(178)) or (inputs(9));
    layer0_outputs(2711) <= not((inputs(38)) or (inputs(55)));
    layer0_outputs(2712) <= (inputs(13)) and not (inputs(92));
    layer0_outputs(2713) <= (inputs(47)) xor (inputs(123));
    layer0_outputs(2714) <= inputs(74);
    layer0_outputs(2715) <= (inputs(124)) or (inputs(14));
    layer0_outputs(2716) <= not(inputs(205)) or (inputs(245));
    layer0_outputs(2717) <= not((inputs(96)) or (inputs(95)));
    layer0_outputs(2718) <= not(inputs(106));
    layer0_outputs(2719) <= not((inputs(41)) or (inputs(153)));
    layer0_outputs(2720) <= not((inputs(154)) or (inputs(37)));
    layer0_outputs(2721) <= (inputs(124)) or (inputs(108));
    layer0_outputs(2722) <= inputs(146);
    layer0_outputs(2723) <= (inputs(42)) or (inputs(185));
    layer0_outputs(2724) <= (inputs(74)) and not (inputs(12));
    layer0_outputs(2725) <= not(inputs(136)) or (inputs(127));
    layer0_outputs(2726) <= not((inputs(240)) or (inputs(101)));
    layer0_outputs(2727) <= inputs(164);
    layer0_outputs(2728) <= not((inputs(127)) xor (inputs(93)));
    layer0_outputs(2729) <= (inputs(244)) or (inputs(164));
    layer0_outputs(2730) <= not((inputs(5)) or (inputs(68)));
    layer0_outputs(2731) <= not(inputs(248));
    layer0_outputs(2732) <= not(inputs(7));
    layer0_outputs(2733) <= not(inputs(199));
    layer0_outputs(2734) <= (inputs(21)) and not (inputs(199));
    layer0_outputs(2735) <= not((inputs(4)) xor (inputs(150)));
    layer0_outputs(2736) <= (inputs(40)) and not (inputs(126));
    layer0_outputs(2737) <= not((inputs(122)) xor (inputs(243)));
    layer0_outputs(2738) <= not((inputs(168)) xor (inputs(143)));
    layer0_outputs(2739) <= (inputs(9)) xor (inputs(127));
    layer0_outputs(2740) <= (inputs(214)) and not (inputs(11));
    layer0_outputs(2741) <= (inputs(61)) and not (inputs(81));
    layer0_outputs(2742) <= (inputs(116)) and not (inputs(245));
    layer0_outputs(2743) <= not(inputs(85)) or (inputs(163));
    layer0_outputs(2744) <= (inputs(202)) and not (inputs(36));
    layer0_outputs(2745) <= (inputs(227)) xor (inputs(91));
    layer0_outputs(2746) <= not(inputs(91)) or (inputs(190));
    layer0_outputs(2747) <= not((inputs(31)) xor (inputs(135)));
    layer0_outputs(2748) <= not((inputs(97)) xor (inputs(157)));
    layer0_outputs(2749) <= not((inputs(212)) xor (inputs(239)));
    layer0_outputs(2750) <= (inputs(232)) or (inputs(55));
    layer0_outputs(2751) <= inputs(103);
    layer0_outputs(2752) <= not(inputs(92));
    layer0_outputs(2753) <= (inputs(90)) xor (inputs(8));
    layer0_outputs(2754) <= (inputs(95)) and not (inputs(65));
    layer0_outputs(2755) <= not((inputs(27)) xor (inputs(248)));
    layer0_outputs(2756) <= not((inputs(112)) and (inputs(18)));
    layer0_outputs(2757) <= not(inputs(76)) or (inputs(252));
    layer0_outputs(2758) <= '1';
    layer0_outputs(2759) <= not(inputs(98)) or (inputs(210));
    layer0_outputs(2760) <= not(inputs(27)) or (inputs(111));
    layer0_outputs(2761) <= (inputs(150)) and not (inputs(93));
    layer0_outputs(2762) <= not(inputs(9));
    layer0_outputs(2763) <= not(inputs(63)) or (inputs(242));
    layer0_outputs(2764) <= inputs(177);
    layer0_outputs(2765) <= (inputs(18)) or (inputs(242));
    layer0_outputs(2766) <= inputs(44);
    layer0_outputs(2767) <= inputs(99);
    layer0_outputs(2768) <= not((inputs(216)) or (inputs(137)));
    layer0_outputs(2769) <= (inputs(26)) and not (inputs(65));
    layer0_outputs(2770) <= not(inputs(202));
    layer0_outputs(2771) <= inputs(235);
    layer0_outputs(2772) <= (inputs(146)) and not (inputs(234));
    layer0_outputs(2773) <= not(inputs(52)) or (inputs(6));
    layer0_outputs(2774) <= inputs(94);
    layer0_outputs(2775) <= inputs(188);
    layer0_outputs(2776) <= not((inputs(181)) xor (inputs(213)));
    layer0_outputs(2777) <= not((inputs(249)) or (inputs(40)));
    layer0_outputs(2778) <= not(inputs(128));
    layer0_outputs(2779) <= inputs(176);
    layer0_outputs(2780) <= (inputs(221)) or (inputs(101));
    layer0_outputs(2781) <= inputs(154);
    layer0_outputs(2782) <= (inputs(78)) xor (inputs(146));
    layer0_outputs(2783) <= inputs(218);
    layer0_outputs(2784) <= not((inputs(115)) xor (inputs(166)));
    layer0_outputs(2785) <= not(inputs(233)) or (inputs(124));
    layer0_outputs(2786) <= not((inputs(161)) xor (inputs(213)));
    layer0_outputs(2787) <= (inputs(90)) and not (inputs(44));
    layer0_outputs(2788) <= '1';
    layer0_outputs(2789) <= inputs(122);
    layer0_outputs(2790) <= not(inputs(180));
    layer0_outputs(2791) <= not(inputs(58));
    layer0_outputs(2792) <= (inputs(37)) and not (inputs(33));
    layer0_outputs(2793) <= not((inputs(28)) xor (inputs(23)));
    layer0_outputs(2794) <= '0';
    layer0_outputs(2795) <= (inputs(74)) or (inputs(158));
    layer0_outputs(2796) <= not(inputs(3)) or (inputs(143));
    layer0_outputs(2797) <= (inputs(51)) xor (inputs(184));
    layer0_outputs(2798) <= (inputs(165)) xor (inputs(16));
    layer0_outputs(2799) <= not(inputs(117));
    layer0_outputs(2800) <= inputs(240);
    layer0_outputs(2801) <= not(inputs(218));
    layer0_outputs(2802) <= not((inputs(104)) or (inputs(82)));
    layer0_outputs(2803) <= not((inputs(14)) or (inputs(32)));
    layer0_outputs(2804) <= (inputs(255)) or (inputs(180));
    layer0_outputs(2805) <= not((inputs(56)) xor (inputs(11)));
    layer0_outputs(2806) <= (inputs(114)) or (inputs(131));
    layer0_outputs(2807) <= not(inputs(122)) or (inputs(90));
    layer0_outputs(2808) <= not(inputs(69));
    layer0_outputs(2809) <= not(inputs(93)) or (inputs(30));
    layer0_outputs(2810) <= '1';
    layer0_outputs(2811) <= (inputs(197)) or (inputs(191));
    layer0_outputs(2812) <= not(inputs(141)) or (inputs(177));
    layer0_outputs(2813) <= not(inputs(54));
    layer0_outputs(2814) <= (inputs(248)) and not (inputs(41));
    layer0_outputs(2815) <= not(inputs(219));
    layer0_outputs(2816) <= inputs(249);
    layer0_outputs(2817) <= inputs(227);
    layer0_outputs(2818) <= not((inputs(241)) or (inputs(4)));
    layer0_outputs(2819) <= not((inputs(134)) and (inputs(69)));
    layer0_outputs(2820) <= (inputs(87)) and not (inputs(79));
    layer0_outputs(2821) <= (inputs(163)) xor (inputs(100));
    layer0_outputs(2822) <= (inputs(246)) and not (inputs(78));
    layer0_outputs(2823) <= (inputs(212)) and not (inputs(107));
    layer0_outputs(2824) <= not((inputs(202)) xor (inputs(105)));
    layer0_outputs(2825) <= not((inputs(33)) xor (inputs(104)));
    layer0_outputs(2826) <= (inputs(209)) xor (inputs(161));
    layer0_outputs(2827) <= inputs(74);
    layer0_outputs(2828) <= (inputs(217)) and not (inputs(187));
    layer0_outputs(2829) <= (inputs(148)) xor (inputs(205));
    layer0_outputs(2830) <= not((inputs(146)) xor (inputs(107)));
    layer0_outputs(2831) <= (inputs(89)) or (inputs(34));
    layer0_outputs(2832) <= inputs(94);
    layer0_outputs(2833) <= inputs(104);
    layer0_outputs(2834) <= (inputs(27)) xor (inputs(149));
    layer0_outputs(2835) <= (inputs(11)) or (inputs(173));
    layer0_outputs(2836) <= not(inputs(26));
    layer0_outputs(2837) <= not((inputs(21)) xor (inputs(135)));
    layer0_outputs(2838) <= (inputs(202)) or (inputs(35));
    layer0_outputs(2839) <= (inputs(185)) xor (inputs(183));
    layer0_outputs(2840) <= not(inputs(124)) or (inputs(44));
    layer0_outputs(2841) <= not((inputs(85)) or (inputs(214)));
    layer0_outputs(2842) <= (inputs(48)) xor (inputs(130));
    layer0_outputs(2843) <= not(inputs(6));
    layer0_outputs(2844) <= not((inputs(11)) or (inputs(40)));
    layer0_outputs(2845) <= not(inputs(77));
    layer0_outputs(2846) <= not((inputs(104)) or (inputs(217)));
    layer0_outputs(2847) <= (inputs(120)) and not (inputs(138));
    layer0_outputs(2848) <= (inputs(161)) and not (inputs(178));
    layer0_outputs(2849) <= '1';
    layer0_outputs(2850) <= (inputs(209)) or (inputs(132));
    layer0_outputs(2851) <= (inputs(140)) and (inputs(12));
    layer0_outputs(2852) <= not((inputs(39)) xor (inputs(249)));
    layer0_outputs(2853) <= not((inputs(208)) xor (inputs(249)));
    layer0_outputs(2854) <= not(inputs(166));
    layer0_outputs(2855) <= not((inputs(152)) or (inputs(250)));
    layer0_outputs(2856) <= (inputs(136)) or (inputs(164));
    layer0_outputs(2857) <= (inputs(91)) and not (inputs(196));
    layer0_outputs(2858) <= (inputs(169)) and not (inputs(25));
    layer0_outputs(2859) <= inputs(233);
    layer0_outputs(2860) <= (inputs(178)) xor (inputs(193));
    layer0_outputs(2861) <= (inputs(215)) or (inputs(31));
    layer0_outputs(2862) <= (inputs(74)) xor (inputs(48));
    layer0_outputs(2863) <= not(inputs(168));
    layer0_outputs(2864) <= not((inputs(8)) or (inputs(151)));
    layer0_outputs(2865) <= not(inputs(66)) or (inputs(80));
    layer0_outputs(2866) <= (inputs(121)) and not (inputs(162));
    layer0_outputs(2867) <= '0';
    layer0_outputs(2868) <= inputs(44);
    layer0_outputs(2869) <= inputs(89);
    layer0_outputs(2870) <= not((inputs(35)) or (inputs(139)));
    layer0_outputs(2871) <= (inputs(66)) and (inputs(227));
    layer0_outputs(2872) <= not(inputs(162)) or (inputs(61));
    layer0_outputs(2873) <= not(inputs(162));
    layer0_outputs(2874) <= (inputs(149)) and not (inputs(189));
    layer0_outputs(2875) <= not((inputs(122)) or (inputs(169)));
    layer0_outputs(2876) <= not(inputs(100));
    layer0_outputs(2877) <= not(inputs(194));
    layer0_outputs(2878) <= not(inputs(152)) or (inputs(4));
    layer0_outputs(2879) <= not((inputs(205)) and (inputs(254)));
    layer0_outputs(2880) <= (inputs(212)) xor (inputs(190));
    layer0_outputs(2881) <= (inputs(155)) or (inputs(207));
    layer0_outputs(2882) <= not(inputs(13)) or (inputs(244));
    layer0_outputs(2883) <= not((inputs(116)) or (inputs(246)));
    layer0_outputs(2884) <= (inputs(116)) xor (inputs(104));
    layer0_outputs(2885) <= (inputs(31)) and not (inputs(96));
    layer0_outputs(2886) <= not((inputs(197)) xor (inputs(71)));
    layer0_outputs(2887) <= not((inputs(99)) or (inputs(20)));
    layer0_outputs(2888) <= (inputs(183)) or (inputs(10));
    layer0_outputs(2889) <= not((inputs(252)) xor (inputs(135)));
    layer0_outputs(2890) <= (inputs(109)) xor (inputs(12));
    layer0_outputs(2891) <= not(inputs(78));
    layer0_outputs(2892) <= (inputs(121)) or (inputs(233));
    layer0_outputs(2893) <= (inputs(202)) and not (inputs(9));
    layer0_outputs(2894) <= not((inputs(88)) xor (inputs(216)));
    layer0_outputs(2895) <= '1';
    layer0_outputs(2896) <= not((inputs(77)) or (inputs(170)));
    layer0_outputs(2897) <= inputs(51);
    layer0_outputs(2898) <= (inputs(91)) xor (inputs(232));
    layer0_outputs(2899) <= inputs(123);
    layer0_outputs(2900) <= not(inputs(40));
    layer0_outputs(2901) <= not((inputs(64)) xor (inputs(65)));
    layer0_outputs(2902) <= inputs(161);
    layer0_outputs(2903) <= not((inputs(180)) or (inputs(222)));
    layer0_outputs(2904) <= not(inputs(193));
    layer0_outputs(2905) <= (inputs(135)) or (inputs(22));
    layer0_outputs(2906) <= not(inputs(17));
    layer0_outputs(2907) <= not((inputs(132)) and (inputs(137)));
    layer0_outputs(2908) <= not((inputs(27)) xor (inputs(12)));
    layer0_outputs(2909) <= (inputs(243)) or (inputs(218));
    layer0_outputs(2910) <= inputs(50);
    layer0_outputs(2911) <= not(inputs(145));
    layer0_outputs(2912) <= not(inputs(217)) or (inputs(130));
    layer0_outputs(2913) <= (inputs(130)) xor (inputs(137));
    layer0_outputs(2914) <= not(inputs(180)) or (inputs(156));
    layer0_outputs(2915) <= not((inputs(88)) xor (inputs(74)));
    layer0_outputs(2916) <= not((inputs(222)) xor (inputs(71)));
    layer0_outputs(2917) <= (inputs(125)) and not (inputs(4));
    layer0_outputs(2918) <= (inputs(115)) xor (inputs(177));
    layer0_outputs(2919) <= (inputs(156)) or (inputs(131));
    layer0_outputs(2920) <= inputs(73);
    layer0_outputs(2921) <= not(inputs(32));
    layer0_outputs(2922) <= not(inputs(139)) or (inputs(237));
    layer0_outputs(2923) <= '1';
    layer0_outputs(2924) <= not((inputs(156)) or (inputs(44)));
    layer0_outputs(2925) <= not(inputs(177));
    layer0_outputs(2926) <= (inputs(147)) and not (inputs(210));
    layer0_outputs(2927) <= not(inputs(185));
    layer0_outputs(2928) <= (inputs(49)) and (inputs(10));
    layer0_outputs(2929) <= not((inputs(57)) xor (inputs(67)));
    layer0_outputs(2930) <= (inputs(27)) or (inputs(219));
    layer0_outputs(2931) <= not((inputs(6)) xor (inputs(132)));
    layer0_outputs(2932) <= (inputs(180)) and not (inputs(35));
    layer0_outputs(2933) <= (inputs(39)) or (inputs(204));
    layer0_outputs(2934) <= not(inputs(9)) or (inputs(210));
    layer0_outputs(2935) <= not(inputs(77)) or (inputs(33));
    layer0_outputs(2936) <= not((inputs(214)) xor (inputs(200)));
    layer0_outputs(2937) <= (inputs(168)) or (inputs(210));
    layer0_outputs(2938) <= (inputs(185)) and not (inputs(80));
    layer0_outputs(2939) <= (inputs(132)) and not (inputs(254));
    layer0_outputs(2940) <= not(inputs(214)) or (inputs(21));
    layer0_outputs(2941) <= not(inputs(239)) or (inputs(35));
    layer0_outputs(2942) <= (inputs(151)) xor (inputs(168));
    layer0_outputs(2943) <= (inputs(252)) and (inputs(130));
    layer0_outputs(2944) <= '1';
    layer0_outputs(2945) <= inputs(56);
    layer0_outputs(2946) <= inputs(57);
    layer0_outputs(2947) <= not(inputs(17)) or (inputs(175));
    layer0_outputs(2948) <= (inputs(152)) and not (inputs(203));
    layer0_outputs(2949) <= not(inputs(255)) or (inputs(214));
    layer0_outputs(2950) <= inputs(199);
    layer0_outputs(2951) <= not((inputs(24)) xor (inputs(207)));
    layer0_outputs(2952) <= not(inputs(218)) or (inputs(111));
    layer0_outputs(2953) <= not((inputs(207)) or (inputs(251)));
    layer0_outputs(2954) <= (inputs(105)) and not (inputs(103));
    layer0_outputs(2955) <= not(inputs(230)) or (inputs(79));
    layer0_outputs(2956) <= (inputs(145)) and not (inputs(222));
    layer0_outputs(2957) <= not(inputs(213)) or (inputs(100));
    layer0_outputs(2958) <= (inputs(75)) and not (inputs(146));
    layer0_outputs(2959) <= (inputs(78)) and not (inputs(158));
    layer0_outputs(2960) <= (inputs(38)) and not (inputs(217));
    layer0_outputs(2961) <= not(inputs(98)) or (inputs(226));
    layer0_outputs(2962) <= not((inputs(110)) or (inputs(78)));
    layer0_outputs(2963) <= not((inputs(18)) xor (inputs(118)));
    layer0_outputs(2964) <= not((inputs(150)) or (inputs(128)));
    layer0_outputs(2965) <= inputs(102);
    layer0_outputs(2966) <= not(inputs(39)) or (inputs(173));
    layer0_outputs(2967) <= (inputs(176)) and not (inputs(124));
    layer0_outputs(2968) <= (inputs(116)) or (inputs(140));
    layer0_outputs(2969) <= not(inputs(253)) or (inputs(142));
    layer0_outputs(2970) <= inputs(115);
    layer0_outputs(2971) <= not((inputs(223)) or (inputs(219)));
    layer0_outputs(2972) <= (inputs(102)) and not (inputs(236));
    layer0_outputs(2973) <= (inputs(89)) or (inputs(21));
    layer0_outputs(2974) <= not(inputs(137));
    layer0_outputs(2975) <= not(inputs(114));
    layer0_outputs(2976) <= (inputs(222)) xor (inputs(170));
    layer0_outputs(2977) <= not((inputs(76)) or (inputs(70)));
    layer0_outputs(2978) <= '1';
    layer0_outputs(2979) <= not(inputs(101));
    layer0_outputs(2980) <= (inputs(162)) or (inputs(17));
    layer0_outputs(2981) <= not(inputs(245)) or (inputs(126));
    layer0_outputs(2982) <= inputs(116);
    layer0_outputs(2983) <= not((inputs(211)) xor (inputs(233)));
    layer0_outputs(2984) <= not((inputs(195)) xor (inputs(51)));
    layer0_outputs(2985) <= not(inputs(250)) or (inputs(0));
    layer0_outputs(2986) <= not(inputs(188));
    layer0_outputs(2987) <= (inputs(121)) xor (inputs(125));
    layer0_outputs(2988) <= not(inputs(103));
    layer0_outputs(2989) <= not(inputs(41)) or (inputs(147));
    layer0_outputs(2990) <= not((inputs(248)) and (inputs(108)));
    layer0_outputs(2991) <= inputs(24);
    layer0_outputs(2992) <= (inputs(3)) and not (inputs(49));
    layer0_outputs(2993) <= not((inputs(36)) or (inputs(180)));
    layer0_outputs(2994) <= (inputs(12)) xor (inputs(150));
    layer0_outputs(2995) <= (inputs(228)) xor (inputs(157));
    layer0_outputs(2996) <= not(inputs(84));
    layer0_outputs(2997) <= (inputs(224)) or (inputs(246));
    layer0_outputs(2998) <= (inputs(78)) and not (inputs(25));
    layer0_outputs(2999) <= not((inputs(112)) xor (inputs(102)));
    layer0_outputs(3000) <= not((inputs(231)) or (inputs(55)));
    layer0_outputs(3001) <= (inputs(233)) xor (inputs(227));
    layer0_outputs(3002) <= not(inputs(182)) or (inputs(236));
    layer0_outputs(3003) <= (inputs(3)) or (inputs(215));
    layer0_outputs(3004) <= (inputs(104)) and not (inputs(235));
    layer0_outputs(3005) <= (inputs(98)) or (inputs(58));
    layer0_outputs(3006) <= not((inputs(104)) xor (inputs(22)));
    layer0_outputs(3007) <= '1';
    layer0_outputs(3008) <= not(inputs(121));
    layer0_outputs(3009) <= not((inputs(143)) and (inputs(174)));
    layer0_outputs(3010) <= not((inputs(250)) and (inputs(49)));
    layer0_outputs(3011) <= (inputs(108)) and not (inputs(177));
    layer0_outputs(3012) <= (inputs(7)) or (inputs(119));
    layer0_outputs(3013) <= not((inputs(155)) xor (inputs(200)));
    layer0_outputs(3014) <= not((inputs(144)) or (inputs(242)));
    layer0_outputs(3015) <= not((inputs(68)) or (inputs(193)));
    layer0_outputs(3016) <= (inputs(183)) or (inputs(66));
    layer0_outputs(3017) <= not(inputs(57)) or (inputs(249));
    layer0_outputs(3018) <= (inputs(182)) and not (inputs(11));
    layer0_outputs(3019) <= not((inputs(26)) or (inputs(137)));
    layer0_outputs(3020) <= (inputs(109)) xor (inputs(242));
    layer0_outputs(3021) <= not((inputs(228)) or (inputs(248)));
    layer0_outputs(3022) <= inputs(179);
    layer0_outputs(3023) <= (inputs(230)) and not (inputs(60));
    layer0_outputs(3024) <= (inputs(71)) xor (inputs(185));
    layer0_outputs(3025) <= not(inputs(56));
    layer0_outputs(3026) <= (inputs(23)) or (inputs(198));
    layer0_outputs(3027) <= '1';
    layer0_outputs(3028) <= not(inputs(180)) or (inputs(114));
    layer0_outputs(3029) <= not((inputs(193)) xor (inputs(188)));
    layer0_outputs(3030) <= not((inputs(70)) xor (inputs(102)));
    layer0_outputs(3031) <= not(inputs(162)) or (inputs(109));
    layer0_outputs(3032) <= not((inputs(111)) or (inputs(100)));
    layer0_outputs(3033) <= not(inputs(255));
    layer0_outputs(3034) <= (inputs(1)) and not (inputs(22));
    layer0_outputs(3035) <= (inputs(195)) xor (inputs(64));
    layer0_outputs(3036) <= not(inputs(155)) or (inputs(251));
    layer0_outputs(3037) <= not(inputs(235));
    layer0_outputs(3038) <= (inputs(168)) xor (inputs(249));
    layer0_outputs(3039) <= (inputs(236)) and not (inputs(43));
    layer0_outputs(3040) <= inputs(168);
    layer0_outputs(3041) <= not(inputs(123));
    layer0_outputs(3042) <= (inputs(30)) or (inputs(233));
    layer0_outputs(3043) <= '1';
    layer0_outputs(3044) <= not((inputs(181)) or (inputs(104)));
    layer0_outputs(3045) <= not((inputs(216)) xor (inputs(204)));
    layer0_outputs(3046) <= not((inputs(158)) xor (inputs(51)));
    layer0_outputs(3047) <= not((inputs(202)) xor (inputs(253)));
    layer0_outputs(3048) <= (inputs(154)) and not (inputs(214));
    layer0_outputs(3049) <= inputs(219);
    layer0_outputs(3050) <= not((inputs(11)) and (inputs(1)));
    layer0_outputs(3051) <= (inputs(91)) and (inputs(54));
    layer0_outputs(3052) <= not((inputs(184)) and (inputs(153)));
    layer0_outputs(3053) <= not((inputs(255)) xor (inputs(89)));
    layer0_outputs(3054) <= (inputs(196)) and not (inputs(159));
    layer0_outputs(3055) <= inputs(73);
    layer0_outputs(3056) <= (inputs(222)) and not (inputs(21));
    layer0_outputs(3057) <= (inputs(91)) or (inputs(149));
    layer0_outputs(3058) <= not((inputs(248)) or (inputs(57)));
    layer0_outputs(3059) <= not((inputs(109)) or (inputs(60)));
    layer0_outputs(3060) <= (inputs(50)) or (inputs(174));
    layer0_outputs(3061) <= (inputs(215)) and not (inputs(129));
    layer0_outputs(3062) <= inputs(203);
    layer0_outputs(3063) <= (inputs(25)) and not (inputs(46));
    layer0_outputs(3064) <= not((inputs(20)) or (inputs(51)));
    layer0_outputs(3065) <= not(inputs(154));
    layer0_outputs(3066) <= not((inputs(14)) xor (inputs(242)));
    layer0_outputs(3067) <= (inputs(146)) or (inputs(54));
    layer0_outputs(3068) <= inputs(241);
    layer0_outputs(3069) <= not(inputs(107));
    layer0_outputs(3070) <= not(inputs(112)) or (inputs(144));
    layer0_outputs(3071) <= not(inputs(183)) or (inputs(231));
    layer0_outputs(3072) <= not(inputs(87)) or (inputs(194));
    layer0_outputs(3073) <= not((inputs(144)) or (inputs(188)));
    layer0_outputs(3074) <= '0';
    layer0_outputs(3075) <= (inputs(167)) and not (inputs(212));
    layer0_outputs(3076) <= not(inputs(123)) or (inputs(97));
    layer0_outputs(3077) <= not((inputs(9)) xor (inputs(235)));
    layer0_outputs(3078) <= inputs(152);
    layer0_outputs(3079) <= (inputs(30)) and not (inputs(254));
    layer0_outputs(3080) <= (inputs(80)) and not (inputs(223));
    layer0_outputs(3081) <= not(inputs(222)) or (inputs(96));
    layer0_outputs(3082) <= not(inputs(248));
    layer0_outputs(3083) <= not((inputs(197)) or (inputs(75)));
    layer0_outputs(3084) <= not((inputs(208)) and (inputs(42)));
    layer0_outputs(3085) <= inputs(124);
    layer0_outputs(3086) <= inputs(172);
    layer0_outputs(3087) <= not((inputs(31)) xor (inputs(153)));
    layer0_outputs(3088) <= not(inputs(104)) or (inputs(88));
    layer0_outputs(3089) <= (inputs(220)) and not (inputs(250));
    layer0_outputs(3090) <= not((inputs(95)) or (inputs(204)));
    layer0_outputs(3091) <= not(inputs(181));
    layer0_outputs(3092) <= (inputs(23)) and not (inputs(236));
    layer0_outputs(3093) <= (inputs(104)) or (inputs(242));
    layer0_outputs(3094) <= not((inputs(184)) xor (inputs(139)));
    layer0_outputs(3095) <= not((inputs(51)) and (inputs(104)));
    layer0_outputs(3096) <= not((inputs(77)) xor (inputs(79)));
    layer0_outputs(3097) <= (inputs(25)) xor (inputs(95));
    layer0_outputs(3098) <= not(inputs(56));
    layer0_outputs(3099) <= '1';
    layer0_outputs(3100) <= (inputs(13)) xor (inputs(120));
    layer0_outputs(3101) <= (inputs(80)) or (inputs(95));
    layer0_outputs(3102) <= not(inputs(196));
    layer0_outputs(3103) <= (inputs(19)) or (inputs(168));
    layer0_outputs(3104) <= not(inputs(15)) or (inputs(111));
    layer0_outputs(3105) <= (inputs(231)) or (inputs(140));
    layer0_outputs(3106) <= (inputs(105)) and not (inputs(60));
    layer0_outputs(3107) <= not((inputs(1)) or (inputs(102)));
    layer0_outputs(3108) <= (inputs(58)) xor (inputs(77));
    layer0_outputs(3109) <= (inputs(205)) or (inputs(167));
    layer0_outputs(3110) <= not((inputs(43)) xor (inputs(219)));
    layer0_outputs(3111) <= not((inputs(159)) xor (inputs(214)));
    layer0_outputs(3112) <= not((inputs(123)) or (inputs(221)));
    layer0_outputs(3113) <= (inputs(167)) or (inputs(68));
    layer0_outputs(3114) <= (inputs(140)) and not (inputs(44));
    layer0_outputs(3115) <= (inputs(106)) xor (inputs(52));
    layer0_outputs(3116) <= not((inputs(221)) xor (inputs(192)));
    layer0_outputs(3117) <= (inputs(215)) and not (inputs(229));
    layer0_outputs(3118) <= not(inputs(78)) or (inputs(174));
    layer0_outputs(3119) <= (inputs(250)) or (inputs(20));
    layer0_outputs(3120) <= inputs(222);
    layer0_outputs(3121) <= (inputs(225)) and not (inputs(188));
    layer0_outputs(3122) <= not((inputs(208)) xor (inputs(155)));
    layer0_outputs(3123) <= '0';
    layer0_outputs(3124) <= not(inputs(105));
    layer0_outputs(3125) <= '1';
    layer0_outputs(3126) <= inputs(40);
    layer0_outputs(3127) <= not((inputs(210)) and (inputs(206)));
    layer0_outputs(3128) <= not((inputs(255)) or (inputs(154)));
    layer0_outputs(3129) <= inputs(133);
    layer0_outputs(3130) <= inputs(76);
    layer0_outputs(3131) <= not(inputs(214)) or (inputs(32));
    layer0_outputs(3132) <= '1';
    layer0_outputs(3133) <= (inputs(96)) or (inputs(186));
    layer0_outputs(3134) <= (inputs(188)) and (inputs(28));
    layer0_outputs(3135) <= (inputs(222)) and not (inputs(209));
    layer0_outputs(3136) <= (inputs(160)) xor (inputs(112));
    layer0_outputs(3137) <= inputs(170);
    layer0_outputs(3138) <= (inputs(93)) or (inputs(17));
    layer0_outputs(3139) <= not((inputs(42)) and (inputs(20)));
    layer0_outputs(3140) <= not((inputs(182)) or (inputs(165)));
    layer0_outputs(3141) <= not(inputs(68));
    layer0_outputs(3142) <= not(inputs(151));
    layer0_outputs(3143) <= (inputs(183)) xor (inputs(223));
    layer0_outputs(3144) <= not(inputs(3)) or (inputs(205));
    layer0_outputs(3145) <= not(inputs(106)) or (inputs(52));
    layer0_outputs(3146) <= not((inputs(181)) or (inputs(17)));
    layer0_outputs(3147) <= not((inputs(99)) xor (inputs(116)));
    layer0_outputs(3148) <= '1';
    layer0_outputs(3149) <= not((inputs(15)) or (inputs(173)));
    layer0_outputs(3150) <= not((inputs(90)) xor (inputs(32)));
    layer0_outputs(3151) <= not(inputs(65)) or (inputs(25));
    layer0_outputs(3152) <= (inputs(222)) xor (inputs(55));
    layer0_outputs(3153) <= (inputs(26)) and not (inputs(229));
    layer0_outputs(3154) <= not(inputs(207));
    layer0_outputs(3155) <= (inputs(92)) xor (inputs(223));
    layer0_outputs(3156) <= not(inputs(138)) or (inputs(77));
    layer0_outputs(3157) <= '0';
    layer0_outputs(3158) <= inputs(135);
    layer0_outputs(3159) <= inputs(107);
    layer0_outputs(3160) <= (inputs(168)) or (inputs(105));
    layer0_outputs(3161) <= not(inputs(197));
    layer0_outputs(3162) <= (inputs(76)) xor (inputs(81));
    layer0_outputs(3163) <= not(inputs(4));
    layer0_outputs(3164) <= inputs(92);
    layer0_outputs(3165) <= (inputs(126)) and not (inputs(24));
    layer0_outputs(3166) <= not((inputs(51)) xor (inputs(92)));
    layer0_outputs(3167) <= (inputs(71)) xor (inputs(218));
    layer0_outputs(3168) <= not((inputs(136)) xor (inputs(63)));
    layer0_outputs(3169) <= inputs(119);
    layer0_outputs(3170) <= (inputs(97)) or (inputs(65));
    layer0_outputs(3171) <= not((inputs(102)) xor (inputs(70)));
    layer0_outputs(3172) <= (inputs(67)) and not (inputs(225));
    layer0_outputs(3173) <= (inputs(242)) or (inputs(189));
    layer0_outputs(3174) <= not((inputs(199)) xor (inputs(234)));
    layer0_outputs(3175) <= (inputs(231)) or (inputs(182));
    layer0_outputs(3176) <= (inputs(80)) or (inputs(58));
    layer0_outputs(3177) <= not(inputs(169));
    layer0_outputs(3178) <= not((inputs(152)) xor (inputs(175)));
    layer0_outputs(3179) <= inputs(117);
    layer0_outputs(3180) <= inputs(133);
    layer0_outputs(3181) <= not(inputs(239));
    layer0_outputs(3182) <= (inputs(209)) xor (inputs(115));
    layer0_outputs(3183) <= (inputs(22)) and (inputs(41));
    layer0_outputs(3184) <= not(inputs(151)) or (inputs(38));
    layer0_outputs(3185) <= inputs(77);
    layer0_outputs(3186) <= not((inputs(64)) or (inputs(193)));
    layer0_outputs(3187) <= not(inputs(178));
    layer0_outputs(3188) <= not((inputs(152)) xor (inputs(95)));
    layer0_outputs(3189) <= not((inputs(103)) xor (inputs(245)));
    layer0_outputs(3190) <= not((inputs(113)) xor (inputs(13)));
    layer0_outputs(3191) <= not((inputs(129)) or (inputs(154)));
    layer0_outputs(3192) <= not(inputs(35)) or (inputs(130));
    layer0_outputs(3193) <= (inputs(135)) xor (inputs(254));
    layer0_outputs(3194) <= (inputs(179)) xor (inputs(253));
    layer0_outputs(3195) <= '1';
    layer0_outputs(3196) <= not((inputs(63)) or (inputs(241)));
    layer0_outputs(3197) <= not(inputs(154)) or (inputs(241));
    layer0_outputs(3198) <= not(inputs(124));
    layer0_outputs(3199) <= (inputs(19)) or (inputs(180));
    layer0_outputs(3200) <= not(inputs(59));
    layer0_outputs(3201) <= not(inputs(149)) or (inputs(128));
    layer0_outputs(3202) <= (inputs(5)) xor (inputs(86));
    layer0_outputs(3203) <= not(inputs(149));
    layer0_outputs(3204) <= (inputs(201)) and not (inputs(161));
    layer0_outputs(3205) <= (inputs(12)) or (inputs(22));
    layer0_outputs(3206) <= not(inputs(229));
    layer0_outputs(3207) <= not(inputs(214)) or (inputs(147));
    layer0_outputs(3208) <= inputs(213);
    layer0_outputs(3209) <= not((inputs(53)) xor (inputs(238)));
    layer0_outputs(3210) <= not(inputs(177)) or (inputs(58));
    layer0_outputs(3211) <= not(inputs(23)) or (inputs(180));
    layer0_outputs(3212) <= not(inputs(73));
    layer0_outputs(3213) <= not(inputs(102)) or (inputs(238));
    layer0_outputs(3214) <= not(inputs(25)) or (inputs(254));
    layer0_outputs(3215) <= (inputs(200)) and not (inputs(221));
    layer0_outputs(3216) <= (inputs(145)) or (inputs(78));
    layer0_outputs(3217) <= inputs(80);
    layer0_outputs(3218) <= (inputs(227)) xor (inputs(234));
    layer0_outputs(3219) <= not((inputs(129)) or (inputs(57)));
    layer0_outputs(3220) <= not((inputs(27)) xor (inputs(143)));
    layer0_outputs(3221) <= not((inputs(124)) or (inputs(202)));
    layer0_outputs(3222) <= (inputs(109)) and (inputs(22));
    layer0_outputs(3223) <= (inputs(46)) or (inputs(156));
    layer0_outputs(3224) <= '0';
    layer0_outputs(3225) <= not(inputs(58)) or (inputs(88));
    layer0_outputs(3226) <= inputs(60);
    layer0_outputs(3227) <= (inputs(125)) xor (inputs(123));
    layer0_outputs(3228) <= not(inputs(218)) or (inputs(28));
    layer0_outputs(3229) <= (inputs(103)) and not (inputs(223));
    layer0_outputs(3230) <= (inputs(42)) and not (inputs(163));
    layer0_outputs(3231) <= inputs(18);
    layer0_outputs(3232) <= not(inputs(88));
    layer0_outputs(3233) <= not(inputs(240));
    layer0_outputs(3234) <= not(inputs(181)) or (inputs(160));
    layer0_outputs(3235) <= (inputs(131)) xor (inputs(225));
    layer0_outputs(3236) <= (inputs(87)) or (inputs(5));
    layer0_outputs(3237) <= not((inputs(0)) and (inputs(21)));
    layer0_outputs(3238) <= (inputs(239)) xor (inputs(196));
    layer0_outputs(3239) <= not((inputs(79)) xor (inputs(195)));
    layer0_outputs(3240) <= '1';
    layer0_outputs(3241) <= (inputs(57)) or (inputs(26));
    layer0_outputs(3242) <= '0';
    layer0_outputs(3243) <= not((inputs(161)) xor (inputs(71)));
    layer0_outputs(3244) <= not(inputs(70));
    layer0_outputs(3245) <= not(inputs(134)) or (inputs(112));
    layer0_outputs(3246) <= (inputs(109)) or (inputs(230));
    layer0_outputs(3247) <= (inputs(130)) and not (inputs(26));
    layer0_outputs(3248) <= (inputs(106)) and not (inputs(61));
    layer0_outputs(3249) <= (inputs(29)) and (inputs(186));
    layer0_outputs(3250) <= not((inputs(32)) or (inputs(230)));
    layer0_outputs(3251) <= not(inputs(45));
    layer0_outputs(3252) <= (inputs(229)) or (inputs(104));
    layer0_outputs(3253) <= inputs(104);
    layer0_outputs(3254) <= not(inputs(147)) or (inputs(198));
    layer0_outputs(3255) <= not((inputs(154)) and (inputs(212)));
    layer0_outputs(3256) <= (inputs(54)) or (inputs(75));
    layer0_outputs(3257) <= not((inputs(201)) or (inputs(23)));
    layer0_outputs(3258) <= not((inputs(145)) and (inputs(70)));
    layer0_outputs(3259) <= (inputs(6)) and not (inputs(249));
    layer0_outputs(3260) <= (inputs(218)) or (inputs(20));
    layer0_outputs(3261) <= inputs(137);
    layer0_outputs(3262) <= (inputs(182)) and not (inputs(219));
    layer0_outputs(3263) <= (inputs(191)) xor (inputs(66));
    layer0_outputs(3264) <= not((inputs(207)) xor (inputs(227)));
    layer0_outputs(3265) <= not((inputs(84)) or (inputs(213)));
    layer0_outputs(3266) <= (inputs(248)) and (inputs(224));
    layer0_outputs(3267) <= (inputs(16)) or (inputs(83));
    layer0_outputs(3268) <= (inputs(132)) xor (inputs(213));
    layer0_outputs(3269) <= not(inputs(155)) or (inputs(129));
    layer0_outputs(3270) <= (inputs(67)) or (inputs(217));
    layer0_outputs(3271) <= (inputs(215)) and (inputs(69));
    layer0_outputs(3272) <= (inputs(112)) and (inputs(254));
    layer0_outputs(3273) <= not(inputs(177)) or (inputs(19));
    layer0_outputs(3274) <= (inputs(201)) xor (inputs(197));
    layer0_outputs(3275) <= not(inputs(135));
    layer0_outputs(3276) <= inputs(0);
    layer0_outputs(3277) <= (inputs(184)) or (inputs(46));
    layer0_outputs(3278) <= not((inputs(101)) or (inputs(20)));
    layer0_outputs(3279) <= (inputs(107)) xor (inputs(140));
    layer0_outputs(3280) <= inputs(242);
    layer0_outputs(3281) <= not((inputs(54)) xor (inputs(163)));
    layer0_outputs(3282) <= (inputs(202)) xor (inputs(42));
    layer0_outputs(3283) <= not(inputs(175));
    layer0_outputs(3284) <= not(inputs(184));
    layer0_outputs(3285) <= not(inputs(109)) or (inputs(11));
    layer0_outputs(3286) <= (inputs(88)) and not (inputs(159));
    layer0_outputs(3287) <= (inputs(56)) and not (inputs(36));
    layer0_outputs(3288) <= inputs(136);
    layer0_outputs(3289) <= not((inputs(113)) and (inputs(98)));
    layer0_outputs(3290) <= inputs(120);
    layer0_outputs(3291) <= not((inputs(204)) or (inputs(43)));
    layer0_outputs(3292) <= not((inputs(212)) xor (inputs(83)));
    layer0_outputs(3293) <= not(inputs(174)) or (inputs(33));
    layer0_outputs(3294) <= not(inputs(191)) or (inputs(10));
    layer0_outputs(3295) <= not((inputs(57)) or (inputs(157)));
    layer0_outputs(3296) <= inputs(117);
    layer0_outputs(3297) <= inputs(137);
    layer0_outputs(3298) <= not(inputs(53)) or (inputs(243));
    layer0_outputs(3299) <= (inputs(234)) and not (inputs(28));
    layer0_outputs(3300) <= not(inputs(130));
    layer0_outputs(3301) <= (inputs(107)) and not (inputs(6));
    layer0_outputs(3302) <= not(inputs(123)) or (inputs(229));
    layer0_outputs(3303) <= not(inputs(61));
    layer0_outputs(3304) <= inputs(16);
    layer0_outputs(3305) <= inputs(127);
    layer0_outputs(3306) <= not((inputs(193)) xor (inputs(66)));
    layer0_outputs(3307) <= (inputs(71)) xor (inputs(0));
    layer0_outputs(3308) <= not(inputs(137));
    layer0_outputs(3309) <= not(inputs(119));
    layer0_outputs(3310) <= inputs(214);
    layer0_outputs(3311) <= (inputs(204)) and not (inputs(99));
    layer0_outputs(3312) <= not(inputs(115));
    layer0_outputs(3313) <= inputs(110);
    layer0_outputs(3314) <= inputs(161);
    layer0_outputs(3315) <= (inputs(211)) or (inputs(195));
    layer0_outputs(3316) <= (inputs(162)) or (inputs(11));
    layer0_outputs(3317) <= inputs(139);
    layer0_outputs(3318) <= not(inputs(192));
    layer0_outputs(3319) <= not(inputs(18)) or (inputs(181));
    layer0_outputs(3320) <= not(inputs(55));
    layer0_outputs(3321) <= (inputs(109)) and not (inputs(127));
    layer0_outputs(3322) <= (inputs(102)) or (inputs(44));
    layer0_outputs(3323) <= (inputs(174)) or (inputs(253));
    layer0_outputs(3324) <= (inputs(60)) and not (inputs(80));
    layer0_outputs(3325) <= not((inputs(26)) and (inputs(7)));
    layer0_outputs(3326) <= (inputs(71)) and not (inputs(192));
    layer0_outputs(3327) <= (inputs(133)) and not (inputs(97));
    layer0_outputs(3328) <= not(inputs(147));
    layer0_outputs(3329) <= (inputs(187)) and not (inputs(18));
    layer0_outputs(3330) <= (inputs(241)) or (inputs(18));
    layer0_outputs(3331) <= '0';
    layer0_outputs(3332) <= (inputs(201)) or (inputs(224));
    layer0_outputs(3333) <= not(inputs(84));
    layer0_outputs(3334) <= not(inputs(89));
    layer0_outputs(3335) <= not(inputs(90)) or (inputs(159));
    layer0_outputs(3336) <= not(inputs(86));
    layer0_outputs(3337) <= not(inputs(84)) or (inputs(29));
    layer0_outputs(3338) <= inputs(225);
    layer0_outputs(3339) <= (inputs(57)) and not (inputs(215));
    layer0_outputs(3340) <= not(inputs(104)) or (inputs(6));
    layer0_outputs(3341) <= not((inputs(225)) xor (inputs(105)));
    layer0_outputs(3342) <= not((inputs(206)) or (inputs(40)));
    layer0_outputs(3343) <= (inputs(193)) and not (inputs(108));
    layer0_outputs(3344) <= not(inputs(169));
    layer0_outputs(3345) <= '1';
    layer0_outputs(3346) <= not(inputs(117)) or (inputs(249));
    layer0_outputs(3347) <= (inputs(111)) xor (inputs(96));
    layer0_outputs(3348) <= not((inputs(24)) xor (inputs(246)));
    layer0_outputs(3349) <= (inputs(159)) and not (inputs(219));
    layer0_outputs(3350) <= (inputs(79)) and not (inputs(249));
    layer0_outputs(3351) <= not((inputs(255)) xor (inputs(85)));
    layer0_outputs(3352) <= not((inputs(27)) xor (inputs(55)));
    layer0_outputs(3353) <= (inputs(25)) or (inputs(71));
    layer0_outputs(3354) <= inputs(217);
    layer0_outputs(3355) <= not((inputs(186)) or (inputs(123)));
    layer0_outputs(3356) <= (inputs(107)) or (inputs(2));
    layer0_outputs(3357) <= (inputs(21)) or (inputs(170));
    layer0_outputs(3358) <= (inputs(26)) and not (inputs(195));
    layer0_outputs(3359) <= (inputs(164)) and (inputs(86));
    layer0_outputs(3360) <= not(inputs(27));
    layer0_outputs(3361) <= (inputs(212)) or (inputs(39));
    layer0_outputs(3362) <= not((inputs(89)) or (inputs(77)));
    layer0_outputs(3363) <= not((inputs(212)) xor (inputs(88)));
    layer0_outputs(3364) <= not(inputs(197));
    layer0_outputs(3365) <= (inputs(188)) and not (inputs(95));
    layer0_outputs(3366) <= not((inputs(97)) or (inputs(173)));
    layer0_outputs(3367) <= not(inputs(59)) or (inputs(5));
    layer0_outputs(3368) <= not((inputs(70)) xor (inputs(87)));
    layer0_outputs(3369) <= not((inputs(38)) xor (inputs(104)));
    layer0_outputs(3370) <= not(inputs(173));
    layer0_outputs(3371) <= (inputs(50)) or (inputs(121));
    layer0_outputs(3372) <= (inputs(146)) and not (inputs(226));
    layer0_outputs(3373) <= (inputs(133)) or (inputs(177));
    layer0_outputs(3374) <= (inputs(48)) and (inputs(223));
    layer0_outputs(3375) <= not(inputs(68));
    layer0_outputs(3376) <= (inputs(134)) and not (inputs(8));
    layer0_outputs(3377) <= (inputs(84)) or (inputs(82));
    layer0_outputs(3378) <= not(inputs(215)) or (inputs(80));
    layer0_outputs(3379) <= (inputs(223)) and not (inputs(43));
    layer0_outputs(3380) <= inputs(244);
    layer0_outputs(3381) <= not(inputs(52)) or (inputs(129));
    layer0_outputs(3382) <= (inputs(98)) or (inputs(123));
    layer0_outputs(3383) <= inputs(43);
    layer0_outputs(3384) <= (inputs(185)) xor (inputs(51));
    layer0_outputs(3385) <= not(inputs(192)) or (inputs(207));
    layer0_outputs(3386) <= (inputs(5)) xor (inputs(112));
    layer0_outputs(3387) <= not(inputs(43)) or (inputs(19));
    layer0_outputs(3388) <= not(inputs(205));
    layer0_outputs(3389) <= (inputs(48)) and not (inputs(83));
    layer0_outputs(3390) <= (inputs(171)) and not (inputs(124));
    layer0_outputs(3391) <= (inputs(49)) xor (inputs(116));
    layer0_outputs(3392) <= not(inputs(99)) or (inputs(227));
    layer0_outputs(3393) <= not((inputs(249)) xor (inputs(121)));
    layer0_outputs(3394) <= not(inputs(58)) or (inputs(126));
    layer0_outputs(3395) <= not(inputs(163));
    layer0_outputs(3396) <= not((inputs(198)) or (inputs(143)));
    layer0_outputs(3397) <= not((inputs(243)) or (inputs(92)));
    layer0_outputs(3398) <= not(inputs(67)) or (inputs(246));
    layer0_outputs(3399) <= (inputs(124)) or (inputs(82));
    layer0_outputs(3400) <= (inputs(186)) or (inputs(36));
    layer0_outputs(3401) <= (inputs(132)) or (inputs(36));
    layer0_outputs(3402) <= (inputs(68)) or (inputs(170));
    layer0_outputs(3403) <= not(inputs(135));
    layer0_outputs(3404) <= not(inputs(136));
    layer0_outputs(3405) <= not((inputs(120)) xor (inputs(109)));
    layer0_outputs(3406) <= '1';
    layer0_outputs(3407) <= not((inputs(130)) and (inputs(3)));
    layer0_outputs(3408) <= not(inputs(122));
    layer0_outputs(3409) <= inputs(24);
    layer0_outputs(3410) <= inputs(120);
    layer0_outputs(3411) <= not(inputs(232)) or (inputs(111));
    layer0_outputs(3412) <= (inputs(74)) xor (inputs(87));
    layer0_outputs(3413) <= (inputs(8)) and (inputs(186));
    layer0_outputs(3414) <= not((inputs(116)) xor (inputs(43)));
    layer0_outputs(3415) <= not(inputs(196));
    layer0_outputs(3416) <= inputs(90);
    layer0_outputs(3417) <= inputs(136);
    layer0_outputs(3418) <= not((inputs(67)) or (inputs(172)));
    layer0_outputs(3419) <= (inputs(121)) or (inputs(62));
    layer0_outputs(3420) <= (inputs(158)) xor (inputs(53));
    layer0_outputs(3421) <= not((inputs(39)) or (inputs(243)));
    layer0_outputs(3422) <= '1';
    layer0_outputs(3423) <= '1';
    layer0_outputs(3424) <= (inputs(116)) and not (inputs(97));
    layer0_outputs(3425) <= inputs(124);
    layer0_outputs(3426) <= not(inputs(8)) or (inputs(222));
    layer0_outputs(3427) <= (inputs(14)) or (inputs(211));
    layer0_outputs(3428) <= (inputs(103)) and not (inputs(77));
    layer0_outputs(3429) <= not((inputs(79)) and (inputs(65)));
    layer0_outputs(3430) <= not(inputs(155));
    layer0_outputs(3431) <= (inputs(225)) and (inputs(60));
    layer0_outputs(3432) <= not(inputs(57));
    layer0_outputs(3433) <= not(inputs(120)) or (inputs(118));
    layer0_outputs(3434) <= (inputs(53)) and not (inputs(23));
    layer0_outputs(3435) <= not(inputs(111)) or (inputs(112));
    layer0_outputs(3436) <= (inputs(92)) and not (inputs(207));
    layer0_outputs(3437) <= not((inputs(187)) xor (inputs(96)));
    layer0_outputs(3438) <= (inputs(71)) xor (inputs(130));
    layer0_outputs(3439) <= not(inputs(80)) or (inputs(146));
    layer0_outputs(3440) <= not(inputs(22));
    layer0_outputs(3441) <= not(inputs(19)) or (inputs(15));
    layer0_outputs(3442) <= not(inputs(165));
    layer0_outputs(3443) <= not((inputs(132)) xor (inputs(211)));
    layer0_outputs(3444) <= (inputs(112)) or (inputs(225));
    layer0_outputs(3445) <= inputs(31);
    layer0_outputs(3446) <= not(inputs(230));
    layer0_outputs(3447) <= not(inputs(56));
    layer0_outputs(3448) <= (inputs(237)) or (inputs(87));
    layer0_outputs(3449) <= '0';
    layer0_outputs(3450) <= inputs(34);
    layer0_outputs(3451) <= (inputs(122)) or (inputs(4));
    layer0_outputs(3452) <= '1';
    layer0_outputs(3453) <= (inputs(162)) or (inputs(143));
    layer0_outputs(3454) <= not((inputs(137)) or (inputs(153)));
    layer0_outputs(3455) <= not(inputs(138));
    layer0_outputs(3456) <= not(inputs(163)) or (inputs(45));
    layer0_outputs(3457) <= '0';
    layer0_outputs(3458) <= not((inputs(171)) or (inputs(178)));
    layer0_outputs(3459) <= (inputs(187)) or (inputs(165));
    layer0_outputs(3460) <= not((inputs(224)) and (inputs(80)));
    layer0_outputs(3461) <= inputs(41);
    layer0_outputs(3462) <= (inputs(134)) and not (inputs(123));
    layer0_outputs(3463) <= not(inputs(108)) or (inputs(78));
    layer0_outputs(3464) <= not((inputs(206)) xor (inputs(246)));
    layer0_outputs(3465) <= not((inputs(0)) or (inputs(71)));
    layer0_outputs(3466) <= not(inputs(105));
    layer0_outputs(3467) <= not((inputs(167)) or (inputs(142)));
    layer0_outputs(3468) <= not(inputs(15));
    layer0_outputs(3469) <= (inputs(186)) xor (inputs(90));
    layer0_outputs(3470) <= (inputs(16)) or (inputs(59));
    layer0_outputs(3471) <= not(inputs(143));
    layer0_outputs(3472) <= not(inputs(164));
    layer0_outputs(3473) <= not(inputs(43));
    layer0_outputs(3474) <= not((inputs(103)) and (inputs(120)));
    layer0_outputs(3475) <= inputs(38);
    layer0_outputs(3476) <= (inputs(57)) and not (inputs(115));
    layer0_outputs(3477) <= not(inputs(186)) or (inputs(19));
    layer0_outputs(3478) <= not((inputs(140)) xor (inputs(48)));
    layer0_outputs(3479) <= (inputs(82)) and not (inputs(178));
    layer0_outputs(3480) <= (inputs(160)) or (inputs(50));
    layer0_outputs(3481) <= not(inputs(138)) or (inputs(90));
    layer0_outputs(3482) <= not((inputs(255)) or (inputs(4)));
    layer0_outputs(3483) <= not(inputs(26)) or (inputs(227));
    layer0_outputs(3484) <= (inputs(70)) xor (inputs(47));
    layer0_outputs(3485) <= not(inputs(169)) or (inputs(255));
    layer0_outputs(3486) <= not((inputs(220)) xor (inputs(232)));
    layer0_outputs(3487) <= not((inputs(3)) and (inputs(98)));
    layer0_outputs(3488) <= not((inputs(51)) and (inputs(29)));
    layer0_outputs(3489) <= not(inputs(53));
    layer0_outputs(3490) <= (inputs(32)) or (inputs(217));
    layer0_outputs(3491) <= inputs(116);
    layer0_outputs(3492) <= not(inputs(150)) or (inputs(161));
    layer0_outputs(3493) <= not(inputs(231));
    layer0_outputs(3494) <= not(inputs(0));
    layer0_outputs(3495) <= (inputs(24)) or (inputs(33));
    layer0_outputs(3496) <= (inputs(191)) and not (inputs(145));
    layer0_outputs(3497) <= (inputs(33)) or (inputs(187));
    layer0_outputs(3498) <= not((inputs(238)) or (inputs(107)));
    layer0_outputs(3499) <= (inputs(141)) xor (inputs(25));
    layer0_outputs(3500) <= inputs(100);
    layer0_outputs(3501) <= not(inputs(140));
    layer0_outputs(3502) <= inputs(76);
    layer0_outputs(3503) <= (inputs(69)) and (inputs(18));
    layer0_outputs(3504) <= not((inputs(162)) or (inputs(233)));
    layer0_outputs(3505) <= not(inputs(24)) or (inputs(89));
    layer0_outputs(3506) <= (inputs(70)) and not (inputs(233));
    layer0_outputs(3507) <= not((inputs(156)) xor (inputs(126)));
    layer0_outputs(3508) <= not(inputs(139));
    layer0_outputs(3509) <= not((inputs(163)) xor (inputs(84)));
    layer0_outputs(3510) <= inputs(71);
    layer0_outputs(3511) <= not(inputs(56));
    layer0_outputs(3512) <= not(inputs(55));
    layer0_outputs(3513) <= not(inputs(183)) or (inputs(66));
    layer0_outputs(3514) <= not((inputs(226)) or (inputs(93)));
    layer0_outputs(3515) <= inputs(132);
    layer0_outputs(3516) <= (inputs(67)) and not (inputs(195));
    layer0_outputs(3517) <= not((inputs(83)) xor (inputs(152)));
    layer0_outputs(3518) <= (inputs(154)) and not (inputs(230));
    layer0_outputs(3519) <= (inputs(80)) and (inputs(208));
    layer0_outputs(3520) <= not(inputs(74));
    layer0_outputs(3521) <= (inputs(252)) xor (inputs(26));
    layer0_outputs(3522) <= not(inputs(214)) or (inputs(159));
    layer0_outputs(3523) <= not((inputs(89)) or (inputs(219)));
    layer0_outputs(3524) <= (inputs(15)) and not (inputs(174));
    layer0_outputs(3525) <= inputs(72);
    layer0_outputs(3526) <= (inputs(200)) and not (inputs(233));
    layer0_outputs(3527) <= (inputs(30)) and (inputs(11));
    layer0_outputs(3528) <= (inputs(92)) or (inputs(228));
    layer0_outputs(3529) <= not((inputs(22)) xor (inputs(165)));
    layer0_outputs(3530) <= not(inputs(92)) or (inputs(252));
    layer0_outputs(3531) <= not((inputs(175)) and (inputs(184)));
    layer0_outputs(3532) <= not(inputs(89));
    layer0_outputs(3533) <= not(inputs(153));
    layer0_outputs(3534) <= not(inputs(135)) or (inputs(85));
    layer0_outputs(3535) <= inputs(121);
    layer0_outputs(3536) <= not(inputs(30)) or (inputs(145));
    layer0_outputs(3537) <= (inputs(155)) and not (inputs(16));
    layer0_outputs(3538) <= not((inputs(144)) xor (inputs(118)));
    layer0_outputs(3539) <= (inputs(138)) and not (inputs(147));
    layer0_outputs(3540) <= not((inputs(68)) and (inputs(193)));
    layer0_outputs(3541) <= not((inputs(246)) or (inputs(78)));
    layer0_outputs(3542) <= (inputs(100)) or (inputs(77));
    layer0_outputs(3543) <= (inputs(210)) xor (inputs(82));
    layer0_outputs(3544) <= (inputs(139)) and not (inputs(171));
    layer0_outputs(3545) <= not((inputs(27)) or (inputs(177)));
    layer0_outputs(3546) <= not(inputs(182)) or (inputs(95));
    layer0_outputs(3547) <= (inputs(105)) and not (inputs(198));
    layer0_outputs(3548) <= (inputs(251)) xor (inputs(29));
    layer0_outputs(3549) <= not(inputs(201));
    layer0_outputs(3550) <= not((inputs(85)) or (inputs(132)));
    layer0_outputs(3551) <= '0';
    layer0_outputs(3552) <= not(inputs(3)) or (inputs(6));
    layer0_outputs(3553) <= not((inputs(26)) and (inputs(97)));
    layer0_outputs(3554) <= (inputs(214)) or (inputs(194));
    layer0_outputs(3555) <= not((inputs(182)) or (inputs(39)));
    layer0_outputs(3556) <= not((inputs(106)) or (inputs(28)));
    layer0_outputs(3557) <= not((inputs(63)) or (inputs(107)));
    layer0_outputs(3558) <= not(inputs(232));
    layer0_outputs(3559) <= not(inputs(27)) or (inputs(176));
    layer0_outputs(3560) <= not((inputs(165)) and (inputs(196)));
    layer0_outputs(3561) <= inputs(215);
    layer0_outputs(3562) <= (inputs(2)) or (inputs(212));
    layer0_outputs(3563) <= (inputs(153)) and not (inputs(23));
    layer0_outputs(3564) <= (inputs(251)) xor (inputs(170));
    layer0_outputs(3565) <= (inputs(161)) and not (inputs(43));
    layer0_outputs(3566) <= '0';
    layer0_outputs(3567) <= not((inputs(63)) xor (inputs(135)));
    layer0_outputs(3568) <= '0';
    layer0_outputs(3569) <= (inputs(120)) or (inputs(46));
    layer0_outputs(3570) <= inputs(99);
    layer0_outputs(3571) <= (inputs(99)) or (inputs(12));
    layer0_outputs(3572) <= (inputs(169)) or (inputs(162));
    layer0_outputs(3573) <= not((inputs(219)) or (inputs(122)));
    layer0_outputs(3574) <= not(inputs(60)) or (inputs(83));
    layer0_outputs(3575) <= not(inputs(91));
    layer0_outputs(3576) <= not((inputs(177)) or (inputs(69)));
    layer0_outputs(3577) <= '0';
    layer0_outputs(3578) <= '0';
    layer0_outputs(3579) <= not((inputs(27)) xor (inputs(102)));
    layer0_outputs(3580) <= not((inputs(129)) xor (inputs(2)));
    layer0_outputs(3581) <= inputs(119);
    layer0_outputs(3582) <= not(inputs(190));
    layer0_outputs(3583) <= not(inputs(181));
    layer0_outputs(3584) <= not((inputs(207)) xor (inputs(123)));
    layer0_outputs(3585) <= (inputs(143)) or (inputs(100));
    layer0_outputs(3586) <= not(inputs(116)) or (inputs(46));
    layer0_outputs(3587) <= (inputs(190)) xor (inputs(254));
    layer0_outputs(3588) <= not((inputs(11)) and (inputs(35)));
    layer0_outputs(3589) <= (inputs(154)) or (inputs(108));
    layer0_outputs(3590) <= '1';
    layer0_outputs(3591) <= not((inputs(170)) and (inputs(85)));
    layer0_outputs(3592) <= (inputs(222)) and not (inputs(81));
    layer0_outputs(3593) <= (inputs(34)) xor (inputs(239));
    layer0_outputs(3594) <= not((inputs(35)) xor (inputs(114)));
    layer0_outputs(3595) <= '0';
    layer0_outputs(3596) <= not(inputs(205));
    layer0_outputs(3597) <= (inputs(185)) or (inputs(161));
    layer0_outputs(3598) <= not(inputs(74)) or (inputs(207));
    layer0_outputs(3599) <= not(inputs(101));
    layer0_outputs(3600) <= not((inputs(175)) xor (inputs(181)));
    layer0_outputs(3601) <= not(inputs(122));
    layer0_outputs(3602) <= inputs(101);
    layer0_outputs(3603) <= (inputs(99)) or (inputs(48));
    layer0_outputs(3604) <= (inputs(76)) or (inputs(216));
    layer0_outputs(3605) <= (inputs(48)) or (inputs(188));
    layer0_outputs(3606) <= (inputs(116)) and not (inputs(233));
    layer0_outputs(3607) <= (inputs(130)) or (inputs(231));
    layer0_outputs(3608) <= not(inputs(152));
    layer0_outputs(3609) <= (inputs(53)) and not (inputs(12));
    layer0_outputs(3610) <= not((inputs(65)) and (inputs(247)));
    layer0_outputs(3611) <= (inputs(68)) and not (inputs(28));
    layer0_outputs(3612) <= (inputs(129)) xor (inputs(169));
    layer0_outputs(3613) <= not((inputs(51)) xor (inputs(236)));
    layer0_outputs(3614) <= not((inputs(104)) xor (inputs(126)));
    layer0_outputs(3615) <= inputs(255);
    layer0_outputs(3616) <= not((inputs(225)) xor (inputs(162)));
    layer0_outputs(3617) <= inputs(33);
    layer0_outputs(3618) <= inputs(121);
    layer0_outputs(3619) <= not((inputs(114)) or (inputs(218)));
    layer0_outputs(3620) <= (inputs(63)) xor (inputs(185));
    layer0_outputs(3621) <= (inputs(237)) or (inputs(2));
    layer0_outputs(3622) <= not((inputs(0)) xor (inputs(205)));
    layer0_outputs(3623) <= (inputs(180)) and not (inputs(143));
    layer0_outputs(3624) <= not(inputs(141)) or (inputs(52));
    layer0_outputs(3625) <= (inputs(57)) and not (inputs(253));
    layer0_outputs(3626) <= (inputs(44)) or (inputs(52));
    layer0_outputs(3627) <= not(inputs(172));
    layer0_outputs(3628) <= not((inputs(118)) xor (inputs(126)));
    layer0_outputs(3629) <= not(inputs(45)) or (inputs(234));
    layer0_outputs(3630) <= not(inputs(215)) or (inputs(150));
    layer0_outputs(3631) <= not(inputs(177));
    layer0_outputs(3632) <= '0';
    layer0_outputs(3633) <= inputs(115);
    layer0_outputs(3634) <= '1';
    layer0_outputs(3635) <= (inputs(9)) and not (inputs(127));
    layer0_outputs(3636) <= (inputs(100)) or (inputs(109));
    layer0_outputs(3637) <= inputs(2);
    layer0_outputs(3638) <= (inputs(253)) and not (inputs(64));
    layer0_outputs(3639) <= (inputs(100)) and not (inputs(206));
    layer0_outputs(3640) <= inputs(101);
    layer0_outputs(3641) <= not(inputs(3));
    layer0_outputs(3642) <= (inputs(212)) xor (inputs(193));
    layer0_outputs(3643) <= (inputs(106)) or (inputs(99));
    layer0_outputs(3644) <= not(inputs(230));
    layer0_outputs(3645) <= not((inputs(74)) or (inputs(39)));
    layer0_outputs(3646) <= not((inputs(63)) xor (inputs(135)));
    layer0_outputs(3647) <= not(inputs(104)) or (inputs(148));
    layer0_outputs(3648) <= (inputs(88)) xor (inputs(76));
    layer0_outputs(3649) <= (inputs(80)) and (inputs(49));
    layer0_outputs(3650) <= (inputs(155)) and not (inputs(248));
    layer0_outputs(3651) <= not(inputs(117)) or (inputs(181));
    layer0_outputs(3652) <= not(inputs(22)) or (inputs(46));
    layer0_outputs(3653) <= not((inputs(49)) and (inputs(97)));
    layer0_outputs(3654) <= inputs(168);
    layer0_outputs(3655) <= (inputs(207)) or (inputs(88));
    layer0_outputs(3656) <= not(inputs(26)) or (inputs(95));
    layer0_outputs(3657) <= not(inputs(152)) or (inputs(158));
    layer0_outputs(3658) <= not((inputs(212)) xor (inputs(153)));
    layer0_outputs(3659) <= not(inputs(41));
    layer0_outputs(3660) <= (inputs(88)) or (inputs(73));
    layer0_outputs(3661) <= inputs(18);
    layer0_outputs(3662) <= inputs(123);
    layer0_outputs(3663) <= (inputs(157)) xor (inputs(207));
    layer0_outputs(3664) <= not(inputs(133));
    layer0_outputs(3665) <= not((inputs(210)) xor (inputs(162)));
    layer0_outputs(3666) <= (inputs(169)) xor (inputs(86));
    layer0_outputs(3667) <= (inputs(118)) or (inputs(246));
    layer0_outputs(3668) <= not((inputs(116)) or (inputs(128)));
    layer0_outputs(3669) <= (inputs(12)) xor (inputs(195));
    layer0_outputs(3670) <= (inputs(172)) and (inputs(158));
    layer0_outputs(3671) <= (inputs(80)) and not (inputs(30));
    layer0_outputs(3672) <= (inputs(85)) and not (inputs(204));
    layer0_outputs(3673) <= not((inputs(129)) or (inputs(98)));
    layer0_outputs(3674) <= inputs(150);
    layer0_outputs(3675) <= not((inputs(160)) or (inputs(195)));
    layer0_outputs(3676) <= (inputs(201)) and (inputs(70));
    layer0_outputs(3677) <= (inputs(16)) xor (inputs(160));
    layer0_outputs(3678) <= not(inputs(103));
    layer0_outputs(3679) <= not(inputs(221)) or (inputs(37));
    layer0_outputs(3680) <= (inputs(82)) xor (inputs(13));
    layer0_outputs(3681) <= not(inputs(150));
    layer0_outputs(3682) <= not(inputs(87));
    layer0_outputs(3683) <= not(inputs(154)) or (inputs(168));
    layer0_outputs(3684) <= not(inputs(196)) or (inputs(53));
    layer0_outputs(3685) <= not((inputs(5)) xor (inputs(71)));
    layer0_outputs(3686) <= not((inputs(59)) xor (inputs(180)));
    layer0_outputs(3687) <= not((inputs(72)) xor (inputs(127)));
    layer0_outputs(3688) <= '1';
    layer0_outputs(3689) <= not(inputs(39));
    layer0_outputs(3690) <= inputs(114);
    layer0_outputs(3691) <= (inputs(255)) and not (inputs(79));
    layer0_outputs(3692) <= not(inputs(125));
    layer0_outputs(3693) <= not(inputs(5));
    layer0_outputs(3694) <= (inputs(198)) and (inputs(151));
    layer0_outputs(3695) <= inputs(173);
    layer0_outputs(3696) <= (inputs(242)) and not (inputs(129));
    layer0_outputs(3697) <= (inputs(3)) and (inputs(96));
    layer0_outputs(3698) <= not(inputs(27));
    layer0_outputs(3699) <= not(inputs(29));
    layer0_outputs(3700) <= not((inputs(200)) or (inputs(77)));
    layer0_outputs(3701) <= inputs(242);
    layer0_outputs(3702) <= (inputs(1)) and not (inputs(210));
    layer0_outputs(3703) <= not((inputs(224)) and (inputs(53)));
    layer0_outputs(3704) <= (inputs(59)) and not (inputs(223));
    layer0_outputs(3705) <= inputs(103);
    layer0_outputs(3706) <= not((inputs(42)) or (inputs(178)));
    layer0_outputs(3707) <= (inputs(114)) or (inputs(176));
    layer0_outputs(3708) <= (inputs(168)) or (inputs(127));
    layer0_outputs(3709) <= not(inputs(218)) or (inputs(48));
    layer0_outputs(3710) <= (inputs(100)) or (inputs(198));
    layer0_outputs(3711) <= '1';
    layer0_outputs(3712) <= not(inputs(218)) or (inputs(83));
    layer0_outputs(3713) <= (inputs(74)) or (inputs(215));
    layer0_outputs(3714) <= (inputs(104)) or (inputs(34));
    layer0_outputs(3715) <= '1';
    layer0_outputs(3716) <= not(inputs(130)) or (inputs(131));
    layer0_outputs(3717) <= inputs(71);
    layer0_outputs(3718) <= (inputs(90)) and not (inputs(96));
    layer0_outputs(3719) <= (inputs(102)) or (inputs(111));
    layer0_outputs(3720) <= inputs(152);
    layer0_outputs(3721) <= inputs(172);
    layer0_outputs(3722) <= inputs(173);
    layer0_outputs(3723) <= (inputs(240)) or (inputs(215));
    layer0_outputs(3724) <= (inputs(170)) xor (inputs(97));
    layer0_outputs(3725) <= (inputs(105)) and not (inputs(230));
    layer0_outputs(3726) <= not(inputs(198)) or (inputs(15));
    layer0_outputs(3727) <= not((inputs(81)) xor (inputs(110)));
    layer0_outputs(3728) <= '1';
    layer0_outputs(3729) <= '0';
    layer0_outputs(3730) <= inputs(39);
    layer0_outputs(3731) <= not((inputs(51)) or (inputs(153)));
    layer0_outputs(3732) <= (inputs(54)) and not (inputs(60));
    layer0_outputs(3733) <= (inputs(56)) and not (inputs(98));
    layer0_outputs(3734) <= (inputs(144)) and not (inputs(216));
    layer0_outputs(3735) <= inputs(233);
    layer0_outputs(3736) <= not(inputs(167)) or (inputs(103));
    layer0_outputs(3737) <= not((inputs(92)) xor (inputs(9)));
    layer0_outputs(3738) <= (inputs(248)) or (inputs(101));
    layer0_outputs(3739) <= not(inputs(41));
    layer0_outputs(3740) <= (inputs(109)) xor (inputs(248));
    layer0_outputs(3741) <= (inputs(174)) and not (inputs(193));
    layer0_outputs(3742) <= not(inputs(31)) or (inputs(229));
    layer0_outputs(3743) <= (inputs(30)) xor (inputs(197));
    layer0_outputs(3744) <= not((inputs(121)) or (inputs(160)));
    layer0_outputs(3745) <= not((inputs(219)) and (inputs(220)));
    layer0_outputs(3746) <= (inputs(107)) or (inputs(214));
    layer0_outputs(3747) <= inputs(218);
    layer0_outputs(3748) <= not(inputs(89)) or (inputs(121));
    layer0_outputs(3749) <= (inputs(128)) and (inputs(218));
    layer0_outputs(3750) <= inputs(166);
    layer0_outputs(3751) <= (inputs(205)) or (inputs(98));
    layer0_outputs(3752) <= not(inputs(77));
    layer0_outputs(3753) <= (inputs(106)) xor (inputs(140));
    layer0_outputs(3754) <= not((inputs(122)) xor (inputs(68)));
    layer0_outputs(3755) <= not((inputs(56)) xor (inputs(187)));
    layer0_outputs(3756) <= not(inputs(243)) or (inputs(231));
    layer0_outputs(3757) <= (inputs(235)) and not (inputs(241));
    layer0_outputs(3758) <= not((inputs(213)) xor (inputs(217)));
    layer0_outputs(3759) <= not(inputs(106));
    layer0_outputs(3760) <= (inputs(25)) and not (inputs(28));
    layer0_outputs(3761) <= not((inputs(155)) xor (inputs(242)));
    layer0_outputs(3762) <= not(inputs(154)) or (inputs(24));
    layer0_outputs(3763) <= inputs(156);
    layer0_outputs(3764) <= not(inputs(214));
    layer0_outputs(3765) <= (inputs(171)) and not (inputs(224));
    layer0_outputs(3766) <= not((inputs(143)) xor (inputs(79)));
    layer0_outputs(3767) <= (inputs(75)) and not (inputs(138));
    layer0_outputs(3768) <= not((inputs(29)) or (inputs(167)));
    layer0_outputs(3769) <= inputs(81);
    layer0_outputs(3770) <= (inputs(114)) xor (inputs(80));
    layer0_outputs(3771) <= (inputs(52)) and not (inputs(238));
    layer0_outputs(3772) <= (inputs(69)) or (inputs(20));
    layer0_outputs(3773) <= not((inputs(25)) or (inputs(44)));
    layer0_outputs(3774) <= not((inputs(37)) and (inputs(185)));
    layer0_outputs(3775) <= not((inputs(122)) or (inputs(10)));
    layer0_outputs(3776) <= not(inputs(183)) or (inputs(87));
    layer0_outputs(3777) <= not((inputs(102)) xor (inputs(116)));
    layer0_outputs(3778) <= not(inputs(164)) or (inputs(87));
    layer0_outputs(3779) <= not((inputs(139)) or (inputs(226)));
    layer0_outputs(3780) <= (inputs(115)) and (inputs(112));
    layer0_outputs(3781) <= not((inputs(121)) xor (inputs(220)));
    layer0_outputs(3782) <= not((inputs(49)) or (inputs(215)));
    layer0_outputs(3783) <= (inputs(116)) xor (inputs(74));
    layer0_outputs(3784) <= (inputs(2)) and not (inputs(220));
    layer0_outputs(3785) <= inputs(213);
    layer0_outputs(3786) <= not((inputs(35)) and (inputs(178)));
    layer0_outputs(3787) <= (inputs(179)) and not (inputs(244));
    layer0_outputs(3788) <= inputs(121);
    layer0_outputs(3789) <= (inputs(125)) xor (inputs(245));
    layer0_outputs(3790) <= not(inputs(158)) or (inputs(222));
    layer0_outputs(3791) <= not((inputs(244)) and (inputs(239)));
    layer0_outputs(3792) <= (inputs(39)) or (inputs(72));
    layer0_outputs(3793) <= not(inputs(150)) or (inputs(174));
    layer0_outputs(3794) <= (inputs(206)) xor (inputs(166));
    layer0_outputs(3795) <= not(inputs(153));
    layer0_outputs(3796) <= inputs(196);
    layer0_outputs(3797) <= inputs(208);
    layer0_outputs(3798) <= not(inputs(173));
    layer0_outputs(3799) <= not((inputs(33)) xor (inputs(180)));
    layer0_outputs(3800) <= (inputs(54)) and not (inputs(146));
    layer0_outputs(3801) <= not(inputs(53));
    layer0_outputs(3802) <= not((inputs(124)) or (inputs(113)));
    layer0_outputs(3803) <= inputs(119);
    layer0_outputs(3804) <= (inputs(250)) or (inputs(242));
    layer0_outputs(3805) <= (inputs(130)) or (inputs(66));
    layer0_outputs(3806) <= not((inputs(160)) xor (inputs(94)));
    layer0_outputs(3807) <= not(inputs(89)) or (inputs(228));
    layer0_outputs(3808) <= not(inputs(123)) or (inputs(110));
    layer0_outputs(3809) <= inputs(52);
    layer0_outputs(3810) <= (inputs(101)) xor (inputs(219));
    layer0_outputs(3811) <= not(inputs(36)) or (inputs(225));
    layer0_outputs(3812) <= inputs(92);
    layer0_outputs(3813) <= (inputs(111)) xor (inputs(56));
    layer0_outputs(3814) <= (inputs(169)) xor (inputs(237));
    layer0_outputs(3815) <= (inputs(152)) and not (inputs(232));
    layer0_outputs(3816) <= not(inputs(147));
    layer0_outputs(3817) <= (inputs(73)) and not (inputs(44));
    layer0_outputs(3818) <= '1';
    layer0_outputs(3819) <= (inputs(6)) and (inputs(169));
    layer0_outputs(3820) <= (inputs(88)) and (inputs(20));
    layer0_outputs(3821) <= not((inputs(230)) xor (inputs(214)));
    layer0_outputs(3822) <= not((inputs(82)) xor (inputs(76)));
    layer0_outputs(3823) <= (inputs(105)) and not (inputs(164));
    layer0_outputs(3824) <= not(inputs(40)) or (inputs(70));
    layer0_outputs(3825) <= (inputs(251)) xor (inputs(75));
    layer0_outputs(3826) <= (inputs(18)) xor (inputs(249));
    layer0_outputs(3827) <= (inputs(2)) and not (inputs(173));
    layer0_outputs(3828) <= (inputs(230)) or (inputs(190));
    layer0_outputs(3829) <= not(inputs(154)) or (inputs(228));
    layer0_outputs(3830) <= not((inputs(179)) or (inputs(209)));
    layer0_outputs(3831) <= not(inputs(71)) or (inputs(117));
    layer0_outputs(3832) <= not((inputs(180)) or (inputs(214)));
    layer0_outputs(3833) <= not((inputs(40)) xor (inputs(255)));
    layer0_outputs(3834) <= (inputs(118)) or (inputs(252));
    layer0_outputs(3835) <= (inputs(74)) and (inputs(195));
    layer0_outputs(3836) <= inputs(115);
    layer0_outputs(3837) <= (inputs(225)) and not (inputs(112));
    layer0_outputs(3838) <= not(inputs(165));
    layer0_outputs(3839) <= inputs(68);
    layer0_outputs(3840) <= (inputs(6)) and not (inputs(191));
    layer0_outputs(3841) <= not(inputs(119)) or (inputs(239));
    layer0_outputs(3842) <= not(inputs(91)) or (inputs(222));
    layer0_outputs(3843) <= (inputs(225)) or (inputs(105));
    layer0_outputs(3844) <= not((inputs(186)) xor (inputs(4)));
    layer0_outputs(3845) <= not((inputs(80)) xor (inputs(217)));
    layer0_outputs(3846) <= (inputs(41)) and (inputs(165));
    layer0_outputs(3847) <= not(inputs(223)) or (inputs(18));
    layer0_outputs(3848) <= (inputs(157)) xor (inputs(103));
    layer0_outputs(3849) <= inputs(188);
    layer0_outputs(3850) <= (inputs(252)) and (inputs(50));
    layer0_outputs(3851) <= not(inputs(118));
    layer0_outputs(3852) <= inputs(195);
    layer0_outputs(3853) <= (inputs(137)) or (inputs(230));
    layer0_outputs(3854) <= inputs(161);
    layer0_outputs(3855) <= not(inputs(2)) or (inputs(229));
    layer0_outputs(3856) <= not((inputs(4)) and (inputs(53)));
    layer0_outputs(3857) <= not((inputs(171)) or (inputs(66)));
    layer0_outputs(3858) <= not((inputs(182)) xor (inputs(9)));
    layer0_outputs(3859) <= (inputs(172)) or (inputs(198));
    layer0_outputs(3860) <= (inputs(101)) and not (inputs(44));
    layer0_outputs(3861) <= not((inputs(205)) xor (inputs(4)));
    layer0_outputs(3862) <= not(inputs(187));
    layer0_outputs(3863) <= (inputs(153)) or (inputs(253));
    layer0_outputs(3864) <= not(inputs(133)) or (inputs(178));
    layer0_outputs(3865) <= not(inputs(184));
    layer0_outputs(3866) <= not((inputs(87)) or (inputs(142)));
    layer0_outputs(3867) <= not((inputs(227)) xor (inputs(228)));
    layer0_outputs(3868) <= '0';
    layer0_outputs(3869) <= (inputs(244)) xor (inputs(65));
    layer0_outputs(3870) <= (inputs(103)) and not (inputs(69));
    layer0_outputs(3871) <= (inputs(197)) and not (inputs(141));
    layer0_outputs(3872) <= not(inputs(168));
    layer0_outputs(3873) <= (inputs(212)) and not (inputs(255));
    layer0_outputs(3874) <= inputs(225);
    layer0_outputs(3875) <= not(inputs(133)) or (inputs(202));
    layer0_outputs(3876) <= not((inputs(109)) or (inputs(222)));
    layer0_outputs(3877) <= not(inputs(246)) or (inputs(192));
    layer0_outputs(3878) <= not(inputs(173)) or (inputs(81));
    layer0_outputs(3879) <= not((inputs(75)) and (inputs(75)));
    layer0_outputs(3880) <= (inputs(54)) or (inputs(197));
    layer0_outputs(3881) <= not(inputs(111)) or (inputs(25));
    layer0_outputs(3882) <= not((inputs(96)) or (inputs(76)));
    layer0_outputs(3883) <= not((inputs(210)) xor (inputs(162)));
    layer0_outputs(3884) <= (inputs(233)) or (inputs(115));
    layer0_outputs(3885) <= (inputs(140)) and not (inputs(129));
    layer0_outputs(3886) <= (inputs(70)) and not (inputs(238));
    layer0_outputs(3887) <= (inputs(76)) and not (inputs(204));
    layer0_outputs(3888) <= not((inputs(4)) xor (inputs(215)));
    layer0_outputs(3889) <= not((inputs(56)) or (inputs(240)));
    layer0_outputs(3890) <= (inputs(94)) or (inputs(201));
    layer0_outputs(3891) <= not(inputs(255)) or (inputs(175));
    layer0_outputs(3892) <= (inputs(39)) xor (inputs(11));
    layer0_outputs(3893) <= (inputs(40)) or (inputs(26));
    layer0_outputs(3894) <= not((inputs(244)) and (inputs(27)));
    layer0_outputs(3895) <= not(inputs(113)) or (inputs(67));
    layer0_outputs(3896) <= not(inputs(202));
    layer0_outputs(3897) <= (inputs(143)) xor (inputs(130));
    layer0_outputs(3898) <= (inputs(213)) xor (inputs(145));
    layer0_outputs(3899) <= inputs(134);
    layer0_outputs(3900) <= not((inputs(209)) and (inputs(21)));
    layer0_outputs(3901) <= inputs(61);
    layer0_outputs(3902) <= (inputs(202)) xor (inputs(153));
    layer0_outputs(3903) <= not((inputs(61)) or (inputs(95)));
    layer0_outputs(3904) <= not(inputs(32)) or (inputs(37));
    layer0_outputs(3905) <= not((inputs(133)) xor (inputs(102)));
    layer0_outputs(3906) <= not(inputs(175));
    layer0_outputs(3907) <= not((inputs(66)) or (inputs(184)));
    layer0_outputs(3908) <= not(inputs(168)) or (inputs(22));
    layer0_outputs(3909) <= not((inputs(238)) and (inputs(251)));
    layer0_outputs(3910) <= '0';
    layer0_outputs(3911) <= not(inputs(34)) or (inputs(158));
    layer0_outputs(3912) <= (inputs(245)) xor (inputs(113));
    layer0_outputs(3913) <= (inputs(140)) or (inputs(241));
    layer0_outputs(3914) <= not(inputs(187));
    layer0_outputs(3915) <= (inputs(108)) and not (inputs(174));
    layer0_outputs(3916) <= (inputs(81)) and not (inputs(16));
    layer0_outputs(3917) <= not(inputs(84));
    layer0_outputs(3918) <= inputs(44);
    layer0_outputs(3919) <= (inputs(191)) or (inputs(194));
    layer0_outputs(3920) <= not(inputs(105)) or (inputs(245));
    layer0_outputs(3921) <= not(inputs(219)) or (inputs(86));
    layer0_outputs(3922) <= (inputs(205)) and not (inputs(98));
    layer0_outputs(3923) <= not((inputs(203)) or (inputs(169)));
    layer0_outputs(3924) <= inputs(152);
    layer0_outputs(3925) <= (inputs(150)) xor (inputs(96));
    layer0_outputs(3926) <= not((inputs(136)) xor (inputs(142)));
    layer0_outputs(3927) <= not(inputs(46));
    layer0_outputs(3928) <= not((inputs(57)) xor (inputs(66)));
    layer0_outputs(3929) <= (inputs(181)) and not (inputs(32));
    layer0_outputs(3930) <= (inputs(140)) and not (inputs(46));
    layer0_outputs(3931) <= not(inputs(119));
    layer0_outputs(3932) <= not(inputs(21)) or (inputs(49));
    layer0_outputs(3933) <= not(inputs(138));
    layer0_outputs(3934) <= not(inputs(141)) or (inputs(193));
    layer0_outputs(3935) <= not(inputs(76));
    layer0_outputs(3936) <= not(inputs(203));
    layer0_outputs(3937) <= (inputs(118)) and not (inputs(65));
    layer0_outputs(3938) <= not(inputs(206));
    layer0_outputs(3939) <= (inputs(72)) and not (inputs(147));
    layer0_outputs(3940) <= not(inputs(45));
    layer0_outputs(3941) <= (inputs(107)) and not (inputs(38));
    layer0_outputs(3942) <= (inputs(190)) or (inputs(156));
    layer0_outputs(3943) <= (inputs(119)) and not (inputs(126));
    layer0_outputs(3944) <= not((inputs(114)) xor (inputs(67)));
    layer0_outputs(3945) <= '0';
    layer0_outputs(3946) <= (inputs(90)) xor (inputs(187));
    layer0_outputs(3947) <= (inputs(121)) xor (inputs(203));
    layer0_outputs(3948) <= not(inputs(67));
    layer0_outputs(3949) <= not((inputs(111)) and (inputs(212)));
    layer0_outputs(3950) <= (inputs(120)) xor (inputs(11));
    layer0_outputs(3951) <= inputs(15);
    layer0_outputs(3952) <= (inputs(48)) xor (inputs(211));
    layer0_outputs(3953) <= not((inputs(46)) or (inputs(132)));
    layer0_outputs(3954) <= (inputs(116)) and not (inputs(251));
    layer0_outputs(3955) <= (inputs(223)) or (inputs(58));
    layer0_outputs(3956) <= (inputs(207)) and not (inputs(47));
    layer0_outputs(3957) <= not(inputs(61));
    layer0_outputs(3958) <= not((inputs(38)) xor (inputs(249)));
    layer0_outputs(3959) <= (inputs(58)) xor (inputs(196));
    layer0_outputs(3960) <= (inputs(246)) xor (inputs(246));
    layer0_outputs(3961) <= not((inputs(241)) and (inputs(5)));
    layer0_outputs(3962) <= not((inputs(248)) or (inputs(173)));
    layer0_outputs(3963) <= (inputs(51)) xor (inputs(58));
    layer0_outputs(3964) <= not((inputs(44)) xor (inputs(100)));
    layer0_outputs(3965) <= (inputs(204)) and not (inputs(128));
    layer0_outputs(3966) <= not(inputs(102));
    layer0_outputs(3967) <= not(inputs(164));
    layer0_outputs(3968) <= (inputs(128)) and not (inputs(122));
    layer0_outputs(3969) <= not(inputs(141));
    layer0_outputs(3970) <= not(inputs(105));
    layer0_outputs(3971) <= (inputs(115)) and not (inputs(38));
    layer0_outputs(3972) <= inputs(204);
    layer0_outputs(3973) <= not((inputs(81)) xor (inputs(3)));
    layer0_outputs(3974) <= (inputs(185)) and (inputs(23));
    layer0_outputs(3975) <= not(inputs(151));
    layer0_outputs(3976) <= not((inputs(14)) and (inputs(240)));
    layer0_outputs(3977) <= not((inputs(85)) xor (inputs(51)));
    layer0_outputs(3978) <= (inputs(8)) or (inputs(217));
    layer0_outputs(3979) <= (inputs(137)) or (inputs(24));
    layer0_outputs(3980) <= (inputs(41)) and not (inputs(92));
    layer0_outputs(3981) <= (inputs(186)) or (inputs(188));
    layer0_outputs(3982) <= (inputs(56)) and not (inputs(26));
    layer0_outputs(3983) <= not((inputs(132)) and (inputs(147)));
    layer0_outputs(3984) <= inputs(138);
    layer0_outputs(3985) <= (inputs(34)) and not (inputs(249));
    layer0_outputs(3986) <= (inputs(170)) and (inputs(178));
    layer0_outputs(3987) <= inputs(91);
    layer0_outputs(3988) <= not((inputs(89)) and (inputs(254)));
    layer0_outputs(3989) <= not(inputs(124));
    layer0_outputs(3990) <= (inputs(231)) or (inputs(51));
    layer0_outputs(3991) <= not(inputs(151)) or (inputs(78));
    layer0_outputs(3992) <= '1';
    layer0_outputs(3993) <= (inputs(20)) and (inputs(84));
    layer0_outputs(3994) <= not(inputs(25));
    layer0_outputs(3995) <= inputs(43);
    layer0_outputs(3996) <= not((inputs(131)) and (inputs(114)));
    layer0_outputs(3997) <= (inputs(212)) xor (inputs(220));
    layer0_outputs(3998) <= not(inputs(204)) or (inputs(124));
    layer0_outputs(3999) <= not(inputs(194)) or (inputs(77));
    layer0_outputs(4000) <= not(inputs(200)) or (inputs(230));
    layer0_outputs(4001) <= inputs(132);
    layer0_outputs(4002) <= not(inputs(124));
    layer0_outputs(4003) <= (inputs(102)) or (inputs(44));
    layer0_outputs(4004) <= not(inputs(2));
    layer0_outputs(4005) <= (inputs(207)) or (inputs(60));
    layer0_outputs(4006) <= not((inputs(51)) or (inputs(238)));
    layer0_outputs(4007) <= (inputs(150)) or (inputs(224));
    layer0_outputs(4008) <= (inputs(188)) and not (inputs(7));
    layer0_outputs(4009) <= not(inputs(168)) or (inputs(187));
    layer0_outputs(4010) <= (inputs(75)) and not (inputs(28));
    layer0_outputs(4011) <= not(inputs(142)) or (inputs(96));
    layer0_outputs(4012) <= not(inputs(219));
    layer0_outputs(4013) <= not((inputs(157)) xor (inputs(17)));
    layer0_outputs(4014) <= not((inputs(62)) or (inputs(29)));
    layer0_outputs(4015) <= (inputs(147)) and not (inputs(208));
    layer0_outputs(4016) <= (inputs(87)) and not (inputs(11));
    layer0_outputs(4017) <= (inputs(67)) xor (inputs(1));
    layer0_outputs(4018) <= (inputs(42)) xor (inputs(177));
    layer0_outputs(4019) <= not((inputs(189)) xor (inputs(20)));
    layer0_outputs(4020) <= (inputs(235)) xor (inputs(7));
    layer0_outputs(4021) <= (inputs(78)) and not (inputs(159));
    layer0_outputs(4022) <= not(inputs(161)) or (inputs(241));
    layer0_outputs(4023) <= not((inputs(229)) or (inputs(241)));
    layer0_outputs(4024) <= (inputs(190)) xor (inputs(69));
    layer0_outputs(4025) <= not(inputs(97)) or (inputs(29));
    layer0_outputs(4026) <= (inputs(186)) xor (inputs(74));
    layer0_outputs(4027) <= not(inputs(12)) or (inputs(175));
    layer0_outputs(4028) <= not((inputs(68)) or (inputs(37)));
    layer0_outputs(4029) <= (inputs(118)) and not (inputs(114));
    layer0_outputs(4030) <= not(inputs(195)) or (inputs(143));
    layer0_outputs(4031) <= inputs(106);
    layer0_outputs(4032) <= (inputs(27)) or (inputs(202));
    layer0_outputs(4033) <= not(inputs(84)) or (inputs(0));
    layer0_outputs(4034) <= not((inputs(138)) or (inputs(222)));
    layer0_outputs(4035) <= not(inputs(121)) or (inputs(240));
    layer0_outputs(4036) <= (inputs(25)) or (inputs(181));
    layer0_outputs(4037) <= not((inputs(102)) or (inputs(125)));
    layer0_outputs(4038) <= not(inputs(233));
    layer0_outputs(4039) <= inputs(135);
    layer0_outputs(4040) <= (inputs(184)) and not (inputs(65));
    layer0_outputs(4041) <= not(inputs(186)) or (inputs(131));
    layer0_outputs(4042) <= inputs(29);
    layer0_outputs(4043) <= (inputs(0)) and not (inputs(48));
    layer0_outputs(4044) <= (inputs(187)) and (inputs(223));
    layer0_outputs(4045) <= not((inputs(138)) xor (inputs(134)));
    layer0_outputs(4046) <= (inputs(49)) and (inputs(146));
    layer0_outputs(4047) <= not((inputs(175)) or (inputs(164)));
    layer0_outputs(4048) <= inputs(167);
    layer0_outputs(4049) <= not(inputs(255));
    layer0_outputs(4050) <= not(inputs(21)) or (inputs(255));
    layer0_outputs(4051) <= inputs(157);
    layer0_outputs(4052) <= '1';
    layer0_outputs(4053) <= not((inputs(74)) xor (inputs(253)));
    layer0_outputs(4054) <= (inputs(169)) and (inputs(173));
    layer0_outputs(4055) <= (inputs(220)) xor (inputs(44));
    layer0_outputs(4056) <= (inputs(56)) or (inputs(181));
    layer0_outputs(4057) <= not(inputs(152));
    layer0_outputs(4058) <= not(inputs(193));
    layer0_outputs(4059) <= not(inputs(169));
    layer0_outputs(4060) <= inputs(233);
    layer0_outputs(4061) <= '1';
    layer0_outputs(4062) <= not((inputs(86)) xor (inputs(213)));
    layer0_outputs(4063) <= not((inputs(243)) xor (inputs(10)));
    layer0_outputs(4064) <= (inputs(94)) and not (inputs(2));
    layer0_outputs(4065) <= (inputs(117)) xor (inputs(220));
    layer0_outputs(4066) <= not(inputs(58));
    layer0_outputs(4067) <= not(inputs(73)) or (inputs(141));
    layer0_outputs(4068) <= not(inputs(74));
    layer0_outputs(4069) <= not((inputs(101)) xor (inputs(224)));
    layer0_outputs(4070) <= not((inputs(224)) or (inputs(150)));
    layer0_outputs(4071) <= not(inputs(194)) or (inputs(76));
    layer0_outputs(4072) <= (inputs(120)) or (inputs(177));
    layer0_outputs(4073) <= inputs(69);
    layer0_outputs(4074) <= (inputs(75)) xor (inputs(154));
    layer0_outputs(4075) <= not((inputs(153)) or (inputs(246)));
    layer0_outputs(4076) <= not(inputs(167));
    layer0_outputs(4077) <= inputs(73);
    layer0_outputs(4078) <= (inputs(255)) xor (inputs(120));
    layer0_outputs(4079) <= '1';
    layer0_outputs(4080) <= (inputs(236)) and (inputs(49));
    layer0_outputs(4081) <= not((inputs(84)) xor (inputs(3)));
    layer0_outputs(4082) <= not((inputs(113)) or (inputs(167)));
    layer0_outputs(4083) <= not((inputs(90)) xor (inputs(247)));
    layer0_outputs(4084) <= not(inputs(216));
    layer0_outputs(4085) <= not(inputs(148));
    layer0_outputs(4086) <= not(inputs(162));
    layer0_outputs(4087) <= not(inputs(202));
    layer0_outputs(4088) <= (inputs(196)) or (inputs(145));
    layer0_outputs(4089) <= not(inputs(58)) or (inputs(215));
    layer0_outputs(4090) <= (inputs(233)) and not (inputs(192));
    layer0_outputs(4091) <= not((inputs(2)) xor (inputs(119)));
    layer0_outputs(4092) <= not((inputs(230)) xor (inputs(51)));
    layer0_outputs(4093) <= not((inputs(176)) or (inputs(167)));
    layer0_outputs(4094) <= not(inputs(221));
    layer0_outputs(4095) <= not(inputs(29));
    layer0_outputs(4096) <= not((inputs(187)) xor (inputs(67)));
    layer0_outputs(4097) <= not((inputs(95)) xor (inputs(204)));
    layer0_outputs(4098) <= not((inputs(220)) xor (inputs(38)));
    layer0_outputs(4099) <= inputs(73);
    layer0_outputs(4100) <= (inputs(233)) and not (inputs(245));
    layer0_outputs(4101) <= not((inputs(117)) or (inputs(21)));
    layer0_outputs(4102) <= (inputs(67)) xor (inputs(24));
    layer0_outputs(4103) <= not((inputs(90)) xor (inputs(245)));
    layer0_outputs(4104) <= inputs(72);
    layer0_outputs(4105) <= (inputs(148)) and not (inputs(14));
    layer0_outputs(4106) <= (inputs(3)) and not (inputs(10));
    layer0_outputs(4107) <= not((inputs(81)) or (inputs(37)));
    layer0_outputs(4108) <= (inputs(0)) or (inputs(141));
    layer0_outputs(4109) <= not((inputs(38)) or (inputs(187)));
    layer0_outputs(4110) <= '0';
    layer0_outputs(4111) <= not((inputs(245)) xor (inputs(153)));
    layer0_outputs(4112) <= (inputs(66)) xor (inputs(132));
    layer0_outputs(4113) <= not(inputs(132)) or (inputs(30));
    layer0_outputs(4114) <= (inputs(91)) and not (inputs(98));
    layer0_outputs(4115) <= (inputs(100)) and not (inputs(182));
    layer0_outputs(4116) <= inputs(119);
    layer0_outputs(4117) <= not((inputs(90)) or (inputs(219)));
    layer0_outputs(4118) <= not(inputs(42));
    layer0_outputs(4119) <= (inputs(151)) and not (inputs(216));
    layer0_outputs(4120) <= '1';
    layer0_outputs(4121) <= (inputs(7)) and not (inputs(12));
    layer0_outputs(4122) <= '0';
    layer0_outputs(4123) <= not((inputs(199)) xor (inputs(213)));
    layer0_outputs(4124) <= (inputs(252)) and (inputs(210));
    layer0_outputs(4125) <= (inputs(233)) or (inputs(81));
    layer0_outputs(4126) <= not(inputs(203)) or (inputs(123));
    layer0_outputs(4127) <= not((inputs(82)) xor (inputs(58)));
    layer0_outputs(4128) <= '0';
    layer0_outputs(4129) <= (inputs(131)) or (inputs(5));
    layer0_outputs(4130) <= not(inputs(119));
    layer0_outputs(4131) <= not((inputs(236)) or (inputs(208)));
    layer0_outputs(4132) <= inputs(178);
    layer0_outputs(4133) <= not(inputs(163));
    layer0_outputs(4134) <= (inputs(91)) xor (inputs(168));
    layer0_outputs(4135) <= not((inputs(110)) xor (inputs(245)));
    layer0_outputs(4136) <= not(inputs(177));
    layer0_outputs(4137) <= '0';
    layer0_outputs(4138) <= not(inputs(87)) or (inputs(4));
    layer0_outputs(4139) <= inputs(209);
    layer0_outputs(4140) <= inputs(90);
    layer0_outputs(4141) <= (inputs(185)) xor (inputs(115));
    layer0_outputs(4142) <= '1';
    layer0_outputs(4143) <= (inputs(98)) or (inputs(197));
    layer0_outputs(4144) <= (inputs(32)) and not (inputs(35));
    layer0_outputs(4145) <= '1';
    layer0_outputs(4146) <= (inputs(118)) or (inputs(163));
    layer0_outputs(4147) <= '1';
    layer0_outputs(4148) <= not(inputs(172)) or (inputs(97));
    layer0_outputs(4149) <= inputs(62);
    layer0_outputs(4150) <= (inputs(153)) and not (inputs(173));
    layer0_outputs(4151) <= not((inputs(253)) or (inputs(244)));
    layer0_outputs(4152) <= (inputs(151)) and not (inputs(100));
    layer0_outputs(4153) <= (inputs(68)) and not (inputs(192));
    layer0_outputs(4154) <= (inputs(59)) xor (inputs(32));
    layer0_outputs(4155) <= not(inputs(83)) or (inputs(171));
    layer0_outputs(4156) <= (inputs(107)) or (inputs(71));
    layer0_outputs(4157) <= (inputs(93)) or (inputs(19));
    layer0_outputs(4158) <= (inputs(248)) xor (inputs(140));
    layer0_outputs(4159) <= not(inputs(74));
    layer0_outputs(4160) <= (inputs(219)) and not (inputs(245));
    layer0_outputs(4161) <= (inputs(218)) xor (inputs(186));
    layer0_outputs(4162) <= (inputs(30)) and not (inputs(97));
    layer0_outputs(4163) <= not((inputs(46)) or (inputs(134)));
    layer0_outputs(4164) <= not(inputs(10));
    layer0_outputs(4165) <= not(inputs(37));
    layer0_outputs(4166) <= not(inputs(237));
    layer0_outputs(4167) <= not(inputs(89)) or (inputs(205));
    layer0_outputs(4168) <= inputs(176);
    layer0_outputs(4169) <= not(inputs(107)) or (inputs(178));
    layer0_outputs(4170) <= inputs(134);
    layer0_outputs(4171) <= (inputs(182)) and not (inputs(23));
    layer0_outputs(4172) <= '1';
    layer0_outputs(4173) <= (inputs(194)) xor (inputs(159));
    layer0_outputs(4174) <= not(inputs(178));
    layer0_outputs(4175) <= (inputs(128)) and not (inputs(147));
    layer0_outputs(4176) <= (inputs(156)) xor (inputs(136));
    layer0_outputs(4177) <= not((inputs(230)) or (inputs(236)));
    layer0_outputs(4178) <= not(inputs(44)) or (inputs(212));
    layer0_outputs(4179) <= not((inputs(62)) xor (inputs(118)));
    layer0_outputs(4180) <= inputs(210);
    layer0_outputs(4181) <= (inputs(70)) xor (inputs(174));
    layer0_outputs(4182) <= not(inputs(152)) or (inputs(208));
    layer0_outputs(4183) <= not(inputs(233)) or (inputs(12));
    layer0_outputs(4184) <= inputs(24);
    layer0_outputs(4185) <= not((inputs(90)) and (inputs(81)));
    layer0_outputs(4186) <= not(inputs(86)) or (inputs(61));
    layer0_outputs(4187) <= inputs(100);
    layer0_outputs(4188) <= not((inputs(221)) xor (inputs(164)));
    layer0_outputs(4189) <= (inputs(193)) or (inputs(223));
    layer0_outputs(4190) <= not((inputs(54)) or (inputs(134)));
    layer0_outputs(4191) <= not((inputs(12)) or (inputs(89)));
    layer0_outputs(4192) <= (inputs(103)) xor (inputs(25));
    layer0_outputs(4193) <= (inputs(121)) and not (inputs(246));
    layer0_outputs(4194) <= not(inputs(248)) or (inputs(157));
    layer0_outputs(4195) <= (inputs(176)) or (inputs(137));
    layer0_outputs(4196) <= (inputs(86)) or (inputs(95));
    layer0_outputs(4197) <= (inputs(25)) or (inputs(87));
    layer0_outputs(4198) <= not((inputs(29)) or (inputs(220)));
    layer0_outputs(4199) <= not((inputs(71)) or (inputs(24)));
    layer0_outputs(4200) <= not((inputs(74)) xor (inputs(252)));
    layer0_outputs(4201) <= (inputs(162)) xor (inputs(142));
    layer0_outputs(4202) <= (inputs(141)) or (inputs(51));
    layer0_outputs(4203) <= inputs(172);
    layer0_outputs(4204) <= not((inputs(238)) xor (inputs(42)));
    layer0_outputs(4205) <= not((inputs(110)) xor (inputs(144)));
    layer0_outputs(4206) <= not(inputs(232));
    layer0_outputs(4207) <= not((inputs(29)) xor (inputs(91)));
    layer0_outputs(4208) <= not(inputs(59));
    layer0_outputs(4209) <= not(inputs(104));
    layer0_outputs(4210) <= not(inputs(56));
    layer0_outputs(4211) <= inputs(213);
    layer0_outputs(4212) <= inputs(13);
    layer0_outputs(4213) <= '1';
    layer0_outputs(4214) <= not(inputs(3));
    layer0_outputs(4215) <= '1';
    layer0_outputs(4216) <= (inputs(143)) xor (inputs(127));
    layer0_outputs(4217) <= (inputs(239)) and not (inputs(22));
    layer0_outputs(4218) <= not(inputs(58)) or (inputs(217));
    layer0_outputs(4219) <= (inputs(194)) or (inputs(249));
    layer0_outputs(4220) <= not(inputs(197)) or (inputs(72));
    layer0_outputs(4221) <= (inputs(4)) xor (inputs(184));
    layer0_outputs(4222) <= not((inputs(97)) or (inputs(248)));
    layer0_outputs(4223) <= not(inputs(62)) or (inputs(37));
    layer0_outputs(4224) <= inputs(214);
    layer0_outputs(4225) <= inputs(193);
    layer0_outputs(4226) <= not(inputs(88)) or (inputs(1));
    layer0_outputs(4227) <= not(inputs(93));
    layer0_outputs(4228) <= not((inputs(145)) xor (inputs(212)));
    layer0_outputs(4229) <= not(inputs(108)) or (inputs(46));
    layer0_outputs(4230) <= not(inputs(17)) or (inputs(178));
    layer0_outputs(4231) <= '0';
    layer0_outputs(4232) <= (inputs(10)) xor (inputs(14));
    layer0_outputs(4233) <= not((inputs(5)) xor (inputs(54)));
    layer0_outputs(4234) <= (inputs(101)) xor (inputs(115));
    layer0_outputs(4235) <= (inputs(76)) or (inputs(52));
    layer0_outputs(4236) <= not(inputs(184));
    layer0_outputs(4237) <= (inputs(222)) or (inputs(239));
    layer0_outputs(4238) <= not(inputs(11));
    layer0_outputs(4239) <= (inputs(219)) and not (inputs(243));
    layer0_outputs(4240) <= not(inputs(151)) or (inputs(236));
    layer0_outputs(4241) <= (inputs(141)) and not (inputs(138));
    layer0_outputs(4242) <= not((inputs(28)) xor (inputs(149)));
    layer0_outputs(4243) <= (inputs(220)) and not (inputs(125));
    layer0_outputs(4244) <= not(inputs(224));
    layer0_outputs(4245) <= (inputs(147)) and not (inputs(238));
    layer0_outputs(4246) <= inputs(22);
    layer0_outputs(4247) <= (inputs(223)) xor (inputs(40));
    layer0_outputs(4248) <= inputs(246);
    layer0_outputs(4249) <= not(inputs(226)) or (inputs(222));
    layer0_outputs(4250) <= not((inputs(72)) or (inputs(110)));
    layer0_outputs(4251) <= not((inputs(167)) or (inputs(125)));
    layer0_outputs(4252) <= not(inputs(76)) or (inputs(150));
    layer0_outputs(4253) <= '1';
    layer0_outputs(4254) <= (inputs(55)) or (inputs(123));
    layer0_outputs(4255) <= '0';
    layer0_outputs(4256) <= (inputs(11)) xor (inputs(222));
    layer0_outputs(4257) <= not(inputs(116));
    layer0_outputs(4258) <= not(inputs(231));
    layer0_outputs(4259) <= (inputs(42)) and not (inputs(159));
    layer0_outputs(4260) <= inputs(88);
    layer0_outputs(4261) <= inputs(222);
    layer0_outputs(4262) <= (inputs(201)) and (inputs(21));
    layer0_outputs(4263) <= (inputs(210)) xor (inputs(67));
    layer0_outputs(4264) <= not(inputs(90)) or (inputs(49));
    layer0_outputs(4265) <= not(inputs(171));
    layer0_outputs(4266) <= not((inputs(37)) xor (inputs(86)));
    layer0_outputs(4267) <= '1';
    layer0_outputs(4268) <= not((inputs(76)) or (inputs(110)));
    layer0_outputs(4269) <= '0';
    layer0_outputs(4270) <= (inputs(173)) or (inputs(114));
    layer0_outputs(4271) <= (inputs(77)) and not (inputs(238));
    layer0_outputs(4272) <= not(inputs(103));
    layer0_outputs(4273) <= (inputs(72)) and not (inputs(47));
    layer0_outputs(4274) <= (inputs(91)) or (inputs(64));
    layer0_outputs(4275) <= (inputs(43)) xor (inputs(191));
    layer0_outputs(4276) <= inputs(8);
    layer0_outputs(4277) <= not((inputs(207)) and (inputs(128)));
    layer0_outputs(4278) <= not((inputs(82)) xor (inputs(35)));
    layer0_outputs(4279) <= '1';
    layer0_outputs(4280) <= not(inputs(59));
    layer0_outputs(4281) <= (inputs(96)) and not (inputs(99));
    layer0_outputs(4282) <= not(inputs(177)) or (inputs(252));
    layer0_outputs(4283) <= (inputs(91)) xor (inputs(179));
    layer0_outputs(4284) <= (inputs(93)) and not (inputs(247));
    layer0_outputs(4285) <= (inputs(133)) or (inputs(127));
    layer0_outputs(4286) <= inputs(145);
    layer0_outputs(4287) <= (inputs(62)) or (inputs(226));
    layer0_outputs(4288) <= not((inputs(8)) xor (inputs(202)));
    layer0_outputs(4289) <= not(inputs(216));
    layer0_outputs(4290) <= not(inputs(136));
    layer0_outputs(4291) <= '0';
    layer0_outputs(4292) <= not((inputs(123)) xor (inputs(106)));
    layer0_outputs(4293) <= (inputs(134)) xor (inputs(213));
    layer0_outputs(4294) <= (inputs(233)) or (inputs(39));
    layer0_outputs(4295) <= not((inputs(221)) or (inputs(203)));
    layer0_outputs(4296) <= inputs(115);
    layer0_outputs(4297) <= (inputs(141)) xor (inputs(255));
    layer0_outputs(4298) <= not(inputs(46));
    layer0_outputs(4299) <= inputs(62);
    layer0_outputs(4300) <= inputs(145);
    layer0_outputs(4301) <= not((inputs(209)) and (inputs(44)));
    layer0_outputs(4302) <= (inputs(214)) xor (inputs(251));
    layer0_outputs(4303) <= not(inputs(154)) or (inputs(143));
    layer0_outputs(4304) <= inputs(18);
    layer0_outputs(4305) <= (inputs(138)) or (inputs(141));
    layer0_outputs(4306) <= (inputs(145)) and (inputs(220));
    layer0_outputs(4307) <= not((inputs(104)) xor (inputs(162)));
    layer0_outputs(4308) <= '1';
    layer0_outputs(4309) <= (inputs(148)) xor (inputs(151));
    layer0_outputs(4310) <= inputs(89);
    layer0_outputs(4311) <= not(inputs(101)) or (inputs(156));
    layer0_outputs(4312) <= not(inputs(119));
    layer0_outputs(4313) <= inputs(151);
    layer0_outputs(4314) <= (inputs(230)) xor (inputs(128));
    layer0_outputs(4315) <= (inputs(42)) and not (inputs(203));
    layer0_outputs(4316) <= (inputs(117)) xor (inputs(255));
    layer0_outputs(4317) <= not((inputs(84)) xor (inputs(110)));
    layer0_outputs(4318) <= not(inputs(203)) or (inputs(223));
    layer0_outputs(4319) <= not((inputs(96)) and (inputs(146)));
    layer0_outputs(4320) <= not(inputs(148));
    layer0_outputs(4321) <= not(inputs(37)) or (inputs(19));
    layer0_outputs(4322) <= (inputs(97)) or (inputs(121));
    layer0_outputs(4323) <= inputs(141);
    layer0_outputs(4324) <= not((inputs(93)) or (inputs(61)));
    layer0_outputs(4325) <= not((inputs(111)) or (inputs(181)));
    layer0_outputs(4326) <= not(inputs(183)) or (inputs(162));
    layer0_outputs(4327) <= not((inputs(215)) or (inputs(146)));
    layer0_outputs(4328) <= not((inputs(216)) or (inputs(246)));
    layer0_outputs(4329) <= (inputs(78)) and not (inputs(30));
    layer0_outputs(4330) <= inputs(89);
    layer0_outputs(4331) <= not((inputs(208)) or (inputs(158)));
    layer0_outputs(4332) <= inputs(67);
    layer0_outputs(4333) <= not((inputs(241)) xor (inputs(64)));
    layer0_outputs(4334) <= (inputs(202)) or (inputs(212));
    layer0_outputs(4335) <= not(inputs(46)) or (inputs(20));
    layer0_outputs(4336) <= not((inputs(17)) or (inputs(202)));
    layer0_outputs(4337) <= (inputs(170)) and not (inputs(234));
    layer0_outputs(4338) <= not((inputs(20)) or (inputs(106)));
    layer0_outputs(4339) <= (inputs(224)) xor (inputs(4));
    layer0_outputs(4340) <= not(inputs(216));
    layer0_outputs(4341) <= inputs(106);
    layer0_outputs(4342) <= (inputs(171)) or (inputs(237));
    layer0_outputs(4343) <= (inputs(91)) and not (inputs(237));
    layer0_outputs(4344) <= (inputs(44)) or (inputs(227));
    layer0_outputs(4345) <= (inputs(6)) xor (inputs(235));
    layer0_outputs(4346) <= (inputs(166)) or (inputs(9));
    layer0_outputs(4347) <= (inputs(153)) or (inputs(78));
    layer0_outputs(4348) <= not(inputs(196));
    layer0_outputs(4349) <= not(inputs(183)) or (inputs(50));
    layer0_outputs(4350) <= inputs(133);
    layer0_outputs(4351) <= (inputs(193)) or (inputs(146));
    layer0_outputs(4352) <= not(inputs(203));
    layer0_outputs(4353) <= not((inputs(101)) xor (inputs(242)));
    layer0_outputs(4354) <= (inputs(1)) and not (inputs(248));
    layer0_outputs(4355) <= not(inputs(171)) or (inputs(64));
    layer0_outputs(4356) <= inputs(76);
    layer0_outputs(4357) <= (inputs(174)) and (inputs(238));
    layer0_outputs(4358) <= not((inputs(32)) or (inputs(197)));
    layer0_outputs(4359) <= not((inputs(1)) or (inputs(236)));
    layer0_outputs(4360) <= inputs(132);
    layer0_outputs(4361) <= not((inputs(63)) or (inputs(187)));
    layer0_outputs(4362) <= not(inputs(216));
    layer0_outputs(4363) <= (inputs(133)) and not (inputs(237));
    layer0_outputs(4364) <= (inputs(93)) or (inputs(55));
    layer0_outputs(4365) <= not(inputs(168)) or (inputs(162));
    layer0_outputs(4366) <= not((inputs(48)) xor (inputs(192)));
    layer0_outputs(4367) <= (inputs(57)) xor (inputs(26));
    layer0_outputs(4368) <= not((inputs(186)) or (inputs(116)));
    layer0_outputs(4369) <= not((inputs(191)) or (inputs(173)));
    layer0_outputs(4370) <= (inputs(123)) and not (inputs(238));
    layer0_outputs(4371) <= not(inputs(210));
    layer0_outputs(4372) <= '1';
    layer0_outputs(4373) <= not(inputs(26)) or (inputs(145));
    layer0_outputs(4374) <= '1';
    layer0_outputs(4375) <= not(inputs(78));
    layer0_outputs(4376) <= (inputs(134)) xor (inputs(124));
    layer0_outputs(4377) <= not(inputs(241)) or (inputs(207));
    layer0_outputs(4378) <= inputs(189);
    layer0_outputs(4379) <= (inputs(194)) xor (inputs(130));
    layer0_outputs(4380) <= '0';
    layer0_outputs(4381) <= (inputs(6)) and (inputs(219));
    layer0_outputs(4382) <= not(inputs(128)) or (inputs(130));
    layer0_outputs(4383) <= (inputs(74)) and not (inputs(194));
    layer0_outputs(4384) <= inputs(68);
    layer0_outputs(4385) <= not(inputs(182));
    layer0_outputs(4386) <= not(inputs(164));
    layer0_outputs(4387) <= '1';
    layer0_outputs(4388) <= not(inputs(56)) or (inputs(178));
    layer0_outputs(4389) <= not((inputs(40)) or (inputs(110)));
    layer0_outputs(4390) <= (inputs(48)) xor (inputs(32));
    layer0_outputs(4391) <= not(inputs(198));
    layer0_outputs(4392) <= not(inputs(132));
    layer0_outputs(4393) <= (inputs(0)) xor (inputs(180));
    layer0_outputs(4394) <= not((inputs(88)) or (inputs(114)));
    layer0_outputs(4395) <= (inputs(122)) xor (inputs(56));
    layer0_outputs(4396) <= not((inputs(18)) or (inputs(153)));
    layer0_outputs(4397) <= not((inputs(101)) or (inputs(2)));
    layer0_outputs(4398) <= not(inputs(166));
    layer0_outputs(4399) <= not((inputs(37)) or (inputs(89)));
    layer0_outputs(4400) <= inputs(210);
    layer0_outputs(4401) <= not(inputs(90));
    layer0_outputs(4402) <= (inputs(71)) xor (inputs(144));
    layer0_outputs(4403) <= not(inputs(108));
    layer0_outputs(4404) <= inputs(104);
    layer0_outputs(4405) <= inputs(119);
    layer0_outputs(4406) <= (inputs(100)) or (inputs(174));
    layer0_outputs(4407) <= (inputs(16)) and not (inputs(83));
    layer0_outputs(4408) <= inputs(163);
    layer0_outputs(4409) <= '0';
    layer0_outputs(4410) <= not(inputs(86));
    layer0_outputs(4411) <= not((inputs(104)) or (inputs(249)));
    layer0_outputs(4412) <= not((inputs(151)) or (inputs(130)));
    layer0_outputs(4413) <= not(inputs(199));
    layer0_outputs(4414) <= not(inputs(245)) or (inputs(104));
    layer0_outputs(4415) <= not((inputs(192)) or (inputs(225)));
    layer0_outputs(4416) <= (inputs(49)) or (inputs(124));
    layer0_outputs(4417) <= (inputs(152)) xor (inputs(222));
    layer0_outputs(4418) <= inputs(188);
    layer0_outputs(4419) <= not(inputs(135)) or (inputs(86));
    layer0_outputs(4420) <= not((inputs(70)) xor (inputs(55)));
    layer0_outputs(4421) <= (inputs(44)) or (inputs(153));
    layer0_outputs(4422) <= not(inputs(69));
    layer0_outputs(4423) <= not(inputs(226)) or (inputs(82));
    layer0_outputs(4424) <= not(inputs(110));
    layer0_outputs(4425) <= inputs(198);
    layer0_outputs(4426) <= inputs(132);
    layer0_outputs(4427) <= not(inputs(45)) or (inputs(165));
    layer0_outputs(4428) <= not((inputs(154)) or (inputs(252)));
    layer0_outputs(4429) <= '0';
    layer0_outputs(4430) <= (inputs(179)) and not (inputs(37));
    layer0_outputs(4431) <= inputs(30);
    layer0_outputs(4432) <= (inputs(55)) and not (inputs(139));
    layer0_outputs(4433) <= not(inputs(166)) or (inputs(233));
    layer0_outputs(4434) <= inputs(212);
    layer0_outputs(4435) <= (inputs(65)) xor (inputs(135));
    layer0_outputs(4436) <= (inputs(174)) xor (inputs(144));
    layer0_outputs(4437) <= not((inputs(243)) xor (inputs(72)));
    layer0_outputs(4438) <= not(inputs(215)) or (inputs(146));
    layer0_outputs(4439) <= not(inputs(174)) or (inputs(53));
    layer0_outputs(4440) <= (inputs(154)) or (inputs(150));
    layer0_outputs(4441) <= (inputs(178)) xor (inputs(143));
    layer0_outputs(4442) <= (inputs(152)) and not (inputs(159));
    layer0_outputs(4443) <= inputs(136);
    layer0_outputs(4444) <= (inputs(156)) or (inputs(154));
    layer0_outputs(4445) <= (inputs(199)) and not (inputs(146));
    layer0_outputs(4446) <= not(inputs(230));
    layer0_outputs(4447) <= '0';
    layer0_outputs(4448) <= '0';
    layer0_outputs(4449) <= not((inputs(239)) or (inputs(76)));
    layer0_outputs(4450) <= (inputs(242)) xor (inputs(251));
    layer0_outputs(4451) <= not(inputs(71)) or (inputs(161));
    layer0_outputs(4452) <= not((inputs(194)) or (inputs(178)));
    layer0_outputs(4453) <= not(inputs(196)) or (inputs(225));
    layer0_outputs(4454) <= '1';
    layer0_outputs(4455) <= (inputs(115)) or (inputs(238));
    layer0_outputs(4456) <= not(inputs(213));
    layer0_outputs(4457) <= (inputs(203)) and not (inputs(30));
    layer0_outputs(4458) <= not((inputs(29)) or (inputs(141)));
    layer0_outputs(4459) <= (inputs(114)) and not (inputs(225));
    layer0_outputs(4460) <= not((inputs(85)) or (inputs(248)));
    layer0_outputs(4461) <= not(inputs(229)) or (inputs(226));
    layer0_outputs(4462) <= not(inputs(147)) or (inputs(39));
    layer0_outputs(4463) <= not((inputs(45)) or (inputs(190)));
    layer0_outputs(4464) <= inputs(226);
    layer0_outputs(4465) <= not((inputs(104)) xor (inputs(157)));
    layer0_outputs(4466) <= (inputs(201)) or (inputs(240));
    layer0_outputs(4467) <= not(inputs(148));
    layer0_outputs(4468) <= inputs(179);
    layer0_outputs(4469) <= not((inputs(43)) or (inputs(111)));
    layer0_outputs(4470) <= inputs(216);
    layer0_outputs(4471) <= not((inputs(215)) or (inputs(103)));
    layer0_outputs(4472) <= '0';
    layer0_outputs(4473) <= (inputs(229)) or (inputs(46));
    layer0_outputs(4474) <= not((inputs(158)) or (inputs(134)));
    layer0_outputs(4475) <= not((inputs(74)) xor (inputs(72)));
    layer0_outputs(4476) <= not(inputs(137));
    layer0_outputs(4477) <= not((inputs(77)) xor (inputs(96)));
    layer0_outputs(4478) <= (inputs(75)) and not (inputs(228));
    layer0_outputs(4479) <= '0';
    layer0_outputs(4480) <= (inputs(75)) xor (inputs(99));
    layer0_outputs(4481) <= not(inputs(84));
    layer0_outputs(4482) <= inputs(199);
    layer0_outputs(4483) <= not(inputs(175));
    layer0_outputs(4484) <= inputs(218);
    layer0_outputs(4485) <= not(inputs(150));
    layer0_outputs(4486) <= not((inputs(133)) xor (inputs(128)));
    layer0_outputs(4487) <= (inputs(133)) and (inputs(164));
    layer0_outputs(4488) <= (inputs(56)) or (inputs(14));
    layer0_outputs(4489) <= (inputs(95)) and not (inputs(78));
    layer0_outputs(4490) <= not(inputs(199));
    layer0_outputs(4491) <= (inputs(76)) and not (inputs(123));
    layer0_outputs(4492) <= (inputs(182)) xor (inputs(245));
    layer0_outputs(4493) <= (inputs(216)) and (inputs(76));
    layer0_outputs(4494) <= inputs(55);
    layer0_outputs(4495) <= not((inputs(225)) xor (inputs(57)));
    layer0_outputs(4496) <= not((inputs(94)) or (inputs(201)));
    layer0_outputs(4497) <= not((inputs(184)) xor (inputs(13)));
    layer0_outputs(4498) <= (inputs(184)) and not (inputs(89));
    layer0_outputs(4499) <= (inputs(181)) and (inputs(11));
    layer0_outputs(4500) <= '1';
    layer0_outputs(4501) <= not(inputs(225)) or (inputs(84));
    layer0_outputs(4502) <= not(inputs(179)) or (inputs(131));
    layer0_outputs(4503) <= not((inputs(7)) or (inputs(201)));
    layer0_outputs(4504) <= not((inputs(34)) xor (inputs(153)));
    layer0_outputs(4505) <= not((inputs(203)) or (inputs(136)));
    layer0_outputs(4506) <= (inputs(57)) or (inputs(1));
    layer0_outputs(4507) <= not(inputs(166)) or (inputs(46));
    layer0_outputs(4508) <= (inputs(154)) xor (inputs(216));
    layer0_outputs(4509) <= '0';
    layer0_outputs(4510) <= (inputs(228)) xor (inputs(230));
    layer0_outputs(4511) <= not((inputs(21)) xor (inputs(158)));
    layer0_outputs(4512) <= inputs(180);
    layer0_outputs(4513) <= not((inputs(155)) or (inputs(156)));
    layer0_outputs(4514) <= (inputs(74)) xor (inputs(198));
    layer0_outputs(4515) <= not((inputs(141)) or (inputs(167)));
    layer0_outputs(4516) <= not(inputs(74));
    layer0_outputs(4517) <= not(inputs(146));
    layer0_outputs(4518) <= not((inputs(99)) or (inputs(18)));
    layer0_outputs(4519) <= (inputs(116)) or (inputs(20));
    layer0_outputs(4520) <= not(inputs(150));
    layer0_outputs(4521) <= (inputs(67)) and not (inputs(43));
    layer0_outputs(4522) <= not(inputs(180)) or (inputs(158));
    layer0_outputs(4523) <= not((inputs(210)) xor (inputs(225)));
    layer0_outputs(4524) <= not((inputs(19)) or (inputs(233)));
    layer0_outputs(4525) <= inputs(154);
    layer0_outputs(4526) <= not(inputs(118)) or (inputs(162));
    layer0_outputs(4527) <= not(inputs(102)) or (inputs(85));
    layer0_outputs(4528) <= (inputs(252)) xor (inputs(116));
    layer0_outputs(4529) <= (inputs(48)) and (inputs(141));
    layer0_outputs(4530) <= '0';
    layer0_outputs(4531) <= not(inputs(131));
    layer0_outputs(4532) <= not(inputs(92)) or (inputs(244));
    layer0_outputs(4533) <= not((inputs(36)) xor (inputs(11)));
    layer0_outputs(4534) <= (inputs(8)) xor (inputs(71));
    layer0_outputs(4535) <= (inputs(136)) and not (inputs(111));
    layer0_outputs(4536) <= '1';
    layer0_outputs(4537) <= (inputs(254)) and not (inputs(250));
    layer0_outputs(4538) <= not(inputs(44));
    layer0_outputs(4539) <= (inputs(201)) xor (inputs(170));
    layer0_outputs(4540) <= not(inputs(106)) or (inputs(205));
    layer0_outputs(4541) <= inputs(167);
    layer0_outputs(4542) <= not(inputs(122)) or (inputs(19));
    layer0_outputs(4543) <= not((inputs(58)) or (inputs(224)));
    layer0_outputs(4544) <= inputs(101);
    layer0_outputs(4545) <= '1';
    layer0_outputs(4546) <= (inputs(226)) xor (inputs(39));
    layer0_outputs(4547) <= not(inputs(72));
    layer0_outputs(4548) <= (inputs(143)) or (inputs(75));
    layer0_outputs(4549) <= (inputs(88)) and not (inputs(106));
    layer0_outputs(4550) <= not(inputs(135));
    layer0_outputs(4551) <= (inputs(36)) or (inputs(220));
    layer0_outputs(4552) <= (inputs(226)) and not (inputs(5));
    layer0_outputs(4553) <= not((inputs(214)) xor (inputs(51)));
    layer0_outputs(4554) <= not((inputs(91)) xor (inputs(236)));
    layer0_outputs(4555) <= not((inputs(42)) or (inputs(100)));
    layer0_outputs(4556) <= not(inputs(144)) or (inputs(161));
    layer0_outputs(4557) <= inputs(188);
    layer0_outputs(4558) <= not((inputs(110)) or (inputs(81)));
    layer0_outputs(4559) <= (inputs(190)) and not (inputs(239));
    layer0_outputs(4560) <= not(inputs(73)) or (inputs(165));
    layer0_outputs(4561) <= not(inputs(40)) or (inputs(239));
    layer0_outputs(4562) <= (inputs(198)) and not (inputs(27));
    layer0_outputs(4563) <= (inputs(86)) and not (inputs(164));
    layer0_outputs(4564) <= '1';
    layer0_outputs(4565) <= (inputs(5)) and not (inputs(187));
    layer0_outputs(4566) <= not((inputs(186)) xor (inputs(33)));
    layer0_outputs(4567) <= not((inputs(223)) xor (inputs(168)));
    layer0_outputs(4568) <= not((inputs(24)) or (inputs(157)));
    layer0_outputs(4569) <= not((inputs(64)) xor (inputs(75)));
    layer0_outputs(4570) <= '0';
    layer0_outputs(4571) <= (inputs(89)) and not (inputs(161));
    layer0_outputs(4572) <= (inputs(119)) xor (inputs(58));
    layer0_outputs(4573) <= not((inputs(71)) xor (inputs(94)));
    layer0_outputs(4574) <= '0';
    layer0_outputs(4575) <= inputs(52);
    layer0_outputs(4576) <= not(inputs(253)) or (inputs(19));
    layer0_outputs(4577) <= inputs(82);
    layer0_outputs(4578) <= inputs(195);
    layer0_outputs(4579) <= (inputs(181)) or (inputs(5));
    layer0_outputs(4580) <= (inputs(50)) or (inputs(1));
    layer0_outputs(4581) <= not(inputs(168)) or (inputs(108));
    layer0_outputs(4582) <= (inputs(228)) or (inputs(185));
    layer0_outputs(4583) <= (inputs(60)) xor (inputs(215));
    layer0_outputs(4584) <= not(inputs(108));
    layer0_outputs(4585) <= not(inputs(153));
    layer0_outputs(4586) <= not((inputs(19)) or (inputs(168)));
    layer0_outputs(4587) <= (inputs(146)) and not (inputs(129));
    layer0_outputs(4588) <= inputs(208);
    layer0_outputs(4589) <= not((inputs(240)) xor (inputs(124)));
    layer0_outputs(4590) <= (inputs(143)) xor (inputs(222));
    layer0_outputs(4591) <= not(inputs(139)) or (inputs(220));
    layer0_outputs(4592) <= (inputs(54)) and not (inputs(190));
    layer0_outputs(4593) <= (inputs(56)) xor (inputs(251));
    layer0_outputs(4594) <= '0';
    layer0_outputs(4595) <= not(inputs(162));
    layer0_outputs(4596) <= not(inputs(204));
    layer0_outputs(4597) <= (inputs(161)) or (inputs(180));
    layer0_outputs(4598) <= not((inputs(112)) or (inputs(218)));
    layer0_outputs(4599) <= (inputs(160)) xor (inputs(70));
    layer0_outputs(4600) <= not((inputs(43)) or (inputs(245)));
    layer0_outputs(4601) <= inputs(121);
    layer0_outputs(4602) <= not(inputs(162));
    layer0_outputs(4603) <= not((inputs(73)) or (inputs(57)));
    layer0_outputs(4604) <= (inputs(16)) or (inputs(71));
    layer0_outputs(4605) <= (inputs(19)) and not (inputs(30));
    layer0_outputs(4606) <= not((inputs(194)) or (inputs(50)));
    layer0_outputs(4607) <= not((inputs(63)) and (inputs(171)));
    layer0_outputs(4608) <= not((inputs(118)) or (inputs(232)));
    layer0_outputs(4609) <= (inputs(118)) xor (inputs(1));
    layer0_outputs(4610) <= not(inputs(128)) or (inputs(7));
    layer0_outputs(4611) <= inputs(185);
    layer0_outputs(4612) <= not((inputs(58)) xor (inputs(161)));
    layer0_outputs(4613) <= not(inputs(77));
    layer0_outputs(4614) <= (inputs(136)) and not (inputs(250));
    layer0_outputs(4615) <= inputs(87);
    layer0_outputs(4616) <= (inputs(99)) or (inputs(191));
    layer0_outputs(4617) <= (inputs(197)) xor (inputs(254));
    layer0_outputs(4618) <= not(inputs(198));
    layer0_outputs(4619) <= '0';
    layer0_outputs(4620) <= inputs(210);
    layer0_outputs(4621) <= (inputs(137)) or (inputs(113));
    layer0_outputs(4622) <= inputs(107);
    layer0_outputs(4623) <= (inputs(51)) xor (inputs(251));
    layer0_outputs(4624) <= (inputs(133)) and not (inputs(165));
    layer0_outputs(4625) <= inputs(124);
    layer0_outputs(4626) <= not(inputs(71));
    layer0_outputs(4627) <= (inputs(139)) or (inputs(129));
    layer0_outputs(4628) <= (inputs(126)) xor (inputs(132));
    layer0_outputs(4629) <= not((inputs(243)) xor (inputs(57)));
    layer0_outputs(4630) <= not((inputs(246)) or (inputs(25)));
    layer0_outputs(4631) <= not(inputs(153)) or (inputs(59));
    layer0_outputs(4632) <= (inputs(167)) and not (inputs(140));
    layer0_outputs(4633) <= (inputs(75)) or (inputs(58));
    layer0_outputs(4634) <= not(inputs(21)) or (inputs(170));
    layer0_outputs(4635) <= not(inputs(172));
    layer0_outputs(4636) <= not(inputs(197));
    layer0_outputs(4637) <= not((inputs(10)) xor (inputs(135)));
    layer0_outputs(4638) <= (inputs(94)) or (inputs(76));
    layer0_outputs(4639) <= not((inputs(161)) xor (inputs(73)));
    layer0_outputs(4640) <= (inputs(162)) or (inputs(243));
    layer0_outputs(4641) <= (inputs(27)) and not (inputs(222));
    layer0_outputs(4642) <= (inputs(89)) xor (inputs(241));
    layer0_outputs(4643) <= (inputs(158)) xor (inputs(84));
    layer0_outputs(4644) <= not(inputs(55)) or (inputs(226));
    layer0_outputs(4645) <= inputs(26);
    layer0_outputs(4646) <= not((inputs(135)) xor (inputs(105)));
    layer0_outputs(4647) <= not(inputs(229));
    layer0_outputs(4648) <= inputs(120);
    layer0_outputs(4649) <= (inputs(149)) and not (inputs(97));
    layer0_outputs(4650) <= (inputs(75)) or (inputs(70));
    layer0_outputs(4651) <= '0';
    layer0_outputs(4652) <= (inputs(134)) and not (inputs(178));
    layer0_outputs(4653) <= (inputs(231)) and (inputs(151));
    layer0_outputs(4654) <= not((inputs(41)) or (inputs(14)));
    layer0_outputs(4655) <= (inputs(132)) xor (inputs(13));
    layer0_outputs(4656) <= not(inputs(188)) or (inputs(231));
    layer0_outputs(4657) <= not((inputs(84)) xor (inputs(49)));
    layer0_outputs(4658) <= not(inputs(229)) or (inputs(31));
    layer0_outputs(4659) <= not(inputs(113));
    layer0_outputs(4660) <= not(inputs(220)) or (inputs(128));
    layer0_outputs(4661) <= (inputs(146)) or (inputs(56));
    layer0_outputs(4662) <= inputs(254);
    layer0_outputs(4663) <= not(inputs(99));
    layer0_outputs(4664) <= not(inputs(134));
    layer0_outputs(4665) <= inputs(93);
    layer0_outputs(4666) <= (inputs(98)) xor (inputs(139));
    layer0_outputs(4667) <= not((inputs(85)) or (inputs(42)));
    layer0_outputs(4668) <= not((inputs(199)) or (inputs(139)));
    layer0_outputs(4669) <= not((inputs(60)) or (inputs(31)));
    layer0_outputs(4670) <= (inputs(93)) and not (inputs(4));
    layer0_outputs(4671) <= not(inputs(240)) or (inputs(234));
    layer0_outputs(4672) <= not(inputs(165));
    layer0_outputs(4673) <= not(inputs(182));
    layer0_outputs(4674) <= inputs(176);
    layer0_outputs(4675) <= (inputs(233)) or (inputs(94));
    layer0_outputs(4676) <= (inputs(29)) xor (inputs(183));
    layer0_outputs(4677) <= (inputs(192)) xor (inputs(47));
    layer0_outputs(4678) <= inputs(141);
    layer0_outputs(4679) <= not((inputs(146)) xor (inputs(230)));
    layer0_outputs(4680) <= not(inputs(66));
    layer0_outputs(4681) <= (inputs(36)) xor (inputs(72));
    layer0_outputs(4682) <= inputs(171);
    layer0_outputs(4683) <= (inputs(175)) or (inputs(36));
    layer0_outputs(4684) <= (inputs(253)) and not (inputs(213));
    layer0_outputs(4685) <= not(inputs(183)) or (inputs(33));
    layer0_outputs(4686) <= not(inputs(173));
    layer0_outputs(4687) <= not(inputs(19));
    layer0_outputs(4688) <= (inputs(103)) xor (inputs(85));
    layer0_outputs(4689) <= (inputs(41)) xor (inputs(68));
    layer0_outputs(4690) <= not(inputs(92));
    layer0_outputs(4691) <= inputs(170);
    layer0_outputs(4692) <= not(inputs(10)) or (inputs(81));
    layer0_outputs(4693) <= not(inputs(164)) or (inputs(145));
    layer0_outputs(4694) <= inputs(49);
    layer0_outputs(4695) <= (inputs(243)) and not (inputs(127));
    layer0_outputs(4696) <= (inputs(210)) or (inputs(120));
    layer0_outputs(4697) <= not((inputs(85)) xor (inputs(176)));
    layer0_outputs(4698) <= inputs(164);
    layer0_outputs(4699) <= (inputs(202)) or (inputs(170));
    layer0_outputs(4700) <= (inputs(249)) xor (inputs(37));
    layer0_outputs(4701) <= (inputs(84)) and not (inputs(80));
    layer0_outputs(4702) <= '1';
    layer0_outputs(4703) <= (inputs(23)) or (inputs(124));
    layer0_outputs(4704) <= not((inputs(144)) or (inputs(148)));
    layer0_outputs(4705) <= not((inputs(32)) xor (inputs(197)));
    layer0_outputs(4706) <= not((inputs(89)) xor (inputs(114)));
    layer0_outputs(4707) <= inputs(80);
    layer0_outputs(4708) <= (inputs(128)) xor (inputs(84));
    layer0_outputs(4709) <= not(inputs(231));
    layer0_outputs(4710) <= not(inputs(61)) or (inputs(113));
    layer0_outputs(4711) <= not((inputs(227)) xor (inputs(115)));
    layer0_outputs(4712) <= not((inputs(8)) xor (inputs(79)));
    layer0_outputs(4713) <= not((inputs(105)) or (inputs(249)));
    layer0_outputs(4714) <= (inputs(175)) xor (inputs(105));
    layer0_outputs(4715) <= (inputs(150)) or (inputs(195));
    layer0_outputs(4716) <= not((inputs(34)) xor (inputs(151)));
    layer0_outputs(4717) <= (inputs(162)) or (inputs(232));
    layer0_outputs(4718) <= (inputs(96)) xor (inputs(143));
    layer0_outputs(4719) <= not(inputs(211)) or (inputs(159));
    layer0_outputs(4720) <= (inputs(101)) xor (inputs(2));
    layer0_outputs(4721) <= inputs(204);
    layer0_outputs(4722) <= not((inputs(208)) xor (inputs(7)));
    layer0_outputs(4723) <= not((inputs(198)) xor (inputs(228)));
    layer0_outputs(4724) <= not(inputs(84));
    layer0_outputs(4725) <= not((inputs(156)) xor (inputs(186)));
    layer0_outputs(4726) <= inputs(182);
    layer0_outputs(4727) <= not((inputs(72)) or (inputs(93)));
    layer0_outputs(4728) <= not(inputs(213));
    layer0_outputs(4729) <= not((inputs(28)) or (inputs(241)));
    layer0_outputs(4730) <= (inputs(237)) xor (inputs(22));
    layer0_outputs(4731) <= (inputs(196)) or (inputs(59));
    layer0_outputs(4732) <= (inputs(131)) xor (inputs(163));
    layer0_outputs(4733) <= not((inputs(151)) xor (inputs(244)));
    layer0_outputs(4734) <= not(inputs(95)) or (inputs(199));
    layer0_outputs(4735) <= inputs(99);
    layer0_outputs(4736) <= (inputs(139)) and not (inputs(252));
    layer0_outputs(4737) <= not((inputs(98)) xor (inputs(223)));
    layer0_outputs(4738) <= inputs(24);
    layer0_outputs(4739) <= not(inputs(115));
    layer0_outputs(4740) <= not(inputs(21)) or (inputs(218));
    layer0_outputs(4741) <= not(inputs(118));
    layer0_outputs(4742) <= (inputs(194)) xor (inputs(68));
    layer0_outputs(4743) <= not(inputs(244));
    layer0_outputs(4744) <= not((inputs(215)) xor (inputs(58)));
    layer0_outputs(4745) <= (inputs(0)) xor (inputs(33));
    layer0_outputs(4746) <= not((inputs(61)) or (inputs(65)));
    layer0_outputs(4747) <= (inputs(52)) xor (inputs(9));
    layer0_outputs(4748) <= '0';
    layer0_outputs(4749) <= not(inputs(232)) or (inputs(126));
    layer0_outputs(4750) <= (inputs(120)) xor (inputs(47));
    layer0_outputs(4751) <= inputs(118);
    layer0_outputs(4752) <= not((inputs(24)) xor (inputs(71)));
    layer0_outputs(4753) <= not((inputs(223)) xor (inputs(3)));
    layer0_outputs(4754) <= not(inputs(166));
    layer0_outputs(4755) <= inputs(242);
    layer0_outputs(4756) <= not((inputs(148)) xor (inputs(255)));
    layer0_outputs(4757) <= not((inputs(53)) and (inputs(142)));
    layer0_outputs(4758) <= not(inputs(190)) or (inputs(75));
    layer0_outputs(4759) <= not(inputs(171)) or (inputs(70));
    layer0_outputs(4760) <= not((inputs(44)) xor (inputs(254)));
    layer0_outputs(4761) <= not(inputs(186)) or (inputs(26));
    layer0_outputs(4762) <= not((inputs(22)) xor (inputs(38)));
    layer0_outputs(4763) <= (inputs(52)) xor (inputs(8));
    layer0_outputs(4764) <= (inputs(169)) xor (inputs(202));
    layer0_outputs(4765) <= '1';
    layer0_outputs(4766) <= not((inputs(127)) xor (inputs(163)));
    layer0_outputs(4767) <= not(inputs(117));
    layer0_outputs(4768) <= not((inputs(140)) or (inputs(249)));
    layer0_outputs(4769) <= not((inputs(176)) xor (inputs(74)));
    layer0_outputs(4770) <= not(inputs(198)) or (inputs(119));
    layer0_outputs(4771) <= inputs(203);
    layer0_outputs(4772) <= not(inputs(219));
    layer0_outputs(4773) <= not((inputs(188)) xor (inputs(62)));
    layer0_outputs(4774) <= (inputs(101)) or (inputs(215));
    layer0_outputs(4775) <= not((inputs(99)) or (inputs(21)));
    layer0_outputs(4776) <= '1';
    layer0_outputs(4777) <= (inputs(212)) or (inputs(220));
    layer0_outputs(4778) <= not((inputs(32)) xor (inputs(29)));
    layer0_outputs(4779) <= not((inputs(119)) or (inputs(162)));
    layer0_outputs(4780) <= (inputs(9)) and not (inputs(89));
    layer0_outputs(4781) <= not(inputs(234));
    layer0_outputs(4782) <= not((inputs(125)) or (inputs(245)));
    layer0_outputs(4783) <= (inputs(170)) xor (inputs(110));
    layer0_outputs(4784) <= '1';
    layer0_outputs(4785) <= not(inputs(103));
    layer0_outputs(4786) <= not((inputs(68)) xor (inputs(1)));
    layer0_outputs(4787) <= not((inputs(37)) or (inputs(185)));
    layer0_outputs(4788) <= not((inputs(15)) or (inputs(99)));
    layer0_outputs(4789) <= not((inputs(49)) xor (inputs(172)));
    layer0_outputs(4790) <= not(inputs(135));
    layer0_outputs(4791) <= '0';
    layer0_outputs(4792) <= not(inputs(173)) or (inputs(204));
    layer0_outputs(4793) <= not(inputs(147)) or (inputs(244));
    layer0_outputs(4794) <= (inputs(151)) or (inputs(252));
    layer0_outputs(4795) <= not(inputs(197));
    layer0_outputs(4796) <= not(inputs(176)) or (inputs(130));
    layer0_outputs(4797) <= not(inputs(107));
    layer0_outputs(4798) <= not((inputs(240)) xor (inputs(6)));
    layer0_outputs(4799) <= '0';
    layer0_outputs(4800) <= (inputs(8)) xor (inputs(38));
    layer0_outputs(4801) <= (inputs(165)) and not (inputs(81));
    layer0_outputs(4802) <= (inputs(56)) and not (inputs(119));
    layer0_outputs(4803) <= (inputs(46)) xor (inputs(48));
    layer0_outputs(4804) <= not(inputs(228));
    layer0_outputs(4805) <= not((inputs(137)) xor (inputs(3)));
    layer0_outputs(4806) <= (inputs(156)) and not (inputs(11));
    layer0_outputs(4807) <= inputs(121);
    layer0_outputs(4808) <= (inputs(185)) and not (inputs(114));
    layer0_outputs(4809) <= '1';
    layer0_outputs(4810) <= inputs(16);
    layer0_outputs(4811) <= (inputs(90)) and not (inputs(192));
    layer0_outputs(4812) <= (inputs(138)) xor (inputs(48));
    layer0_outputs(4813) <= (inputs(69)) or (inputs(188));
    layer0_outputs(4814) <= not(inputs(234));
    layer0_outputs(4815) <= inputs(102);
    layer0_outputs(4816) <= (inputs(94)) and not (inputs(221));
    layer0_outputs(4817) <= (inputs(135)) and not (inputs(131));
    layer0_outputs(4818) <= not(inputs(111));
    layer0_outputs(4819) <= (inputs(12)) and not (inputs(6));
    layer0_outputs(4820) <= not((inputs(10)) and (inputs(141)));
    layer0_outputs(4821) <= (inputs(163)) or (inputs(172));
    layer0_outputs(4822) <= not(inputs(72)) or (inputs(52));
    layer0_outputs(4823) <= inputs(107);
    layer0_outputs(4824) <= not(inputs(92));
    layer0_outputs(4825) <= (inputs(155)) and not (inputs(110));
    layer0_outputs(4826) <= not(inputs(252)) or (inputs(5));
    layer0_outputs(4827) <= (inputs(138)) or (inputs(118));
    layer0_outputs(4828) <= not((inputs(227)) or (inputs(99)));
    layer0_outputs(4829) <= (inputs(151)) or (inputs(22));
    layer0_outputs(4830) <= (inputs(69)) and not (inputs(11));
    layer0_outputs(4831) <= inputs(131);
    layer0_outputs(4832) <= (inputs(200)) and not (inputs(128));
    layer0_outputs(4833) <= (inputs(142)) or (inputs(136));
    layer0_outputs(4834) <= (inputs(220)) or (inputs(223));
    layer0_outputs(4835) <= (inputs(225)) xor (inputs(67));
    layer0_outputs(4836) <= not(inputs(82));
    layer0_outputs(4837) <= (inputs(146)) xor (inputs(175));
    layer0_outputs(4838) <= not((inputs(180)) or (inputs(96)));
    layer0_outputs(4839) <= (inputs(92)) and not (inputs(13));
    layer0_outputs(4840) <= inputs(221);
    layer0_outputs(4841) <= not((inputs(28)) xor (inputs(194)));
    layer0_outputs(4842) <= not((inputs(202)) or (inputs(248)));
    layer0_outputs(4843) <= (inputs(134)) and not (inputs(36));
    layer0_outputs(4844) <= not(inputs(165));
    layer0_outputs(4845) <= not(inputs(177)) or (inputs(184));
    layer0_outputs(4846) <= (inputs(211)) and not (inputs(47));
    layer0_outputs(4847) <= inputs(75);
    layer0_outputs(4848) <= inputs(71);
    layer0_outputs(4849) <= (inputs(173)) and not (inputs(254));
    layer0_outputs(4850) <= (inputs(135)) or (inputs(77));
    layer0_outputs(4851) <= (inputs(7)) xor (inputs(104));
    layer0_outputs(4852) <= not((inputs(202)) or (inputs(100)));
    layer0_outputs(4853) <= (inputs(234)) and (inputs(210));
    layer0_outputs(4854) <= inputs(27);
    layer0_outputs(4855) <= '1';
    layer0_outputs(4856) <= (inputs(204)) or (inputs(195));
    layer0_outputs(4857) <= (inputs(106)) or (inputs(238));
    layer0_outputs(4858) <= not(inputs(89));
    layer0_outputs(4859) <= not(inputs(16));
    layer0_outputs(4860) <= (inputs(106)) xor (inputs(131));
    layer0_outputs(4861) <= not(inputs(87));
    layer0_outputs(4862) <= inputs(125);
    layer0_outputs(4863) <= (inputs(201)) and (inputs(55));
    layer0_outputs(4864) <= not((inputs(200)) or (inputs(24)));
    layer0_outputs(4865) <= not(inputs(26)) or (inputs(2));
    layer0_outputs(4866) <= not(inputs(40));
    layer0_outputs(4867) <= '0';
    layer0_outputs(4868) <= (inputs(87)) xor (inputs(159));
    layer0_outputs(4869) <= (inputs(67)) and not (inputs(207));
    layer0_outputs(4870) <= not(inputs(217)) or (inputs(111));
    layer0_outputs(4871) <= not((inputs(198)) and (inputs(9)));
    layer0_outputs(4872) <= not(inputs(91));
    layer0_outputs(4873) <= not((inputs(213)) or (inputs(81)));
    layer0_outputs(4874) <= (inputs(186)) or (inputs(39));
    layer0_outputs(4875) <= not((inputs(255)) or (inputs(148)));
    layer0_outputs(4876) <= not(inputs(40)) or (inputs(252));
    layer0_outputs(4877) <= (inputs(229)) and not (inputs(193));
    layer0_outputs(4878) <= not(inputs(115)) or (inputs(37));
    layer0_outputs(4879) <= (inputs(199)) xor (inputs(168));
    layer0_outputs(4880) <= inputs(167);
    layer0_outputs(4881) <= inputs(131);
    layer0_outputs(4882) <= (inputs(186)) or (inputs(12));
    layer0_outputs(4883) <= not((inputs(212)) xor (inputs(188)));
    layer0_outputs(4884) <= not(inputs(135)) or (inputs(179));
    layer0_outputs(4885) <= not(inputs(183)) or (inputs(130));
    layer0_outputs(4886) <= (inputs(83)) xor (inputs(67));
    layer0_outputs(4887) <= not((inputs(7)) and (inputs(160)));
    layer0_outputs(4888) <= inputs(100);
    layer0_outputs(4889) <= inputs(123);
    layer0_outputs(4890) <= not((inputs(152)) or (inputs(176)));
    layer0_outputs(4891) <= inputs(209);
    layer0_outputs(4892) <= (inputs(86)) and not (inputs(10));
    layer0_outputs(4893) <= not((inputs(244)) and (inputs(77)));
    layer0_outputs(4894) <= not((inputs(101)) xor (inputs(73)));
    layer0_outputs(4895) <= not(inputs(229));
    layer0_outputs(4896) <= not((inputs(155)) or (inputs(7)));
    layer0_outputs(4897) <= not(inputs(253)) or (inputs(231));
    layer0_outputs(4898) <= (inputs(228)) and not (inputs(11));
    layer0_outputs(4899) <= not(inputs(184));
    layer0_outputs(4900) <= (inputs(80)) and not (inputs(9));
    layer0_outputs(4901) <= not((inputs(86)) or (inputs(199)));
    layer0_outputs(4902) <= (inputs(16)) and not (inputs(26));
    layer0_outputs(4903) <= not(inputs(154)) or (inputs(191));
    layer0_outputs(4904) <= not((inputs(240)) and (inputs(16)));
    layer0_outputs(4905) <= '0';
    layer0_outputs(4906) <= not((inputs(173)) or (inputs(60)));
    layer0_outputs(4907) <= not((inputs(98)) or (inputs(255)));
    layer0_outputs(4908) <= '0';
    layer0_outputs(4909) <= not(inputs(166));
    layer0_outputs(4910) <= (inputs(57)) xor (inputs(237));
    layer0_outputs(4911) <= inputs(40);
    layer0_outputs(4912) <= not(inputs(208)) or (inputs(19));
    layer0_outputs(4913) <= not(inputs(182));
    layer0_outputs(4914) <= not(inputs(65)) or (inputs(220));
    layer0_outputs(4915) <= inputs(60);
    layer0_outputs(4916) <= (inputs(71)) xor (inputs(192));
    layer0_outputs(4917) <= inputs(153);
    layer0_outputs(4918) <= '1';
    layer0_outputs(4919) <= (inputs(78)) xor (inputs(241));
    layer0_outputs(4920) <= (inputs(27)) or (inputs(231));
    layer0_outputs(4921) <= not(inputs(102)) or (inputs(227));
    layer0_outputs(4922) <= not((inputs(223)) or (inputs(22)));
    layer0_outputs(4923) <= (inputs(150)) and not (inputs(253));
    layer0_outputs(4924) <= (inputs(153)) and not (inputs(247));
    layer0_outputs(4925) <= inputs(41);
    layer0_outputs(4926) <= not((inputs(142)) and (inputs(246)));
    layer0_outputs(4927) <= inputs(19);
    layer0_outputs(4928) <= (inputs(176)) and (inputs(108));
    layer0_outputs(4929) <= not(inputs(182));
    layer0_outputs(4930) <= inputs(46);
    layer0_outputs(4931) <= '1';
    layer0_outputs(4932) <= not((inputs(87)) or (inputs(84)));
    layer0_outputs(4933) <= not(inputs(215)) or (inputs(253));
    layer0_outputs(4934) <= inputs(52);
    layer0_outputs(4935) <= not(inputs(103));
    layer0_outputs(4936) <= not((inputs(121)) and (inputs(159)));
    layer0_outputs(4937) <= not((inputs(22)) or (inputs(222)));
    layer0_outputs(4938) <= not(inputs(133));
    layer0_outputs(4939) <= not(inputs(212));
    layer0_outputs(4940) <= not((inputs(109)) xor (inputs(176)));
    layer0_outputs(4941) <= not(inputs(167)) or (inputs(154));
    layer0_outputs(4942) <= (inputs(237)) and not (inputs(149));
    layer0_outputs(4943) <= not(inputs(247));
    layer0_outputs(4944) <= inputs(195);
    layer0_outputs(4945) <= (inputs(146)) xor (inputs(89));
    layer0_outputs(4946) <= not((inputs(146)) or (inputs(161)));
    layer0_outputs(4947) <= inputs(232);
    layer0_outputs(4948) <= not((inputs(154)) xor (inputs(183)));
    layer0_outputs(4949) <= not(inputs(174));
    layer0_outputs(4950) <= (inputs(203)) or (inputs(121));
    layer0_outputs(4951) <= '1';
    layer0_outputs(4952) <= (inputs(94)) xor (inputs(172));
    layer0_outputs(4953) <= not((inputs(53)) or (inputs(37)));
    layer0_outputs(4954) <= (inputs(85)) and not (inputs(60));
    layer0_outputs(4955) <= inputs(230);
    layer0_outputs(4956) <= (inputs(44)) or (inputs(115));
    layer0_outputs(4957) <= not((inputs(21)) or (inputs(181)));
    layer0_outputs(4958) <= '0';
    layer0_outputs(4959) <= not(inputs(137)) or (inputs(42));
    layer0_outputs(4960) <= not((inputs(169)) or (inputs(122)));
    layer0_outputs(4961) <= not(inputs(135));
    layer0_outputs(4962) <= not((inputs(203)) or (inputs(210)));
    layer0_outputs(4963) <= inputs(171);
    layer0_outputs(4964) <= not(inputs(216)) or (inputs(208));
    layer0_outputs(4965) <= not(inputs(51));
    layer0_outputs(4966) <= '0';
    layer0_outputs(4967) <= not((inputs(117)) xor (inputs(30)));
    layer0_outputs(4968) <= '0';
    layer0_outputs(4969) <= not(inputs(250));
    layer0_outputs(4970) <= inputs(179);
    layer0_outputs(4971) <= '0';
    layer0_outputs(4972) <= (inputs(77)) xor (inputs(213));
    layer0_outputs(4973) <= not(inputs(217));
    layer0_outputs(4974) <= not((inputs(227)) and (inputs(5)));
    layer0_outputs(4975) <= not(inputs(148)) or (inputs(22));
    layer0_outputs(4976) <= (inputs(136)) and not (inputs(28));
    layer0_outputs(4977) <= not((inputs(57)) or (inputs(147)));
    layer0_outputs(4978) <= (inputs(115)) xor (inputs(8));
    layer0_outputs(4979) <= '0';
    layer0_outputs(4980) <= (inputs(53)) and not (inputs(48));
    layer0_outputs(4981) <= (inputs(75)) and not (inputs(171));
    layer0_outputs(4982) <= not((inputs(73)) xor (inputs(46)));
    layer0_outputs(4983) <= '0';
    layer0_outputs(4984) <= not(inputs(5)) or (inputs(16));
    layer0_outputs(4985) <= not((inputs(55)) xor (inputs(153)));
    layer0_outputs(4986) <= not(inputs(219)) or (inputs(64));
    layer0_outputs(4987) <= not((inputs(116)) or (inputs(142)));
    layer0_outputs(4988) <= (inputs(194)) xor (inputs(250));
    layer0_outputs(4989) <= not(inputs(71));
    layer0_outputs(4990) <= not(inputs(1)) or (inputs(228));
    layer0_outputs(4991) <= (inputs(88)) and not (inputs(115));
    layer0_outputs(4992) <= not(inputs(161));
    layer0_outputs(4993) <= (inputs(233)) and not (inputs(80));
    layer0_outputs(4994) <= not((inputs(138)) or (inputs(221)));
    layer0_outputs(4995) <= not(inputs(132)) or (inputs(227));
    layer0_outputs(4996) <= not(inputs(122));
    layer0_outputs(4997) <= not(inputs(92));
    layer0_outputs(4998) <= '0';
    layer0_outputs(4999) <= (inputs(233)) xor (inputs(74));
    layer0_outputs(5000) <= not(inputs(4));
    layer0_outputs(5001) <= not((inputs(180)) or (inputs(63)));
    layer0_outputs(5002) <= (inputs(122)) and not (inputs(166));
    layer0_outputs(5003) <= inputs(153);
    layer0_outputs(5004) <= (inputs(81)) and (inputs(143));
    layer0_outputs(5005) <= (inputs(54)) and not (inputs(82));
    layer0_outputs(5006) <= not(inputs(165)) or (inputs(139));
    layer0_outputs(5007) <= not(inputs(168));
    layer0_outputs(5008) <= not((inputs(28)) or (inputs(73)));
    layer0_outputs(5009) <= not((inputs(137)) xor (inputs(68)));
    layer0_outputs(5010) <= (inputs(37)) or (inputs(108));
    layer0_outputs(5011) <= '1';
    layer0_outputs(5012) <= (inputs(178)) xor (inputs(69));
    layer0_outputs(5013) <= not(inputs(110));
    layer0_outputs(5014) <= not(inputs(154)) or (inputs(61));
    layer0_outputs(5015) <= '1';
    layer0_outputs(5016) <= (inputs(50)) xor (inputs(241));
    layer0_outputs(5017) <= (inputs(129)) xor (inputs(187));
    layer0_outputs(5018) <= not((inputs(87)) or (inputs(131)));
    layer0_outputs(5019) <= (inputs(151)) and not (inputs(191));
    layer0_outputs(5020) <= (inputs(160)) xor (inputs(132));
    layer0_outputs(5021) <= (inputs(139)) xor (inputs(188));
    layer0_outputs(5022) <= (inputs(253)) and not (inputs(163));
    layer0_outputs(5023) <= inputs(223);
    layer0_outputs(5024) <= not((inputs(105)) xor (inputs(162)));
    layer0_outputs(5025) <= (inputs(133)) and not (inputs(197));
    layer0_outputs(5026) <= not(inputs(125));
    layer0_outputs(5027) <= not(inputs(243));
    layer0_outputs(5028) <= not((inputs(190)) or (inputs(242)));
    layer0_outputs(5029) <= (inputs(110)) and (inputs(222));
    layer0_outputs(5030) <= not((inputs(131)) or (inputs(122)));
    layer0_outputs(5031) <= not(inputs(196)) or (inputs(128));
    layer0_outputs(5032) <= inputs(198);
    layer0_outputs(5033) <= not((inputs(33)) or (inputs(174)));
    layer0_outputs(5034) <= not(inputs(70)) or (inputs(45));
    layer0_outputs(5035) <= not((inputs(245)) xor (inputs(110)));
    layer0_outputs(5036) <= not(inputs(29)) or (inputs(124));
    layer0_outputs(5037) <= not(inputs(24));
    layer0_outputs(5038) <= not((inputs(26)) xor (inputs(166)));
    layer0_outputs(5039) <= (inputs(49)) and not (inputs(129));
    layer0_outputs(5040) <= not(inputs(115)) or (inputs(192));
    layer0_outputs(5041) <= (inputs(97)) xor (inputs(138));
    layer0_outputs(5042) <= not(inputs(125)) or (inputs(240));
    layer0_outputs(5043) <= inputs(5);
    layer0_outputs(5044) <= '1';
    layer0_outputs(5045) <= not(inputs(100));
    layer0_outputs(5046) <= not((inputs(172)) or (inputs(195)));
    layer0_outputs(5047) <= not((inputs(8)) xor (inputs(44)));
    layer0_outputs(5048) <= '1';
    layer0_outputs(5049) <= inputs(94);
    layer0_outputs(5050) <= not((inputs(52)) xor (inputs(114)));
    layer0_outputs(5051) <= not((inputs(221)) xor (inputs(171)));
    layer0_outputs(5052) <= inputs(172);
    layer0_outputs(5053) <= (inputs(227)) xor (inputs(68));
    layer0_outputs(5054) <= (inputs(9)) xor (inputs(117));
    layer0_outputs(5055) <= not(inputs(170)) or (inputs(221));
    layer0_outputs(5056) <= (inputs(197)) and not (inputs(40));
    layer0_outputs(5057) <= inputs(196);
    layer0_outputs(5058) <= not(inputs(100));
    layer0_outputs(5059) <= '0';
    layer0_outputs(5060) <= not((inputs(254)) or (inputs(92)));
    layer0_outputs(5061) <= (inputs(27)) and not (inputs(203));
    layer0_outputs(5062) <= (inputs(211)) or (inputs(104));
    layer0_outputs(5063) <= (inputs(47)) or (inputs(217));
    layer0_outputs(5064) <= (inputs(74)) xor (inputs(111));
    layer0_outputs(5065) <= (inputs(103)) or (inputs(82));
    layer0_outputs(5066) <= (inputs(66)) and (inputs(80));
    layer0_outputs(5067) <= not(inputs(172));
    layer0_outputs(5068) <= inputs(93);
    layer0_outputs(5069) <= '1';
    layer0_outputs(5070) <= (inputs(159)) and (inputs(27));
    layer0_outputs(5071) <= not((inputs(160)) and (inputs(53)));
    layer0_outputs(5072) <= not(inputs(169));
    layer0_outputs(5073) <= not(inputs(103)) or (inputs(221));
    layer0_outputs(5074) <= not(inputs(40));
    layer0_outputs(5075) <= inputs(42);
    layer0_outputs(5076) <= not(inputs(68)) or (inputs(223));
    layer0_outputs(5077) <= not(inputs(226));
    layer0_outputs(5078) <= (inputs(174)) and not (inputs(235));
    layer0_outputs(5079) <= (inputs(120)) and not (inputs(143));
    layer0_outputs(5080) <= inputs(228);
    layer0_outputs(5081) <= not((inputs(93)) or (inputs(30)));
    layer0_outputs(5082) <= (inputs(138)) and not (inputs(69));
    layer0_outputs(5083) <= (inputs(120)) and not (inputs(26));
    layer0_outputs(5084) <= (inputs(109)) and not (inputs(255));
    layer0_outputs(5085) <= inputs(94);
    layer0_outputs(5086) <= '1';
    layer0_outputs(5087) <= not(inputs(160)) or (inputs(31));
    layer0_outputs(5088) <= inputs(246);
    layer0_outputs(5089) <= (inputs(134)) and not (inputs(104));
    layer0_outputs(5090) <= not(inputs(172));
    layer0_outputs(5091) <= (inputs(32)) or (inputs(10));
    layer0_outputs(5092) <= (inputs(23)) or (inputs(226));
    layer0_outputs(5093) <= inputs(40);
    layer0_outputs(5094) <= (inputs(171)) and not (inputs(229));
    layer0_outputs(5095) <= not(inputs(82)) or (inputs(211));
    layer0_outputs(5096) <= not(inputs(210)) or (inputs(204));
    layer0_outputs(5097) <= (inputs(214)) or (inputs(50));
    layer0_outputs(5098) <= not(inputs(113)) or (inputs(205));
    layer0_outputs(5099) <= '1';
    layer0_outputs(5100) <= not(inputs(42));
    layer0_outputs(5101) <= (inputs(26)) xor (inputs(107));
    layer0_outputs(5102) <= inputs(9);
    layer0_outputs(5103) <= inputs(199);
    layer0_outputs(5104) <= (inputs(24)) xor (inputs(226));
    layer0_outputs(5105) <= not((inputs(227)) or (inputs(236)));
    layer0_outputs(5106) <= (inputs(236)) or (inputs(75));
    layer0_outputs(5107) <= (inputs(166)) and not (inputs(106));
    layer0_outputs(5108) <= (inputs(47)) xor (inputs(164));
    layer0_outputs(5109) <= '0';
    layer0_outputs(5110) <= not((inputs(216)) or (inputs(197)));
    layer0_outputs(5111) <= inputs(140);
    layer0_outputs(5112) <= '1';
    layer0_outputs(5113) <= not(inputs(155)) or (inputs(53));
    layer0_outputs(5114) <= (inputs(83)) and not (inputs(226));
    layer0_outputs(5115) <= (inputs(43)) xor (inputs(31));
    layer0_outputs(5116) <= (inputs(87)) or (inputs(209));
    layer0_outputs(5117) <= not((inputs(92)) xor (inputs(116)));
    layer0_outputs(5118) <= (inputs(180)) and not (inputs(33));
    layer0_outputs(5119) <= not(inputs(203));
    layer0_outputs(5120) <= (inputs(178)) or (inputs(34));
    layer0_outputs(5121) <= not(inputs(169));
    layer0_outputs(5122) <= inputs(29);
    layer0_outputs(5123) <= '0';
    layer0_outputs(5124) <= '1';
    layer0_outputs(5125) <= (inputs(189)) xor (inputs(1));
    layer0_outputs(5126) <= not((inputs(109)) or (inputs(21)));
    layer0_outputs(5127) <= inputs(205);
    layer0_outputs(5128) <= (inputs(72)) or (inputs(234));
    layer0_outputs(5129) <= '0';
    layer0_outputs(5130) <= (inputs(139)) and not (inputs(235));
    layer0_outputs(5131) <= not(inputs(84)) or (inputs(203));
    layer0_outputs(5132) <= not(inputs(218));
    layer0_outputs(5133) <= not(inputs(51)) or (inputs(12));
    layer0_outputs(5134) <= inputs(233);
    layer0_outputs(5135) <= not(inputs(72)) or (inputs(113));
    layer0_outputs(5136) <= (inputs(211)) and not (inputs(200));
    layer0_outputs(5137) <= inputs(91);
    layer0_outputs(5138) <= not(inputs(153));
    layer0_outputs(5139) <= (inputs(48)) xor (inputs(182));
    layer0_outputs(5140) <= (inputs(179)) and not (inputs(224));
    layer0_outputs(5141) <= (inputs(51)) xor (inputs(162));
    layer0_outputs(5142) <= (inputs(6)) or (inputs(183));
    layer0_outputs(5143) <= '0';
    layer0_outputs(5144) <= (inputs(193)) or (inputs(68));
    layer0_outputs(5145) <= not(inputs(105)) or (inputs(222));
    layer0_outputs(5146) <= '1';
    layer0_outputs(5147) <= not(inputs(39));
    layer0_outputs(5148) <= '1';
    layer0_outputs(5149) <= (inputs(69)) or (inputs(201));
    layer0_outputs(5150) <= (inputs(2)) and (inputs(158));
    layer0_outputs(5151) <= not(inputs(90));
    layer0_outputs(5152) <= not(inputs(87)) or (inputs(227));
    layer0_outputs(5153) <= inputs(111);
    layer0_outputs(5154) <= (inputs(164)) or (inputs(125));
    layer0_outputs(5155) <= not(inputs(135));
    layer0_outputs(5156) <= not((inputs(204)) xor (inputs(74)));
    layer0_outputs(5157) <= not((inputs(9)) xor (inputs(202)));
    layer0_outputs(5158) <= not(inputs(68)) or (inputs(26));
    layer0_outputs(5159) <= (inputs(192)) and (inputs(24));
    layer0_outputs(5160) <= not(inputs(199));
    layer0_outputs(5161) <= not(inputs(207));
    layer0_outputs(5162) <= (inputs(52)) and not (inputs(44));
    layer0_outputs(5163) <= (inputs(108)) and (inputs(239));
    layer0_outputs(5164) <= not(inputs(225)) or (inputs(250));
    layer0_outputs(5165) <= '1';
    layer0_outputs(5166) <= (inputs(211)) and not (inputs(177));
    layer0_outputs(5167) <= (inputs(204)) xor (inputs(171));
    layer0_outputs(5168) <= not(inputs(181));
    layer0_outputs(5169) <= (inputs(104)) xor (inputs(225));
    layer0_outputs(5170) <= not(inputs(101));
    layer0_outputs(5171) <= not((inputs(227)) and (inputs(233)));
    layer0_outputs(5172) <= inputs(109);
    layer0_outputs(5173) <= (inputs(219)) or (inputs(128));
    layer0_outputs(5174) <= '0';
    layer0_outputs(5175) <= not((inputs(146)) and (inputs(238)));
    layer0_outputs(5176) <= not((inputs(169)) or (inputs(188)));
    layer0_outputs(5177) <= not((inputs(69)) xor (inputs(188)));
    layer0_outputs(5178) <= not(inputs(164));
    layer0_outputs(5179) <= not(inputs(101));
    layer0_outputs(5180) <= not((inputs(85)) or (inputs(110)));
    layer0_outputs(5181) <= not((inputs(199)) or (inputs(205)));
    layer0_outputs(5182) <= '0';
    layer0_outputs(5183) <= inputs(198);
    layer0_outputs(5184) <= not((inputs(173)) or (inputs(127)));
    layer0_outputs(5185) <= (inputs(155)) and not (inputs(82));
    layer0_outputs(5186) <= not(inputs(213)) or (inputs(224));
    layer0_outputs(5187) <= inputs(41);
    layer0_outputs(5188) <= (inputs(99)) or (inputs(120));
    layer0_outputs(5189) <= not(inputs(36));
    layer0_outputs(5190) <= (inputs(77)) or (inputs(151));
    layer0_outputs(5191) <= '1';
    layer0_outputs(5192) <= not((inputs(61)) xor (inputs(183)));
    layer0_outputs(5193) <= (inputs(169)) and not (inputs(162));
    layer0_outputs(5194) <= not(inputs(8)) or (inputs(95));
    layer0_outputs(5195) <= not((inputs(210)) or (inputs(149)));
    layer0_outputs(5196) <= (inputs(9)) xor (inputs(237));
    layer0_outputs(5197) <= '1';
    layer0_outputs(5198) <= (inputs(194)) or (inputs(179));
    layer0_outputs(5199) <= inputs(24);
    layer0_outputs(5200) <= (inputs(92)) or (inputs(230));
    layer0_outputs(5201) <= not((inputs(115)) or (inputs(85)));
    layer0_outputs(5202) <= (inputs(54)) and not (inputs(115));
    layer0_outputs(5203) <= (inputs(112)) or (inputs(164));
    layer0_outputs(5204) <= (inputs(188)) xor (inputs(154));
    layer0_outputs(5205) <= (inputs(192)) and not (inputs(144));
    layer0_outputs(5206) <= inputs(17);
    layer0_outputs(5207) <= (inputs(233)) and not (inputs(79));
    layer0_outputs(5208) <= inputs(181);
    layer0_outputs(5209) <= (inputs(243)) or (inputs(40));
    layer0_outputs(5210) <= inputs(111);
    layer0_outputs(5211) <= not(inputs(170)) or (inputs(67));
    layer0_outputs(5212) <= not((inputs(18)) xor (inputs(101)));
    layer0_outputs(5213) <= not((inputs(1)) and (inputs(210)));
    layer0_outputs(5214) <= not((inputs(34)) xor (inputs(154)));
    layer0_outputs(5215) <= inputs(38);
    layer0_outputs(5216) <= inputs(91);
    layer0_outputs(5217) <= not((inputs(5)) xor (inputs(205)));
    layer0_outputs(5218) <= not((inputs(0)) xor (inputs(238)));
    layer0_outputs(5219) <= not(inputs(39)) or (inputs(253));
    layer0_outputs(5220) <= (inputs(212)) or (inputs(58));
    layer0_outputs(5221) <= not((inputs(254)) and (inputs(249)));
    layer0_outputs(5222) <= (inputs(90)) xor (inputs(159));
    layer0_outputs(5223) <= not((inputs(242)) xor (inputs(239)));
    layer0_outputs(5224) <= inputs(207);
    layer0_outputs(5225) <= (inputs(98)) or (inputs(91));
    layer0_outputs(5226) <= not((inputs(59)) xor (inputs(75)));
    layer0_outputs(5227) <= not((inputs(240)) or (inputs(224)));
    layer0_outputs(5228) <= (inputs(137)) xor (inputs(109));
    layer0_outputs(5229) <= not(inputs(55)) or (inputs(230));
    layer0_outputs(5230) <= not(inputs(206));
    layer0_outputs(5231) <= not((inputs(69)) xor (inputs(56)));
    layer0_outputs(5232) <= inputs(168);
    layer0_outputs(5233) <= not(inputs(35)) or (inputs(29));
    layer0_outputs(5234) <= not((inputs(87)) or (inputs(87)));
    layer0_outputs(5235) <= (inputs(82)) and (inputs(14));
    layer0_outputs(5236) <= (inputs(65)) or (inputs(190));
    layer0_outputs(5237) <= not(inputs(105));
    layer0_outputs(5238) <= not(inputs(216)) or (inputs(209));
    layer0_outputs(5239) <= not((inputs(215)) or (inputs(145)));
    layer0_outputs(5240) <= inputs(54);
    layer0_outputs(5241) <= (inputs(59)) xor (inputs(77));
    layer0_outputs(5242) <= not(inputs(72));
    layer0_outputs(5243) <= (inputs(42)) and not (inputs(224));
    layer0_outputs(5244) <= (inputs(152)) and not (inputs(187));
    layer0_outputs(5245) <= not(inputs(115)) or (inputs(50));
    layer0_outputs(5246) <= (inputs(171)) and (inputs(159));
    layer0_outputs(5247) <= not(inputs(13)) or (inputs(145));
    layer0_outputs(5248) <= (inputs(156)) or (inputs(127));
    layer0_outputs(5249) <= inputs(163);
    layer0_outputs(5250) <= not(inputs(23));
    layer0_outputs(5251) <= not((inputs(234)) or (inputs(253)));
    layer0_outputs(5252) <= not(inputs(213));
    layer0_outputs(5253) <= not(inputs(61));
    layer0_outputs(5254) <= (inputs(67)) and not (inputs(159));
    layer0_outputs(5255) <= (inputs(195)) or (inputs(179));
    layer0_outputs(5256) <= not((inputs(82)) or (inputs(230)));
    layer0_outputs(5257) <= not(inputs(132)) or (inputs(23));
    layer0_outputs(5258) <= not((inputs(11)) or (inputs(114)));
    layer0_outputs(5259) <= not((inputs(57)) or (inputs(18)));
    layer0_outputs(5260) <= not((inputs(166)) or (inputs(149)));
    layer0_outputs(5261) <= not(inputs(157));
    layer0_outputs(5262) <= not((inputs(165)) or (inputs(67)));
    layer0_outputs(5263) <= not((inputs(183)) or (inputs(159)));
    layer0_outputs(5264) <= inputs(21);
    layer0_outputs(5265) <= not(inputs(89)) or (inputs(26));
    layer0_outputs(5266) <= not(inputs(122)) or (inputs(205));
    layer0_outputs(5267) <= not((inputs(219)) xor (inputs(226)));
    layer0_outputs(5268) <= (inputs(73)) or (inputs(137));
    layer0_outputs(5269) <= not((inputs(241)) or (inputs(100)));
    layer0_outputs(5270) <= not(inputs(166)) or (inputs(228));
    layer0_outputs(5271) <= '0';
    layer0_outputs(5272) <= not((inputs(110)) or (inputs(37)));
    layer0_outputs(5273) <= not((inputs(74)) or (inputs(94)));
    layer0_outputs(5274) <= not(inputs(93));
    layer0_outputs(5275) <= (inputs(100)) xor (inputs(205));
    layer0_outputs(5276) <= (inputs(106)) or (inputs(106));
    layer0_outputs(5277) <= not((inputs(52)) xor (inputs(181)));
    layer0_outputs(5278) <= inputs(86);
    layer0_outputs(5279) <= (inputs(157)) and (inputs(108));
    layer0_outputs(5280) <= (inputs(25)) or (inputs(166));
    layer0_outputs(5281) <= not(inputs(42));
    layer0_outputs(5282) <= not(inputs(72)) or (inputs(180));
    layer0_outputs(5283) <= inputs(160);
    layer0_outputs(5284) <= (inputs(198)) xor (inputs(254));
    layer0_outputs(5285) <= (inputs(98)) and not (inputs(250));
    layer0_outputs(5286) <= (inputs(22)) and (inputs(50));
    layer0_outputs(5287) <= not(inputs(55)) or (inputs(161));
    layer0_outputs(5288) <= inputs(163);
    layer0_outputs(5289) <= (inputs(84)) or (inputs(3));
    layer0_outputs(5290) <= not(inputs(44)) or (inputs(131));
    layer0_outputs(5291) <= not((inputs(171)) or (inputs(64)));
    layer0_outputs(5292) <= (inputs(205)) xor (inputs(93));
    layer0_outputs(5293) <= not((inputs(131)) xor (inputs(41)));
    layer0_outputs(5294) <= (inputs(186)) xor (inputs(25));
    layer0_outputs(5295) <= (inputs(68)) or (inputs(62));
    layer0_outputs(5296) <= not(inputs(220)) or (inputs(199));
    layer0_outputs(5297) <= (inputs(164)) and not (inputs(113));
    layer0_outputs(5298) <= (inputs(28)) and not (inputs(246));
    layer0_outputs(5299) <= (inputs(121)) or (inputs(158));
    layer0_outputs(5300) <= (inputs(168)) xor (inputs(10));
    layer0_outputs(5301) <= not((inputs(239)) or (inputs(176)));
    layer0_outputs(5302) <= (inputs(189)) or (inputs(43));
    layer0_outputs(5303) <= not((inputs(104)) xor (inputs(247)));
    layer0_outputs(5304) <= not((inputs(189)) or (inputs(56)));
    layer0_outputs(5305) <= (inputs(112)) xor (inputs(156));
    layer0_outputs(5306) <= inputs(212);
    layer0_outputs(5307) <= (inputs(213)) or (inputs(215));
    layer0_outputs(5308) <= (inputs(255)) xor (inputs(220));
    layer0_outputs(5309) <= not((inputs(2)) and (inputs(192)));
    layer0_outputs(5310) <= not((inputs(22)) xor (inputs(171)));
    layer0_outputs(5311) <= not(inputs(86)) or (inputs(81));
    layer0_outputs(5312) <= (inputs(49)) and (inputs(241));
    layer0_outputs(5313) <= not(inputs(122)) or (inputs(4));
    layer0_outputs(5314) <= inputs(132);
    layer0_outputs(5315) <= not((inputs(146)) xor (inputs(209)));
    layer0_outputs(5316) <= (inputs(213)) or (inputs(46));
    layer0_outputs(5317) <= not((inputs(5)) or (inputs(213)));
    layer0_outputs(5318) <= (inputs(53)) xor (inputs(121));
    layer0_outputs(5319) <= not(inputs(90)) or (inputs(173));
    layer0_outputs(5320) <= (inputs(224)) and (inputs(23));
    layer0_outputs(5321) <= inputs(151);
    layer0_outputs(5322) <= not(inputs(91)) or (inputs(197));
    layer0_outputs(5323) <= not((inputs(74)) xor (inputs(105)));
    layer0_outputs(5324) <= (inputs(35)) and not (inputs(205));
    layer0_outputs(5325) <= inputs(236);
    layer0_outputs(5326) <= inputs(194);
    layer0_outputs(5327) <= inputs(244);
    layer0_outputs(5328) <= (inputs(91)) xor (inputs(168));
    layer0_outputs(5329) <= not(inputs(214)) or (inputs(37));
    layer0_outputs(5330) <= inputs(109);
    layer0_outputs(5331) <= inputs(174);
    layer0_outputs(5332) <= inputs(70);
    layer0_outputs(5333) <= (inputs(232)) or (inputs(243));
    layer0_outputs(5334) <= not((inputs(201)) and (inputs(188)));
    layer0_outputs(5335) <= inputs(52);
    layer0_outputs(5336) <= inputs(70);
    layer0_outputs(5337) <= (inputs(108)) and not (inputs(26));
    layer0_outputs(5338) <= inputs(162);
    layer0_outputs(5339) <= (inputs(191)) and not (inputs(83));
    layer0_outputs(5340) <= '0';
    layer0_outputs(5341) <= (inputs(203)) and (inputs(42));
    layer0_outputs(5342) <= not((inputs(190)) xor (inputs(90)));
    layer0_outputs(5343) <= not(inputs(235)) or (inputs(252));
    layer0_outputs(5344) <= inputs(202);
    layer0_outputs(5345) <= (inputs(252)) and not (inputs(225));
    layer0_outputs(5346) <= inputs(80);
    layer0_outputs(5347) <= (inputs(61)) and not (inputs(158));
    layer0_outputs(5348) <= (inputs(84)) xor (inputs(115));
    layer0_outputs(5349) <= not(inputs(231)) or (inputs(61));
    layer0_outputs(5350) <= not((inputs(211)) xor (inputs(38)));
    layer0_outputs(5351) <= not((inputs(101)) xor (inputs(72)));
    layer0_outputs(5352) <= not(inputs(103));
    layer0_outputs(5353) <= not(inputs(231)) or (inputs(162));
    layer0_outputs(5354) <= (inputs(78)) xor (inputs(98));
    layer0_outputs(5355) <= not((inputs(194)) or (inputs(42)));
    layer0_outputs(5356) <= not((inputs(182)) or (inputs(240)));
    layer0_outputs(5357) <= (inputs(93)) or (inputs(64));
    layer0_outputs(5358) <= not((inputs(3)) or (inputs(163)));
    layer0_outputs(5359) <= not((inputs(6)) and (inputs(217)));
    layer0_outputs(5360) <= inputs(215);
    layer0_outputs(5361) <= not(inputs(106));
    layer0_outputs(5362) <= (inputs(16)) or (inputs(82));
    layer0_outputs(5363) <= (inputs(102)) and not (inputs(247));
    layer0_outputs(5364) <= (inputs(153)) xor (inputs(228));
    layer0_outputs(5365) <= (inputs(141)) and not (inputs(129));
    layer0_outputs(5366) <= inputs(12);
    layer0_outputs(5367) <= not(inputs(36));
    layer0_outputs(5368) <= not((inputs(20)) xor (inputs(200)));
    layer0_outputs(5369) <= (inputs(214)) and not (inputs(87));
    layer0_outputs(5370) <= inputs(103);
    layer0_outputs(5371) <= (inputs(213)) or (inputs(185));
    layer0_outputs(5372) <= not(inputs(74));
    layer0_outputs(5373) <= (inputs(213)) and not (inputs(26));
    layer0_outputs(5374) <= not(inputs(58)) or (inputs(130));
    layer0_outputs(5375) <= '0';
    layer0_outputs(5376) <= (inputs(237)) or (inputs(214));
    layer0_outputs(5377) <= not((inputs(122)) or (inputs(129)));
    layer0_outputs(5378) <= (inputs(73)) and not (inputs(213));
    layer0_outputs(5379) <= not(inputs(240));
    layer0_outputs(5380) <= not(inputs(40));
    layer0_outputs(5381) <= inputs(141);
    layer0_outputs(5382) <= inputs(250);
    layer0_outputs(5383) <= not((inputs(34)) or (inputs(226)));
    layer0_outputs(5384) <= not((inputs(239)) or (inputs(71)));
    layer0_outputs(5385) <= (inputs(142)) xor (inputs(129));
    layer0_outputs(5386) <= not(inputs(129));
    layer0_outputs(5387) <= (inputs(245)) xor (inputs(226));
    layer0_outputs(5388) <= not((inputs(155)) or (inputs(194)));
    layer0_outputs(5389) <= not((inputs(15)) xor (inputs(230)));
    layer0_outputs(5390) <= inputs(77);
    layer0_outputs(5391) <= not(inputs(208));
    layer0_outputs(5392) <= not(inputs(209));
    layer0_outputs(5393) <= not((inputs(48)) and (inputs(156)));
    layer0_outputs(5394) <= not((inputs(5)) or (inputs(25)));
    layer0_outputs(5395) <= not((inputs(231)) or (inputs(187)));
    layer0_outputs(5396) <= not(inputs(205));
    layer0_outputs(5397) <= not((inputs(173)) or (inputs(172)));
    layer0_outputs(5398) <= inputs(5);
    layer0_outputs(5399) <= (inputs(176)) or (inputs(10));
    layer0_outputs(5400) <= not((inputs(17)) xor (inputs(197)));
    layer0_outputs(5401) <= (inputs(36)) and (inputs(192));
    layer0_outputs(5402) <= not((inputs(2)) xor (inputs(134)));
    layer0_outputs(5403) <= not((inputs(79)) xor (inputs(40)));
    layer0_outputs(5404) <= '0';
    layer0_outputs(5405) <= not(inputs(138)) or (inputs(126));
    layer0_outputs(5406) <= not(inputs(127)) or (inputs(14));
    layer0_outputs(5407) <= not((inputs(136)) xor (inputs(143)));
    layer0_outputs(5408) <= (inputs(54)) or (inputs(122));
    layer0_outputs(5409) <= not((inputs(211)) or (inputs(131)));
    layer0_outputs(5410) <= (inputs(87)) xor (inputs(63));
    layer0_outputs(5411) <= (inputs(184)) and (inputs(86));
    layer0_outputs(5412) <= not((inputs(71)) or (inputs(99)));
    layer0_outputs(5413) <= not(inputs(195));
    layer0_outputs(5414) <= not(inputs(124));
    layer0_outputs(5415) <= not((inputs(12)) or (inputs(124)));
    layer0_outputs(5416) <= (inputs(75)) or (inputs(17));
    layer0_outputs(5417) <= not((inputs(179)) or (inputs(217)));
    layer0_outputs(5418) <= inputs(89);
    layer0_outputs(5419) <= not((inputs(125)) or (inputs(207)));
    layer0_outputs(5420) <= (inputs(217)) or (inputs(95));
    layer0_outputs(5421) <= (inputs(50)) or (inputs(77));
    layer0_outputs(5422) <= not((inputs(254)) and (inputs(202)));
    layer0_outputs(5423) <= (inputs(166)) xor (inputs(241));
    layer0_outputs(5424) <= (inputs(196)) and not (inputs(51));
    layer0_outputs(5425) <= not(inputs(230)) or (inputs(173));
    layer0_outputs(5426) <= inputs(117);
    layer0_outputs(5427) <= not(inputs(90));
    layer0_outputs(5428) <= (inputs(95)) or (inputs(124));
    layer0_outputs(5429) <= not(inputs(40));
    layer0_outputs(5430) <= not((inputs(214)) or (inputs(91)));
    layer0_outputs(5431) <= (inputs(203)) and (inputs(185));
    layer0_outputs(5432) <= not((inputs(205)) xor (inputs(63)));
    layer0_outputs(5433) <= (inputs(55)) or (inputs(17));
    layer0_outputs(5434) <= inputs(94);
    layer0_outputs(5435) <= not(inputs(132));
    layer0_outputs(5436) <= '1';
    layer0_outputs(5437) <= not((inputs(104)) or (inputs(121)));
    layer0_outputs(5438) <= (inputs(221)) and not (inputs(128));
    layer0_outputs(5439) <= (inputs(230)) and not (inputs(161));
    layer0_outputs(5440) <= not(inputs(123)) or (inputs(145));
    layer0_outputs(5441) <= not((inputs(157)) xor (inputs(18)));
    layer0_outputs(5442) <= (inputs(133)) and not (inputs(162));
    layer0_outputs(5443) <= (inputs(199)) and (inputs(217));
    layer0_outputs(5444) <= not(inputs(20)) or (inputs(95));
    layer0_outputs(5445) <= not((inputs(241)) and (inputs(136)));
    layer0_outputs(5446) <= inputs(76);
    layer0_outputs(5447) <= (inputs(199)) and not (inputs(98));
    layer0_outputs(5448) <= not(inputs(96));
    layer0_outputs(5449) <= not((inputs(204)) xor (inputs(108)));
    layer0_outputs(5450) <= not(inputs(9));
    layer0_outputs(5451) <= (inputs(52)) xor (inputs(157));
    layer0_outputs(5452) <= not(inputs(145));
    layer0_outputs(5453) <= not(inputs(151));
    layer0_outputs(5454) <= (inputs(199)) and not (inputs(47));
    layer0_outputs(5455) <= (inputs(88)) and not (inputs(62));
    layer0_outputs(5456) <= not((inputs(59)) xor (inputs(177)));
    layer0_outputs(5457) <= not(inputs(143)) or (inputs(128));
    layer0_outputs(5458) <= (inputs(165)) or (inputs(224));
    layer0_outputs(5459) <= (inputs(55)) and not (inputs(141));
    layer0_outputs(5460) <= not((inputs(66)) xor (inputs(75)));
    layer0_outputs(5461) <= not((inputs(245)) xor (inputs(197)));
    layer0_outputs(5462) <= not(inputs(170));
    layer0_outputs(5463) <= '0';
    layer0_outputs(5464) <= not((inputs(37)) or (inputs(95)));
    layer0_outputs(5465) <= not(inputs(72));
    layer0_outputs(5466) <= not(inputs(169)) or (inputs(253));
    layer0_outputs(5467) <= '1';
    layer0_outputs(5468) <= inputs(216);
    layer0_outputs(5469) <= '0';
    layer0_outputs(5470) <= inputs(43);
    layer0_outputs(5471) <= inputs(195);
    layer0_outputs(5472) <= not((inputs(233)) or (inputs(137)));
    layer0_outputs(5473) <= inputs(132);
    layer0_outputs(5474) <= inputs(139);
    layer0_outputs(5475) <= (inputs(170)) and not (inputs(3));
    layer0_outputs(5476) <= not((inputs(110)) or (inputs(149)));
    layer0_outputs(5477) <= (inputs(222)) and (inputs(252));
    layer0_outputs(5478) <= not(inputs(103)) or (inputs(232));
    layer0_outputs(5479) <= not(inputs(192)) or (inputs(24));
    layer0_outputs(5480) <= not((inputs(133)) or (inputs(180)));
    layer0_outputs(5481) <= (inputs(20)) xor (inputs(119));
    layer0_outputs(5482) <= not(inputs(132));
    layer0_outputs(5483) <= not((inputs(27)) xor (inputs(229)));
    layer0_outputs(5484) <= not(inputs(202)) or (inputs(236));
    layer0_outputs(5485) <= not(inputs(65));
    layer0_outputs(5486) <= (inputs(184)) and not (inputs(135));
    layer0_outputs(5487) <= (inputs(74)) xor (inputs(246));
    layer0_outputs(5488) <= inputs(49);
    layer0_outputs(5489) <= (inputs(213)) or (inputs(241));
    layer0_outputs(5490) <= not(inputs(215)) or (inputs(202));
    layer0_outputs(5491) <= not(inputs(20));
    layer0_outputs(5492) <= (inputs(178)) or (inputs(134));
    layer0_outputs(5493) <= (inputs(185)) or (inputs(201));
    layer0_outputs(5494) <= not(inputs(161)) or (inputs(58));
    layer0_outputs(5495) <= not(inputs(133)) or (inputs(235));
    layer0_outputs(5496) <= not(inputs(30));
    layer0_outputs(5497) <= not(inputs(75));
    layer0_outputs(5498) <= (inputs(88)) xor (inputs(252));
    layer0_outputs(5499) <= not(inputs(50)) or (inputs(186));
    layer0_outputs(5500) <= not(inputs(213));
    layer0_outputs(5501) <= (inputs(190)) xor (inputs(152));
    layer0_outputs(5502) <= not((inputs(40)) or (inputs(4)));
    layer0_outputs(5503) <= (inputs(106)) xor (inputs(98));
    layer0_outputs(5504) <= not((inputs(21)) xor (inputs(134)));
    layer0_outputs(5505) <= (inputs(126)) or (inputs(74));
    layer0_outputs(5506) <= not((inputs(81)) or (inputs(134)));
    layer0_outputs(5507) <= inputs(90);
    layer0_outputs(5508) <= (inputs(39)) xor (inputs(105));
    layer0_outputs(5509) <= not((inputs(69)) or (inputs(212)));
    layer0_outputs(5510) <= not((inputs(22)) xor (inputs(214)));
    layer0_outputs(5511) <= not(inputs(148)) or (inputs(227));
    layer0_outputs(5512) <= not((inputs(117)) xor (inputs(31)));
    layer0_outputs(5513) <= not((inputs(208)) xor (inputs(66)));
    layer0_outputs(5514) <= not(inputs(180));
    layer0_outputs(5515) <= not((inputs(88)) xor (inputs(224)));
    layer0_outputs(5516) <= not((inputs(71)) and (inputs(221)));
    layer0_outputs(5517) <= (inputs(196)) and not (inputs(149));
    layer0_outputs(5518) <= not(inputs(136)) or (inputs(212));
    layer0_outputs(5519) <= not(inputs(48));
    layer0_outputs(5520) <= not((inputs(199)) and (inputs(132)));
    layer0_outputs(5521) <= not(inputs(213)) or (inputs(229));
    layer0_outputs(5522) <= not(inputs(188));
    layer0_outputs(5523) <= inputs(121);
    layer0_outputs(5524) <= not((inputs(110)) or (inputs(109)));
    layer0_outputs(5525) <= (inputs(96)) xor (inputs(146));
    layer0_outputs(5526) <= inputs(55);
    layer0_outputs(5527) <= not(inputs(141)) or (inputs(138));
    layer0_outputs(5528) <= not(inputs(122));
    layer0_outputs(5529) <= (inputs(91)) or (inputs(170));
    layer0_outputs(5530) <= '1';
    layer0_outputs(5531) <= '0';
    layer0_outputs(5532) <= inputs(55);
    layer0_outputs(5533) <= inputs(179);
    layer0_outputs(5534) <= inputs(86);
    layer0_outputs(5535) <= (inputs(123)) and not (inputs(42));
    layer0_outputs(5536) <= not((inputs(153)) xor (inputs(175)));
    layer0_outputs(5537) <= (inputs(66)) or (inputs(247));
    layer0_outputs(5538) <= inputs(57);
    layer0_outputs(5539) <= '1';
    layer0_outputs(5540) <= not(inputs(149));
    layer0_outputs(5541) <= not(inputs(232));
    layer0_outputs(5542) <= not(inputs(99)) or (inputs(202));
    layer0_outputs(5543) <= not((inputs(232)) or (inputs(233)));
    layer0_outputs(5544) <= not((inputs(4)) or (inputs(12)));
    layer0_outputs(5545) <= not((inputs(66)) or (inputs(211)));
    layer0_outputs(5546) <= '0';
    layer0_outputs(5547) <= (inputs(141)) or (inputs(26));
    layer0_outputs(5548) <= not(inputs(195));
    layer0_outputs(5549) <= inputs(131);
    layer0_outputs(5550) <= not(inputs(83)) or (inputs(164));
    layer0_outputs(5551) <= not(inputs(172));
    layer0_outputs(5552) <= (inputs(255)) and not (inputs(83));
    layer0_outputs(5553) <= not((inputs(189)) or (inputs(47)));
    layer0_outputs(5554) <= inputs(140);
    layer0_outputs(5555) <= (inputs(245)) and not (inputs(34));
    layer0_outputs(5556) <= inputs(203);
    layer0_outputs(5557) <= not((inputs(153)) or (inputs(30)));
    layer0_outputs(5558) <= (inputs(38)) or (inputs(72));
    layer0_outputs(5559) <= inputs(54);
    layer0_outputs(5560) <= '1';
    layer0_outputs(5561) <= (inputs(154)) and not (inputs(108));
    layer0_outputs(5562) <= not((inputs(39)) or (inputs(65)));
    layer0_outputs(5563) <= (inputs(59)) and not (inputs(111));
    layer0_outputs(5564) <= not((inputs(148)) and (inputs(213)));
    layer0_outputs(5565) <= (inputs(41)) xor (inputs(48));
    layer0_outputs(5566) <= not(inputs(177));
    layer0_outputs(5567) <= (inputs(85)) or (inputs(22));
    layer0_outputs(5568) <= not((inputs(144)) or (inputs(148)));
    layer0_outputs(5569) <= '0';
    layer0_outputs(5570) <= (inputs(206)) or (inputs(165));
    layer0_outputs(5571) <= (inputs(183)) xor (inputs(181));
    layer0_outputs(5572) <= not(inputs(183));
    layer0_outputs(5573) <= not(inputs(88));
    layer0_outputs(5574) <= not((inputs(192)) or (inputs(201)));
    layer0_outputs(5575) <= (inputs(18)) and not (inputs(70));
    layer0_outputs(5576) <= not(inputs(5)) or (inputs(111));
    layer0_outputs(5577) <= (inputs(52)) and not (inputs(211));
    layer0_outputs(5578) <= (inputs(158)) or (inputs(190));
    layer0_outputs(5579) <= not(inputs(165));
    layer0_outputs(5580) <= not((inputs(130)) xor (inputs(121)));
    layer0_outputs(5581) <= not(inputs(92));
    layer0_outputs(5582) <= not(inputs(208));
    layer0_outputs(5583) <= (inputs(147)) and not (inputs(13));
    layer0_outputs(5584) <= (inputs(236)) and not (inputs(162));
    layer0_outputs(5585) <= not((inputs(49)) xor (inputs(189)));
    layer0_outputs(5586) <= not((inputs(171)) or (inputs(210)));
    layer0_outputs(5587) <= not(inputs(101)) or (inputs(151));
    layer0_outputs(5588) <= inputs(138);
    layer0_outputs(5589) <= not(inputs(47));
    layer0_outputs(5590) <= (inputs(250)) or (inputs(20));
    layer0_outputs(5591) <= '0';
    layer0_outputs(5592) <= (inputs(205)) or (inputs(56));
    layer0_outputs(5593) <= inputs(199);
    layer0_outputs(5594) <= (inputs(97)) xor (inputs(235));
    layer0_outputs(5595) <= (inputs(129)) and not (inputs(253));
    layer0_outputs(5596) <= '0';
    layer0_outputs(5597) <= (inputs(181)) or (inputs(166));
    layer0_outputs(5598) <= (inputs(238)) or (inputs(199));
    layer0_outputs(5599) <= not(inputs(68)) or (inputs(2));
    layer0_outputs(5600) <= (inputs(182)) or (inputs(180));
    layer0_outputs(5601) <= (inputs(218)) and not (inputs(126));
    layer0_outputs(5602) <= (inputs(17)) xor (inputs(183));
    layer0_outputs(5603) <= (inputs(55)) or (inputs(180));
    layer0_outputs(5604) <= not((inputs(32)) or (inputs(130)));
    layer0_outputs(5605) <= inputs(111);
    layer0_outputs(5606) <= (inputs(213)) or (inputs(223));
    layer0_outputs(5607) <= inputs(119);
    layer0_outputs(5608) <= inputs(211);
    layer0_outputs(5609) <= not((inputs(73)) or (inputs(181)));
    layer0_outputs(5610) <= (inputs(141)) xor (inputs(33));
    layer0_outputs(5611) <= '1';
    layer0_outputs(5612) <= not((inputs(1)) or (inputs(193)));
    layer0_outputs(5613) <= (inputs(69)) and not (inputs(177));
    layer0_outputs(5614) <= (inputs(155)) or (inputs(164));
    layer0_outputs(5615) <= not(inputs(252));
    layer0_outputs(5616) <= (inputs(147)) or (inputs(167));
    layer0_outputs(5617) <= not((inputs(198)) xor (inputs(72)));
    layer0_outputs(5618) <= not(inputs(153));
    layer0_outputs(5619) <= not(inputs(69)) or (inputs(144));
    layer0_outputs(5620) <= not(inputs(77));
    layer0_outputs(5621) <= not(inputs(138)) or (inputs(151));
    layer0_outputs(5622) <= (inputs(109)) and (inputs(235));
    layer0_outputs(5623) <= inputs(39);
    layer0_outputs(5624) <= not(inputs(187)) or (inputs(33));
    layer0_outputs(5625) <= not(inputs(28)) or (inputs(176));
    layer0_outputs(5626) <= not(inputs(15));
    layer0_outputs(5627) <= inputs(103);
    layer0_outputs(5628) <= not(inputs(221)) or (inputs(173));
    layer0_outputs(5629) <= not(inputs(226));
    layer0_outputs(5630) <= (inputs(7)) xor (inputs(139));
    layer0_outputs(5631) <= (inputs(125)) xor (inputs(69));
    layer0_outputs(5632) <= not(inputs(231));
    layer0_outputs(5633) <= (inputs(25)) xor (inputs(68));
    layer0_outputs(5634) <= inputs(61);
    layer0_outputs(5635) <= (inputs(179)) and not (inputs(96));
    layer0_outputs(5636) <= not((inputs(198)) xor (inputs(60)));
    layer0_outputs(5637) <= inputs(163);
    layer0_outputs(5638) <= inputs(100);
    layer0_outputs(5639) <= (inputs(2)) or (inputs(115));
    layer0_outputs(5640) <= (inputs(209)) and not (inputs(226));
    layer0_outputs(5641) <= (inputs(226)) and not (inputs(33));
    layer0_outputs(5642) <= not(inputs(201)) or (inputs(221));
    layer0_outputs(5643) <= (inputs(188)) and not (inputs(137));
    layer0_outputs(5644) <= not((inputs(200)) and (inputs(14)));
    layer0_outputs(5645) <= not(inputs(55)) or (inputs(8));
    layer0_outputs(5646) <= inputs(203);
    layer0_outputs(5647) <= not((inputs(36)) xor (inputs(11)));
    layer0_outputs(5648) <= '1';
    layer0_outputs(5649) <= '1';
    layer0_outputs(5650) <= not(inputs(248)) or (inputs(34));
    layer0_outputs(5651) <= '1';
    layer0_outputs(5652) <= not(inputs(33));
    layer0_outputs(5653) <= inputs(137);
    layer0_outputs(5654) <= not((inputs(153)) or (inputs(178)));
    layer0_outputs(5655) <= (inputs(46)) and not (inputs(11));
    layer0_outputs(5656) <= (inputs(136)) or (inputs(239));
    layer0_outputs(5657) <= not(inputs(64));
    layer0_outputs(5658) <= (inputs(101)) or (inputs(208));
    layer0_outputs(5659) <= (inputs(50)) xor (inputs(103));
    layer0_outputs(5660) <= (inputs(181)) or (inputs(191));
    layer0_outputs(5661) <= inputs(27);
    layer0_outputs(5662) <= not((inputs(215)) xor (inputs(49)));
    layer0_outputs(5663) <= (inputs(158)) and (inputs(21));
    layer0_outputs(5664) <= not(inputs(175));
    layer0_outputs(5665) <= not((inputs(211)) xor (inputs(17)));
    layer0_outputs(5666) <= inputs(133);
    layer0_outputs(5667) <= not(inputs(32)) or (inputs(49));
    layer0_outputs(5668) <= '1';
    layer0_outputs(5669) <= '1';
    layer0_outputs(5670) <= not(inputs(106)) or (inputs(171));
    layer0_outputs(5671) <= (inputs(111)) or (inputs(150));
    layer0_outputs(5672) <= not((inputs(185)) or (inputs(159)));
    layer0_outputs(5673) <= inputs(73);
    layer0_outputs(5674) <= not((inputs(248)) or (inputs(103)));
    layer0_outputs(5675) <= inputs(15);
    layer0_outputs(5676) <= not(inputs(230));
    layer0_outputs(5677) <= (inputs(219)) or (inputs(219));
    layer0_outputs(5678) <= (inputs(180)) and not (inputs(109));
    layer0_outputs(5679) <= inputs(43);
    layer0_outputs(5680) <= not(inputs(168)) or (inputs(189));
    layer0_outputs(5681) <= not(inputs(37));
    layer0_outputs(5682) <= not((inputs(193)) or (inputs(187)));
    layer0_outputs(5683) <= (inputs(200)) or (inputs(36));
    layer0_outputs(5684) <= not(inputs(225)) or (inputs(46));
    layer0_outputs(5685) <= not((inputs(208)) xor (inputs(141)));
    layer0_outputs(5686) <= not((inputs(61)) xor (inputs(12)));
    layer0_outputs(5687) <= (inputs(170)) and not (inputs(2));
    layer0_outputs(5688) <= (inputs(23)) or (inputs(115));
    layer0_outputs(5689) <= (inputs(198)) or (inputs(110));
    layer0_outputs(5690) <= (inputs(85)) and not (inputs(35));
    layer0_outputs(5691) <= (inputs(25)) or (inputs(35));
    layer0_outputs(5692) <= (inputs(117)) and not (inputs(222));
    layer0_outputs(5693) <= (inputs(110)) xor (inputs(35));
    layer0_outputs(5694) <= (inputs(209)) or (inputs(17));
    layer0_outputs(5695) <= (inputs(248)) or (inputs(95));
    layer0_outputs(5696) <= not((inputs(227)) or (inputs(206)));
    layer0_outputs(5697) <= not(inputs(192));
    layer0_outputs(5698) <= (inputs(177)) and not (inputs(75));
    layer0_outputs(5699) <= inputs(54);
    layer0_outputs(5700) <= not(inputs(175)) or (inputs(45));
    layer0_outputs(5701) <= (inputs(97)) and (inputs(246));
    layer0_outputs(5702) <= (inputs(127)) and (inputs(217));
    layer0_outputs(5703) <= not((inputs(87)) or (inputs(150)));
    layer0_outputs(5704) <= (inputs(65)) or (inputs(154));
    layer0_outputs(5705) <= not((inputs(75)) or (inputs(230)));
    layer0_outputs(5706) <= not(inputs(90)) or (inputs(92));
    layer0_outputs(5707) <= not(inputs(187)) or (inputs(7));
    layer0_outputs(5708) <= inputs(71);
    layer0_outputs(5709) <= (inputs(219)) or (inputs(133));
    layer0_outputs(5710) <= (inputs(40)) or (inputs(146));
    layer0_outputs(5711) <= (inputs(234)) or (inputs(223));
    layer0_outputs(5712) <= not(inputs(228));
    layer0_outputs(5713) <= (inputs(183)) and not (inputs(175));
    layer0_outputs(5714) <= not((inputs(138)) xor (inputs(154)));
    layer0_outputs(5715) <= (inputs(155)) and not (inputs(131));
    layer0_outputs(5716) <= not((inputs(38)) or (inputs(83)));
    layer0_outputs(5717) <= (inputs(102)) xor (inputs(81));
    layer0_outputs(5718) <= inputs(132);
    layer0_outputs(5719) <= not(inputs(206));
    layer0_outputs(5720) <= (inputs(67)) xor (inputs(15));
    layer0_outputs(5721) <= not(inputs(99)) or (inputs(142));
    layer0_outputs(5722) <= not((inputs(148)) or (inputs(16)));
    layer0_outputs(5723) <= not(inputs(67)) or (inputs(223));
    layer0_outputs(5724) <= inputs(224);
    layer0_outputs(5725) <= inputs(55);
    layer0_outputs(5726) <= not(inputs(84)) or (inputs(30));
    layer0_outputs(5727) <= (inputs(13)) and not (inputs(204));
    layer0_outputs(5728) <= (inputs(190)) or (inputs(120));
    layer0_outputs(5729) <= inputs(182);
    layer0_outputs(5730) <= not(inputs(235));
    layer0_outputs(5731) <= (inputs(85)) or (inputs(184));
    layer0_outputs(5732) <= not((inputs(116)) or (inputs(75)));
    layer0_outputs(5733) <= (inputs(31)) xor (inputs(7));
    layer0_outputs(5734) <= (inputs(196)) or (inputs(209));
    layer0_outputs(5735) <= not(inputs(24)) or (inputs(109));
    layer0_outputs(5736) <= not((inputs(168)) or (inputs(98)));
    layer0_outputs(5737) <= (inputs(150)) and not (inputs(210));
    layer0_outputs(5738) <= (inputs(154)) or (inputs(241));
    layer0_outputs(5739) <= not(inputs(109));
    layer0_outputs(5740) <= inputs(82);
    layer0_outputs(5741) <= '1';
    layer0_outputs(5742) <= not((inputs(131)) and (inputs(226)));
    layer0_outputs(5743) <= (inputs(63)) xor (inputs(21));
    layer0_outputs(5744) <= not((inputs(146)) or (inputs(40)));
    layer0_outputs(5745) <= not(inputs(200));
    layer0_outputs(5746) <= not((inputs(114)) or (inputs(236)));
    layer0_outputs(5747) <= (inputs(38)) or (inputs(104));
    layer0_outputs(5748) <= not(inputs(218));
    layer0_outputs(5749) <= (inputs(78)) and (inputs(189));
    layer0_outputs(5750) <= not((inputs(248)) or (inputs(247)));
    layer0_outputs(5751) <= (inputs(93)) or (inputs(116));
    layer0_outputs(5752) <= not((inputs(151)) or (inputs(203)));
    layer0_outputs(5753) <= not((inputs(238)) and (inputs(76)));
    layer0_outputs(5754) <= not((inputs(108)) xor (inputs(76)));
    layer0_outputs(5755) <= inputs(61);
    layer0_outputs(5756) <= not(inputs(151));
    layer0_outputs(5757) <= (inputs(137)) and not (inputs(126));
    layer0_outputs(5758) <= not((inputs(153)) or (inputs(34)));
    layer0_outputs(5759) <= (inputs(229)) or (inputs(107));
    layer0_outputs(5760) <= (inputs(149)) or (inputs(166));
    layer0_outputs(5761) <= not(inputs(102)) or (inputs(48));
    layer0_outputs(5762) <= (inputs(36)) and not (inputs(145));
    layer0_outputs(5763) <= inputs(28);
    layer0_outputs(5764) <= (inputs(206)) or (inputs(89));
    layer0_outputs(5765) <= (inputs(209)) xor (inputs(236));
    layer0_outputs(5766) <= not((inputs(49)) or (inputs(137)));
    layer0_outputs(5767) <= (inputs(160)) or (inputs(232));
    layer0_outputs(5768) <= not(inputs(137)) or (inputs(157));
    layer0_outputs(5769) <= '1';
    layer0_outputs(5770) <= (inputs(234)) and not (inputs(208));
    layer0_outputs(5771) <= '1';
    layer0_outputs(5772) <= inputs(144);
    layer0_outputs(5773) <= not(inputs(202));
    layer0_outputs(5774) <= (inputs(41)) or (inputs(200));
    layer0_outputs(5775) <= not((inputs(46)) xor (inputs(227)));
    layer0_outputs(5776) <= inputs(197);
    layer0_outputs(5777) <= not((inputs(164)) or (inputs(95)));
    layer0_outputs(5778) <= (inputs(9)) and not (inputs(193));
    layer0_outputs(5779) <= inputs(165);
    layer0_outputs(5780) <= not(inputs(30));
    layer0_outputs(5781) <= not(inputs(48));
    layer0_outputs(5782) <= '0';
    layer0_outputs(5783) <= not((inputs(53)) and (inputs(197)));
    layer0_outputs(5784) <= not(inputs(97));
    layer0_outputs(5785) <= not(inputs(114)) or (inputs(43));
    layer0_outputs(5786) <= inputs(176);
    layer0_outputs(5787) <= (inputs(126)) xor (inputs(40));
    layer0_outputs(5788) <= inputs(108);
    layer0_outputs(5789) <= (inputs(204)) xor (inputs(167));
    layer0_outputs(5790) <= (inputs(238)) xor (inputs(55));
    layer0_outputs(5791) <= inputs(249);
    layer0_outputs(5792) <= inputs(162);
    layer0_outputs(5793) <= (inputs(70)) or (inputs(234));
    layer0_outputs(5794) <= not((inputs(73)) xor (inputs(221)));
    layer0_outputs(5795) <= (inputs(124)) xor (inputs(4));
    layer0_outputs(5796) <= (inputs(239)) and not (inputs(47));
    layer0_outputs(5797) <= (inputs(201)) and not (inputs(70));
    layer0_outputs(5798) <= (inputs(62)) xor (inputs(19));
    layer0_outputs(5799) <= not(inputs(36)) or (inputs(136));
    layer0_outputs(5800) <= (inputs(143)) and not (inputs(247));
    layer0_outputs(5801) <= inputs(228);
    layer0_outputs(5802) <= inputs(83);
    layer0_outputs(5803) <= not((inputs(227)) xor (inputs(186)));
    layer0_outputs(5804) <= (inputs(51)) and not (inputs(234));
    layer0_outputs(5805) <= (inputs(49)) and (inputs(4));
    layer0_outputs(5806) <= (inputs(124)) or (inputs(24));
    layer0_outputs(5807) <= not((inputs(131)) or (inputs(58)));
    layer0_outputs(5808) <= not(inputs(158)) or (inputs(191));
    layer0_outputs(5809) <= '0';
    layer0_outputs(5810) <= (inputs(234)) and not (inputs(127));
    layer0_outputs(5811) <= not((inputs(181)) xor (inputs(204)));
    layer0_outputs(5812) <= not((inputs(72)) xor (inputs(213)));
    layer0_outputs(5813) <= (inputs(228)) xor (inputs(139));
    layer0_outputs(5814) <= not(inputs(59)) or (inputs(159));
    layer0_outputs(5815) <= not(inputs(142)) or (inputs(66));
    layer0_outputs(5816) <= inputs(187);
    layer0_outputs(5817) <= (inputs(18)) or (inputs(240));
    layer0_outputs(5818) <= (inputs(43)) xor (inputs(53));
    layer0_outputs(5819) <= (inputs(218)) and not (inputs(125));
    layer0_outputs(5820) <= (inputs(43)) or (inputs(219));
    layer0_outputs(5821) <= (inputs(50)) or (inputs(87));
    layer0_outputs(5822) <= (inputs(36)) xor (inputs(68));
    layer0_outputs(5823) <= not((inputs(219)) xor (inputs(206)));
    layer0_outputs(5824) <= (inputs(95)) or (inputs(133));
    layer0_outputs(5825) <= not(inputs(56)) or (inputs(96));
    layer0_outputs(5826) <= not(inputs(134)) or (inputs(226));
    layer0_outputs(5827) <= (inputs(4)) and not (inputs(192));
    layer0_outputs(5828) <= not((inputs(198)) xor (inputs(204)));
    layer0_outputs(5829) <= not((inputs(41)) and (inputs(59)));
    layer0_outputs(5830) <= not((inputs(168)) or (inputs(17)));
    layer0_outputs(5831) <= (inputs(62)) and not (inputs(30));
    layer0_outputs(5832) <= (inputs(200)) and not (inputs(225));
    layer0_outputs(5833) <= not(inputs(118));
    layer0_outputs(5834) <= not(inputs(150)) or (inputs(228));
    layer0_outputs(5835) <= (inputs(8)) or (inputs(82));
    layer0_outputs(5836) <= not(inputs(149)) or (inputs(193));
    layer0_outputs(5837) <= not((inputs(130)) xor (inputs(185)));
    layer0_outputs(5838) <= (inputs(84)) and not (inputs(180));
    layer0_outputs(5839) <= not((inputs(64)) xor (inputs(159)));
    layer0_outputs(5840) <= not(inputs(127)) or (inputs(8));
    layer0_outputs(5841) <= (inputs(211)) or (inputs(144));
    layer0_outputs(5842) <= not(inputs(95)) or (inputs(223));
    layer0_outputs(5843) <= not(inputs(209)) or (inputs(111));
    layer0_outputs(5844) <= not(inputs(164));
    layer0_outputs(5845) <= (inputs(210)) or (inputs(50));
    layer0_outputs(5846) <= not((inputs(223)) xor (inputs(87)));
    layer0_outputs(5847) <= not(inputs(215)) or (inputs(127));
    layer0_outputs(5848) <= (inputs(135)) or (inputs(252));
    layer0_outputs(5849) <= (inputs(52)) or (inputs(224));
    layer0_outputs(5850) <= (inputs(26)) or (inputs(26));
    layer0_outputs(5851) <= (inputs(112)) or (inputs(235));
    layer0_outputs(5852) <= not(inputs(62));
    layer0_outputs(5853) <= (inputs(242)) and not (inputs(64));
    layer0_outputs(5854) <= not((inputs(3)) xor (inputs(162)));
    layer0_outputs(5855) <= (inputs(125)) or (inputs(134));
    layer0_outputs(5856) <= not((inputs(63)) or (inputs(60)));
    layer0_outputs(5857) <= not((inputs(114)) or (inputs(166)));
    layer0_outputs(5858) <= (inputs(212)) or (inputs(60));
    layer0_outputs(5859) <= not((inputs(28)) xor (inputs(219)));
    layer0_outputs(5860) <= (inputs(124)) xor (inputs(117));
    layer0_outputs(5861) <= (inputs(71)) and not (inputs(5));
    layer0_outputs(5862) <= not(inputs(175));
    layer0_outputs(5863) <= (inputs(84)) and not (inputs(248));
    layer0_outputs(5864) <= inputs(118);
    layer0_outputs(5865) <= not(inputs(73));
    layer0_outputs(5866) <= not(inputs(192)) or (inputs(33));
    layer0_outputs(5867) <= (inputs(203)) and not (inputs(250));
    layer0_outputs(5868) <= '0';
    layer0_outputs(5869) <= not(inputs(242)) or (inputs(15));
    layer0_outputs(5870) <= not(inputs(39)) or (inputs(225));
    layer0_outputs(5871) <= not((inputs(9)) or (inputs(101)));
    layer0_outputs(5872) <= (inputs(17)) xor (inputs(135));
    layer0_outputs(5873) <= not((inputs(205)) xor (inputs(11)));
    layer0_outputs(5874) <= inputs(97);
    layer0_outputs(5875) <= (inputs(52)) and (inputs(149));
    layer0_outputs(5876) <= inputs(229);
    layer0_outputs(5877) <= not(inputs(60)) or (inputs(64));
    layer0_outputs(5878) <= not((inputs(13)) xor (inputs(99)));
    layer0_outputs(5879) <= not(inputs(18));
    layer0_outputs(5880) <= inputs(156);
    layer0_outputs(5881) <= not((inputs(195)) xor (inputs(236)));
    layer0_outputs(5882) <= '0';
    layer0_outputs(5883) <= (inputs(103)) xor (inputs(70));
    layer0_outputs(5884) <= not((inputs(194)) xor (inputs(19)));
    layer0_outputs(5885) <= not(inputs(117)) or (inputs(114));
    layer0_outputs(5886) <= (inputs(70)) xor (inputs(183));
    layer0_outputs(5887) <= '1';
    layer0_outputs(5888) <= (inputs(101)) and not (inputs(248));
    layer0_outputs(5889) <= inputs(215);
    layer0_outputs(5890) <= (inputs(170)) and not (inputs(62));
    layer0_outputs(5891) <= (inputs(49)) xor (inputs(59));
    layer0_outputs(5892) <= inputs(123);
    layer0_outputs(5893) <= (inputs(38)) and not (inputs(175));
    layer0_outputs(5894) <= not(inputs(91)) or (inputs(235));
    layer0_outputs(5895) <= not((inputs(246)) xor (inputs(200)));
    layer0_outputs(5896) <= not((inputs(55)) or (inputs(68)));
    layer0_outputs(5897) <= not(inputs(16));
    layer0_outputs(5898) <= inputs(122);
    layer0_outputs(5899) <= (inputs(231)) or (inputs(129));
    layer0_outputs(5900) <= inputs(58);
    layer0_outputs(5901) <= not(inputs(135));
    layer0_outputs(5902) <= (inputs(108)) and not (inputs(25));
    layer0_outputs(5903) <= (inputs(30)) xor (inputs(217));
    layer0_outputs(5904) <= not(inputs(106));
    layer0_outputs(5905) <= not(inputs(164)) or (inputs(144));
    layer0_outputs(5906) <= '1';
    layer0_outputs(5907) <= not((inputs(207)) xor (inputs(232)));
    layer0_outputs(5908) <= inputs(137);
    layer0_outputs(5909) <= inputs(124);
    layer0_outputs(5910) <= (inputs(79)) or (inputs(117));
    layer0_outputs(5911) <= not(inputs(188)) or (inputs(223));
    layer0_outputs(5912) <= (inputs(41)) or (inputs(93));
    layer0_outputs(5913) <= not((inputs(36)) or (inputs(18)));
    layer0_outputs(5914) <= not(inputs(85));
    layer0_outputs(5915) <= (inputs(48)) xor (inputs(237));
    layer0_outputs(5916) <= inputs(85);
    layer0_outputs(5917) <= inputs(132);
    layer0_outputs(5918) <= not((inputs(105)) or (inputs(189)));
    layer0_outputs(5919) <= (inputs(18)) xor (inputs(160));
    layer0_outputs(5920) <= (inputs(253)) or (inputs(83));
    layer0_outputs(5921) <= inputs(247);
    layer0_outputs(5922) <= (inputs(42)) and not (inputs(250));
    layer0_outputs(5923) <= not(inputs(163)) or (inputs(65));
    layer0_outputs(5924) <= (inputs(146)) and not (inputs(7));
    layer0_outputs(5925) <= not((inputs(116)) xor (inputs(109)));
    layer0_outputs(5926) <= inputs(117);
    layer0_outputs(5927) <= not((inputs(84)) xor (inputs(229)));
    layer0_outputs(5928) <= (inputs(59)) and not (inputs(208));
    layer0_outputs(5929) <= '0';
    layer0_outputs(5930) <= (inputs(194)) and (inputs(81));
    layer0_outputs(5931) <= (inputs(252)) and (inputs(163));
    layer0_outputs(5932) <= (inputs(104)) or (inputs(27));
    layer0_outputs(5933) <= (inputs(23)) xor (inputs(18));
    layer0_outputs(5934) <= not((inputs(218)) xor (inputs(71)));
    layer0_outputs(5935) <= not(inputs(252)) or (inputs(23));
    layer0_outputs(5936) <= (inputs(235)) xor (inputs(18));
    layer0_outputs(5937) <= not((inputs(126)) or (inputs(116)));
    layer0_outputs(5938) <= '0';
    layer0_outputs(5939) <= (inputs(140)) or (inputs(114));
    layer0_outputs(5940) <= inputs(17);
    layer0_outputs(5941) <= not((inputs(125)) xor (inputs(226)));
    layer0_outputs(5942) <= '0';
    layer0_outputs(5943) <= inputs(202);
    layer0_outputs(5944) <= (inputs(114)) and not (inputs(125));
    layer0_outputs(5945) <= (inputs(252)) and not (inputs(128));
    layer0_outputs(5946) <= not(inputs(19));
    layer0_outputs(5947) <= (inputs(88)) xor (inputs(131));
    layer0_outputs(5948) <= not(inputs(120)) or (inputs(101));
    layer0_outputs(5949) <= not(inputs(26));
    layer0_outputs(5950) <= not((inputs(127)) and (inputs(41)));
    layer0_outputs(5951) <= inputs(85);
    layer0_outputs(5952) <= (inputs(115)) xor (inputs(100));
    layer0_outputs(5953) <= (inputs(127)) and not (inputs(2));
    layer0_outputs(5954) <= (inputs(83)) and not (inputs(174));
    layer0_outputs(5955) <= (inputs(3)) or (inputs(171));
    layer0_outputs(5956) <= not(inputs(214));
    layer0_outputs(5957) <= (inputs(126)) and not (inputs(158));
    layer0_outputs(5958) <= (inputs(163)) and not (inputs(253));
    layer0_outputs(5959) <= inputs(131);
    layer0_outputs(5960) <= (inputs(231)) and not (inputs(128));
    layer0_outputs(5961) <= inputs(25);
    layer0_outputs(5962) <= (inputs(89)) and not (inputs(87));
    layer0_outputs(5963) <= not((inputs(168)) xor (inputs(107)));
    layer0_outputs(5964) <= not(inputs(246)) or (inputs(160));
    layer0_outputs(5965) <= not((inputs(7)) xor (inputs(5)));
    layer0_outputs(5966) <= not((inputs(210)) or (inputs(6)));
    layer0_outputs(5967) <= (inputs(60)) xor (inputs(222));
    layer0_outputs(5968) <= (inputs(129)) and not (inputs(112));
    layer0_outputs(5969) <= not(inputs(90));
    layer0_outputs(5970) <= not(inputs(21));
    layer0_outputs(5971) <= (inputs(157)) or (inputs(114));
    layer0_outputs(5972) <= (inputs(148)) and not (inputs(0));
    layer0_outputs(5973) <= (inputs(253)) or (inputs(155));
    layer0_outputs(5974) <= not(inputs(153));
    layer0_outputs(5975) <= inputs(218);
    layer0_outputs(5976) <= not((inputs(188)) or (inputs(56)));
    layer0_outputs(5977) <= (inputs(9)) or (inputs(112));
    layer0_outputs(5978) <= (inputs(207)) and not (inputs(251));
    layer0_outputs(5979) <= inputs(72);
    layer0_outputs(5980) <= (inputs(157)) and not (inputs(192));
    layer0_outputs(5981) <= (inputs(129)) and not (inputs(174));
    layer0_outputs(5982) <= (inputs(229)) xor (inputs(34));
    layer0_outputs(5983) <= '0';
    layer0_outputs(5984) <= not(inputs(168));
    layer0_outputs(5985) <= not(inputs(149));
    layer0_outputs(5986) <= not(inputs(52)) or (inputs(125));
    layer0_outputs(5987) <= not(inputs(183));
    layer0_outputs(5988) <= not(inputs(5)) or (inputs(7));
    layer0_outputs(5989) <= (inputs(148)) or (inputs(86));
    layer0_outputs(5990) <= inputs(150);
    layer0_outputs(5991) <= not(inputs(120));
    layer0_outputs(5992) <= not((inputs(172)) or (inputs(183)));
    layer0_outputs(5993) <= inputs(39);
    layer0_outputs(5994) <= (inputs(73)) or (inputs(67));
    layer0_outputs(5995) <= not((inputs(72)) or (inputs(124)));
    layer0_outputs(5996) <= inputs(241);
    layer0_outputs(5997) <= not((inputs(125)) xor (inputs(193)));
    layer0_outputs(5998) <= (inputs(240)) or (inputs(100));
    layer0_outputs(5999) <= not(inputs(107)) or (inputs(63));
    layer0_outputs(6000) <= not((inputs(16)) and (inputs(193)));
    layer0_outputs(6001) <= (inputs(148)) or (inputs(158));
    layer0_outputs(6002) <= inputs(118);
    layer0_outputs(6003) <= not((inputs(216)) or (inputs(241)));
    layer0_outputs(6004) <= not((inputs(238)) or (inputs(0)));
    layer0_outputs(6005) <= '0';
    layer0_outputs(6006) <= not(inputs(235)) or (inputs(28));
    layer0_outputs(6007) <= (inputs(18)) or (inputs(52));
    layer0_outputs(6008) <= inputs(182);
    layer0_outputs(6009) <= (inputs(69)) xor (inputs(14));
    layer0_outputs(6010) <= (inputs(202)) or (inputs(19));
    layer0_outputs(6011) <= (inputs(204)) or (inputs(21));
    layer0_outputs(6012) <= (inputs(71)) and not (inputs(193));
    layer0_outputs(6013) <= (inputs(154)) and (inputs(178));
    layer0_outputs(6014) <= not((inputs(20)) or (inputs(172)));
    layer0_outputs(6015) <= not(inputs(140));
    layer0_outputs(6016) <= (inputs(31)) and (inputs(22));
    layer0_outputs(6017) <= not((inputs(187)) or (inputs(204)));
    layer0_outputs(6018) <= (inputs(242)) and not (inputs(112));
    layer0_outputs(6019) <= not((inputs(226)) xor (inputs(125)));
    layer0_outputs(6020) <= inputs(168);
    layer0_outputs(6021) <= inputs(206);
    layer0_outputs(6022) <= inputs(215);
    layer0_outputs(6023) <= not((inputs(143)) and (inputs(197)));
    layer0_outputs(6024) <= not(inputs(137));
    layer0_outputs(6025) <= '0';
    layer0_outputs(6026) <= '1';
    layer0_outputs(6027) <= (inputs(96)) xor (inputs(123));
    layer0_outputs(6028) <= (inputs(21)) and not (inputs(143));
    layer0_outputs(6029) <= not((inputs(126)) or (inputs(240)));
    layer0_outputs(6030) <= not((inputs(233)) or (inputs(127)));
    layer0_outputs(6031) <= (inputs(101)) and not (inputs(91));
    layer0_outputs(6032) <= inputs(108);
    layer0_outputs(6033) <= inputs(61);
    layer0_outputs(6034) <= not((inputs(224)) or (inputs(240)));
    layer0_outputs(6035) <= (inputs(250)) xor (inputs(219));
    layer0_outputs(6036) <= not(inputs(26));
    layer0_outputs(6037) <= (inputs(229)) or (inputs(20));
    layer0_outputs(6038) <= not(inputs(188)) or (inputs(11));
    layer0_outputs(6039) <= (inputs(165)) or (inputs(37));
    layer0_outputs(6040) <= not((inputs(87)) or (inputs(246)));
    layer0_outputs(6041) <= (inputs(211)) and (inputs(193));
    layer0_outputs(6042) <= (inputs(162)) or (inputs(92));
    layer0_outputs(6043) <= not(inputs(104));
    layer0_outputs(6044) <= not((inputs(157)) xor (inputs(95)));
    layer0_outputs(6045) <= (inputs(17)) xor (inputs(70));
    layer0_outputs(6046) <= inputs(232);
    layer0_outputs(6047) <= inputs(147);
    layer0_outputs(6048) <= (inputs(196)) and (inputs(65));
    layer0_outputs(6049) <= (inputs(101)) and not (inputs(92));
    layer0_outputs(6050) <= not((inputs(101)) or (inputs(11)));
    layer0_outputs(6051) <= (inputs(145)) xor (inputs(124));
    layer0_outputs(6052) <= '1';
    layer0_outputs(6053) <= (inputs(244)) xor (inputs(130));
    layer0_outputs(6054) <= (inputs(88)) or (inputs(109));
    layer0_outputs(6055) <= not(inputs(1));
    layer0_outputs(6056) <= (inputs(229)) xor (inputs(139));
    layer0_outputs(6057) <= (inputs(51)) and not (inputs(22));
    layer0_outputs(6058) <= inputs(106);
    layer0_outputs(6059) <= (inputs(6)) and not (inputs(23));
    layer0_outputs(6060) <= not((inputs(192)) or (inputs(39)));
    layer0_outputs(6061) <= (inputs(175)) and (inputs(124));
    layer0_outputs(6062) <= not((inputs(106)) xor (inputs(250)));
    layer0_outputs(6063) <= (inputs(198)) xor (inputs(129));
    layer0_outputs(6064) <= inputs(26);
    layer0_outputs(6065) <= not(inputs(25));
    layer0_outputs(6066) <= (inputs(45)) or (inputs(114));
    layer0_outputs(6067) <= not((inputs(150)) xor (inputs(213)));
    layer0_outputs(6068) <= (inputs(131)) and (inputs(174));
    layer0_outputs(6069) <= not((inputs(182)) xor (inputs(104)));
    layer0_outputs(6070) <= '1';
    layer0_outputs(6071) <= (inputs(191)) or (inputs(115));
    layer0_outputs(6072) <= inputs(92);
    layer0_outputs(6073) <= not((inputs(65)) or (inputs(171)));
    layer0_outputs(6074) <= not((inputs(113)) xor (inputs(185)));
    layer0_outputs(6075) <= not(inputs(202));
    layer0_outputs(6076) <= not(inputs(134));
    layer0_outputs(6077) <= (inputs(173)) xor (inputs(181));
    layer0_outputs(6078) <= not((inputs(105)) and (inputs(183)));
    layer0_outputs(6079) <= not((inputs(213)) xor (inputs(182)));
    layer0_outputs(6080) <= not(inputs(170));
    layer0_outputs(6081) <= not(inputs(44));
    layer0_outputs(6082) <= not(inputs(133)) or (inputs(72));
    layer0_outputs(6083) <= (inputs(138)) xor (inputs(7));
    layer0_outputs(6084) <= (inputs(169)) xor (inputs(202));
    layer0_outputs(6085) <= not(inputs(4)) or (inputs(113));
    layer0_outputs(6086) <= not(inputs(182)) or (inputs(179));
    layer0_outputs(6087) <= not(inputs(132));
    layer0_outputs(6088) <= (inputs(210)) and not (inputs(12));
    layer0_outputs(6089) <= not(inputs(131)) or (inputs(231));
    layer0_outputs(6090) <= not((inputs(125)) xor (inputs(155)));
    layer0_outputs(6091) <= (inputs(26)) xor (inputs(167));
    layer0_outputs(6092) <= not((inputs(209)) xor (inputs(143)));
    layer0_outputs(6093) <= not((inputs(252)) xor (inputs(239)));
    layer0_outputs(6094) <= inputs(201);
    layer0_outputs(6095) <= '1';
    layer0_outputs(6096) <= (inputs(209)) or (inputs(182));
    layer0_outputs(6097) <= (inputs(134)) and not (inputs(19));
    layer0_outputs(6098) <= not(inputs(148)) or (inputs(247));
    layer0_outputs(6099) <= (inputs(236)) and not (inputs(51));
    layer0_outputs(6100) <= not(inputs(153)) or (inputs(80));
    layer0_outputs(6101) <= not((inputs(207)) or (inputs(152)));
    layer0_outputs(6102) <= not(inputs(241));
    layer0_outputs(6103) <= not((inputs(55)) xor (inputs(84)));
    layer0_outputs(6104) <= '1';
    layer0_outputs(6105) <= (inputs(195)) xor (inputs(158));
    layer0_outputs(6106) <= not(inputs(46));
    layer0_outputs(6107) <= not(inputs(55));
    layer0_outputs(6108) <= (inputs(123)) or (inputs(153));
    layer0_outputs(6109) <= inputs(93);
    layer0_outputs(6110) <= (inputs(249)) and not (inputs(221));
    layer0_outputs(6111) <= (inputs(96)) or (inputs(166));
    layer0_outputs(6112) <= (inputs(216)) or (inputs(156));
    layer0_outputs(6113) <= not((inputs(131)) xor (inputs(80)));
    layer0_outputs(6114) <= not(inputs(90)) or (inputs(29));
    layer0_outputs(6115) <= not((inputs(172)) xor (inputs(111)));
    layer0_outputs(6116) <= (inputs(251)) and not (inputs(53));
    layer0_outputs(6117) <= inputs(96);
    layer0_outputs(6118) <= inputs(119);
    layer0_outputs(6119) <= not(inputs(111)) or (inputs(30));
    layer0_outputs(6120) <= not(inputs(2));
    layer0_outputs(6121) <= (inputs(185)) and not (inputs(91));
    layer0_outputs(6122) <= not((inputs(173)) or (inputs(82)));
    layer0_outputs(6123) <= not((inputs(61)) or (inputs(140)));
    layer0_outputs(6124) <= '1';
    layer0_outputs(6125) <= not((inputs(141)) or (inputs(48)));
    layer0_outputs(6126) <= (inputs(38)) or (inputs(82));
    layer0_outputs(6127) <= not(inputs(24));
    layer0_outputs(6128) <= (inputs(91)) or (inputs(26));
    layer0_outputs(6129) <= (inputs(239)) xor (inputs(68));
    layer0_outputs(6130) <= (inputs(238)) or (inputs(132));
    layer0_outputs(6131) <= not((inputs(170)) xor (inputs(35)));
    layer0_outputs(6132) <= not((inputs(63)) xor (inputs(25)));
    layer0_outputs(6133) <= not(inputs(120));
    layer0_outputs(6134) <= not(inputs(137)) or (inputs(119));
    layer0_outputs(6135) <= not((inputs(65)) or (inputs(32)));
    layer0_outputs(6136) <= (inputs(111)) or (inputs(126));
    layer0_outputs(6137) <= (inputs(157)) or (inputs(246));
    layer0_outputs(6138) <= not((inputs(137)) or (inputs(121)));
    layer0_outputs(6139) <= (inputs(131)) and not (inputs(13));
    layer0_outputs(6140) <= (inputs(98)) xor (inputs(248));
    layer0_outputs(6141) <= not((inputs(237)) xor (inputs(195)));
    layer0_outputs(6142) <= not(inputs(75)) or (inputs(148));
    layer0_outputs(6143) <= (inputs(75)) or (inputs(33));
    layer0_outputs(6144) <= (inputs(102)) and not (inputs(27));
    layer0_outputs(6145) <= not((inputs(141)) xor (inputs(77)));
    layer0_outputs(6146) <= not((inputs(242)) xor (inputs(128)));
    layer0_outputs(6147) <= not((inputs(112)) or (inputs(0)));
    layer0_outputs(6148) <= not((inputs(1)) and (inputs(34)));
    layer0_outputs(6149) <= (inputs(23)) xor (inputs(221));
    layer0_outputs(6150) <= not(inputs(136));
    layer0_outputs(6151) <= (inputs(215)) and not (inputs(16));
    layer0_outputs(6152) <= not((inputs(76)) or (inputs(61)));
    layer0_outputs(6153) <= (inputs(55)) and not (inputs(116));
    layer0_outputs(6154) <= inputs(182);
    layer0_outputs(6155) <= inputs(6);
    layer0_outputs(6156) <= not(inputs(111));
    layer0_outputs(6157) <= not(inputs(103));
    layer0_outputs(6158) <= (inputs(173)) xor (inputs(196));
    layer0_outputs(6159) <= not((inputs(182)) xor (inputs(162)));
    layer0_outputs(6160) <= inputs(179);
    layer0_outputs(6161) <= not((inputs(13)) xor (inputs(152)));
    layer0_outputs(6162) <= not(inputs(239)) or (inputs(203));
    layer0_outputs(6163) <= not((inputs(88)) or (inputs(112)));
    layer0_outputs(6164) <= not(inputs(100)) or (inputs(225));
    layer0_outputs(6165) <= (inputs(227)) xor (inputs(123));
    layer0_outputs(6166) <= (inputs(120)) or (inputs(217));
    layer0_outputs(6167) <= not(inputs(194)) or (inputs(139));
    layer0_outputs(6168) <= not(inputs(182)) or (inputs(80));
    layer0_outputs(6169) <= (inputs(196)) and not (inputs(179));
    layer0_outputs(6170) <= (inputs(2)) or (inputs(111));
    layer0_outputs(6171) <= (inputs(156)) and not (inputs(128));
    layer0_outputs(6172) <= not(inputs(185));
    layer0_outputs(6173) <= (inputs(78)) or (inputs(167));
    layer0_outputs(6174) <= not((inputs(14)) xor (inputs(141)));
    layer0_outputs(6175) <= (inputs(189)) or (inputs(56));
    layer0_outputs(6176) <= not((inputs(227)) and (inputs(1)));
    layer0_outputs(6177) <= not((inputs(43)) or (inputs(152)));
    layer0_outputs(6178) <= not((inputs(222)) or (inputs(236)));
    layer0_outputs(6179) <= (inputs(159)) and not (inputs(44));
    layer0_outputs(6180) <= not((inputs(216)) xor (inputs(58)));
    layer0_outputs(6181) <= (inputs(190)) or (inputs(151));
    layer0_outputs(6182) <= (inputs(54)) or (inputs(121));
    layer0_outputs(6183) <= not((inputs(239)) xor (inputs(250)));
    layer0_outputs(6184) <= inputs(141);
    layer0_outputs(6185) <= inputs(120);
    layer0_outputs(6186) <= '1';
    layer0_outputs(6187) <= inputs(60);
    layer0_outputs(6188) <= not(inputs(43)) or (inputs(77));
    layer0_outputs(6189) <= not(inputs(154)) or (inputs(39));
    layer0_outputs(6190) <= (inputs(13)) or (inputs(181));
    layer0_outputs(6191) <= not(inputs(168)) or (inputs(249));
    layer0_outputs(6192) <= (inputs(99)) and not (inputs(255));
    layer0_outputs(6193) <= (inputs(166)) or (inputs(156));
    layer0_outputs(6194) <= (inputs(161)) xor (inputs(220));
    layer0_outputs(6195) <= not(inputs(199));
    layer0_outputs(6196) <= (inputs(242)) xor (inputs(255));
    layer0_outputs(6197) <= (inputs(67)) and not (inputs(32));
    layer0_outputs(6198) <= not((inputs(32)) or (inputs(31)));
    layer0_outputs(6199) <= inputs(158);
    layer0_outputs(6200) <= not(inputs(92));
    layer0_outputs(6201) <= not(inputs(103));
    layer0_outputs(6202) <= not((inputs(91)) and (inputs(204)));
    layer0_outputs(6203) <= not((inputs(230)) xor (inputs(145)));
    layer0_outputs(6204) <= not(inputs(113));
    layer0_outputs(6205) <= (inputs(132)) xor (inputs(133));
    layer0_outputs(6206) <= (inputs(235)) and not (inputs(1));
    layer0_outputs(6207) <= '0';
    layer0_outputs(6208) <= not(inputs(152));
    layer0_outputs(6209) <= not((inputs(166)) or (inputs(220)));
    layer0_outputs(6210) <= not((inputs(165)) or (inputs(246)));
    layer0_outputs(6211) <= not(inputs(245)) or (inputs(29));
    layer0_outputs(6212) <= not((inputs(40)) or (inputs(147)));
    layer0_outputs(6213) <= not(inputs(22));
    layer0_outputs(6214) <= inputs(134);
    layer0_outputs(6215) <= not(inputs(57));
    layer0_outputs(6216) <= not(inputs(41)) or (inputs(250));
    layer0_outputs(6217) <= (inputs(106)) or (inputs(138));
    layer0_outputs(6218) <= (inputs(72)) and (inputs(160));
    layer0_outputs(6219) <= (inputs(156)) or (inputs(102));
    layer0_outputs(6220) <= not(inputs(157)) or (inputs(96));
    layer0_outputs(6221) <= (inputs(126)) xor (inputs(250));
    layer0_outputs(6222) <= (inputs(216)) and not (inputs(234));
    layer0_outputs(6223) <= not((inputs(134)) or (inputs(175)));
    layer0_outputs(6224) <= inputs(133);
    layer0_outputs(6225) <= not((inputs(74)) xor (inputs(185)));
    layer0_outputs(6226) <= not(inputs(232));
    layer0_outputs(6227) <= not(inputs(201)) or (inputs(113));
    layer0_outputs(6228) <= (inputs(165)) or (inputs(148));
    layer0_outputs(6229) <= '0';
    layer0_outputs(6230) <= (inputs(33)) or (inputs(173));
    layer0_outputs(6231) <= not((inputs(198)) xor (inputs(198)));
    layer0_outputs(6232) <= not((inputs(130)) or (inputs(147)));
    layer0_outputs(6233) <= (inputs(93)) or (inputs(215));
    layer0_outputs(6234) <= (inputs(29)) and not (inputs(252));
    layer0_outputs(6235) <= not((inputs(203)) xor (inputs(247)));
    layer0_outputs(6236) <= not(inputs(196));
    layer0_outputs(6237) <= inputs(110);
    layer0_outputs(6238) <= not(inputs(116)) or (inputs(215));
    layer0_outputs(6239) <= not(inputs(99)) or (inputs(173));
    layer0_outputs(6240) <= (inputs(102)) xor (inputs(12));
    layer0_outputs(6241) <= not(inputs(194)) or (inputs(33));
    layer0_outputs(6242) <= (inputs(214)) or (inputs(5));
    layer0_outputs(6243) <= not((inputs(235)) or (inputs(4)));
    layer0_outputs(6244) <= inputs(1);
    layer0_outputs(6245) <= not(inputs(131)) or (inputs(169));
    layer0_outputs(6246) <= not((inputs(107)) xor (inputs(179)));
    layer0_outputs(6247) <= inputs(70);
    layer0_outputs(6248) <= inputs(62);
    layer0_outputs(6249) <= not((inputs(121)) and (inputs(152)));
    layer0_outputs(6250) <= (inputs(168)) and not (inputs(34));
    layer0_outputs(6251) <= not((inputs(142)) or (inputs(84)));
    layer0_outputs(6252) <= inputs(132);
    layer0_outputs(6253) <= not((inputs(213)) xor (inputs(26)));
    layer0_outputs(6254) <= (inputs(179)) or (inputs(90));
    layer0_outputs(6255) <= (inputs(94)) xor (inputs(57));
    layer0_outputs(6256) <= not(inputs(186));
    layer0_outputs(6257) <= not(inputs(35)) or (inputs(63));
    layer0_outputs(6258) <= not(inputs(229));
    layer0_outputs(6259) <= not((inputs(122)) xor (inputs(31)));
    layer0_outputs(6260) <= not((inputs(186)) or (inputs(102)));
    layer0_outputs(6261) <= inputs(181);
    layer0_outputs(6262) <= '0';
    layer0_outputs(6263) <= not(inputs(133)) or (inputs(38));
    layer0_outputs(6264) <= (inputs(105)) or (inputs(64));
    layer0_outputs(6265) <= (inputs(116)) and not (inputs(47));
    layer0_outputs(6266) <= not(inputs(36));
    layer0_outputs(6267) <= (inputs(202)) and not (inputs(52));
    layer0_outputs(6268) <= (inputs(160)) xor (inputs(249));
    layer0_outputs(6269) <= (inputs(105)) xor (inputs(83));
    layer0_outputs(6270) <= (inputs(216)) or (inputs(35));
    layer0_outputs(6271) <= inputs(77);
    layer0_outputs(6272) <= (inputs(133)) and not (inputs(222));
    layer0_outputs(6273) <= inputs(89);
    layer0_outputs(6274) <= not(inputs(31)) or (inputs(177));
    layer0_outputs(6275) <= (inputs(118)) and not (inputs(112));
    layer0_outputs(6276) <= not(inputs(16)) or (inputs(44));
    layer0_outputs(6277) <= not((inputs(69)) xor (inputs(41)));
    layer0_outputs(6278) <= '1';
    layer0_outputs(6279) <= not((inputs(102)) and (inputs(167)));
    layer0_outputs(6280) <= (inputs(186)) and not (inputs(174));
    layer0_outputs(6281) <= (inputs(212)) or (inputs(148));
    layer0_outputs(6282) <= not(inputs(196));
    layer0_outputs(6283) <= not((inputs(97)) or (inputs(14)));
    layer0_outputs(6284) <= (inputs(157)) and not (inputs(211));
    layer0_outputs(6285) <= not(inputs(13)) or (inputs(247));
    layer0_outputs(6286) <= inputs(130);
    layer0_outputs(6287) <= not(inputs(212));
    layer0_outputs(6288) <= not(inputs(187)) or (inputs(209));
    layer0_outputs(6289) <= not(inputs(117)) or (inputs(39));
    layer0_outputs(6290) <= inputs(232);
    layer0_outputs(6291) <= (inputs(145)) xor (inputs(105));
    layer0_outputs(6292) <= not((inputs(164)) xor (inputs(181)));
    layer0_outputs(6293) <= (inputs(61)) xor (inputs(225));
    layer0_outputs(6294) <= not(inputs(250)) or (inputs(131));
    layer0_outputs(6295) <= not((inputs(172)) or (inputs(37)));
    layer0_outputs(6296) <= inputs(152);
    layer0_outputs(6297) <= not(inputs(69)) or (inputs(60));
    layer0_outputs(6298) <= (inputs(253)) or (inputs(219));
    layer0_outputs(6299) <= (inputs(180)) xor (inputs(61));
    layer0_outputs(6300) <= (inputs(100)) or (inputs(80));
    layer0_outputs(6301) <= (inputs(110)) xor (inputs(190));
    layer0_outputs(6302) <= not((inputs(254)) xor (inputs(106)));
    layer0_outputs(6303) <= inputs(142);
    layer0_outputs(6304) <= not((inputs(58)) xor (inputs(127)));
    layer0_outputs(6305) <= (inputs(254)) or (inputs(161));
    layer0_outputs(6306) <= not((inputs(47)) or (inputs(140)));
    layer0_outputs(6307) <= (inputs(25)) or (inputs(189));
    layer0_outputs(6308) <= not((inputs(48)) xor (inputs(205)));
    layer0_outputs(6309) <= not((inputs(213)) or (inputs(76)));
    layer0_outputs(6310) <= (inputs(82)) and not (inputs(47));
    layer0_outputs(6311) <= inputs(136);
    layer0_outputs(6312) <= not((inputs(177)) xor (inputs(66)));
    layer0_outputs(6313) <= (inputs(231)) or (inputs(247));
    layer0_outputs(6314) <= not((inputs(47)) xor (inputs(105)));
    layer0_outputs(6315) <= not((inputs(124)) or (inputs(93)));
    layer0_outputs(6316) <= (inputs(182)) and not (inputs(123));
    layer0_outputs(6317) <= (inputs(117)) or (inputs(33));
    layer0_outputs(6318) <= not((inputs(39)) or (inputs(255)));
    layer0_outputs(6319) <= (inputs(62)) or (inputs(216));
    layer0_outputs(6320) <= '1';
    layer0_outputs(6321) <= not((inputs(43)) xor (inputs(38)));
    layer0_outputs(6322) <= (inputs(66)) or (inputs(213));
    layer0_outputs(6323) <= not((inputs(73)) xor (inputs(3)));
    layer0_outputs(6324) <= (inputs(186)) xor (inputs(204));
    layer0_outputs(6325) <= not((inputs(16)) xor (inputs(173)));
    layer0_outputs(6326) <= not(inputs(216));
    layer0_outputs(6327) <= not(inputs(150));
    layer0_outputs(6328) <= not((inputs(250)) or (inputs(0)));
    layer0_outputs(6329) <= not(inputs(71)) or (inputs(50));
    layer0_outputs(6330) <= '0';
    layer0_outputs(6331) <= (inputs(123)) and not (inputs(64));
    layer0_outputs(6332) <= inputs(124);
    layer0_outputs(6333) <= inputs(102);
    layer0_outputs(6334) <= (inputs(127)) or (inputs(165));
    layer0_outputs(6335) <= (inputs(1)) and (inputs(249));
    layer0_outputs(6336) <= not(inputs(98));
    layer0_outputs(6337) <= not(inputs(102)) or (inputs(48));
    layer0_outputs(6338) <= '1';
    layer0_outputs(6339) <= (inputs(111)) and not (inputs(44));
    layer0_outputs(6340) <= not((inputs(6)) and (inputs(47)));
    layer0_outputs(6341) <= not(inputs(208));
    layer0_outputs(6342) <= not((inputs(25)) and (inputs(254)));
    layer0_outputs(6343) <= (inputs(60)) xor (inputs(63));
    layer0_outputs(6344) <= not(inputs(20)) or (inputs(4));
    layer0_outputs(6345) <= not((inputs(147)) xor (inputs(34)));
    layer0_outputs(6346) <= (inputs(24)) and not (inputs(82));
    layer0_outputs(6347) <= not(inputs(107));
    layer0_outputs(6348) <= not(inputs(238)) or (inputs(214));
    layer0_outputs(6349) <= (inputs(66)) and not (inputs(236));
    layer0_outputs(6350) <= inputs(57);
    layer0_outputs(6351) <= not((inputs(3)) xor (inputs(155)));
    layer0_outputs(6352) <= not((inputs(194)) xor (inputs(71)));
    layer0_outputs(6353) <= (inputs(26)) and (inputs(245));
    layer0_outputs(6354) <= not(inputs(26));
    layer0_outputs(6355) <= inputs(61);
    layer0_outputs(6356) <= not((inputs(195)) or (inputs(205)));
    layer0_outputs(6357) <= '0';
    layer0_outputs(6358) <= (inputs(185)) and not (inputs(145));
    layer0_outputs(6359) <= not((inputs(235)) or (inputs(24)));
    layer0_outputs(6360) <= inputs(149);
    layer0_outputs(6361) <= inputs(138);
    layer0_outputs(6362) <= not((inputs(196)) or (inputs(74)));
    layer0_outputs(6363) <= (inputs(55)) and not (inputs(172));
    layer0_outputs(6364) <= not(inputs(248));
    layer0_outputs(6365) <= not(inputs(57));
    layer0_outputs(6366) <= not(inputs(56));
    layer0_outputs(6367) <= not(inputs(102)) or (inputs(33));
    layer0_outputs(6368) <= (inputs(38)) and (inputs(246));
    layer0_outputs(6369) <= inputs(182);
    layer0_outputs(6370) <= (inputs(252)) or (inputs(160));
    layer0_outputs(6371) <= not(inputs(198)) or (inputs(203));
    layer0_outputs(6372) <= not((inputs(69)) or (inputs(46)));
    layer0_outputs(6373) <= (inputs(77)) and not (inputs(66));
    layer0_outputs(6374) <= (inputs(214)) or (inputs(108));
    layer0_outputs(6375) <= not(inputs(164)) or (inputs(236));
    layer0_outputs(6376) <= (inputs(220)) xor (inputs(69));
    layer0_outputs(6377) <= (inputs(100)) and not (inputs(211));
    layer0_outputs(6378) <= (inputs(117)) and not (inputs(50));
    layer0_outputs(6379) <= not(inputs(163)) or (inputs(80));
    layer0_outputs(6380) <= (inputs(243)) or (inputs(120));
    layer0_outputs(6381) <= not((inputs(74)) or (inputs(36)));
    layer0_outputs(6382) <= not(inputs(141));
    layer0_outputs(6383) <= '1';
    layer0_outputs(6384) <= inputs(217);
    layer0_outputs(6385) <= inputs(17);
    layer0_outputs(6386) <= not((inputs(210)) or (inputs(101)));
    layer0_outputs(6387) <= (inputs(216)) xor (inputs(239));
    layer0_outputs(6388) <= not((inputs(181)) or (inputs(143)));
    layer0_outputs(6389) <= (inputs(182)) xor (inputs(130));
    layer0_outputs(6390) <= not(inputs(202)) or (inputs(22));
    layer0_outputs(6391) <= (inputs(213)) and not (inputs(171));
    layer0_outputs(6392) <= not(inputs(73)) or (inputs(245));
    layer0_outputs(6393) <= (inputs(100)) or (inputs(80));
    layer0_outputs(6394) <= not(inputs(67)) or (inputs(177));
    layer0_outputs(6395) <= not(inputs(100));
    layer0_outputs(6396) <= not(inputs(80)) or (inputs(95));
    layer0_outputs(6397) <= not(inputs(230));
    layer0_outputs(6398) <= not(inputs(25));
    layer0_outputs(6399) <= (inputs(214)) and not (inputs(240));
    layer0_outputs(6400) <= not(inputs(41)) or (inputs(129));
    layer0_outputs(6401) <= not(inputs(100)) or (inputs(18));
    layer0_outputs(6402) <= (inputs(228)) xor (inputs(160));
    layer0_outputs(6403) <= (inputs(43)) or (inputs(132));
    layer0_outputs(6404) <= not(inputs(120)) or (inputs(45));
    layer0_outputs(6405) <= (inputs(247)) or (inputs(195));
    layer0_outputs(6406) <= (inputs(26)) xor (inputs(220));
    layer0_outputs(6407) <= (inputs(172)) xor (inputs(41));
    layer0_outputs(6408) <= (inputs(126)) or (inputs(161));
    layer0_outputs(6409) <= inputs(202);
    layer0_outputs(6410) <= inputs(194);
    layer0_outputs(6411) <= (inputs(105)) and not (inputs(158));
    layer0_outputs(6412) <= (inputs(160)) or (inputs(35));
    layer0_outputs(6413) <= (inputs(168)) and not (inputs(184));
    layer0_outputs(6414) <= not((inputs(214)) xor (inputs(241)));
    layer0_outputs(6415) <= not(inputs(206)) or (inputs(211));
    layer0_outputs(6416) <= inputs(40);
    layer0_outputs(6417) <= not((inputs(117)) or (inputs(52)));
    layer0_outputs(6418) <= not((inputs(245)) xor (inputs(156)));
    layer0_outputs(6419) <= not((inputs(211)) xor (inputs(98)));
    layer0_outputs(6420) <= not((inputs(214)) or (inputs(234)));
    layer0_outputs(6421) <= not(inputs(22)) or (inputs(190));
    layer0_outputs(6422) <= not((inputs(144)) or (inputs(206)));
    layer0_outputs(6423) <= not(inputs(138)) or (inputs(242));
    layer0_outputs(6424) <= not((inputs(83)) or (inputs(181)));
    layer0_outputs(6425) <= (inputs(88)) and not (inputs(242));
    layer0_outputs(6426) <= (inputs(41)) or (inputs(212));
    layer0_outputs(6427) <= not((inputs(80)) xor (inputs(14)));
    layer0_outputs(6428) <= not((inputs(5)) and (inputs(212)));
    layer0_outputs(6429) <= not(inputs(14));
    layer0_outputs(6430) <= not(inputs(150));
    layer0_outputs(6431) <= not(inputs(176)) or (inputs(13));
    layer0_outputs(6432) <= (inputs(61)) and not (inputs(39));
    layer0_outputs(6433) <= (inputs(4)) or (inputs(126));
    layer0_outputs(6434) <= '1';
    layer0_outputs(6435) <= not((inputs(91)) or (inputs(144)));
    layer0_outputs(6436) <= (inputs(176)) or (inputs(178));
    layer0_outputs(6437) <= not(inputs(149)) or (inputs(210));
    layer0_outputs(6438) <= not((inputs(194)) or (inputs(219)));
    layer0_outputs(6439) <= not(inputs(109)) or (inputs(13));
    layer0_outputs(6440) <= inputs(109);
    layer0_outputs(6441) <= not(inputs(88));
    layer0_outputs(6442) <= not(inputs(85)) or (inputs(16));
    layer0_outputs(6443) <= not(inputs(54));
    layer0_outputs(6444) <= (inputs(77)) or (inputs(147));
    layer0_outputs(6445) <= (inputs(192)) xor (inputs(179));
    layer0_outputs(6446) <= not(inputs(182));
    layer0_outputs(6447) <= inputs(107);
    layer0_outputs(6448) <= not(inputs(82)) or (inputs(18));
    layer0_outputs(6449) <= not((inputs(69)) or (inputs(20)));
    layer0_outputs(6450) <= (inputs(185)) or (inputs(50));
    layer0_outputs(6451) <= not(inputs(150)) or (inputs(16));
    layer0_outputs(6452) <= (inputs(209)) or (inputs(197));
    layer0_outputs(6453) <= not((inputs(0)) or (inputs(66)));
    layer0_outputs(6454) <= (inputs(224)) xor (inputs(206));
    layer0_outputs(6455) <= not((inputs(167)) xor (inputs(21)));
    layer0_outputs(6456) <= inputs(80);
    layer0_outputs(6457) <= (inputs(26)) xor (inputs(155));
    layer0_outputs(6458) <= inputs(232);
    layer0_outputs(6459) <= (inputs(216)) and not (inputs(249));
    layer0_outputs(6460) <= not(inputs(179)) or (inputs(220));
    layer0_outputs(6461) <= (inputs(205)) or (inputs(206));
    layer0_outputs(6462) <= (inputs(140)) and (inputs(132));
    layer0_outputs(6463) <= not((inputs(165)) xor (inputs(33)));
    layer0_outputs(6464) <= (inputs(207)) xor (inputs(206));
    layer0_outputs(6465) <= not(inputs(198));
    layer0_outputs(6466) <= (inputs(133)) and not (inputs(14));
    layer0_outputs(6467) <= not((inputs(252)) xor (inputs(169)));
    layer0_outputs(6468) <= not(inputs(195)) or (inputs(228));
    layer0_outputs(6469) <= not((inputs(192)) and (inputs(217)));
    layer0_outputs(6470) <= inputs(135);
    layer0_outputs(6471) <= inputs(171);
    layer0_outputs(6472) <= (inputs(73)) and not (inputs(27));
    layer0_outputs(6473) <= inputs(152);
    layer0_outputs(6474) <= inputs(84);
    layer0_outputs(6475) <= (inputs(228)) or (inputs(67));
    layer0_outputs(6476) <= not((inputs(156)) or (inputs(78)));
    layer0_outputs(6477) <= not((inputs(233)) or (inputs(226)));
    layer0_outputs(6478) <= not(inputs(228));
    layer0_outputs(6479) <= (inputs(251)) xor (inputs(244));
    layer0_outputs(6480) <= not((inputs(134)) xor (inputs(209)));
    layer0_outputs(6481) <= not((inputs(105)) xor (inputs(108)));
    layer0_outputs(6482) <= (inputs(71)) and not (inputs(229));
    layer0_outputs(6483) <= inputs(230);
    layer0_outputs(6484) <= not(inputs(184)) or (inputs(207));
    layer0_outputs(6485) <= not((inputs(27)) or (inputs(70)));
    layer0_outputs(6486) <= not(inputs(135));
    layer0_outputs(6487) <= '1';
    layer0_outputs(6488) <= (inputs(16)) or (inputs(181));
    layer0_outputs(6489) <= inputs(101);
    layer0_outputs(6490) <= not(inputs(163));
    layer0_outputs(6491) <= not((inputs(225)) or (inputs(170)));
    layer0_outputs(6492) <= (inputs(225)) xor (inputs(139));
    layer0_outputs(6493) <= not((inputs(145)) and (inputs(226)));
    layer0_outputs(6494) <= (inputs(106)) xor (inputs(252));
    layer0_outputs(6495) <= (inputs(210)) or (inputs(68));
    layer0_outputs(6496) <= not(inputs(39));
    layer0_outputs(6497) <= not(inputs(150)) or (inputs(78));
    layer0_outputs(6498) <= inputs(151);
    layer0_outputs(6499) <= inputs(199);
    layer0_outputs(6500) <= not(inputs(94));
    layer0_outputs(6501) <= not((inputs(103)) or (inputs(178)));
    layer0_outputs(6502) <= not(inputs(74));
    layer0_outputs(6503) <= (inputs(133)) xor (inputs(16));
    layer0_outputs(6504) <= (inputs(245)) xor (inputs(24));
    layer0_outputs(6505) <= (inputs(106)) and not (inputs(237));
    layer0_outputs(6506) <= not((inputs(34)) xor (inputs(227)));
    layer0_outputs(6507) <= not(inputs(135));
    layer0_outputs(6508) <= '1';
    layer0_outputs(6509) <= (inputs(37)) and not (inputs(237));
    layer0_outputs(6510) <= (inputs(67)) or (inputs(122));
    layer0_outputs(6511) <= not(inputs(71)) or (inputs(140));
    layer0_outputs(6512) <= (inputs(103)) and not (inputs(205));
    layer0_outputs(6513) <= not((inputs(182)) or (inputs(238)));
    layer0_outputs(6514) <= not((inputs(194)) and (inputs(15)));
    layer0_outputs(6515) <= not(inputs(68));
    layer0_outputs(6516) <= not(inputs(183)) or (inputs(35));
    layer0_outputs(6517) <= inputs(166);
    layer0_outputs(6518) <= not(inputs(63)) or (inputs(160));
    layer0_outputs(6519) <= not((inputs(76)) xor (inputs(209)));
    layer0_outputs(6520) <= not((inputs(33)) and (inputs(220)));
    layer0_outputs(6521) <= not(inputs(62)) or (inputs(77));
    layer0_outputs(6522) <= (inputs(103)) and not (inputs(209));
    layer0_outputs(6523) <= not(inputs(133)) or (inputs(4));
    layer0_outputs(6524) <= (inputs(110)) and not (inputs(16));
    layer0_outputs(6525) <= (inputs(79)) and not (inputs(110));
    layer0_outputs(6526) <= (inputs(70)) and (inputs(219));
    layer0_outputs(6527) <= not((inputs(62)) or (inputs(183)));
    layer0_outputs(6528) <= not(inputs(57));
    layer0_outputs(6529) <= not((inputs(194)) xor (inputs(171)));
    layer0_outputs(6530) <= not((inputs(253)) or (inputs(65)));
    layer0_outputs(6531) <= inputs(110);
    layer0_outputs(6532) <= '0';
    layer0_outputs(6533) <= inputs(134);
    layer0_outputs(6534) <= not(inputs(156)) or (inputs(99));
    layer0_outputs(6535) <= not((inputs(172)) and (inputs(2)));
    layer0_outputs(6536) <= inputs(50);
    layer0_outputs(6537) <= '0';
    layer0_outputs(6538) <= (inputs(124)) xor (inputs(246));
    layer0_outputs(6539) <= (inputs(165)) or (inputs(164));
    layer0_outputs(6540) <= (inputs(239)) and not (inputs(0));
    layer0_outputs(6541) <= not(inputs(83));
    layer0_outputs(6542) <= inputs(56);
    layer0_outputs(6543) <= not(inputs(216)) or (inputs(142));
    layer0_outputs(6544) <= (inputs(151)) and not (inputs(77));
    layer0_outputs(6545) <= (inputs(218)) and not (inputs(177));
    layer0_outputs(6546) <= (inputs(58)) and not (inputs(24));
    layer0_outputs(6547) <= inputs(119);
    layer0_outputs(6548) <= (inputs(83)) or (inputs(50));
    layer0_outputs(6549) <= (inputs(103)) and not (inputs(64));
    layer0_outputs(6550) <= not((inputs(147)) or (inputs(37)));
    layer0_outputs(6551) <= not(inputs(152));
    layer0_outputs(6552) <= (inputs(161)) and not (inputs(1));
    layer0_outputs(6553) <= not(inputs(155)) or (inputs(15));
    layer0_outputs(6554) <= not((inputs(108)) xor (inputs(78)));
    layer0_outputs(6555) <= (inputs(12)) and (inputs(0));
    layer0_outputs(6556) <= (inputs(238)) and (inputs(171));
    layer0_outputs(6557) <= not(inputs(120));
    layer0_outputs(6558) <= (inputs(205)) or (inputs(174));
    layer0_outputs(6559) <= not((inputs(21)) xor (inputs(23)));
    layer0_outputs(6560) <= not((inputs(150)) or (inputs(83)));
    layer0_outputs(6561) <= not(inputs(141));
    layer0_outputs(6562) <= inputs(184);
    layer0_outputs(6563) <= (inputs(153)) and not (inputs(253));
    layer0_outputs(6564) <= not(inputs(7));
    layer0_outputs(6565) <= (inputs(136)) and not (inputs(19));
    layer0_outputs(6566) <= inputs(176);
    layer0_outputs(6567) <= not((inputs(144)) or (inputs(12)));
    layer0_outputs(6568) <= (inputs(14)) xor (inputs(8));
    layer0_outputs(6569) <= (inputs(107)) or (inputs(228));
    layer0_outputs(6570) <= inputs(21);
    layer0_outputs(6571) <= not(inputs(123)) or (inputs(137));
    layer0_outputs(6572) <= (inputs(91)) or (inputs(222));
    layer0_outputs(6573) <= not((inputs(42)) or (inputs(142)));
    layer0_outputs(6574) <= not((inputs(246)) and (inputs(60)));
    layer0_outputs(6575) <= not((inputs(3)) or (inputs(182)));
    layer0_outputs(6576) <= (inputs(176)) xor (inputs(47));
    layer0_outputs(6577) <= (inputs(185)) or (inputs(25));
    layer0_outputs(6578) <= not(inputs(202));
    layer0_outputs(6579) <= not(inputs(164));
    layer0_outputs(6580) <= (inputs(163)) or (inputs(194));
    layer0_outputs(6581) <= (inputs(185)) and not (inputs(52));
    layer0_outputs(6582) <= (inputs(193)) xor (inputs(47));
    layer0_outputs(6583) <= not((inputs(34)) or (inputs(105)));
    layer0_outputs(6584) <= (inputs(51)) and (inputs(77));
    layer0_outputs(6585) <= (inputs(215)) xor (inputs(190));
    layer0_outputs(6586) <= not(inputs(125));
    layer0_outputs(6587) <= (inputs(231)) or (inputs(54));
    layer0_outputs(6588) <= (inputs(167)) and not (inputs(222));
    layer0_outputs(6589) <= (inputs(78)) or (inputs(167));
    layer0_outputs(6590) <= not((inputs(202)) or (inputs(181)));
    layer0_outputs(6591) <= (inputs(28)) and not (inputs(9));
    layer0_outputs(6592) <= (inputs(90)) and not (inputs(23));
    layer0_outputs(6593) <= (inputs(180)) and not (inputs(67));
    layer0_outputs(6594) <= not((inputs(147)) or (inputs(42)));
    layer0_outputs(6595) <= not((inputs(82)) or (inputs(174)));
    layer0_outputs(6596) <= not(inputs(18)) or (inputs(161));
    layer0_outputs(6597) <= not((inputs(134)) or (inputs(209)));
    layer0_outputs(6598) <= not(inputs(213)) or (inputs(51));
    layer0_outputs(6599) <= (inputs(163)) xor (inputs(235));
    layer0_outputs(6600) <= (inputs(162)) or (inputs(163));
    layer0_outputs(6601) <= (inputs(22)) and not (inputs(175));
    layer0_outputs(6602) <= not(inputs(137)) or (inputs(166));
    layer0_outputs(6603) <= (inputs(74)) xor (inputs(184));
    layer0_outputs(6604) <= (inputs(126)) and not (inputs(89));
    layer0_outputs(6605) <= not(inputs(140)) or (inputs(234));
    layer0_outputs(6606) <= not(inputs(174));
    layer0_outputs(6607) <= (inputs(172)) xor (inputs(92));
    layer0_outputs(6608) <= not((inputs(169)) or (inputs(179)));
    layer0_outputs(6609) <= (inputs(192)) xor (inputs(116));
    layer0_outputs(6610) <= not(inputs(91)) or (inputs(221));
    layer0_outputs(6611) <= (inputs(241)) xor (inputs(217));
    layer0_outputs(6612) <= (inputs(189)) or (inputs(30));
    layer0_outputs(6613) <= (inputs(233)) and not (inputs(245));
    layer0_outputs(6614) <= not(inputs(51)) or (inputs(51));
    layer0_outputs(6615) <= inputs(252);
    layer0_outputs(6616) <= '1';
    layer0_outputs(6617) <= (inputs(119)) and not (inputs(241));
    layer0_outputs(6618) <= (inputs(28)) xor (inputs(46));
    layer0_outputs(6619) <= (inputs(116)) or (inputs(61));
    layer0_outputs(6620) <= not(inputs(130)) or (inputs(14));
    layer0_outputs(6621) <= (inputs(96)) xor (inputs(58));
    layer0_outputs(6622) <= inputs(181);
    layer0_outputs(6623) <= (inputs(88)) and not (inputs(179));
    layer0_outputs(6624) <= not((inputs(82)) xor (inputs(71)));
    layer0_outputs(6625) <= not(inputs(78));
    layer0_outputs(6626) <= not(inputs(85));
    layer0_outputs(6627) <= (inputs(248)) or (inputs(41));
    layer0_outputs(6628) <= not((inputs(0)) and (inputs(214)));
    layer0_outputs(6629) <= not(inputs(125)) or (inputs(220));
    layer0_outputs(6630) <= not(inputs(96)) or (inputs(208));
    layer0_outputs(6631) <= (inputs(76)) and not (inputs(15));
    layer0_outputs(6632) <= not(inputs(216));
    layer0_outputs(6633) <= not(inputs(165));
    layer0_outputs(6634) <= not(inputs(128));
    layer0_outputs(6635) <= (inputs(195)) and not (inputs(192));
    layer0_outputs(6636) <= inputs(229);
    layer0_outputs(6637) <= not((inputs(93)) xor (inputs(245)));
    layer0_outputs(6638) <= (inputs(26)) or (inputs(210));
    layer0_outputs(6639) <= (inputs(2)) xor (inputs(189));
    layer0_outputs(6640) <= (inputs(217)) xor (inputs(101));
    layer0_outputs(6641) <= (inputs(62)) and not (inputs(22));
    layer0_outputs(6642) <= inputs(85);
    layer0_outputs(6643) <= not(inputs(0));
    layer0_outputs(6644) <= (inputs(158)) and (inputs(125));
    layer0_outputs(6645) <= (inputs(142)) and not (inputs(250));
    layer0_outputs(6646) <= (inputs(190)) or (inputs(6));
    layer0_outputs(6647) <= not(inputs(90));
    layer0_outputs(6648) <= not((inputs(211)) and (inputs(114)));
    layer0_outputs(6649) <= not((inputs(157)) xor (inputs(196)));
    layer0_outputs(6650) <= (inputs(192)) xor (inputs(142));
    layer0_outputs(6651) <= not((inputs(147)) or (inputs(9)));
    layer0_outputs(6652) <= (inputs(243)) and not (inputs(219));
    layer0_outputs(6653) <= (inputs(141)) and not (inputs(217));
    layer0_outputs(6654) <= (inputs(91)) xor (inputs(92));
    layer0_outputs(6655) <= not((inputs(217)) and (inputs(78)));
    layer0_outputs(6656) <= not((inputs(6)) xor (inputs(133)));
    layer0_outputs(6657) <= not(inputs(187));
    layer0_outputs(6658) <= not(inputs(114));
    layer0_outputs(6659) <= inputs(49);
    layer0_outputs(6660) <= (inputs(195)) and not (inputs(239));
    layer0_outputs(6661) <= inputs(3);
    layer0_outputs(6662) <= not(inputs(122));
    layer0_outputs(6663) <= inputs(166);
    layer0_outputs(6664) <= not((inputs(89)) or (inputs(126)));
    layer0_outputs(6665) <= not((inputs(34)) or (inputs(17)));
    layer0_outputs(6666) <= not((inputs(142)) or (inputs(12)));
    layer0_outputs(6667) <= (inputs(1)) or (inputs(168));
    layer0_outputs(6668) <= '0';
    layer0_outputs(6669) <= '0';
    layer0_outputs(6670) <= (inputs(76)) or (inputs(124));
    layer0_outputs(6671) <= (inputs(149)) xor (inputs(19));
    layer0_outputs(6672) <= not(inputs(62));
    layer0_outputs(6673) <= '0';
    layer0_outputs(6674) <= (inputs(237)) and not (inputs(95));
    layer0_outputs(6675) <= not(inputs(182));
    layer0_outputs(6676) <= (inputs(55)) xor (inputs(105));
    layer0_outputs(6677) <= not((inputs(237)) or (inputs(198)));
    layer0_outputs(6678) <= not(inputs(209));
    layer0_outputs(6679) <= (inputs(191)) or (inputs(27));
    layer0_outputs(6680) <= not(inputs(183)) or (inputs(226));
    layer0_outputs(6681) <= not(inputs(31)) or (inputs(190));
    layer0_outputs(6682) <= inputs(174);
    layer0_outputs(6683) <= not(inputs(99)) or (inputs(93));
    layer0_outputs(6684) <= (inputs(122)) and not (inputs(7));
    layer0_outputs(6685) <= (inputs(63)) and not (inputs(29));
    layer0_outputs(6686) <= inputs(118);
    layer0_outputs(6687) <= inputs(114);
    layer0_outputs(6688) <= not(inputs(115)) or (inputs(254));
    layer0_outputs(6689) <= not((inputs(156)) and (inputs(108)));
    layer0_outputs(6690) <= not(inputs(72));
    layer0_outputs(6691) <= (inputs(156)) or (inputs(197));
    layer0_outputs(6692) <= (inputs(254)) and not (inputs(209));
    layer0_outputs(6693) <= not((inputs(6)) or (inputs(93)));
    layer0_outputs(6694) <= (inputs(206)) xor (inputs(139));
    layer0_outputs(6695) <= not(inputs(181));
    layer0_outputs(6696) <= not(inputs(134));
    layer0_outputs(6697) <= (inputs(203)) or (inputs(33));
    layer0_outputs(6698) <= not((inputs(66)) and (inputs(189)));
    layer0_outputs(6699) <= '1';
    layer0_outputs(6700) <= (inputs(200)) xor (inputs(70));
    layer0_outputs(6701) <= (inputs(70)) and not (inputs(242));
    layer0_outputs(6702) <= not(inputs(140)) or (inputs(239));
    layer0_outputs(6703) <= not(inputs(153)) or (inputs(56));
    layer0_outputs(6704) <= not(inputs(154));
    layer0_outputs(6705) <= (inputs(13)) xor (inputs(174));
    layer0_outputs(6706) <= (inputs(187)) or (inputs(41));
    layer0_outputs(6707) <= inputs(9);
    layer0_outputs(6708) <= not((inputs(214)) or (inputs(248)));
    layer0_outputs(6709) <= not(inputs(170)) or (inputs(205));
    layer0_outputs(6710) <= (inputs(10)) and not (inputs(34));
    layer0_outputs(6711) <= '0';
    layer0_outputs(6712) <= (inputs(192)) and (inputs(127));
    layer0_outputs(6713) <= not(inputs(232));
    layer0_outputs(6714) <= (inputs(119)) xor (inputs(76));
    layer0_outputs(6715) <= not((inputs(42)) or (inputs(247)));
    layer0_outputs(6716) <= not((inputs(234)) or (inputs(19)));
    layer0_outputs(6717) <= not(inputs(178));
    layer0_outputs(6718) <= (inputs(198)) xor (inputs(82));
    layer0_outputs(6719) <= not(inputs(15));
    layer0_outputs(6720) <= not((inputs(78)) or (inputs(77)));
    layer0_outputs(6721) <= (inputs(242)) and not (inputs(113));
    layer0_outputs(6722) <= inputs(183);
    layer0_outputs(6723) <= not((inputs(81)) or (inputs(185)));
    layer0_outputs(6724) <= inputs(120);
    layer0_outputs(6725) <= (inputs(111)) or (inputs(67));
    layer0_outputs(6726) <= not((inputs(32)) or (inputs(228)));
    layer0_outputs(6727) <= not(inputs(26));
    layer0_outputs(6728) <= not(inputs(116));
    layer0_outputs(6729) <= (inputs(120)) or (inputs(11));
    layer0_outputs(6730) <= (inputs(186)) and not (inputs(128));
    layer0_outputs(6731) <= (inputs(146)) and not (inputs(174));
    layer0_outputs(6732) <= not((inputs(68)) or (inputs(40)));
    layer0_outputs(6733) <= not((inputs(211)) xor (inputs(247)));
    layer0_outputs(6734) <= not((inputs(39)) or (inputs(10)));
    layer0_outputs(6735) <= not(inputs(252)) or (inputs(209));
    layer0_outputs(6736) <= not(inputs(120)) or (inputs(14));
    layer0_outputs(6737) <= (inputs(124)) xor (inputs(182));
    layer0_outputs(6738) <= (inputs(125)) xor (inputs(191));
    layer0_outputs(6739) <= not(inputs(106));
    layer0_outputs(6740) <= (inputs(151)) and not (inputs(137));
    layer0_outputs(6741) <= (inputs(173)) and not (inputs(44));
    layer0_outputs(6742) <= not(inputs(155)) or (inputs(100));
    layer0_outputs(6743) <= not((inputs(62)) or (inputs(219)));
    layer0_outputs(6744) <= inputs(229);
    layer0_outputs(6745) <= (inputs(95)) and not (inputs(38));
    layer0_outputs(6746) <= (inputs(163)) xor (inputs(189));
    layer0_outputs(6747) <= (inputs(165)) and not (inputs(98));
    layer0_outputs(6748) <= not(inputs(151)) or (inputs(148));
    layer0_outputs(6749) <= (inputs(171)) or (inputs(185));
    layer0_outputs(6750) <= not((inputs(82)) or (inputs(165)));
    layer0_outputs(6751) <= not(inputs(103));
    layer0_outputs(6752) <= not((inputs(21)) or (inputs(171)));
    layer0_outputs(6753) <= not((inputs(234)) xor (inputs(25)));
    layer0_outputs(6754) <= (inputs(137)) and not (inputs(225));
    layer0_outputs(6755) <= '1';
    layer0_outputs(6756) <= not(inputs(22));
    layer0_outputs(6757) <= inputs(137);
    layer0_outputs(6758) <= not((inputs(191)) or (inputs(10)));
    layer0_outputs(6759) <= not((inputs(38)) xor (inputs(231)));
    layer0_outputs(6760) <= not(inputs(19)) or (inputs(20));
    layer0_outputs(6761) <= not(inputs(93));
    layer0_outputs(6762) <= not(inputs(43)) or (inputs(66));
    layer0_outputs(6763) <= not(inputs(38)) or (inputs(31));
    layer0_outputs(6764) <= (inputs(68)) and not (inputs(14));
    layer0_outputs(6765) <= not(inputs(43));
    layer0_outputs(6766) <= (inputs(123)) and not (inputs(15));
    layer0_outputs(6767) <= inputs(40);
    layer0_outputs(6768) <= (inputs(239)) xor (inputs(219));
    layer0_outputs(6769) <= '0';
    layer0_outputs(6770) <= not(inputs(243)) or (inputs(179));
    layer0_outputs(6771) <= (inputs(63)) xor (inputs(24));
    layer0_outputs(6772) <= inputs(244);
    layer0_outputs(6773) <= not((inputs(143)) xor (inputs(34)));
    layer0_outputs(6774) <= not((inputs(80)) or (inputs(16)));
    layer0_outputs(6775) <= inputs(132);
    layer0_outputs(6776) <= '1';
    layer0_outputs(6777) <= (inputs(79)) or (inputs(88));
    layer0_outputs(6778) <= not((inputs(32)) and (inputs(158)));
    layer0_outputs(6779) <= (inputs(10)) and (inputs(17));
    layer0_outputs(6780) <= not((inputs(66)) or (inputs(199)));
    layer0_outputs(6781) <= not((inputs(47)) xor (inputs(22)));
    layer0_outputs(6782) <= (inputs(164)) xor (inputs(247));
    layer0_outputs(6783) <= (inputs(201)) and not (inputs(85));
    layer0_outputs(6784) <= not(inputs(177));
    layer0_outputs(6785) <= (inputs(209)) or (inputs(75));
    layer0_outputs(6786) <= (inputs(96)) and (inputs(144));
    layer0_outputs(6787) <= not((inputs(70)) xor (inputs(34)));
    layer0_outputs(6788) <= inputs(3);
    layer0_outputs(6789) <= inputs(47);
    layer0_outputs(6790) <= not(inputs(0)) or (inputs(63));
    layer0_outputs(6791) <= not((inputs(156)) and (inputs(59)));
    layer0_outputs(6792) <= not((inputs(6)) xor (inputs(179)));
    layer0_outputs(6793) <= (inputs(125)) and not (inputs(37));
    layer0_outputs(6794) <= not(inputs(198)) or (inputs(13));
    layer0_outputs(6795) <= (inputs(139)) and (inputs(169));
    layer0_outputs(6796) <= '0';
    layer0_outputs(6797) <= inputs(70);
    layer0_outputs(6798) <= not((inputs(178)) and (inputs(232)));
    layer0_outputs(6799) <= (inputs(169)) xor (inputs(184));
    layer0_outputs(6800) <= not(inputs(43));
    layer0_outputs(6801) <= (inputs(178)) or (inputs(179));
    layer0_outputs(6802) <= inputs(150);
    layer0_outputs(6803) <= (inputs(134)) xor (inputs(2));
    layer0_outputs(6804) <= not(inputs(162));
    layer0_outputs(6805) <= (inputs(46)) or (inputs(159));
    layer0_outputs(6806) <= (inputs(57)) and not (inputs(131));
    layer0_outputs(6807) <= not(inputs(68));
    layer0_outputs(6808) <= not((inputs(202)) or (inputs(244)));
    layer0_outputs(6809) <= not(inputs(103)) or (inputs(66));
    layer0_outputs(6810) <= inputs(96);
    layer0_outputs(6811) <= not(inputs(150)) or (inputs(167));
    layer0_outputs(6812) <= not(inputs(2));
    layer0_outputs(6813) <= (inputs(120)) and not (inputs(172));
    layer0_outputs(6814) <= inputs(148);
    layer0_outputs(6815) <= not(inputs(42));
    layer0_outputs(6816) <= (inputs(129)) and (inputs(93));
    layer0_outputs(6817) <= '0';
    layer0_outputs(6818) <= not((inputs(243)) or (inputs(160)));
    layer0_outputs(6819) <= not((inputs(22)) and (inputs(220)));
    layer0_outputs(6820) <= not((inputs(145)) xor (inputs(148)));
    layer0_outputs(6821) <= not(inputs(178));
    layer0_outputs(6822) <= (inputs(233)) and not (inputs(45));
    layer0_outputs(6823) <= not((inputs(227)) and (inputs(141)));
    layer0_outputs(6824) <= (inputs(159)) or (inputs(197));
    layer0_outputs(6825) <= (inputs(200)) and not (inputs(239));
    layer0_outputs(6826) <= not((inputs(159)) xor (inputs(6)));
    layer0_outputs(6827) <= (inputs(101)) and not (inputs(172));
    layer0_outputs(6828) <= '1';
    layer0_outputs(6829) <= not(inputs(94)) or (inputs(97));
    layer0_outputs(6830) <= not((inputs(228)) or (inputs(147)));
    layer0_outputs(6831) <= not((inputs(40)) xor (inputs(238)));
    layer0_outputs(6832) <= not((inputs(196)) or (inputs(8)));
    layer0_outputs(6833) <= not(inputs(79)) or (inputs(82));
    layer0_outputs(6834) <= (inputs(31)) and not (inputs(239));
    layer0_outputs(6835) <= not((inputs(50)) or (inputs(133)));
    layer0_outputs(6836) <= (inputs(133)) xor (inputs(78));
    layer0_outputs(6837) <= not((inputs(168)) or (inputs(118)));
    layer0_outputs(6838) <= (inputs(224)) and not (inputs(237));
    layer0_outputs(6839) <= not(inputs(112));
    layer0_outputs(6840) <= inputs(39);
    layer0_outputs(6841) <= not((inputs(198)) and (inputs(139)));
    layer0_outputs(6842) <= '0';
    layer0_outputs(6843) <= (inputs(52)) xor (inputs(190));
    layer0_outputs(6844) <= not(inputs(152)) or (inputs(203));
    layer0_outputs(6845) <= not(inputs(220)) or (inputs(43));
    layer0_outputs(6846) <= not((inputs(147)) or (inputs(160)));
    layer0_outputs(6847) <= (inputs(176)) xor (inputs(172));
    layer0_outputs(6848) <= not(inputs(10)) or (inputs(94));
    layer0_outputs(6849) <= not(inputs(175)) or (inputs(194));
    layer0_outputs(6850) <= not(inputs(185)) or (inputs(251));
    layer0_outputs(6851) <= not(inputs(59)) or (inputs(207));
    layer0_outputs(6852) <= (inputs(200)) and not (inputs(33));
    layer0_outputs(6853) <= not(inputs(32));
    layer0_outputs(6854) <= inputs(16);
    layer0_outputs(6855) <= not(inputs(74));
    layer0_outputs(6856) <= '1';
    layer0_outputs(6857) <= (inputs(99)) and (inputs(128));
    layer0_outputs(6858) <= (inputs(128)) xor (inputs(191));
    layer0_outputs(6859) <= not((inputs(117)) xor (inputs(244)));
    layer0_outputs(6860) <= not(inputs(94)) or (inputs(238));
    layer0_outputs(6861) <= (inputs(171)) or (inputs(180));
    layer0_outputs(6862) <= inputs(200);
    layer0_outputs(6863) <= not(inputs(79)) or (inputs(115));
    layer0_outputs(6864) <= (inputs(147)) and not (inputs(240));
    layer0_outputs(6865) <= not((inputs(154)) or (inputs(19)));
    layer0_outputs(6866) <= not((inputs(219)) and (inputs(172)));
    layer0_outputs(6867) <= (inputs(199)) and not (inputs(93));
    layer0_outputs(6868) <= not((inputs(223)) or (inputs(194)));
    layer0_outputs(6869) <= not(inputs(131)) or (inputs(192));
    layer0_outputs(6870) <= (inputs(223)) and (inputs(69));
    layer0_outputs(6871) <= (inputs(108)) and not (inputs(19));
    layer0_outputs(6872) <= not((inputs(48)) or (inputs(117)));
    layer0_outputs(6873) <= (inputs(139)) or (inputs(30));
    layer0_outputs(6874) <= not((inputs(4)) and (inputs(16)));
    layer0_outputs(6875) <= not((inputs(192)) or (inputs(41)));
    layer0_outputs(6876) <= '1';
    layer0_outputs(6877) <= not(inputs(70));
    layer0_outputs(6878) <= not((inputs(140)) and (inputs(77)));
    layer0_outputs(6879) <= inputs(182);
    layer0_outputs(6880) <= not(inputs(38));
    layer0_outputs(6881) <= not(inputs(103));
    layer0_outputs(6882) <= not((inputs(20)) and (inputs(108)));
    layer0_outputs(6883) <= inputs(118);
    layer0_outputs(6884) <= not((inputs(241)) or (inputs(126)));
    layer0_outputs(6885) <= not((inputs(159)) and (inputs(225)));
    layer0_outputs(6886) <= not(inputs(155)) or (inputs(43));
    layer0_outputs(6887) <= not((inputs(128)) xor (inputs(206)));
    layer0_outputs(6888) <= (inputs(227)) or (inputs(88));
    layer0_outputs(6889) <= (inputs(116)) or (inputs(219));
    layer0_outputs(6890) <= '1';
    layer0_outputs(6891) <= (inputs(62)) xor (inputs(227));
    layer0_outputs(6892) <= (inputs(116)) and not (inputs(191));
    layer0_outputs(6893) <= inputs(140);
    layer0_outputs(6894) <= not((inputs(213)) and (inputs(42)));
    layer0_outputs(6895) <= (inputs(125)) or (inputs(185));
    layer0_outputs(6896) <= not((inputs(18)) and (inputs(112)));
    layer0_outputs(6897) <= (inputs(1)) and (inputs(221));
    layer0_outputs(6898) <= not(inputs(81));
    layer0_outputs(6899) <= not(inputs(43)) or (inputs(62));
    layer0_outputs(6900) <= inputs(113);
    layer0_outputs(6901) <= not(inputs(178)) or (inputs(212));
    layer0_outputs(6902) <= inputs(54);
    layer0_outputs(6903) <= '0';
    layer0_outputs(6904) <= not(inputs(239)) or (inputs(77));
    layer0_outputs(6905) <= not((inputs(34)) xor (inputs(206)));
    layer0_outputs(6906) <= (inputs(64)) and not (inputs(89));
    layer0_outputs(6907) <= not((inputs(140)) or (inputs(35)));
    layer0_outputs(6908) <= not((inputs(15)) xor (inputs(56)));
    layer0_outputs(6909) <= not(inputs(231));
    layer0_outputs(6910) <= '0';
    layer0_outputs(6911) <= not(inputs(199));
    layer0_outputs(6912) <= inputs(76);
    layer0_outputs(6913) <= not((inputs(255)) or (inputs(78)));
    layer0_outputs(6914) <= (inputs(45)) and not (inputs(40));
    layer0_outputs(6915) <= not(inputs(34));
    layer0_outputs(6916) <= not(inputs(200)) or (inputs(214));
    layer0_outputs(6917) <= not((inputs(33)) or (inputs(183)));
    layer0_outputs(6918) <= not(inputs(60));
    layer0_outputs(6919) <= (inputs(81)) or (inputs(211));
    layer0_outputs(6920) <= '1';
    layer0_outputs(6921) <= (inputs(211)) and not (inputs(101));
    layer0_outputs(6922) <= (inputs(36)) xor (inputs(243));
    layer0_outputs(6923) <= not((inputs(7)) and (inputs(123)));
    layer0_outputs(6924) <= '0';
    layer0_outputs(6925) <= inputs(73);
    layer0_outputs(6926) <= inputs(57);
    layer0_outputs(6927) <= (inputs(234)) and not (inputs(190));
    layer0_outputs(6928) <= (inputs(153)) or (inputs(249));
    layer0_outputs(6929) <= not((inputs(121)) xor (inputs(162)));
    layer0_outputs(6930) <= not(inputs(184));
    layer0_outputs(6931) <= not(inputs(158));
    layer0_outputs(6932) <= not((inputs(230)) or (inputs(136)));
    layer0_outputs(6933) <= not(inputs(117));
    layer0_outputs(6934) <= not((inputs(211)) xor (inputs(163)));
    layer0_outputs(6935) <= not(inputs(194)) or (inputs(246));
    layer0_outputs(6936) <= not(inputs(91));
    layer0_outputs(6937) <= inputs(85);
    layer0_outputs(6938) <= (inputs(15)) or (inputs(179));
    layer0_outputs(6939) <= (inputs(184)) or (inputs(234));
    layer0_outputs(6940) <= (inputs(200)) and not (inputs(189));
    layer0_outputs(6941) <= not((inputs(187)) xor (inputs(180)));
    layer0_outputs(6942) <= (inputs(57)) or (inputs(204));
    layer0_outputs(6943) <= not(inputs(164)) or (inputs(176));
    layer0_outputs(6944) <= (inputs(239)) xor (inputs(52));
    layer0_outputs(6945) <= not((inputs(57)) xor (inputs(186)));
    layer0_outputs(6946) <= '0';
    layer0_outputs(6947) <= (inputs(127)) xor (inputs(151));
    layer0_outputs(6948) <= not(inputs(232)) or (inputs(50));
    layer0_outputs(6949) <= (inputs(175)) and not (inputs(178));
    layer0_outputs(6950) <= (inputs(108)) or (inputs(230));
    layer0_outputs(6951) <= (inputs(85)) and not (inputs(184));
    layer0_outputs(6952) <= not((inputs(166)) xor (inputs(25)));
    layer0_outputs(6953) <= (inputs(133)) and not (inputs(109));
    layer0_outputs(6954) <= not(inputs(101));
    layer0_outputs(6955) <= (inputs(102)) or (inputs(83));
    layer0_outputs(6956) <= (inputs(240)) or (inputs(4));
    layer0_outputs(6957) <= not(inputs(36));
    layer0_outputs(6958) <= not((inputs(33)) xor (inputs(141)));
    layer0_outputs(6959) <= not(inputs(132));
    layer0_outputs(6960) <= not((inputs(60)) and (inputs(94)));
    layer0_outputs(6961) <= (inputs(79)) xor (inputs(52));
    layer0_outputs(6962) <= not((inputs(99)) and (inputs(97)));
    layer0_outputs(6963) <= (inputs(22)) or (inputs(164));
    layer0_outputs(6964) <= not(inputs(209));
    layer0_outputs(6965) <= not(inputs(255));
    layer0_outputs(6966) <= inputs(157);
    layer0_outputs(6967) <= not((inputs(229)) or (inputs(227)));
    layer0_outputs(6968) <= not((inputs(142)) xor (inputs(100)));
    layer0_outputs(6969) <= not(inputs(189)) or (inputs(29));
    layer0_outputs(6970) <= not((inputs(82)) xor (inputs(208)));
    layer0_outputs(6971) <= not((inputs(219)) or (inputs(1)));
    layer0_outputs(6972) <= inputs(217);
    layer0_outputs(6973) <= not(inputs(80));
    layer0_outputs(6974) <= (inputs(16)) and (inputs(190));
    layer0_outputs(6975) <= not(inputs(76));
    layer0_outputs(6976) <= not(inputs(38)) or (inputs(188));
    layer0_outputs(6977) <= inputs(246);
    layer0_outputs(6978) <= (inputs(59)) xor (inputs(16));
    layer0_outputs(6979) <= not(inputs(224));
    layer0_outputs(6980) <= not(inputs(149));
    layer0_outputs(6981) <= not((inputs(196)) xor (inputs(246)));
    layer0_outputs(6982) <= (inputs(184)) or (inputs(207));
    layer0_outputs(6983) <= '1';
    layer0_outputs(6984) <= (inputs(132)) or (inputs(200));
    layer0_outputs(6985) <= inputs(50);
    layer0_outputs(6986) <= (inputs(240)) and not (inputs(185));
    layer0_outputs(6987) <= not((inputs(42)) and (inputs(216)));
    layer0_outputs(6988) <= not(inputs(232));
    layer0_outputs(6989) <= (inputs(41)) or (inputs(47));
    layer0_outputs(6990) <= (inputs(140)) and not (inputs(101));
    layer0_outputs(6991) <= not((inputs(68)) xor (inputs(12)));
    layer0_outputs(6992) <= not((inputs(9)) xor (inputs(92)));
    layer0_outputs(6993) <= '0';
    layer0_outputs(6994) <= not(inputs(95)) or (inputs(28));
    layer0_outputs(6995) <= (inputs(31)) xor (inputs(137));
    layer0_outputs(6996) <= (inputs(223)) or (inputs(212));
    layer0_outputs(6997) <= not((inputs(99)) xor (inputs(86)));
    layer0_outputs(6998) <= not(inputs(88));
    layer0_outputs(6999) <= not((inputs(200)) or (inputs(95)));
    layer0_outputs(7000) <= (inputs(97)) and (inputs(184));
    layer0_outputs(7001) <= not(inputs(109));
    layer0_outputs(7002) <= not(inputs(87)) or (inputs(189));
    layer0_outputs(7003) <= (inputs(135)) and not (inputs(63));
    layer0_outputs(7004) <= (inputs(195)) xor (inputs(195));
    layer0_outputs(7005) <= not(inputs(8)) or (inputs(42));
    layer0_outputs(7006) <= (inputs(134)) and not (inputs(238));
    layer0_outputs(7007) <= not(inputs(38));
    layer0_outputs(7008) <= (inputs(220)) or (inputs(139));
    layer0_outputs(7009) <= not(inputs(242));
    layer0_outputs(7010) <= (inputs(151)) or (inputs(205));
    layer0_outputs(7011) <= '0';
    layer0_outputs(7012) <= not(inputs(136)) or (inputs(63));
    layer0_outputs(7013) <= (inputs(216)) or (inputs(227));
    layer0_outputs(7014) <= not((inputs(160)) and (inputs(142)));
    layer0_outputs(7015) <= not((inputs(37)) or (inputs(181)));
    layer0_outputs(7016) <= (inputs(20)) xor (inputs(10));
    layer0_outputs(7017) <= (inputs(84)) and not (inputs(128));
    layer0_outputs(7018) <= not(inputs(189)) or (inputs(239));
    layer0_outputs(7019) <= (inputs(149)) and (inputs(99));
    layer0_outputs(7020) <= (inputs(129)) xor (inputs(79));
    layer0_outputs(7021) <= not(inputs(7)) or (inputs(32));
    layer0_outputs(7022) <= not((inputs(62)) xor (inputs(84)));
    layer0_outputs(7023) <= (inputs(233)) xor (inputs(24));
    layer0_outputs(7024) <= (inputs(143)) and (inputs(3));
    layer0_outputs(7025) <= not((inputs(182)) xor (inputs(165)));
    layer0_outputs(7026) <= inputs(220);
    layer0_outputs(7027) <= not(inputs(238));
    layer0_outputs(7028) <= (inputs(141)) and not (inputs(109));
    layer0_outputs(7029) <= not((inputs(50)) or (inputs(50)));
    layer0_outputs(7030) <= (inputs(252)) xor (inputs(194));
    layer0_outputs(7031) <= inputs(188);
    layer0_outputs(7032) <= inputs(10);
    layer0_outputs(7033) <= '1';
    layer0_outputs(7034) <= inputs(246);
    layer0_outputs(7035) <= inputs(58);
    layer0_outputs(7036) <= not(inputs(138)) or (inputs(36));
    layer0_outputs(7037) <= not((inputs(5)) and (inputs(64)));
    layer0_outputs(7038) <= not(inputs(2)) or (inputs(48));
    layer0_outputs(7039) <= not(inputs(218));
    layer0_outputs(7040) <= '0';
    layer0_outputs(7041) <= '1';
    layer0_outputs(7042) <= (inputs(47)) and (inputs(206));
    layer0_outputs(7043) <= not(inputs(120)) or (inputs(174));
    layer0_outputs(7044) <= (inputs(219)) xor (inputs(194));
    layer0_outputs(7045) <= inputs(118);
    layer0_outputs(7046) <= not((inputs(15)) or (inputs(28)));
    layer0_outputs(7047) <= not(inputs(116));
    layer0_outputs(7048) <= not(inputs(119)) or (inputs(2));
    layer0_outputs(7049) <= not((inputs(93)) or (inputs(109)));
    layer0_outputs(7050) <= not(inputs(88));
    layer0_outputs(7051) <= '0';
    layer0_outputs(7052) <= inputs(241);
    layer0_outputs(7053) <= inputs(230);
    layer0_outputs(7054) <= inputs(150);
    layer0_outputs(7055) <= inputs(180);
    layer0_outputs(7056) <= not((inputs(66)) or (inputs(253)));
    layer0_outputs(7057) <= (inputs(217)) and not (inputs(208));
    layer0_outputs(7058) <= (inputs(26)) and not (inputs(193));
    layer0_outputs(7059) <= (inputs(149)) and not (inputs(82));
    layer0_outputs(7060) <= not((inputs(191)) or (inputs(149)));
    layer0_outputs(7061) <= (inputs(122)) or (inputs(64));
    layer0_outputs(7062) <= not(inputs(3)) or (inputs(65));
    layer0_outputs(7063) <= inputs(9);
    layer0_outputs(7064) <= not((inputs(205)) or (inputs(94)));
    layer0_outputs(7065) <= not((inputs(126)) and (inputs(19)));
    layer0_outputs(7066) <= (inputs(180)) and not (inputs(81));
    layer0_outputs(7067) <= (inputs(214)) and not (inputs(7));
    layer0_outputs(7068) <= not((inputs(55)) xor (inputs(43)));
    layer0_outputs(7069) <= not((inputs(11)) or (inputs(170)));
    layer0_outputs(7070) <= inputs(1);
    layer0_outputs(7071) <= not((inputs(254)) and (inputs(35)));
    layer0_outputs(7072) <= inputs(199);
    layer0_outputs(7073) <= not((inputs(110)) or (inputs(225)));
    layer0_outputs(7074) <= not(inputs(59)) or (inputs(228));
    layer0_outputs(7075) <= not((inputs(54)) xor (inputs(3)));
    layer0_outputs(7076) <= not((inputs(58)) xor (inputs(129)));
    layer0_outputs(7077) <= '1';
    layer0_outputs(7078) <= (inputs(102)) xor (inputs(235));
    layer0_outputs(7079) <= (inputs(79)) xor (inputs(144));
    layer0_outputs(7080) <= inputs(93);
    layer0_outputs(7081) <= (inputs(227)) xor (inputs(199));
    layer0_outputs(7082) <= (inputs(115)) and not (inputs(119));
    layer0_outputs(7083) <= '0';
    layer0_outputs(7084) <= (inputs(52)) or (inputs(81));
    layer0_outputs(7085) <= (inputs(166)) xor (inputs(49));
    layer0_outputs(7086) <= (inputs(64)) xor (inputs(213));
    layer0_outputs(7087) <= (inputs(153)) and not (inputs(183));
    layer0_outputs(7088) <= (inputs(17)) and not (inputs(10));
    layer0_outputs(7089) <= not(inputs(52)) or (inputs(133));
    layer0_outputs(7090) <= not((inputs(37)) or (inputs(31)));
    layer0_outputs(7091) <= (inputs(75)) and not (inputs(186));
    layer0_outputs(7092) <= not(inputs(202)) or (inputs(237));
    layer0_outputs(7093) <= not((inputs(171)) or (inputs(10)));
    layer0_outputs(7094) <= (inputs(171)) and (inputs(53));
    layer0_outputs(7095) <= not((inputs(218)) xor (inputs(75)));
    layer0_outputs(7096) <= not((inputs(145)) xor (inputs(70)));
    layer0_outputs(7097) <= '1';
    layer0_outputs(7098) <= not(inputs(93)) or (inputs(35));
    layer0_outputs(7099) <= not((inputs(170)) or (inputs(126)));
    layer0_outputs(7100) <= not(inputs(232));
    layer0_outputs(7101) <= (inputs(189)) and not (inputs(21));
    layer0_outputs(7102) <= not((inputs(191)) xor (inputs(217)));
    layer0_outputs(7103) <= (inputs(144)) and not (inputs(239));
    layer0_outputs(7104) <= '0';
    layer0_outputs(7105) <= (inputs(129)) and not (inputs(112));
    layer0_outputs(7106) <= inputs(235);
    layer0_outputs(7107) <= (inputs(99)) and not (inputs(31));
    layer0_outputs(7108) <= (inputs(25)) and (inputs(65));
    layer0_outputs(7109) <= (inputs(101)) and not (inputs(39));
    layer0_outputs(7110) <= (inputs(29)) or (inputs(131));
    layer0_outputs(7111) <= (inputs(168)) and not (inputs(162));
    layer0_outputs(7112) <= (inputs(114)) or (inputs(76));
    layer0_outputs(7113) <= not(inputs(7));
    layer0_outputs(7114) <= not((inputs(218)) or (inputs(48)));
    layer0_outputs(7115) <= not((inputs(191)) or (inputs(189)));
    layer0_outputs(7116) <= not(inputs(7));
    layer0_outputs(7117) <= inputs(17);
    layer0_outputs(7118) <= (inputs(174)) xor (inputs(235));
    layer0_outputs(7119) <= '1';
    layer0_outputs(7120) <= not(inputs(53)) or (inputs(238));
    layer0_outputs(7121) <= (inputs(91)) or (inputs(146));
    layer0_outputs(7122) <= inputs(14);
    layer0_outputs(7123) <= not(inputs(132)) or (inputs(251));
    layer0_outputs(7124) <= not(inputs(6)) or (inputs(19));
    layer0_outputs(7125) <= not((inputs(230)) or (inputs(143)));
    layer0_outputs(7126) <= (inputs(211)) xor (inputs(125));
    layer0_outputs(7127) <= '1';
    layer0_outputs(7128) <= not(inputs(167));
    layer0_outputs(7129) <= '1';
    layer0_outputs(7130) <= not((inputs(198)) xor (inputs(25)));
    layer0_outputs(7131) <= (inputs(37)) xor (inputs(189));
    layer0_outputs(7132) <= not(inputs(56)) or (inputs(144));
    layer0_outputs(7133) <= inputs(32);
    layer0_outputs(7134) <= not((inputs(117)) xor (inputs(160)));
    layer0_outputs(7135) <= not((inputs(207)) xor (inputs(88)));
    layer0_outputs(7136) <= (inputs(200)) and not (inputs(61));
    layer0_outputs(7137) <= not((inputs(130)) or (inputs(45)));
    layer0_outputs(7138) <= inputs(189);
    layer0_outputs(7139) <= (inputs(197)) or (inputs(60));
    layer0_outputs(7140) <= (inputs(247)) xor (inputs(230));
    layer0_outputs(7141) <= (inputs(125)) or (inputs(108));
    layer0_outputs(7142) <= not((inputs(5)) or (inputs(50)));
    layer0_outputs(7143) <= not(inputs(107));
    layer0_outputs(7144) <= inputs(6);
    layer0_outputs(7145) <= inputs(154);
    layer0_outputs(7146) <= not(inputs(219)) or (inputs(188));
    layer0_outputs(7147) <= (inputs(114)) and not (inputs(97));
    layer0_outputs(7148) <= not(inputs(178));
    layer0_outputs(7149) <= not((inputs(4)) and (inputs(87)));
    layer0_outputs(7150) <= (inputs(254)) xor (inputs(155));
    layer0_outputs(7151) <= not(inputs(209));
    layer0_outputs(7152) <= not(inputs(130));
    layer0_outputs(7153) <= inputs(145);
    layer0_outputs(7154) <= inputs(180);
    layer0_outputs(7155) <= inputs(228);
    layer0_outputs(7156) <= '0';
    layer0_outputs(7157) <= not((inputs(5)) or (inputs(186)));
    layer0_outputs(7158) <= (inputs(225)) xor (inputs(198));
    layer0_outputs(7159) <= not(inputs(44)) or (inputs(159));
    layer0_outputs(7160) <= not(inputs(152)) or (inputs(19));
    layer0_outputs(7161) <= not(inputs(230));
    layer0_outputs(7162) <= '1';
    layer0_outputs(7163) <= not((inputs(228)) or (inputs(2)));
    layer0_outputs(7164) <= not(inputs(22)) or (inputs(8));
    layer0_outputs(7165) <= not((inputs(206)) xor (inputs(9)));
    layer0_outputs(7166) <= inputs(2);
    layer0_outputs(7167) <= (inputs(34)) or (inputs(121));
    layer0_outputs(7168) <= (inputs(72)) and not (inputs(94));
    layer0_outputs(7169) <= (inputs(194)) xor (inputs(150));
    layer0_outputs(7170) <= (inputs(20)) or (inputs(134));
    layer0_outputs(7171) <= not((inputs(133)) or (inputs(45)));
    layer0_outputs(7172) <= not(inputs(54)) or (inputs(150));
    layer0_outputs(7173) <= (inputs(202)) or (inputs(93));
    layer0_outputs(7174) <= not((inputs(235)) or (inputs(93)));
    layer0_outputs(7175) <= (inputs(38)) xor (inputs(96));
    layer0_outputs(7176) <= not(inputs(55)) or (inputs(2));
    layer0_outputs(7177) <= not((inputs(77)) or (inputs(75)));
    layer0_outputs(7178) <= not((inputs(253)) xor (inputs(203)));
    layer0_outputs(7179) <= (inputs(168)) and not (inputs(228));
    layer0_outputs(7180) <= not(inputs(78));
    layer0_outputs(7181) <= not((inputs(52)) xor (inputs(102)));
    layer0_outputs(7182) <= not((inputs(205)) xor (inputs(187)));
    layer0_outputs(7183) <= (inputs(214)) and not (inputs(252));
    layer0_outputs(7184) <= (inputs(95)) xor (inputs(58));
    layer0_outputs(7185) <= '1';
    layer0_outputs(7186) <= not((inputs(164)) and (inputs(175)));
    layer0_outputs(7187) <= not(inputs(138));
    layer0_outputs(7188) <= '0';
    layer0_outputs(7189) <= inputs(129);
    layer0_outputs(7190) <= (inputs(134)) or (inputs(32));
    layer0_outputs(7191) <= (inputs(48)) and not (inputs(110));
    layer0_outputs(7192) <= not(inputs(40)) or (inputs(203));
    layer0_outputs(7193) <= '0';
    layer0_outputs(7194) <= '1';
    layer0_outputs(7195) <= (inputs(244)) and not (inputs(242));
    layer0_outputs(7196) <= not(inputs(25));
    layer0_outputs(7197) <= inputs(130);
    layer0_outputs(7198) <= not(inputs(37));
    layer0_outputs(7199) <= (inputs(177)) xor (inputs(164));
    layer0_outputs(7200) <= inputs(52);
    layer0_outputs(7201) <= not((inputs(141)) and (inputs(66)));
    layer0_outputs(7202) <= (inputs(166)) and not (inputs(60));
    layer0_outputs(7203) <= (inputs(87)) or (inputs(235));
    layer0_outputs(7204) <= not((inputs(177)) or (inputs(128)));
    layer0_outputs(7205) <= not(inputs(69));
    layer0_outputs(7206) <= not((inputs(178)) or (inputs(177)));
    layer0_outputs(7207) <= inputs(40);
    layer0_outputs(7208) <= inputs(207);
    layer0_outputs(7209) <= inputs(128);
    layer0_outputs(7210) <= (inputs(251)) and not (inputs(239));
    layer0_outputs(7211) <= (inputs(123)) and not (inputs(73));
    layer0_outputs(7212) <= (inputs(223)) and not (inputs(107));
    layer0_outputs(7213) <= inputs(72);
    layer0_outputs(7214) <= (inputs(51)) or (inputs(110));
    layer0_outputs(7215) <= not(inputs(168)) or (inputs(219));
    layer0_outputs(7216) <= inputs(92);
    layer0_outputs(7217) <= inputs(207);
    layer0_outputs(7218) <= not((inputs(72)) xor (inputs(13)));
    layer0_outputs(7219) <= (inputs(120)) and not (inputs(228));
    layer0_outputs(7220) <= not(inputs(141));
    layer0_outputs(7221) <= not(inputs(153)) or (inputs(212));
    layer0_outputs(7222) <= not(inputs(200)) or (inputs(29));
    layer0_outputs(7223) <= not((inputs(212)) xor (inputs(7)));
    layer0_outputs(7224) <= (inputs(249)) and (inputs(79));
    layer0_outputs(7225) <= not((inputs(65)) or (inputs(171)));
    layer0_outputs(7226) <= (inputs(190)) and not (inputs(0));
    layer0_outputs(7227) <= not((inputs(176)) or (inputs(207)));
    layer0_outputs(7228) <= (inputs(218)) and not (inputs(232));
    layer0_outputs(7229) <= (inputs(188)) or (inputs(60));
    layer0_outputs(7230) <= not((inputs(131)) xor (inputs(206)));
    layer0_outputs(7231) <= not((inputs(19)) or (inputs(52)));
    layer0_outputs(7232) <= inputs(160);
    layer0_outputs(7233) <= not(inputs(72));
    layer0_outputs(7234) <= (inputs(177)) xor (inputs(73));
    layer0_outputs(7235) <= not(inputs(154)) or (inputs(164));
    layer0_outputs(7236) <= not(inputs(134)) or (inputs(67));
    layer0_outputs(7237) <= (inputs(175)) or (inputs(133));
    layer0_outputs(7238) <= not((inputs(130)) and (inputs(250)));
    layer0_outputs(7239) <= not(inputs(184)) or (inputs(204));
    layer0_outputs(7240) <= (inputs(18)) xor (inputs(212));
    layer0_outputs(7241) <= (inputs(121)) and not (inputs(237));
    layer0_outputs(7242) <= not(inputs(219)) or (inputs(23));
    layer0_outputs(7243) <= (inputs(85)) or (inputs(137));
    layer0_outputs(7244) <= (inputs(125)) or (inputs(107));
    layer0_outputs(7245) <= not(inputs(108)) or (inputs(249));
    layer0_outputs(7246) <= inputs(168);
    layer0_outputs(7247) <= (inputs(178)) xor (inputs(110));
    layer0_outputs(7248) <= not(inputs(246)) or (inputs(248));
    layer0_outputs(7249) <= (inputs(17)) xor (inputs(182));
    layer0_outputs(7250) <= not(inputs(171));
    layer0_outputs(7251) <= inputs(74);
    layer0_outputs(7252) <= (inputs(141)) or (inputs(163));
    layer0_outputs(7253) <= '0';
    layer0_outputs(7254) <= not((inputs(33)) xor (inputs(125)));
    layer0_outputs(7255) <= (inputs(72)) or (inputs(247));
    layer0_outputs(7256) <= not((inputs(131)) or (inputs(144)));
    layer0_outputs(7257) <= not(inputs(18));
    layer0_outputs(7258) <= (inputs(193)) or (inputs(90));
    layer0_outputs(7259) <= (inputs(123)) and not (inputs(237));
    layer0_outputs(7260) <= not(inputs(181)) or (inputs(141));
    layer0_outputs(7261) <= (inputs(135)) xor (inputs(19));
    layer0_outputs(7262) <= not((inputs(2)) xor (inputs(193)));
    layer0_outputs(7263) <= (inputs(129)) or (inputs(113));
    layer0_outputs(7264) <= (inputs(116)) and not (inputs(39));
    layer0_outputs(7265) <= not(inputs(30)) or (inputs(75));
    layer0_outputs(7266) <= not(inputs(138)) or (inputs(126));
    layer0_outputs(7267) <= not((inputs(79)) or (inputs(59)));
    layer0_outputs(7268) <= inputs(213);
    layer0_outputs(7269) <= not(inputs(196));
    layer0_outputs(7270) <= not((inputs(119)) xor (inputs(173)));
    layer0_outputs(7271) <= inputs(21);
    layer0_outputs(7272) <= not(inputs(231)) or (inputs(66));
    layer0_outputs(7273) <= inputs(87);
    layer0_outputs(7274) <= inputs(231);
    layer0_outputs(7275) <= '0';
    layer0_outputs(7276) <= not(inputs(20));
    layer0_outputs(7277) <= not(inputs(168)) or (inputs(242));
    layer0_outputs(7278) <= not(inputs(254));
    layer0_outputs(7279) <= not(inputs(131));
    layer0_outputs(7280) <= not((inputs(249)) xor (inputs(103)));
    layer0_outputs(7281) <= not(inputs(136)) or (inputs(224));
    layer0_outputs(7282) <= inputs(105);
    layer0_outputs(7283) <= not(inputs(79)) or (inputs(180));
    layer0_outputs(7284) <= not(inputs(131));
    layer0_outputs(7285) <= (inputs(207)) and not (inputs(240));
    layer0_outputs(7286) <= not(inputs(99));
    layer0_outputs(7287) <= inputs(104);
    layer0_outputs(7288) <= not((inputs(12)) xor (inputs(125)));
    layer0_outputs(7289) <= '0';
    layer0_outputs(7290) <= inputs(201);
    layer0_outputs(7291) <= not(inputs(89)) or (inputs(44));
    layer0_outputs(7292) <= inputs(172);
    layer0_outputs(7293) <= inputs(89);
    layer0_outputs(7294) <= inputs(112);
    layer0_outputs(7295) <= not(inputs(64));
    layer0_outputs(7296) <= not((inputs(148)) xor (inputs(221)));
    layer0_outputs(7297) <= not((inputs(130)) xor (inputs(118)));
    layer0_outputs(7298) <= inputs(124);
    layer0_outputs(7299) <= not((inputs(15)) xor (inputs(166)));
    layer0_outputs(7300) <= inputs(163);
    layer0_outputs(7301) <= (inputs(224)) and not (inputs(248));
    layer0_outputs(7302) <= not((inputs(143)) and (inputs(144)));
    layer0_outputs(7303) <= not((inputs(69)) xor (inputs(124)));
    layer0_outputs(7304) <= (inputs(231)) or (inputs(127));
    layer0_outputs(7305) <= (inputs(147)) or (inputs(250));
    layer0_outputs(7306) <= not(inputs(138)) or (inputs(243));
    layer0_outputs(7307) <= not((inputs(21)) or (inputs(166)));
    layer0_outputs(7308) <= (inputs(151)) xor (inputs(14));
    layer0_outputs(7309) <= not(inputs(155));
    layer0_outputs(7310) <= not(inputs(61));
    layer0_outputs(7311) <= inputs(110);
    layer0_outputs(7312) <= not(inputs(22)) or (inputs(114));
    layer0_outputs(7313) <= inputs(38);
    layer0_outputs(7314) <= not(inputs(29));
    layer0_outputs(7315) <= not(inputs(45));
    layer0_outputs(7316) <= (inputs(37)) or (inputs(53));
    layer0_outputs(7317) <= (inputs(89)) xor (inputs(19));
    layer0_outputs(7318) <= '1';
    layer0_outputs(7319) <= (inputs(11)) and not (inputs(208));
    layer0_outputs(7320) <= (inputs(39)) and not (inputs(13));
    layer0_outputs(7321) <= not(inputs(148));
    layer0_outputs(7322) <= (inputs(18)) and not (inputs(239));
    layer0_outputs(7323) <= (inputs(202)) and not (inputs(126));
    layer0_outputs(7324) <= (inputs(31)) and not (inputs(49));
    layer0_outputs(7325) <= not((inputs(30)) or (inputs(115)));
    layer0_outputs(7326) <= not((inputs(32)) xor (inputs(212)));
    layer0_outputs(7327) <= not(inputs(24));
    layer0_outputs(7328) <= (inputs(171)) or (inputs(41));
    layer0_outputs(7329) <= (inputs(144)) and (inputs(41));
    layer0_outputs(7330) <= not((inputs(61)) or (inputs(41)));
    layer0_outputs(7331) <= inputs(196);
    layer0_outputs(7332) <= inputs(138);
    layer0_outputs(7333) <= (inputs(57)) or (inputs(178));
    layer0_outputs(7334) <= not((inputs(201)) xor (inputs(43)));
    layer0_outputs(7335) <= not(inputs(141));
    layer0_outputs(7336) <= (inputs(53)) xor (inputs(98));
    layer0_outputs(7337) <= (inputs(30)) or (inputs(27));
    layer0_outputs(7338) <= inputs(234);
    layer0_outputs(7339) <= not((inputs(188)) xor (inputs(8)));
    layer0_outputs(7340) <= inputs(120);
    layer0_outputs(7341) <= inputs(98);
    layer0_outputs(7342) <= not((inputs(135)) or (inputs(51)));
    layer0_outputs(7343) <= not(inputs(233));
    layer0_outputs(7344) <= (inputs(152)) and not (inputs(81));
    layer0_outputs(7345) <= not(inputs(202)) or (inputs(83));
    layer0_outputs(7346) <= not(inputs(24)) or (inputs(208));
    layer0_outputs(7347) <= inputs(149);
    layer0_outputs(7348) <= not(inputs(233));
    layer0_outputs(7349) <= (inputs(164)) and not (inputs(9));
    layer0_outputs(7350) <= (inputs(185)) and not (inputs(128));
    layer0_outputs(7351) <= (inputs(201)) and not (inputs(23));
    layer0_outputs(7352) <= not(inputs(20));
    layer0_outputs(7353) <= not((inputs(199)) xor (inputs(58)));
    layer0_outputs(7354) <= (inputs(109)) xor (inputs(214));
    layer0_outputs(7355) <= (inputs(224)) or (inputs(89));
    layer0_outputs(7356) <= not(inputs(71)) or (inputs(240));
    layer0_outputs(7357) <= not((inputs(23)) xor (inputs(140)));
    layer0_outputs(7358) <= (inputs(211)) or (inputs(28));
    layer0_outputs(7359) <= inputs(88);
    layer0_outputs(7360) <= not((inputs(48)) or (inputs(157)));
    layer0_outputs(7361) <= not(inputs(83)) or (inputs(130));
    layer0_outputs(7362) <= not((inputs(107)) or (inputs(137)));
    layer0_outputs(7363) <= (inputs(209)) or (inputs(105));
    layer0_outputs(7364) <= (inputs(56)) or (inputs(219));
    layer0_outputs(7365) <= not((inputs(88)) or (inputs(66)));
    layer0_outputs(7366) <= not(inputs(106)) or (inputs(7));
    layer0_outputs(7367) <= (inputs(39)) xor (inputs(245));
    layer0_outputs(7368) <= (inputs(31)) and not (inputs(26));
    layer0_outputs(7369) <= not(inputs(174)) or (inputs(246));
    layer0_outputs(7370) <= not((inputs(120)) xor (inputs(224)));
    layer0_outputs(7371) <= not(inputs(70)) or (inputs(254));
    layer0_outputs(7372) <= not(inputs(183)) or (inputs(96));
    layer0_outputs(7373) <= not(inputs(240));
    layer0_outputs(7374) <= (inputs(85)) xor (inputs(80));
    layer0_outputs(7375) <= not((inputs(76)) and (inputs(108)));
    layer0_outputs(7376) <= (inputs(16)) or (inputs(24));
    layer0_outputs(7377) <= '0';
    layer0_outputs(7378) <= (inputs(36)) xor (inputs(134));
    layer0_outputs(7379) <= inputs(33);
    layer0_outputs(7380) <= not((inputs(48)) xor (inputs(35)));
    layer0_outputs(7381) <= not((inputs(99)) or (inputs(242)));
    layer0_outputs(7382) <= (inputs(209)) or (inputs(179));
    layer0_outputs(7383) <= (inputs(37)) xor (inputs(237));
    layer0_outputs(7384) <= '0';
    layer0_outputs(7385) <= (inputs(113)) xor (inputs(154));
    layer0_outputs(7386) <= '1';
    layer0_outputs(7387) <= not(inputs(86)) or (inputs(157));
    layer0_outputs(7388) <= not(inputs(169));
    layer0_outputs(7389) <= (inputs(174)) xor (inputs(228));
    layer0_outputs(7390) <= (inputs(249)) and not (inputs(47));
    layer0_outputs(7391) <= inputs(170);
    layer0_outputs(7392) <= (inputs(108)) and not (inputs(36));
    layer0_outputs(7393) <= inputs(72);
    layer0_outputs(7394) <= (inputs(184)) and not (inputs(145));
    layer0_outputs(7395) <= inputs(118);
    layer0_outputs(7396) <= not(inputs(127));
    layer0_outputs(7397) <= (inputs(134)) or (inputs(6));
    layer0_outputs(7398) <= '0';
    layer0_outputs(7399) <= not(inputs(254)) or (inputs(174));
    layer0_outputs(7400) <= not(inputs(204));
    layer0_outputs(7401) <= not((inputs(189)) or (inputs(182)));
    layer0_outputs(7402) <= inputs(74);
    layer0_outputs(7403) <= (inputs(156)) xor (inputs(50));
    layer0_outputs(7404) <= not(inputs(47)) or (inputs(13));
    layer0_outputs(7405) <= inputs(158);
    layer0_outputs(7406) <= not(inputs(179));
    layer0_outputs(7407) <= inputs(13);
    layer0_outputs(7408) <= not(inputs(104));
    layer0_outputs(7409) <= not(inputs(98)) or (inputs(148));
    layer0_outputs(7410) <= not(inputs(118));
    layer0_outputs(7411) <= inputs(43);
    layer0_outputs(7412) <= (inputs(231)) xor (inputs(161));
    layer0_outputs(7413) <= '0';
    layer0_outputs(7414) <= '0';
    layer0_outputs(7415) <= not((inputs(87)) and (inputs(45)));
    layer0_outputs(7416) <= (inputs(102)) or (inputs(99));
    layer0_outputs(7417) <= (inputs(235)) or (inputs(215));
    layer0_outputs(7418) <= '1';
    layer0_outputs(7419) <= not((inputs(153)) xor (inputs(65)));
    layer0_outputs(7420) <= (inputs(224)) xor (inputs(232));
    layer0_outputs(7421) <= inputs(101);
    layer0_outputs(7422) <= (inputs(186)) and not (inputs(32));
    layer0_outputs(7423) <= not((inputs(191)) xor (inputs(96)));
    layer0_outputs(7424) <= not((inputs(111)) xor (inputs(136)));
    layer0_outputs(7425) <= not((inputs(6)) or (inputs(101)));
    layer0_outputs(7426) <= (inputs(78)) and not (inputs(245));
    layer0_outputs(7427) <= inputs(166);
    layer0_outputs(7428) <= inputs(195);
    layer0_outputs(7429) <= (inputs(244)) xor (inputs(73));
    layer0_outputs(7430) <= not((inputs(234)) or (inputs(123)));
    layer0_outputs(7431) <= (inputs(170)) and not (inputs(35));
    layer0_outputs(7432) <= not((inputs(0)) xor (inputs(117)));
    layer0_outputs(7433) <= not(inputs(119));
    layer0_outputs(7434) <= not(inputs(65));
    layer0_outputs(7435) <= (inputs(56)) or (inputs(38));
    layer0_outputs(7436) <= not(inputs(23));
    layer0_outputs(7437) <= not((inputs(231)) or (inputs(28)));
    layer0_outputs(7438) <= (inputs(183)) and not (inputs(139));
    layer0_outputs(7439) <= '1';
    layer0_outputs(7440) <= not((inputs(12)) and (inputs(36)));
    layer0_outputs(7441) <= inputs(115);
    layer0_outputs(7442) <= inputs(45);
    layer0_outputs(7443) <= (inputs(123)) and not (inputs(190));
    layer0_outputs(7444) <= (inputs(83)) and not (inputs(246));
    layer0_outputs(7445) <= not(inputs(197)) or (inputs(192));
    layer0_outputs(7446) <= not(inputs(23)) or (inputs(49));
    layer0_outputs(7447) <= inputs(83);
    layer0_outputs(7448) <= (inputs(128)) or (inputs(109));
    layer0_outputs(7449) <= (inputs(102)) xor (inputs(247));
    layer0_outputs(7450) <= inputs(26);
    layer0_outputs(7451) <= (inputs(165)) and not (inputs(112));
    layer0_outputs(7452) <= not((inputs(245)) xor (inputs(181)));
    layer0_outputs(7453) <= (inputs(242)) xor (inputs(215));
    layer0_outputs(7454) <= not(inputs(45)) or (inputs(72));
    layer0_outputs(7455) <= (inputs(143)) and not (inputs(222));
    layer0_outputs(7456) <= not((inputs(207)) and (inputs(2)));
    layer0_outputs(7457) <= inputs(112);
    layer0_outputs(7458) <= not((inputs(86)) xor (inputs(230)));
    layer0_outputs(7459) <= not(inputs(127));
    layer0_outputs(7460) <= not((inputs(12)) xor (inputs(193)));
    layer0_outputs(7461) <= not(inputs(110)) or (inputs(130));
    layer0_outputs(7462) <= (inputs(183)) and not (inputs(246));
    layer0_outputs(7463) <= (inputs(50)) and not (inputs(0));
    layer0_outputs(7464) <= (inputs(35)) xor (inputs(50));
    layer0_outputs(7465) <= (inputs(107)) or (inputs(217));
    layer0_outputs(7466) <= '0';
    layer0_outputs(7467) <= (inputs(198)) xor (inputs(199));
    layer0_outputs(7468) <= inputs(51);
    layer0_outputs(7469) <= (inputs(71)) and (inputs(187));
    layer0_outputs(7470) <= not((inputs(209)) or (inputs(23)));
    layer0_outputs(7471) <= not((inputs(50)) or (inputs(105)));
    layer0_outputs(7472) <= not(inputs(104));
    layer0_outputs(7473) <= (inputs(207)) xor (inputs(94));
    layer0_outputs(7474) <= not(inputs(37)) or (inputs(4));
    layer0_outputs(7475) <= (inputs(236)) and not (inputs(47));
    layer0_outputs(7476) <= not((inputs(173)) or (inputs(71)));
    layer0_outputs(7477) <= not(inputs(83));
    layer0_outputs(7478) <= inputs(188);
    layer0_outputs(7479) <= not((inputs(85)) xor (inputs(80)));
    layer0_outputs(7480) <= not(inputs(152)) or (inputs(149));
    layer0_outputs(7481) <= inputs(153);
    layer0_outputs(7482) <= not(inputs(199));
    layer0_outputs(7483) <= not(inputs(24));
    layer0_outputs(7484) <= (inputs(15)) xor (inputs(95));
    layer0_outputs(7485) <= (inputs(7)) and not (inputs(246));
    layer0_outputs(7486) <= inputs(52);
    layer0_outputs(7487) <= not(inputs(167));
    layer0_outputs(7488) <= not((inputs(5)) xor (inputs(71)));
    layer0_outputs(7489) <= not((inputs(68)) or (inputs(164)));
    layer0_outputs(7490) <= not((inputs(211)) or (inputs(90)));
    layer0_outputs(7491) <= not((inputs(41)) or (inputs(158)));
    layer0_outputs(7492) <= not((inputs(149)) or (inputs(102)));
    layer0_outputs(7493) <= not(inputs(60)) or (inputs(193));
    layer0_outputs(7494) <= (inputs(91)) and not (inputs(18));
    layer0_outputs(7495) <= not(inputs(90));
    layer0_outputs(7496) <= (inputs(90)) or (inputs(129));
    layer0_outputs(7497) <= not(inputs(74));
    layer0_outputs(7498) <= inputs(69);
    layer0_outputs(7499) <= not((inputs(99)) xor (inputs(77)));
    layer0_outputs(7500) <= (inputs(85)) and not (inputs(9));
    layer0_outputs(7501) <= '1';
    layer0_outputs(7502) <= not(inputs(61)) or (inputs(35));
    layer0_outputs(7503) <= inputs(89);
    layer0_outputs(7504) <= not(inputs(210));
    layer0_outputs(7505) <= not((inputs(84)) or (inputs(49)));
    layer0_outputs(7506) <= not((inputs(209)) xor (inputs(57)));
    layer0_outputs(7507) <= not((inputs(77)) xor (inputs(183)));
    layer0_outputs(7508) <= inputs(108);
    layer0_outputs(7509) <= not((inputs(232)) or (inputs(78)));
    layer0_outputs(7510) <= inputs(122);
    layer0_outputs(7511) <= (inputs(75)) xor (inputs(216));
    layer0_outputs(7512) <= not(inputs(207));
    layer0_outputs(7513) <= not(inputs(157)) or (inputs(95));
    layer0_outputs(7514) <= inputs(127);
    layer0_outputs(7515) <= (inputs(141)) or (inputs(52));
    layer0_outputs(7516) <= (inputs(66)) and not (inputs(228));
    layer0_outputs(7517) <= not((inputs(57)) xor (inputs(171)));
    layer0_outputs(7518) <= not(inputs(109));
    layer0_outputs(7519) <= not((inputs(193)) xor (inputs(68)));
    layer0_outputs(7520) <= not(inputs(226)) or (inputs(16));
    layer0_outputs(7521) <= not(inputs(39)) or (inputs(12));
    layer0_outputs(7522) <= inputs(161);
    layer0_outputs(7523) <= (inputs(228)) xor (inputs(100));
    layer0_outputs(7524) <= not(inputs(66));
    layer0_outputs(7525) <= not((inputs(37)) or (inputs(167)));
    layer0_outputs(7526) <= inputs(119);
    layer0_outputs(7527) <= not(inputs(218)) or (inputs(58));
    layer0_outputs(7528) <= (inputs(237)) xor (inputs(111));
    layer0_outputs(7529) <= not(inputs(157)) or (inputs(30));
    layer0_outputs(7530) <= (inputs(203)) xor (inputs(140));
    layer0_outputs(7531) <= (inputs(53)) and not (inputs(233));
    layer0_outputs(7532) <= (inputs(244)) and not (inputs(248));
    layer0_outputs(7533) <= not((inputs(201)) xor (inputs(206)));
    layer0_outputs(7534) <= (inputs(63)) and (inputs(8));
    layer0_outputs(7535) <= not(inputs(217));
    layer0_outputs(7536) <= (inputs(102)) and not (inputs(31));
    layer0_outputs(7537) <= '1';
    layer0_outputs(7538) <= (inputs(0)) xor (inputs(170));
    layer0_outputs(7539) <= not((inputs(88)) xor (inputs(146)));
    layer0_outputs(7540) <= '1';
    layer0_outputs(7541) <= (inputs(188)) xor (inputs(7));
    layer0_outputs(7542) <= not((inputs(41)) or (inputs(232)));
    layer0_outputs(7543) <= not((inputs(142)) or (inputs(176)));
    layer0_outputs(7544) <= inputs(223);
    layer0_outputs(7545) <= (inputs(185)) and not (inputs(247));
    layer0_outputs(7546) <= not(inputs(137)) or (inputs(89));
    layer0_outputs(7547) <= (inputs(172)) or (inputs(70));
    layer0_outputs(7548) <= not((inputs(27)) or (inputs(159)));
    layer0_outputs(7549) <= (inputs(156)) or (inputs(145));
    layer0_outputs(7550) <= not((inputs(159)) or (inputs(152)));
    layer0_outputs(7551) <= not((inputs(89)) or (inputs(212)));
    layer0_outputs(7552) <= not(inputs(131));
    layer0_outputs(7553) <= not(inputs(138)) or (inputs(133));
    layer0_outputs(7554) <= not(inputs(118)) or (inputs(233));
    layer0_outputs(7555) <= '0';
    layer0_outputs(7556) <= (inputs(78)) xor (inputs(133));
    layer0_outputs(7557) <= not((inputs(25)) or (inputs(170)));
    layer0_outputs(7558) <= not(inputs(110));
    layer0_outputs(7559) <= (inputs(87)) and not (inputs(211));
    layer0_outputs(7560) <= not((inputs(134)) and (inputs(13)));
    layer0_outputs(7561) <= not(inputs(85)) or (inputs(246));
    layer0_outputs(7562) <= not((inputs(70)) xor (inputs(91)));
    layer0_outputs(7563) <= not(inputs(193));
    layer0_outputs(7564) <= not((inputs(55)) xor (inputs(224)));
    layer0_outputs(7565) <= not((inputs(252)) or (inputs(24)));
    layer0_outputs(7566) <= not(inputs(255)) or (inputs(118));
    layer0_outputs(7567) <= inputs(116);
    layer0_outputs(7568) <= not(inputs(36));
    layer0_outputs(7569) <= inputs(122);
    layer0_outputs(7570) <= (inputs(19)) xor (inputs(204));
    layer0_outputs(7571) <= not((inputs(243)) or (inputs(152)));
    layer0_outputs(7572) <= not(inputs(213));
    layer0_outputs(7573) <= (inputs(49)) and (inputs(142));
    layer0_outputs(7574) <= not((inputs(249)) and (inputs(129)));
    layer0_outputs(7575) <= not(inputs(233));
    layer0_outputs(7576) <= not((inputs(162)) or (inputs(218)));
    layer0_outputs(7577) <= (inputs(235)) or (inputs(123));
    layer0_outputs(7578) <= (inputs(231)) xor (inputs(174));
    layer0_outputs(7579) <= inputs(92);
    layer0_outputs(7580) <= inputs(1);
    layer0_outputs(7581) <= not(inputs(52)) or (inputs(10));
    layer0_outputs(7582) <= not(inputs(100)) or (inputs(210));
    layer0_outputs(7583) <= not(inputs(60)) or (inputs(210));
    layer0_outputs(7584) <= (inputs(151)) and not (inputs(75));
    layer0_outputs(7585) <= '1';
    layer0_outputs(7586) <= not((inputs(160)) xor (inputs(83)));
    layer0_outputs(7587) <= (inputs(134)) and not (inputs(64));
    layer0_outputs(7588) <= (inputs(160)) xor (inputs(39));
    layer0_outputs(7589) <= not(inputs(172)) or (inputs(241));
    layer0_outputs(7590) <= inputs(87);
    layer0_outputs(7591) <= not((inputs(250)) xor (inputs(242)));
    layer0_outputs(7592) <= (inputs(254)) and not (inputs(153));
    layer0_outputs(7593) <= not((inputs(237)) or (inputs(229)));
    layer0_outputs(7594) <= inputs(122);
    layer0_outputs(7595) <= not(inputs(153));
    layer0_outputs(7596) <= (inputs(107)) and not (inputs(242));
    layer0_outputs(7597) <= inputs(162);
    layer0_outputs(7598) <= (inputs(182)) xor (inputs(40));
    layer0_outputs(7599) <= inputs(156);
    layer0_outputs(7600) <= (inputs(87)) xor (inputs(193));
    layer0_outputs(7601) <= (inputs(245)) xor (inputs(81));
    layer0_outputs(7602) <= (inputs(221)) and not (inputs(39));
    layer0_outputs(7603) <= not(inputs(74));
    layer0_outputs(7604) <= not(inputs(163));
    layer0_outputs(7605) <= not((inputs(141)) xor (inputs(173)));
    layer0_outputs(7606) <= '1';
    layer0_outputs(7607) <= not((inputs(227)) xor (inputs(143)));
    layer0_outputs(7608) <= inputs(226);
    layer0_outputs(7609) <= not(inputs(215)) or (inputs(183));
    layer0_outputs(7610) <= inputs(109);
    layer0_outputs(7611) <= (inputs(69)) or (inputs(82));
    layer0_outputs(7612) <= (inputs(225)) and not (inputs(169));
    layer0_outputs(7613) <= inputs(93);
    layer0_outputs(7614) <= (inputs(236)) or (inputs(112));
    layer0_outputs(7615) <= not((inputs(197)) or (inputs(230)));
    layer0_outputs(7616) <= not((inputs(226)) and (inputs(153)));
    layer0_outputs(7617) <= (inputs(15)) and (inputs(2));
    layer0_outputs(7618) <= inputs(58);
    layer0_outputs(7619) <= inputs(225);
    layer0_outputs(7620) <= (inputs(176)) and not (inputs(116));
    layer0_outputs(7621) <= (inputs(56)) xor (inputs(224));
    layer0_outputs(7622) <= not((inputs(151)) or (inputs(6)));
    layer0_outputs(7623) <= not((inputs(59)) and (inputs(59)));
    layer0_outputs(7624) <= not((inputs(119)) or (inputs(16)));
    layer0_outputs(7625) <= not(inputs(49)) or (inputs(192));
    layer0_outputs(7626) <= not((inputs(182)) or (inputs(18)));
    layer0_outputs(7627) <= not(inputs(181));
    layer0_outputs(7628) <= (inputs(28)) or (inputs(150));
    layer0_outputs(7629) <= inputs(171);
    layer0_outputs(7630) <= (inputs(19)) or (inputs(140));
    layer0_outputs(7631) <= not((inputs(131)) and (inputs(31)));
    layer0_outputs(7632) <= (inputs(12)) and not (inputs(211));
    layer0_outputs(7633) <= not((inputs(58)) xor (inputs(49)));
    layer0_outputs(7634) <= (inputs(98)) xor (inputs(55));
    layer0_outputs(7635) <= not((inputs(200)) or (inputs(51)));
    layer0_outputs(7636) <= (inputs(186)) or (inputs(130));
    layer0_outputs(7637) <= not((inputs(198)) or (inputs(69)));
    layer0_outputs(7638) <= '1';
    layer0_outputs(7639) <= not((inputs(250)) or (inputs(187)));
    layer0_outputs(7640) <= inputs(209);
    layer0_outputs(7641) <= not((inputs(67)) or (inputs(36)));
    layer0_outputs(7642) <= not(inputs(134));
    layer0_outputs(7643) <= inputs(174);
    layer0_outputs(7644) <= (inputs(76)) and not (inputs(128));
    layer0_outputs(7645) <= not(inputs(79)) or (inputs(62));
    layer0_outputs(7646) <= (inputs(227)) or (inputs(117));
    layer0_outputs(7647) <= not((inputs(29)) xor (inputs(140)));
    layer0_outputs(7648) <= not(inputs(169));
    layer0_outputs(7649) <= (inputs(221)) and (inputs(17));
    layer0_outputs(7650) <= (inputs(186)) and not (inputs(84));
    layer0_outputs(7651) <= inputs(167);
    layer0_outputs(7652) <= '1';
    layer0_outputs(7653) <= (inputs(203)) and not (inputs(162));
    layer0_outputs(7654) <= not((inputs(116)) xor (inputs(28)));
    layer0_outputs(7655) <= not((inputs(132)) xor (inputs(15)));
    layer0_outputs(7656) <= not((inputs(172)) and (inputs(207)));
    layer0_outputs(7657) <= inputs(125);
    layer0_outputs(7658) <= inputs(222);
    layer0_outputs(7659) <= inputs(40);
    layer0_outputs(7660) <= inputs(12);
    layer0_outputs(7661) <= not((inputs(42)) or (inputs(22)));
    layer0_outputs(7662) <= not((inputs(149)) xor (inputs(187)));
    layer0_outputs(7663) <= inputs(114);
    layer0_outputs(7664) <= (inputs(63)) and (inputs(19));
    layer0_outputs(7665) <= (inputs(184)) and not (inputs(109));
    layer0_outputs(7666) <= (inputs(56)) or (inputs(78));
    layer0_outputs(7667) <= not((inputs(36)) and (inputs(246)));
    layer0_outputs(7668) <= not(inputs(149)) or (inputs(229));
    layer0_outputs(7669) <= not(inputs(29)) or (inputs(112));
    layer0_outputs(7670) <= not(inputs(145)) or (inputs(29));
    layer0_outputs(7671) <= (inputs(104)) or (inputs(115));
    layer0_outputs(7672) <= (inputs(234)) and not (inputs(59));
    layer0_outputs(7673) <= not((inputs(156)) or (inputs(56)));
    layer0_outputs(7674) <= inputs(159);
    layer0_outputs(7675) <= '0';
    layer0_outputs(7676) <= (inputs(93)) or (inputs(125));
    layer0_outputs(7677) <= '1';
    layer0_outputs(7678) <= not(inputs(160)) or (inputs(245));
    layer0_outputs(7679) <= inputs(100);
    layer0_outputs(7680) <= not(inputs(163)) or (inputs(33));
    layer0_outputs(7681) <= inputs(159);
    layer0_outputs(7682) <= (inputs(246)) xor (inputs(203));
    layer0_outputs(7683) <= not((inputs(175)) or (inputs(122)));
    layer0_outputs(7684) <= '0';
    layer0_outputs(7685) <= not(inputs(105)) or (inputs(236));
    layer0_outputs(7686) <= not(inputs(146)) or (inputs(204));
    layer0_outputs(7687) <= inputs(38);
    layer0_outputs(7688) <= not((inputs(172)) xor (inputs(211)));
    layer0_outputs(7689) <= (inputs(87)) and not (inputs(150));
    layer0_outputs(7690) <= (inputs(48)) xor (inputs(61));
    layer0_outputs(7691) <= (inputs(66)) and not (inputs(23));
    layer0_outputs(7692) <= (inputs(49)) xor (inputs(132));
    layer0_outputs(7693) <= (inputs(67)) and not (inputs(221));
    layer0_outputs(7694) <= not(inputs(220)) or (inputs(155));
    layer0_outputs(7695) <= not(inputs(153)) or (inputs(126));
    layer0_outputs(7696) <= not(inputs(216)) or (inputs(11));
    layer0_outputs(7697) <= not(inputs(159));
    layer0_outputs(7698) <= not((inputs(27)) xor (inputs(233)));
    layer0_outputs(7699) <= (inputs(108)) or (inputs(66));
    layer0_outputs(7700) <= not(inputs(132)) or (inputs(162));
    layer0_outputs(7701) <= not(inputs(92)) or (inputs(98));
    layer0_outputs(7702) <= (inputs(16)) and not (inputs(124));
    layer0_outputs(7703) <= not(inputs(121));
    layer0_outputs(7704) <= (inputs(160)) or (inputs(249));
    layer0_outputs(7705) <= (inputs(190)) or (inputs(29));
    layer0_outputs(7706) <= (inputs(88)) xor (inputs(30));
    layer0_outputs(7707) <= (inputs(21)) and not (inputs(176));
    layer0_outputs(7708) <= not((inputs(123)) or (inputs(112)));
    layer0_outputs(7709) <= (inputs(7)) or (inputs(95));
    layer0_outputs(7710) <= not((inputs(210)) and (inputs(250)));
    layer0_outputs(7711) <= (inputs(29)) xor (inputs(136));
    layer0_outputs(7712) <= (inputs(14)) and not (inputs(142));
    layer0_outputs(7713) <= not((inputs(24)) and (inputs(28)));
    layer0_outputs(7714) <= '0';
    layer0_outputs(7715) <= inputs(232);
    layer0_outputs(7716) <= inputs(83);
    layer0_outputs(7717) <= inputs(236);
    layer0_outputs(7718) <= not(inputs(52)) or (inputs(244));
    layer0_outputs(7719) <= not(inputs(23)) or (inputs(31));
    layer0_outputs(7720) <= not((inputs(8)) xor (inputs(154)));
    layer0_outputs(7721) <= not(inputs(149)) or (inputs(167));
    layer0_outputs(7722) <= inputs(56);
    layer0_outputs(7723) <= (inputs(56)) and not (inputs(168));
    layer0_outputs(7724) <= (inputs(71)) and not (inputs(168));
    layer0_outputs(7725) <= not(inputs(62));
    layer0_outputs(7726) <= (inputs(135)) xor (inputs(165));
    layer0_outputs(7727) <= not((inputs(113)) or (inputs(23)));
    layer0_outputs(7728) <= not((inputs(37)) or (inputs(167)));
    layer0_outputs(7729) <= not(inputs(214)) or (inputs(15));
    layer0_outputs(7730) <= not(inputs(53));
    layer0_outputs(7731) <= (inputs(243)) xor (inputs(238));
    layer0_outputs(7732) <= not(inputs(137)) or (inputs(241));
    layer0_outputs(7733) <= not((inputs(21)) xor (inputs(52)));
    layer0_outputs(7734) <= not(inputs(69)) or (inputs(77));
    layer0_outputs(7735) <= not((inputs(46)) or (inputs(38)));
    layer0_outputs(7736) <= not(inputs(161)) or (inputs(32));
    layer0_outputs(7737) <= (inputs(35)) xor (inputs(246));
    layer0_outputs(7738) <= inputs(71);
    layer0_outputs(7739) <= inputs(23);
    layer0_outputs(7740) <= inputs(221);
    layer0_outputs(7741) <= (inputs(226)) xor (inputs(94));
    layer0_outputs(7742) <= (inputs(53)) and not (inputs(55));
    layer0_outputs(7743) <= (inputs(62)) and not (inputs(36));
    layer0_outputs(7744) <= not(inputs(198)) or (inputs(194));
    layer0_outputs(7745) <= not(inputs(199));
    layer0_outputs(7746) <= not(inputs(59)) or (inputs(182));
    layer0_outputs(7747) <= not((inputs(181)) or (inputs(9)));
    layer0_outputs(7748) <= (inputs(39)) xor (inputs(69));
    layer0_outputs(7749) <= (inputs(85)) or (inputs(183));
    layer0_outputs(7750) <= not((inputs(35)) and (inputs(222)));
    layer0_outputs(7751) <= not((inputs(113)) and (inputs(49)));
    layer0_outputs(7752) <= (inputs(200)) or (inputs(100));
    layer0_outputs(7753) <= (inputs(159)) and not (inputs(253));
    layer0_outputs(7754) <= inputs(89);
    layer0_outputs(7755) <= '1';
    layer0_outputs(7756) <= inputs(219);
    layer0_outputs(7757) <= (inputs(86)) and not (inputs(51));
    layer0_outputs(7758) <= (inputs(57)) xor (inputs(12));
    layer0_outputs(7759) <= not(inputs(77));
    layer0_outputs(7760) <= not((inputs(212)) or (inputs(206)));
    layer0_outputs(7761) <= not((inputs(102)) xor (inputs(253)));
    layer0_outputs(7762) <= not(inputs(168));
    layer0_outputs(7763) <= inputs(3);
    layer0_outputs(7764) <= not(inputs(251));
    layer0_outputs(7765) <= not((inputs(33)) xor (inputs(196)));
    layer0_outputs(7766) <= (inputs(157)) or (inputs(125));
    layer0_outputs(7767) <= (inputs(31)) and not (inputs(145));
    layer0_outputs(7768) <= not((inputs(35)) or (inputs(230)));
    layer0_outputs(7769) <= (inputs(146)) or (inputs(174));
    layer0_outputs(7770) <= inputs(214);
    layer0_outputs(7771) <= not((inputs(136)) or (inputs(244)));
    layer0_outputs(7772) <= not(inputs(20)) or (inputs(116));
    layer0_outputs(7773) <= (inputs(216)) or (inputs(30));
    layer0_outputs(7774) <= not(inputs(251));
    layer0_outputs(7775) <= inputs(226);
    layer0_outputs(7776) <= '0';
    layer0_outputs(7777) <= not(inputs(131)) or (inputs(234));
    layer0_outputs(7778) <= not((inputs(148)) or (inputs(32)));
    layer0_outputs(7779) <= not(inputs(217));
    layer0_outputs(7780) <= not(inputs(192));
    layer0_outputs(7781) <= inputs(242);
    layer0_outputs(7782) <= inputs(247);
    layer0_outputs(7783) <= not((inputs(99)) xor (inputs(175)));
    layer0_outputs(7784) <= (inputs(226)) or (inputs(154));
    layer0_outputs(7785) <= (inputs(199)) and not (inputs(62));
    layer0_outputs(7786) <= not((inputs(36)) or (inputs(131)));
    layer0_outputs(7787) <= (inputs(167)) and not (inputs(60));
    layer0_outputs(7788) <= not((inputs(130)) or (inputs(183)));
    layer0_outputs(7789) <= not(inputs(196));
    layer0_outputs(7790) <= not(inputs(101)) or (inputs(105));
    layer0_outputs(7791) <= not((inputs(133)) xor (inputs(165)));
    layer0_outputs(7792) <= (inputs(153)) and not (inputs(38));
    layer0_outputs(7793) <= not((inputs(178)) xor (inputs(137)));
    layer0_outputs(7794) <= inputs(141);
    layer0_outputs(7795) <= inputs(195);
    layer0_outputs(7796) <= inputs(78);
    layer0_outputs(7797) <= inputs(24);
    layer0_outputs(7798) <= not((inputs(59)) or (inputs(96)));
    layer0_outputs(7799) <= inputs(74);
    layer0_outputs(7800) <= not(inputs(119)) or (inputs(159));
    layer0_outputs(7801) <= not(inputs(169)) or (inputs(181));
    layer0_outputs(7802) <= not(inputs(107)) or (inputs(62));
    layer0_outputs(7803) <= (inputs(25)) and not (inputs(25));
    layer0_outputs(7804) <= not((inputs(161)) xor (inputs(72)));
    layer0_outputs(7805) <= '1';
    layer0_outputs(7806) <= (inputs(24)) or (inputs(187));
    layer0_outputs(7807) <= not((inputs(159)) or (inputs(18)));
    layer0_outputs(7808) <= (inputs(144)) or (inputs(79));
    layer0_outputs(7809) <= inputs(163);
    layer0_outputs(7810) <= '1';
    layer0_outputs(7811) <= (inputs(170)) xor (inputs(118));
    layer0_outputs(7812) <= not(inputs(197)) or (inputs(149));
    layer0_outputs(7813) <= (inputs(109)) or (inputs(229));
    layer0_outputs(7814) <= inputs(115);
    layer0_outputs(7815) <= not((inputs(174)) xor (inputs(242)));
    layer0_outputs(7816) <= '1';
    layer0_outputs(7817) <= not(inputs(149));
    layer0_outputs(7818) <= not(inputs(118)) or (inputs(226));
    layer0_outputs(7819) <= not((inputs(165)) xor (inputs(95)));
    layer0_outputs(7820) <= not(inputs(189));
    layer0_outputs(7821) <= not((inputs(204)) and (inputs(234)));
    layer0_outputs(7822) <= not(inputs(83));
    layer0_outputs(7823) <= inputs(82);
    layer0_outputs(7824) <= (inputs(203)) and not (inputs(250));
    layer0_outputs(7825) <= '1';
    layer0_outputs(7826) <= (inputs(125)) or (inputs(74));
    layer0_outputs(7827) <= not((inputs(150)) xor (inputs(18)));
    layer0_outputs(7828) <= (inputs(11)) xor (inputs(228));
    layer0_outputs(7829) <= not(inputs(84)) or (inputs(190));
    layer0_outputs(7830) <= (inputs(119)) or (inputs(102));
    layer0_outputs(7831) <= not((inputs(90)) xor (inputs(185)));
    layer0_outputs(7832) <= not((inputs(222)) xor (inputs(230)));
    layer0_outputs(7833) <= inputs(176);
    layer0_outputs(7834) <= inputs(158);
    layer0_outputs(7835) <= (inputs(202)) and not (inputs(159));
    layer0_outputs(7836) <= (inputs(107)) and not (inputs(16));
    layer0_outputs(7837) <= (inputs(58)) and not (inputs(131));
    layer0_outputs(7838) <= not((inputs(180)) or (inputs(49)));
    layer0_outputs(7839) <= not(inputs(246)) or (inputs(144));
    layer0_outputs(7840) <= (inputs(31)) and (inputs(16));
    layer0_outputs(7841) <= not((inputs(116)) or (inputs(131)));
    layer0_outputs(7842) <= not((inputs(146)) or (inputs(119)));
    layer0_outputs(7843) <= inputs(158);
    layer0_outputs(7844) <= inputs(157);
    layer0_outputs(7845) <= not(inputs(73));
    layer0_outputs(7846) <= not((inputs(134)) or (inputs(111)));
    layer0_outputs(7847) <= not((inputs(186)) xor (inputs(43)));
    layer0_outputs(7848) <= not(inputs(247)) or (inputs(68));
    layer0_outputs(7849) <= not(inputs(9));
    layer0_outputs(7850) <= not((inputs(247)) and (inputs(239)));
    layer0_outputs(7851) <= not(inputs(238)) or (inputs(252));
    layer0_outputs(7852) <= inputs(139);
    layer0_outputs(7853) <= not(inputs(191)) or (inputs(251));
    layer0_outputs(7854) <= not(inputs(133));
    layer0_outputs(7855) <= inputs(51);
    layer0_outputs(7856) <= not(inputs(199)) or (inputs(213));
    layer0_outputs(7857) <= (inputs(241)) or (inputs(21));
    layer0_outputs(7858) <= inputs(211);
    layer0_outputs(7859) <= (inputs(109)) or (inputs(201));
    layer0_outputs(7860) <= (inputs(46)) or (inputs(185));
    layer0_outputs(7861) <= not((inputs(19)) xor (inputs(154)));
    layer0_outputs(7862) <= not(inputs(39)) or (inputs(131));
    layer0_outputs(7863) <= not((inputs(136)) xor (inputs(237)));
    layer0_outputs(7864) <= '1';
    layer0_outputs(7865) <= (inputs(178)) and not (inputs(126));
    layer0_outputs(7866) <= not((inputs(182)) or (inputs(67)));
    layer0_outputs(7867) <= not(inputs(116));
    layer0_outputs(7868) <= (inputs(210)) or (inputs(93));
    layer0_outputs(7869) <= (inputs(39)) xor (inputs(10));
    layer0_outputs(7870) <= not(inputs(119)) or (inputs(190));
    layer0_outputs(7871) <= inputs(73);
    layer0_outputs(7872) <= not((inputs(86)) or (inputs(94)));
    layer0_outputs(7873) <= (inputs(8)) xor (inputs(167));
    layer0_outputs(7874) <= '1';
    layer0_outputs(7875) <= not(inputs(73));
    layer0_outputs(7876) <= (inputs(1)) xor (inputs(108));
    layer0_outputs(7877) <= not((inputs(35)) xor (inputs(102)));
    layer0_outputs(7878) <= (inputs(103)) and not (inputs(219));
    layer0_outputs(7879) <= inputs(38);
    layer0_outputs(7880) <= (inputs(86)) and not (inputs(124));
    layer0_outputs(7881) <= not((inputs(57)) xor (inputs(10)));
    layer0_outputs(7882) <= not((inputs(37)) or (inputs(109)));
    layer0_outputs(7883) <= (inputs(199)) xor (inputs(16));
    layer0_outputs(7884) <= not(inputs(183)) or (inputs(225));
    layer0_outputs(7885) <= not((inputs(244)) and (inputs(52)));
    layer0_outputs(7886) <= (inputs(153)) or (inputs(236));
    layer0_outputs(7887) <= (inputs(186)) and not (inputs(93));
    layer0_outputs(7888) <= not((inputs(227)) xor (inputs(129)));
    layer0_outputs(7889) <= not((inputs(131)) xor (inputs(104)));
    layer0_outputs(7890) <= not(inputs(34));
    layer0_outputs(7891) <= inputs(165);
    layer0_outputs(7892) <= inputs(39);
    layer0_outputs(7893) <= inputs(165);
    layer0_outputs(7894) <= not(inputs(101));
    layer0_outputs(7895) <= not(inputs(124)) or (inputs(177));
    layer0_outputs(7896) <= (inputs(167)) or (inputs(194));
    layer0_outputs(7897) <= (inputs(197)) or (inputs(207));
    layer0_outputs(7898) <= not(inputs(200));
    layer0_outputs(7899) <= (inputs(222)) or (inputs(209));
    layer0_outputs(7900) <= (inputs(154)) and (inputs(233));
    layer0_outputs(7901) <= (inputs(61)) or (inputs(67));
    layer0_outputs(7902) <= not((inputs(200)) xor (inputs(184)));
    layer0_outputs(7903) <= not((inputs(34)) or (inputs(117)));
    layer0_outputs(7904) <= inputs(197);
    layer0_outputs(7905) <= not(inputs(149)) or (inputs(231));
    layer0_outputs(7906) <= not((inputs(52)) or (inputs(122)));
    layer0_outputs(7907) <= not(inputs(231)) or (inputs(44));
    layer0_outputs(7908) <= (inputs(94)) xor (inputs(226));
    layer0_outputs(7909) <= not(inputs(149));
    layer0_outputs(7910) <= not(inputs(94)) or (inputs(236));
    layer0_outputs(7911) <= (inputs(242)) or (inputs(139));
    layer0_outputs(7912) <= not((inputs(78)) xor (inputs(85)));
    layer0_outputs(7913) <= not((inputs(151)) xor (inputs(206)));
    layer0_outputs(7914) <= (inputs(173)) xor (inputs(255));
    layer0_outputs(7915) <= (inputs(75)) or (inputs(155));
    layer0_outputs(7916) <= not(inputs(105)) or (inputs(237));
    layer0_outputs(7917) <= not(inputs(173)) or (inputs(129));
    layer0_outputs(7918) <= not((inputs(161)) or (inputs(214)));
    layer0_outputs(7919) <= not(inputs(107));
    layer0_outputs(7920) <= (inputs(71)) or (inputs(50));
    layer0_outputs(7921) <= not((inputs(107)) and (inputs(16)));
    layer0_outputs(7922) <= not(inputs(42));
    layer0_outputs(7923) <= not((inputs(233)) xor (inputs(90)));
    layer0_outputs(7924) <= '1';
    layer0_outputs(7925) <= inputs(60);
    layer0_outputs(7926) <= (inputs(139)) xor (inputs(102));
    layer0_outputs(7927) <= (inputs(22)) and not (inputs(3));
    layer0_outputs(7928) <= (inputs(70)) xor (inputs(210));
    layer0_outputs(7929) <= not(inputs(103));
    layer0_outputs(7930) <= '0';
    layer0_outputs(7931) <= not(inputs(118));
    layer0_outputs(7932) <= (inputs(122)) xor (inputs(154));
    layer0_outputs(7933) <= not((inputs(52)) or (inputs(146)));
    layer0_outputs(7934) <= not((inputs(210)) or (inputs(93)));
    layer0_outputs(7935) <= (inputs(30)) and not (inputs(176));
    layer0_outputs(7936) <= (inputs(37)) xor (inputs(54));
    layer0_outputs(7937) <= (inputs(21)) xor (inputs(152));
    layer0_outputs(7938) <= not((inputs(224)) and (inputs(240)));
    layer0_outputs(7939) <= (inputs(138)) and not (inputs(188));
    layer0_outputs(7940) <= not(inputs(41));
    layer0_outputs(7941) <= (inputs(27)) and not (inputs(222));
    layer0_outputs(7942) <= inputs(136);
    layer0_outputs(7943) <= '0';
    layer0_outputs(7944) <= (inputs(101)) and not (inputs(242));
    layer0_outputs(7945) <= inputs(124);
    layer0_outputs(7946) <= not(inputs(43));
    layer0_outputs(7947) <= not(inputs(47)) or (inputs(91));
    layer0_outputs(7948) <= (inputs(11)) or (inputs(189));
    layer0_outputs(7949) <= not((inputs(20)) xor (inputs(177)));
    layer0_outputs(7950) <= (inputs(238)) xor (inputs(235));
    layer0_outputs(7951) <= (inputs(18)) and (inputs(241));
    layer0_outputs(7952) <= '0';
    layer0_outputs(7953) <= (inputs(245)) and (inputs(66));
    layer0_outputs(7954) <= not((inputs(93)) xor (inputs(248)));
    layer0_outputs(7955) <= not((inputs(66)) or (inputs(67)));
    layer0_outputs(7956) <= not(inputs(58)) or (inputs(218));
    layer0_outputs(7957) <= '0';
    layer0_outputs(7958) <= not(inputs(29));
    layer0_outputs(7959) <= not(inputs(232)) or (inputs(249));
    layer0_outputs(7960) <= (inputs(178)) and not (inputs(4));
    layer0_outputs(7961) <= not((inputs(198)) or (inputs(97)));
    layer0_outputs(7962) <= (inputs(107)) or (inputs(84));
    layer0_outputs(7963) <= (inputs(111)) and (inputs(14));
    layer0_outputs(7964) <= not((inputs(147)) or (inputs(235)));
    layer0_outputs(7965) <= not(inputs(170));
    layer0_outputs(7966) <= not(inputs(43)) or (inputs(155));
    layer0_outputs(7967) <= (inputs(157)) and not (inputs(0));
    layer0_outputs(7968) <= not(inputs(124)) or (inputs(176));
    layer0_outputs(7969) <= not(inputs(252)) or (inputs(55));
    layer0_outputs(7970) <= (inputs(227)) and (inputs(115));
    layer0_outputs(7971) <= (inputs(78)) or (inputs(53));
    layer0_outputs(7972) <= (inputs(115)) and not (inputs(98));
    layer0_outputs(7973) <= not(inputs(88));
    layer0_outputs(7974) <= inputs(201);
    layer0_outputs(7975) <= inputs(118);
    layer0_outputs(7976) <= (inputs(162)) and (inputs(171));
    layer0_outputs(7977) <= not(inputs(213)) or (inputs(195));
    layer0_outputs(7978) <= not((inputs(217)) xor (inputs(251)));
    layer0_outputs(7979) <= (inputs(9)) xor (inputs(172));
    layer0_outputs(7980) <= not(inputs(142));
    layer0_outputs(7981) <= (inputs(16)) and not (inputs(46));
    layer0_outputs(7982) <= inputs(229);
    layer0_outputs(7983) <= inputs(17);
    layer0_outputs(7984) <= (inputs(15)) or (inputs(46));
    layer0_outputs(7985) <= (inputs(173)) xor (inputs(63));
    layer0_outputs(7986) <= (inputs(194)) or (inputs(64));
    layer0_outputs(7987) <= inputs(58);
    layer0_outputs(7988) <= (inputs(68)) and not (inputs(131));
    layer0_outputs(7989) <= not((inputs(23)) or (inputs(62)));
    layer0_outputs(7990) <= not((inputs(27)) and (inputs(80)));
    layer0_outputs(7991) <= not(inputs(252));
    layer0_outputs(7992) <= not(inputs(108)) or (inputs(65));
    layer0_outputs(7993) <= (inputs(78)) and (inputs(71));
    layer0_outputs(7994) <= not((inputs(202)) or (inputs(19)));
    layer0_outputs(7995) <= '1';
    layer0_outputs(7996) <= inputs(186);
    layer0_outputs(7997) <= (inputs(69)) and not (inputs(96));
    layer0_outputs(7998) <= inputs(174);
    layer0_outputs(7999) <= not((inputs(27)) xor (inputs(28)));
    layer0_outputs(8000) <= inputs(117);
    layer0_outputs(8001) <= not((inputs(66)) or (inputs(147)));
    layer0_outputs(8002) <= (inputs(66)) and not (inputs(97));
    layer0_outputs(8003) <= not(inputs(151));
    layer0_outputs(8004) <= (inputs(117)) or (inputs(60));
    layer0_outputs(8005) <= not(inputs(62));
    layer0_outputs(8006) <= not(inputs(182));
    layer0_outputs(8007) <= (inputs(15)) and (inputs(205));
    layer0_outputs(8008) <= inputs(101);
    layer0_outputs(8009) <= (inputs(24)) xor (inputs(13));
    layer0_outputs(8010) <= not(inputs(183));
    layer0_outputs(8011) <= not(inputs(250)) or (inputs(126));
    layer0_outputs(8012) <= not((inputs(219)) xor (inputs(190)));
    layer0_outputs(8013) <= not(inputs(15)) or (inputs(131));
    layer0_outputs(8014) <= (inputs(55)) or (inputs(30));
    layer0_outputs(8015) <= not(inputs(106)) or (inputs(250));
    layer0_outputs(8016) <= (inputs(135)) or (inputs(246));
    layer0_outputs(8017) <= (inputs(45)) and not (inputs(7));
    layer0_outputs(8018) <= not((inputs(51)) and (inputs(207)));
    layer0_outputs(8019) <= not(inputs(189));
    layer0_outputs(8020) <= (inputs(44)) and not (inputs(50));
    layer0_outputs(8021) <= (inputs(137)) and not (inputs(62));
    layer0_outputs(8022) <= not(inputs(80)) or (inputs(28));
    layer0_outputs(8023) <= inputs(118);
    layer0_outputs(8024) <= (inputs(83)) xor (inputs(207));
    layer0_outputs(8025) <= inputs(88);
    layer0_outputs(8026) <= not(inputs(113));
    layer0_outputs(8027) <= not((inputs(29)) or (inputs(130)));
    layer0_outputs(8028) <= (inputs(108)) and not (inputs(134));
    layer0_outputs(8029) <= inputs(102);
    layer0_outputs(8030) <= inputs(15);
    layer0_outputs(8031) <= (inputs(89)) and not (inputs(117));
    layer0_outputs(8032) <= inputs(89);
    layer0_outputs(8033) <= (inputs(30)) xor (inputs(82));
    layer0_outputs(8034) <= not((inputs(221)) and (inputs(46)));
    layer0_outputs(8035) <= inputs(84);
    layer0_outputs(8036) <= (inputs(23)) xor (inputs(3));
    layer0_outputs(8037) <= not((inputs(102)) and (inputs(240)));
    layer0_outputs(8038) <= '1';
    layer0_outputs(8039) <= not((inputs(23)) xor (inputs(119)));
    layer0_outputs(8040) <= (inputs(97)) xor (inputs(142));
    layer0_outputs(8041) <= not(inputs(199)) or (inputs(197));
    layer0_outputs(8042) <= not((inputs(110)) or (inputs(63)));
    layer0_outputs(8043) <= not((inputs(59)) or (inputs(130)));
    layer0_outputs(8044) <= not(inputs(228));
    layer0_outputs(8045) <= not((inputs(120)) xor (inputs(135)));
    layer0_outputs(8046) <= (inputs(222)) and not (inputs(79));
    layer0_outputs(8047) <= '0';
    layer0_outputs(8048) <= not(inputs(1));
    layer0_outputs(8049) <= (inputs(62)) or (inputs(196));
    layer0_outputs(8050) <= (inputs(178)) xor (inputs(11));
    layer0_outputs(8051) <= (inputs(220)) xor (inputs(207));
    layer0_outputs(8052) <= (inputs(101)) and not (inputs(6));
    layer0_outputs(8053) <= not((inputs(117)) or (inputs(126)));
    layer0_outputs(8054) <= not(inputs(231)) or (inputs(34));
    layer0_outputs(8055) <= (inputs(80)) xor (inputs(183));
    layer0_outputs(8056) <= not(inputs(71)) or (inputs(170));
    layer0_outputs(8057) <= '1';
    layer0_outputs(8058) <= (inputs(92)) and not (inputs(175));
    layer0_outputs(8059) <= (inputs(104)) xor (inputs(239));
    layer0_outputs(8060) <= not(inputs(136));
    layer0_outputs(8061) <= not(inputs(152)) or (inputs(77));
    layer0_outputs(8062) <= not(inputs(58));
    layer0_outputs(8063) <= not(inputs(5));
    layer0_outputs(8064) <= inputs(215);
    layer0_outputs(8065) <= (inputs(72)) and not (inputs(195));
    layer0_outputs(8066) <= (inputs(44)) or (inputs(61));
    layer0_outputs(8067) <= (inputs(251)) and (inputs(226));
    layer0_outputs(8068) <= inputs(76);
    layer0_outputs(8069) <= (inputs(38)) xor (inputs(6));
    layer0_outputs(8070) <= (inputs(198)) and not (inputs(14));
    layer0_outputs(8071) <= not(inputs(145)) or (inputs(248));
    layer0_outputs(8072) <= not(inputs(184)) or (inputs(73));
    layer0_outputs(8073) <= (inputs(23)) or (inputs(168));
    layer0_outputs(8074) <= inputs(190);
    layer0_outputs(8075) <= not(inputs(123));
    layer0_outputs(8076) <= not(inputs(15)) or (inputs(156));
    layer0_outputs(8077) <= '0';
    layer0_outputs(8078) <= (inputs(85)) and not (inputs(128));
    layer0_outputs(8079) <= inputs(104);
    layer0_outputs(8080) <= (inputs(225)) and not (inputs(61));
    layer0_outputs(8081) <= not(inputs(167)) or (inputs(170));
    layer0_outputs(8082) <= not(inputs(105));
    layer0_outputs(8083) <= not((inputs(158)) xor (inputs(139)));
    layer0_outputs(8084) <= not(inputs(109)) or (inputs(14));
    layer0_outputs(8085) <= not(inputs(13));
    layer0_outputs(8086) <= (inputs(86)) xor (inputs(85));
    layer0_outputs(8087) <= (inputs(165)) and not (inputs(9));
    layer0_outputs(8088) <= not((inputs(68)) or (inputs(181)));
    layer0_outputs(8089) <= (inputs(241)) xor (inputs(54));
    layer0_outputs(8090) <= inputs(38);
    layer0_outputs(8091) <= '0';
    layer0_outputs(8092) <= (inputs(213)) and not (inputs(4));
    layer0_outputs(8093) <= not(inputs(96));
    layer0_outputs(8094) <= (inputs(92)) and (inputs(118));
    layer0_outputs(8095) <= (inputs(142)) or (inputs(235));
    layer0_outputs(8096) <= (inputs(197)) or (inputs(193));
    layer0_outputs(8097) <= not(inputs(135));
    layer0_outputs(8098) <= (inputs(168)) and not (inputs(104));
    layer0_outputs(8099) <= inputs(255);
    layer0_outputs(8100) <= inputs(106);
    layer0_outputs(8101) <= (inputs(238)) and not (inputs(127));
    layer0_outputs(8102) <= not((inputs(90)) xor (inputs(216)));
    layer0_outputs(8103) <= '0';
    layer0_outputs(8104) <= (inputs(196)) or (inputs(141));
    layer0_outputs(8105) <= not(inputs(174)) or (inputs(174));
    layer0_outputs(8106) <= not((inputs(63)) and (inputs(180)));
    layer0_outputs(8107) <= not(inputs(58));
    layer0_outputs(8108) <= not(inputs(77)) or (inputs(160));
    layer0_outputs(8109) <= '1';
    layer0_outputs(8110) <= not(inputs(144));
    layer0_outputs(8111) <= (inputs(113)) or (inputs(81));
    layer0_outputs(8112) <= inputs(157);
    layer0_outputs(8113) <= not(inputs(181)) or (inputs(247));
    layer0_outputs(8114) <= not(inputs(104));
    layer0_outputs(8115) <= (inputs(76)) or (inputs(244));
    layer0_outputs(8116) <= (inputs(117)) or (inputs(46));
    layer0_outputs(8117) <= inputs(242);
    layer0_outputs(8118) <= (inputs(138)) xor (inputs(18));
    layer0_outputs(8119) <= inputs(215);
    layer0_outputs(8120) <= (inputs(157)) or (inputs(124));
    layer0_outputs(8121) <= '1';
    layer0_outputs(8122) <= (inputs(59)) or (inputs(174));
    layer0_outputs(8123) <= not(inputs(43));
    layer0_outputs(8124) <= not(inputs(67)) or (inputs(177));
    layer0_outputs(8125) <= (inputs(87)) or (inputs(156));
    layer0_outputs(8126) <= (inputs(157)) or (inputs(206));
    layer0_outputs(8127) <= not((inputs(104)) or (inputs(31)));
    layer0_outputs(8128) <= (inputs(70)) and not (inputs(112));
    layer0_outputs(8129) <= inputs(232);
    layer0_outputs(8130) <= inputs(78);
    layer0_outputs(8131) <= (inputs(200)) and not (inputs(85));
    layer0_outputs(8132) <= '1';
    layer0_outputs(8133) <= not((inputs(206)) or (inputs(233)));
    layer0_outputs(8134) <= not((inputs(104)) or (inputs(107)));
    layer0_outputs(8135) <= not((inputs(71)) and (inputs(145)));
    layer0_outputs(8136) <= (inputs(156)) or (inputs(12));
    layer0_outputs(8137) <= (inputs(59)) or (inputs(12));
    layer0_outputs(8138) <= not(inputs(156)) or (inputs(127));
    layer0_outputs(8139) <= (inputs(153)) or (inputs(230));
    layer0_outputs(8140) <= not(inputs(250));
    layer0_outputs(8141) <= (inputs(52)) or (inputs(121));
    layer0_outputs(8142) <= not(inputs(154));
    layer0_outputs(8143) <= not((inputs(8)) or (inputs(104)));
    layer0_outputs(8144) <= (inputs(255)) xor (inputs(27));
    layer0_outputs(8145) <= not(inputs(184)) or (inputs(84));
    layer0_outputs(8146) <= (inputs(2)) xor (inputs(134));
    layer0_outputs(8147) <= not(inputs(7)) or (inputs(67));
    layer0_outputs(8148) <= inputs(142);
    layer0_outputs(8149) <= (inputs(249)) or (inputs(165));
    layer0_outputs(8150) <= (inputs(125)) and not (inputs(220));
    layer0_outputs(8151) <= not(inputs(58));
    layer0_outputs(8152) <= not((inputs(24)) xor (inputs(142)));
    layer0_outputs(8153) <= not(inputs(166)) or (inputs(63));
    layer0_outputs(8154) <= (inputs(64)) and not (inputs(3));
    layer0_outputs(8155) <= (inputs(69)) xor (inputs(6));
    layer0_outputs(8156) <= (inputs(70)) and not (inputs(117));
    layer0_outputs(8157) <= not(inputs(117));
    layer0_outputs(8158) <= not(inputs(0));
    layer0_outputs(8159) <= not((inputs(41)) or (inputs(6)));
    layer0_outputs(8160) <= (inputs(142)) and (inputs(133));
    layer0_outputs(8161) <= not((inputs(47)) xor (inputs(151)));
    layer0_outputs(8162) <= not(inputs(163)) or (inputs(216));
    layer0_outputs(8163) <= (inputs(35)) or (inputs(143));
    layer0_outputs(8164) <= (inputs(35)) and not (inputs(124));
    layer0_outputs(8165) <= not((inputs(200)) or (inputs(157)));
    layer0_outputs(8166) <= not(inputs(164));
    layer0_outputs(8167) <= inputs(85);
    layer0_outputs(8168) <= not(inputs(240)) or (inputs(177));
    layer0_outputs(8169) <= inputs(119);
    layer0_outputs(8170) <= not((inputs(123)) xor (inputs(17)));
    layer0_outputs(8171) <= (inputs(119)) or (inputs(100));
    layer0_outputs(8172) <= (inputs(241)) and not (inputs(110));
    layer0_outputs(8173) <= not(inputs(216)) or (inputs(160));
    layer0_outputs(8174) <= not((inputs(157)) xor (inputs(46)));
    layer0_outputs(8175) <= (inputs(87)) and not (inputs(28));
    layer0_outputs(8176) <= (inputs(54)) xor (inputs(56));
    layer0_outputs(8177) <= not(inputs(120)) or (inputs(49));
    layer0_outputs(8178) <= (inputs(242)) xor (inputs(48));
    layer0_outputs(8179) <= (inputs(185)) and (inputs(187));
    layer0_outputs(8180) <= not((inputs(130)) or (inputs(137)));
    layer0_outputs(8181) <= inputs(200);
    layer0_outputs(8182) <= '0';
    layer0_outputs(8183) <= (inputs(8)) or (inputs(172));
    layer0_outputs(8184) <= (inputs(74)) and not (inputs(32));
    layer0_outputs(8185) <= (inputs(202)) xor (inputs(2));
    layer0_outputs(8186) <= not(inputs(184)) or (inputs(129));
    layer0_outputs(8187) <= (inputs(242)) xor (inputs(139));
    layer0_outputs(8188) <= not(inputs(240));
    layer0_outputs(8189) <= not((inputs(78)) or (inputs(203)));
    layer0_outputs(8190) <= (inputs(15)) and not (inputs(203));
    layer0_outputs(8191) <= '1';
    layer0_outputs(8192) <= (inputs(124)) xor (inputs(6));
    layer0_outputs(8193) <= (inputs(118)) or (inputs(94));
    layer0_outputs(8194) <= '0';
    layer0_outputs(8195) <= (inputs(126)) and (inputs(10));
    layer0_outputs(8196) <= (inputs(166)) xor (inputs(28));
    layer0_outputs(8197) <= not(inputs(24)) or (inputs(254));
    layer0_outputs(8198) <= (inputs(128)) xor (inputs(130));
    layer0_outputs(8199) <= (inputs(56)) xor (inputs(182));
    layer0_outputs(8200) <= inputs(82);
    layer0_outputs(8201) <= not((inputs(123)) or (inputs(107)));
    layer0_outputs(8202) <= (inputs(227)) or (inputs(51));
    layer0_outputs(8203) <= (inputs(38)) and not (inputs(204));
    layer0_outputs(8204) <= inputs(187);
    layer0_outputs(8205) <= inputs(36);
    layer0_outputs(8206) <= not(inputs(122)) or (inputs(60));
    layer0_outputs(8207) <= (inputs(218)) xor (inputs(209));
    layer0_outputs(8208) <= inputs(181);
    layer0_outputs(8209) <= not((inputs(92)) or (inputs(50)));
    layer0_outputs(8210) <= (inputs(86)) or (inputs(31));
    layer0_outputs(8211) <= not(inputs(201));
    layer0_outputs(8212) <= not(inputs(40)) or (inputs(195));
    layer0_outputs(8213) <= not(inputs(122)) or (inputs(97));
    layer0_outputs(8214) <= (inputs(123)) and not (inputs(216));
    layer0_outputs(8215) <= not((inputs(0)) or (inputs(231)));
    layer0_outputs(8216) <= not((inputs(15)) or (inputs(77)));
    layer0_outputs(8217) <= not(inputs(159)) or (inputs(208));
    layer0_outputs(8218) <= not((inputs(29)) and (inputs(50)));
    layer0_outputs(8219) <= (inputs(174)) and (inputs(146));
    layer0_outputs(8220) <= not(inputs(170)) or (inputs(252));
    layer0_outputs(8221) <= (inputs(228)) and not (inputs(228));
    layer0_outputs(8222) <= not(inputs(60)) or (inputs(174));
    layer0_outputs(8223) <= (inputs(78)) and not (inputs(208));
    layer0_outputs(8224) <= (inputs(234)) and (inputs(52));
    layer0_outputs(8225) <= not(inputs(164));
    layer0_outputs(8226) <= inputs(64);
    layer0_outputs(8227) <= (inputs(45)) xor (inputs(85));
    layer0_outputs(8228) <= not(inputs(201)) or (inputs(8));
    layer0_outputs(8229) <= (inputs(91)) and not (inputs(247));
    layer0_outputs(8230) <= not(inputs(70));
    layer0_outputs(8231) <= (inputs(86)) and not (inputs(30));
    layer0_outputs(8232) <= not((inputs(138)) or (inputs(154)));
    layer0_outputs(8233) <= inputs(27);
    layer0_outputs(8234) <= (inputs(186)) and not (inputs(84));
    layer0_outputs(8235) <= (inputs(53)) or (inputs(176));
    layer0_outputs(8236) <= (inputs(34)) xor (inputs(115));
    layer0_outputs(8237) <= inputs(179);
    layer0_outputs(8238) <= not((inputs(89)) or (inputs(95)));
    layer0_outputs(8239) <= (inputs(112)) or (inputs(59));
    layer0_outputs(8240) <= not(inputs(198)) or (inputs(95));
    layer0_outputs(8241) <= not(inputs(135)) or (inputs(64));
    layer0_outputs(8242) <= inputs(106);
    layer0_outputs(8243) <= not((inputs(108)) or (inputs(224)));
    layer0_outputs(8244) <= (inputs(211)) and (inputs(12));
    layer0_outputs(8245) <= not(inputs(103));
    layer0_outputs(8246) <= not(inputs(29)) or (inputs(156));
    layer0_outputs(8247) <= (inputs(82)) xor (inputs(23));
    layer0_outputs(8248) <= (inputs(25)) or (inputs(185));
    layer0_outputs(8249) <= (inputs(133)) and not (inputs(97));
    layer0_outputs(8250) <= (inputs(112)) xor (inputs(83));
    layer0_outputs(8251) <= not(inputs(151));
    layer0_outputs(8252) <= not(inputs(79));
    layer0_outputs(8253) <= (inputs(239)) and (inputs(154));
    layer0_outputs(8254) <= (inputs(126)) or (inputs(170));
    layer0_outputs(8255) <= (inputs(231)) or (inputs(29));
    layer0_outputs(8256) <= not((inputs(83)) xor (inputs(111)));
    layer0_outputs(8257) <= (inputs(231)) xor (inputs(27));
    layer0_outputs(8258) <= (inputs(20)) or (inputs(93));
    layer0_outputs(8259) <= '1';
    layer0_outputs(8260) <= not(inputs(86)) or (inputs(173));
    layer0_outputs(8261) <= not(inputs(21));
    layer0_outputs(8262) <= inputs(199);
    layer0_outputs(8263) <= not(inputs(72));
    layer0_outputs(8264) <= (inputs(161)) xor (inputs(173));
    layer0_outputs(8265) <= not((inputs(244)) xor (inputs(228)));
    layer0_outputs(8266) <= (inputs(3)) or (inputs(179));
    layer0_outputs(8267) <= (inputs(141)) and not (inputs(143));
    layer0_outputs(8268) <= not((inputs(130)) xor (inputs(64)));
    layer0_outputs(8269) <= not((inputs(150)) xor (inputs(157)));
    layer0_outputs(8270) <= not((inputs(148)) xor (inputs(117)));
    layer0_outputs(8271) <= (inputs(101)) or (inputs(26));
    layer0_outputs(8272) <= inputs(121);
    layer0_outputs(8273) <= not(inputs(73));
    layer0_outputs(8274) <= '0';
    layer0_outputs(8275) <= (inputs(251)) or (inputs(162));
    layer0_outputs(8276) <= inputs(140);
    layer0_outputs(8277) <= not((inputs(202)) and (inputs(78)));
    layer0_outputs(8278) <= (inputs(208)) or (inputs(215));
    layer0_outputs(8279) <= inputs(7);
    layer0_outputs(8280) <= '0';
    layer0_outputs(8281) <= (inputs(146)) or (inputs(53));
    layer0_outputs(8282) <= (inputs(226)) or (inputs(172));
    layer0_outputs(8283) <= (inputs(110)) and not (inputs(127));
    layer0_outputs(8284) <= (inputs(84)) and not (inputs(125));
    layer0_outputs(8285) <= inputs(84);
    layer0_outputs(8286) <= not(inputs(95));
    layer0_outputs(8287) <= (inputs(159)) or (inputs(139));
    layer0_outputs(8288) <= not(inputs(47));
    layer0_outputs(8289) <= not(inputs(139));
    layer0_outputs(8290) <= (inputs(197)) and not (inputs(131));
    layer0_outputs(8291) <= (inputs(110)) and not (inputs(240));
    layer0_outputs(8292) <= inputs(156);
    layer0_outputs(8293) <= not((inputs(14)) xor (inputs(168)));
    layer0_outputs(8294) <= inputs(185);
    layer0_outputs(8295) <= not((inputs(238)) xor (inputs(238)));
    layer0_outputs(8296) <= (inputs(223)) or (inputs(155));
    layer0_outputs(8297) <= not((inputs(181)) xor (inputs(166)));
    layer0_outputs(8298) <= (inputs(54)) or (inputs(192));
    layer0_outputs(8299) <= inputs(220);
    layer0_outputs(8300) <= (inputs(167)) and not (inputs(111));
    layer0_outputs(8301) <= not(inputs(167));
    layer0_outputs(8302) <= (inputs(232)) and (inputs(207));
    layer0_outputs(8303) <= not((inputs(81)) or (inputs(117)));
    layer0_outputs(8304) <= not((inputs(194)) or (inputs(81)));
    layer0_outputs(8305) <= not((inputs(27)) or (inputs(189)));
    layer0_outputs(8306) <= not(inputs(60));
    layer0_outputs(8307) <= not(inputs(182));
    layer0_outputs(8308) <= inputs(55);
    layer0_outputs(8309) <= not(inputs(153));
    layer0_outputs(8310) <= (inputs(208)) or (inputs(24));
    layer0_outputs(8311) <= (inputs(248)) and (inputs(28));
    layer0_outputs(8312) <= not(inputs(29));
    layer0_outputs(8313) <= not(inputs(203)) or (inputs(61));
    layer0_outputs(8314) <= not((inputs(235)) or (inputs(123)));
    layer0_outputs(8315) <= not(inputs(103)) or (inputs(96));
    layer0_outputs(8316) <= '0';
    layer0_outputs(8317) <= not(inputs(136));
    layer0_outputs(8318) <= not((inputs(4)) or (inputs(109)));
    layer0_outputs(8319) <= (inputs(222)) and not (inputs(3));
    layer0_outputs(8320) <= not(inputs(21)) or (inputs(222));
    layer0_outputs(8321) <= not(inputs(26));
    layer0_outputs(8322) <= not(inputs(147));
    layer0_outputs(8323) <= (inputs(157)) and (inputs(129));
    layer0_outputs(8324) <= not((inputs(129)) or (inputs(196)));
    layer0_outputs(8325) <= not((inputs(164)) or (inputs(88)));
    layer0_outputs(8326) <= (inputs(47)) and (inputs(108));
    layer0_outputs(8327) <= not(inputs(215)) or (inputs(226));
    layer0_outputs(8328) <= (inputs(151)) or (inputs(116));
    layer0_outputs(8329) <= (inputs(76)) and (inputs(76));
    layer0_outputs(8330) <= (inputs(69)) xor (inputs(187));
    layer0_outputs(8331) <= not((inputs(140)) xor (inputs(209)));
    layer0_outputs(8332) <= inputs(200);
    layer0_outputs(8333) <= not(inputs(172)) or (inputs(108));
    layer0_outputs(8334) <= (inputs(190)) xor (inputs(197));
    layer0_outputs(8335) <= not(inputs(230)) or (inputs(1));
    layer0_outputs(8336) <= not(inputs(124));
    layer0_outputs(8337) <= '1';
    layer0_outputs(8338) <= (inputs(237)) or (inputs(6));
    layer0_outputs(8339) <= not(inputs(86));
    layer0_outputs(8340) <= inputs(106);
    layer0_outputs(8341) <= (inputs(244)) xor (inputs(198));
    layer0_outputs(8342) <= not(inputs(137)) or (inputs(99));
    layer0_outputs(8343) <= (inputs(46)) or (inputs(48));
    layer0_outputs(8344) <= (inputs(48)) and not (inputs(114));
    layer0_outputs(8345) <= not(inputs(73)) or (inputs(200));
    layer0_outputs(8346) <= inputs(105);
    layer0_outputs(8347) <= (inputs(151)) and not (inputs(178));
    layer0_outputs(8348) <= not(inputs(133));
    layer0_outputs(8349) <= not(inputs(236));
    layer0_outputs(8350) <= (inputs(173)) and not (inputs(22));
    layer0_outputs(8351) <= not(inputs(119));
    layer0_outputs(8352) <= inputs(66);
    layer0_outputs(8353) <= not((inputs(109)) or (inputs(253)));
    layer0_outputs(8354) <= not(inputs(148));
    layer0_outputs(8355) <= not((inputs(209)) xor (inputs(182)));
    layer0_outputs(8356) <= not(inputs(154)) or (inputs(206));
    layer0_outputs(8357) <= (inputs(78)) xor (inputs(3));
    layer0_outputs(8358) <= not((inputs(254)) and (inputs(240)));
    layer0_outputs(8359) <= not(inputs(240)) or (inputs(217));
    layer0_outputs(8360) <= not((inputs(45)) and (inputs(8)));
    layer0_outputs(8361) <= not(inputs(165)) or (inputs(81));
    layer0_outputs(8362) <= (inputs(14)) and (inputs(162));
    layer0_outputs(8363) <= not((inputs(207)) xor (inputs(213)));
    layer0_outputs(8364) <= (inputs(172)) xor (inputs(79));
    layer0_outputs(8365) <= '1';
    layer0_outputs(8366) <= not(inputs(6)) or (inputs(121));
    layer0_outputs(8367) <= (inputs(137)) and not (inputs(69));
    layer0_outputs(8368) <= not(inputs(142));
    layer0_outputs(8369) <= not((inputs(215)) and (inputs(102)));
    layer0_outputs(8370) <= inputs(2);
    layer0_outputs(8371) <= not(inputs(197));
    layer0_outputs(8372) <= not((inputs(231)) or (inputs(123)));
    layer0_outputs(8373) <= inputs(163);
    layer0_outputs(8374) <= not((inputs(248)) or (inputs(138)));
    layer0_outputs(8375) <= inputs(77);
    layer0_outputs(8376) <= '0';
    layer0_outputs(8377) <= not(inputs(106));
    layer0_outputs(8378) <= (inputs(101)) and not (inputs(40));
    layer0_outputs(8379) <= (inputs(1)) and (inputs(214));
    layer0_outputs(8380) <= not(inputs(59));
    layer0_outputs(8381) <= (inputs(37)) xor (inputs(157));
    layer0_outputs(8382) <= (inputs(142)) or (inputs(103));
    layer0_outputs(8383) <= not((inputs(231)) xor (inputs(26)));
    layer0_outputs(8384) <= (inputs(138)) and not (inputs(194));
    layer0_outputs(8385) <= not((inputs(40)) or (inputs(197)));
    layer0_outputs(8386) <= not((inputs(222)) or (inputs(243)));
    layer0_outputs(8387) <= inputs(204);
    layer0_outputs(8388) <= (inputs(170)) and not (inputs(25));
    layer0_outputs(8389) <= (inputs(216)) and not (inputs(229));
    layer0_outputs(8390) <= not(inputs(223));
    layer0_outputs(8391) <= not(inputs(57));
    layer0_outputs(8392) <= not((inputs(32)) xor (inputs(31)));
    layer0_outputs(8393) <= not(inputs(116)) or (inputs(144));
    layer0_outputs(8394) <= not(inputs(54)) or (inputs(176));
    layer0_outputs(8395) <= not((inputs(225)) xor (inputs(38)));
    layer0_outputs(8396) <= (inputs(95)) xor (inputs(26));
    layer0_outputs(8397) <= (inputs(154)) and not (inputs(208));
    layer0_outputs(8398) <= inputs(56);
    layer0_outputs(8399) <= not((inputs(127)) xor (inputs(86)));
    layer0_outputs(8400) <= not((inputs(23)) or (inputs(83)));
    layer0_outputs(8401) <= (inputs(143)) or (inputs(154));
    layer0_outputs(8402) <= inputs(29);
    layer0_outputs(8403) <= not((inputs(54)) xor (inputs(175)));
    layer0_outputs(8404) <= (inputs(237)) xor (inputs(209));
    layer0_outputs(8405) <= (inputs(191)) xor (inputs(36));
    layer0_outputs(8406) <= inputs(165);
    layer0_outputs(8407) <= not((inputs(79)) or (inputs(83)));
    layer0_outputs(8408) <= '1';
    layer0_outputs(8409) <= not(inputs(101));
    layer0_outputs(8410) <= (inputs(44)) and not (inputs(174));
    layer0_outputs(8411) <= not(inputs(200));
    layer0_outputs(8412) <= not(inputs(140)) or (inputs(122));
    layer0_outputs(8413) <= not((inputs(210)) or (inputs(35)));
    layer0_outputs(8414) <= inputs(148);
    layer0_outputs(8415) <= not((inputs(108)) or (inputs(34)));
    layer0_outputs(8416) <= (inputs(176)) and not (inputs(146));
    layer0_outputs(8417) <= not((inputs(205)) xor (inputs(191)));
    layer0_outputs(8418) <= (inputs(190)) and (inputs(161));
    layer0_outputs(8419) <= inputs(204);
    layer0_outputs(8420) <= (inputs(20)) and (inputs(6));
    layer0_outputs(8421) <= (inputs(133)) or (inputs(235));
    layer0_outputs(8422) <= (inputs(68)) and not (inputs(204));
    layer0_outputs(8423) <= (inputs(233)) xor (inputs(189));
    layer0_outputs(8424) <= not(inputs(53)) or (inputs(207));
    layer0_outputs(8425) <= not(inputs(214));
    layer0_outputs(8426) <= not(inputs(251)) or (inputs(86));
    layer0_outputs(8427) <= inputs(144);
    layer0_outputs(8428) <= not((inputs(172)) and (inputs(243)));
    layer0_outputs(8429) <= inputs(3);
    layer0_outputs(8430) <= (inputs(94)) or (inputs(123));
    layer0_outputs(8431) <= not(inputs(171));
    layer0_outputs(8432) <= not(inputs(73)) or (inputs(204));
    layer0_outputs(8433) <= (inputs(45)) or (inputs(63));
    layer0_outputs(8434) <= not((inputs(76)) xor (inputs(124)));
    layer0_outputs(8435) <= inputs(186);
    layer0_outputs(8436) <= not(inputs(118));
    layer0_outputs(8437) <= '0';
    layer0_outputs(8438) <= '0';
    layer0_outputs(8439) <= inputs(87);
    layer0_outputs(8440) <= (inputs(56)) or (inputs(232));
    layer0_outputs(8441) <= (inputs(101)) or (inputs(19));
    layer0_outputs(8442) <= not((inputs(178)) xor (inputs(141)));
    layer0_outputs(8443) <= (inputs(30)) and (inputs(177));
    layer0_outputs(8444) <= (inputs(236)) xor (inputs(143));
    layer0_outputs(8445) <= (inputs(206)) or (inputs(77));
    layer0_outputs(8446) <= not(inputs(61)) or (inputs(224));
    layer0_outputs(8447) <= not(inputs(188));
    layer0_outputs(8448) <= (inputs(86)) and (inputs(84));
    layer0_outputs(8449) <= not((inputs(141)) or (inputs(42)));
    layer0_outputs(8450) <= not((inputs(244)) or (inputs(81)));
    layer0_outputs(8451) <= (inputs(165)) and not (inputs(89));
    layer0_outputs(8452) <= (inputs(100)) or (inputs(168));
    layer0_outputs(8453) <= not(inputs(212));
    layer0_outputs(8454) <= inputs(11);
    layer0_outputs(8455) <= inputs(169);
    layer0_outputs(8456) <= (inputs(101)) or (inputs(113));
    layer0_outputs(8457) <= (inputs(30)) xor (inputs(222));
    layer0_outputs(8458) <= inputs(135);
    layer0_outputs(8459) <= (inputs(247)) and not (inputs(48));
    layer0_outputs(8460) <= (inputs(236)) and not (inputs(255));
    layer0_outputs(8461) <= inputs(117);
    layer0_outputs(8462) <= (inputs(127)) or (inputs(180));
    layer0_outputs(8463) <= inputs(242);
    layer0_outputs(8464) <= not(inputs(185));
    layer0_outputs(8465) <= not(inputs(72)) or (inputs(205));
    layer0_outputs(8466) <= inputs(179);
    layer0_outputs(8467) <= inputs(252);
    layer0_outputs(8468) <= not(inputs(56)) or (inputs(175));
    layer0_outputs(8469) <= (inputs(140)) and not (inputs(82));
    layer0_outputs(8470) <= (inputs(105)) and not (inputs(84));
    layer0_outputs(8471) <= inputs(99);
    layer0_outputs(8472) <= inputs(120);
    layer0_outputs(8473) <= (inputs(185)) xor (inputs(244));
    layer0_outputs(8474) <= not((inputs(254)) xor (inputs(164)));
    layer0_outputs(8475) <= not((inputs(188)) xor (inputs(122)));
    layer0_outputs(8476) <= not((inputs(218)) xor (inputs(231)));
    layer0_outputs(8477) <= not((inputs(100)) or (inputs(122)));
    layer0_outputs(8478) <= not(inputs(189)) or (inputs(24));
    layer0_outputs(8479) <= not(inputs(137));
    layer0_outputs(8480) <= (inputs(119)) and not (inputs(131));
    layer0_outputs(8481) <= (inputs(108)) or (inputs(157));
    layer0_outputs(8482) <= not((inputs(142)) or (inputs(157)));
    layer0_outputs(8483) <= inputs(117);
    layer0_outputs(8484) <= not((inputs(86)) or (inputs(125)));
    layer0_outputs(8485) <= '1';
    layer0_outputs(8486) <= '0';
    layer0_outputs(8487) <= inputs(56);
    layer0_outputs(8488) <= (inputs(109)) or (inputs(40));
    layer0_outputs(8489) <= not((inputs(172)) or (inputs(163)));
    layer0_outputs(8490) <= (inputs(191)) and not (inputs(107));
    layer0_outputs(8491) <= not((inputs(72)) or (inputs(64)));
    layer0_outputs(8492) <= not((inputs(102)) xor (inputs(103)));
    layer0_outputs(8493) <= (inputs(13)) and not (inputs(13));
    layer0_outputs(8494) <= not((inputs(63)) or (inputs(161)));
    layer0_outputs(8495) <= inputs(102);
    layer0_outputs(8496) <= (inputs(20)) and not (inputs(62));
    layer0_outputs(8497) <= not(inputs(142));
    layer0_outputs(8498) <= not(inputs(138));
    layer0_outputs(8499) <= not(inputs(73));
    layer0_outputs(8500) <= not(inputs(101)) or (inputs(179));
    layer0_outputs(8501) <= inputs(44);
    layer0_outputs(8502) <= not(inputs(4));
    layer0_outputs(8503) <= not((inputs(191)) or (inputs(101)));
    layer0_outputs(8504) <= (inputs(245)) and not (inputs(5));
    layer0_outputs(8505) <= not((inputs(86)) or (inputs(83)));
    layer0_outputs(8506) <= (inputs(153)) or (inputs(152));
    layer0_outputs(8507) <= not(inputs(86));
    layer0_outputs(8508) <= not((inputs(234)) or (inputs(97)));
    layer0_outputs(8509) <= (inputs(169)) xor (inputs(140));
    layer0_outputs(8510) <= (inputs(227)) xor (inputs(54));
    layer0_outputs(8511) <= (inputs(59)) and not (inputs(0));
    layer0_outputs(8512) <= not(inputs(183));
    layer0_outputs(8513) <= not(inputs(72));
    layer0_outputs(8514) <= not((inputs(143)) and (inputs(110)));
    layer0_outputs(8515) <= not(inputs(190)) or (inputs(192));
    layer0_outputs(8516) <= not(inputs(114)) or (inputs(96));
    layer0_outputs(8517) <= (inputs(120)) and not (inputs(5));
    layer0_outputs(8518) <= inputs(172);
    layer0_outputs(8519) <= (inputs(94)) and (inputs(25));
    layer0_outputs(8520) <= inputs(178);
    layer0_outputs(8521) <= (inputs(172)) xor (inputs(123));
    layer0_outputs(8522) <= inputs(59);
    layer0_outputs(8523) <= not(inputs(149)) or (inputs(93));
    layer0_outputs(8524) <= inputs(142);
    layer0_outputs(8525) <= not((inputs(178)) xor (inputs(128)));
    layer0_outputs(8526) <= not((inputs(40)) xor (inputs(164)));
    layer0_outputs(8527) <= (inputs(124)) and not (inputs(240));
    layer0_outputs(8528) <= not(inputs(209)) or (inputs(251));
    layer0_outputs(8529) <= inputs(233);
    layer0_outputs(8530) <= not(inputs(136));
    layer0_outputs(8531) <= inputs(126);
    layer0_outputs(8532) <= inputs(162);
    layer0_outputs(8533) <= inputs(225);
    layer0_outputs(8534) <= (inputs(182)) xor (inputs(210));
    layer0_outputs(8535) <= not((inputs(237)) xor (inputs(201)));
    layer0_outputs(8536) <= not((inputs(214)) xor (inputs(46)));
    layer0_outputs(8537) <= inputs(162);
    layer0_outputs(8538) <= not((inputs(51)) xor (inputs(185)));
    layer0_outputs(8539) <= inputs(102);
    layer0_outputs(8540) <= (inputs(169)) xor (inputs(49));
    layer0_outputs(8541) <= '0';
    layer0_outputs(8542) <= not((inputs(212)) xor (inputs(155)));
    layer0_outputs(8543) <= (inputs(2)) xor (inputs(216));
    layer0_outputs(8544) <= not(inputs(163));
    layer0_outputs(8545) <= (inputs(112)) or (inputs(55));
    layer0_outputs(8546) <= '0';
    layer0_outputs(8547) <= (inputs(193)) or (inputs(98));
    layer0_outputs(8548) <= not((inputs(207)) xor (inputs(148)));
    layer0_outputs(8549) <= (inputs(121)) or (inputs(191));
    layer0_outputs(8550) <= (inputs(203)) and not (inputs(227));
    layer0_outputs(8551) <= not(inputs(5));
    layer0_outputs(8552) <= '1';
    layer0_outputs(8553) <= (inputs(168)) and not (inputs(92));
    layer0_outputs(8554) <= (inputs(222)) xor (inputs(171));
    layer0_outputs(8555) <= (inputs(25)) or (inputs(183));
    layer0_outputs(8556) <= (inputs(211)) and not (inputs(23));
    layer0_outputs(8557) <= not(inputs(179));
    layer0_outputs(8558) <= not((inputs(80)) xor (inputs(170)));
    layer0_outputs(8559) <= (inputs(159)) and (inputs(159));
    layer0_outputs(8560) <= '1';
    layer0_outputs(8561) <= inputs(120);
    layer0_outputs(8562) <= (inputs(192)) or (inputs(150));
    layer0_outputs(8563) <= not((inputs(231)) or (inputs(200)));
    layer0_outputs(8564) <= (inputs(47)) xor (inputs(105));
    layer0_outputs(8565) <= not(inputs(88)) or (inputs(98));
    layer0_outputs(8566) <= inputs(165);
    layer0_outputs(8567) <= (inputs(175)) or (inputs(81));
    layer0_outputs(8568) <= not(inputs(113)) or (inputs(238));
    layer0_outputs(8569) <= '0';
    layer0_outputs(8570) <= not((inputs(98)) and (inputs(1)));
    layer0_outputs(8571) <= (inputs(103)) and not (inputs(158));
    layer0_outputs(8572) <= inputs(174);
    layer0_outputs(8573) <= inputs(250);
    layer0_outputs(8574) <= not(inputs(156)) or (inputs(236));
    layer0_outputs(8575) <= not((inputs(176)) or (inputs(90)));
    layer0_outputs(8576) <= not(inputs(108)) or (inputs(125));
    layer0_outputs(8577) <= (inputs(241)) and (inputs(36));
    layer0_outputs(8578) <= inputs(106);
    layer0_outputs(8579) <= not((inputs(42)) or (inputs(155)));
    layer0_outputs(8580) <= not((inputs(184)) or (inputs(67)));
    layer0_outputs(8581) <= not(inputs(195));
    layer0_outputs(8582) <= (inputs(56)) and not (inputs(193));
    layer0_outputs(8583) <= (inputs(168)) and not (inputs(111));
    layer0_outputs(8584) <= not((inputs(91)) or (inputs(178)));
    layer0_outputs(8585) <= not((inputs(145)) xor (inputs(123)));
    layer0_outputs(8586) <= (inputs(125)) or (inputs(235));
    layer0_outputs(8587) <= not(inputs(50)) or (inputs(11));
    layer0_outputs(8588) <= (inputs(218)) xor (inputs(7));
    layer0_outputs(8589) <= not(inputs(27));
    layer0_outputs(8590) <= (inputs(69)) xor (inputs(155));
    layer0_outputs(8591) <= '1';
    layer0_outputs(8592) <= not(inputs(9));
    layer0_outputs(8593) <= (inputs(206)) or (inputs(253));
    layer0_outputs(8594) <= (inputs(1)) and (inputs(62));
    layer0_outputs(8595) <= not(inputs(221)) or (inputs(30));
    layer0_outputs(8596) <= inputs(204);
    layer0_outputs(8597) <= not(inputs(75)) or (inputs(126));
    layer0_outputs(8598) <= inputs(35);
    layer0_outputs(8599) <= inputs(147);
    layer0_outputs(8600) <= (inputs(116)) xor (inputs(17));
    layer0_outputs(8601) <= (inputs(157)) xor (inputs(39));
    layer0_outputs(8602) <= (inputs(103)) and not (inputs(148));
    layer0_outputs(8603) <= (inputs(105)) and not (inputs(251));
    layer0_outputs(8604) <= inputs(103);
    layer0_outputs(8605) <= not((inputs(184)) or (inputs(23)));
    layer0_outputs(8606) <= (inputs(87)) and not (inputs(177));
    layer0_outputs(8607) <= inputs(58);
    layer0_outputs(8608) <= not((inputs(98)) or (inputs(169)));
    layer0_outputs(8609) <= not(inputs(164)) or (inputs(236));
    layer0_outputs(8610) <= not(inputs(33));
    layer0_outputs(8611) <= not((inputs(233)) or (inputs(244)));
    layer0_outputs(8612) <= not(inputs(149));
    layer0_outputs(8613) <= (inputs(186)) and not (inputs(236));
    layer0_outputs(8614) <= not(inputs(102));
    layer0_outputs(8615) <= (inputs(74)) or (inputs(133));
    layer0_outputs(8616) <= inputs(196);
    layer0_outputs(8617) <= inputs(123);
    layer0_outputs(8618) <= (inputs(41)) xor (inputs(53));
    layer0_outputs(8619) <= (inputs(228)) and not (inputs(192));
    layer0_outputs(8620) <= (inputs(153)) and not (inputs(80));
    layer0_outputs(8621) <= (inputs(201)) xor (inputs(248));
    layer0_outputs(8622) <= (inputs(63)) xor (inputs(171));
    layer0_outputs(8623) <= not((inputs(171)) xor (inputs(239)));
    layer0_outputs(8624) <= not((inputs(250)) and (inputs(225)));
    layer0_outputs(8625) <= (inputs(191)) or (inputs(81));
    layer0_outputs(8626) <= not(inputs(71));
    layer0_outputs(8627) <= (inputs(13)) and not (inputs(50));
    layer0_outputs(8628) <= not((inputs(194)) or (inputs(105)));
    layer0_outputs(8629) <= not(inputs(105));
    layer0_outputs(8630) <= not((inputs(205)) xor (inputs(193)));
    layer0_outputs(8631) <= not(inputs(181)) or (inputs(228));
    layer0_outputs(8632) <= not(inputs(59));
    layer0_outputs(8633) <= inputs(26);
    layer0_outputs(8634) <= inputs(132);
    layer0_outputs(8635) <= not(inputs(187)) or (inputs(32));
    layer0_outputs(8636) <= (inputs(115)) and not (inputs(244));
    layer0_outputs(8637) <= not(inputs(18));
    layer0_outputs(8638) <= not((inputs(10)) or (inputs(157)));
    layer0_outputs(8639) <= not(inputs(166));
    layer0_outputs(8640) <= not(inputs(241)) or (inputs(65));
    layer0_outputs(8641) <= not((inputs(179)) xor (inputs(9)));
    layer0_outputs(8642) <= inputs(231);
    layer0_outputs(8643) <= inputs(180);
    layer0_outputs(8644) <= inputs(216);
    layer0_outputs(8645) <= (inputs(91)) or (inputs(143));
    layer0_outputs(8646) <= not((inputs(16)) xor (inputs(51)));
    layer0_outputs(8647) <= not((inputs(0)) xor (inputs(49)));
    layer0_outputs(8648) <= not((inputs(216)) or (inputs(241)));
    layer0_outputs(8649) <= (inputs(159)) and not (inputs(3));
    layer0_outputs(8650) <= not(inputs(16)) or (inputs(94));
    layer0_outputs(8651) <= (inputs(60)) or (inputs(178));
    layer0_outputs(8652) <= inputs(56);
    layer0_outputs(8653) <= not((inputs(92)) or (inputs(188)));
    layer0_outputs(8654) <= not((inputs(203)) or (inputs(96)));
    layer0_outputs(8655) <= not((inputs(215)) xor (inputs(238)));
    layer0_outputs(8656) <= inputs(124);
    layer0_outputs(8657) <= (inputs(224)) and not (inputs(204));
    layer0_outputs(8658) <= not(inputs(106)) or (inputs(93));
    layer0_outputs(8659) <= not((inputs(205)) or (inputs(93)));
    layer0_outputs(8660) <= not((inputs(53)) xor (inputs(218)));
    layer0_outputs(8661) <= inputs(55);
    layer0_outputs(8662) <= inputs(39);
    layer0_outputs(8663) <= (inputs(2)) xor (inputs(240));
    layer0_outputs(8664) <= (inputs(53)) xor (inputs(212));
    layer0_outputs(8665) <= inputs(200);
    layer0_outputs(8666) <= not(inputs(136));
    layer0_outputs(8667) <= not((inputs(139)) or (inputs(44)));
    layer0_outputs(8668) <= (inputs(148)) and not (inputs(207));
    layer0_outputs(8669) <= (inputs(218)) and (inputs(63));
    layer0_outputs(8670) <= not(inputs(60));
    layer0_outputs(8671) <= inputs(154);
    layer0_outputs(8672) <= not(inputs(119)) or (inputs(89));
    layer0_outputs(8673) <= not(inputs(15));
    layer0_outputs(8674) <= not(inputs(66)) or (inputs(64));
    layer0_outputs(8675) <= not((inputs(17)) xor (inputs(254)));
    layer0_outputs(8676) <= not((inputs(199)) xor (inputs(13)));
    layer0_outputs(8677) <= (inputs(40)) and not (inputs(99));
    layer0_outputs(8678) <= (inputs(246)) and not (inputs(236));
    layer0_outputs(8679) <= inputs(133);
    layer0_outputs(8680) <= inputs(100);
    layer0_outputs(8681) <= (inputs(139)) xor (inputs(53));
    layer0_outputs(8682) <= not((inputs(125)) or (inputs(83)));
    layer0_outputs(8683) <= not(inputs(243));
    layer0_outputs(8684) <= (inputs(70)) or (inputs(236));
    layer0_outputs(8685) <= (inputs(196)) and not (inputs(129));
    layer0_outputs(8686) <= not((inputs(208)) xor (inputs(138)));
    layer0_outputs(8687) <= (inputs(149)) and not (inputs(146));
    layer0_outputs(8688) <= not(inputs(64));
    layer0_outputs(8689) <= (inputs(72)) or (inputs(191));
    layer0_outputs(8690) <= not((inputs(137)) xor (inputs(140)));
    layer0_outputs(8691) <= (inputs(209)) and not (inputs(12));
    layer0_outputs(8692) <= (inputs(214)) and (inputs(170));
    layer0_outputs(8693) <= inputs(156);
    layer0_outputs(8694) <= inputs(189);
    layer0_outputs(8695) <= not((inputs(34)) and (inputs(1)));
    layer0_outputs(8696) <= not(inputs(50));
    layer0_outputs(8697) <= (inputs(169)) and not (inputs(19));
    layer0_outputs(8698) <= inputs(167);
    layer0_outputs(8699) <= (inputs(170)) and not (inputs(69));
    layer0_outputs(8700) <= not((inputs(112)) or (inputs(173)));
    layer0_outputs(8701) <= (inputs(83)) and not (inputs(74));
    layer0_outputs(8702) <= not((inputs(8)) xor (inputs(56)));
    layer0_outputs(8703) <= inputs(24);
    layer0_outputs(8704) <= not(inputs(60));
    layer0_outputs(8705) <= not(inputs(108));
    layer0_outputs(8706) <= '0';
    layer0_outputs(8707) <= not((inputs(232)) xor (inputs(14)));
    layer0_outputs(8708) <= (inputs(217)) and not (inputs(64));
    layer0_outputs(8709) <= not((inputs(31)) or (inputs(221)));
    layer0_outputs(8710) <= not(inputs(182));
    layer0_outputs(8711) <= inputs(184);
    layer0_outputs(8712) <= not(inputs(197)) or (inputs(242));
    layer0_outputs(8713) <= '0';
    layer0_outputs(8714) <= (inputs(146)) or (inputs(144));
    layer0_outputs(8715) <= (inputs(148)) and not (inputs(227));
    layer0_outputs(8716) <= not((inputs(213)) xor (inputs(166)));
    layer0_outputs(8717) <= (inputs(66)) or (inputs(255));
    layer0_outputs(8718) <= not(inputs(229));
    layer0_outputs(8719) <= '0';
    layer0_outputs(8720) <= (inputs(35)) xor (inputs(75));
    layer0_outputs(8721) <= (inputs(125)) or (inputs(255));
    layer0_outputs(8722) <= not(inputs(253));
    layer0_outputs(8723) <= not(inputs(202));
    layer0_outputs(8724) <= '1';
    layer0_outputs(8725) <= not((inputs(43)) or (inputs(18)));
    layer0_outputs(8726) <= not(inputs(105)) or (inputs(40));
    layer0_outputs(8727) <= not(inputs(16)) or (inputs(37));
    layer0_outputs(8728) <= '1';
    layer0_outputs(8729) <= (inputs(95)) or (inputs(86));
    layer0_outputs(8730) <= not(inputs(96)) or (inputs(8));
    layer0_outputs(8731) <= not((inputs(118)) xor (inputs(93)));
    layer0_outputs(8732) <= not(inputs(131));
    layer0_outputs(8733) <= not(inputs(205)) or (inputs(20));
    layer0_outputs(8734) <= not(inputs(108));
    layer0_outputs(8735) <= not(inputs(204)) or (inputs(46));
    layer0_outputs(8736) <= not(inputs(221)) or (inputs(110));
    layer0_outputs(8737) <= (inputs(215)) xor (inputs(221));
    layer0_outputs(8738) <= (inputs(131)) and not (inputs(5));
    layer0_outputs(8739) <= not(inputs(198)) or (inputs(170));
    layer0_outputs(8740) <= not((inputs(149)) or (inputs(142)));
    layer0_outputs(8741) <= not((inputs(116)) and (inputs(114)));
    layer0_outputs(8742) <= not(inputs(73));
    layer0_outputs(8743) <= inputs(35);
    layer0_outputs(8744) <= inputs(76);
    layer0_outputs(8745) <= '0';
    layer0_outputs(8746) <= not((inputs(247)) or (inputs(165)));
    layer0_outputs(8747) <= not(inputs(139)) or (inputs(245));
    layer0_outputs(8748) <= not(inputs(42));
    layer0_outputs(8749) <= not((inputs(99)) xor (inputs(33)));
    layer0_outputs(8750) <= not((inputs(25)) and (inputs(134)));
    layer0_outputs(8751) <= not(inputs(117));
    layer0_outputs(8752) <= (inputs(162)) and (inputs(245));
    layer0_outputs(8753) <= (inputs(126)) and not (inputs(48));
    layer0_outputs(8754) <= (inputs(51)) or (inputs(59));
    layer0_outputs(8755) <= not(inputs(139));
    layer0_outputs(8756) <= (inputs(39)) xor (inputs(156));
    layer0_outputs(8757) <= (inputs(170)) xor (inputs(220));
    layer0_outputs(8758) <= (inputs(226)) or (inputs(220));
    layer0_outputs(8759) <= '1';
    layer0_outputs(8760) <= not(inputs(24)) or (inputs(59));
    layer0_outputs(8761) <= (inputs(76)) or (inputs(203));
    layer0_outputs(8762) <= not(inputs(155)) or (inputs(61));
    layer0_outputs(8763) <= inputs(102);
    layer0_outputs(8764) <= (inputs(23)) or (inputs(40));
    layer0_outputs(8765) <= not(inputs(119));
    layer0_outputs(8766) <= not(inputs(38));
    layer0_outputs(8767) <= '0';
    layer0_outputs(8768) <= (inputs(245)) and not (inputs(9));
    layer0_outputs(8769) <= not(inputs(12)) or (inputs(29));
    layer0_outputs(8770) <= (inputs(138)) and not (inputs(163));
    layer0_outputs(8771) <= not(inputs(56));
    layer0_outputs(8772) <= (inputs(30)) or (inputs(132));
    layer0_outputs(8773) <= not(inputs(147)) or (inputs(97));
    layer0_outputs(8774) <= not((inputs(187)) xor (inputs(8)));
    layer0_outputs(8775) <= not((inputs(115)) or (inputs(252)));
    layer0_outputs(8776) <= inputs(72);
    layer0_outputs(8777) <= not((inputs(240)) xor (inputs(216)));
    layer0_outputs(8778) <= inputs(6);
    layer0_outputs(8779) <= not(inputs(189));
    layer0_outputs(8780) <= (inputs(122)) and not (inputs(65));
    layer0_outputs(8781) <= not(inputs(158));
    layer0_outputs(8782) <= (inputs(139)) xor (inputs(65));
    layer0_outputs(8783) <= (inputs(98)) xor (inputs(82));
    layer0_outputs(8784) <= (inputs(148)) xor (inputs(109));
    layer0_outputs(8785) <= (inputs(98)) and not (inputs(234));
    layer0_outputs(8786) <= not(inputs(33)) or (inputs(50));
    layer0_outputs(8787) <= inputs(75);
    layer0_outputs(8788) <= not(inputs(93));
    layer0_outputs(8789) <= not(inputs(89));
    layer0_outputs(8790) <= not(inputs(99));
    layer0_outputs(8791) <= (inputs(193)) xor (inputs(114));
    layer0_outputs(8792) <= not((inputs(67)) xor (inputs(28)));
    layer0_outputs(8793) <= not(inputs(87));
    layer0_outputs(8794) <= not(inputs(46));
    layer0_outputs(8795) <= (inputs(141)) and not (inputs(11));
    layer0_outputs(8796) <= inputs(7);
    layer0_outputs(8797) <= inputs(114);
    layer0_outputs(8798) <= inputs(139);
    layer0_outputs(8799) <= (inputs(187)) xor (inputs(117));
    layer0_outputs(8800) <= '1';
    layer0_outputs(8801) <= not(inputs(215));
    layer0_outputs(8802) <= not(inputs(248));
    layer0_outputs(8803) <= inputs(135);
    layer0_outputs(8804) <= not(inputs(197));
    layer0_outputs(8805) <= not(inputs(131)) or (inputs(246));
    layer0_outputs(8806) <= not(inputs(35));
    layer0_outputs(8807) <= inputs(137);
    layer0_outputs(8808) <= not(inputs(246));
    layer0_outputs(8809) <= (inputs(198)) and not (inputs(160));
    layer0_outputs(8810) <= not((inputs(40)) or (inputs(7)));
    layer0_outputs(8811) <= not((inputs(39)) xor (inputs(244)));
    layer0_outputs(8812) <= not(inputs(253)) or (inputs(143));
    layer0_outputs(8813) <= inputs(30);
    layer0_outputs(8814) <= (inputs(62)) or (inputs(157));
    layer0_outputs(8815) <= '1';
    layer0_outputs(8816) <= (inputs(180)) and not (inputs(81));
    layer0_outputs(8817) <= not(inputs(74));
    layer0_outputs(8818) <= not((inputs(87)) xor (inputs(97)));
    layer0_outputs(8819) <= not((inputs(151)) xor (inputs(11)));
    layer0_outputs(8820) <= not(inputs(15));
    layer0_outputs(8821) <= '0';
    layer0_outputs(8822) <= not(inputs(74));
    layer0_outputs(8823) <= not(inputs(157));
    layer0_outputs(8824) <= not((inputs(170)) or (inputs(181)));
    layer0_outputs(8825) <= not(inputs(194)) or (inputs(233));
    layer0_outputs(8826) <= (inputs(205)) xor (inputs(15));
    layer0_outputs(8827) <= not((inputs(105)) xor (inputs(190)));
    layer0_outputs(8828) <= (inputs(114)) and (inputs(80));
    layer0_outputs(8829) <= '1';
    layer0_outputs(8830) <= not((inputs(46)) xor (inputs(43)));
    layer0_outputs(8831) <= not((inputs(39)) or (inputs(125)));
    layer0_outputs(8832) <= '0';
    layer0_outputs(8833) <= (inputs(93)) or (inputs(198));
    layer0_outputs(8834) <= not(inputs(91));
    layer0_outputs(8835) <= (inputs(224)) or (inputs(208));
    layer0_outputs(8836) <= not(inputs(231)) or (inputs(41));
    layer0_outputs(8837) <= (inputs(253)) and not (inputs(115));
    layer0_outputs(8838) <= (inputs(178)) or (inputs(164));
    layer0_outputs(8839) <= inputs(94);
    layer0_outputs(8840) <= not((inputs(182)) xor (inputs(238)));
    layer0_outputs(8841) <= not(inputs(162)) or (inputs(210));
    layer0_outputs(8842) <= (inputs(239)) xor (inputs(223));
    layer0_outputs(8843) <= inputs(93);
    layer0_outputs(8844) <= not(inputs(160)) or (inputs(231));
    layer0_outputs(8845) <= not((inputs(130)) or (inputs(92)));
    layer0_outputs(8846) <= not(inputs(216)) or (inputs(199));
    layer0_outputs(8847) <= not(inputs(88)) or (inputs(5));
    layer0_outputs(8848) <= inputs(106);
    layer0_outputs(8849) <= (inputs(104)) or (inputs(228));
    layer0_outputs(8850) <= (inputs(20)) or (inputs(131));
    layer0_outputs(8851) <= (inputs(157)) or (inputs(54));
    layer0_outputs(8852) <= not(inputs(203)) or (inputs(228));
    layer0_outputs(8853) <= not(inputs(57));
    layer0_outputs(8854) <= (inputs(158)) and not (inputs(145));
    layer0_outputs(8855) <= (inputs(111)) and (inputs(147));
    layer0_outputs(8856) <= '1';
    layer0_outputs(8857) <= not((inputs(84)) or (inputs(62)));
    layer0_outputs(8858) <= (inputs(151)) and not (inputs(54));
    layer0_outputs(8859) <= inputs(201);
    layer0_outputs(8860) <= (inputs(85)) and not (inputs(151));
    layer0_outputs(8861) <= not((inputs(243)) and (inputs(95)));
    layer0_outputs(8862) <= inputs(199);
    layer0_outputs(8863) <= '0';
    layer0_outputs(8864) <= not((inputs(99)) or (inputs(140)));
    layer0_outputs(8865) <= not(inputs(73)) or (inputs(15));
    layer0_outputs(8866) <= not(inputs(111)) or (inputs(209));
    layer0_outputs(8867) <= not((inputs(37)) or (inputs(52)));
    layer0_outputs(8868) <= not(inputs(101));
    layer0_outputs(8869) <= not(inputs(101));
    layer0_outputs(8870) <= not(inputs(242));
    layer0_outputs(8871) <= inputs(9);
    layer0_outputs(8872) <= not(inputs(118)) or (inputs(2));
    layer0_outputs(8873) <= not((inputs(161)) or (inputs(127)));
    layer0_outputs(8874) <= not(inputs(185)) or (inputs(97));
    layer0_outputs(8875) <= not(inputs(242));
    layer0_outputs(8876) <= (inputs(218)) and not (inputs(158));
    layer0_outputs(8877) <= (inputs(247)) and not (inputs(193));
    layer0_outputs(8878) <= not((inputs(7)) or (inputs(121)));
    layer0_outputs(8879) <= not(inputs(148));
    layer0_outputs(8880) <= not(inputs(148));
    layer0_outputs(8881) <= (inputs(185)) or (inputs(215));
    layer0_outputs(8882) <= (inputs(14)) and not (inputs(129));
    layer0_outputs(8883) <= (inputs(72)) and not (inputs(147));
    layer0_outputs(8884) <= not(inputs(135)) or (inputs(244));
    layer0_outputs(8885) <= not(inputs(124));
    layer0_outputs(8886) <= not(inputs(180)) or (inputs(28));
    layer0_outputs(8887) <= not((inputs(193)) xor (inputs(78)));
    layer0_outputs(8888) <= not(inputs(205)) or (inputs(235));
    layer0_outputs(8889) <= (inputs(213)) and not (inputs(172));
    layer0_outputs(8890) <= inputs(4);
    layer0_outputs(8891) <= not((inputs(175)) or (inputs(37)));
    layer0_outputs(8892) <= not((inputs(92)) xor (inputs(193)));
    layer0_outputs(8893) <= not(inputs(76));
    layer0_outputs(8894) <= inputs(104);
    layer0_outputs(8895) <= not(inputs(137)) or (inputs(94));
    layer0_outputs(8896) <= (inputs(96)) and not (inputs(236));
    layer0_outputs(8897) <= inputs(138);
    layer0_outputs(8898) <= not((inputs(41)) or (inputs(140)));
    layer0_outputs(8899) <= (inputs(33)) or (inputs(171));
    layer0_outputs(8900) <= (inputs(86)) and not (inputs(27));
    layer0_outputs(8901) <= not((inputs(14)) or (inputs(118)));
    layer0_outputs(8902) <= not((inputs(231)) or (inputs(6)));
    layer0_outputs(8903) <= not(inputs(124));
    layer0_outputs(8904) <= (inputs(249)) and not (inputs(3));
    layer0_outputs(8905) <= (inputs(146)) xor (inputs(44));
    layer0_outputs(8906) <= inputs(27);
    layer0_outputs(8907) <= inputs(214);
    layer0_outputs(8908) <= (inputs(54)) xor (inputs(57));
    layer0_outputs(8909) <= (inputs(40)) and not (inputs(64));
    layer0_outputs(8910) <= (inputs(8)) or (inputs(76));
    layer0_outputs(8911) <= not(inputs(84)) or (inputs(23));
    layer0_outputs(8912) <= not((inputs(255)) and (inputs(50)));
    layer0_outputs(8913) <= (inputs(88)) or (inputs(248));
    layer0_outputs(8914) <= (inputs(176)) or (inputs(209));
    layer0_outputs(8915) <= not(inputs(92));
    layer0_outputs(8916) <= '1';
    layer0_outputs(8917) <= '0';
    layer0_outputs(8918) <= (inputs(28)) and (inputs(81));
    layer0_outputs(8919) <= (inputs(213)) and not (inputs(180));
    layer0_outputs(8920) <= not((inputs(61)) and (inputs(33)));
    layer0_outputs(8921) <= not((inputs(231)) or (inputs(135)));
    layer0_outputs(8922) <= not((inputs(193)) or (inputs(208)));
    layer0_outputs(8923) <= (inputs(9)) and not (inputs(178));
    layer0_outputs(8924) <= not((inputs(97)) or (inputs(231)));
    layer0_outputs(8925) <= not(inputs(118));
    layer0_outputs(8926) <= not((inputs(145)) xor (inputs(14)));
    layer0_outputs(8927) <= (inputs(74)) and not (inputs(19));
    layer0_outputs(8928) <= not((inputs(248)) or (inputs(220)));
    layer0_outputs(8929) <= not((inputs(248)) and (inputs(127)));
    layer0_outputs(8930) <= (inputs(37)) and not (inputs(62));
    layer0_outputs(8931) <= not(inputs(234));
    layer0_outputs(8932) <= inputs(37);
    layer0_outputs(8933) <= not(inputs(216));
    layer0_outputs(8934) <= '0';
    layer0_outputs(8935) <= not(inputs(44));
    layer0_outputs(8936) <= (inputs(72)) xor (inputs(41));
    layer0_outputs(8937) <= not((inputs(102)) xor (inputs(32)));
    layer0_outputs(8938) <= inputs(185);
    layer0_outputs(8939) <= not(inputs(167)) or (inputs(113));
    layer0_outputs(8940) <= (inputs(73)) and not (inputs(30));
    layer0_outputs(8941) <= inputs(179);
    layer0_outputs(8942) <= not(inputs(101));
    layer0_outputs(8943) <= (inputs(165)) or (inputs(108));
    layer0_outputs(8944) <= (inputs(58)) and not (inputs(161));
    layer0_outputs(8945) <= not((inputs(126)) xor (inputs(38)));
    layer0_outputs(8946) <= (inputs(132)) or (inputs(187));
    layer0_outputs(8947) <= not((inputs(151)) or (inputs(239)));
    layer0_outputs(8948) <= not((inputs(196)) or (inputs(155)));
    layer0_outputs(8949) <= not(inputs(84));
    layer0_outputs(8950) <= (inputs(158)) and not (inputs(160));
    layer0_outputs(8951) <= inputs(217);
    layer0_outputs(8952) <= not(inputs(117));
    layer0_outputs(8953) <= '0';
    layer0_outputs(8954) <= (inputs(103)) and not (inputs(224));
    layer0_outputs(8955) <= not(inputs(199));
    layer0_outputs(8956) <= inputs(136);
    layer0_outputs(8957) <= (inputs(101)) and not (inputs(22));
    layer0_outputs(8958) <= inputs(128);
    layer0_outputs(8959) <= not(inputs(120));
    layer0_outputs(8960) <= not((inputs(42)) xor (inputs(7)));
    layer0_outputs(8961) <= not(inputs(49)) or (inputs(35));
    layer0_outputs(8962) <= inputs(232);
    layer0_outputs(8963) <= inputs(106);
    layer0_outputs(8964) <= not(inputs(143)) or (inputs(175));
    layer0_outputs(8965) <= not(inputs(2));
    layer0_outputs(8966) <= (inputs(217)) xor (inputs(88));
    layer0_outputs(8967) <= not(inputs(91));
    layer0_outputs(8968) <= not(inputs(228));
    layer0_outputs(8969) <= not((inputs(0)) xor (inputs(124)));
    layer0_outputs(8970) <= not((inputs(17)) xor (inputs(85)));
    layer0_outputs(8971) <= not(inputs(71)) or (inputs(246));
    layer0_outputs(8972) <= '0';
    layer0_outputs(8973) <= (inputs(179)) and not (inputs(251));
    layer0_outputs(8974) <= not(inputs(123));
    layer0_outputs(8975) <= (inputs(28)) xor (inputs(120));
    layer0_outputs(8976) <= (inputs(40)) xor (inputs(96));
    layer0_outputs(8977) <= not((inputs(76)) xor (inputs(26)));
    layer0_outputs(8978) <= (inputs(56)) or (inputs(171));
    layer0_outputs(8979) <= not((inputs(68)) and (inputs(238)));
    layer0_outputs(8980) <= (inputs(210)) or (inputs(53));
    layer0_outputs(8981) <= inputs(245);
    layer0_outputs(8982) <= not((inputs(94)) or (inputs(100)));
    layer0_outputs(8983) <= inputs(225);
    layer0_outputs(8984) <= (inputs(45)) xor (inputs(23));
    layer0_outputs(8985) <= (inputs(176)) and not (inputs(97));
    layer0_outputs(8986) <= not(inputs(126)) or (inputs(76));
    layer0_outputs(8987) <= inputs(115);
    layer0_outputs(8988) <= not(inputs(218)) or (inputs(160));
    layer0_outputs(8989) <= (inputs(50)) and (inputs(146));
    layer0_outputs(8990) <= not(inputs(221));
    layer0_outputs(8991) <= (inputs(205)) xor (inputs(180));
    layer0_outputs(8992) <= (inputs(246)) and not (inputs(28));
    layer0_outputs(8993) <= not((inputs(181)) xor (inputs(163)));
    layer0_outputs(8994) <= (inputs(42)) or (inputs(32));
    layer0_outputs(8995) <= (inputs(236)) xor (inputs(166));
    layer0_outputs(8996) <= inputs(188);
    layer0_outputs(8997) <= '0';
    layer0_outputs(8998) <= '0';
    layer0_outputs(8999) <= (inputs(184)) and not (inputs(76));
    layer0_outputs(9000) <= not((inputs(112)) xor (inputs(149)));
    layer0_outputs(9001) <= (inputs(143)) and not (inputs(176));
    layer0_outputs(9002) <= (inputs(243)) and not (inputs(67));
    layer0_outputs(9003) <= inputs(122);
    layer0_outputs(9004) <= not(inputs(9)) or (inputs(4));
    layer0_outputs(9005) <= (inputs(104)) xor (inputs(255));
    layer0_outputs(9006) <= not((inputs(37)) xor (inputs(225)));
    layer0_outputs(9007) <= not((inputs(174)) or (inputs(156)));
    layer0_outputs(9008) <= '1';
    layer0_outputs(9009) <= not((inputs(150)) or (inputs(244)));
    layer0_outputs(9010) <= inputs(235);
    layer0_outputs(9011) <= inputs(104);
    layer0_outputs(9012) <= not((inputs(102)) or (inputs(123)));
    layer0_outputs(9013) <= not(inputs(136)) or (inputs(13));
    layer0_outputs(9014) <= not(inputs(187));
    layer0_outputs(9015) <= not(inputs(159)) or (inputs(129));
    layer0_outputs(9016) <= inputs(119);
    layer0_outputs(9017) <= not(inputs(149)) or (inputs(24));
    layer0_outputs(9018) <= not((inputs(27)) or (inputs(154)));
    layer0_outputs(9019) <= '0';
    layer0_outputs(9020) <= not(inputs(167)) or (inputs(42));
    layer0_outputs(9021) <= (inputs(47)) xor (inputs(76));
    layer0_outputs(9022) <= not(inputs(120));
    layer0_outputs(9023) <= '1';
    layer0_outputs(9024) <= (inputs(134)) xor (inputs(54));
    layer0_outputs(9025) <= (inputs(149)) xor (inputs(145));
    layer0_outputs(9026) <= not((inputs(133)) xor (inputs(146)));
    layer0_outputs(9027) <= not(inputs(105));
    layer0_outputs(9028) <= not(inputs(25)) or (inputs(145));
    layer0_outputs(9029) <= (inputs(149)) or (inputs(126));
    layer0_outputs(9030) <= (inputs(118)) and not (inputs(192));
    layer0_outputs(9031) <= not(inputs(150)) or (inputs(13));
    layer0_outputs(9032) <= inputs(121);
    layer0_outputs(9033) <= not(inputs(89));
    layer0_outputs(9034) <= (inputs(186)) or (inputs(187));
    layer0_outputs(9035) <= not((inputs(57)) or (inputs(166)));
    layer0_outputs(9036) <= not(inputs(8));
    layer0_outputs(9037) <= not((inputs(162)) xor (inputs(154)));
    layer0_outputs(9038) <= (inputs(215)) and not (inputs(60));
    layer0_outputs(9039) <= not(inputs(144));
    layer0_outputs(9040) <= not(inputs(34)) or (inputs(3));
    layer0_outputs(9041) <= not((inputs(125)) or (inputs(20)));
    layer0_outputs(9042) <= not((inputs(134)) xor (inputs(80)));
    layer0_outputs(9043) <= not((inputs(11)) or (inputs(74)));
    layer0_outputs(9044) <= not((inputs(80)) xor (inputs(235)));
    layer0_outputs(9045) <= not((inputs(49)) xor (inputs(88)));
    layer0_outputs(9046) <= not(inputs(244));
    layer0_outputs(9047) <= (inputs(0)) or (inputs(151));
    layer0_outputs(9048) <= (inputs(139)) and not (inputs(240));
    layer0_outputs(9049) <= not(inputs(8));
    layer0_outputs(9050) <= (inputs(230)) and (inputs(41));
    layer0_outputs(9051) <= not(inputs(249)) or (inputs(89));
    layer0_outputs(9052) <= (inputs(42)) and not (inputs(159));
    layer0_outputs(9053) <= inputs(135);
    layer0_outputs(9054) <= (inputs(100)) and not (inputs(157));
    layer0_outputs(9055) <= not((inputs(208)) or (inputs(68)));
    layer0_outputs(9056) <= (inputs(109)) or (inputs(184));
    layer0_outputs(9057) <= (inputs(146)) xor (inputs(226));
    layer0_outputs(9058) <= not(inputs(230)) or (inputs(156));
    layer0_outputs(9059) <= (inputs(203)) and not (inputs(224));
    layer0_outputs(9060) <= not(inputs(124));
    layer0_outputs(9061) <= not((inputs(188)) or (inputs(135)));
    layer0_outputs(9062) <= inputs(216);
    layer0_outputs(9063) <= not(inputs(230)) or (inputs(148));
    layer0_outputs(9064) <= not((inputs(190)) xor (inputs(83)));
    layer0_outputs(9065) <= (inputs(197)) and not (inputs(249));
    layer0_outputs(9066) <= not((inputs(158)) xor (inputs(222)));
    layer0_outputs(9067) <= not((inputs(23)) and (inputs(242)));
    layer0_outputs(9068) <= not((inputs(173)) or (inputs(139)));
    layer0_outputs(9069) <= not((inputs(27)) xor (inputs(72)));
    layer0_outputs(9070) <= inputs(200);
    layer0_outputs(9071) <= (inputs(53)) xor (inputs(84));
    layer0_outputs(9072) <= (inputs(123)) or (inputs(159));
    layer0_outputs(9073) <= (inputs(216)) or (inputs(243));
    layer0_outputs(9074) <= not(inputs(86)) or (inputs(16));
    layer0_outputs(9075) <= inputs(152);
    layer0_outputs(9076) <= not(inputs(239));
    layer0_outputs(9077) <= (inputs(59)) and not (inputs(235));
    layer0_outputs(9078) <= inputs(52);
    layer0_outputs(9079) <= (inputs(74)) or (inputs(31));
    layer0_outputs(9080) <= not(inputs(17)) or (inputs(194));
    layer0_outputs(9081) <= not(inputs(140)) or (inputs(41));
    layer0_outputs(9082) <= not((inputs(14)) or (inputs(58)));
    layer0_outputs(9083) <= not((inputs(127)) or (inputs(158)));
    layer0_outputs(9084) <= (inputs(175)) and not (inputs(241));
    layer0_outputs(9085) <= not((inputs(240)) xor (inputs(106)));
    layer0_outputs(9086) <= not(inputs(94));
    layer0_outputs(9087) <= '1';
    layer0_outputs(9088) <= (inputs(8)) or (inputs(236));
    layer0_outputs(9089) <= inputs(52);
    layer0_outputs(9090) <= (inputs(9)) and not (inputs(209));
    layer0_outputs(9091) <= not(inputs(77)) or (inputs(194));
    layer0_outputs(9092) <= not(inputs(99)) or (inputs(222));
    layer0_outputs(9093) <= not(inputs(77));
    layer0_outputs(9094) <= not(inputs(213)) or (inputs(210));
    layer0_outputs(9095) <= inputs(41);
    layer0_outputs(9096) <= not(inputs(120));
    layer0_outputs(9097) <= inputs(7);
    layer0_outputs(9098) <= (inputs(87)) and not (inputs(209));
    layer0_outputs(9099) <= not(inputs(153)) or (inputs(248));
    layer0_outputs(9100) <= '1';
    layer0_outputs(9101) <= inputs(61);
    layer0_outputs(9102) <= '1';
    layer0_outputs(9103) <= (inputs(35)) xor (inputs(164));
    layer0_outputs(9104) <= (inputs(232)) and not (inputs(203));
    layer0_outputs(9105) <= (inputs(20)) xor (inputs(127));
    layer0_outputs(9106) <= (inputs(105)) or (inputs(220));
    layer0_outputs(9107) <= inputs(23);
    layer0_outputs(9108) <= not(inputs(80));
    layer0_outputs(9109) <= not(inputs(184)) or (inputs(18));
    layer0_outputs(9110) <= not(inputs(100)) or (inputs(128));
    layer0_outputs(9111) <= (inputs(57)) and not (inputs(96));
    layer0_outputs(9112) <= not((inputs(222)) xor (inputs(148)));
    layer0_outputs(9113) <= inputs(166);
    layer0_outputs(9114) <= inputs(183);
    layer0_outputs(9115) <= (inputs(8)) or (inputs(118));
    layer0_outputs(9116) <= not((inputs(4)) or (inputs(41)));
    layer0_outputs(9117) <= (inputs(229)) and not (inputs(222));
    layer0_outputs(9118) <= not((inputs(209)) xor (inputs(92)));
    layer0_outputs(9119) <= not(inputs(128)) or (inputs(0));
    layer0_outputs(9120) <= not((inputs(143)) or (inputs(55)));
    layer0_outputs(9121) <= (inputs(186)) and not (inputs(115));
    layer0_outputs(9122) <= not((inputs(192)) xor (inputs(248)));
    layer0_outputs(9123) <= inputs(78);
    layer0_outputs(9124) <= not((inputs(68)) xor (inputs(159)));
    layer0_outputs(9125) <= (inputs(40)) or (inputs(187));
    layer0_outputs(9126) <= not(inputs(113));
    layer0_outputs(9127) <= not(inputs(15)) or (inputs(83));
    layer0_outputs(9128) <= not(inputs(31)) or (inputs(3));
    layer0_outputs(9129) <= not((inputs(34)) or (inputs(118)));
    layer0_outputs(9130) <= not(inputs(135));
    layer0_outputs(9131) <= (inputs(11)) or (inputs(213));
    layer0_outputs(9132) <= not((inputs(77)) or (inputs(21)));
    layer0_outputs(9133) <= (inputs(176)) and not (inputs(210));
    layer0_outputs(9134) <= '0';
    layer0_outputs(9135) <= not((inputs(235)) xor (inputs(237)));
    layer0_outputs(9136) <= (inputs(210)) xor (inputs(126));
    layer0_outputs(9137) <= not(inputs(247));
    layer0_outputs(9138) <= not(inputs(168));
    layer0_outputs(9139) <= not((inputs(213)) or (inputs(220)));
    layer0_outputs(9140) <= (inputs(2)) and not (inputs(82));
    layer0_outputs(9141) <= inputs(32);
    layer0_outputs(9142) <= inputs(229);
    layer0_outputs(9143) <= inputs(127);
    layer0_outputs(9144) <= (inputs(8)) or (inputs(119));
    layer0_outputs(9145) <= not((inputs(112)) xor (inputs(56)));
    layer0_outputs(9146) <= inputs(177);
    layer0_outputs(9147) <= (inputs(241)) and not (inputs(34));
    layer0_outputs(9148) <= inputs(227);
    layer0_outputs(9149) <= not((inputs(222)) and (inputs(19)));
    layer0_outputs(9150) <= inputs(251);
    layer0_outputs(9151) <= (inputs(174)) and (inputs(113));
    layer0_outputs(9152) <= inputs(56);
    layer0_outputs(9153) <= not((inputs(158)) and (inputs(25)));
    layer0_outputs(9154) <= (inputs(204)) xor (inputs(90));
    layer0_outputs(9155) <= not(inputs(135)) or (inputs(211));
    layer0_outputs(9156) <= (inputs(17)) and not (inputs(14));
    layer0_outputs(9157) <= not(inputs(211)) or (inputs(11));
    layer0_outputs(9158) <= not((inputs(186)) xor (inputs(28)));
    layer0_outputs(9159) <= (inputs(216)) xor (inputs(211));
    layer0_outputs(9160) <= not((inputs(167)) or (inputs(191)));
    layer0_outputs(9161) <= inputs(219);
    layer0_outputs(9162) <= not(inputs(88));
    layer0_outputs(9163) <= inputs(159);
    layer0_outputs(9164) <= (inputs(79)) and (inputs(176));
    layer0_outputs(9165) <= inputs(141);
    layer0_outputs(9166) <= not((inputs(67)) or (inputs(6)));
    layer0_outputs(9167) <= not((inputs(108)) xor (inputs(137)));
    layer0_outputs(9168) <= not((inputs(179)) or (inputs(159)));
    layer0_outputs(9169) <= (inputs(234)) and not (inputs(83));
    layer0_outputs(9170) <= not((inputs(0)) xor (inputs(234)));
    layer0_outputs(9171) <= not(inputs(68)) or (inputs(201));
    layer0_outputs(9172) <= (inputs(206)) or (inputs(179));
    layer0_outputs(9173) <= (inputs(245)) or (inputs(3));
    layer0_outputs(9174) <= not((inputs(81)) and (inputs(63)));
    layer0_outputs(9175) <= (inputs(237)) and (inputs(220));
    layer0_outputs(9176) <= inputs(107);
    layer0_outputs(9177) <= inputs(177);
    layer0_outputs(9178) <= not(inputs(55)) or (inputs(104));
    layer0_outputs(9179) <= not((inputs(78)) xor (inputs(113)));
    layer0_outputs(9180) <= inputs(118);
    layer0_outputs(9181) <= inputs(121);
    layer0_outputs(9182) <= (inputs(60)) xor (inputs(215));
    layer0_outputs(9183) <= not((inputs(69)) or (inputs(153)));
    layer0_outputs(9184) <= (inputs(71)) and not (inputs(218));
    layer0_outputs(9185) <= (inputs(89)) and not (inputs(114));
    layer0_outputs(9186) <= inputs(68);
    layer0_outputs(9187) <= not(inputs(171));
    layer0_outputs(9188) <= not(inputs(181));
    layer0_outputs(9189) <= inputs(77);
    layer0_outputs(9190) <= (inputs(102)) or (inputs(163));
    layer0_outputs(9191) <= not((inputs(85)) or (inputs(14)));
    layer0_outputs(9192) <= not(inputs(201));
    layer0_outputs(9193) <= (inputs(157)) and (inputs(244));
    layer0_outputs(9194) <= not(inputs(116));
    layer0_outputs(9195) <= not(inputs(196));
    layer0_outputs(9196) <= not((inputs(166)) or (inputs(116)));
    layer0_outputs(9197) <= inputs(140);
    layer0_outputs(9198) <= inputs(87);
    layer0_outputs(9199) <= not(inputs(80)) or (inputs(157));
    layer0_outputs(9200) <= not(inputs(134)) or (inputs(219));
    layer0_outputs(9201) <= not(inputs(117));
    layer0_outputs(9202) <= not(inputs(175));
    layer0_outputs(9203) <= (inputs(139)) and (inputs(189));
    layer0_outputs(9204) <= (inputs(55)) xor (inputs(89));
    layer0_outputs(9205) <= (inputs(123)) xor (inputs(78));
    layer0_outputs(9206) <= not(inputs(137)) or (inputs(208));
    layer0_outputs(9207) <= (inputs(170)) xor (inputs(10));
    layer0_outputs(9208) <= (inputs(44)) or (inputs(89));
    layer0_outputs(9209) <= inputs(58);
    layer0_outputs(9210) <= (inputs(118)) or (inputs(37));
    layer0_outputs(9211) <= not(inputs(116));
    layer0_outputs(9212) <= not((inputs(86)) and (inputs(152)));
    layer0_outputs(9213) <= not(inputs(184)) or (inputs(93));
    layer0_outputs(9214) <= inputs(166);
    layer0_outputs(9215) <= not(inputs(104));
    layer0_outputs(9216) <= not(inputs(164));
    layer0_outputs(9217) <= '1';
    layer0_outputs(9218) <= not((inputs(103)) xor (inputs(73)));
    layer0_outputs(9219) <= not((inputs(197)) xor (inputs(227)));
    layer0_outputs(9220) <= (inputs(3)) or (inputs(130));
    layer0_outputs(9221) <= not((inputs(221)) or (inputs(214)));
    layer0_outputs(9222) <= inputs(66);
    layer0_outputs(9223) <= not((inputs(168)) or (inputs(53)));
    layer0_outputs(9224) <= not((inputs(68)) xor (inputs(243)));
    layer0_outputs(9225) <= inputs(53);
    layer0_outputs(9226) <= not((inputs(49)) or (inputs(105)));
    layer0_outputs(9227) <= (inputs(149)) and not (inputs(7));
    layer0_outputs(9228) <= (inputs(232)) xor (inputs(96));
    layer0_outputs(9229) <= not(inputs(30)) or (inputs(215));
    layer0_outputs(9230) <= inputs(147);
    layer0_outputs(9231) <= (inputs(58)) xor (inputs(107));
    layer0_outputs(9232) <= not(inputs(72));
    layer0_outputs(9233) <= (inputs(126)) or (inputs(167));
    layer0_outputs(9234) <= not(inputs(89));
    layer0_outputs(9235) <= not(inputs(217));
    layer0_outputs(9236) <= (inputs(5)) xor (inputs(38));
    layer0_outputs(9237) <= not(inputs(222));
    layer0_outputs(9238) <= not((inputs(40)) xor (inputs(58)));
    layer0_outputs(9239) <= not(inputs(199));
    layer0_outputs(9240) <= not(inputs(134)) or (inputs(28));
    layer0_outputs(9241) <= not((inputs(142)) and (inputs(46)));
    layer0_outputs(9242) <= inputs(64);
    layer0_outputs(9243) <= (inputs(187)) xor (inputs(75));
    layer0_outputs(9244) <= not(inputs(57));
    layer0_outputs(9245) <= inputs(167);
    layer0_outputs(9246) <= not(inputs(179));
    layer0_outputs(9247) <= not((inputs(43)) xor (inputs(0)));
    layer0_outputs(9248) <= not((inputs(66)) xor (inputs(15)));
    layer0_outputs(9249) <= (inputs(89)) and not (inputs(225));
    layer0_outputs(9250) <= not((inputs(155)) and (inputs(17)));
    layer0_outputs(9251) <= not((inputs(171)) or (inputs(241)));
    layer0_outputs(9252) <= not(inputs(138));
    layer0_outputs(9253) <= '0';
    layer0_outputs(9254) <= inputs(197);
    layer0_outputs(9255) <= not(inputs(54));
    layer0_outputs(9256) <= inputs(170);
    layer0_outputs(9257) <= (inputs(8)) or (inputs(28));
    layer0_outputs(9258) <= not((inputs(53)) or (inputs(122)));
    layer0_outputs(9259) <= (inputs(204)) or (inputs(196));
    layer0_outputs(9260) <= inputs(223);
    layer0_outputs(9261) <= not(inputs(89));
    layer0_outputs(9262) <= inputs(185);
    layer0_outputs(9263) <= (inputs(140)) and not (inputs(94));
    layer0_outputs(9264) <= not(inputs(223)) or (inputs(225));
    layer0_outputs(9265) <= not((inputs(52)) or (inputs(194)));
    layer0_outputs(9266) <= (inputs(133)) and not (inputs(219));
    layer0_outputs(9267) <= (inputs(254)) and not (inputs(158));
    layer0_outputs(9268) <= inputs(7);
    layer0_outputs(9269) <= inputs(164);
    layer0_outputs(9270) <= not((inputs(146)) xor (inputs(196)));
    layer0_outputs(9271) <= not(inputs(121)) or (inputs(45));
    layer0_outputs(9272) <= (inputs(81)) and not (inputs(110));
    layer0_outputs(9273) <= '0';
    layer0_outputs(9274) <= not(inputs(173)) or (inputs(251));
    layer0_outputs(9275) <= inputs(163);
    layer0_outputs(9276) <= (inputs(123)) or (inputs(179));
    layer0_outputs(9277) <= not((inputs(217)) and (inputs(17)));
    layer0_outputs(9278) <= not((inputs(88)) or (inputs(5)));
    layer0_outputs(9279) <= (inputs(242)) and not (inputs(192));
    layer0_outputs(9280) <= (inputs(132)) or (inputs(16));
    layer0_outputs(9281) <= (inputs(218)) xor (inputs(214));
    layer0_outputs(9282) <= not(inputs(104));
    layer0_outputs(9283) <= inputs(70);
    layer0_outputs(9284) <= not(inputs(0));
    layer0_outputs(9285) <= not(inputs(189));
    layer0_outputs(9286) <= inputs(224);
    layer0_outputs(9287) <= not(inputs(136));
    layer0_outputs(9288) <= not(inputs(206));
    layer0_outputs(9289) <= not(inputs(187));
    layer0_outputs(9290) <= not((inputs(24)) or (inputs(11)));
    layer0_outputs(9291) <= not(inputs(190));
    layer0_outputs(9292) <= not(inputs(44)) or (inputs(7));
    layer0_outputs(9293) <= not(inputs(15));
    layer0_outputs(9294) <= not((inputs(51)) or (inputs(108)));
    layer0_outputs(9295) <= not((inputs(254)) and (inputs(143)));
    layer0_outputs(9296) <= not((inputs(63)) and (inputs(211)));
    layer0_outputs(9297) <= not(inputs(97)) or (inputs(157));
    layer0_outputs(9298) <= not(inputs(191)) or (inputs(36));
    layer0_outputs(9299) <= not(inputs(73));
    layer0_outputs(9300) <= not((inputs(202)) or (inputs(149)));
    layer0_outputs(9301) <= (inputs(66)) or (inputs(69));
    layer0_outputs(9302) <= (inputs(251)) xor (inputs(62));
    layer0_outputs(9303) <= not((inputs(241)) xor (inputs(151)));
    layer0_outputs(9304) <= not(inputs(147)) or (inputs(12));
    layer0_outputs(9305) <= (inputs(53)) xor (inputs(103));
    layer0_outputs(9306) <= not((inputs(139)) or (inputs(25)));
    layer0_outputs(9307) <= (inputs(53)) or (inputs(232));
    layer0_outputs(9308) <= (inputs(138)) or (inputs(241));
    layer0_outputs(9309) <= not((inputs(47)) and (inputs(223)));
    layer0_outputs(9310) <= inputs(136);
    layer0_outputs(9311) <= (inputs(108)) and not (inputs(128));
    layer0_outputs(9312) <= not((inputs(211)) xor (inputs(33)));
    layer0_outputs(9313) <= (inputs(168)) and not (inputs(162));
    layer0_outputs(9314) <= inputs(126);
    layer0_outputs(9315) <= '1';
    layer0_outputs(9316) <= not(inputs(142));
    layer0_outputs(9317) <= inputs(166);
    layer0_outputs(9318) <= not((inputs(130)) xor (inputs(147)));
    layer0_outputs(9319) <= not((inputs(84)) xor (inputs(70)));
    layer0_outputs(9320) <= (inputs(163)) or (inputs(209));
    layer0_outputs(9321) <= not((inputs(207)) xor (inputs(154)));
    layer0_outputs(9322) <= inputs(118);
    layer0_outputs(9323) <= (inputs(137)) and not (inputs(5));
    layer0_outputs(9324) <= not((inputs(27)) and (inputs(111)));
    layer0_outputs(9325) <= (inputs(40)) and not (inputs(100));
    layer0_outputs(9326) <= inputs(23);
    layer0_outputs(9327) <= (inputs(26)) and not (inputs(30));
    layer0_outputs(9328) <= (inputs(122)) or (inputs(203));
    layer0_outputs(9329) <= (inputs(110)) or (inputs(62));
    layer0_outputs(9330) <= (inputs(147)) or (inputs(117));
    layer0_outputs(9331) <= inputs(236);
    layer0_outputs(9332) <= not(inputs(140));
    layer0_outputs(9333) <= (inputs(171)) or (inputs(6));
    layer0_outputs(9334) <= inputs(231);
    layer0_outputs(9335) <= not((inputs(194)) or (inputs(55)));
    layer0_outputs(9336) <= (inputs(5)) xor (inputs(193));
    layer0_outputs(9337) <= (inputs(26)) or (inputs(20));
    layer0_outputs(9338) <= inputs(255);
    layer0_outputs(9339) <= (inputs(54)) or (inputs(167));
    layer0_outputs(9340) <= (inputs(9)) xor (inputs(216));
    layer0_outputs(9341) <= (inputs(150)) and not (inputs(160));
    layer0_outputs(9342) <= inputs(153);
    layer0_outputs(9343) <= (inputs(69)) xor (inputs(162));
    layer0_outputs(9344) <= not((inputs(111)) and (inputs(118)));
    layer0_outputs(9345) <= (inputs(138)) or (inputs(101));
    layer0_outputs(9346) <= inputs(141);
    layer0_outputs(9347) <= not(inputs(158));
    layer0_outputs(9348) <= inputs(104);
    layer0_outputs(9349) <= (inputs(86)) or (inputs(231));
    layer0_outputs(9350) <= '1';
    layer0_outputs(9351) <= not(inputs(149)) or (inputs(157));
    layer0_outputs(9352) <= '0';
    layer0_outputs(9353) <= (inputs(138)) xor (inputs(16));
    layer0_outputs(9354) <= not((inputs(147)) xor (inputs(134)));
    layer0_outputs(9355) <= (inputs(67)) and not (inputs(77));
    layer0_outputs(9356) <= (inputs(67)) or (inputs(50));
    layer0_outputs(9357) <= not((inputs(78)) xor (inputs(38)));
    layer0_outputs(9358) <= not(inputs(238)) or (inputs(49));
    layer0_outputs(9359) <= not((inputs(82)) or (inputs(162)));
    layer0_outputs(9360) <= not((inputs(147)) xor (inputs(34)));
    layer0_outputs(9361) <= not(inputs(181)) or (inputs(124));
    layer0_outputs(9362) <= (inputs(134)) and not (inputs(65));
    layer0_outputs(9363) <= not(inputs(148));
    layer0_outputs(9364) <= (inputs(205)) and not (inputs(20));
    layer0_outputs(9365) <= not((inputs(9)) xor (inputs(42)));
    layer0_outputs(9366) <= not((inputs(119)) or (inputs(241)));
    layer0_outputs(9367) <= not(inputs(195)) or (inputs(228));
    layer0_outputs(9368) <= not(inputs(140));
    layer0_outputs(9369) <= not(inputs(85));
    layer0_outputs(9370) <= (inputs(218)) xor (inputs(105));
    layer0_outputs(9371) <= not((inputs(62)) xor (inputs(66)));
    layer0_outputs(9372) <= inputs(87);
    layer0_outputs(9373) <= not((inputs(102)) or (inputs(23)));
    layer0_outputs(9374) <= not((inputs(66)) or (inputs(239)));
    layer0_outputs(9375) <= (inputs(215)) xor (inputs(220));
    layer0_outputs(9376) <= not(inputs(101)) or (inputs(98));
    layer0_outputs(9377) <= (inputs(167)) xor (inputs(237));
    layer0_outputs(9378) <= (inputs(249)) and not (inputs(144));
    layer0_outputs(9379) <= not(inputs(170));
    layer0_outputs(9380) <= not(inputs(134));
    layer0_outputs(9381) <= inputs(245);
    layer0_outputs(9382) <= (inputs(68)) and not (inputs(141));
    layer0_outputs(9383) <= (inputs(192)) and not (inputs(43));
    layer0_outputs(9384) <= not(inputs(41)) or (inputs(99));
    layer0_outputs(9385) <= not(inputs(138));
    layer0_outputs(9386) <= (inputs(188)) or (inputs(208));
    layer0_outputs(9387) <= inputs(227);
    layer0_outputs(9388) <= (inputs(14)) xor (inputs(186));
    layer0_outputs(9389) <= inputs(180);
    layer0_outputs(9390) <= inputs(131);
    layer0_outputs(9391) <= '1';
    layer0_outputs(9392) <= not(inputs(167));
    layer0_outputs(9393) <= not(inputs(106));
    layer0_outputs(9394) <= (inputs(210)) and not (inputs(4));
    layer0_outputs(9395) <= (inputs(24)) xor (inputs(115));
    layer0_outputs(9396) <= (inputs(66)) xor (inputs(3));
    layer0_outputs(9397) <= (inputs(24)) and not (inputs(17));
    layer0_outputs(9398) <= (inputs(12)) xor (inputs(150));
    layer0_outputs(9399) <= (inputs(14)) or (inputs(63));
    layer0_outputs(9400) <= not(inputs(13));
    layer0_outputs(9401) <= not((inputs(17)) or (inputs(200)));
    layer0_outputs(9402) <= inputs(217);
    layer0_outputs(9403) <= not(inputs(148)) or (inputs(195));
    layer0_outputs(9404) <= inputs(211);
    layer0_outputs(9405) <= (inputs(34)) xor (inputs(69));
    layer0_outputs(9406) <= not((inputs(215)) or (inputs(97)));
    layer0_outputs(9407) <= (inputs(118)) and not (inputs(229));
    layer0_outputs(9408) <= not((inputs(164)) xor (inputs(70)));
    layer0_outputs(9409) <= (inputs(201)) or (inputs(21));
    layer0_outputs(9410) <= (inputs(46)) and not (inputs(59));
    layer0_outputs(9411) <= inputs(234);
    layer0_outputs(9412) <= not(inputs(109));
    layer0_outputs(9413) <= not((inputs(38)) xor (inputs(103)));
    layer0_outputs(9414) <= (inputs(151)) xor (inputs(30));
    layer0_outputs(9415) <= not(inputs(122)) or (inputs(239));
    layer0_outputs(9416) <= inputs(121);
    layer0_outputs(9417) <= (inputs(185)) xor (inputs(156));
    layer0_outputs(9418) <= not(inputs(87));
    layer0_outputs(9419) <= (inputs(69)) and not (inputs(234));
    layer0_outputs(9420) <= inputs(252);
    layer0_outputs(9421) <= inputs(167);
    layer0_outputs(9422) <= not((inputs(165)) or (inputs(17)));
    layer0_outputs(9423) <= (inputs(87)) and not (inputs(253));
    layer0_outputs(9424) <= not(inputs(145)) or (inputs(250));
    layer0_outputs(9425) <= (inputs(198)) and not (inputs(44));
    layer0_outputs(9426) <= not((inputs(210)) xor (inputs(32)));
    layer0_outputs(9427) <= not((inputs(200)) or (inputs(233)));
    layer0_outputs(9428) <= not((inputs(220)) xor (inputs(190)));
    layer0_outputs(9429) <= inputs(205);
    layer0_outputs(9430) <= (inputs(55)) and not (inputs(190));
    layer0_outputs(9431) <= (inputs(64)) xor (inputs(215));
    layer0_outputs(9432) <= not(inputs(205));
    layer0_outputs(9433) <= (inputs(227)) or (inputs(128));
    layer0_outputs(9434) <= (inputs(199)) and not (inputs(231));
    layer0_outputs(9435) <= (inputs(184)) and not (inputs(230));
    layer0_outputs(9436) <= not(inputs(59)) or (inputs(21));
    layer0_outputs(9437) <= inputs(208);
    layer0_outputs(9438) <= (inputs(48)) or (inputs(172));
    layer0_outputs(9439) <= not((inputs(253)) and (inputs(111)));
    layer0_outputs(9440) <= not(inputs(225));
    layer0_outputs(9441) <= (inputs(197)) xor (inputs(120));
    layer0_outputs(9442) <= (inputs(51)) and (inputs(240));
    layer0_outputs(9443) <= not((inputs(58)) or (inputs(98)));
    layer0_outputs(9444) <= not(inputs(185));
    layer0_outputs(9445) <= (inputs(183)) xor (inputs(92));
    layer0_outputs(9446) <= (inputs(157)) or (inputs(181));
    layer0_outputs(9447) <= inputs(172);
    layer0_outputs(9448) <= inputs(123);
    layer0_outputs(9449) <= not(inputs(160)) or (inputs(198));
    layer0_outputs(9450) <= not((inputs(164)) or (inputs(149)));
    layer0_outputs(9451) <= not((inputs(194)) or (inputs(42)));
    layer0_outputs(9452) <= (inputs(243)) xor (inputs(228));
    layer0_outputs(9453) <= not(inputs(103));
    layer0_outputs(9454) <= (inputs(200)) and not (inputs(64));
    layer0_outputs(9455) <= inputs(53);
    layer0_outputs(9456) <= not((inputs(230)) xor (inputs(144)));
    layer0_outputs(9457) <= (inputs(214)) or (inputs(106));
    layer0_outputs(9458) <= '1';
    layer0_outputs(9459) <= '0';
    layer0_outputs(9460) <= (inputs(103)) and not (inputs(26));
    layer0_outputs(9461) <= not(inputs(60)) or (inputs(33));
    layer0_outputs(9462) <= '1';
    layer0_outputs(9463) <= not(inputs(155));
    layer0_outputs(9464) <= not((inputs(206)) or (inputs(68)));
    layer0_outputs(9465) <= inputs(171);
    layer0_outputs(9466) <= (inputs(80)) or (inputs(226));
    layer0_outputs(9467) <= not(inputs(51)) or (inputs(108));
    layer0_outputs(9468) <= not((inputs(129)) xor (inputs(53)));
    layer0_outputs(9469) <= (inputs(222)) or (inputs(38));
    layer0_outputs(9470) <= not((inputs(91)) xor (inputs(21)));
    layer0_outputs(9471) <= (inputs(245)) or (inputs(205));
    layer0_outputs(9472) <= not((inputs(158)) and (inputs(24)));
    layer0_outputs(9473) <= not((inputs(63)) or (inputs(142)));
    layer0_outputs(9474) <= not(inputs(112));
    layer0_outputs(9475) <= inputs(227);
    layer0_outputs(9476) <= inputs(199);
    layer0_outputs(9477) <= (inputs(106)) and not (inputs(82));
    layer0_outputs(9478) <= not(inputs(80)) or (inputs(169));
    layer0_outputs(9479) <= (inputs(36)) xor (inputs(215));
    layer0_outputs(9480) <= (inputs(242)) xor (inputs(129));
    layer0_outputs(9481) <= inputs(24);
    layer0_outputs(9482) <= not(inputs(3)) or (inputs(15));
    layer0_outputs(9483) <= (inputs(143)) or (inputs(76));
    layer0_outputs(9484) <= (inputs(144)) and (inputs(148));
    layer0_outputs(9485) <= '1';
    layer0_outputs(9486) <= (inputs(198)) xor (inputs(30));
    layer0_outputs(9487) <= not(inputs(20));
    layer0_outputs(9488) <= not((inputs(70)) or (inputs(112)));
    layer0_outputs(9489) <= not(inputs(199));
    layer0_outputs(9490) <= (inputs(209)) or (inputs(41));
    layer0_outputs(9491) <= not(inputs(138));
    layer0_outputs(9492) <= not(inputs(87));
    layer0_outputs(9493) <= not((inputs(72)) or (inputs(63)));
    layer0_outputs(9494) <= (inputs(153)) or (inputs(108));
    layer0_outputs(9495) <= not((inputs(199)) or (inputs(194)));
    layer0_outputs(9496) <= (inputs(247)) or (inputs(103));
    layer0_outputs(9497) <= not((inputs(45)) or (inputs(177)));
    layer0_outputs(9498) <= not((inputs(34)) and (inputs(244)));
    layer0_outputs(9499) <= not((inputs(178)) xor (inputs(136)));
    layer0_outputs(9500) <= not((inputs(25)) or (inputs(178)));
    layer0_outputs(9501) <= inputs(208);
    layer0_outputs(9502) <= not((inputs(116)) or (inputs(42)));
    layer0_outputs(9503) <= (inputs(31)) or (inputs(183));
    layer0_outputs(9504) <= '1';
    layer0_outputs(9505) <= inputs(26);
    layer0_outputs(9506) <= inputs(109);
    layer0_outputs(9507) <= not(inputs(153)) or (inputs(26));
    layer0_outputs(9508) <= (inputs(164)) xor (inputs(227));
    layer0_outputs(9509) <= inputs(216);
    layer0_outputs(9510) <= not(inputs(214)) or (inputs(111));
    layer0_outputs(9511) <= not(inputs(206)) or (inputs(184));
    layer0_outputs(9512) <= not(inputs(24)) or (inputs(144));
    layer0_outputs(9513) <= (inputs(35)) xor (inputs(82));
    layer0_outputs(9514) <= (inputs(253)) xor (inputs(233));
    layer0_outputs(9515) <= not((inputs(120)) or (inputs(83)));
    layer0_outputs(9516) <= (inputs(148)) and not (inputs(88));
    layer0_outputs(9517) <= inputs(150);
    layer0_outputs(9518) <= (inputs(56)) and not (inputs(209));
    layer0_outputs(9519) <= inputs(28);
    layer0_outputs(9520) <= not(inputs(164)) or (inputs(236));
    layer0_outputs(9521) <= (inputs(140)) and not (inputs(17));
    layer0_outputs(9522) <= not(inputs(214)) or (inputs(29));
    layer0_outputs(9523) <= inputs(56);
    layer0_outputs(9524) <= (inputs(89)) and not (inputs(237));
    layer0_outputs(9525) <= not((inputs(237)) xor (inputs(187)));
    layer0_outputs(9526) <= (inputs(121)) and not (inputs(188));
    layer0_outputs(9527) <= not((inputs(231)) xor (inputs(233)));
    layer0_outputs(9528) <= not((inputs(70)) or (inputs(179)));
    layer0_outputs(9529) <= not(inputs(79)) or (inputs(178));
    layer0_outputs(9530) <= not((inputs(102)) and (inputs(199)));
    layer0_outputs(9531) <= (inputs(25)) xor (inputs(210));
    layer0_outputs(9532) <= (inputs(195)) or (inputs(236));
    layer0_outputs(9533) <= (inputs(153)) or (inputs(49));
    layer0_outputs(9534) <= (inputs(61)) or (inputs(194));
    layer0_outputs(9535) <= not(inputs(28));
    layer0_outputs(9536) <= (inputs(82)) xor (inputs(189));
    layer0_outputs(9537) <= not((inputs(6)) or (inputs(75)));
    layer0_outputs(9538) <= (inputs(45)) and not (inputs(254));
    layer0_outputs(9539) <= (inputs(230)) xor (inputs(44));
    layer0_outputs(9540) <= '1';
    layer0_outputs(9541) <= '1';
    layer0_outputs(9542) <= not(inputs(118)) or (inputs(224));
    layer0_outputs(9543) <= inputs(27);
    layer0_outputs(9544) <= (inputs(141)) and not (inputs(194));
    layer0_outputs(9545) <= not(inputs(196)) or (inputs(52));
    layer0_outputs(9546) <= not((inputs(218)) xor (inputs(199)));
    layer0_outputs(9547) <= not((inputs(237)) or (inputs(122)));
    layer0_outputs(9548) <= not((inputs(98)) xor (inputs(30)));
    layer0_outputs(9549) <= not((inputs(250)) or (inputs(62)));
    layer0_outputs(9550) <= not((inputs(243)) xor (inputs(23)));
    layer0_outputs(9551) <= not(inputs(248)) or (inputs(62));
    layer0_outputs(9552) <= not(inputs(96));
    layer0_outputs(9553) <= not((inputs(225)) or (inputs(95)));
    layer0_outputs(9554) <= not((inputs(103)) or (inputs(197)));
    layer0_outputs(9555) <= not(inputs(86)) or (inputs(79));
    layer0_outputs(9556) <= not(inputs(216));
    layer0_outputs(9557) <= not((inputs(41)) xor (inputs(62)));
    layer0_outputs(9558) <= (inputs(24)) and (inputs(78));
    layer0_outputs(9559) <= (inputs(183)) xor (inputs(210));
    layer0_outputs(9560) <= (inputs(176)) or (inputs(16));
    layer0_outputs(9561) <= inputs(174);
    layer0_outputs(9562) <= not(inputs(202)) or (inputs(237));
    layer0_outputs(9563) <= not(inputs(205)) or (inputs(80));
    layer0_outputs(9564) <= not(inputs(139));
    layer0_outputs(9565) <= (inputs(200)) and not (inputs(239));
    layer0_outputs(9566) <= not(inputs(66));
    layer0_outputs(9567) <= (inputs(187)) or (inputs(162));
    layer0_outputs(9568) <= (inputs(234)) or (inputs(241));
    layer0_outputs(9569) <= inputs(200);
    layer0_outputs(9570) <= not((inputs(148)) or (inputs(87)));
    layer0_outputs(9571) <= (inputs(82)) and not (inputs(192));
    layer0_outputs(9572) <= not((inputs(88)) and (inputs(130)));
    layer0_outputs(9573) <= not((inputs(132)) xor (inputs(83)));
    layer0_outputs(9574) <= not(inputs(105)) or (inputs(11));
    layer0_outputs(9575) <= (inputs(91)) xor (inputs(41));
    layer0_outputs(9576) <= not(inputs(101)) or (inputs(234));
    layer0_outputs(9577) <= not(inputs(241));
    layer0_outputs(9578) <= not((inputs(237)) and (inputs(45)));
    layer0_outputs(9579) <= not((inputs(94)) or (inputs(19)));
    layer0_outputs(9580) <= (inputs(11)) and (inputs(234));
    layer0_outputs(9581) <= not(inputs(182));
    layer0_outputs(9582) <= (inputs(244)) and not (inputs(13));
    layer0_outputs(9583) <= not((inputs(53)) or (inputs(13)));
    layer0_outputs(9584) <= '0';
    layer0_outputs(9585) <= (inputs(102)) and not (inputs(226));
    layer0_outputs(9586) <= (inputs(203)) or (inputs(93));
    layer0_outputs(9587) <= (inputs(165)) xor (inputs(236));
    layer0_outputs(9588) <= not((inputs(141)) or (inputs(131)));
    layer0_outputs(9589) <= (inputs(221)) or (inputs(176));
    layer0_outputs(9590) <= not((inputs(189)) xor (inputs(123)));
    layer0_outputs(9591) <= (inputs(244)) and not (inputs(130));
    layer0_outputs(9592) <= (inputs(101)) and not (inputs(251));
    layer0_outputs(9593) <= (inputs(165)) or (inputs(150));
    layer0_outputs(9594) <= (inputs(132)) and not (inputs(21));
    layer0_outputs(9595) <= not(inputs(86));
    layer0_outputs(9596) <= inputs(237);
    layer0_outputs(9597) <= not((inputs(14)) and (inputs(157)));
    layer0_outputs(9598) <= (inputs(218)) xor (inputs(57));
    layer0_outputs(9599) <= (inputs(151)) xor (inputs(66));
    layer0_outputs(9600) <= inputs(150);
    layer0_outputs(9601) <= not(inputs(208));
    layer0_outputs(9602) <= (inputs(224)) xor (inputs(252));
    layer0_outputs(9603) <= (inputs(168)) and not (inputs(212));
    layer0_outputs(9604) <= not(inputs(212)) or (inputs(208));
    layer0_outputs(9605) <= not((inputs(211)) xor (inputs(39)));
    layer0_outputs(9606) <= not((inputs(150)) xor (inputs(90)));
    layer0_outputs(9607) <= not(inputs(10)) or (inputs(93));
    layer0_outputs(9608) <= (inputs(158)) and not (inputs(158));
    layer0_outputs(9609) <= not((inputs(46)) and (inputs(113)));
    layer0_outputs(9610) <= inputs(180);
    layer0_outputs(9611) <= not((inputs(44)) xor (inputs(77)));
    layer0_outputs(9612) <= (inputs(158)) or (inputs(180));
    layer0_outputs(9613) <= (inputs(138)) or (inputs(237));
    layer0_outputs(9614) <= (inputs(4)) xor (inputs(166));
    layer0_outputs(9615) <= (inputs(205)) and (inputs(237));
    layer0_outputs(9616) <= not(inputs(133));
    layer0_outputs(9617) <= (inputs(113)) or (inputs(125));
    layer0_outputs(9618) <= not((inputs(166)) or (inputs(142)));
    layer0_outputs(9619) <= inputs(40);
    layer0_outputs(9620) <= (inputs(8)) or (inputs(103));
    layer0_outputs(9621) <= not((inputs(80)) and (inputs(44)));
    layer0_outputs(9622) <= (inputs(193)) and not (inputs(183));
    layer0_outputs(9623) <= (inputs(83)) xor (inputs(220));
    layer0_outputs(9624) <= (inputs(103)) and not (inputs(231));
    layer0_outputs(9625) <= (inputs(157)) or (inputs(191));
    layer0_outputs(9626) <= not((inputs(179)) or (inputs(162)));
    layer0_outputs(9627) <= (inputs(213)) or (inputs(174));
    layer0_outputs(9628) <= (inputs(109)) xor (inputs(144));
    layer0_outputs(9629) <= inputs(158);
    layer0_outputs(9630) <= (inputs(64)) xor (inputs(109));
    layer0_outputs(9631) <= not((inputs(207)) and (inputs(216)));
    layer0_outputs(9632) <= inputs(171);
    layer0_outputs(9633) <= (inputs(223)) or (inputs(156));
    layer0_outputs(9634) <= (inputs(54)) or (inputs(247));
    layer0_outputs(9635) <= not((inputs(185)) or (inputs(171)));
    layer0_outputs(9636) <= inputs(160);
    layer0_outputs(9637) <= not((inputs(253)) and (inputs(126)));
    layer0_outputs(9638) <= not(inputs(38)) or (inputs(236));
    layer0_outputs(9639) <= (inputs(144)) and (inputs(52));
    layer0_outputs(9640) <= not((inputs(114)) or (inputs(51)));
    layer0_outputs(9641) <= not(inputs(215));
    layer0_outputs(9642) <= (inputs(47)) or (inputs(97));
    layer0_outputs(9643) <= not(inputs(137));
    layer0_outputs(9644) <= (inputs(17)) and not (inputs(17));
    layer0_outputs(9645) <= not((inputs(173)) or (inputs(171)));
    layer0_outputs(9646) <= (inputs(130)) and not (inputs(62));
    layer0_outputs(9647) <= not(inputs(79));
    layer0_outputs(9648) <= not((inputs(144)) and (inputs(130)));
    layer0_outputs(9649) <= not(inputs(106)) or (inputs(59));
    layer0_outputs(9650) <= inputs(171);
    layer0_outputs(9651) <= inputs(162);
    layer0_outputs(9652) <= (inputs(166)) and not (inputs(226));
    layer0_outputs(9653) <= '0';
    layer0_outputs(9654) <= (inputs(6)) xor (inputs(0));
    layer0_outputs(9655) <= inputs(107);
    layer0_outputs(9656) <= (inputs(48)) or (inputs(102));
    layer0_outputs(9657) <= not(inputs(198)) or (inputs(189));
    layer0_outputs(9658) <= not(inputs(225)) or (inputs(169));
    layer0_outputs(9659) <= inputs(186);
    layer0_outputs(9660) <= (inputs(90)) and not (inputs(249));
    layer0_outputs(9661) <= not((inputs(94)) xor (inputs(200)));
    layer0_outputs(9662) <= not((inputs(255)) xor (inputs(70)));
    layer0_outputs(9663) <= not((inputs(68)) xor (inputs(170)));
    layer0_outputs(9664) <= (inputs(81)) and not (inputs(254));
    layer0_outputs(9665) <= not((inputs(53)) xor (inputs(144)));
    layer0_outputs(9666) <= (inputs(252)) and not (inputs(7));
    layer0_outputs(9667) <= inputs(106);
    layer0_outputs(9668) <= not(inputs(15));
    layer0_outputs(9669) <= not((inputs(136)) and (inputs(65)));
    layer0_outputs(9670) <= (inputs(51)) and (inputs(27));
    layer0_outputs(9671) <= not((inputs(40)) or (inputs(56)));
    layer0_outputs(9672) <= (inputs(126)) and not (inputs(221));
    layer0_outputs(9673) <= not(inputs(197));
    layer0_outputs(9674) <= not(inputs(39));
    layer0_outputs(9675) <= not(inputs(113)) or (inputs(160));
    layer0_outputs(9676) <= not(inputs(79));
    layer0_outputs(9677) <= not((inputs(249)) or (inputs(168)));
    layer0_outputs(9678) <= not(inputs(197)) or (inputs(210));
    layer0_outputs(9679) <= not(inputs(13)) or (inputs(86));
    layer0_outputs(9680) <= (inputs(24)) and not (inputs(241));
    layer0_outputs(9681) <= not((inputs(216)) or (inputs(249)));
    layer0_outputs(9682) <= not((inputs(244)) xor (inputs(105)));
    layer0_outputs(9683) <= not(inputs(153)) or (inputs(166));
    layer0_outputs(9684) <= (inputs(184)) and not (inputs(78));
    layer0_outputs(9685) <= not(inputs(139));
    layer0_outputs(9686) <= '0';
    layer0_outputs(9687) <= (inputs(74)) xor (inputs(123));
    layer0_outputs(9688) <= not(inputs(173));
    layer0_outputs(9689) <= '0';
    layer0_outputs(9690) <= not(inputs(94));
    layer0_outputs(9691) <= (inputs(4)) or (inputs(133));
    layer0_outputs(9692) <= inputs(230);
    layer0_outputs(9693) <= not(inputs(229)) or (inputs(202));
    layer0_outputs(9694) <= not(inputs(149)) or (inputs(57));
    layer0_outputs(9695) <= not((inputs(48)) or (inputs(215)));
    layer0_outputs(9696) <= inputs(216);
    layer0_outputs(9697) <= not((inputs(50)) or (inputs(170)));
    layer0_outputs(9698) <= (inputs(180)) and not (inputs(235));
    layer0_outputs(9699) <= (inputs(107)) xor (inputs(13));
    layer0_outputs(9700) <= not(inputs(229)) or (inputs(243));
    layer0_outputs(9701) <= not(inputs(120));
    layer0_outputs(9702) <= '1';
    layer0_outputs(9703) <= (inputs(148)) and not (inputs(231));
    layer0_outputs(9704) <= not(inputs(119)) or (inputs(190));
    layer0_outputs(9705) <= not(inputs(65)) or (inputs(106));
    layer0_outputs(9706) <= (inputs(107)) and not (inputs(22));
    layer0_outputs(9707) <= not(inputs(62)) or (inputs(209));
    layer0_outputs(9708) <= (inputs(212)) xor (inputs(105));
    layer0_outputs(9709) <= (inputs(181)) or (inputs(58));
    layer0_outputs(9710) <= not(inputs(103)) or (inputs(127));
    layer0_outputs(9711) <= not((inputs(166)) or (inputs(97)));
    layer0_outputs(9712) <= (inputs(170)) or (inputs(188));
    layer0_outputs(9713) <= not((inputs(82)) xor (inputs(5)));
    layer0_outputs(9714) <= not((inputs(133)) or (inputs(214)));
    layer0_outputs(9715) <= (inputs(27)) or (inputs(41));
    layer0_outputs(9716) <= not((inputs(134)) or (inputs(148)));
    layer0_outputs(9717) <= (inputs(54)) xor (inputs(42));
    layer0_outputs(9718) <= not(inputs(138));
    layer0_outputs(9719) <= not(inputs(211)) or (inputs(15));
    layer0_outputs(9720) <= not((inputs(169)) xor (inputs(43)));
    layer0_outputs(9721) <= not((inputs(237)) xor (inputs(83)));
    layer0_outputs(9722) <= not(inputs(165)) or (inputs(129));
    layer0_outputs(9723) <= (inputs(139)) or (inputs(50));
    layer0_outputs(9724) <= not((inputs(136)) or (inputs(112)));
    layer0_outputs(9725) <= (inputs(40)) or (inputs(136));
    layer0_outputs(9726) <= not(inputs(229));
    layer0_outputs(9727) <= not(inputs(147));
    layer0_outputs(9728) <= not((inputs(145)) xor (inputs(61)));
    layer0_outputs(9729) <= not(inputs(22));
    layer0_outputs(9730) <= not((inputs(69)) xor (inputs(250)));
    layer0_outputs(9731) <= not(inputs(194)) or (inputs(75));
    layer0_outputs(9732) <= not(inputs(254));
    layer0_outputs(9733) <= not((inputs(223)) and (inputs(108)));
    layer0_outputs(9734) <= (inputs(254)) xor (inputs(221));
    layer0_outputs(9735) <= (inputs(41)) xor (inputs(57));
    layer0_outputs(9736) <= (inputs(18)) and not (inputs(65));
    layer0_outputs(9737) <= not(inputs(121)) or (inputs(179));
    layer0_outputs(9738) <= not((inputs(29)) and (inputs(142)));
    layer0_outputs(9739) <= (inputs(122)) and not (inputs(137));
    layer0_outputs(9740) <= not(inputs(85)) or (inputs(45));
    layer0_outputs(9741) <= inputs(192);
    layer0_outputs(9742) <= (inputs(129)) and (inputs(34));
    layer0_outputs(9743) <= (inputs(33)) xor (inputs(206));
    layer0_outputs(9744) <= not((inputs(54)) or (inputs(178)));
    layer0_outputs(9745) <= not(inputs(103)) or (inputs(112));
    layer0_outputs(9746) <= not(inputs(37));
    layer0_outputs(9747) <= (inputs(57)) xor (inputs(46));
    layer0_outputs(9748) <= inputs(181);
    layer0_outputs(9749) <= (inputs(33)) and not (inputs(158));
    layer0_outputs(9750) <= not(inputs(108));
    layer0_outputs(9751) <= not((inputs(75)) and (inputs(43)));
    layer0_outputs(9752) <= not(inputs(229));
    layer0_outputs(9753) <= not((inputs(64)) or (inputs(38)));
    layer0_outputs(9754) <= not((inputs(191)) xor (inputs(60)));
    layer0_outputs(9755) <= inputs(43);
    layer0_outputs(9756) <= inputs(141);
    layer0_outputs(9757) <= not(inputs(63));
    layer0_outputs(9758) <= not(inputs(220)) or (inputs(247));
    layer0_outputs(9759) <= (inputs(45)) and not (inputs(234));
    layer0_outputs(9760) <= '0';
    layer0_outputs(9761) <= inputs(189);
    layer0_outputs(9762) <= (inputs(217)) and not (inputs(81));
    layer0_outputs(9763) <= not(inputs(113));
    layer0_outputs(9764) <= '1';
    layer0_outputs(9765) <= (inputs(232)) or (inputs(111));
    layer0_outputs(9766) <= (inputs(229)) and not (inputs(20));
    layer0_outputs(9767) <= inputs(183);
    layer0_outputs(9768) <= inputs(65);
    layer0_outputs(9769) <= (inputs(52)) xor (inputs(161));
    layer0_outputs(9770) <= not(inputs(212)) or (inputs(141));
    layer0_outputs(9771) <= not((inputs(29)) or (inputs(230)));
    layer0_outputs(9772) <= (inputs(84)) and not (inputs(79));
    layer0_outputs(9773) <= inputs(255);
    layer0_outputs(9774) <= not(inputs(111));
    layer0_outputs(9775) <= not(inputs(100));
    layer0_outputs(9776) <= (inputs(149)) or (inputs(172));
    layer0_outputs(9777) <= not(inputs(42)) or (inputs(31));
    layer0_outputs(9778) <= not((inputs(197)) xor (inputs(187)));
    layer0_outputs(9779) <= not((inputs(189)) or (inputs(222)));
    layer0_outputs(9780) <= (inputs(206)) xor (inputs(8));
    layer0_outputs(9781) <= not(inputs(161)) or (inputs(11));
    layer0_outputs(9782) <= (inputs(85)) and not (inputs(185));
    layer0_outputs(9783) <= not(inputs(194)) or (inputs(161));
    layer0_outputs(9784) <= (inputs(28)) xor (inputs(33));
    layer0_outputs(9785) <= inputs(103);
    layer0_outputs(9786) <= (inputs(98)) and not (inputs(238));
    layer0_outputs(9787) <= (inputs(75)) or (inputs(15));
    layer0_outputs(9788) <= (inputs(118)) or (inputs(79));
    layer0_outputs(9789) <= not(inputs(201));
    layer0_outputs(9790) <= (inputs(63)) and not (inputs(112));
    layer0_outputs(9791) <= (inputs(166)) and not (inputs(34));
    layer0_outputs(9792) <= (inputs(21)) and not (inputs(91));
    layer0_outputs(9793) <= not((inputs(151)) or (inputs(248)));
    layer0_outputs(9794) <= not(inputs(156)) or (inputs(240));
    layer0_outputs(9795) <= not((inputs(186)) or (inputs(40)));
    layer0_outputs(9796) <= (inputs(69)) xor (inputs(202));
    layer0_outputs(9797) <= inputs(102);
    layer0_outputs(9798) <= not(inputs(195));
    layer0_outputs(9799) <= (inputs(155)) xor (inputs(131));
    layer0_outputs(9800) <= not((inputs(77)) xor (inputs(222)));
    layer0_outputs(9801) <= (inputs(60)) or (inputs(117));
    layer0_outputs(9802) <= not(inputs(136));
    layer0_outputs(9803) <= (inputs(197)) and (inputs(48));
    layer0_outputs(9804) <= not(inputs(139));
    layer0_outputs(9805) <= (inputs(173)) and (inputs(132));
    layer0_outputs(9806) <= (inputs(57)) and not (inputs(195));
    layer0_outputs(9807) <= (inputs(170)) and not (inputs(114));
    layer0_outputs(9808) <= (inputs(32)) or (inputs(114));
    layer0_outputs(9809) <= (inputs(208)) xor (inputs(47));
    layer0_outputs(9810) <= not(inputs(206));
    layer0_outputs(9811) <= not((inputs(189)) xor (inputs(23)));
    layer0_outputs(9812) <= not(inputs(94)) or (inputs(130));
    layer0_outputs(9813) <= '1';
    layer0_outputs(9814) <= inputs(181);
    layer0_outputs(9815) <= not((inputs(121)) xor (inputs(154)));
    layer0_outputs(9816) <= not(inputs(104)) or (inputs(164));
    layer0_outputs(9817) <= (inputs(232)) or (inputs(124));
    layer0_outputs(9818) <= (inputs(32)) or (inputs(175));
    layer0_outputs(9819) <= not(inputs(155));
    layer0_outputs(9820) <= not((inputs(232)) xor (inputs(5)));
    layer0_outputs(9821) <= not((inputs(154)) or (inputs(22)));
    layer0_outputs(9822) <= (inputs(228)) and not (inputs(206));
    layer0_outputs(9823) <= inputs(201);
    layer0_outputs(9824) <= not(inputs(44)) or (inputs(112));
    layer0_outputs(9825) <= (inputs(102)) or (inputs(44));
    layer0_outputs(9826) <= (inputs(88)) and not (inputs(82));
    layer0_outputs(9827) <= not(inputs(42)) or (inputs(75));
    layer0_outputs(9828) <= not(inputs(90)) or (inputs(163));
    layer0_outputs(9829) <= (inputs(39)) and not (inputs(95));
    layer0_outputs(9830) <= (inputs(168)) and not (inputs(28));
    layer0_outputs(9831) <= not(inputs(230));
    layer0_outputs(9832) <= not(inputs(182));
    layer0_outputs(9833) <= (inputs(1)) or (inputs(149));
    layer0_outputs(9834) <= '0';
    layer0_outputs(9835) <= not(inputs(100));
    layer0_outputs(9836) <= (inputs(166)) and not (inputs(98));
    layer0_outputs(9837) <= not((inputs(42)) or (inputs(84)));
    layer0_outputs(9838) <= not((inputs(136)) or (inputs(124)));
    layer0_outputs(9839) <= not(inputs(89)) or (inputs(33));
    layer0_outputs(9840) <= inputs(249);
    layer0_outputs(9841) <= not((inputs(35)) or (inputs(54)));
    layer0_outputs(9842) <= (inputs(54)) xor (inputs(140));
    layer0_outputs(9843) <= (inputs(129)) and not (inputs(22));
    layer0_outputs(9844) <= not((inputs(63)) or (inputs(90)));
    layer0_outputs(9845) <= not((inputs(63)) xor (inputs(14)));
    layer0_outputs(9846) <= not(inputs(1)) or (inputs(35));
    layer0_outputs(9847) <= not((inputs(241)) or (inputs(137)));
    layer0_outputs(9848) <= inputs(220);
    layer0_outputs(9849) <= not(inputs(181));
    layer0_outputs(9850) <= not((inputs(46)) xor (inputs(88)));
    layer0_outputs(9851) <= not((inputs(130)) or (inputs(117)));
    layer0_outputs(9852) <= not((inputs(232)) or (inputs(24)));
    layer0_outputs(9853) <= (inputs(139)) and not (inputs(244));
    layer0_outputs(9854) <= not((inputs(197)) and (inputs(192)));
    layer0_outputs(9855) <= not((inputs(192)) xor (inputs(226)));
    layer0_outputs(9856) <= (inputs(231)) and not (inputs(173));
    layer0_outputs(9857) <= inputs(253);
    layer0_outputs(9858) <= (inputs(249)) or (inputs(67));
    layer0_outputs(9859) <= not(inputs(164)) or (inputs(145));
    layer0_outputs(9860) <= (inputs(8)) and not (inputs(62));
    layer0_outputs(9861) <= (inputs(229)) or (inputs(190));
    layer0_outputs(9862) <= (inputs(115)) or (inputs(212));
    layer0_outputs(9863) <= (inputs(0)) and not (inputs(86));
    layer0_outputs(9864) <= (inputs(205)) xor (inputs(45));
    layer0_outputs(9865) <= inputs(140);
    layer0_outputs(9866) <= not((inputs(185)) or (inputs(28)));
    layer0_outputs(9867) <= (inputs(70)) xor (inputs(205));
    layer0_outputs(9868) <= inputs(73);
    layer0_outputs(9869) <= inputs(171);
    layer0_outputs(9870) <= not(inputs(199)) or (inputs(114));
    layer0_outputs(9871) <= not((inputs(164)) or (inputs(78)));
    layer0_outputs(9872) <= not(inputs(215));
    layer0_outputs(9873) <= not((inputs(215)) and (inputs(5)));
    layer0_outputs(9874) <= not((inputs(197)) or (inputs(93)));
    layer0_outputs(9875) <= not((inputs(202)) or (inputs(146)));
    layer0_outputs(9876) <= not(inputs(135)) or (inputs(10));
    layer0_outputs(9877) <= not(inputs(90)) or (inputs(125));
    layer0_outputs(9878) <= (inputs(172)) xor (inputs(18));
    layer0_outputs(9879) <= not((inputs(65)) or (inputs(211)));
    layer0_outputs(9880) <= (inputs(201)) and not (inputs(225));
    layer0_outputs(9881) <= (inputs(90)) or (inputs(74));
    layer0_outputs(9882) <= (inputs(60)) or (inputs(100));
    layer0_outputs(9883) <= not((inputs(197)) xor (inputs(189)));
    layer0_outputs(9884) <= not(inputs(61));
    layer0_outputs(9885) <= not(inputs(172));
    layer0_outputs(9886) <= inputs(165);
    layer0_outputs(9887) <= not((inputs(14)) or (inputs(146)));
    layer0_outputs(9888) <= (inputs(159)) xor (inputs(156));
    layer0_outputs(9889) <= not((inputs(231)) xor (inputs(212)));
    layer0_outputs(9890) <= not(inputs(182)) or (inputs(77));
    layer0_outputs(9891) <= not(inputs(19));
    layer0_outputs(9892) <= (inputs(147)) or (inputs(83));
    layer0_outputs(9893) <= not(inputs(50));
    layer0_outputs(9894) <= not(inputs(151)) or (inputs(10));
    layer0_outputs(9895) <= (inputs(99)) and not (inputs(248));
    layer0_outputs(9896) <= (inputs(160)) and not (inputs(238));
    layer0_outputs(9897) <= (inputs(30)) xor (inputs(27));
    layer0_outputs(9898) <= inputs(188);
    layer0_outputs(9899) <= (inputs(121)) and not (inputs(9));
    layer0_outputs(9900) <= (inputs(136)) and not (inputs(174));
    layer0_outputs(9901) <= (inputs(217)) and not (inputs(114));
    layer0_outputs(9902) <= not(inputs(146));
    layer0_outputs(9903) <= (inputs(196)) or (inputs(146));
    layer0_outputs(9904) <= (inputs(144)) xor (inputs(154));
    layer0_outputs(9905) <= inputs(15);
    layer0_outputs(9906) <= not(inputs(28));
    layer0_outputs(9907) <= inputs(175);
    layer0_outputs(9908) <= not(inputs(175));
    layer0_outputs(9909) <= (inputs(233)) and (inputs(134));
    layer0_outputs(9910) <= not((inputs(218)) or (inputs(31)));
    layer0_outputs(9911) <= not(inputs(105));
    layer0_outputs(9912) <= not((inputs(166)) or (inputs(186)));
    layer0_outputs(9913) <= not(inputs(14));
    layer0_outputs(9914) <= not(inputs(56)) or (inputs(139));
    layer0_outputs(9915) <= not((inputs(57)) or (inputs(132)));
    layer0_outputs(9916) <= (inputs(188)) and not (inputs(23));
    layer0_outputs(9917) <= not(inputs(56));
    layer0_outputs(9918) <= (inputs(90)) and not (inputs(193));
    layer0_outputs(9919) <= not((inputs(67)) and (inputs(89)));
    layer0_outputs(9920) <= not(inputs(149));
    layer0_outputs(9921) <= inputs(92);
    layer0_outputs(9922) <= (inputs(13)) or (inputs(146));
    layer0_outputs(9923) <= not(inputs(50)) or (inputs(226));
    layer0_outputs(9924) <= not(inputs(125));
    layer0_outputs(9925) <= not(inputs(103)) or (inputs(1));
    layer0_outputs(9926) <= (inputs(142)) and not (inputs(142));
    layer0_outputs(9927) <= inputs(223);
    layer0_outputs(9928) <= (inputs(253)) and not (inputs(227));
    layer0_outputs(9929) <= (inputs(191)) or (inputs(151));
    layer0_outputs(9930) <= not((inputs(174)) or (inputs(180)));
    layer0_outputs(9931) <= not((inputs(157)) and (inputs(184)));
    layer0_outputs(9932) <= not(inputs(57)) or (inputs(145));
    layer0_outputs(9933) <= (inputs(91)) and not (inputs(131));
    layer0_outputs(9934) <= (inputs(148)) or (inputs(142));
    layer0_outputs(9935) <= not(inputs(247)) or (inputs(47));
    layer0_outputs(9936) <= (inputs(6)) xor (inputs(42));
    layer0_outputs(9937) <= inputs(227);
    layer0_outputs(9938) <= (inputs(206)) and not (inputs(219));
    layer0_outputs(9939) <= inputs(216);
    layer0_outputs(9940) <= not(inputs(231));
    layer0_outputs(9941) <= '0';
    layer0_outputs(9942) <= (inputs(208)) and not (inputs(128));
    layer0_outputs(9943) <= inputs(144);
    layer0_outputs(9944) <= not(inputs(214)) or (inputs(102));
    layer0_outputs(9945) <= (inputs(17)) xor (inputs(135));
    layer0_outputs(9946) <= not(inputs(10)) or (inputs(235));
    layer0_outputs(9947) <= not(inputs(101)) or (inputs(233));
    layer0_outputs(9948) <= '0';
    layer0_outputs(9949) <= (inputs(64)) and not (inputs(43));
    layer0_outputs(9950) <= (inputs(248)) and not (inputs(176));
    layer0_outputs(9951) <= (inputs(239)) or (inputs(148));
    layer0_outputs(9952) <= (inputs(118)) and not (inputs(127));
    layer0_outputs(9953) <= not(inputs(62)) or (inputs(157));
    layer0_outputs(9954) <= (inputs(65)) or (inputs(58));
    layer0_outputs(9955) <= not((inputs(159)) or (inputs(77)));
    layer0_outputs(9956) <= not(inputs(152)) or (inputs(18));
    layer0_outputs(9957) <= not(inputs(179));
    layer0_outputs(9958) <= (inputs(41)) xor (inputs(72));
    layer0_outputs(9959) <= (inputs(191)) or (inputs(12));
    layer0_outputs(9960) <= not(inputs(30)) or (inputs(10));
    layer0_outputs(9961) <= '0';
    layer0_outputs(9962) <= not(inputs(84)) or (inputs(230));
    layer0_outputs(9963) <= not(inputs(38)) or (inputs(237));
    layer0_outputs(9964) <= inputs(170);
    layer0_outputs(9965) <= inputs(180);
    layer0_outputs(9966) <= '1';
    layer0_outputs(9967) <= (inputs(138)) or (inputs(85));
    layer0_outputs(9968) <= not(inputs(135));
    layer0_outputs(9969) <= not((inputs(83)) or (inputs(174)));
    layer0_outputs(9970) <= (inputs(52)) and not (inputs(255));
    layer0_outputs(9971) <= not(inputs(121)) or (inputs(189));
    layer0_outputs(9972) <= not((inputs(100)) or (inputs(150)));
    layer0_outputs(9973) <= not((inputs(45)) and (inputs(37)));
    layer0_outputs(9974) <= not(inputs(160));
    layer0_outputs(9975) <= inputs(164);
    layer0_outputs(9976) <= not(inputs(162));
    layer0_outputs(9977) <= not((inputs(213)) or (inputs(160)));
    layer0_outputs(9978) <= not((inputs(211)) or (inputs(186)));
    layer0_outputs(9979) <= (inputs(189)) and not (inputs(50));
    layer0_outputs(9980) <= (inputs(232)) or (inputs(104));
    layer0_outputs(9981) <= not(inputs(199));
    layer0_outputs(9982) <= not((inputs(195)) xor (inputs(220)));
    layer0_outputs(9983) <= not(inputs(178)) or (inputs(245));
    layer0_outputs(9984) <= (inputs(139)) and not (inputs(248));
    layer0_outputs(9985) <= (inputs(60)) and not (inputs(249));
    layer0_outputs(9986) <= not(inputs(240));
    layer0_outputs(9987) <= (inputs(157)) xor (inputs(186));
    layer0_outputs(9988) <= not(inputs(231));
    layer0_outputs(9989) <= not(inputs(181));
    layer0_outputs(9990) <= (inputs(71)) and not (inputs(191));
    layer0_outputs(9991) <= (inputs(142)) xor (inputs(166));
    layer0_outputs(9992) <= not(inputs(231));
    layer0_outputs(9993) <= inputs(134);
    layer0_outputs(9994) <= (inputs(135)) xor (inputs(43));
    layer0_outputs(9995) <= (inputs(163)) xor (inputs(198));
    layer0_outputs(9996) <= '1';
    layer0_outputs(9997) <= (inputs(240)) and not (inputs(35));
    layer0_outputs(9998) <= (inputs(155)) and not (inputs(230));
    layer0_outputs(9999) <= (inputs(36)) xor (inputs(146));
    layer0_outputs(10000) <= inputs(195);
    layer0_outputs(10001) <= (inputs(184)) and not (inputs(178));
    layer0_outputs(10002) <= inputs(90);
    layer0_outputs(10003) <= not(inputs(104));
    layer0_outputs(10004) <= inputs(100);
    layer0_outputs(10005) <= inputs(229);
    layer0_outputs(10006) <= (inputs(15)) and not (inputs(130));
    layer0_outputs(10007) <= not((inputs(139)) or (inputs(215)));
    layer0_outputs(10008) <= not(inputs(234));
    layer0_outputs(10009) <= (inputs(252)) and (inputs(208));
    layer0_outputs(10010) <= (inputs(229)) and not (inputs(66));
    layer0_outputs(10011) <= not((inputs(48)) or (inputs(182)));
    layer0_outputs(10012) <= '1';
    layer0_outputs(10013) <= not(inputs(0)) or (inputs(99));
    layer0_outputs(10014) <= (inputs(130)) xor (inputs(109));
    layer0_outputs(10015) <= not((inputs(13)) xor (inputs(172)));
    layer0_outputs(10016) <= (inputs(223)) and not (inputs(45));
    layer0_outputs(10017) <= not((inputs(243)) or (inputs(108)));
    layer0_outputs(10018) <= not((inputs(1)) or (inputs(116)));
    layer0_outputs(10019) <= not((inputs(179)) xor (inputs(31)));
    layer0_outputs(10020) <= (inputs(135)) and not (inputs(31));
    layer0_outputs(10021) <= not(inputs(41)) or (inputs(32));
    layer0_outputs(10022) <= (inputs(17)) or (inputs(71));
    layer0_outputs(10023) <= (inputs(93)) xor (inputs(13));
    layer0_outputs(10024) <= (inputs(175)) xor (inputs(161));
    layer0_outputs(10025) <= not(inputs(86)) or (inputs(146));
    layer0_outputs(10026) <= (inputs(21)) xor (inputs(150));
    layer0_outputs(10027) <= not(inputs(120));
    layer0_outputs(10028) <= (inputs(91)) or (inputs(94));
    layer0_outputs(10029) <= inputs(213);
    layer0_outputs(10030) <= not((inputs(178)) and (inputs(142)));
    layer0_outputs(10031) <= (inputs(87)) and not (inputs(37));
    layer0_outputs(10032) <= not(inputs(119));
    layer0_outputs(10033) <= (inputs(189)) or (inputs(140));
    layer0_outputs(10034) <= not(inputs(107));
    layer0_outputs(10035) <= not((inputs(44)) xor (inputs(218)));
    layer0_outputs(10036) <= (inputs(234)) or (inputs(91));
    layer0_outputs(10037) <= not(inputs(153));
    layer0_outputs(10038) <= (inputs(86)) xor (inputs(229));
    layer0_outputs(10039) <= (inputs(137)) and not (inputs(81));
    layer0_outputs(10040) <= (inputs(59)) and not (inputs(208));
    layer0_outputs(10041) <= not((inputs(117)) xor (inputs(209)));
    layer0_outputs(10042) <= not(inputs(140)) or (inputs(229));
    layer0_outputs(10043) <= inputs(86);
    layer0_outputs(10044) <= (inputs(27)) and not (inputs(160));
    layer0_outputs(10045) <= not((inputs(121)) or (inputs(190)));
    layer0_outputs(10046) <= (inputs(62)) and (inputs(159));
    layer0_outputs(10047) <= (inputs(214)) or (inputs(93));
    layer0_outputs(10048) <= not(inputs(193));
    layer0_outputs(10049) <= (inputs(235)) and not (inputs(59));
    layer0_outputs(10050) <= inputs(202);
    layer0_outputs(10051) <= (inputs(107)) and not (inputs(196));
    layer0_outputs(10052) <= not(inputs(88));
    layer0_outputs(10053) <= (inputs(131)) xor (inputs(166));
    layer0_outputs(10054) <= not(inputs(161));
    layer0_outputs(10055) <= not(inputs(181)) or (inputs(220));
    layer0_outputs(10056) <= (inputs(218)) or (inputs(104));
    layer0_outputs(10057) <= not((inputs(159)) or (inputs(83)));
    layer0_outputs(10058) <= '0';
    layer0_outputs(10059) <= not(inputs(36)) or (inputs(113));
    layer0_outputs(10060) <= (inputs(186)) or (inputs(134));
    layer0_outputs(10061) <= not(inputs(218)) or (inputs(49));
    layer0_outputs(10062) <= not(inputs(168));
    layer0_outputs(10063) <= inputs(106);
    layer0_outputs(10064) <= inputs(154);
    layer0_outputs(10065) <= not((inputs(116)) xor (inputs(212)));
    layer0_outputs(10066) <= not((inputs(209)) or (inputs(204)));
    layer0_outputs(10067) <= not(inputs(77));
    layer0_outputs(10068) <= not(inputs(154)) or (inputs(25));
    layer0_outputs(10069) <= not(inputs(228));
    layer0_outputs(10070) <= (inputs(217)) and (inputs(112));
    layer0_outputs(10071) <= (inputs(129)) xor (inputs(110));
    layer0_outputs(10072) <= not((inputs(54)) or (inputs(150)));
    layer0_outputs(10073) <= not(inputs(180)) or (inputs(34));
    layer0_outputs(10074) <= not((inputs(109)) or (inputs(218)));
    layer0_outputs(10075) <= not(inputs(119));
    layer0_outputs(10076) <= (inputs(61)) or (inputs(226));
    layer0_outputs(10077) <= (inputs(115)) or (inputs(100));
    layer0_outputs(10078) <= (inputs(117)) or (inputs(150));
    layer0_outputs(10079) <= (inputs(126)) and not (inputs(130));
    layer0_outputs(10080) <= (inputs(72)) or (inputs(96));
    layer0_outputs(10081) <= (inputs(155)) and not (inputs(91));
    layer0_outputs(10082) <= '1';
    layer0_outputs(10083) <= not((inputs(123)) or (inputs(155)));
    layer0_outputs(10084) <= (inputs(61)) and not (inputs(5));
    layer0_outputs(10085) <= '0';
    layer0_outputs(10086) <= not((inputs(15)) and (inputs(43)));
    layer0_outputs(10087) <= not(inputs(55));
    layer0_outputs(10088) <= (inputs(241)) and (inputs(194));
    layer0_outputs(10089) <= inputs(216);
    layer0_outputs(10090) <= (inputs(215)) and not (inputs(243));
    layer0_outputs(10091) <= not(inputs(228)) or (inputs(32));
    layer0_outputs(10092) <= (inputs(14)) xor (inputs(224));
    layer0_outputs(10093) <= (inputs(140)) and not (inputs(236));
    layer0_outputs(10094) <= not(inputs(60)) or (inputs(194));
    layer0_outputs(10095) <= '0';
    layer0_outputs(10096) <= not((inputs(12)) or (inputs(212)));
    layer0_outputs(10097) <= not(inputs(75)) or (inputs(7));
    layer0_outputs(10098) <= not((inputs(251)) or (inputs(234)));
    layer0_outputs(10099) <= not((inputs(103)) xor (inputs(157)));
    layer0_outputs(10100) <= (inputs(187)) or (inputs(172));
    layer0_outputs(10101) <= not(inputs(95));
    layer0_outputs(10102) <= inputs(246);
    layer0_outputs(10103) <= (inputs(232)) or (inputs(55));
    layer0_outputs(10104) <= (inputs(30)) and not (inputs(108));
    layer0_outputs(10105) <= (inputs(101)) or (inputs(148));
    layer0_outputs(10106) <= (inputs(171)) or (inputs(158));
    layer0_outputs(10107) <= (inputs(46)) or (inputs(248));
    layer0_outputs(10108) <= not(inputs(207)) or (inputs(127));
    layer0_outputs(10109) <= (inputs(105)) xor (inputs(32));
    layer0_outputs(10110) <= (inputs(151)) and not (inputs(166));
    layer0_outputs(10111) <= (inputs(214)) or (inputs(146));
    layer0_outputs(10112) <= '0';
    layer0_outputs(10113) <= (inputs(205)) and not (inputs(247));
    layer0_outputs(10114) <= not(inputs(119));
    layer0_outputs(10115) <= not(inputs(109)) or (inputs(1));
    layer0_outputs(10116) <= not((inputs(156)) or (inputs(143)));
    layer0_outputs(10117) <= not(inputs(84)) or (inputs(207));
    layer0_outputs(10118) <= not(inputs(80));
    layer0_outputs(10119) <= not(inputs(135)) or (inputs(5));
    layer0_outputs(10120) <= not(inputs(7));
    layer0_outputs(10121) <= '0';
    layer0_outputs(10122) <= (inputs(189)) and not (inputs(7));
    layer0_outputs(10123) <= inputs(188);
    layer0_outputs(10124) <= not(inputs(74));
    layer0_outputs(10125) <= (inputs(91)) or (inputs(67));
    layer0_outputs(10126) <= inputs(196);
    layer0_outputs(10127) <= (inputs(27)) or (inputs(32));
    layer0_outputs(10128) <= (inputs(141)) or (inputs(181));
    layer0_outputs(10129) <= (inputs(122)) or (inputs(194));
    layer0_outputs(10130) <= '1';
    layer0_outputs(10131) <= inputs(200);
    layer0_outputs(10132) <= not((inputs(195)) or (inputs(252)));
    layer0_outputs(10133) <= not(inputs(255));
    layer0_outputs(10134) <= inputs(168);
    layer0_outputs(10135) <= (inputs(217)) or (inputs(68));
    layer0_outputs(10136) <= not((inputs(167)) or (inputs(173)));
    layer0_outputs(10137) <= inputs(153);
    layer0_outputs(10138) <= not(inputs(229));
    layer0_outputs(10139) <= (inputs(208)) xor (inputs(215));
    layer0_outputs(10140) <= (inputs(122)) or (inputs(61));
    layer0_outputs(10141) <= not((inputs(252)) or (inputs(229)));
    layer0_outputs(10142) <= not(inputs(63));
    layer0_outputs(10143) <= inputs(147);
    layer0_outputs(10144) <= (inputs(101)) and not (inputs(30));
    layer0_outputs(10145) <= (inputs(99)) xor (inputs(13));
    layer0_outputs(10146) <= '0';
    layer0_outputs(10147) <= not(inputs(31)) or (inputs(131));
    layer0_outputs(10148) <= (inputs(113)) and (inputs(136));
    layer0_outputs(10149) <= not(inputs(118));
    layer0_outputs(10150) <= not(inputs(96)) or (inputs(30));
    layer0_outputs(10151) <= not((inputs(100)) or (inputs(159)));
    layer0_outputs(10152) <= inputs(48);
    layer0_outputs(10153) <= not((inputs(212)) xor (inputs(233)));
    layer0_outputs(10154) <= not((inputs(12)) xor (inputs(69)));
    layer0_outputs(10155) <= not((inputs(199)) xor (inputs(230)));
    layer0_outputs(10156) <= not((inputs(205)) xor (inputs(199)));
    layer0_outputs(10157) <= not((inputs(82)) or (inputs(167)));
    layer0_outputs(10158) <= (inputs(212)) or (inputs(230));
    layer0_outputs(10159) <= (inputs(228)) or (inputs(210));
    layer0_outputs(10160) <= not((inputs(137)) or (inputs(27)));
    layer0_outputs(10161) <= not((inputs(185)) and (inputs(198)));
    layer0_outputs(10162) <= (inputs(100)) or (inputs(205));
    layer0_outputs(10163) <= not((inputs(37)) xor (inputs(18)));
    layer0_outputs(10164) <= (inputs(49)) xor (inputs(189));
    layer0_outputs(10165) <= not(inputs(181));
    layer0_outputs(10166) <= not((inputs(181)) xor (inputs(36)));
    layer0_outputs(10167) <= (inputs(213)) or (inputs(60));
    layer0_outputs(10168) <= not(inputs(230));
    layer0_outputs(10169) <= not(inputs(217));
    layer0_outputs(10170) <= '1';
    layer0_outputs(10171) <= not(inputs(153)) or (inputs(115));
    layer0_outputs(10172) <= (inputs(0)) or (inputs(150));
    layer0_outputs(10173) <= (inputs(95)) or (inputs(54));
    layer0_outputs(10174) <= not((inputs(228)) and (inputs(189)));
    layer0_outputs(10175) <= inputs(199);
    layer0_outputs(10176) <= not((inputs(160)) or (inputs(252)));
    layer0_outputs(10177) <= (inputs(185)) and not (inputs(189));
    layer0_outputs(10178) <= inputs(61);
    layer0_outputs(10179) <= not((inputs(87)) xor (inputs(147)));
    layer0_outputs(10180) <= '0';
    layer0_outputs(10181) <= inputs(132);
    layer0_outputs(10182) <= not((inputs(224)) or (inputs(252)));
    layer0_outputs(10183) <= not(inputs(181));
    layer0_outputs(10184) <= inputs(151);
    layer0_outputs(10185) <= (inputs(52)) and not (inputs(192));
    layer0_outputs(10186) <= not(inputs(173)) or (inputs(218));
    layer0_outputs(10187) <= not((inputs(184)) xor (inputs(55)));
    layer0_outputs(10188) <= (inputs(226)) xor (inputs(146));
    layer0_outputs(10189) <= (inputs(102)) and not (inputs(97));
    layer0_outputs(10190) <= (inputs(4)) or (inputs(198));
    layer0_outputs(10191) <= inputs(40);
    layer0_outputs(10192) <= inputs(148);
    layer0_outputs(10193) <= (inputs(33)) and not (inputs(1));
    layer0_outputs(10194) <= inputs(7);
    layer0_outputs(10195) <= not((inputs(207)) or (inputs(33)));
    layer0_outputs(10196) <= inputs(249);
    layer0_outputs(10197) <= not((inputs(10)) and (inputs(64)));
    layer0_outputs(10198) <= not(inputs(173));
    layer0_outputs(10199) <= (inputs(254)) and (inputs(43));
    layer0_outputs(10200) <= inputs(42);
    layer0_outputs(10201) <= (inputs(116)) and not (inputs(14));
    layer0_outputs(10202) <= (inputs(205)) xor (inputs(174));
    layer0_outputs(10203) <= inputs(94);
    layer0_outputs(10204) <= (inputs(171)) or (inputs(73));
    layer0_outputs(10205) <= not((inputs(192)) xor (inputs(138)));
    layer0_outputs(10206) <= (inputs(88)) and not (inputs(161));
    layer0_outputs(10207) <= not(inputs(133));
    layer0_outputs(10208) <= not((inputs(48)) and (inputs(246)));
    layer0_outputs(10209) <= inputs(202);
    layer0_outputs(10210) <= (inputs(129)) and not (inputs(251));
    layer0_outputs(10211) <= not((inputs(57)) xor (inputs(10)));
    layer0_outputs(10212) <= (inputs(164)) and (inputs(23));
    layer0_outputs(10213) <= (inputs(36)) or (inputs(104));
    layer0_outputs(10214) <= (inputs(70)) and not (inputs(20));
    layer0_outputs(10215) <= not(inputs(27)) or (inputs(237));
    layer0_outputs(10216) <= '1';
    layer0_outputs(10217) <= not(inputs(226));
    layer0_outputs(10218) <= (inputs(200)) or (inputs(238));
    layer0_outputs(10219) <= inputs(170);
    layer0_outputs(10220) <= (inputs(197)) and not (inputs(93));
    layer0_outputs(10221) <= not(inputs(75));
    layer0_outputs(10222) <= not(inputs(109));
    layer0_outputs(10223) <= not(inputs(139)) or (inputs(164));
    layer0_outputs(10224) <= not((inputs(112)) xor (inputs(199)));
    layer0_outputs(10225) <= not(inputs(80));
    layer0_outputs(10226) <= not((inputs(117)) xor (inputs(18)));
    layer0_outputs(10227) <= (inputs(37)) xor (inputs(231));
    layer0_outputs(10228) <= inputs(37);
    layer0_outputs(10229) <= not(inputs(169)) or (inputs(219));
    layer0_outputs(10230) <= not(inputs(92)) or (inputs(81));
    layer0_outputs(10231) <= not((inputs(254)) or (inputs(158)));
    layer0_outputs(10232) <= (inputs(131)) or (inputs(223));
    layer0_outputs(10233) <= (inputs(196)) or (inputs(190));
    layer0_outputs(10234) <= (inputs(147)) or (inputs(38));
    layer0_outputs(10235) <= not((inputs(0)) or (inputs(140)));
    layer0_outputs(10236) <= not((inputs(86)) or (inputs(181)));
    layer0_outputs(10237) <= not((inputs(247)) xor (inputs(102)));
    layer0_outputs(10238) <= not((inputs(200)) xor (inputs(216)));
    layer0_outputs(10239) <= '0';
    outputs(0) <= (layer0_outputs(5076)) and not (layer0_outputs(5838));
    outputs(1) <= (layer0_outputs(7252)) and not (layer0_outputs(8310));
    outputs(2) <= (layer0_outputs(6041)) or (layer0_outputs(2449));
    outputs(3) <= not(layer0_outputs(1720));
    outputs(4) <= not(layer0_outputs(4807));
    outputs(5) <= not(layer0_outputs(1296));
    outputs(6) <= not((layer0_outputs(3142)) xor (layer0_outputs(6826)));
    outputs(7) <= (layer0_outputs(8140)) xor (layer0_outputs(2453));
    outputs(8) <= layer0_outputs(1904);
    outputs(9) <= not(layer0_outputs(3979));
    outputs(10) <= not(layer0_outputs(5415));
    outputs(11) <= (layer0_outputs(991)) and not (layer0_outputs(3098));
    outputs(12) <= not(layer0_outputs(6282));
    outputs(13) <= not((layer0_outputs(3535)) xor (layer0_outputs(6402)));
    outputs(14) <= not((layer0_outputs(1783)) xor (layer0_outputs(9080)));
    outputs(15) <= layer0_outputs(1353);
    outputs(16) <= not(layer0_outputs(2344));
    outputs(17) <= not(layer0_outputs(2362));
    outputs(18) <= not((layer0_outputs(9835)) and (layer0_outputs(366)));
    outputs(19) <= not(layer0_outputs(5713)) or (layer0_outputs(1630));
    outputs(20) <= not(layer0_outputs(1165));
    outputs(21) <= not((layer0_outputs(5931)) or (layer0_outputs(3101)));
    outputs(22) <= (layer0_outputs(2216)) and not (layer0_outputs(4677));
    outputs(23) <= not(layer0_outputs(636));
    outputs(24) <= '1';
    outputs(25) <= not(layer0_outputs(514));
    outputs(26) <= not((layer0_outputs(7825)) xor (layer0_outputs(2112)));
    outputs(27) <= layer0_outputs(1446);
    outputs(28) <= (layer0_outputs(3279)) xor (layer0_outputs(2172));
    outputs(29) <= layer0_outputs(2240);
    outputs(30) <= layer0_outputs(8527);
    outputs(31) <= not((layer0_outputs(3762)) xor (layer0_outputs(5326)));
    outputs(32) <= (layer0_outputs(9731)) and not (layer0_outputs(4347));
    outputs(33) <= (layer0_outputs(3425)) and (layer0_outputs(9254));
    outputs(34) <= (layer0_outputs(10233)) and not (layer0_outputs(9376));
    outputs(35) <= not((layer0_outputs(8448)) and (layer0_outputs(7847)));
    outputs(36) <= not(layer0_outputs(5317));
    outputs(37) <= layer0_outputs(595);
    outputs(38) <= not(layer0_outputs(8853));
    outputs(39) <= not(layer0_outputs(4391));
    outputs(40) <= not(layer0_outputs(4037));
    outputs(41) <= not((layer0_outputs(2710)) and (layer0_outputs(6605)));
    outputs(42) <= not(layer0_outputs(6114));
    outputs(43) <= layer0_outputs(6948);
    outputs(44) <= not(layer0_outputs(8870)) or (layer0_outputs(9388));
    outputs(45) <= layer0_outputs(1821);
    outputs(46) <= not(layer0_outputs(6470));
    outputs(47) <= (layer0_outputs(5233)) and (layer0_outputs(9055));
    outputs(48) <= not(layer0_outputs(9599));
    outputs(49) <= (layer0_outputs(5208)) or (layer0_outputs(7424));
    outputs(50) <= not(layer0_outputs(452));
    outputs(51) <= not(layer0_outputs(7412));
    outputs(52) <= layer0_outputs(1301);
    outputs(53) <= not(layer0_outputs(1320));
    outputs(54) <= not(layer0_outputs(4949)) or (layer0_outputs(1293));
    outputs(55) <= not(layer0_outputs(6878));
    outputs(56) <= not((layer0_outputs(5739)) and (layer0_outputs(8899)));
    outputs(57) <= not(layer0_outputs(5257));
    outputs(58) <= (layer0_outputs(8781)) xor (layer0_outputs(8994));
    outputs(59) <= not((layer0_outputs(9463)) xor (layer0_outputs(3182)));
    outputs(60) <= (layer0_outputs(7377)) or (layer0_outputs(7963));
    outputs(61) <= not(layer0_outputs(3076)) or (layer0_outputs(4613));
    outputs(62) <= (layer0_outputs(9500)) and not (layer0_outputs(5085));
    outputs(63) <= layer0_outputs(7066);
    outputs(64) <= layer0_outputs(7370);
    outputs(65) <= layer0_outputs(6525);
    outputs(66) <= layer0_outputs(7216);
    outputs(67) <= (layer0_outputs(7800)) and not (layer0_outputs(5374));
    outputs(68) <= not(layer0_outputs(6820));
    outputs(69) <= not(layer0_outputs(9075));
    outputs(70) <= not((layer0_outputs(6092)) xor (layer0_outputs(3556)));
    outputs(71) <= not(layer0_outputs(9318));
    outputs(72) <= not((layer0_outputs(7398)) or (layer0_outputs(2519)));
    outputs(73) <= (layer0_outputs(9653)) or (layer0_outputs(7342));
    outputs(74) <= not((layer0_outputs(789)) and (layer0_outputs(3053)));
    outputs(75) <= (layer0_outputs(5776)) and not (layer0_outputs(2496));
    outputs(76) <= not(layer0_outputs(9536));
    outputs(77) <= (layer0_outputs(7959)) and (layer0_outputs(1388));
    outputs(78) <= (layer0_outputs(1441)) and not (layer0_outputs(3600));
    outputs(79) <= (layer0_outputs(2192)) and (layer0_outputs(88));
    outputs(80) <= not(layer0_outputs(4242));
    outputs(81) <= layer0_outputs(2831);
    outputs(82) <= layer0_outputs(6793);
    outputs(83) <= not(layer0_outputs(10110));
    outputs(84) <= not(layer0_outputs(1629));
    outputs(85) <= layer0_outputs(3753);
    outputs(86) <= (layer0_outputs(9519)) xor (layer0_outputs(8908));
    outputs(87) <= (layer0_outputs(3055)) or (layer0_outputs(6222));
    outputs(88) <= (layer0_outputs(208)) or (layer0_outputs(2215));
    outputs(89) <= layer0_outputs(6551);
    outputs(90) <= not(layer0_outputs(9616));
    outputs(91) <= not(layer0_outputs(6120)) or (layer0_outputs(1234));
    outputs(92) <= not((layer0_outputs(9174)) xor (layer0_outputs(1767)));
    outputs(93) <= (layer0_outputs(4910)) or (layer0_outputs(8187));
    outputs(94) <= not(layer0_outputs(3089));
    outputs(95) <= layer0_outputs(7244);
    outputs(96) <= not(layer0_outputs(812)) or (layer0_outputs(8182));
    outputs(97) <= not((layer0_outputs(9383)) or (layer0_outputs(9035)));
    outputs(98) <= not((layer0_outputs(807)) xor (layer0_outputs(3850)));
    outputs(99) <= not(layer0_outputs(3163)) or (layer0_outputs(5505));
    outputs(100) <= not((layer0_outputs(7556)) xor (layer0_outputs(5261)));
    outputs(101) <= not((layer0_outputs(4421)) or (layer0_outputs(2549)));
    outputs(102) <= (layer0_outputs(4445)) or (layer0_outputs(1146));
    outputs(103) <= not((layer0_outputs(1305)) xor (layer0_outputs(8059)));
    outputs(104) <= layer0_outputs(6134);
    outputs(105) <= (layer0_outputs(7967)) and not (layer0_outputs(4405));
    outputs(106) <= (layer0_outputs(9272)) or (layer0_outputs(5292));
    outputs(107) <= (layer0_outputs(2507)) xor (layer0_outputs(9400));
    outputs(108) <= not((layer0_outputs(7901)) and (layer0_outputs(2085)));
    outputs(109) <= not(layer0_outputs(3183));
    outputs(110) <= (layer0_outputs(6686)) or (layer0_outputs(2563));
    outputs(111) <= not(layer0_outputs(3714));
    outputs(112) <= not(layer0_outputs(1933));
    outputs(113) <= layer0_outputs(6773);
    outputs(114) <= not((layer0_outputs(348)) xor (layer0_outputs(109)));
    outputs(115) <= layer0_outputs(2969);
    outputs(116) <= not(layer0_outputs(9762));
    outputs(117) <= not(layer0_outputs(6041));
    outputs(118) <= not(layer0_outputs(1912));
    outputs(119) <= not(layer0_outputs(7017));
    outputs(120) <= (layer0_outputs(9635)) xor (layer0_outputs(103));
    outputs(121) <= layer0_outputs(8521);
    outputs(122) <= layer0_outputs(682);
    outputs(123) <= not(layer0_outputs(9581));
    outputs(124) <= layer0_outputs(7251);
    outputs(125) <= not(layer0_outputs(9870));
    outputs(126) <= not(layer0_outputs(6311));
    outputs(127) <= layer0_outputs(8359);
    outputs(128) <= not((layer0_outputs(1525)) xor (layer0_outputs(5295)));
    outputs(129) <= not(layer0_outputs(7171));
    outputs(130) <= (layer0_outputs(4914)) and not (layer0_outputs(8129));
    outputs(131) <= not((layer0_outputs(4368)) or (layer0_outputs(2161)));
    outputs(132) <= not(layer0_outputs(9414));
    outputs(133) <= (layer0_outputs(2607)) and not (layer0_outputs(8713));
    outputs(134) <= not(layer0_outputs(9332)) or (layer0_outputs(4889));
    outputs(135) <= not((layer0_outputs(6512)) xor (layer0_outputs(9435)));
    outputs(136) <= (layer0_outputs(9358)) and not (layer0_outputs(5793));
    outputs(137) <= layer0_outputs(8254);
    outputs(138) <= not((layer0_outputs(4493)) or (layer0_outputs(10113)));
    outputs(139) <= not(layer0_outputs(7495));
    outputs(140) <= not((layer0_outputs(1879)) and (layer0_outputs(879)));
    outputs(141) <= not(layer0_outputs(9678));
    outputs(142) <= not((layer0_outputs(4577)) or (layer0_outputs(8066)));
    outputs(143) <= not(layer0_outputs(7673));
    outputs(144) <= not((layer0_outputs(717)) or (layer0_outputs(5954)));
    outputs(145) <= layer0_outputs(7257);
    outputs(146) <= not((layer0_outputs(5869)) xor (layer0_outputs(2817)));
    outputs(147) <= not((layer0_outputs(2596)) xor (layer0_outputs(10068)));
    outputs(148) <= layer0_outputs(539);
    outputs(149) <= layer0_outputs(6572);
    outputs(150) <= not(layer0_outputs(96)) or (layer0_outputs(2951));
    outputs(151) <= not(layer0_outputs(8919));
    outputs(152) <= '0';
    outputs(153) <= layer0_outputs(5729);
    outputs(154) <= layer0_outputs(2798);
    outputs(155) <= not(layer0_outputs(2395));
    outputs(156) <= (layer0_outputs(6321)) and not (layer0_outputs(2929));
    outputs(157) <= (layer0_outputs(6940)) xor (layer0_outputs(7405));
    outputs(158) <= layer0_outputs(6932);
    outputs(159) <= layer0_outputs(3403);
    outputs(160) <= (layer0_outputs(9590)) xor (layer0_outputs(1185));
    outputs(161) <= not((layer0_outputs(4625)) xor (layer0_outputs(6596)));
    outputs(162) <= (layer0_outputs(3470)) or (layer0_outputs(249));
    outputs(163) <= not(layer0_outputs(8975));
    outputs(164) <= not((layer0_outputs(5588)) xor (layer0_outputs(9460)));
    outputs(165) <= not(layer0_outputs(1291)) or (layer0_outputs(3606));
    outputs(166) <= not((layer0_outputs(9826)) xor (layer0_outputs(5911)));
    outputs(167) <= not((layer0_outputs(9520)) xor (layer0_outputs(2368)));
    outputs(168) <= not((layer0_outputs(5238)) and (layer0_outputs(3414)));
    outputs(169) <= (layer0_outputs(1698)) and not (layer0_outputs(8415));
    outputs(170) <= layer0_outputs(3393);
    outputs(171) <= layer0_outputs(3841);
    outputs(172) <= layer0_outputs(4599);
    outputs(173) <= not(layer0_outputs(7603));
    outputs(174) <= (layer0_outputs(5130)) xor (layer0_outputs(2149));
    outputs(175) <= (layer0_outputs(2451)) xor (layer0_outputs(8435));
    outputs(176) <= not(layer0_outputs(2204));
    outputs(177) <= layer0_outputs(8104);
    outputs(178) <= not(layer0_outputs(9989));
    outputs(179) <= not(layer0_outputs(7099)) or (layer0_outputs(6357));
    outputs(180) <= (layer0_outputs(1761)) or (layer0_outputs(2000));
    outputs(181) <= not(layer0_outputs(7747));
    outputs(182) <= not((layer0_outputs(2054)) and (layer0_outputs(3343)));
    outputs(183) <= not(layer0_outputs(3367));
    outputs(184) <= layer0_outputs(6775);
    outputs(185) <= (layer0_outputs(6160)) and (layer0_outputs(8400));
    outputs(186) <= not((layer0_outputs(3019)) xor (layer0_outputs(7566)));
    outputs(187) <= not((layer0_outputs(8724)) and (layer0_outputs(2944)));
    outputs(188) <= layer0_outputs(4245);
    outputs(189) <= not(layer0_outputs(3579));
    outputs(190) <= layer0_outputs(7160);
    outputs(191) <= layer0_outputs(7703);
    outputs(192) <= layer0_outputs(469);
    outputs(193) <= not((layer0_outputs(3453)) xor (layer0_outputs(4966)));
    outputs(194) <= (layer0_outputs(1045)) and (layer0_outputs(1880));
    outputs(195) <= not(layer0_outputs(8325));
    outputs(196) <= layer0_outputs(729);
    outputs(197) <= layer0_outputs(8921);
    outputs(198) <= not((layer0_outputs(5352)) xor (layer0_outputs(46)));
    outputs(199) <= (layer0_outputs(3019)) or (layer0_outputs(7776));
    outputs(200) <= layer0_outputs(7508);
    outputs(201) <= not(layer0_outputs(1843));
    outputs(202) <= not(layer0_outputs(2516));
    outputs(203) <= layer0_outputs(9814);
    outputs(204) <= not(layer0_outputs(452));
    outputs(205) <= not((layer0_outputs(6758)) and (layer0_outputs(6245)));
    outputs(206) <= (layer0_outputs(7283)) and not (layer0_outputs(8151));
    outputs(207) <= not(layer0_outputs(4601));
    outputs(208) <= not((layer0_outputs(6121)) or (layer0_outputs(4838)));
    outputs(209) <= not((layer0_outputs(8056)) xor (layer0_outputs(4609)));
    outputs(210) <= not((layer0_outputs(8123)) xor (layer0_outputs(8845)));
    outputs(211) <= not(layer0_outputs(2359));
    outputs(212) <= (layer0_outputs(710)) xor (layer0_outputs(2713));
    outputs(213) <= (layer0_outputs(7263)) xor (layer0_outputs(9213));
    outputs(214) <= not(layer0_outputs(7262)) or (layer0_outputs(7788));
    outputs(215) <= (layer0_outputs(4802)) xor (layer0_outputs(8719));
    outputs(216) <= not(layer0_outputs(4963)) or (layer0_outputs(4483));
    outputs(217) <= '0';
    outputs(218) <= (layer0_outputs(6655)) and (layer0_outputs(8373));
    outputs(219) <= not((layer0_outputs(6774)) xor (layer0_outputs(892)));
    outputs(220) <= not(layer0_outputs(2115)) or (layer0_outputs(7600));
    outputs(221) <= layer0_outputs(1845);
    outputs(222) <= not(layer0_outputs(10185));
    outputs(223) <= not(layer0_outputs(8805));
    outputs(224) <= layer0_outputs(9184);
    outputs(225) <= layer0_outputs(1835);
    outputs(226) <= (layer0_outputs(7624)) xor (layer0_outputs(1489));
    outputs(227) <= not(layer0_outputs(9348));
    outputs(228) <= not(layer0_outputs(5067)) or (layer0_outputs(4470));
    outputs(229) <= layer0_outputs(1577);
    outputs(230) <= (layer0_outputs(2267)) xor (layer0_outputs(7764));
    outputs(231) <= layer0_outputs(8175);
    outputs(232) <= (layer0_outputs(794)) and not (layer0_outputs(9945));
    outputs(233) <= layer0_outputs(3275);
    outputs(234) <= layer0_outputs(2972);
    outputs(235) <= not(layer0_outputs(7848));
    outputs(236) <= not(layer0_outputs(1336));
    outputs(237) <= layer0_outputs(4478);
    outputs(238) <= (layer0_outputs(7104)) or (layer0_outputs(140));
    outputs(239) <= layer0_outputs(9223);
    outputs(240) <= (layer0_outputs(9779)) xor (layer0_outputs(2938));
    outputs(241) <= not(layer0_outputs(3684));
    outputs(242) <= layer0_outputs(5256);
    outputs(243) <= not((layer0_outputs(6598)) or (layer0_outputs(3221)));
    outputs(244) <= (layer0_outputs(10188)) or (layer0_outputs(4956));
    outputs(245) <= not(layer0_outputs(8865));
    outputs(246) <= not(layer0_outputs(1605));
    outputs(247) <= layer0_outputs(8440);
    outputs(248) <= not(layer0_outputs(9075));
    outputs(249) <= not(layer0_outputs(6757));
    outputs(250) <= layer0_outputs(2704);
    outputs(251) <= not(layer0_outputs(4995));
    outputs(252) <= not(layer0_outputs(7789)) or (layer0_outputs(9038));
    outputs(253) <= layer0_outputs(39);
    outputs(254) <= layer0_outputs(2382);
    outputs(255) <= layer0_outputs(1407);
    outputs(256) <= layer0_outputs(9823);
    outputs(257) <= layer0_outputs(8271);
    outputs(258) <= not(layer0_outputs(10129)) or (layer0_outputs(9477));
    outputs(259) <= not((layer0_outputs(1135)) xor (layer0_outputs(7818)));
    outputs(260) <= (layer0_outputs(3996)) and not (layer0_outputs(5872));
    outputs(261) <= (layer0_outputs(6042)) xor (layer0_outputs(5408));
    outputs(262) <= (layer0_outputs(8565)) xor (layer0_outputs(8640));
    outputs(263) <= not(layer0_outputs(6439));
    outputs(264) <= not(layer0_outputs(9970));
    outputs(265) <= (layer0_outputs(10005)) xor (layer0_outputs(8032));
    outputs(266) <= layer0_outputs(9969);
    outputs(267) <= layer0_outputs(6583);
    outputs(268) <= layer0_outputs(3487);
    outputs(269) <= not(layer0_outputs(2942));
    outputs(270) <= not((layer0_outputs(2041)) xor (layer0_outputs(9771)));
    outputs(271) <= not(layer0_outputs(5837));
    outputs(272) <= (layer0_outputs(1350)) xor (layer0_outputs(462));
    outputs(273) <= layer0_outputs(3608);
    outputs(274) <= not(layer0_outputs(4851));
    outputs(275) <= (layer0_outputs(6909)) xor (layer0_outputs(9088));
    outputs(276) <= layer0_outputs(9457);
    outputs(277) <= (layer0_outputs(1890)) xor (layer0_outputs(3997));
    outputs(278) <= layer0_outputs(8946);
    outputs(279) <= not((layer0_outputs(8748)) xor (layer0_outputs(10117)));
    outputs(280) <= not((layer0_outputs(4803)) xor (layer0_outputs(6475)));
    outputs(281) <= not((layer0_outputs(2680)) xor (layer0_outputs(6726)));
    outputs(282) <= (layer0_outputs(7018)) and (layer0_outputs(957));
    outputs(283) <= '1';
    outputs(284) <= (layer0_outputs(5652)) and (layer0_outputs(6423));
    outputs(285) <= layer0_outputs(9497);
    outputs(286) <= (layer0_outputs(5581)) xor (layer0_outputs(3329));
    outputs(287) <= layer0_outputs(2270);
    outputs(288) <= layer0_outputs(6150);
    outputs(289) <= not(layer0_outputs(6382));
    outputs(290) <= (layer0_outputs(1487)) and not (layer0_outputs(6544));
    outputs(291) <= (layer0_outputs(3064)) and not (layer0_outputs(755));
    outputs(292) <= not((layer0_outputs(9550)) xor (layer0_outputs(8349)));
    outputs(293) <= (layer0_outputs(3137)) and not (layer0_outputs(7044));
    outputs(294) <= layer0_outputs(8270);
    outputs(295) <= (layer0_outputs(8188)) and (layer0_outputs(9263));
    outputs(296) <= layer0_outputs(195);
    outputs(297) <= layer0_outputs(9747);
    outputs(298) <= '1';
    outputs(299) <= not(layer0_outputs(5501));
    outputs(300) <= (layer0_outputs(628)) or (layer0_outputs(8117));
    outputs(301) <= not((layer0_outputs(5029)) or (layer0_outputs(6841)));
    outputs(302) <= (layer0_outputs(9841)) and not (layer0_outputs(1707));
    outputs(303) <= layer0_outputs(726);
    outputs(304) <= layer0_outputs(1147);
    outputs(305) <= layer0_outputs(2053);
    outputs(306) <= not((layer0_outputs(6066)) xor (layer0_outputs(4920)));
    outputs(307) <= not((layer0_outputs(9980)) or (layer0_outputs(6028)));
    outputs(308) <= (layer0_outputs(3999)) and not (layer0_outputs(9173));
    outputs(309) <= not(layer0_outputs(5836));
    outputs(310) <= not(layer0_outputs(976));
    outputs(311) <= not((layer0_outputs(3306)) or (layer0_outputs(7867)));
    outputs(312) <= (layer0_outputs(9319)) xor (layer0_outputs(9857));
    outputs(313) <= not(layer0_outputs(2110)) or (layer0_outputs(9867));
    outputs(314) <= layer0_outputs(3178);
    outputs(315) <= not((layer0_outputs(5442)) xor (layer0_outputs(5013)));
    outputs(316) <= not(layer0_outputs(3799));
    outputs(317) <= not((layer0_outputs(8139)) or (layer0_outputs(8196)));
    outputs(318) <= not((layer0_outputs(3551)) xor (layer0_outputs(7669)));
    outputs(319) <= not(layer0_outputs(9750)) or (layer0_outputs(549));
    outputs(320) <= '1';
    outputs(321) <= layer0_outputs(1647);
    outputs(322) <= (layer0_outputs(7378)) xor (layer0_outputs(5695));
    outputs(323) <= (layer0_outputs(2645)) and not (layer0_outputs(8783));
    outputs(324) <= (layer0_outputs(6816)) or (layer0_outputs(9662));
    outputs(325) <= not(layer0_outputs(1854));
    outputs(326) <= (layer0_outputs(7287)) xor (layer0_outputs(492));
    outputs(327) <= (layer0_outputs(9065)) or (layer0_outputs(3051));
    outputs(328) <= not(layer0_outputs(190));
    outputs(329) <= not(layer0_outputs(5169));
    outputs(330) <= layer0_outputs(4585);
    outputs(331) <= not(layer0_outputs(7356));
    outputs(332) <= not((layer0_outputs(763)) xor (layer0_outputs(2515)));
    outputs(333) <= not(layer0_outputs(7489));
    outputs(334) <= not((layer0_outputs(661)) xor (layer0_outputs(9221)));
    outputs(335) <= not(layer0_outputs(8937));
    outputs(336) <= not(layer0_outputs(3422)) or (layer0_outputs(2861));
    outputs(337) <= not(layer0_outputs(8512)) or (layer0_outputs(8026));
    outputs(338) <= (layer0_outputs(4151)) xor (layer0_outputs(5696));
    outputs(339) <= not(layer0_outputs(5465));
    outputs(340) <= not(layer0_outputs(8141));
    outputs(341) <= layer0_outputs(8229);
    outputs(342) <= layer0_outputs(10157);
    outputs(343) <= (layer0_outputs(5693)) and not (layer0_outputs(3580));
    outputs(344) <= not((layer0_outputs(10035)) xor (layer0_outputs(5483)));
    outputs(345) <= not(layer0_outputs(2430));
    outputs(346) <= not(layer0_outputs(1952));
    outputs(347) <= (layer0_outputs(1858)) and not (layer0_outputs(3044));
    outputs(348) <= not(layer0_outputs(10224));
    outputs(349) <= (layer0_outputs(1545)) and not (layer0_outputs(4314));
    outputs(350) <= not((layer0_outputs(2953)) xor (layer0_outputs(236)));
    outputs(351) <= not(layer0_outputs(1703));
    outputs(352) <= not(layer0_outputs(3816));
    outputs(353) <= (layer0_outputs(9718)) and not (layer0_outputs(9144));
    outputs(354) <= not(layer0_outputs(6420)) or (layer0_outputs(5454));
    outputs(355) <= (layer0_outputs(18)) and not (layer0_outputs(4237));
    outputs(356) <= (layer0_outputs(1899)) and not (layer0_outputs(9543));
    outputs(357) <= layer0_outputs(8459);
    outputs(358) <= (layer0_outputs(644)) or (layer0_outputs(575));
    outputs(359) <= not(layer0_outputs(8549));
    outputs(360) <= not(layer0_outputs(8698));
    outputs(361) <= layer0_outputs(1187);
    outputs(362) <= not((layer0_outputs(5198)) xor (layer0_outputs(4864)));
    outputs(363) <= (layer0_outputs(2050)) and not (layer0_outputs(4569));
    outputs(364) <= not(layer0_outputs(5885));
    outputs(365) <= not(layer0_outputs(6629)) or (layer0_outputs(5694));
    outputs(366) <= not((layer0_outputs(8336)) and (layer0_outputs(3888)));
    outputs(367) <= not(layer0_outputs(8926)) or (layer0_outputs(9889));
    outputs(368) <= (layer0_outputs(3454)) and not (layer0_outputs(1751));
    outputs(369) <= (layer0_outputs(1345)) xor (layer0_outputs(1536));
    outputs(370) <= (layer0_outputs(4092)) and not (layer0_outputs(5414));
    outputs(371) <= not(layer0_outputs(6659)) or (layer0_outputs(7195));
    outputs(372) <= (layer0_outputs(5598)) and not (layer0_outputs(3295));
    outputs(373) <= not((layer0_outputs(7477)) xor (layer0_outputs(4249)));
    outputs(374) <= not(layer0_outputs(4039));
    outputs(375) <= not((layer0_outputs(6015)) and (layer0_outputs(2756)));
    outputs(376) <= layer0_outputs(5756);
    outputs(377) <= layer0_outputs(10040);
    outputs(378) <= not(layer0_outputs(7476));
    outputs(379) <= layer0_outputs(4655);
    outputs(380) <= not((layer0_outputs(2295)) xor (layer0_outputs(3122)));
    outputs(381) <= not(layer0_outputs(4513)) or (layer0_outputs(5210));
    outputs(382) <= not(layer0_outputs(4474));
    outputs(383) <= not((layer0_outputs(5707)) xor (layer0_outputs(9740)));
    outputs(384) <= not((layer0_outputs(835)) xor (layer0_outputs(3610)));
    outputs(385) <= layer0_outputs(10205);
    outputs(386) <= layer0_outputs(3954);
    outputs(387) <= not(layer0_outputs(824));
    outputs(388) <= not(layer0_outputs(5757));
    outputs(389) <= layer0_outputs(6585);
    outputs(390) <= not((layer0_outputs(1184)) or (layer0_outputs(3378)));
    outputs(391) <= not(layer0_outputs(602));
    outputs(392) <= layer0_outputs(8335);
    outputs(393) <= not(layer0_outputs(4705));
    outputs(394) <= not(layer0_outputs(5144));
    outputs(395) <= not((layer0_outputs(576)) xor (layer0_outputs(104)));
    outputs(396) <= (layer0_outputs(1001)) and (layer0_outputs(4136));
    outputs(397) <= (layer0_outputs(7208)) or (layer0_outputs(4646));
    outputs(398) <= layer0_outputs(5795);
    outputs(399) <= not((layer0_outputs(2011)) and (layer0_outputs(3624)));
    outputs(400) <= not((layer0_outputs(6904)) xor (layer0_outputs(8672)));
    outputs(401) <= layer0_outputs(1006);
    outputs(402) <= not(layer0_outputs(6980));
    outputs(403) <= layer0_outputs(8237);
    outputs(404) <= not((layer0_outputs(8890)) xor (layer0_outputs(1172)));
    outputs(405) <= not(layer0_outputs(7245));
    outputs(406) <= not(layer0_outputs(2094));
    outputs(407) <= not(layer0_outputs(9081));
    outputs(408) <= not((layer0_outputs(4030)) xor (layer0_outputs(918)));
    outputs(409) <= not(layer0_outputs(7476)) or (layer0_outputs(6674));
    outputs(410) <= not((layer0_outputs(8437)) xor (layer0_outputs(4062)));
    outputs(411) <= layer0_outputs(8161);
    outputs(412) <= layer0_outputs(8604);
    outputs(413) <= not(layer0_outputs(4664)) or (layer0_outputs(5059));
    outputs(414) <= (layer0_outputs(9846)) and (layer0_outputs(9207));
    outputs(415) <= not(layer0_outputs(9850));
    outputs(416) <= layer0_outputs(2309);
    outputs(417) <= not(layer0_outputs(5366));
    outputs(418) <= not((layer0_outputs(7276)) and (layer0_outputs(5879)));
    outputs(419) <= (layer0_outputs(1238)) or (layer0_outputs(7343));
    outputs(420) <= not((layer0_outputs(3255)) and (layer0_outputs(3198)));
    outputs(421) <= layer0_outputs(34);
    outputs(422) <= layer0_outputs(5432);
    outputs(423) <= not(layer0_outputs(7176)) or (layer0_outputs(2729));
    outputs(424) <= not((layer0_outputs(7336)) or (layer0_outputs(1068)));
    outputs(425) <= not((layer0_outputs(369)) and (layer0_outputs(8415)));
    outputs(426) <= not(layer0_outputs(6011));
    outputs(427) <= (layer0_outputs(2531)) and not (layer0_outputs(3708));
    outputs(428) <= (layer0_outputs(392)) and not (layer0_outputs(3980));
    outputs(429) <= not((layer0_outputs(1439)) xor (layer0_outputs(9549)));
    outputs(430) <= not(layer0_outputs(3654));
    outputs(431) <= (layer0_outputs(9744)) xor (layer0_outputs(9213));
    outputs(432) <= not(layer0_outputs(6964)) or (layer0_outputs(7466));
    outputs(433) <= not((layer0_outputs(3276)) xor (layer0_outputs(6531)));
    outputs(434) <= (layer0_outputs(7719)) and (layer0_outputs(4321));
    outputs(435) <= not(layer0_outputs(4673));
    outputs(436) <= layer0_outputs(5458);
    outputs(437) <= (layer0_outputs(3314)) and not (layer0_outputs(5059));
    outputs(438) <= not((layer0_outputs(2589)) xor (layer0_outputs(651)));
    outputs(439) <= not((layer0_outputs(9608)) xor (layer0_outputs(6007)));
    outputs(440) <= not(layer0_outputs(7777));
    outputs(441) <= not((layer0_outputs(1347)) or (layer0_outputs(8243)));
    outputs(442) <= not(layer0_outputs(6791)) or (layer0_outputs(6333));
    outputs(443) <= layer0_outputs(3408);
    outputs(444) <= (layer0_outputs(8102)) or (layer0_outputs(9333));
    outputs(445) <= layer0_outputs(6785);
    outputs(446) <= not(layer0_outputs(2492));
    outputs(447) <= not(layer0_outputs(8561));
    outputs(448) <= not((layer0_outputs(3948)) xor (layer0_outputs(3291)));
    outputs(449) <= not(layer0_outputs(9714));
    outputs(450) <= not(layer0_outputs(9957));
    outputs(451) <= layer0_outputs(6208);
    outputs(452) <= not(layer0_outputs(4443));
    outputs(453) <= not(layer0_outputs(980)) or (layer0_outputs(192));
    outputs(454) <= not(layer0_outputs(5060)) or (layer0_outputs(8644));
    outputs(455) <= layer0_outputs(9287);
    outputs(456) <= (layer0_outputs(9277)) xor (layer0_outputs(2520));
    outputs(457) <= not(layer0_outputs(4770));
    outputs(458) <= not((layer0_outputs(7124)) xor (layer0_outputs(8398)));
    outputs(459) <= not((layer0_outputs(5512)) and (layer0_outputs(8682)));
    outputs(460) <= layer0_outputs(8966);
    outputs(461) <= not((layer0_outputs(6920)) xor (layer0_outputs(1791)));
    outputs(462) <= not(layer0_outputs(1021));
    outputs(463) <= layer0_outputs(4679);
    outputs(464) <= (layer0_outputs(8990)) and (layer0_outputs(6050));
    outputs(465) <= not(layer0_outputs(6637));
    outputs(466) <= layer0_outputs(2807);
    outputs(467) <= layer0_outputs(6560);
    outputs(468) <= not(layer0_outputs(10020));
    outputs(469) <= not(layer0_outputs(3102));
    outputs(470) <= not((layer0_outputs(1660)) xor (layer0_outputs(8394)));
    outputs(471) <= not(layer0_outputs(1249)) or (layer0_outputs(3696));
    outputs(472) <= not(layer0_outputs(1037));
    outputs(473) <= not(layer0_outputs(998));
    outputs(474) <= (layer0_outputs(7209)) xor (layer0_outputs(1648));
    outputs(475) <= (layer0_outputs(7090)) or (layer0_outputs(5063));
    outputs(476) <= layer0_outputs(1537);
    outputs(477) <= (layer0_outputs(9436)) xor (layer0_outputs(8063));
    outputs(478) <= not(layer0_outputs(4417));
    outputs(479) <= not(layer0_outputs(1389));
    outputs(480) <= not(layer0_outputs(1249));
    outputs(481) <= not(layer0_outputs(10039));
    outputs(482) <= (layer0_outputs(1527)) and not (layer0_outputs(2336));
    outputs(483) <= not(layer0_outputs(6282));
    outputs(484) <= not(layer0_outputs(1776)) or (layer0_outputs(5005));
    outputs(485) <= layer0_outputs(7281);
    outputs(486) <= (layer0_outputs(9940)) and (layer0_outputs(10218));
    outputs(487) <= layer0_outputs(2016);
    outputs(488) <= not(layer0_outputs(8642));
    outputs(489) <= layer0_outputs(8688);
    outputs(490) <= not(layer0_outputs(6830));
    outputs(491) <= not(layer0_outputs(8322)) or (layer0_outputs(1196));
    outputs(492) <= layer0_outputs(8715);
    outputs(493) <= not((layer0_outputs(2098)) xor (layer0_outputs(5265)));
    outputs(494) <= not(layer0_outputs(4995)) or (layer0_outputs(3236));
    outputs(495) <= layer0_outputs(8120);
    outputs(496) <= not(layer0_outputs(7308));
    outputs(497) <= layer0_outputs(4363);
    outputs(498) <= layer0_outputs(5989);
    outputs(499) <= not((layer0_outputs(985)) xor (layer0_outputs(3999)));
    outputs(500) <= (layer0_outputs(763)) and not (layer0_outputs(3751));
    outputs(501) <= layer0_outputs(2887);
    outputs(502) <= not(layer0_outputs(258));
    outputs(503) <= not((layer0_outputs(7058)) xor (layer0_outputs(408)));
    outputs(504) <= not(layer0_outputs(1922));
    outputs(505) <= not(layer0_outputs(1137));
    outputs(506) <= (layer0_outputs(4333)) xor (layer0_outputs(4618));
    outputs(507) <= layer0_outputs(6746);
    outputs(508) <= layer0_outputs(6024);
    outputs(509) <= (layer0_outputs(4660)) and not (layer0_outputs(8303));
    outputs(510) <= layer0_outputs(7683);
    outputs(511) <= (layer0_outputs(1865)) and not (layer0_outputs(2830));
    outputs(512) <= layer0_outputs(5425);
    outputs(513) <= layer0_outputs(9544);
    outputs(514) <= not(layer0_outputs(4289));
    outputs(515) <= layer0_outputs(5054);
    outputs(516) <= (layer0_outputs(557)) or (layer0_outputs(5087));
    outputs(517) <= not(layer0_outputs(9900));
    outputs(518) <= not((layer0_outputs(6236)) xor (layer0_outputs(4409)));
    outputs(519) <= not((layer0_outputs(3630)) xor (layer0_outputs(3667)));
    outputs(520) <= not(layer0_outputs(4440));
    outputs(521) <= layer0_outputs(1363);
    outputs(522) <= layer0_outputs(6462);
    outputs(523) <= (layer0_outputs(1254)) xor (layer0_outputs(4125));
    outputs(524) <= not((layer0_outputs(2136)) xor (layer0_outputs(4595)));
    outputs(525) <= not((layer0_outputs(10188)) xor (layer0_outputs(9764)));
    outputs(526) <= not((layer0_outputs(5152)) xor (layer0_outputs(1282)));
    outputs(527) <= (layer0_outputs(4630)) xor (layer0_outputs(6173));
    outputs(528) <= not(layer0_outputs(5629)) or (layer0_outputs(7725));
    outputs(529) <= not(layer0_outputs(1392));
    outputs(530) <= layer0_outputs(1484);
    outputs(531) <= (layer0_outputs(8637)) xor (layer0_outputs(9017));
    outputs(532) <= layer0_outputs(162);
    outputs(533) <= (layer0_outputs(7555)) or (layer0_outputs(4652));
    outputs(534) <= (layer0_outputs(3930)) and not (layer0_outputs(9401));
    outputs(535) <= layer0_outputs(8878);
    outputs(536) <= layer0_outputs(4241);
    outputs(537) <= (layer0_outputs(6393)) or (layer0_outputs(943));
    outputs(538) <= not((layer0_outputs(8925)) xor (layer0_outputs(9197)));
    outputs(539) <= (layer0_outputs(8382)) xor (layer0_outputs(4064));
    outputs(540) <= layer0_outputs(5528);
    outputs(541) <= not(layer0_outputs(2657));
    outputs(542) <= (layer0_outputs(3485)) xor (layer0_outputs(135));
    outputs(543) <= layer0_outputs(2134);
    outputs(544) <= (layer0_outputs(7872)) xor (layer0_outputs(4882));
    outputs(545) <= layer0_outputs(1758);
    outputs(546) <= (layer0_outputs(3685)) xor (layer0_outputs(4874));
    outputs(547) <= (layer0_outputs(7263)) xor (layer0_outputs(8125));
    outputs(548) <= (layer0_outputs(8392)) xor (layer0_outputs(5221));
    outputs(549) <= (layer0_outputs(5584)) xor (layer0_outputs(4420));
    outputs(550) <= not(layer0_outputs(2385));
    outputs(551) <= not((layer0_outputs(6625)) xor (layer0_outputs(6758)));
    outputs(552) <= (layer0_outputs(6056)) or (layer0_outputs(6782));
    outputs(553) <= (layer0_outputs(7530)) and not (layer0_outputs(7612));
    outputs(554) <= (layer0_outputs(8231)) and not (layer0_outputs(9808));
    outputs(555) <= layer0_outputs(1151);
    outputs(556) <= layer0_outputs(1173);
    outputs(557) <= not(layer0_outputs(1124));
    outputs(558) <= layer0_outputs(453);
    outputs(559) <= (layer0_outputs(5691)) xor (layer0_outputs(3982));
    outputs(560) <= not(layer0_outputs(7481));
    outputs(561) <= '1';
    outputs(562) <= not(layer0_outputs(391)) or (layer0_outputs(703));
    outputs(563) <= layer0_outputs(5084);
    outputs(564) <= not(layer0_outputs(7917)) or (layer0_outputs(2211));
    outputs(565) <= not(layer0_outputs(10222));
    outputs(566) <= not(layer0_outputs(770));
    outputs(567) <= not(layer0_outputs(9554));
    outputs(568) <= layer0_outputs(1403);
    outputs(569) <= (layer0_outputs(9356)) xor (layer0_outputs(8014));
    outputs(570) <= not(layer0_outputs(6273)) or (layer0_outputs(1558));
    outputs(571) <= not(layer0_outputs(5126));
    outputs(572) <= not(layer0_outputs(2648));
    outputs(573) <= (layer0_outputs(8543)) or (layer0_outputs(943));
    outputs(574) <= not(layer0_outputs(3048));
    outputs(575) <= (layer0_outputs(7563)) xor (layer0_outputs(6724));
    outputs(576) <= not((layer0_outputs(9003)) xor (layer0_outputs(5082)));
    outputs(577) <= layer0_outputs(240);
    outputs(578) <= not((layer0_outputs(10059)) xor (layer0_outputs(6962)));
    outputs(579) <= not(layer0_outputs(1708));
    outputs(580) <= layer0_outputs(8293);
    outputs(581) <= not((layer0_outputs(6140)) or (layer0_outputs(1868)));
    outputs(582) <= (layer0_outputs(3768)) and not (layer0_outputs(6687));
    outputs(583) <= (layer0_outputs(6457)) and not (layer0_outputs(8423));
    outputs(584) <= (layer0_outputs(7373)) xor (layer0_outputs(1782));
    outputs(585) <= (layer0_outputs(8653)) xor (layer0_outputs(4303));
    outputs(586) <= layer0_outputs(3647);
    outputs(587) <= not(layer0_outputs(56));
    outputs(588) <= (layer0_outputs(772)) or (layer0_outputs(736));
    outputs(589) <= not(layer0_outputs(126));
    outputs(590) <= layer0_outputs(2293);
    outputs(591) <= not((layer0_outputs(6689)) and (layer0_outputs(5941)));
    outputs(592) <= layer0_outputs(182);
    outputs(593) <= layer0_outputs(5307);
    outputs(594) <= not(layer0_outputs(4940)) or (layer0_outputs(4121));
    outputs(595) <= not(layer0_outputs(6253));
    outputs(596) <= not((layer0_outputs(7701)) xor (layer0_outputs(3101)));
    outputs(597) <= (layer0_outputs(9679)) xor (layer0_outputs(4739));
    outputs(598) <= not(layer0_outputs(2553));
    outputs(599) <= not(layer0_outputs(10222));
    outputs(600) <= not((layer0_outputs(3780)) xor (layer0_outputs(6166)));
    outputs(601) <= not(layer0_outputs(8503)) or (layer0_outputs(2656));
    outputs(602) <= layer0_outputs(8545);
    outputs(603) <= not(layer0_outputs(1746));
    outputs(604) <= not((layer0_outputs(6089)) and (layer0_outputs(5977)));
    outputs(605) <= not(layer0_outputs(5168));
    outputs(606) <= (layer0_outputs(9765)) xor (layer0_outputs(6146));
    outputs(607) <= not(layer0_outputs(5527));
    outputs(608) <= layer0_outputs(1410);
    outputs(609) <= (layer0_outputs(9793)) and not (layer0_outputs(3160));
    outputs(610) <= not(layer0_outputs(7669)) or (layer0_outputs(519));
    outputs(611) <= not(layer0_outputs(7647));
    outputs(612) <= not((layer0_outputs(7552)) and (layer0_outputs(824)));
    outputs(613) <= not(layer0_outputs(3140));
    outputs(614) <= layer0_outputs(1749);
    outputs(615) <= not((layer0_outputs(8963)) xor (layer0_outputs(7008)));
    outputs(616) <= not(layer0_outputs(9411)) or (layer0_outputs(852));
    outputs(617) <= (layer0_outputs(9295)) and not (layer0_outputs(6009));
    outputs(618) <= not(layer0_outputs(4167)) or (layer0_outputs(8692));
    outputs(619) <= layer0_outputs(4790);
    outputs(620) <= not((layer0_outputs(904)) xor (layer0_outputs(7120)));
    outputs(621) <= not((layer0_outputs(7005)) and (layer0_outputs(3198)));
    outputs(622) <= (layer0_outputs(2186)) and not (layer0_outputs(1570));
    outputs(623) <= not(layer0_outputs(3111));
    outputs(624) <= not((layer0_outputs(564)) xor (layer0_outputs(9185)));
    outputs(625) <= not(layer0_outputs(2566));
    outputs(626) <= layer0_outputs(5883);
    outputs(627) <= layer0_outputs(1683);
    outputs(628) <= not(layer0_outputs(2937));
    outputs(629) <= layer0_outputs(569);
    outputs(630) <= (layer0_outputs(7519)) and (layer0_outputs(5128));
    outputs(631) <= (layer0_outputs(1514)) xor (layer0_outputs(874));
    outputs(632) <= layer0_outputs(6738);
    outputs(633) <= not(layer0_outputs(1935)) or (layer0_outputs(6070));
    outputs(634) <= not(layer0_outputs(6245)) or (layer0_outputs(4197));
    outputs(635) <= (layer0_outputs(237)) and (layer0_outputs(5539));
    outputs(636) <= not(layer0_outputs(4443));
    outputs(637) <= not(layer0_outputs(7941));
    outputs(638) <= layer0_outputs(3188);
    outputs(639) <= layer0_outputs(2480);
    outputs(640) <= not(layer0_outputs(9408));
    outputs(641) <= not((layer0_outputs(7697)) and (layer0_outputs(6200)));
    outputs(642) <= not((layer0_outputs(8703)) xor (layer0_outputs(4704)));
    outputs(643) <= not(layer0_outputs(2408));
    outputs(644) <= layer0_outputs(10143);
    outputs(645) <= not((layer0_outputs(9112)) or (layer0_outputs(7147)));
    outputs(646) <= layer0_outputs(7292);
    outputs(647) <= not(layer0_outputs(4188));
    outputs(648) <= not(layer0_outputs(7570));
    outputs(649) <= not(layer0_outputs(2266));
    outputs(650) <= (layer0_outputs(4870)) xor (layer0_outputs(6797));
    outputs(651) <= (layer0_outputs(5209)) xor (layer0_outputs(10063));
    outputs(652) <= not(layer0_outputs(10228));
    outputs(653) <= '1';
    outputs(654) <= (layer0_outputs(3691)) xor (layer0_outputs(1283));
    outputs(655) <= not(layer0_outputs(1318));
    outputs(656) <= not(layer0_outputs(2017));
    outputs(657) <= not(layer0_outputs(4271)) or (layer0_outputs(9807));
    outputs(658) <= not((layer0_outputs(983)) and (layer0_outputs(926)));
    outputs(659) <= not(layer0_outputs(4308)) or (layer0_outputs(6800));
    outputs(660) <= not(layer0_outputs(3252));
    outputs(661) <= (layer0_outputs(3524)) xor (layer0_outputs(6930));
    outputs(662) <= not(layer0_outputs(8050));
    outputs(663) <= (layer0_outputs(9069)) xor (layer0_outputs(5856));
    outputs(664) <= not(layer0_outputs(5232));
    outputs(665) <= not(layer0_outputs(1065));
    outputs(666) <= not(layer0_outputs(3598));
    outputs(667) <= (layer0_outputs(243)) xor (layer0_outputs(9488));
    outputs(668) <= not((layer0_outputs(5081)) and (layer0_outputs(1194)));
    outputs(669) <= layer0_outputs(3130);
    outputs(670) <= (layer0_outputs(5629)) xor (layer0_outputs(9093));
    outputs(671) <= not((layer0_outputs(3728)) and (layer0_outputs(752)));
    outputs(672) <= not(layer0_outputs(3707));
    outputs(673) <= layer0_outputs(7987);
    outputs(674) <= not(layer0_outputs(5199));
    outputs(675) <= not((layer0_outputs(9489)) and (layer0_outputs(7604)));
    outputs(676) <= not(layer0_outputs(6959));
    outputs(677) <= layer0_outputs(5428);
    outputs(678) <= not(layer0_outputs(1127));
    outputs(679) <= layer0_outputs(3502);
    outputs(680) <= (layer0_outputs(5222)) and not (layer0_outputs(133));
    outputs(681) <= (layer0_outputs(5428)) or (layer0_outputs(9984));
    outputs(682) <= not(layer0_outputs(9141));
    outputs(683) <= layer0_outputs(6868);
    outputs(684) <= (layer0_outputs(3406)) xor (layer0_outputs(2292));
    outputs(685) <= not(layer0_outputs(3146));
    outputs(686) <= layer0_outputs(2007);
    outputs(687) <= not(layer0_outputs(5655)) or (layer0_outputs(703));
    outputs(688) <= not((layer0_outputs(1907)) xor (layer0_outputs(1786)));
    outputs(689) <= (layer0_outputs(731)) and (layer0_outputs(8621));
    outputs(690) <= layer0_outputs(5557);
    outputs(691) <= not(layer0_outputs(10011));
    outputs(692) <= not(layer0_outputs(5342));
    outputs(693) <= (layer0_outputs(8479)) xor (layer0_outputs(7384));
    outputs(694) <= not(layer0_outputs(5321));
    outputs(695) <= not(layer0_outputs(5409));
    outputs(696) <= not((layer0_outputs(3387)) xor (layer0_outputs(1254)));
    outputs(697) <= layer0_outputs(5377);
    outputs(698) <= not((layer0_outputs(5)) and (layer0_outputs(2966)));
    outputs(699) <= not(layer0_outputs(1556)) or (layer0_outputs(9943));
    outputs(700) <= layer0_outputs(8765);
    outputs(701) <= layer0_outputs(1840);
    outputs(702) <= (layer0_outputs(1447)) xor (layer0_outputs(7917));
    outputs(703) <= not(layer0_outputs(7410));
    outputs(704) <= '1';
    outputs(705) <= not((layer0_outputs(3950)) xor (layer0_outputs(9822)));
    outputs(706) <= layer0_outputs(4258);
    outputs(707) <= (layer0_outputs(8180)) and (layer0_outputs(294));
    outputs(708) <= (layer0_outputs(1779)) xor (layer0_outputs(203));
    outputs(709) <= not((layer0_outputs(10129)) xor (layer0_outputs(9180)));
    outputs(710) <= not(layer0_outputs(4727));
    outputs(711) <= layer0_outputs(5084);
    outputs(712) <= (layer0_outputs(6207)) xor (layer0_outputs(8977));
    outputs(713) <= not((layer0_outputs(7578)) xor (layer0_outputs(5607)));
    outputs(714) <= layer0_outputs(8094);
    outputs(715) <= not(layer0_outputs(315));
    outputs(716) <= (layer0_outputs(6461)) xor (layer0_outputs(6299));
    outputs(717) <= (layer0_outputs(2875)) xor (layer0_outputs(1286));
    outputs(718) <= not((layer0_outputs(9543)) xor (layer0_outputs(10166)));
    outputs(719) <= not((layer0_outputs(1556)) and (layer0_outputs(105)));
    outputs(720) <= (layer0_outputs(131)) xor (layer0_outputs(9729));
    outputs(721) <= not(layer0_outputs(3838)) or (layer0_outputs(132));
    outputs(722) <= layer0_outputs(3662);
    outputs(723) <= layer0_outputs(3623);
    outputs(724) <= not((layer0_outputs(5061)) xor (layer0_outputs(742)));
    outputs(725) <= not(layer0_outputs(3682));
    outputs(726) <= (layer0_outputs(475)) or (layer0_outputs(8981));
    outputs(727) <= not((layer0_outputs(2116)) xor (layer0_outputs(273)));
    outputs(728) <= (layer0_outputs(2672)) xor (layer0_outputs(3007));
    outputs(729) <= not(layer0_outputs(1107)) or (layer0_outputs(7300));
    outputs(730) <= (layer0_outputs(9820)) or (layer0_outputs(2498));
    outputs(731) <= (layer0_outputs(9407)) xor (layer0_outputs(5289));
    outputs(732) <= not(layer0_outputs(9705)) or (layer0_outputs(2754));
    outputs(733) <= (layer0_outputs(8370)) xor (layer0_outputs(987));
    outputs(734) <= not(layer0_outputs(3833)) or (layer0_outputs(2498));
    outputs(735) <= not((layer0_outputs(6970)) xor (layer0_outputs(8970)));
    outputs(736) <= (layer0_outputs(6542)) and not (layer0_outputs(7693));
    outputs(737) <= layer0_outputs(7264);
    outputs(738) <= not(layer0_outputs(6559)) or (layer0_outputs(2281));
    outputs(739) <= not(layer0_outputs(4833));
    outputs(740) <= layer0_outputs(3576);
    outputs(741) <= (layer0_outputs(392)) and (layer0_outputs(5453));
    outputs(742) <= not(layer0_outputs(7195)) or (layer0_outputs(7038));
    outputs(743) <= (layer0_outputs(755)) xor (layer0_outputs(3189));
    outputs(744) <= not(layer0_outputs(1599)) or (layer0_outputs(8230));
    outputs(745) <= (layer0_outputs(5056)) or (layer0_outputs(3614));
    outputs(746) <= (layer0_outputs(5237)) and not (layer0_outputs(9414));
    outputs(747) <= not(layer0_outputs(10018)) or (layer0_outputs(9423));
    outputs(748) <= layer0_outputs(9252);
    outputs(749) <= not(layer0_outputs(5956)) or (layer0_outputs(7091));
    outputs(750) <= not(layer0_outputs(4671)) or (layer0_outputs(797));
    outputs(751) <= (layer0_outputs(2333)) xor (layer0_outputs(4322));
    outputs(752) <= (layer0_outputs(2713)) xor (layer0_outputs(9410));
    outputs(753) <= not(layer0_outputs(5511));
    outputs(754) <= not(layer0_outputs(843)) or (layer0_outputs(3484));
    outputs(755) <= not(layer0_outputs(6980)) or (layer0_outputs(6769));
    outputs(756) <= layer0_outputs(3994);
    outputs(757) <= not(layer0_outputs(3038));
    outputs(758) <= (layer0_outputs(6445)) xor (layer0_outputs(1262));
    outputs(759) <= not(layer0_outputs(6379));
    outputs(760) <= layer0_outputs(3179);
    outputs(761) <= not(layer0_outputs(9692));
    outputs(762) <= layer0_outputs(1792);
    outputs(763) <= not(layer0_outputs(9288)) or (layer0_outputs(10002));
    outputs(764) <= not(layer0_outputs(5169)) or (layer0_outputs(188));
    outputs(765) <= layer0_outputs(5902);
    outputs(766) <= (layer0_outputs(2580)) and not (layer0_outputs(10113));
    outputs(767) <= layer0_outputs(4583);
    outputs(768) <= layer0_outputs(1126);
    outputs(769) <= not((layer0_outputs(6092)) and (layer0_outputs(1082)));
    outputs(770) <= not(layer0_outputs(9416));
    outputs(771) <= layer0_outputs(386);
    outputs(772) <= not(layer0_outputs(5271));
    outputs(773) <= not(layer0_outputs(4672)) or (layer0_outputs(8744));
    outputs(774) <= not(layer0_outputs(8502)) or (layer0_outputs(5681));
    outputs(775) <= (layer0_outputs(3588)) xor (layer0_outputs(310));
    outputs(776) <= layer0_outputs(2470);
    outputs(777) <= not((layer0_outputs(4484)) xor (layer0_outputs(6851)));
    outputs(778) <= not(layer0_outputs(5144));
    outputs(779) <= not(layer0_outputs(5506)) or (layer0_outputs(9491));
    outputs(780) <= not(layer0_outputs(5252));
    outputs(781) <= layer0_outputs(9506);
    outputs(782) <= not((layer0_outputs(4503)) and (layer0_outputs(1423)));
    outputs(783) <= not((layer0_outputs(9917)) xor (layer0_outputs(7985)));
    outputs(784) <= not(layer0_outputs(2227));
    outputs(785) <= layer0_outputs(7056);
    outputs(786) <= layer0_outputs(1268);
    outputs(787) <= not(layer0_outputs(1722));
    outputs(788) <= layer0_outputs(9230);
    outputs(789) <= layer0_outputs(5734);
    outputs(790) <= not(layer0_outputs(718));
    outputs(791) <= not((layer0_outputs(7495)) and (layer0_outputs(7994)));
    outputs(792) <= (layer0_outputs(6982)) xor (layer0_outputs(5904));
    outputs(793) <= not(layer0_outputs(3049));
    outputs(794) <= not(layer0_outputs(2549));
    outputs(795) <= layer0_outputs(8582);
    outputs(796) <= layer0_outputs(9625);
    outputs(797) <= not(layer0_outputs(1481)) or (layer0_outputs(860));
    outputs(798) <= (layer0_outputs(6283)) and (layer0_outputs(6602));
    outputs(799) <= (layer0_outputs(6101)) xor (layer0_outputs(3169));
    outputs(800) <= layer0_outputs(1568);
    outputs(801) <= layer0_outputs(3718);
    outputs(802) <= (layer0_outputs(2616)) xor (layer0_outputs(4187));
    outputs(803) <= layer0_outputs(974);
    outputs(804) <= layer0_outputs(4059);
    outputs(805) <= layer0_outputs(8389);
    outputs(806) <= (layer0_outputs(9640)) xor (layer0_outputs(9050));
    outputs(807) <= layer0_outputs(7698);
    outputs(808) <= (layer0_outputs(1802)) xor (layer0_outputs(6361));
    outputs(809) <= (layer0_outputs(2388)) and not (layer0_outputs(378));
    outputs(810) <= not((layer0_outputs(6198)) xor (layer0_outputs(3438)));
    outputs(811) <= not(layer0_outputs(9066)) or (layer0_outputs(2886));
    outputs(812) <= not((layer0_outputs(2202)) xor (layer0_outputs(9424)));
    outputs(813) <= not(layer0_outputs(1735));
    outputs(814) <= layer0_outputs(9521);
    outputs(815) <= not(layer0_outputs(9310));
    outputs(816) <= layer0_outputs(4224);
    outputs(817) <= not(layer0_outputs(1035));
    outputs(818) <= layer0_outputs(1006);
    outputs(819) <= not(layer0_outputs(8410));
    outputs(820) <= not((layer0_outputs(2465)) xor (layer0_outputs(6377)));
    outputs(821) <= (layer0_outputs(3382)) xor (layer0_outputs(9878));
    outputs(822) <= not(layer0_outputs(1195));
    outputs(823) <= not(layer0_outputs(848));
    outputs(824) <= (layer0_outputs(1104)) xor (layer0_outputs(5003));
    outputs(825) <= not((layer0_outputs(6033)) or (layer0_outputs(4078)));
    outputs(826) <= layer0_outputs(7928);
    outputs(827) <= (layer0_outputs(5116)) and not (layer0_outputs(2402));
    outputs(828) <= layer0_outputs(1096);
    outputs(829) <= (layer0_outputs(440)) xor (layer0_outputs(1486));
    outputs(830) <= not((layer0_outputs(5810)) xor (layer0_outputs(3664)));
    outputs(831) <= not(layer0_outputs(1333)) or (layer0_outputs(4678));
    outputs(832) <= not(layer0_outputs(8864));
    outputs(833) <= not(layer0_outputs(251)) or (layer0_outputs(9855));
    outputs(834) <= not(layer0_outputs(4636));
    outputs(835) <= not(layer0_outputs(5564)) or (layer0_outputs(7395));
    outputs(836) <= layer0_outputs(1220);
    outputs(837) <= not((layer0_outputs(7267)) and (layer0_outputs(1418)));
    outputs(838) <= not(layer0_outputs(6246));
    outputs(839) <= not(layer0_outputs(2040));
    outputs(840) <= not((layer0_outputs(6219)) xor (layer0_outputs(1391)));
    outputs(841) <= not((layer0_outputs(8581)) and (layer0_outputs(3239)));
    outputs(842) <= not(layer0_outputs(7651));
    outputs(843) <= not(layer0_outputs(4590));
    outputs(844) <= layer0_outputs(6334);
    outputs(845) <= layer0_outputs(8292);
    outputs(846) <= not((layer0_outputs(7548)) xor (layer0_outputs(9237)));
    outputs(847) <= layer0_outputs(8003);
    outputs(848) <= (layer0_outputs(5411)) xor (layer0_outputs(7507));
    outputs(849) <= layer0_outputs(7550);
    outputs(850) <= (layer0_outputs(1726)) and (layer0_outputs(9013));
    outputs(851) <= not(layer0_outputs(2484)) or (layer0_outputs(738));
    outputs(852) <= (layer0_outputs(1102)) and not (layer0_outputs(3692));
    outputs(853) <= '0';
    outputs(854) <= (layer0_outputs(5913)) and (layer0_outputs(5389));
    outputs(855) <= not(layer0_outputs(10207));
    outputs(856) <= not(layer0_outputs(3171));
    outputs(857) <= not((layer0_outputs(5221)) and (layer0_outputs(5871)));
    outputs(858) <= layer0_outputs(3164);
    outputs(859) <= (layer0_outputs(3734)) xor (layer0_outputs(9598));
    outputs(860) <= layer0_outputs(6360);
    outputs(861) <= not(layer0_outputs(2441)) or (layer0_outputs(6032));
    outputs(862) <= layer0_outputs(7141);
    outputs(863) <= layer0_outputs(8161);
    outputs(864) <= layer0_outputs(10190);
    outputs(865) <= not((layer0_outputs(1643)) or (layer0_outputs(7753)));
    outputs(866) <= layer0_outputs(1501);
    outputs(867) <= (layer0_outputs(7799)) and not (layer0_outputs(1242));
    outputs(868) <= '1';
    outputs(869) <= not((layer0_outputs(8298)) xor (layer0_outputs(1642)));
    outputs(870) <= not(layer0_outputs(5277)) or (layer0_outputs(2124));
    outputs(871) <= (layer0_outputs(3481)) and not (layer0_outputs(111));
    outputs(872) <= (layer0_outputs(2470)) and not (layer0_outputs(9053));
    outputs(873) <= layer0_outputs(1168);
    outputs(874) <= layer0_outputs(1102);
    outputs(875) <= not(layer0_outputs(5156));
    outputs(876) <= (layer0_outputs(99)) and not (layer0_outputs(9996));
    outputs(877) <= (layer0_outputs(3592)) xor (layer0_outputs(5236));
    outputs(878) <= not(layer0_outputs(9763)) or (layer0_outputs(246));
    outputs(879) <= not(layer0_outputs(9368));
    outputs(880) <= not(layer0_outputs(4940)) or (layer0_outputs(4383));
    outputs(881) <= not(layer0_outputs(2660));
    outputs(882) <= not((layer0_outputs(5822)) or (layer0_outputs(3618)));
    outputs(883) <= layer0_outputs(6144);
    outputs(884) <= layer0_outputs(2055);
    outputs(885) <= layer0_outputs(6407);
    outputs(886) <= layer0_outputs(372);
    outputs(887) <= not(layer0_outputs(1397));
    outputs(888) <= not(layer0_outputs(554));
    outputs(889) <= layer0_outputs(864);
    outputs(890) <= not(layer0_outputs(532)) or (layer0_outputs(8787));
    outputs(891) <= not((layer0_outputs(2877)) xor (layer0_outputs(307)));
    outputs(892) <= layer0_outputs(8660);
    outputs(893) <= not(layer0_outputs(6441));
    outputs(894) <= (layer0_outputs(1366)) or (layer0_outputs(4015));
    outputs(895) <= (layer0_outputs(2816)) or (layer0_outputs(2647));
    outputs(896) <= not((layer0_outputs(5194)) and (layer0_outputs(3397)));
    outputs(897) <= layer0_outputs(5355);
    outputs(898) <= layer0_outputs(4786);
    outputs(899) <= not(layer0_outputs(3838)) or (layer0_outputs(10083));
    outputs(900) <= not(layer0_outputs(8647)) or (layer0_outputs(8530));
    outputs(901) <= not(layer0_outputs(10145));
    outputs(902) <= (layer0_outputs(1564)) xor (layer0_outputs(8311));
    outputs(903) <= not(layer0_outputs(7375)) or (layer0_outputs(9528));
    outputs(904) <= layer0_outputs(4045);
    outputs(905) <= not((layer0_outputs(4992)) xor (layer0_outputs(6161)));
    outputs(906) <= layer0_outputs(1858);
    outputs(907) <= not(layer0_outputs(2491));
    outputs(908) <= not((layer0_outputs(531)) or (layer0_outputs(4069)));
    outputs(909) <= not(layer0_outputs(6882)) or (layer0_outputs(170));
    outputs(910) <= not(layer0_outputs(1235));
    outputs(911) <= not(layer0_outputs(8449));
    outputs(912) <= not(layer0_outputs(8879)) or (layer0_outputs(621));
    outputs(913) <= not(layer0_outputs(2088));
    outputs(914) <= not((layer0_outputs(8548)) or (layer0_outputs(9442)));
    outputs(915) <= (layer0_outputs(2865)) xor (layer0_outputs(9066));
    outputs(916) <= layer0_outputs(6759);
    outputs(917) <= not(layer0_outputs(4797));
    outputs(918) <= not(layer0_outputs(1984));
    outputs(919) <= not(layer0_outputs(4623));
    outputs(920) <= layer0_outputs(4093);
    outputs(921) <= not(layer0_outputs(209));
    outputs(922) <= (layer0_outputs(6818)) and not (layer0_outputs(3042));
    outputs(923) <= layer0_outputs(3117);
    outputs(924) <= (layer0_outputs(5332)) and (layer0_outputs(4019));
    outputs(925) <= (layer0_outputs(9703)) and not (layer0_outputs(8275));
    outputs(926) <= (layer0_outputs(8749)) and (layer0_outputs(1038));
    outputs(927) <= not(layer0_outputs(3150));
    outputs(928) <= not(layer0_outputs(3632));
    outputs(929) <= not(layer0_outputs(6520)) or (layer0_outputs(4482));
    outputs(930) <= not(layer0_outputs(9858));
    outputs(931) <= not(layer0_outputs(7804)) or (layer0_outputs(3942));
    outputs(932) <= (layer0_outputs(8600)) xor (layer0_outputs(3862));
    outputs(933) <= not(layer0_outputs(3462));
    outputs(934) <= not(layer0_outputs(6363));
    outputs(935) <= '1';
    outputs(936) <= not(layer0_outputs(1112)) or (layer0_outputs(7714));
    outputs(937) <= not((layer0_outputs(8932)) or (layer0_outputs(8412)));
    outputs(938) <= (layer0_outputs(3898)) or (layer0_outputs(8133));
    outputs(939) <= not(layer0_outputs(4955));
    outputs(940) <= not(layer0_outputs(9920));
    outputs(941) <= layer0_outputs(10205);
    outputs(942) <= not((layer0_outputs(1554)) xor (layer0_outputs(6716)));
    outputs(943) <= (layer0_outputs(9449)) and (layer0_outputs(9454));
    outputs(944) <= not((layer0_outputs(693)) or (layer0_outputs(6794)));
    outputs(945) <= (layer0_outputs(7351)) or (layer0_outputs(3734));
    outputs(946) <= layer0_outputs(1761);
    outputs(947) <= not(layer0_outputs(9005));
    outputs(948) <= layer0_outputs(4832);
    outputs(949) <= not(layer0_outputs(3336));
    outputs(950) <= layer0_outputs(5714);
    outputs(951) <= not(layer0_outputs(1655));
    outputs(952) <= not((layer0_outputs(461)) xor (layer0_outputs(6768)));
    outputs(953) <= (layer0_outputs(2859)) xor (layer0_outputs(7907));
    outputs(954) <= not(layer0_outputs(6049));
    outputs(955) <= '1';
    outputs(956) <= (layer0_outputs(353)) and not (layer0_outputs(674));
    outputs(957) <= (layer0_outputs(3088)) and not (layer0_outputs(3161));
    outputs(958) <= not(layer0_outputs(1638));
    outputs(959) <= layer0_outputs(3941);
    outputs(960) <= layer0_outputs(7349);
    outputs(961) <= layer0_outputs(4733);
    outputs(962) <= layer0_outputs(5330);
    outputs(963) <= layer0_outputs(8278);
    outputs(964) <= (layer0_outputs(8401)) and not (layer0_outputs(838));
    outputs(965) <= layer0_outputs(5183);
    outputs(966) <= layer0_outputs(2319);
    outputs(967) <= (layer0_outputs(8987)) or (layer0_outputs(10093));
    outputs(968) <= not(layer0_outputs(2789));
    outputs(969) <= layer0_outputs(7168);
    outputs(970) <= layer0_outputs(1788);
    outputs(971) <= not((layer0_outputs(1719)) or (layer0_outputs(1130)));
    outputs(972) <= layer0_outputs(6691);
    outputs(973) <= layer0_outputs(2541);
    outputs(974) <= not(layer0_outputs(2954));
    outputs(975) <= not(layer0_outputs(9725));
    outputs(976) <= (layer0_outputs(7565)) xor (layer0_outputs(4983));
    outputs(977) <= layer0_outputs(9683);
    outputs(978) <= (layer0_outputs(905)) and (layer0_outputs(3008));
    outputs(979) <= not(layer0_outputs(9522));
    outputs(980) <= not(layer0_outputs(30));
    outputs(981) <= not(layer0_outputs(6995));
    outputs(982) <= not(layer0_outputs(7068));
    outputs(983) <= (layer0_outputs(732)) and (layer0_outputs(1769));
    outputs(984) <= not(layer0_outputs(1676));
    outputs(985) <= not(layer0_outputs(2830));
    outputs(986) <= not((layer0_outputs(9147)) xor (layer0_outputs(7340)));
    outputs(987) <= '1';
    outputs(988) <= (layer0_outputs(9171)) and not (layer0_outputs(5685));
    outputs(989) <= not(layer0_outputs(3285));
    outputs(990) <= (layer0_outputs(5451)) or (layer0_outputs(9910));
    outputs(991) <= layer0_outputs(8679);
    outputs(992) <= not(layer0_outputs(4218));
    outputs(993) <= layer0_outputs(9425);
    outputs(994) <= (layer0_outputs(5736)) and (layer0_outputs(5861));
    outputs(995) <= not(layer0_outputs(7010));
    outputs(996) <= not((layer0_outputs(9359)) xor (layer0_outputs(3392)));
    outputs(997) <= layer0_outputs(6455);
    outputs(998) <= not(layer0_outputs(3557));
    outputs(999) <= not(layer0_outputs(385));
    outputs(1000) <= (layer0_outputs(1678)) xor (layer0_outputs(2920));
    outputs(1001) <= layer0_outputs(1280);
    outputs(1002) <= not(layer0_outputs(8506));
    outputs(1003) <= (layer0_outputs(1321)) xor (layer0_outputs(7153));
    outputs(1004) <= not((layer0_outputs(496)) xor (layer0_outputs(2447)));
    outputs(1005) <= layer0_outputs(3341);
    outputs(1006) <= not(layer0_outputs(5956));
    outputs(1007) <= layer0_outputs(5637);
    outputs(1008) <= layer0_outputs(2918);
    outputs(1009) <= not(layer0_outputs(3075));
    outputs(1010) <= not(layer0_outputs(2487)) or (layer0_outputs(7174));
    outputs(1011) <= not((layer0_outputs(1057)) or (layer0_outputs(5061)));
    outputs(1012) <= (layer0_outputs(7952)) xor (layer0_outputs(319));
    outputs(1013) <= layer0_outputs(7852);
    outputs(1014) <= (layer0_outputs(4427)) xor (layer0_outputs(9778));
    outputs(1015) <= (layer0_outputs(6836)) xor (layer0_outputs(9395));
    outputs(1016) <= not((layer0_outputs(5211)) or (layer0_outputs(6080)));
    outputs(1017) <= (layer0_outputs(7550)) and (layer0_outputs(7553));
    outputs(1018) <= not((layer0_outputs(2225)) xor (layer0_outputs(4092)));
    outputs(1019) <= layer0_outputs(2238);
    outputs(1020) <= (layer0_outputs(1814)) xor (layer0_outputs(9562));
    outputs(1021) <= (layer0_outputs(9320)) and not (layer0_outputs(9501));
    outputs(1022) <= not((layer0_outputs(5543)) xor (layer0_outputs(6328)));
    outputs(1023) <= layer0_outputs(8060);
    outputs(1024) <= (layer0_outputs(9035)) and not (layer0_outputs(296));
    outputs(1025) <= not((layer0_outputs(4851)) xor (layer0_outputs(6188)));
    outputs(1026) <= '0';
    outputs(1027) <= not((layer0_outputs(3185)) or (layer0_outputs(2627)));
    outputs(1028) <= (layer0_outputs(4056)) and (layer0_outputs(9068));
    outputs(1029) <= not(layer0_outputs(1609)) or (layer0_outputs(472));
    outputs(1030) <= not((layer0_outputs(6248)) or (layer0_outputs(8061)));
    outputs(1031) <= not((layer0_outputs(3023)) or (layer0_outputs(6869)));
    outputs(1032) <= (layer0_outputs(351)) xor (layer0_outputs(1670));
    outputs(1033) <= (layer0_outputs(7063)) and (layer0_outputs(3623));
    outputs(1034) <= not(layer0_outputs(7480));
    outputs(1035) <= not(layer0_outputs(5529));
    outputs(1036) <= layer0_outputs(212);
    outputs(1037) <= not((layer0_outputs(8465)) xor (layer0_outputs(8963)));
    outputs(1038) <= (layer0_outputs(5725)) xor (layer0_outputs(6703));
    outputs(1039) <= not((layer0_outputs(1607)) or (layer0_outputs(548)));
    outputs(1040) <= (layer0_outputs(8038)) and not (layer0_outputs(8421));
    outputs(1041) <= layer0_outputs(538);
    outputs(1042) <= (layer0_outputs(5595)) and not (layer0_outputs(207));
    outputs(1043) <= not(layer0_outputs(1569));
    outputs(1044) <= '0';
    outputs(1045) <= (layer0_outputs(9464)) and not (layer0_outputs(3012));
    outputs(1046) <= not((layer0_outputs(9586)) or (layer0_outputs(6995)));
    outputs(1047) <= not(layer0_outputs(8301));
    outputs(1048) <= not((layer0_outputs(707)) xor (layer0_outputs(6086)));
    outputs(1049) <= layer0_outputs(8199);
    outputs(1050) <= layer0_outputs(142);
    outputs(1051) <= not((layer0_outputs(8091)) or (layer0_outputs(6285)));
    outputs(1052) <= (layer0_outputs(3760)) and not (layer0_outputs(6612));
    outputs(1053) <= not((layer0_outputs(8811)) and (layer0_outputs(7780)));
    outputs(1054) <= (layer0_outputs(1342)) and not (layer0_outputs(1908));
    outputs(1055) <= not((layer0_outputs(3876)) or (layer0_outputs(1671)));
    outputs(1056) <= not(layer0_outputs(2932));
    outputs(1057) <= not((layer0_outputs(7748)) or (layer0_outputs(4580)));
    outputs(1058) <= (layer0_outputs(7854)) and not (layer0_outputs(8643));
    outputs(1059) <= not((layer0_outputs(2659)) or (layer0_outputs(3317)));
    outputs(1060) <= (layer0_outputs(6778)) and not (layer0_outputs(3152));
    outputs(1061) <= (layer0_outputs(1801)) and not (layer0_outputs(8071));
    outputs(1062) <= not(layer0_outputs(316));
    outputs(1063) <= (layer0_outputs(1279)) or (layer0_outputs(7117));
    outputs(1064) <= (layer0_outputs(3069)) and (layer0_outputs(10195));
    outputs(1065) <= layer0_outputs(4532);
    outputs(1066) <= layer0_outputs(8558);
    outputs(1067) <= not(layer0_outputs(5617));
    outputs(1068) <= (layer0_outputs(535)) and (layer0_outputs(816));
    outputs(1069) <= layer0_outputs(1839);
    outputs(1070) <= layer0_outputs(4134);
    outputs(1071) <= not((layer0_outputs(4796)) or (layer0_outputs(3709)));
    outputs(1072) <= not((layer0_outputs(3376)) xor (layer0_outputs(143)));
    outputs(1073) <= layer0_outputs(5057);
    outputs(1074) <= (layer0_outputs(9734)) and not (layer0_outputs(6397));
    outputs(1075) <= not((layer0_outputs(6180)) xor (layer0_outputs(2814)));
    outputs(1076) <= (layer0_outputs(5392)) and (layer0_outputs(8002));
    outputs(1077) <= layer0_outputs(4750);
    outputs(1078) <= not((layer0_outputs(6681)) or (layer0_outputs(9848)));
    outputs(1079) <= not((layer0_outputs(2785)) xor (layer0_outputs(5313)));
    outputs(1080) <= (layer0_outputs(2344)) and (layer0_outputs(6437));
    outputs(1081) <= (layer0_outputs(9784)) and not (layer0_outputs(9887));
    outputs(1082) <= not(layer0_outputs(773));
    outputs(1083) <= not((layer0_outputs(5507)) or (layer0_outputs(1072)));
    outputs(1084) <= (layer0_outputs(8967)) and (layer0_outputs(5848));
    outputs(1085) <= not((layer0_outputs(2881)) or (layer0_outputs(4963)));
    outputs(1086) <= (layer0_outputs(5562)) xor (layer0_outputs(1526));
    outputs(1087) <= layer0_outputs(391);
    outputs(1088) <= (layer0_outputs(9239)) xor (layer0_outputs(4128));
    outputs(1089) <= '0';
    outputs(1090) <= (layer0_outputs(522)) and (layer0_outputs(6107));
    outputs(1091) <= not((layer0_outputs(7159)) xor (layer0_outputs(866)));
    outputs(1092) <= not(layer0_outputs(1450));
    outputs(1093) <= layer0_outputs(3775);
    outputs(1094) <= not((layer0_outputs(4669)) xor (layer0_outputs(2564)));
    outputs(1095) <= not((layer0_outputs(10063)) or (layer0_outputs(1008)));
    outputs(1096) <= layer0_outputs(6997);
    outputs(1097) <= (layer0_outputs(9146)) xor (layer0_outputs(8952));
    outputs(1098) <= (layer0_outputs(2231)) and not (layer0_outputs(3121));
    outputs(1099) <= (layer0_outputs(9528)) and (layer0_outputs(4377));
    outputs(1100) <= (layer0_outputs(3630)) and (layer0_outputs(4674));
    outputs(1101) <= (layer0_outputs(5647)) and (layer0_outputs(365));
    outputs(1102) <= layer0_outputs(5480);
    outputs(1103) <= (layer0_outputs(3693)) and not (layer0_outputs(6725));
    outputs(1104) <= (layer0_outputs(4774)) xor (layer0_outputs(3104));
    outputs(1105) <= (layer0_outputs(2002)) and (layer0_outputs(7219));
    outputs(1106) <= (layer0_outputs(5299)) and (layer0_outputs(374));
    outputs(1107) <= not(layer0_outputs(2727));
    outputs(1108) <= (layer0_outputs(2271)) xor (layer0_outputs(6215));
    outputs(1109) <= not((layer0_outputs(8940)) xor (layer0_outputs(1400)));
    outputs(1110) <= layer0_outputs(6623);
    outputs(1111) <= not((layer0_outputs(9027)) or (layer0_outputs(9280)));
    outputs(1112) <= not((layer0_outputs(6374)) xor (layer0_outputs(7598)));
    outputs(1113) <= (layer0_outputs(10065)) and not (layer0_outputs(4478));
    outputs(1114) <= not(layer0_outputs(1898));
    outputs(1115) <= not(layer0_outputs(6348));
    outputs(1116) <= layer0_outputs(5624);
    outputs(1117) <= (layer0_outputs(9639)) and not (layer0_outputs(9390));
    outputs(1118) <= not(layer0_outputs(1508));
    outputs(1119) <= (layer0_outputs(5508)) and not (layer0_outputs(1873));
    outputs(1120) <= '0';
    outputs(1121) <= not(layer0_outputs(8143));
    outputs(1122) <= (layer0_outputs(2067)) xor (layer0_outputs(1941));
    outputs(1123) <= not(layer0_outputs(1565));
    outputs(1124) <= layer0_outputs(4626);
    outputs(1125) <= (layer0_outputs(762)) and not (layer0_outputs(9968));
    outputs(1126) <= not(layer0_outputs(6951));
    outputs(1127) <= not((layer0_outputs(9960)) or (layer0_outputs(8572)));
    outputs(1128) <= not((layer0_outputs(3005)) or (layer0_outputs(7664)));
    outputs(1129) <= (layer0_outputs(10149)) and not (layer0_outputs(1966));
    outputs(1130) <= '0';
    outputs(1131) <= (layer0_outputs(6825)) xor (layer0_outputs(4504));
    outputs(1132) <= not(layer0_outputs(7128));
    outputs(1133) <= (layer0_outputs(8915)) xor (layer0_outputs(9125));
    outputs(1134) <= (layer0_outputs(3806)) xor (layer0_outputs(9967));
    outputs(1135) <= '0';
    outputs(1136) <= not((layer0_outputs(8022)) and (layer0_outputs(4692)));
    outputs(1137) <= not((layer0_outputs(1451)) or (layer0_outputs(2195)));
    outputs(1138) <= not(layer0_outputs(5990));
    outputs(1139) <= '0';
    outputs(1140) <= not((layer0_outputs(2276)) or (layer0_outputs(9506)));
    outputs(1141) <= not(layer0_outputs(9130));
    outputs(1142) <= not(layer0_outputs(8610));
    outputs(1143) <= not((layer0_outputs(181)) or (layer0_outputs(4732)));
    outputs(1144) <= not((layer0_outputs(743)) or (layer0_outputs(9067)));
    outputs(1145) <= (layer0_outputs(9221)) and not (layer0_outputs(1008));
    outputs(1146) <= not((layer0_outputs(8283)) or (layer0_outputs(2802)));
    outputs(1147) <= '0';
    outputs(1148) <= (layer0_outputs(3158)) and not (layer0_outputs(4112));
    outputs(1149) <= (layer0_outputs(7904)) xor (layer0_outputs(3287));
    outputs(1150) <= not(layer0_outputs(6503));
    outputs(1151) <= not(layer0_outputs(5955));
    outputs(1152) <= not(layer0_outputs(7080));
    outputs(1153) <= (layer0_outputs(6910)) and not (layer0_outputs(5406));
    outputs(1154) <= not((layer0_outputs(2035)) xor (layer0_outputs(1075)));
    outputs(1155) <= layer0_outputs(8742);
    outputs(1156) <= layer0_outputs(9370);
    outputs(1157) <= not((layer0_outputs(2453)) xor (layer0_outputs(3484)));
    outputs(1158) <= layer0_outputs(267);
    outputs(1159) <= not((layer0_outputs(1945)) or (layer0_outputs(10050)));
    outputs(1160) <= not((layer0_outputs(662)) xor (layer0_outputs(3045)));
    outputs(1161) <= (layer0_outputs(4246)) and (layer0_outputs(4456));
    outputs(1162) <= (layer0_outputs(8393)) and not (layer0_outputs(6037));
    outputs(1163) <= layer0_outputs(4549);
    outputs(1164) <= not(layer0_outputs(8516));
    outputs(1165) <= (layer0_outputs(5040)) and not (layer0_outputs(6045));
    outputs(1166) <= layer0_outputs(8911);
    outputs(1167) <= layer0_outputs(2737);
    outputs(1168) <= not((layer0_outputs(8771)) or (layer0_outputs(9111)));
    outputs(1169) <= (layer0_outputs(7474)) and (layer0_outputs(3290));
    outputs(1170) <= (layer0_outputs(9810)) and not (layer0_outputs(9281));
    outputs(1171) <= (layer0_outputs(8216)) and not (layer0_outputs(10132));
    outputs(1172) <= not((layer0_outputs(7315)) xor (layer0_outputs(2977)));
    outputs(1173) <= (layer0_outputs(3244)) and not (layer0_outputs(7045));
    outputs(1174) <= '0';
    outputs(1175) <= not(layer0_outputs(3494)) or (layer0_outputs(3266));
    outputs(1176) <= layer0_outputs(6676);
    outputs(1177) <= (layer0_outputs(7003)) and not (layer0_outputs(6686));
    outputs(1178) <= not((layer0_outputs(7291)) or (layer0_outputs(3495)));
    outputs(1179) <= not(layer0_outputs(4052));
    outputs(1180) <= not(layer0_outputs(748));
    outputs(1181) <= not((layer0_outputs(3765)) or (layer0_outputs(2917)));
    outputs(1182) <= not(layer0_outputs(5380));
    outputs(1183) <= (layer0_outputs(49)) xor (layer0_outputs(997));
    outputs(1184) <= (layer0_outputs(7452)) xor (layer0_outputs(781));
    outputs(1185) <= (layer0_outputs(487)) and not (layer0_outputs(1430));
    outputs(1186) <= (layer0_outputs(900)) and not (layer0_outputs(9094));
    outputs(1187) <= not((layer0_outputs(3650)) xor (layer0_outputs(2282)));
    outputs(1188) <= not(layer0_outputs(373));
    outputs(1189) <= not((layer0_outputs(3068)) or (layer0_outputs(7656)));
    outputs(1190) <= (layer0_outputs(6337)) xor (layer0_outputs(4180));
    outputs(1191) <= (layer0_outputs(7462)) and not (layer0_outputs(1015));
    outputs(1192) <= (layer0_outputs(9326)) and (layer0_outputs(5077));
    outputs(1193) <= (layer0_outputs(9074)) and (layer0_outputs(155));
    outputs(1194) <= not((layer0_outputs(69)) xor (layer0_outputs(3225)));
    outputs(1195) <= (layer0_outputs(4775)) and not (layer0_outputs(3549));
    outputs(1196) <= not((layer0_outputs(7966)) or (layer0_outputs(7752)));
    outputs(1197) <= (layer0_outputs(6838)) and not (layer0_outputs(8057));
    outputs(1198) <= not(layer0_outputs(1851));
    outputs(1199) <= layer0_outputs(3725);
    outputs(1200) <= not((layer0_outputs(7020)) or (layer0_outputs(4290)));
    outputs(1201) <= layer0_outputs(4960);
    outputs(1202) <= not((layer0_outputs(2758)) or (layer0_outputs(2971)));
    outputs(1203) <= (layer0_outputs(8920)) and not (layer0_outputs(3257));
    outputs(1204) <= not((layer0_outputs(6085)) or (layer0_outputs(6562)));
    outputs(1205) <= (layer0_outputs(5180)) and not (layer0_outputs(585));
    outputs(1206) <= not((layer0_outputs(863)) or (layer0_outputs(1005)));
    outputs(1207) <= layer0_outputs(6062);
    outputs(1208) <= not((layer0_outputs(9054)) or (layer0_outputs(8866)));
    outputs(1209) <= layer0_outputs(9606);
    outputs(1210) <= layer0_outputs(3782);
    outputs(1211) <= not((layer0_outputs(9934)) or (layer0_outputs(5680)));
    outputs(1212) <= (layer0_outputs(5739)) and not (layer0_outputs(8126));
    outputs(1213) <= not((layer0_outputs(3595)) or (layer0_outputs(1335)));
    outputs(1214) <= layer0_outputs(5323);
    outputs(1215) <= (layer0_outputs(6472)) xor (layer0_outputs(6187));
    outputs(1216) <= (layer0_outputs(6270)) xor (layer0_outputs(2091));
    outputs(1217) <= (layer0_outputs(5055)) xor (layer0_outputs(3751));
    outputs(1218) <= not((layer0_outputs(9698)) or (layer0_outputs(1202)));
    outputs(1219) <= not(layer0_outputs(2824));
    outputs(1220) <= not((layer0_outputs(6944)) or (layer0_outputs(6001)));
    outputs(1221) <= (layer0_outputs(8008)) xor (layer0_outputs(238));
    outputs(1222) <= (layer0_outputs(8328)) or (layer0_outputs(8244));
    outputs(1223) <= not((layer0_outputs(9724)) and (layer0_outputs(5950)));
    outputs(1224) <= (layer0_outputs(7198)) and not (layer0_outputs(3491));
    outputs(1225) <= not((layer0_outputs(5127)) or (layer0_outputs(9457)));
    outputs(1226) <= layer0_outputs(7720);
    outputs(1227) <= (layer0_outputs(9217)) xor (layer0_outputs(3236));
    outputs(1228) <= (layer0_outputs(6211)) and not (layer0_outputs(4836));
    outputs(1229) <= (layer0_outputs(3897)) and not (layer0_outputs(3073));
    outputs(1230) <= not(layer0_outputs(548));
    outputs(1231) <= '0';
    outputs(1232) <= layer0_outputs(8474);
    outputs(1233) <= (layer0_outputs(4664)) xor (layer0_outputs(3741));
    outputs(1234) <= (layer0_outputs(6979)) and not (layer0_outputs(6892));
    outputs(1235) <= layer0_outputs(251);
    outputs(1236) <= not((layer0_outputs(954)) and (layer0_outputs(3261)));
    outputs(1237) <= (layer0_outputs(3078)) xor (layer0_outputs(7110));
    outputs(1238) <= layer0_outputs(9240);
    outputs(1239) <= not((layer0_outputs(7934)) xor (layer0_outputs(5195)));
    outputs(1240) <= not((layer0_outputs(7139)) xor (layer0_outputs(6411)));
    outputs(1241) <= not((layer0_outputs(2044)) xor (layer0_outputs(5824)));
    outputs(1242) <= (layer0_outputs(1949)) and not (layer0_outputs(444));
    outputs(1243) <= (layer0_outputs(3826)) and (layer0_outputs(3471));
    outputs(1244) <= (layer0_outputs(507)) and not (layer0_outputs(5840));
    outputs(1245) <= not((layer0_outputs(5888)) xor (layer0_outputs(3185)));
    outputs(1246) <= '0';
    outputs(1247) <= layer0_outputs(4005);
    outputs(1248) <= layer0_outputs(1201);
    outputs(1249) <= (layer0_outputs(4773)) and not (layer0_outputs(6506));
    outputs(1250) <= not(layer0_outputs(8430));
    outputs(1251) <= layer0_outputs(2823);
    outputs(1252) <= (layer0_outputs(7069)) and (layer0_outputs(5045));
    outputs(1253) <= not((layer0_outputs(7345)) xor (layer0_outputs(750)));
    outputs(1254) <= layer0_outputs(6550);
    outputs(1255) <= not((layer0_outputs(6647)) xor (layer0_outputs(203)));
    outputs(1256) <= layer0_outputs(7271);
    outputs(1257) <= (layer0_outputs(6145)) and not (layer0_outputs(578));
    outputs(1258) <= not((layer0_outputs(3338)) or (layer0_outputs(8085)));
    outputs(1259) <= not((layer0_outputs(8562)) xor (layer0_outputs(9808)));
    outputs(1260) <= (layer0_outputs(7745)) and not (layer0_outputs(8009));
    outputs(1261) <= layer0_outputs(2157);
    outputs(1262) <= not((layer0_outputs(9036)) and (layer0_outputs(8177)));
    outputs(1263) <= not(layer0_outputs(7973));
    outputs(1264) <= not((layer0_outputs(8052)) or (layer0_outputs(6488)));
    outputs(1265) <= not(layer0_outputs(7915));
    outputs(1266) <= layer0_outputs(4935);
    outputs(1267) <= not((layer0_outputs(5294)) xor (layer0_outputs(4076)));
    outputs(1268) <= (layer0_outputs(7558)) and not (layer0_outputs(2279));
    outputs(1269) <= not((layer0_outputs(10047)) or (layer0_outputs(2918)));
    outputs(1270) <= not((layer0_outputs(3810)) or (layer0_outputs(8782)));
    outputs(1271) <= (layer0_outputs(1474)) and not (layer0_outputs(4717));
    outputs(1272) <= layer0_outputs(5136);
    outputs(1273) <= layer0_outputs(8016);
    outputs(1274) <= not(layer0_outputs(4735)) or (layer0_outputs(1682));
    outputs(1275) <= (layer0_outputs(8480)) xor (layer0_outputs(3796));
    outputs(1276) <= not(layer0_outputs(22));
    outputs(1277) <= not((layer0_outputs(5111)) xor (layer0_outputs(7405)));
    outputs(1278) <= '0';
    outputs(1279) <= layer0_outputs(807);
    outputs(1280) <= layer0_outputs(9559);
    outputs(1281) <= layer0_outputs(6877);
    outputs(1282) <= (layer0_outputs(6396)) xor (layer0_outputs(279));
    outputs(1283) <= layer0_outputs(291);
    outputs(1284) <= layer0_outputs(2145);
    outputs(1285) <= not((layer0_outputs(5336)) or (layer0_outputs(7431)));
    outputs(1286) <= layer0_outputs(2214);
    outputs(1287) <= (layer0_outputs(3212)) and not (layer0_outputs(9869));
    outputs(1288) <= layer0_outputs(6886);
    outputs(1289) <= layer0_outputs(6323);
    outputs(1290) <= (layer0_outputs(6295)) and not (layer0_outputs(4698));
    outputs(1291) <= (layer0_outputs(9871)) and not (layer0_outputs(8058));
    outputs(1292) <= (layer0_outputs(6417)) and (layer0_outputs(3412));
    outputs(1293) <= not(layer0_outputs(6516));
    outputs(1294) <= layer0_outputs(3918);
    outputs(1295) <= layer0_outputs(2572);
    outputs(1296) <= (layer0_outputs(4127)) and not (layer0_outputs(7008));
    outputs(1297) <= not((layer0_outputs(1396)) xor (layer0_outputs(530)));
    outputs(1298) <= layer0_outputs(2813);
    outputs(1299) <= (layer0_outputs(6169)) and not (layer0_outputs(4488));
    outputs(1300) <= layer0_outputs(3354);
    outputs(1301) <= not(layer0_outputs(1538));
    outputs(1302) <= (layer0_outputs(6726)) xor (layer0_outputs(7883));
    outputs(1303) <= (layer0_outputs(194)) xor (layer0_outputs(9494));
    outputs(1304) <= '0';
    outputs(1305) <= (layer0_outputs(9697)) and not (layer0_outputs(3717));
    outputs(1306) <= (layer0_outputs(2600)) and not (layer0_outputs(2106));
    outputs(1307) <= (layer0_outputs(10220)) and not (layer0_outputs(515));
    outputs(1308) <= (layer0_outputs(2828)) and not (layer0_outputs(3927));
    outputs(1309) <= not((layer0_outputs(2550)) or (layer0_outputs(4057)));
    outputs(1310) <= layer0_outputs(7553);
    outputs(1311) <= layer0_outputs(953);
    outputs(1312) <= (layer0_outputs(6062)) and not (layer0_outputs(4888));
    outputs(1313) <= (layer0_outputs(4835)) and (layer0_outputs(7162));
    outputs(1314) <= (layer0_outputs(5364)) xor (layer0_outputs(2471));
    outputs(1315) <= (layer0_outputs(2095)) and not (layer0_outputs(4232));
    outputs(1316) <= (layer0_outputs(8586)) and (layer0_outputs(2635));
    outputs(1317) <= layer0_outputs(2956);
    outputs(1318) <= (layer0_outputs(6316)) xor (layer0_outputs(3413));
    outputs(1319) <= not(layer0_outputs(101));
    outputs(1320) <= (layer0_outputs(7797)) and not (layer0_outputs(4071));
    outputs(1321) <= layer0_outputs(2379);
    outputs(1322) <= not((layer0_outputs(9787)) or (layer0_outputs(6300)));
    outputs(1323) <= (layer0_outputs(6580)) xor (layer0_outputs(1434));
    outputs(1324) <= not((layer0_outputs(3235)) or (layer0_outputs(7939)));
    outputs(1325) <= (layer0_outputs(1526)) xor (layer0_outputs(7842));
    outputs(1326) <= layer0_outputs(171);
    outputs(1327) <= (layer0_outputs(7546)) and (layer0_outputs(8858));
    outputs(1328) <= (layer0_outputs(7990)) and (layer0_outputs(5226));
    outputs(1329) <= not((layer0_outputs(6074)) xor (layer0_outputs(3533)));
    outputs(1330) <= layer0_outputs(3209);
    outputs(1331) <= (layer0_outputs(5517)) and not (layer0_outputs(793));
    outputs(1332) <= (layer0_outputs(9475)) and not (layer0_outputs(911));
    outputs(1333) <= not(layer0_outputs(9287));
    outputs(1334) <= (layer0_outputs(7029)) and not (layer0_outputs(6920));
    outputs(1335) <= layer0_outputs(4071);
    outputs(1336) <= (layer0_outputs(5524)) and (layer0_outputs(6485));
    outputs(1337) <= not((layer0_outputs(4043)) or (layer0_outputs(1524)));
    outputs(1338) <= (layer0_outputs(4513)) and (layer0_outputs(4301));
    outputs(1339) <= '0';
    outputs(1340) <= not(layer0_outputs(2522));
    outputs(1341) <= not(layer0_outputs(8210));
    outputs(1342) <= layer0_outputs(8007);
    outputs(1343) <= layer0_outputs(8201);
    outputs(1344) <= layer0_outputs(4404);
    outputs(1345) <= (layer0_outputs(5440)) and not (layer0_outputs(1840));
    outputs(1346) <= not((layer0_outputs(9034)) or (layer0_outputs(8819)));
    outputs(1347) <= not(layer0_outputs(6374));
    outputs(1348) <= (layer0_outputs(7286)) and not (layer0_outputs(8441));
    outputs(1349) <= (layer0_outputs(9705)) and not (layer0_outputs(3433));
    outputs(1350) <= (layer0_outputs(5807)) and (layer0_outputs(7474));
    outputs(1351) <= (layer0_outputs(1730)) or (layer0_outputs(6529));
    outputs(1352) <= not(layer0_outputs(4089));
    outputs(1353) <= (layer0_outputs(1491)) and not (layer0_outputs(3059));
    outputs(1354) <= (layer0_outputs(9220)) and not (layer0_outputs(5404));
    outputs(1355) <= (layer0_outputs(6698)) and not (layer0_outputs(6335));
    outputs(1356) <= layer0_outputs(7877);
    outputs(1357) <= layer0_outputs(3265);
    outputs(1358) <= (layer0_outputs(8722)) and not (layer0_outputs(5600));
    outputs(1359) <= (layer0_outputs(7437)) and not (layer0_outputs(2848));
    outputs(1360) <= (layer0_outputs(2782)) xor (layer0_outputs(901));
    outputs(1361) <= (layer0_outputs(5067)) and not (layer0_outputs(8445));
    outputs(1362) <= '0';
    outputs(1363) <= '0';
    outputs(1364) <= (layer0_outputs(2868)) and not (layer0_outputs(1437));
    outputs(1365) <= '0';
    outputs(1366) <= (layer0_outputs(357)) and (layer0_outputs(3190));
    outputs(1367) <= (layer0_outputs(7247)) and not (layer0_outputs(749));
    outputs(1368) <= not(layer0_outputs(144));
    outputs(1369) <= '0';
    outputs(1370) <= layer0_outputs(10187);
    outputs(1371) <= (layer0_outputs(4452)) and not (layer0_outputs(3902));
    outputs(1372) <= (layer0_outputs(1027)) and (layer0_outputs(9194));
    outputs(1373) <= (layer0_outputs(4574)) and not (layer0_outputs(8607));
    outputs(1374) <= not(layer0_outputs(1745));
    outputs(1375) <= (layer0_outputs(6061)) and not (layer0_outputs(855));
    outputs(1376) <= not((layer0_outputs(1700)) xor (layer0_outputs(9602)));
    outputs(1377) <= not(layer0_outputs(5216));
    outputs(1378) <= (layer0_outputs(660)) and not (layer0_outputs(10111));
    outputs(1379) <= (layer0_outputs(1748)) xor (layer0_outputs(9609));
    outputs(1380) <= not(layer0_outputs(564));
    outputs(1381) <= not(layer0_outputs(1160));
    outputs(1382) <= not(layer0_outputs(2012));
    outputs(1383) <= (layer0_outputs(7557)) and (layer0_outputs(2030));
    outputs(1384) <= layer0_outputs(6223);
    outputs(1385) <= (layer0_outputs(2862)) xor (layer0_outputs(4402));
    outputs(1386) <= not(layer0_outputs(2571));
    outputs(1387) <= (layer0_outputs(4674)) and not (layer0_outputs(6769));
    outputs(1388) <= (layer0_outputs(3106)) xor (layer0_outputs(7465));
    outputs(1389) <= (layer0_outputs(9656)) xor (layer0_outputs(2305));
    outputs(1390) <= layer0_outputs(148);
    outputs(1391) <= (layer0_outputs(4476)) and not (layer0_outputs(8958));
    outputs(1392) <= layer0_outputs(8548);
    outputs(1393) <= not(layer0_outputs(1427)) or (layer0_outputs(6076));
    outputs(1394) <= (layer0_outputs(949)) and (layer0_outputs(9440));
    outputs(1395) <= not(layer0_outputs(6733));
    outputs(1396) <= (layer0_outputs(7236)) and not (layer0_outputs(4350));
    outputs(1397) <= not((layer0_outputs(7625)) or (layer0_outputs(6060)));
    outputs(1398) <= (layer0_outputs(5117)) and not (layer0_outputs(4407));
    outputs(1399) <= (layer0_outputs(6104)) and (layer0_outputs(5259));
    outputs(1400) <= not((layer0_outputs(3892)) xor (layer0_outputs(1431)));
    outputs(1401) <= (layer0_outputs(10178)) and not (layer0_outputs(3697));
    outputs(1402) <= (layer0_outputs(3969)) xor (layer0_outputs(9343));
    outputs(1403) <= not(layer0_outputs(6108));
    outputs(1404) <= (layer0_outputs(8297)) and not (layer0_outputs(3515));
    outputs(1405) <= not((layer0_outputs(7530)) xor (layer0_outputs(868)));
    outputs(1406) <= not(layer0_outputs(5165));
    outputs(1407) <= layer0_outputs(2677);
    outputs(1408) <= layer0_outputs(3355);
    outputs(1409) <= not(layer0_outputs(4170));
    outputs(1410) <= (layer0_outputs(3465)) and (layer0_outputs(6658));
    outputs(1411) <= (layer0_outputs(7598)) xor (layer0_outputs(6088));
    outputs(1412) <= not((layer0_outputs(3747)) or (layer0_outputs(4806)));
    outputs(1413) <= '0';
    outputs(1414) <= (layer0_outputs(304)) xor (layer0_outputs(3224));
    outputs(1415) <= not((layer0_outputs(7657)) xor (layer0_outputs(6422)));
    outputs(1416) <= layer0_outputs(6626);
    outputs(1417) <= (layer0_outputs(8999)) and not (layer0_outputs(6494));
    outputs(1418) <= not(layer0_outputs(2915));
    outputs(1419) <= (layer0_outputs(7231)) and (layer0_outputs(2026));
    outputs(1420) <= layer0_outputs(6442);
    outputs(1421) <= not((layer0_outputs(1453)) or (layer0_outputs(9631)));
    outputs(1422) <= (layer0_outputs(7631)) and not (layer0_outputs(7393));
    outputs(1423) <= not((layer0_outputs(10124)) xor (layer0_outputs(6090)));
    outputs(1424) <= (layer0_outputs(6705)) xor (layer0_outputs(9491));
    outputs(1425) <= (layer0_outputs(7310)) and not (layer0_outputs(6143));
    outputs(1426) <= layer0_outputs(5030);
    outputs(1427) <= (layer0_outputs(7601)) and (layer0_outputs(7172));
    outputs(1428) <= (layer0_outputs(10161)) and (layer0_outputs(8383));
    outputs(1429) <= not((layer0_outputs(3478)) xor (layer0_outputs(6381)));
    outputs(1430) <= not((layer0_outputs(37)) xor (layer0_outputs(5696)));
    outputs(1431) <= (layer0_outputs(2978)) and not (layer0_outputs(5635));
    outputs(1432) <= not(layer0_outputs(4475));
    outputs(1433) <= (layer0_outputs(457)) xor (layer0_outputs(8390));
    outputs(1434) <= not((layer0_outputs(6212)) xor (layer0_outputs(2260)));
    outputs(1435) <= (layer0_outputs(7595)) and (layer0_outputs(9718));
    outputs(1436) <= not(layer0_outputs(53));
    outputs(1437) <= (layer0_outputs(6971)) and (layer0_outputs(8314));
    outputs(1438) <= layer0_outputs(8627);
    outputs(1439) <= not(layer0_outputs(3634));
    outputs(1440) <= not(layer0_outputs(6736));
    outputs(1441) <= not(layer0_outputs(4293));
    outputs(1442) <= (layer0_outputs(2552)) and not (layer0_outputs(9116));
    outputs(1443) <= not(layer0_outputs(6942));
    outputs(1444) <= '0';
    outputs(1445) <= (layer0_outputs(6128)) xor (layer0_outputs(252));
    outputs(1446) <= not((layer0_outputs(9135)) xor (layer0_outputs(3796)));
    outputs(1447) <= (layer0_outputs(9468)) and (layer0_outputs(8824));
    outputs(1448) <= not((layer0_outputs(7354)) xor (layer0_outputs(1722)));
    outputs(1449) <= (layer0_outputs(7309)) and (layer0_outputs(3784));
    outputs(1450) <= not((layer0_outputs(654)) xor (layer0_outputs(1033)));
    outputs(1451) <= not((layer0_outputs(8959)) xor (layer0_outputs(2541)));
    outputs(1452) <= not(layer0_outputs(9096));
    outputs(1453) <= layer0_outputs(1296);
    outputs(1454) <= (layer0_outputs(7212)) xor (layer0_outputs(7965));
    outputs(1455) <= layer0_outputs(1210);
    outputs(1456) <= not((layer0_outputs(9438)) or (layer0_outputs(4011)));
    outputs(1457) <= not(layer0_outputs(7267));
    outputs(1458) <= layer0_outputs(7855);
    outputs(1459) <= layer0_outputs(6067);
    outputs(1460) <= not((layer0_outputs(8147)) or (layer0_outputs(2210)));
    outputs(1461) <= (layer0_outputs(3923)) and not (layer0_outputs(5408));
    outputs(1462) <= (layer0_outputs(9852)) and not (layer0_outputs(10123));
    outputs(1463) <= (layer0_outputs(2441)) and (layer0_outputs(306));
    outputs(1464) <= (layer0_outputs(5728)) or (layer0_outputs(3835));
    outputs(1465) <= not(layer0_outputs(6748));
    outputs(1466) <= not(layer0_outputs(5492));
    outputs(1467) <= not(layer0_outputs(5112));
    outputs(1468) <= (layer0_outputs(8995)) and not (layer0_outputs(5275));
    outputs(1469) <= (layer0_outputs(3119)) or (layer0_outputs(1056));
    outputs(1470) <= layer0_outputs(6597);
    outputs(1471) <= not((layer0_outputs(8784)) or (layer0_outputs(6653)));
    outputs(1472) <= (layer0_outputs(4308)) and not (layer0_outputs(2837));
    outputs(1473) <= not((layer0_outputs(1222)) or (layer0_outputs(5012)));
    outputs(1474) <= not((layer0_outputs(2998)) or (layer0_outputs(8378)));
    outputs(1475) <= (layer0_outputs(10017)) and not (layer0_outputs(9109));
    outputs(1476) <= not((layer0_outputs(1655)) or (layer0_outputs(7541)));
    outputs(1477) <= not(layer0_outputs(3518));
    outputs(1478) <= not(layer0_outputs(6097));
    outputs(1479) <= not(layer0_outputs(9691));
    outputs(1480) <= (layer0_outputs(4007)) xor (layer0_outputs(7789));
    outputs(1481) <= (layer0_outputs(2768)) and (layer0_outputs(4853));
    outputs(1482) <= not(layer0_outputs(4500));
    outputs(1483) <= not((layer0_outputs(6058)) or (layer0_outputs(6844)));
    outputs(1484) <= (layer0_outputs(5392)) and not (layer0_outputs(7868));
    outputs(1485) <= layer0_outputs(7025);
    outputs(1486) <= layer0_outputs(8020);
    outputs(1487) <= (layer0_outputs(2268)) and not (layer0_outputs(7051));
    outputs(1488) <= not(layer0_outputs(7408));
    outputs(1489) <= (layer0_outputs(1637)) xor (layer0_outputs(8954));
    outputs(1490) <= layer0_outputs(6235);
    outputs(1491) <= not((layer0_outputs(99)) xor (layer0_outputs(567)));
    outputs(1492) <= not((layer0_outputs(6373)) or (layer0_outputs(1747)));
    outputs(1493) <= not((layer0_outputs(942)) or (layer0_outputs(1257)));
    outputs(1494) <= not(layer0_outputs(3006));
    outputs(1495) <= (layer0_outputs(3878)) and (layer0_outputs(8655));
    outputs(1496) <= not((layer0_outputs(10014)) or (layer0_outputs(8231)));
    outputs(1497) <= (layer0_outputs(9771)) and not (layer0_outputs(7547));
    outputs(1498) <= (layer0_outputs(8552)) and not (layer0_outputs(9545));
    outputs(1499) <= layer0_outputs(1349);
    outputs(1500) <= not(layer0_outputs(9190));
    outputs(1501) <= not((layer0_outputs(6036)) or (layer0_outputs(3931)));
    outputs(1502) <= layer0_outputs(642);
    outputs(1503) <= not((layer0_outputs(7611)) xor (layer0_outputs(9951)));
    outputs(1504) <= (layer0_outputs(3811)) and not (layer0_outputs(533));
    outputs(1505) <= not((layer0_outputs(2636)) or (layer0_outputs(2156)));
    outputs(1506) <= (layer0_outputs(3084)) and not (layer0_outputs(1143));
    outputs(1507) <= not(layer0_outputs(9486));
    outputs(1508) <= layer0_outputs(1176);
    outputs(1509) <= layer0_outputs(4648);
    outputs(1510) <= layer0_outputs(9129);
    outputs(1511) <= not(layer0_outputs(5614));
    outputs(1512) <= not(layer0_outputs(5507));
    outputs(1513) <= not((layer0_outputs(10112)) xor (layer0_outputs(6782)));
    outputs(1514) <= '0';
    outputs(1515) <= (layer0_outputs(6004)) and (layer0_outputs(577));
    outputs(1516) <= not(layer0_outputs(2864));
    outputs(1517) <= layer0_outputs(2039);
    outputs(1518) <= (layer0_outputs(345)) and (layer0_outputs(6911));
    outputs(1519) <= not(layer0_outputs(7913));
    outputs(1520) <= (layer0_outputs(1330)) and (layer0_outputs(2894));
    outputs(1521) <= not(layer0_outputs(4293));
    outputs(1522) <= not((layer0_outputs(1622)) xor (layer0_outputs(8619)));
    outputs(1523) <= not(layer0_outputs(8725));
    outputs(1524) <= (layer0_outputs(4078)) and not (layer0_outputs(7252));
    outputs(1525) <= not((layer0_outputs(667)) or (layer0_outputs(9419)));
    outputs(1526) <= (layer0_outputs(10048)) xor (layer0_outputs(3024));
    outputs(1527) <= not((layer0_outputs(6228)) or (layer0_outputs(84)));
    outputs(1528) <= (layer0_outputs(9861)) xor (layer0_outputs(7093));
    outputs(1529) <= not(layer0_outputs(1510));
    outputs(1530) <= (layer0_outputs(4926)) and not (layer0_outputs(9739));
    outputs(1531) <= (layer0_outputs(7445)) xor (layer0_outputs(3823));
    outputs(1532) <= layer0_outputs(2847);
    outputs(1533) <= layer0_outputs(6369);
    outputs(1534) <= not(layer0_outputs(9751));
    outputs(1535) <= layer0_outputs(4741);
    outputs(1536) <= (layer0_outputs(4088)) xor (layer0_outputs(6590));
    outputs(1537) <= layer0_outputs(10156);
    outputs(1538) <= not(layer0_outputs(3561));
    outputs(1539) <= not(layer0_outputs(7277));
    outputs(1540) <= layer0_outputs(9555);
    outputs(1541) <= layer0_outputs(887);
    outputs(1542) <= not((layer0_outputs(678)) xor (layer0_outputs(8599)));
    outputs(1543) <= not(layer0_outputs(3845));
    outputs(1544) <= layer0_outputs(5226);
    outputs(1545) <= layer0_outputs(6013);
    outputs(1546) <= not((layer0_outputs(1860)) or (layer0_outputs(2146)));
    outputs(1547) <= layer0_outputs(1960);
    outputs(1548) <= not(layer0_outputs(5614));
    outputs(1549) <= not(layer0_outputs(5855));
    outputs(1550) <= not((layer0_outputs(5547)) or (layer0_outputs(1431)));
    outputs(1551) <= layer0_outputs(1210);
    outputs(1552) <= layer0_outputs(8698);
    outputs(1553) <= layer0_outputs(84);
    outputs(1554) <= not((layer0_outputs(7764)) or (layer0_outputs(2921)));
    outputs(1555) <= '0';
    outputs(1556) <= not(layer0_outputs(4290));
    outputs(1557) <= (layer0_outputs(4614)) and (layer0_outputs(2436));
    outputs(1558) <= (layer0_outputs(281)) and not (layer0_outputs(2320));
    outputs(1559) <= not((layer0_outputs(2690)) or (layer0_outputs(2266)));
    outputs(1560) <= (layer0_outputs(3827)) and not (layer0_outputs(1982));
    outputs(1561) <= not((layer0_outputs(7870)) or (layer0_outputs(10202)));
    outputs(1562) <= (layer0_outputs(5859)) and (layer0_outputs(1310));
    outputs(1563) <= not((layer0_outputs(6638)) or (layer0_outputs(9499)));
    outputs(1564) <= (layer0_outputs(3269)) and not (layer0_outputs(416));
    outputs(1565) <= not((layer0_outputs(5987)) or (layer0_outputs(9541)));
    outputs(1566) <= not(layer0_outputs(2761)) or (layer0_outputs(4852));
    outputs(1567) <= (layer0_outputs(7744)) xor (layer0_outputs(9622));
    outputs(1568) <= layer0_outputs(6653);
    outputs(1569) <= (layer0_outputs(9108)) and not (layer0_outputs(8456));
    outputs(1570) <= layer0_outputs(1580);
    outputs(1571) <= (layer0_outputs(8948)) and not (layer0_outputs(7997));
    outputs(1572) <= (layer0_outputs(6142)) and not (layer0_outputs(6281));
    outputs(1573) <= (layer0_outputs(4070)) and (layer0_outputs(221));
    outputs(1574) <= (layer0_outputs(9380)) and not (layer0_outputs(7215));
    outputs(1575) <= (layer0_outputs(593)) and not (layer0_outputs(6002));
    outputs(1576) <= layer0_outputs(6172);
    outputs(1577) <= not(layer0_outputs(4209));
    outputs(1578) <= layer0_outputs(9364);
    outputs(1579) <= not((layer0_outputs(8702)) xor (layer0_outputs(8458)));
    outputs(1580) <= not(layer0_outputs(10100));
    outputs(1581) <= layer0_outputs(3121);
    outputs(1582) <= (layer0_outputs(1715)) and (layer0_outputs(5039));
    outputs(1583) <= (layer0_outputs(4353)) and not (layer0_outputs(6592));
    outputs(1584) <= (layer0_outputs(2668)) xor (layer0_outputs(4142));
    outputs(1585) <= (layer0_outputs(7312)) and not (layer0_outputs(6112));
    outputs(1586) <= (layer0_outputs(5400)) xor (layer0_outputs(4630));
    outputs(1587) <= (layer0_outputs(221)) and not (layer0_outputs(7199));
    outputs(1588) <= (layer0_outputs(9262)) xor (layer0_outputs(8589));
    outputs(1589) <= not(layer0_outputs(1063));
    outputs(1590) <= not(layer0_outputs(6981));
    outputs(1591) <= (layer0_outputs(7953)) and not (layer0_outputs(4858));
    outputs(1592) <= (layer0_outputs(8311)) xor (layer0_outputs(6110));
    outputs(1593) <= not(layer0_outputs(9275));
    outputs(1594) <= (layer0_outputs(7101)) and not (layer0_outputs(5344));
    outputs(1595) <= not(layer0_outputs(9276));
    outputs(1596) <= (layer0_outputs(2418)) and not (layer0_outputs(9160));
    outputs(1597) <= not((layer0_outputs(8381)) or (layer0_outputs(467)));
    outputs(1598) <= not((layer0_outputs(1227)) or (layer0_outputs(6678)));
    outputs(1599) <= (layer0_outputs(6811)) and not (layer0_outputs(10060));
    outputs(1600) <= not(layer0_outputs(1395));
    outputs(1601) <= not(layer0_outputs(2131));
    outputs(1602) <= not(layer0_outputs(9030));
    outputs(1603) <= not((layer0_outputs(4757)) or (layer0_outputs(5391)));
    outputs(1604) <= layer0_outputs(6947);
    outputs(1605) <= not(layer0_outputs(8114));
    outputs(1606) <= (layer0_outputs(7108)) and (layer0_outputs(3014));
    outputs(1607) <= not(layer0_outputs(5194)) or (layer0_outputs(5841));
    outputs(1608) <= (layer0_outputs(5618)) and not (layer0_outputs(7350));
    outputs(1609) <= layer0_outputs(2654);
    outputs(1610) <= '0';
    outputs(1611) <= (layer0_outputs(6307)) and not (layer0_outputs(8257));
    outputs(1612) <= layer0_outputs(1248);
    outputs(1613) <= '0';
    outputs(1614) <= not((layer0_outputs(1961)) or (layer0_outputs(6966)));
    outputs(1615) <= not((layer0_outputs(6276)) or (layer0_outputs(3609)));
    outputs(1616) <= (layer0_outputs(5540)) and not (layer0_outputs(5109));
    outputs(1617) <= not(layer0_outputs(1962));
    outputs(1618) <= layer0_outputs(10041);
    outputs(1619) <= not((layer0_outputs(2186)) xor (layer0_outputs(698)));
    outputs(1620) <= not((layer0_outputs(6315)) xor (layer0_outputs(3599)));
    outputs(1621) <= not((layer0_outputs(9709)) xor (layer0_outputs(9897)));
    outputs(1622) <= (layer0_outputs(290)) and not (layer0_outputs(3656));
    outputs(1623) <= not(layer0_outputs(3613)) or (layer0_outputs(3347));
    outputs(1624) <= layer0_outputs(5045);
    outputs(1625) <= '0';
    outputs(1626) <= layer0_outputs(7377);
    outputs(1627) <= (layer0_outputs(972)) and (layer0_outputs(8166));
    outputs(1628) <= not(layer0_outputs(5812));
    outputs(1629) <= (layer0_outputs(9144)) and not (layer0_outputs(8646));
    outputs(1630) <= (layer0_outputs(6394)) and (layer0_outputs(4584));
    outputs(1631) <= not(layer0_outputs(5738));
    outputs(1632) <= '0';
    outputs(1633) <= not(layer0_outputs(1472)) or (layer0_outputs(8662));
    outputs(1634) <= not((layer0_outputs(3909)) or (layer0_outputs(7313)));
    outputs(1635) <= not((layer0_outputs(6046)) xor (layer0_outputs(4908)));
    outputs(1636) <= layer0_outputs(1747);
    outputs(1637) <= not(layer0_outputs(737));
    outputs(1638) <= not((layer0_outputs(4708)) xor (layer0_outputs(1346)));
    outputs(1639) <= (layer0_outputs(6807)) and not (layer0_outputs(6136));
    outputs(1640) <= (layer0_outputs(10009)) and (layer0_outputs(175));
    outputs(1641) <= (layer0_outputs(4738)) xor (layer0_outputs(9847));
    outputs(1642) <= layer0_outputs(30);
    outputs(1643) <= (layer0_outputs(4725)) and (layer0_outputs(4427));
    outputs(1644) <= not((layer0_outputs(1117)) or (layer0_outputs(7055)));
    outputs(1645) <= layer0_outputs(1651);
    outputs(1646) <= (layer0_outputs(8582)) and not (layer0_outputs(525));
    outputs(1647) <= layer0_outputs(5929);
    outputs(1648) <= (layer0_outputs(3761)) xor (layer0_outputs(788));
    outputs(1649) <= not(layer0_outputs(3202));
    outputs(1650) <= (layer0_outputs(10207)) and (layer0_outputs(393));
    outputs(1651) <= (layer0_outputs(9106)) xor (layer0_outputs(3807));
    outputs(1652) <= not((layer0_outputs(4534)) or (layer0_outputs(257)));
    outputs(1653) <= (layer0_outputs(7733)) and (layer0_outputs(4979));
    outputs(1654) <= (layer0_outputs(7522)) xor (layer0_outputs(6555));
    outputs(1655) <= (layer0_outputs(9326)) xor (layer0_outputs(1430));
    outputs(1656) <= not(layer0_outputs(556));
    outputs(1657) <= layer0_outputs(1923);
    outputs(1658) <= (layer0_outputs(120)) and (layer0_outputs(7341));
    outputs(1659) <= (layer0_outputs(7514)) and not (layer0_outputs(2350));
    outputs(1660) <= layer0_outputs(6608);
    outputs(1661) <= (layer0_outputs(1204)) xor (layer0_outputs(4965));
    outputs(1662) <= (layer0_outputs(2375)) xor (layer0_outputs(5253));
    outputs(1663) <= (layer0_outputs(6880)) and not (layer0_outputs(3715));
    outputs(1664) <= not((layer0_outputs(6587)) or (layer0_outputs(4161)));
    outputs(1665) <= layer0_outputs(16);
    outputs(1666) <= (layer0_outputs(7903)) and not (layer0_outputs(6670));
    outputs(1667) <= not((layer0_outputs(5335)) or (layer0_outputs(7646)));
    outputs(1668) <= not((layer0_outputs(2074)) xor (layer0_outputs(9099)));
    outputs(1669) <= not((layer0_outputs(6376)) or (layer0_outputs(10232)));
    outputs(1670) <= layer0_outputs(9570);
    outputs(1671) <= layer0_outputs(600);
    outputs(1672) <= '0';
    outputs(1673) <= (layer0_outputs(3455)) and (layer0_outputs(272));
    outputs(1674) <= (layer0_outputs(2567)) xor (layer0_outputs(4896));
    outputs(1675) <= (layer0_outputs(6190)) and not (layer0_outputs(3807));
    outputs(1676) <= not(layer0_outputs(712)) or (layer0_outputs(6714));
    outputs(1677) <= (layer0_outputs(8290)) and not (layer0_outputs(4655));
    outputs(1678) <= (layer0_outputs(5097)) xor (layer0_outputs(9112));
    outputs(1679) <= not(layer0_outputs(6508));
    outputs(1680) <= not(layer0_outputs(8540));
    outputs(1681) <= (layer0_outputs(1101)) and not (layer0_outputs(9776));
    outputs(1682) <= (layer0_outputs(2625)) and not (layer0_outputs(1538));
    outputs(1683) <= not(layer0_outputs(1966));
    outputs(1684) <= layer0_outputs(3274);
    outputs(1685) <= not((layer0_outputs(8272)) or (layer0_outputs(8654)));
    outputs(1686) <= (layer0_outputs(8220)) and not (layer0_outputs(185));
    outputs(1687) <= not((layer0_outputs(102)) or (layer0_outputs(9865)));
    outputs(1688) <= (layer0_outputs(7489)) and not (layer0_outputs(955));
    outputs(1689) <= (layer0_outputs(634)) xor (layer0_outputs(6414));
    outputs(1690) <= (layer0_outputs(7317)) and not (layer0_outputs(3572));
    outputs(1691) <= not((layer0_outputs(1797)) or (layer0_outputs(5206)));
    outputs(1692) <= (layer0_outputs(4647)) and not (layer0_outputs(3883));
    outputs(1693) <= not(layer0_outputs(5303));
    outputs(1694) <= (layer0_outputs(5446)) xor (layer0_outputs(6777));
    outputs(1695) <= not((layer0_outputs(8233)) xor (layer0_outputs(8799)));
    outputs(1696) <= layer0_outputs(9714);
    outputs(1697) <= not(layer0_outputs(2631));
    outputs(1698) <= (layer0_outputs(534)) and not (layer0_outputs(5813));
    outputs(1699) <= layer0_outputs(5587);
    outputs(1700) <= not(layer0_outputs(5228));
    outputs(1701) <= (layer0_outputs(8167)) xor (layer0_outputs(3806));
    outputs(1702) <= (layer0_outputs(8705)) xor (layer0_outputs(5672));
    outputs(1703) <= (layer0_outputs(3192)) and not (layer0_outputs(1329));
    outputs(1704) <= (layer0_outputs(6371)) and (layer0_outputs(9332));
    outputs(1705) <= (layer0_outputs(7157)) and not (layer0_outputs(7878));
    outputs(1706) <= (layer0_outputs(2383)) and not (layer0_outputs(3220));
    outputs(1707) <= not(layer0_outputs(4924));
    outputs(1708) <= layer0_outputs(2667);
    outputs(1709) <= not((layer0_outputs(3485)) xor (layer0_outputs(5735)));
    outputs(1710) <= (layer0_outputs(1879)) and not (layer0_outputs(1574));
    outputs(1711) <= not((layer0_outputs(7843)) or (layer0_outputs(3014)));
    outputs(1712) <= not(layer0_outputs(8681));
    outputs(1713) <= not((layer0_outputs(10191)) xor (layer0_outputs(4066)));
    outputs(1714) <= (layer0_outputs(9242)) xor (layer0_outputs(8450));
    outputs(1715) <= (layer0_outputs(2236)) and not (layer0_outputs(865));
    outputs(1716) <= (layer0_outputs(8647)) xor (layer0_outputs(7223));
    outputs(1717) <= not((layer0_outputs(1119)) xor (layer0_outputs(3779)));
    outputs(1718) <= (layer0_outputs(6477)) xor (layer0_outputs(9097));
    outputs(1719) <= (layer0_outputs(1578)) and (layer0_outputs(6293));
    outputs(1720) <= not((layer0_outputs(5140)) or (layer0_outputs(8204)));
    outputs(1721) <= not((layer0_outputs(1620)) and (layer0_outputs(6804)));
    outputs(1722) <= not(layer0_outputs(312));
    outputs(1723) <= (layer0_outputs(7688)) and (layer0_outputs(2558));
    outputs(1724) <= not((layer0_outputs(2891)) xor (layer0_outputs(5974)));
    outputs(1725) <= layer0_outputs(999);
    outputs(1726) <= (layer0_outputs(4434)) xor (layer0_outputs(232));
    outputs(1727) <= not((layer0_outputs(2199)) or (layer0_outputs(4912)));
    outputs(1728) <= (layer0_outputs(9525)) and (layer0_outputs(1919));
    outputs(1729) <= (layer0_outputs(995)) xor (layer0_outputs(10237));
    outputs(1730) <= not((layer0_outputs(5290)) xor (layer0_outputs(8025)));
    outputs(1731) <= (layer0_outputs(6102)) and (layer0_outputs(2291));
    outputs(1732) <= (layer0_outputs(9510)) and not (layer0_outputs(4952));
    outputs(1733) <= not(layer0_outputs(7724));
    outputs(1734) <= not(layer0_outputs(1074));
    outputs(1735) <= not((layer0_outputs(2421)) or (layer0_outputs(6406)));
    outputs(1736) <= (layer0_outputs(5274)) and not (layer0_outputs(6674));
    outputs(1737) <= not(layer0_outputs(6826));
    outputs(1738) <= not((layer0_outputs(5200)) or (layer0_outputs(4623)));
    outputs(1739) <= not((layer0_outputs(4174)) xor (layer0_outputs(10138)));
    outputs(1740) <= not((layer0_outputs(5578)) or (layer0_outputs(2582)));
    outputs(1741) <= (layer0_outputs(3000)) xor (layer0_outputs(2692));
    outputs(1742) <= layer0_outputs(9641);
    outputs(1743) <= (layer0_outputs(4727)) and (layer0_outputs(7641));
    outputs(1744) <= not((layer0_outputs(9755)) xor (layer0_outputs(478)));
    outputs(1745) <= (layer0_outputs(825)) and not (layer0_outputs(581));
    outputs(1746) <= layer0_outputs(6943);
    outputs(1747) <= layer0_outputs(7615);
    outputs(1748) <= layer0_outputs(8663);
    outputs(1749) <= (layer0_outputs(4152)) and not (layer0_outputs(8384));
    outputs(1750) <= not((layer0_outputs(8522)) xor (layer0_outputs(5132)));
    outputs(1751) <= not((layer0_outputs(2827)) xor (layer0_outputs(647)));
    outputs(1752) <= layer0_outputs(4059);
    outputs(1753) <= not((layer0_outputs(7766)) or (layer0_outputs(4772)));
    outputs(1754) <= not(layer0_outputs(1351));
    outputs(1755) <= not(layer0_outputs(2438));
    outputs(1756) <= layer0_outputs(4494);
    outputs(1757) <= (layer0_outputs(4008)) xor (layer0_outputs(293));
    outputs(1758) <= layer0_outputs(5306);
    outputs(1759) <= '0';
    outputs(1760) <= layer0_outputs(6296);
    outputs(1761) <= (layer0_outputs(9601)) and (layer0_outputs(8970));
    outputs(1762) <= (layer0_outputs(959)) or (layer0_outputs(6355));
    outputs(1763) <= (layer0_outputs(8579)) and not (layer0_outputs(7924));
    outputs(1764) <= layer0_outputs(2600);
    outputs(1765) <= (layer0_outputs(9711)) xor (layer0_outputs(9601));
    outputs(1766) <= (layer0_outputs(9225)) xor (layer0_outputs(8751));
    outputs(1767) <= (layer0_outputs(2909)) and not (layer0_outputs(6129));
    outputs(1768) <= not(layer0_outputs(9276));
    outputs(1769) <= (layer0_outputs(4257)) and not (layer0_outputs(3184));
    outputs(1770) <= not((layer0_outputs(4599)) or (layer0_outputs(9476)));
    outputs(1771) <= (layer0_outputs(9775)) and (layer0_outputs(2231));
    outputs(1772) <= not(layer0_outputs(5950));
    outputs(1773) <= layer0_outputs(7817);
    outputs(1774) <= (layer0_outputs(3857)) and not (layer0_outputs(1848));
    outputs(1775) <= (layer0_outputs(6259)) and not (layer0_outputs(359));
    outputs(1776) <= layer0_outputs(1);
    outputs(1777) <= (layer0_outputs(73)) and (layer0_outputs(5906));
    outputs(1778) <= not((layer0_outputs(8965)) xor (layer0_outputs(2209)));
    outputs(1779) <= layer0_outputs(9885);
    outputs(1780) <= not(layer0_outputs(3643));
    outputs(1781) <= (layer0_outputs(5591)) and (layer0_outputs(6008));
    outputs(1782) <= layer0_outputs(7096);
    outputs(1783) <= (layer0_outputs(4689)) xor (layer0_outputs(5464));
    outputs(1784) <= not(layer0_outputs(4093));
    outputs(1785) <= not((layer0_outputs(4974)) or (layer0_outputs(186)));
    outputs(1786) <= (layer0_outputs(4028)) and not (layer0_outputs(8437));
    outputs(1787) <= not(layer0_outputs(2574));
    outputs(1788) <= layer0_outputs(2869);
    outputs(1789) <= layer0_outputs(3410);
    outputs(1790) <= (layer0_outputs(2869)) xor (layer0_outputs(7740));
    outputs(1791) <= layer0_outputs(8584);
    outputs(1792) <= not(layer0_outputs(9682));
    outputs(1793) <= not(layer0_outputs(3746));
    outputs(1794) <= layer0_outputs(7714);
    outputs(1795) <= (layer0_outputs(3892)) and not (layer0_outputs(3299));
    outputs(1796) <= (layer0_outputs(4179)) and (layer0_outputs(7033));
    outputs(1797) <= '0';
    outputs(1798) <= (layer0_outputs(2207)) and not (layer0_outputs(6749));
    outputs(1799) <= layer0_outputs(5999);
    outputs(1800) <= (layer0_outputs(7097)) and not (layer0_outputs(1390));
    outputs(1801) <= (layer0_outputs(6605)) and not (layer0_outputs(6281));
    outputs(1802) <= (layer0_outputs(3788)) xor (layer0_outputs(5433));
    outputs(1803) <= (layer0_outputs(4486)) and not (layer0_outputs(5570));
    outputs(1804) <= (layer0_outputs(6073)) and not (layer0_outputs(442));
    outputs(1805) <= layer0_outputs(7983);
    outputs(1806) <= layer0_outputs(9716);
    outputs(1807) <= not((layer0_outputs(5891)) xor (layer0_outputs(8485)));
    outputs(1808) <= not((layer0_outputs(867)) xor (layer0_outputs(6978)));
    outputs(1809) <= (layer0_outputs(2214)) and (layer0_outputs(5259));
    outputs(1810) <= (layer0_outputs(9688)) and (layer0_outputs(10));
    outputs(1811) <= not(layer0_outputs(2248));
    outputs(1812) <= not((layer0_outputs(10175)) xor (layer0_outputs(9883)));
    outputs(1813) <= (layer0_outputs(9070)) xor (layer0_outputs(5007));
    outputs(1814) <= not(layer0_outputs(2053));
    outputs(1815) <= not((layer0_outputs(2041)) or (layer0_outputs(2669)));
    outputs(1816) <= layer0_outputs(4805);
    outputs(1817) <= layer0_outputs(9652);
    outputs(1818) <= not(layer0_outputs(2846));
    outputs(1819) <= not((layer0_outputs(3420)) or (layer0_outputs(1669)));
    outputs(1820) <= (layer0_outputs(1443)) xor (layer0_outputs(2771));
    outputs(1821) <= not(layer0_outputs(6894));
    outputs(1822) <= '0';
    outputs(1823) <= (layer0_outputs(8820)) and not (layer0_outputs(6440));
    outputs(1824) <= (layer0_outputs(2088)) and (layer0_outputs(8201));
    outputs(1825) <= not(layer0_outputs(10027));
    outputs(1826) <= not(layer0_outputs(1905)) or (layer0_outputs(324));
    outputs(1827) <= (layer0_outputs(282)) and (layer0_outputs(6375));
    outputs(1828) <= (layer0_outputs(3199)) xor (layer0_outputs(8180));
    outputs(1829) <= not(layer0_outputs(7487));
    outputs(1830) <= not(layer0_outputs(9256));
    outputs(1831) <= not((layer0_outputs(7677)) or (layer0_outputs(882)));
    outputs(1832) <= '0';
    outputs(1833) <= (layer0_outputs(5619)) and not (layer0_outputs(9625));
    outputs(1834) <= not((layer0_outputs(1828)) or (layer0_outputs(8235)));
    outputs(1835) <= not((layer0_outputs(7132)) or (layer0_outputs(5740)));
    outputs(1836) <= not((layer0_outputs(628)) xor (layer0_outputs(435)));
    outputs(1837) <= (layer0_outputs(4183)) and not (layer0_outputs(3272));
    outputs(1838) <= (layer0_outputs(5283)) and not (layer0_outputs(1474));
    outputs(1839) <= not((layer0_outputs(7419)) xor (layer0_outputs(8417)));
    outputs(1840) <= (layer0_outputs(8710)) xor (layer0_outputs(975));
    outputs(1841) <= not((layer0_outputs(5388)) or (layer0_outputs(1685)));
    outputs(1842) <= (layer0_outputs(517)) and (layer0_outputs(9183));
    outputs(1843) <= (layer0_outputs(1704)) and (layer0_outputs(8264));
    outputs(1844) <= not(layer0_outputs(1083));
    outputs(1845) <= not((layer0_outputs(3148)) or (layer0_outputs(5664)));
    outputs(1846) <= '0';
    outputs(1847) <= (layer0_outputs(744)) and not (layer0_outputs(9130));
    outputs(1848) <= layer0_outputs(3959);
    outputs(1849) <= (layer0_outputs(3297)) xor (layer0_outputs(1343));
    outputs(1850) <= not((layer0_outputs(5167)) xor (layer0_outputs(1270)));
    outputs(1851) <= not((layer0_outputs(6059)) xor (layer0_outputs(9140)));
    outputs(1852) <= layer0_outputs(5405);
    outputs(1853) <= not(layer0_outputs(56));
    outputs(1854) <= (layer0_outputs(7036)) and (layer0_outputs(2922));
    outputs(1855) <= not((layer0_outputs(8261)) or (layer0_outputs(8996)));
    outputs(1856) <= not(layer0_outputs(5407));
    outputs(1857) <= (layer0_outputs(7371)) and not (layer0_outputs(3168));
    outputs(1858) <= not((layer0_outputs(2851)) or (layer0_outputs(7936)));
    outputs(1859) <= layer0_outputs(6857);
    outputs(1860) <= (layer0_outputs(9274)) and (layer0_outputs(6223));
    outputs(1861) <= layer0_outputs(3444);
    outputs(1862) <= not((layer0_outputs(2639)) xor (layer0_outputs(4453)));
    outputs(1863) <= not((layer0_outputs(497)) or (layer0_outputs(6171)));
    outputs(1864) <= not(layer0_outputs(6334));
    outputs(1865) <= (layer0_outputs(1680)) and (layer0_outputs(4987));
    outputs(1866) <= layer0_outputs(112);
    outputs(1867) <= (layer0_outputs(2668)) xor (layer0_outputs(6264));
    outputs(1868) <= (layer0_outputs(8427)) and not (layer0_outputs(9151));
    outputs(1869) <= not(layer0_outputs(1140));
    outputs(1870) <= (layer0_outputs(2431)) and not (layer0_outputs(2142));
    outputs(1871) <= not(layer0_outputs(287));
    outputs(1872) <= not(layer0_outputs(4858));
    outputs(1873) <= not(layer0_outputs(6012));
    outputs(1874) <= (layer0_outputs(3066)) and not (layer0_outputs(3105));
    outputs(1875) <= not(layer0_outputs(7050));
    outputs(1876) <= (layer0_outputs(5794)) and (layer0_outputs(9750));
    outputs(1877) <= (layer0_outputs(7840)) and not (layer0_outputs(6879));
    outputs(1878) <= not((layer0_outputs(2857)) or (layer0_outputs(4819)));
    outputs(1879) <= (layer0_outputs(3579)) and not (layer0_outputs(5159));
    outputs(1880) <= not(layer0_outputs(4562));
    outputs(1881) <= not((layer0_outputs(8081)) or (layer0_outputs(9169)));
    outputs(1882) <= (layer0_outputs(8267)) and not (layer0_outputs(6613));
    outputs(1883) <= (layer0_outputs(1733)) and (layer0_outputs(6449));
    outputs(1884) <= not(layer0_outputs(7922));
    outputs(1885) <= not((layer0_outputs(9849)) xor (layer0_outputs(7471)));
    outputs(1886) <= (layer0_outputs(8013)) and not (layer0_outputs(4638));
    outputs(1887) <= not(layer0_outputs(2254));
    outputs(1888) <= layer0_outputs(387);
    outputs(1889) <= (layer0_outputs(2065)) and not (layer0_outputs(7427));
    outputs(1890) <= (layer0_outputs(6672)) and not (layer0_outputs(4146));
    outputs(1891) <= not(layer0_outputs(200));
    outputs(1892) <= (layer0_outputs(7088)) and not (layer0_outputs(4371));
    outputs(1893) <= not(layer0_outputs(6153));
    outputs(1894) <= layer0_outputs(6380);
    outputs(1895) <= not((layer0_outputs(187)) or (layer0_outputs(3)));
    outputs(1896) <= not((layer0_outputs(5899)) or (layer0_outputs(8807)));
    outputs(1897) <= not((layer0_outputs(8855)) or (layer0_outputs(6170)));
    outputs(1898) <= (layer0_outputs(44)) xor (layer0_outputs(1424));
    outputs(1899) <= not(layer0_outputs(8128));
    outputs(1900) <= layer0_outputs(8474);
    outputs(1901) <= (layer0_outputs(6693)) and not (layer0_outputs(3600));
    outputs(1902) <= (layer0_outputs(8303)) and not (layer0_outputs(8652));
    outputs(1903) <= (layer0_outputs(8568)) xor (layer0_outputs(6918));
    outputs(1904) <= (layer0_outputs(3823)) xor (layer0_outputs(6327));
    outputs(1905) <= not((layer0_outputs(9282)) or (layer0_outputs(10064)));
    outputs(1906) <= (layer0_outputs(3457)) and not (layer0_outputs(1975));
    outputs(1907) <= (layer0_outputs(10200)) xor (layer0_outputs(2797));
    outputs(1908) <= not((layer0_outputs(3210)) xor (layer0_outputs(3576)));
    outputs(1909) <= '0';
    outputs(1910) <= '0';
    outputs(1911) <= layer0_outputs(7275);
    outputs(1912) <= layer0_outputs(4403);
    outputs(1913) <= not((layer0_outputs(1557)) or (layer0_outputs(5268)));
    outputs(1914) <= (layer0_outputs(3821)) and (layer0_outputs(3601));
    outputs(1915) <= (layer0_outputs(9373)) and not (layer0_outputs(1857));
    outputs(1916) <= (layer0_outputs(3527)) and (layer0_outputs(3077));
    outputs(1917) <= not(layer0_outputs(6275));
    outputs(1918) <= not(layer0_outputs(3736));
    outputs(1919) <= (layer0_outputs(464)) and (layer0_outputs(7647));
    outputs(1920) <= not((layer0_outputs(2511)) xor (layer0_outputs(4282)));
    outputs(1921) <= (layer0_outputs(3729)) and not (layer0_outputs(1171));
    outputs(1922) <= (layer0_outputs(8361)) xor (layer0_outputs(2892));
    outputs(1923) <= not((layer0_outputs(6061)) xor (layer0_outputs(846)));
    outputs(1924) <= not(layer0_outputs(1386));
    outputs(1925) <= not(layer0_outputs(2585));
    outputs(1926) <= not((layer0_outputs(2860)) or (layer0_outputs(9330)));
    outputs(1927) <= not((layer0_outputs(729)) xor (layer0_outputs(4053)));
    outputs(1928) <= not((layer0_outputs(1532)) or (layer0_outputs(7087)));
    outputs(1929) <= not((layer0_outputs(3862)) xor (layer0_outputs(7934)));
    outputs(1930) <= (layer0_outputs(5009)) xor (layer0_outputs(3674));
    outputs(1931) <= (layer0_outputs(5353)) and (layer0_outputs(2425));
    outputs(1932) <= (layer0_outputs(7463)) xor (layer0_outputs(4547));
    outputs(1933) <= (layer0_outputs(1287)) xor (layer0_outputs(6718));
    outputs(1934) <= not(layer0_outputs(4305));
    outputs(1935) <= (layer0_outputs(4497)) xor (layer0_outputs(8510));
    outputs(1936) <= not((layer0_outputs(4519)) or (layer0_outputs(9896)));
    outputs(1937) <= (layer0_outputs(9870)) xor (layer0_outputs(2557));
    outputs(1938) <= (layer0_outputs(7955)) and (layer0_outputs(8648));
    outputs(1939) <= not(layer0_outputs(5539));
    outputs(1940) <= not(layer0_outputs(727));
    outputs(1941) <= (layer0_outputs(1406)) and not (layer0_outputs(83));
    outputs(1942) <= not(layer0_outputs(8838));
    outputs(1943) <= not(layer0_outputs(1115));
    outputs(1944) <= (layer0_outputs(915)) xor (layer0_outputs(7995));
    outputs(1945) <= (layer0_outputs(6950)) xor (layer0_outputs(8673));
    outputs(1946) <= not(layer0_outputs(3589));
    outputs(1947) <= layer0_outputs(3355);
    outputs(1948) <= not((layer0_outputs(3882)) or (layer0_outputs(7238)));
    outputs(1949) <= not((layer0_outputs(1637)) xor (layer0_outputs(4388)));
    outputs(1950) <= not((layer0_outputs(4334)) or (layer0_outputs(9552)));
    outputs(1951) <= (layer0_outputs(858)) xor (layer0_outputs(1272));
    outputs(1952) <= (layer0_outputs(6915)) and (layer0_outputs(5004));
    outputs(1953) <= not((layer0_outputs(1900)) or (layer0_outputs(2212)));
    outputs(1954) <= layer0_outputs(8434);
    outputs(1955) <= (layer0_outputs(3956)) and (layer0_outputs(4451));
    outputs(1956) <= not(layer0_outputs(6052));
    outputs(1957) <= not((layer0_outputs(2068)) or (layer0_outputs(6454)));
    outputs(1958) <= (layer0_outputs(7554)) and not (layer0_outputs(8620));
    outputs(1959) <= (layer0_outputs(1812)) xor (layer0_outputs(4840));
    outputs(1960) <= (layer0_outputs(2625)) and (layer0_outputs(2245));
    outputs(1961) <= layer0_outputs(5342);
    outputs(1962) <= not(layer0_outputs(4941));
    outputs(1963) <= layer0_outputs(3509);
    outputs(1964) <= not(layer0_outputs(1240));
    outputs(1965) <= (layer0_outputs(3958)) and not (layer0_outputs(390));
    outputs(1966) <= layer0_outputs(9444);
    outputs(1967) <= not((layer0_outputs(9115)) or (layer0_outputs(9311)));
    outputs(1968) <= (layer0_outputs(1457)) xor (layer0_outputs(7736));
    outputs(1969) <= not(layer0_outputs(4581));
    outputs(1970) <= '0';
    outputs(1971) <= (layer0_outputs(2047)) xor (layer0_outputs(1387));
    outputs(1972) <= (layer0_outputs(1303)) and not (layer0_outputs(8469));
    outputs(1973) <= layer0_outputs(4608);
    outputs(1974) <= not((layer0_outputs(712)) or (layer0_outputs(7962)));
    outputs(1975) <= not(layer0_outputs(4036));
    outputs(1976) <= not((layer0_outputs(4999)) or (layer0_outputs(10121)));
    outputs(1977) <= layer0_outputs(866);
    outputs(1978) <= layer0_outputs(3595);
    outputs(1979) <= not((layer0_outputs(2111)) or (layer0_outputs(98)));
    outputs(1980) <= layer0_outputs(1710);
    outputs(1981) <= (layer0_outputs(5142)) and (layer0_outputs(7777));
    outputs(1982) <= (layer0_outputs(2338)) and not (layer0_outputs(468));
    outputs(1983) <= not((layer0_outputs(2855)) xor (layer0_outputs(8066)));
    outputs(1984) <= not((layer0_outputs(4367)) or (layer0_outputs(707)));
    outputs(1985) <= not((layer0_outputs(4043)) or (layer0_outputs(10036)));
    outputs(1986) <= layer0_outputs(2699);
    outputs(1987) <= (layer0_outputs(3550)) and not (layer0_outputs(9205));
    outputs(1988) <= (layer0_outputs(1180)) and (layer0_outputs(2169));
    outputs(1989) <= (layer0_outputs(8708)) xor (layer0_outputs(1661));
    outputs(1990) <= (layer0_outputs(7744)) and not (layer0_outputs(8724));
    outputs(1991) <= not(layer0_outputs(8851));
    outputs(1992) <= (layer0_outputs(2586)) and not (layer0_outputs(3282));
    outputs(1993) <= (layer0_outputs(6301)) and not (layer0_outputs(8048));
    outputs(1994) <= layer0_outputs(6635);
    outputs(1995) <= not((layer0_outputs(6825)) or (layer0_outputs(4008)));
    outputs(1996) <= (layer0_outputs(7589)) and (layer0_outputs(9268));
    outputs(1997) <= (layer0_outputs(8315)) xor (layer0_outputs(878));
    outputs(1998) <= not(layer0_outputs(9049));
    outputs(1999) <= layer0_outputs(4392);
    outputs(2000) <= (layer0_outputs(9246)) and not (layer0_outputs(9776));
    outputs(2001) <= layer0_outputs(722);
    outputs(2002) <= (layer0_outputs(10152)) and not (layer0_outputs(572));
    outputs(2003) <= not((layer0_outputs(9816)) or (layer0_outputs(7173)));
    outputs(2004) <= layer0_outputs(6565);
    outputs(2005) <= (layer0_outputs(7743)) xor (layer0_outputs(4169));
    outputs(2006) <= not(layer0_outputs(8060));
    outputs(2007) <= layer0_outputs(6553);
    outputs(2008) <= not((layer0_outputs(733)) or (layer0_outputs(3022)));
    outputs(2009) <= (layer0_outputs(6336)) and not (layer0_outputs(2859));
    outputs(2010) <= not(layer0_outputs(8634));
    outputs(2011) <= not(layer0_outputs(3061));
    outputs(2012) <= not(layer0_outputs(1844));
    outputs(2013) <= layer0_outputs(5565);
    outputs(2014) <= layer0_outputs(318);
    outputs(2015) <= (layer0_outputs(9831)) and not (layer0_outputs(8081));
    outputs(2016) <= not((layer0_outputs(3021)) and (layer0_outputs(9292)));
    outputs(2017) <= not((layer0_outputs(3429)) or (layer0_outputs(2430)));
    outputs(2018) <= not((layer0_outputs(4064)) or (layer0_outputs(1863)));
    outputs(2019) <= not((layer0_outputs(1940)) xor (layer0_outputs(3845)));
    outputs(2020) <= not(layer0_outputs(7926));
    outputs(2021) <= not((layer0_outputs(4204)) xor (layer0_outputs(9864)));
    outputs(2022) <= not(layer0_outputs(7995));
    outputs(2023) <= not((layer0_outputs(4018)) or (layer0_outputs(5293)));
    outputs(2024) <= not(layer0_outputs(3984));
    outputs(2025) <= not((layer0_outputs(7634)) xor (layer0_outputs(8739)));
    outputs(2026) <= not((layer0_outputs(10204)) or (layer0_outputs(2387)));
    outputs(2027) <= (layer0_outputs(8887)) and not (layer0_outputs(4809));
    outputs(2028) <= not(layer0_outputs(5534));
    outputs(2029) <= not(layer0_outputs(8697));
    outputs(2030) <= (layer0_outputs(4613)) and (layer0_outputs(4502));
    outputs(2031) <= (layer0_outputs(6443)) and not (layer0_outputs(7607));
    outputs(2032) <= layer0_outputs(4266);
    outputs(2033) <= (layer0_outputs(9437)) and not (layer0_outputs(10014));
    outputs(2034) <= (layer0_outputs(1353)) and not (layer0_outputs(1010));
    outputs(2035) <= (layer0_outputs(7955)) and not (layer0_outputs(4411));
    outputs(2036) <= (layer0_outputs(5938)) and not (layer0_outputs(4747));
    outputs(2037) <= not(layer0_outputs(9210));
    outputs(2038) <= not(layer0_outputs(5684));
    outputs(2039) <= layer0_outputs(10237);
    outputs(2040) <= not(layer0_outputs(5360));
    outputs(2041) <= not((layer0_outputs(6298)) xor (layer0_outputs(5943)));
    outputs(2042) <= not((layer0_outputs(5637)) or (layer0_outputs(1808)));
    outputs(2043) <= layer0_outputs(9204);
    outputs(2044) <= not((layer0_outputs(761)) xor (layer0_outputs(9311)));
    outputs(2045) <= not((layer0_outputs(1734)) or (layer0_outputs(4818)));
    outputs(2046) <= not(layer0_outputs(2514));
    outputs(2047) <= (layer0_outputs(1699)) and not (layer0_outputs(536));
    outputs(2048) <= not((layer0_outputs(5835)) and (layer0_outputs(9251)));
    outputs(2049) <= not(layer0_outputs(1786)) or (layer0_outputs(3087));
    outputs(2050) <= not((layer0_outputs(9680)) xor (layer0_outputs(1479)));
    outputs(2051) <= (layer0_outputs(8494)) xor (layer0_outputs(3123));
    outputs(2052) <= layer0_outputs(8419);
    outputs(2053) <= not(layer0_outputs(6979)) or (layer0_outputs(9908));
    outputs(2054) <= not(layer0_outputs(4528));
    outputs(2055) <= not(layer0_outputs(872));
    outputs(2056) <= layer0_outputs(3902);
    outputs(2057) <= (layer0_outputs(3311)) or (layer0_outputs(2363));
    outputs(2058) <= layer0_outputs(9184);
    outputs(2059) <= not(layer0_outputs(3132)) or (layer0_outputs(1357));
    outputs(2060) <= (layer0_outputs(3574)) xor (layer0_outputs(7579));
    outputs(2061) <= not((layer0_outputs(6391)) or (layer0_outputs(7657)));
    outputs(2062) <= not(layer0_outputs(5049));
    outputs(2063) <= not((layer0_outputs(8316)) and (layer0_outputs(2774)));
    outputs(2064) <= (layer0_outputs(1627)) xor (layer0_outputs(4874));
    outputs(2065) <= not(layer0_outputs(4398));
    outputs(2066) <= (layer0_outputs(8262)) or (layer0_outputs(2614));
    outputs(2067) <= layer0_outputs(1889);
    outputs(2068) <= not(layer0_outputs(4993));
    outputs(2069) <= '1';
    outputs(2070) <= (layer0_outputs(6157)) xor (layer0_outputs(6353));
    outputs(2071) <= not(layer0_outputs(8478));
    outputs(2072) <= layer0_outputs(8751);
    outputs(2073) <= not(layer0_outputs(7734));
    outputs(2074) <= not((layer0_outputs(4517)) xor (layer0_outputs(455)));
    outputs(2075) <= not(layer0_outputs(9678));
    outputs(2076) <= not(layer0_outputs(10148));
    outputs(2077) <= (layer0_outputs(3559)) xor (layer0_outputs(7728));
    outputs(2078) <= not(layer0_outputs(9020));
    outputs(2079) <= not(layer0_outputs(5189)) or (layer0_outputs(7596));
    outputs(2080) <= layer0_outputs(5760);
    outputs(2081) <= (layer0_outputs(6815)) or (layer0_outputs(979));
    outputs(2082) <= layer0_outputs(7761);
    outputs(2083) <= not(layer0_outputs(4358)) or (layer0_outputs(6316));
    outputs(2084) <= not(layer0_outputs(2526));
    outputs(2085) <= not(layer0_outputs(240));
    outputs(2086) <= not((layer0_outputs(8954)) and (layer0_outputs(10231)));
    outputs(2087) <= layer0_outputs(9995);
    outputs(2088) <= not((layer0_outputs(8704)) xor (layer0_outputs(9661)));
    outputs(2089) <= layer0_outputs(9728);
    outputs(2090) <= layer0_outputs(4753);
    outputs(2091) <= not(layer0_outputs(7671));
    outputs(2092) <= not(layer0_outputs(1885));
    outputs(2093) <= not(layer0_outputs(6951));
    outputs(2094) <= not(layer0_outputs(8844)) or (layer0_outputs(549));
    outputs(2095) <= not((layer0_outputs(8674)) and (layer0_outputs(6665)));
    outputs(2096) <= not(layer0_outputs(3385)) or (layer0_outputs(3730));
    outputs(2097) <= (layer0_outputs(7165)) xor (layer0_outputs(5640));
    outputs(2098) <= layer0_outputs(9502);
    outputs(2099) <= not(layer0_outputs(7692));
    outputs(2100) <= layer0_outputs(1478);
    outputs(2101) <= (layer0_outputs(6087)) or (layer0_outputs(3144));
    outputs(2102) <= (layer0_outputs(6385)) xor (layer0_outputs(9977));
    outputs(2103) <= not((layer0_outputs(3318)) and (layer0_outputs(3135)));
    outputs(2104) <= (layer0_outputs(1490)) and not (layer0_outputs(9834));
    outputs(2105) <= layer0_outputs(1575);
    outputs(2106) <= layer0_outputs(4091);
    outputs(2107) <= not(layer0_outputs(3090));
    outputs(2108) <= not(layer0_outputs(782));
    outputs(2109) <= (layer0_outputs(1341)) xor (layer0_outputs(2905));
    outputs(2110) <= not(layer0_outputs(6608));
    outputs(2111) <= (layer0_outputs(2630)) or (layer0_outputs(8344));
    outputs(2112) <= not(layer0_outputs(2060)) or (layer0_outputs(9582));
    outputs(2113) <= not((layer0_outputs(2782)) xor (layer0_outputs(7765)));
    outputs(2114) <= not(layer0_outputs(4685));
    outputs(2115) <= not((layer0_outputs(6771)) and (layer0_outputs(2843)));
    outputs(2116) <= not(layer0_outputs(2779)) or (layer0_outputs(897));
    outputs(2117) <= (layer0_outputs(2726)) or (layer0_outputs(6785));
    outputs(2118) <= layer0_outputs(6713);
    outputs(2119) <= not(layer0_outputs(4331)) or (layer0_outputs(778));
    outputs(2120) <= layer0_outputs(5179);
    outputs(2121) <= layer0_outputs(9767);
    outputs(2122) <= layer0_outputs(534);
    outputs(2123) <= layer0_outputs(7410);
    outputs(2124) <= not((layer0_outputs(7409)) and (layer0_outputs(7269)));
    outputs(2125) <= (layer0_outputs(5577)) and (layer0_outputs(8331));
    outputs(2126) <= not(layer0_outputs(2605)) or (layer0_outputs(1927));
    outputs(2127) <= not(layer0_outputs(9033)) or (layer0_outputs(1133));
    outputs(2128) <= not(layer0_outputs(5464)) or (layer0_outputs(5488));
    outputs(2129) <= not((layer0_outputs(2153)) or (layer0_outputs(2929)));
    outputs(2130) <= layer0_outputs(913);
    outputs(2131) <= not(layer0_outputs(8811));
    outputs(2132) <= not(layer0_outputs(5314));
    outputs(2133) <= not(layer0_outputs(2716)) or (layer0_outputs(601));
    outputs(2134) <= (layer0_outputs(6114)) xor (layer0_outputs(2546));
    outputs(2135) <= not(layer0_outputs(3913));
    outputs(2136) <= not(layer0_outputs(8630)) or (layer0_outputs(775));
    outputs(2137) <= not(layer0_outputs(5551));
    outputs(2138) <= layer0_outputs(4608);
    outputs(2139) <= not((layer0_outputs(1060)) or (layer0_outputs(7866)));
    outputs(2140) <= not(layer0_outputs(6411)) or (layer0_outputs(5556));
    outputs(2141) <= not(layer0_outputs(2257)) or (layer0_outputs(5912));
    outputs(2142) <= not(layer0_outputs(984)) or (layer0_outputs(3400));
    outputs(2143) <= not((layer0_outputs(4030)) and (layer0_outputs(4815)));
    outputs(2144) <= layer0_outputs(2199);
    outputs(2145) <= layer0_outputs(7918);
    outputs(2146) <= not(layer0_outputs(4948)) or (layer0_outputs(9589));
    outputs(2147) <= not(layer0_outputs(3627));
    outputs(2148) <= (layer0_outputs(8520)) or (layer0_outputs(6070));
    outputs(2149) <= not(layer0_outputs(2774));
    outputs(2150) <= (layer0_outputs(6410)) or (layer0_outputs(8885));
    outputs(2151) <= layer0_outputs(4715);
    outputs(2152) <= layer0_outputs(1559);
    outputs(2153) <= (layer0_outputs(1342)) or (layer0_outputs(6021));
    outputs(2154) <= not(layer0_outputs(1667)) or (layer0_outputs(1300));
    outputs(2155) <= layer0_outputs(9441);
    outputs(2156) <= not(layer0_outputs(5489));
    outputs(2157) <= not(layer0_outputs(4096));
    outputs(2158) <= layer0_outputs(1437);
    outputs(2159) <= not((layer0_outputs(9014)) and (layer0_outputs(3801)));
    outputs(2160) <= not((layer0_outputs(6713)) and (layer0_outputs(3201)));
    outputs(2161) <= (layer0_outputs(8902)) and (layer0_outputs(6350));
    outputs(2162) <= layer0_outputs(653);
    outputs(2163) <= (layer0_outputs(3018)) xor (layer0_outputs(7298));
    outputs(2164) <= (layer0_outputs(3217)) xor (layer0_outputs(8580));
    outputs(2165) <= (layer0_outputs(2840)) and (layer0_outputs(9421));
    outputs(2166) <= layer0_outputs(73);
    outputs(2167) <= (layer0_outputs(2636)) and not (layer0_outputs(526));
    outputs(2168) <= layer0_outputs(8732);
    outputs(2169) <= not(layer0_outputs(8945));
    outputs(2170) <= not(layer0_outputs(6192));
    outputs(2171) <= not((layer0_outputs(3776)) and (layer0_outputs(5884)));
    outputs(2172) <= not(layer0_outputs(622)) or (layer0_outputs(6841));
    outputs(2173) <= not(layer0_outputs(5080));
    outputs(2174) <= (layer0_outputs(10140)) xor (layer0_outputs(3150));
    outputs(2175) <= layer0_outputs(2198);
    outputs(2176) <= not(layer0_outputs(1600)) or (layer0_outputs(140));
    outputs(2177) <= not(layer0_outputs(5347));
    outputs(2178) <= (layer0_outputs(2304)) xor (layer0_outputs(8065));
    outputs(2179) <= not(layer0_outputs(11));
    outputs(2180) <= not(layer0_outputs(566)) or (layer0_outputs(5740));
    outputs(2181) <= (layer0_outputs(5743)) or (layer0_outputs(8183));
    outputs(2182) <= layer0_outputs(1810);
    outputs(2183) <= (layer0_outputs(5187)) and (layer0_outputs(4230));
    outputs(2184) <= not(layer0_outputs(2076));
    outputs(2185) <= layer0_outputs(2838);
    outputs(2186) <= not(layer0_outputs(7679));
    outputs(2187) <= not(layer0_outputs(4887)) or (layer0_outputs(6790));
    outputs(2188) <= (layer0_outputs(145)) xor (layer0_outputs(3481));
    outputs(2189) <= (layer0_outputs(3577)) or (layer0_outputs(9438));
    outputs(2190) <= layer0_outputs(3591);
    outputs(2191) <= layer0_outputs(1573);
    outputs(2192) <= not(layer0_outputs(2684));
    outputs(2193) <= not(layer0_outputs(8332)) or (layer0_outputs(9600));
    outputs(2194) <= not(layer0_outputs(2439)) or (layer0_outputs(5488));
    outputs(2195) <= layer0_outputs(8147);
    outputs(2196) <= layer0_outputs(8909);
    outputs(2197) <= not(layer0_outputs(2145)) or (layer0_outputs(1515));
    outputs(2198) <= not(layer0_outputs(10198));
    outputs(2199) <= layer0_outputs(4119);
    outputs(2200) <= (layer0_outputs(512)) xor (layer0_outputs(1183));
    outputs(2201) <= not(layer0_outputs(4003));
    outputs(2202) <= layer0_outputs(3199);
    outputs(2203) <= layer0_outputs(7084);
    outputs(2204) <= layer0_outputs(3493);
    outputs(2205) <= not((layer0_outputs(8490)) xor (layer0_outputs(7491)));
    outputs(2206) <= not((layer0_outputs(7050)) xor (layer0_outputs(2341)));
    outputs(2207) <= not(layer0_outputs(5624));
    outputs(2208) <= layer0_outputs(5625);
    outputs(2209) <= not(layer0_outputs(477)) or (layer0_outputs(9059));
    outputs(2210) <= (layer0_outputs(9574)) and not (layer0_outputs(5899));
    outputs(2211) <= not((layer0_outputs(3383)) and (layer0_outputs(5803)));
    outputs(2212) <= not(layer0_outputs(5654));
    outputs(2213) <= not(layer0_outputs(6067)) or (layer0_outputs(2646));
    outputs(2214) <= not(layer0_outputs(2362));
    outputs(2215) <= layer0_outputs(4576);
    outputs(2216) <= (layer0_outputs(6964)) xor (layer0_outputs(10047));
    outputs(2217) <= not(layer0_outputs(5097));
    outputs(2218) <= not((layer0_outputs(3709)) xor (layer0_outputs(7977)));
    outputs(2219) <= (layer0_outputs(3069)) xor (layer0_outputs(1337));
    outputs(2220) <= (layer0_outputs(8591)) and (layer0_outputs(7159));
    outputs(2221) <= (layer0_outputs(8473)) or (layer0_outputs(8320));
    outputs(2222) <= not(layer0_outputs(3253));
    outputs(2223) <= (layer0_outputs(2825)) and (layer0_outputs(2241));
    outputs(2224) <= layer0_outputs(4471);
    outputs(2225) <= not((layer0_outputs(1453)) xor (layer0_outputs(79)));
    outputs(2226) <= not((layer0_outputs(4633)) xor (layer0_outputs(4925)));
    outputs(2227) <= not((layer0_outputs(3215)) xor (layer0_outputs(6972)));
    outputs(2228) <= not((layer0_outputs(5707)) or (layer0_outputs(3424)));
    outputs(2229) <= layer0_outputs(9804);
    outputs(2230) <= not(layer0_outputs(3456));
    outputs(2231) <= layer0_outputs(8351);
    outputs(2232) <= not(layer0_outputs(3100));
    outputs(2233) <= not((layer0_outputs(6384)) or (layer0_outputs(868)));
    outputs(2234) <= not((layer0_outputs(3082)) and (layer0_outputs(7860)));
    outputs(2235) <= (layer0_outputs(7320)) or (layer0_outputs(3263));
    outputs(2236) <= layer0_outputs(3339);
    outputs(2237) <= not(layer0_outputs(925));
    outputs(2238) <= not((layer0_outputs(26)) or (layer0_outputs(1751)));
    outputs(2239) <= not(layer0_outputs(3342));
    outputs(2240) <= not(layer0_outputs(4884));
    outputs(2241) <= layer0_outputs(3174);
    outputs(2242) <= layer0_outputs(6902);
    outputs(2243) <= not((layer0_outputs(7166)) or (layer0_outputs(3585)));
    outputs(2244) <= not(layer0_outputs(7067));
    outputs(2245) <= not(layer0_outputs(6724));
    outputs(2246) <= not((layer0_outputs(9236)) xor (layer0_outputs(9358)));
    outputs(2247) <= (layer0_outputs(1555)) or (layer0_outputs(3449));
    outputs(2248) <= (layer0_outputs(4081)) xor (layer0_outputs(4318));
    outputs(2249) <= not(layer0_outputs(9308));
    outputs(2250) <= not((layer0_outputs(4076)) or (layer0_outputs(10084)));
    outputs(2251) <= (layer0_outputs(7100)) xor (layer0_outputs(5182));
    outputs(2252) <= layer0_outputs(2124);
    outputs(2253) <= (layer0_outputs(7250)) xor (layer0_outputs(2858));
    outputs(2254) <= not((layer0_outputs(9190)) xor (layer0_outputs(5120)));
    outputs(2255) <= layer0_outputs(9925);
    outputs(2256) <= not(layer0_outputs(1013));
    outputs(2257) <= not(layer0_outputs(7296));
    outputs(2258) <= not((layer0_outputs(1632)) xor (layer0_outputs(1215)));
    outputs(2259) <= not(layer0_outputs(2806));
    outputs(2260) <= (layer0_outputs(1056)) or (layer0_outputs(994));
    outputs(2261) <= (layer0_outputs(6209)) xor (layer0_outputs(4833));
    outputs(2262) <= (layer0_outputs(4557)) and (layer0_outputs(4289));
    outputs(2263) <= layer0_outputs(7297);
    outputs(2264) <= (layer0_outputs(9250)) and not (layer0_outputs(10062));
    outputs(2265) <= not((layer0_outputs(5724)) or (layer0_outputs(101)));
    outputs(2266) <= layer0_outputs(6200);
    outputs(2267) <= layer0_outputs(6175);
    outputs(2268) <= layer0_outputs(3934);
    outputs(2269) <= (layer0_outputs(4222)) xor (layer0_outputs(6721));
    outputs(2270) <= (layer0_outputs(9296)) xor (layer0_outputs(1782));
    outputs(2271) <= not(layer0_outputs(5031));
    outputs(2272) <= (layer0_outputs(7174)) and (layer0_outputs(6003));
    outputs(2273) <= layer0_outputs(2096);
    outputs(2274) <= not(layer0_outputs(4819));
    outputs(2275) <= not(layer0_outputs(3091));
    outputs(2276) <= not((layer0_outputs(4956)) xor (layer0_outputs(7715)));
    outputs(2277) <= not((layer0_outputs(5246)) or (layer0_outputs(10089)));
    outputs(2278) <= not(layer0_outputs(367)) or (layer0_outputs(795));
    outputs(2279) <= (layer0_outputs(4291)) xor (layer0_outputs(9264));
    outputs(2280) <= not(layer0_outputs(2033)) or (layer0_outputs(626));
    outputs(2281) <= not(layer0_outputs(9340));
    outputs(2282) <= not(layer0_outputs(5205));
    outputs(2283) <= not(layer0_outputs(308));
    outputs(2284) <= not(layer0_outputs(2855)) or (layer0_outputs(7767));
    outputs(2285) <= (layer0_outputs(4980)) xor (layer0_outputs(4173));
    outputs(2286) <= not(layer0_outputs(10167));
    outputs(2287) <= layer0_outputs(7561);
    outputs(2288) <= not(layer0_outputs(6613));
    outputs(2289) <= layer0_outputs(3809);
    outputs(2290) <= layer0_outputs(1509);
    outputs(2291) <= (layer0_outputs(3483)) or (layer0_outputs(6780));
    outputs(2292) <= layer0_outputs(4134);
    outputs(2293) <= (layer0_outputs(6824)) and (layer0_outputs(3711));
    outputs(2294) <= not(layer0_outputs(364));
    outputs(2295) <= not((layer0_outputs(4145)) and (layer0_outputs(1345)));
    outputs(2296) <= (layer0_outputs(6702)) xor (layer0_outputs(9896));
    outputs(2297) <= (layer0_outputs(1623)) or (layer0_outputs(9962));
    outputs(2298) <= not((layer0_outputs(6875)) xor (layer0_outputs(8376)));
    outputs(2299) <= layer0_outputs(8237);
    outputs(2300) <= not(layer0_outputs(1763));
    outputs(2301) <= not((layer0_outputs(8832)) xor (layer0_outputs(934)));
    outputs(2302) <= not(layer0_outputs(1151)) or (layer0_outputs(779));
    outputs(2303) <= (layer0_outputs(302)) and not (layer0_outputs(2970));
    outputs(2304) <= layer0_outputs(7509);
    outputs(2305) <= (layer0_outputs(1990)) xor (layer0_outputs(650));
    outputs(2306) <= (layer0_outputs(5381)) or (layer0_outputs(8542));
    outputs(2307) <= not(layer0_outputs(7828));
    outputs(2308) <= (layer0_outputs(8856)) xor (layer0_outputs(9159));
    outputs(2309) <= not(layer0_outputs(5354));
    outputs(2310) <= layer0_outputs(9612);
    outputs(2311) <= not(layer0_outputs(2229));
    outputs(2312) <= layer0_outputs(7043);
    outputs(2313) <= (layer0_outputs(2355)) and (layer0_outputs(133));
    outputs(2314) <= layer0_outputs(2895);
    outputs(2315) <= (layer0_outputs(298)) or (layer0_outputs(4933));
    outputs(2316) <= not(layer0_outputs(2621)) or (layer0_outputs(151));
    outputs(2317) <= layer0_outputs(9417);
    outputs(2318) <= (layer0_outputs(3505)) xor (layer0_outputs(7862));
    outputs(2319) <= (layer0_outputs(9297)) xor (layer0_outputs(6952));
    outputs(2320) <= (layer0_outputs(6487)) and (layer0_outputs(4257));
    outputs(2321) <= not(layer0_outputs(214));
    outputs(2322) <= (layer0_outputs(2494)) xor (layer0_outputs(6438));
    outputs(2323) <= not((layer0_outputs(2415)) and (layer0_outputs(5536)));
    outputs(2324) <= (layer0_outputs(1142)) xor (layer0_outputs(3365));
    outputs(2325) <= not(layer0_outputs(5534));
    outputs(2326) <= not((layer0_outputs(3229)) or (layer0_outputs(1542)));
    outputs(2327) <= not(layer0_outputs(1836)) or (layer0_outputs(8419));
    outputs(2328) <= not(layer0_outputs(2970));
    outputs(2329) <= not(layer0_outputs(3467));
    outputs(2330) <= (layer0_outputs(6322)) xor (layer0_outputs(2022));
    outputs(2331) <= (layer0_outputs(3867)) and not (layer0_outputs(4877));
    outputs(2332) <= not(layer0_outputs(7804));
    outputs(2333) <= not(layer0_outputs(3322));
    outputs(2334) <= not(layer0_outputs(6468));
    outputs(2335) <= (layer0_outputs(220)) and not (layer0_outputs(5553));
    outputs(2336) <= not(layer0_outputs(3560)) or (layer0_outputs(2799));
    outputs(2337) <= not(layer0_outputs(9989));
    outputs(2338) <= layer0_outputs(8655);
    outputs(2339) <= (layer0_outputs(7059)) or (layer0_outputs(1887));
    outputs(2340) <= not((layer0_outputs(7786)) and (layer0_outputs(4232)));
    outputs(2341) <= not(layer0_outputs(5666));
    outputs(2342) <= layer0_outputs(9113);
    outputs(2343) <= not(layer0_outputs(8247));
    outputs(2344) <= not(layer0_outputs(7813));
    outputs(2345) <= not(layer0_outputs(9766));
    outputs(2346) <= not((layer0_outputs(9117)) or (layer0_outputs(3844)));
    outputs(2347) <= (layer0_outputs(2437)) xor (layer0_outputs(9346));
    outputs(2348) <= not((layer0_outputs(8988)) xor (layer0_outputs(3722)));
    outputs(2349) <= (layer0_outputs(5364)) and not (layer0_outputs(3469));
    outputs(2350) <= (layer0_outputs(8312)) and (layer0_outputs(3152));
    outputs(2351) <= not(layer0_outputs(7567));
    outputs(2352) <= not(layer0_outputs(7649)) or (layer0_outputs(6949));
    outputs(2353) <= (layer0_outputs(4521)) or (layer0_outputs(4682));
    outputs(2354) <= not(layer0_outputs(8313)) or (layer0_outputs(4837));
    outputs(2355) <= (layer0_outputs(241)) xor (layer0_outputs(2044));
    outputs(2356) <= (layer0_outputs(4074)) xor (layer0_outputs(4726));
    outputs(2357) <= not(layer0_outputs(5831));
    outputs(2358) <= layer0_outputs(3692);
    outputs(2359) <= layer0_outputs(8087);
    outputs(2360) <= layer0_outputs(8614);
    outputs(2361) <= not((layer0_outputs(2866)) and (layer0_outputs(5041)));
    outputs(2362) <= not((layer0_outputs(7733)) and (layer0_outputs(4758)));
    outputs(2363) <= (layer0_outputs(5746)) and not (layer0_outputs(8313));
    outputs(2364) <= layer0_outputs(7047);
    outputs(2365) <= not(layer0_outputs(3395)) or (layer0_outputs(2943));
    outputs(2366) <= not(layer0_outputs(10008)) or (layer0_outputs(2537));
    outputs(2367) <= not((layer0_outputs(7710)) xor (layer0_outputs(95)));
    outputs(2368) <= not(layer0_outputs(5508));
    outputs(2369) <= (layer0_outputs(9567)) and (layer0_outputs(9026));
    outputs(2370) <= layer0_outputs(5058);
    outputs(2371) <= (layer0_outputs(3587)) or (layer0_outputs(27));
    outputs(2372) <= (layer0_outputs(1623)) xor (layer0_outputs(1179));
    outputs(2373) <= not(layer0_outputs(2346));
    outputs(2374) <= not((layer0_outputs(8027)) xor (layer0_outputs(3781)));
    outputs(2375) <= not(layer0_outputs(9496));
    outputs(2376) <= not(layer0_outputs(3043)) or (layer0_outputs(297));
    outputs(2377) <= not(layer0_outputs(5751));
    outputs(2378) <= (layer0_outputs(2677)) and not (layer0_outputs(6443));
    outputs(2379) <= not(layer0_outputs(5147));
    outputs(2380) <= (layer0_outputs(767)) xor (layer0_outputs(2753));
    outputs(2381) <= not(layer0_outputs(6459));
    outputs(2382) <= not(layer0_outputs(8766));
    outputs(2383) <= not(layer0_outputs(2982));
    outputs(2384) <= layer0_outputs(537);
    outputs(2385) <= not(layer0_outputs(3954));
    outputs(2386) <= (layer0_outputs(1969)) and (layer0_outputs(3895));
    outputs(2387) <= not((layer0_outputs(938)) or (layer0_outputs(8086)));
    outputs(2388) <= not(layer0_outputs(1346));
    outputs(2389) <= not(layer0_outputs(2700));
    outputs(2390) <= layer0_outputs(35);
    outputs(2391) <= not((layer0_outputs(2734)) or (layer0_outputs(4720)));
    outputs(2392) <= not(layer0_outputs(2632)) or (layer0_outputs(2686));
    outputs(2393) <= not((layer0_outputs(5493)) xor (layer0_outputs(6338)));
    outputs(2394) <= (layer0_outputs(514)) and not (layer0_outputs(5135));
    outputs(2395) <= not(layer0_outputs(8951));
    outputs(2396) <= not(layer0_outputs(873)) or (layer0_outputs(8784));
    outputs(2397) <= layer0_outputs(1626);
    outputs(2398) <= (layer0_outputs(4428)) xor (layer0_outputs(4413));
    outputs(2399) <= not(layer0_outputs(2777));
    outputs(2400) <= not(layer0_outputs(5511));
    outputs(2401) <= not(layer0_outputs(5365));
    outputs(2402) <= not((layer0_outputs(500)) xor (layer0_outputs(1153)));
    outputs(2403) <= (layer0_outputs(4304)) xor (layer0_outputs(3357));
    outputs(2404) <= not((layer0_outputs(4144)) xor (layer0_outputs(3854)));
    outputs(2405) <= not((layer0_outputs(3580)) and (layer0_outputs(146)));
    outputs(2406) <= (layer0_outputs(7593)) and not (layer0_outputs(3138));
    outputs(2407) <= not((layer0_outputs(1047)) and (layer0_outputs(3716)));
    outputs(2408) <= not((layer0_outputs(9083)) and (layer0_outputs(7265)));
    outputs(2409) <= not(layer0_outputs(7075)) or (layer0_outputs(5288));
    outputs(2410) <= layer0_outputs(76);
    outputs(2411) <= not(layer0_outputs(10145));
    outputs(2412) <= layer0_outputs(756);
    outputs(2413) <= not(layer0_outputs(5383)) or (layer0_outputs(9789));
    outputs(2414) <= not(layer0_outputs(4262)) or (layer0_outputs(4153));
    outputs(2415) <= (layer0_outputs(5787)) and not (layer0_outputs(3490));
    outputs(2416) <= not((layer0_outputs(9569)) and (layer0_outputs(7967)));
    outputs(2417) <= (layer0_outputs(5993)) xor (layer0_outputs(10219));
    outputs(2418) <= layer0_outputs(3309);
    outputs(2419) <= (layer0_outputs(10025)) and (layer0_outputs(7190));
    outputs(2420) <= layer0_outputs(8872);
    outputs(2421) <= not((layer0_outputs(4187)) and (layer0_outputs(2658)));
    outputs(2422) <= not(layer0_outputs(6676));
    outputs(2423) <= not(layer0_outputs(3932)) or (layer0_outputs(9095));
    outputs(2424) <= (layer0_outputs(2073)) and (layer0_outputs(9637));
    outputs(2425) <= not(layer0_outputs(8285));
    outputs(2426) <= not(layer0_outputs(4369));
    outputs(2427) <= layer0_outputs(8643);
    outputs(2428) <= not((layer0_outputs(6891)) xor (layer0_outputs(1442)));
    outputs(2429) <= layer0_outputs(6250);
    outputs(2430) <= not(layer0_outputs(7525));
    outputs(2431) <= not((layer0_outputs(1222)) and (layer0_outputs(1521)));
    outputs(2432) <= layer0_outputs(1946);
    outputs(2433) <= not(layer0_outputs(924));
    outputs(2434) <= not(layer0_outputs(2711)) or (layer0_outputs(2980));
    outputs(2435) <= (layer0_outputs(1754)) xor (layer0_outputs(1069));
    outputs(2436) <= (layer0_outputs(10220)) or (layer0_outputs(8429));
    outputs(2437) <= not((layer0_outputs(198)) and (layer0_outputs(8043)));
    outputs(2438) <= (layer0_outputs(431)) xor (layer0_outputs(6662));
    outputs(2439) <= (layer0_outputs(1638)) or (layer0_outputs(8164));
    outputs(2440) <= layer0_outputs(6727);
    outputs(2441) <= not(layer0_outputs(5484)) or (layer0_outputs(9355));
    outputs(2442) <= not((layer0_outputs(2398)) or (layer0_outputs(2719)));
    outputs(2443) <= not(layer0_outputs(5046));
    outputs(2444) <= not(layer0_outputs(5986));
    outputs(2445) <= (layer0_outputs(6844)) or (layer0_outputs(5456));
    outputs(2446) <= not(layer0_outputs(625));
    outputs(2447) <= (layer0_outputs(2459)) xor (layer0_outputs(5660));
    outputs(2448) <= layer0_outputs(1223);
    outputs(2449) <= (layer0_outputs(8892)) and not (layer0_outputs(10011));
    outputs(2450) <= layer0_outputs(9527);
    outputs(2451) <= layer0_outputs(9814);
    outputs(2452) <= layer0_outputs(2533);
    outputs(2453) <= layer0_outputs(8697);
    outputs(2454) <= not(layer0_outputs(7004)) or (layer0_outputs(8704));
    outputs(2455) <= not(layer0_outputs(7735)) or (layer0_outputs(2676));
    outputs(2456) <= (layer0_outputs(6719)) and not (layer0_outputs(420));
    outputs(2457) <= not((layer0_outputs(5690)) and (layer0_outputs(2049)));
    outputs(2458) <= not(layer0_outputs(3848));
    outputs(2459) <= (layer0_outputs(7716)) and (layer0_outputs(5457));
    outputs(2460) <= layer0_outputs(2013);
    outputs(2461) <= not((layer0_outputs(2764)) xor (layer0_outputs(7963)));
    outputs(2462) <= not(layer0_outputs(10072));
    outputs(2463) <= layer0_outputs(6203);
    outputs(2464) <= (layer0_outputs(47)) or (layer0_outputs(7498));
    outputs(2465) <= layer0_outputs(3678);
    outputs(2466) <= layer0_outputs(4330);
    outputs(2467) <= layer0_outputs(401);
    outputs(2468) <= not((layer0_outputs(7126)) or (layer0_outputs(5051)));
    outputs(2469) <= not(layer0_outputs(4609)) or (layer0_outputs(257));
    outputs(2470) <= not(layer0_outputs(7455)) or (layer0_outputs(1691));
    outputs(2471) <= not((layer0_outputs(8067)) xor (layer0_outputs(7940)));
    outputs(2472) <= not(layer0_outputs(102));
    outputs(2473) <= (layer0_outputs(7486)) and not (layer0_outputs(1116));
    outputs(2474) <= layer0_outputs(4785);
    outputs(2475) <= not(layer0_outputs(3421)) or (layer0_outputs(5143));
    outputs(2476) <= layer0_outputs(3586);
    outputs(2477) <= (layer0_outputs(4075)) or (layer0_outputs(2860));
    outputs(2478) <= not((layer0_outputs(7750)) and (layer0_outputs(7871)));
    outputs(2479) <= not(layer0_outputs(9666)) or (layer0_outputs(2934));
    outputs(2480) <= layer0_outputs(4715);
    outputs(2481) <= (layer0_outputs(9868)) xor (layer0_outputs(7006));
    outputs(2482) <= (layer0_outputs(6196)) or (layer0_outputs(8288));
    outputs(2483) <= not(layer0_outputs(9384)) or (layer0_outputs(980));
    outputs(2484) <= (layer0_outputs(2762)) and not (layer0_outputs(499));
    outputs(2485) <= layer0_outputs(4562);
    outputs(2486) <= (layer0_outputs(6386)) and not (layer0_outputs(7219));
    outputs(2487) <= layer0_outputs(5239);
    outputs(2488) <= not((layer0_outputs(1739)) or (layer0_outputs(6031)));
    outputs(2489) <= layer0_outputs(10169);
    outputs(2490) <= not((layer0_outputs(9489)) xor (layer0_outputs(3701)));
    outputs(2491) <= not((layer0_outputs(745)) and (layer0_outputs(6256)));
    outputs(2492) <= (layer0_outputs(4195)) xor (layer0_outputs(2395));
    outputs(2493) <= not(layer0_outputs(2917));
    outputs(2494) <= layer0_outputs(7184);
    outputs(2495) <= (layer0_outputs(3269)) and not (layer0_outputs(2456));
    outputs(2496) <= layer0_outputs(7432);
    outputs(2497) <= layer0_outputs(4597);
    outputs(2498) <= layer0_outputs(2666);
    outputs(2499) <= not((layer0_outputs(3546)) xor (layer0_outputs(8144)));
    outputs(2500) <= not(layer0_outputs(4129));
    outputs(2501) <= layer0_outputs(7256);
    outputs(2502) <= not((layer0_outputs(3010)) xor (layer0_outputs(8200)));
    outputs(2503) <= layer0_outputs(877);
    outputs(2504) <= not(layer0_outputs(3526));
    outputs(2505) <= not((layer0_outputs(9822)) xor (layer0_outputs(871)));
    outputs(2506) <= layer0_outputs(5616);
    outputs(2507) <= (layer0_outputs(10173)) and not (layer0_outputs(4426));
    outputs(2508) <= (layer0_outputs(3443)) xor (layer0_outputs(9912));
    outputs(2509) <= (layer0_outputs(4215)) xor (layer0_outputs(8006));
    outputs(2510) <= not(layer0_outputs(1326)) or (layer0_outputs(4319));
    outputs(2511) <= (layer0_outputs(1417)) or (layer0_outputs(5354));
    outputs(2512) <= not(layer0_outputs(2400)) or (layer0_outputs(8462));
    outputs(2513) <= not(layer0_outputs(168));
    outputs(2514) <= not(layer0_outputs(6649)) or (layer0_outputs(9484));
    outputs(2515) <= not((layer0_outputs(5682)) or (layer0_outputs(1846)));
    outputs(2516) <= not(layer0_outputs(6118));
    outputs(2517) <= (layer0_outputs(6137)) or (layer0_outputs(6989));
    outputs(2518) <= (layer0_outputs(485)) xor (layer0_outputs(7713));
    outputs(2519) <= not(layer0_outputs(665)) or (layer0_outputs(8556));
    outputs(2520) <= (layer0_outputs(823)) or (layer0_outputs(5010));
    outputs(2521) <= not((layer0_outputs(1227)) and (layer0_outputs(1505)));
    outputs(2522) <= not(layer0_outputs(1847)) or (layer0_outputs(9906));
    outputs(2523) <= (layer0_outputs(2877)) xor (layer0_outputs(9665));
    outputs(2524) <= (layer0_outputs(7302)) and not (layer0_outputs(5333));
    outputs(2525) <= not((layer0_outputs(692)) xor (layer0_outputs(5907)));
    outputs(2526) <= layer0_outputs(9987);
    outputs(2527) <= not(layer0_outputs(7416));
    outputs(2528) <= layer0_outputs(9987);
    outputs(2529) <= (layer0_outputs(5521)) or (layer0_outputs(8959));
    outputs(2530) <= (layer0_outputs(10150)) or (layer0_outputs(2953));
    outputs(2531) <= not(layer0_outputs(7312)) or (layer0_outputs(2353));
    outputs(2532) <= layer0_outputs(9710);
    outputs(2533) <= not((layer0_outputs(5007)) or (layer0_outputs(10180)));
    outputs(2534) <= (layer0_outputs(9092)) and not (layer0_outputs(1203));
    outputs(2535) <= (layer0_outputs(1455)) xor (layer0_outputs(372));
    outputs(2536) <= not((layer0_outputs(9131)) and (layer0_outputs(8605)));
    outputs(2537) <= not((layer0_outputs(7868)) or (layer0_outputs(8370)));
    outputs(2538) <= not(layer0_outputs(10104));
    outputs(2539) <= not(layer0_outputs(2033));
    outputs(2540) <= layer0_outputs(1136);
    outputs(2541) <= not(layer0_outputs(3333)) or (layer0_outputs(3632));
    outputs(2542) <= not((layer0_outputs(8995)) xor (layer0_outputs(9685)));
    outputs(2543) <= not(layer0_outputs(3252));
    outputs(2544) <= not((layer0_outputs(1307)) xor (layer0_outputs(7200)));
    outputs(2545) <= not(layer0_outputs(2524));
    outputs(2546) <= not((layer0_outputs(1299)) xor (layer0_outputs(4123)));
    outputs(2547) <= not((layer0_outputs(6400)) and (layer0_outputs(8124)));
    outputs(2548) <= layer0_outputs(3732);
    outputs(2549) <= not(layer0_outputs(5031));
    outputs(2550) <= layer0_outputs(988);
    outputs(2551) <= not(layer0_outputs(5486));
    outputs(2552) <= not(layer0_outputs(3639));
    outputs(2553) <= not((layer0_outputs(1029)) xor (layer0_outputs(4268)));
    outputs(2554) <= not(layer0_outputs(4090));
    outputs(2555) <= not((layer0_outputs(5085)) or (layer0_outputs(2146)));
    outputs(2556) <= layer0_outputs(6253);
    outputs(2557) <= not(layer0_outputs(7060)) or (layer0_outputs(8761));
    outputs(2558) <= not(layer0_outputs(5439));
    outputs(2559) <= (layer0_outputs(9029)) and not (layer0_outputs(4975));
    outputs(2560) <= not((layer0_outputs(5229)) and (layer0_outputs(6717)));
    outputs(2561) <= (layer0_outputs(153)) or (layer0_outputs(7305));
    outputs(2562) <= not(layer0_outputs(1042));
    outputs(2563) <= not(layer0_outputs(2378));
    outputs(2564) <= not((layer0_outputs(5052)) xor (layer0_outputs(825)));
    outputs(2565) <= not((layer0_outputs(3765)) xor (layer0_outputs(7222)));
    outputs(2566) <= not((layer0_outputs(3232)) and (layer0_outputs(7906)));
    outputs(2567) <= not((layer0_outputs(1344)) xor (layer0_outputs(7601)));
    outputs(2568) <= not((layer0_outputs(8228)) xor (layer0_outputs(7548)));
    outputs(2569) <= not(layer0_outputs(1266));
    outputs(2570) <= not((layer0_outputs(3468)) and (layer0_outputs(6502)));
    outputs(2571) <= not((layer0_outputs(2580)) xor (layer0_outputs(8365)));
    outputs(2572) <= not((layer0_outputs(4171)) xor (layer0_outputs(1820)));
    outputs(2573) <= not(layer0_outputs(318));
    outputs(2574) <= (layer0_outputs(1178)) or (layer0_outputs(8218));
    outputs(2575) <= layer0_outputs(4002);
    outputs(2576) <= (layer0_outputs(7249)) or (layer0_outputs(1748));
    outputs(2577) <= not((layer0_outputs(615)) or (layer0_outputs(2440)));
    outputs(2578) <= (layer0_outputs(5185)) xor (layer0_outputs(2702));
    outputs(2579) <= not(layer0_outputs(3998));
    outputs(2580) <= not(layer0_outputs(3233)) or (layer0_outputs(4848));
    outputs(2581) <= not((layer0_outputs(8250)) xor (layer0_outputs(6235)));
    outputs(2582) <= layer0_outputs(6338);
    outputs(2583) <= layer0_outputs(8535);
    outputs(2584) <= not(layer0_outputs(9795)) or (layer0_outputs(1712));
    outputs(2585) <= not(layer0_outputs(9663));
    outputs(2586) <= not((layer0_outputs(138)) xor (layer0_outputs(2194)));
    outputs(2587) <= (layer0_outputs(2593)) and not (layer0_outputs(1709));
    outputs(2588) <= not((layer0_outputs(8549)) and (layer0_outputs(1612)));
    outputs(2589) <= layer0_outputs(1636);
    outputs(2590) <= (layer0_outputs(3531)) xor (layer0_outputs(9815));
    outputs(2591) <= (layer0_outputs(518)) and (layer0_outputs(384));
    outputs(2592) <= layer0_outputs(1578);
    outputs(2593) <= (layer0_outputs(7503)) or (layer0_outputs(4748));
    outputs(2594) <= not(layer0_outputs(5645));
    outputs(2595) <= not(layer0_outputs(7218));
    outputs(2596) <= (layer0_outputs(939)) and not (layer0_outputs(462));
    outputs(2597) <= (layer0_outputs(1341)) xor (layer0_outputs(8146));
    outputs(2598) <= (layer0_outputs(1017)) xor (layer0_outputs(1675));
    outputs(2599) <= (layer0_outputs(8040)) and not (layer0_outputs(5763));
    outputs(2600) <= (layer0_outputs(8308)) and not (layer0_outputs(3467));
    outputs(2601) <= layer0_outputs(6473);
    outputs(2602) <= not(layer0_outputs(6017)) or (layer0_outputs(6615));
    outputs(2603) <= '1';
    outputs(2604) <= not((layer0_outputs(6197)) xor (layer0_outputs(880)));
    outputs(2605) <= not(layer0_outputs(3373));
    outputs(2606) <= not(layer0_outputs(1672));
    outputs(2607) <= not(layer0_outputs(7395));
    outputs(2608) <= (layer0_outputs(2983)) and not (layer0_outputs(7706));
    outputs(2609) <= not(layer0_outputs(8515)) or (layer0_outputs(8318));
    outputs(2610) <= (layer0_outputs(4766)) xor (layer0_outputs(7635));
    outputs(2611) <= not(layer0_outputs(9768)) or (layer0_outputs(1425));
    outputs(2612) <= not((layer0_outputs(6333)) xor (layer0_outputs(10127)));
    outputs(2613) <= not((layer0_outputs(3268)) and (layer0_outputs(8841)));
    outputs(2614) <= not(layer0_outputs(7119)) or (layer0_outputs(4201));
    outputs(2615) <= layer0_outputs(2599);
    outputs(2616) <= not(layer0_outputs(9431)) or (layer0_outputs(1179));
    outputs(2617) <= not((layer0_outputs(4355)) or (layer0_outputs(2141)));
    outputs(2618) <= layer0_outputs(4119);
    outputs(2619) <= (layer0_outputs(3251)) and not (layer0_outputs(9281));
    outputs(2620) <= (layer0_outputs(3976)) or (layer0_outputs(563));
    outputs(2621) <= not((layer0_outputs(5176)) or (layer0_outputs(6591)));
    outputs(2622) <= not((layer0_outputs(4492)) xor (layer0_outputs(3879)));
    outputs(2623) <= not(layer0_outputs(10186));
    outputs(2624) <= not(layer0_outputs(3597)) or (layer0_outputs(5094));
    outputs(2625) <= not((layer0_outputs(4654)) and (layer0_outputs(7875)));
    outputs(2626) <= layer0_outputs(3368);
    outputs(2627) <= layer0_outputs(4123);
    outputs(2628) <= not(layer0_outputs(2058));
    outputs(2629) <= layer0_outputs(5451);
    outputs(2630) <= not((layer0_outputs(1693)) or (layer0_outputs(5892)));
    outputs(2631) <= (layer0_outputs(2143)) and (layer0_outputs(844));
    outputs(2632) <= not(layer0_outputs(6905)) or (layer0_outputs(3874));
    outputs(2633) <= not(layer0_outputs(1302)) or (layer0_outputs(6082));
    outputs(2634) <= not(layer0_outputs(1763));
    outputs(2635) <= layer0_outputs(9546);
    outputs(2636) <= layer0_outputs(7761);
    outputs(2637) <= layer0_outputs(1824);
    outputs(2638) <= layer0_outputs(3972);
    outputs(2639) <= layer0_outputs(2021);
    outputs(2640) <= (layer0_outputs(8104)) xor (layer0_outputs(8984));
    outputs(2641) <= not((layer0_outputs(1767)) xor (layer0_outputs(9044)));
    outputs(2642) <= not((layer0_outputs(1566)) xor (layer0_outputs(9379)));
    outputs(2643) <= not((layer0_outputs(2721)) and (layer0_outputs(5461)));
    outputs(2644) <= not(layer0_outputs(1174)) or (layer0_outputs(2517));
    outputs(2645) <= (layer0_outputs(2244)) or (layer0_outputs(4394));
    outputs(2646) <= layer0_outputs(4604);
    outputs(2647) <= not(layer0_outputs(8472));
    outputs(2648) <= (layer0_outputs(8411)) or (layer0_outputs(1864));
    outputs(2649) <= layer0_outputs(700);
    outputs(2650) <= layer0_outputs(9354);
    outputs(2651) <= layer0_outputs(1781);
    outputs(2652) <= not(layer0_outputs(6549));
    outputs(2653) <= layer0_outputs(7531);
    outputs(2654) <= (layer0_outputs(609)) or (layer0_outputs(8507));
    outputs(2655) <= not(layer0_outputs(433));
    outputs(2656) <= (layer0_outputs(9441)) or (layer0_outputs(7687));
    outputs(2657) <= not(layer0_outputs(5654)) or (layer0_outputs(2931));
    outputs(2658) <= not(layer0_outputs(5307));
    outputs(2659) <= not(layer0_outputs(7307));
    outputs(2660) <= (layer0_outputs(6244)) or (layer0_outputs(7135));
    outputs(2661) <= (layer0_outputs(1774)) xor (layer0_outputs(8800));
    outputs(2662) <= (layer0_outputs(3213)) or (layer0_outputs(7188));
    outputs(2663) <= (layer0_outputs(3877)) and not (layer0_outputs(5285));
    outputs(2664) <= layer0_outputs(7509);
    outputs(2665) <= not(layer0_outputs(427)) or (layer0_outputs(2423));
    outputs(2666) <= (layer0_outputs(9903)) or (layer0_outputs(5958));
    outputs(2667) <= (layer0_outputs(2745)) xor (layer0_outputs(1064));
    outputs(2668) <= (layer0_outputs(8143)) and (layer0_outputs(1608));
    outputs(2669) <= layer0_outputs(4378);
    outputs(2670) <= not(layer0_outputs(7417)) or (layer0_outputs(2109));
    outputs(2671) <= not(layer0_outputs(3016));
    outputs(2672) <= (layer0_outputs(9128)) or (layer0_outputs(5698));
    outputs(2673) <= not(layer0_outputs(6883));
    outputs(2674) <= not(layer0_outputs(3790));
    outputs(2675) <= not(layer0_outputs(8394)) or (layer0_outputs(10016));
    outputs(2676) <= layer0_outputs(8476);
    outputs(2677) <= not((layer0_outputs(7605)) xor (layer0_outputs(7044)));
    outputs(2678) <= not(layer0_outputs(4452)) or (layer0_outputs(1979));
    outputs(2679) <= (layer0_outputs(5208)) or (layer0_outputs(8051));
    outputs(2680) <= layer0_outputs(2188);
    outputs(2681) <= not(layer0_outputs(9746));
    outputs(2682) <= (layer0_outputs(9689)) or (layer0_outputs(5300));
    outputs(2683) <= not(layer0_outputs(3491));
    outputs(2684) <= (layer0_outputs(6925)) xor (layer0_outputs(5220));
    outputs(2685) <= layer0_outputs(9214);
    outputs(2686) <= (layer0_outputs(3062)) and not (layer0_outputs(4349));
    outputs(2687) <= not(layer0_outputs(5548));
    outputs(2688) <= not(layer0_outputs(9195));
    outputs(2689) <= (layer0_outputs(1992)) and (layer0_outputs(867));
    outputs(2690) <= not((layer0_outputs(4135)) xor (layer0_outputs(3802)));
    outputs(2691) <= layer0_outputs(5095);
    outputs(2692) <= not(layer0_outputs(206));
    outputs(2693) <= layer0_outputs(1295);
    outputs(2694) <= not(layer0_outputs(6016)) or (layer0_outputs(4011));
    outputs(2695) <= not(layer0_outputs(1269)) or (layer0_outputs(6536));
    outputs(2696) <= not(layer0_outputs(2584));
    outputs(2697) <= not((layer0_outputs(5224)) xor (layer0_outputs(2651)));
    outputs(2698) <= not(layer0_outputs(8971));
    outputs(2699) <= not((layer0_outputs(6095)) xor (layer0_outputs(4208)));
    outputs(2700) <= not(layer0_outputs(1320));
    outputs(2701) <= not(layer0_outputs(2504)) or (layer0_outputs(7809));
    outputs(2702) <= not((layer0_outputs(7820)) and (layer0_outputs(8171)));
    outputs(2703) <= not((layer0_outputs(7301)) or (layer0_outputs(10193)));
    outputs(2704) <= not(layer0_outputs(4962)) or (layer0_outputs(7336));
    outputs(2705) <= not(layer0_outputs(8255));
    outputs(2706) <= not((layer0_outputs(2196)) or (layer0_outputs(2394)));
    outputs(2707) <= layer0_outputs(4465);
    outputs(2708) <= layer0_outputs(6090);
    outputs(2709) <= not(layer0_outputs(1360));
    outputs(2710) <= not(layer0_outputs(7053));
    outputs(2711) <= layer0_outputs(9836);
    outputs(2712) <= not(layer0_outputs(8852)) or (layer0_outputs(4539));
    outputs(2713) <= not(layer0_outputs(6393));
    outputs(2714) <= not(layer0_outputs(786));
    outputs(2715) <= (layer0_outputs(2437)) and not (layer0_outputs(3203));
    outputs(2716) <= layer0_outputs(2933);
    outputs(2717) <= layer0_outputs(1636);
    outputs(2718) <= layer0_outputs(6001);
    outputs(2719) <= not(layer0_outputs(9859)) or (layer0_outputs(2510));
    outputs(2720) <= layer0_outputs(7929);
    outputs(2721) <= not(layer0_outputs(1793));
    outputs(2722) <= layer0_outputs(610);
    outputs(2723) <= (layer0_outputs(1236)) or (layer0_outputs(1787));
    outputs(2724) <= layer0_outputs(4938);
    outputs(2725) <= (layer0_outputs(8277)) or (layer0_outputs(5839));
    outputs(2726) <= not((layer0_outputs(1759)) xor (layer0_outputs(2976)));
    outputs(2727) <= not(layer0_outputs(2872));
    outputs(2728) <= (layer0_outputs(6944)) xor (layer0_outputs(1370));
    outputs(2729) <= layer0_outputs(1202);
    outputs(2730) <= layer0_outputs(8050);
    outputs(2731) <= (layer0_outputs(6954)) and not (layer0_outputs(5858));
    outputs(2732) <= (layer0_outputs(8681)) and not (layer0_outputs(2322));
    outputs(2733) <= not((layer0_outputs(6453)) and (layer0_outputs(8882)));
    outputs(2734) <= (layer0_outputs(1075)) and (layer0_outputs(6093));
    outputs(2735) <= (layer0_outputs(2476)) xor (layer0_outputs(1482));
    outputs(2736) <= not((layer0_outputs(3747)) and (layer0_outputs(4685)));
    outputs(2737) <= not(layer0_outputs(3515)) or (layer0_outputs(3787));
    outputs(2738) <= not(layer0_outputs(9882));
    outputs(2739) <= (layer0_outputs(6111)) and not (layer0_outputs(5898));
    outputs(2740) <= not((layer0_outputs(1950)) xor (layer0_outputs(474)));
    outputs(2741) <= not(layer0_outputs(9160));
    outputs(2742) <= not(layer0_outputs(3177));
    outputs(2743) <= layer0_outputs(7381);
    outputs(2744) <= (layer0_outputs(8917)) xor (layer0_outputs(2642));
    outputs(2745) <= not(layer0_outputs(2161));
    outputs(2746) <= not((layer0_outputs(8840)) or (layer0_outputs(1479)));
    outputs(2747) <= (layer0_outputs(9923)) and (layer0_outputs(4865));
    outputs(2748) <= not(layer0_outputs(6325));
    outputs(2749) <= not((layer0_outputs(3596)) and (layer0_outputs(9168)));
    outputs(2750) <= (layer0_outputs(2427)) xor (layer0_outputs(8314));
    outputs(2751) <= (layer0_outputs(4329)) xor (layer0_outputs(505));
    outputs(2752) <= layer0_outputs(4506);
    outputs(2753) <= not(layer0_outputs(5832));
    outputs(2754) <= layer0_outputs(10172);
    outputs(2755) <= not(layer0_outputs(103));
    outputs(2756) <= not(layer0_outputs(4240));
    outputs(2757) <= not(layer0_outputs(3335));
    outputs(2758) <= not((layer0_outputs(4725)) and (layer0_outputs(1519)));
    outputs(2759) <= layer0_outputs(4632);
    outputs(2760) <= layer0_outputs(6727);
    outputs(2761) <= '1';
    outputs(2762) <= (layer0_outputs(9099)) xor (layer0_outputs(7365));
    outputs(2763) <= (layer0_outputs(7996)) or (layer0_outputs(5991));
    outputs(2764) <= not((layer0_outputs(2062)) xor (layer0_outputs(8641)));
    outputs(2765) <= (layer0_outputs(9539)) xor (layer0_outputs(5754));
    outputs(2766) <= not(layer0_outputs(3512));
    outputs(2767) <= not(layer0_outputs(5751));
    outputs(2768) <= layer0_outputs(878);
    outputs(2769) <= not((layer0_outputs(9978)) and (layer0_outputs(1664)));
    outputs(2770) <= not((layer0_outputs(3804)) and (layer0_outputs(7524)));
    outputs(2771) <= not(layer0_outputs(643));
    outputs(2772) <= not((layer0_outputs(973)) or (layer0_outputs(6836)));
    outputs(2773) <= (layer0_outputs(3660)) and (layer0_outputs(2757));
    outputs(2774) <= not(layer0_outputs(4762)) or (layer0_outputs(6796));
    outputs(2775) <= not(layer0_outputs(1775)) or (layer0_outputs(7305));
    outputs(2776) <= not((layer0_outputs(5409)) xor (layer0_outputs(3189)));
    outputs(2777) <= (layer0_outputs(1158)) xor (layer0_outputs(9668));
    outputs(2778) <= not(layer0_outputs(82)) or (layer0_outputs(2328));
    outputs(2779) <= not(layer0_outputs(7013));
    outputs(2780) <= layer0_outputs(6039);
    outputs(2781) <= (layer0_outputs(8153)) xor (layer0_outputs(5516));
    outputs(2782) <= not(layer0_outputs(10163)) or (layer0_outputs(4587));
    outputs(2783) <= not(layer0_outputs(4815));
    outputs(2784) <= not(layer0_outputs(8003));
    outputs(2785) <= layer0_outputs(5240);
    outputs(2786) <= not((layer0_outputs(9382)) xor (layer0_outputs(5086)));
    outputs(2787) <= not((layer0_outputs(7144)) xor (layer0_outputs(6163)));
    outputs(2788) <= (layer0_outputs(7505)) or (layer0_outputs(1676));
    outputs(2789) <= (layer0_outputs(2530)) xor (layer0_outputs(8544));
    outputs(2790) <= not(layer0_outputs(4831));
    outputs(2791) <= layer0_outputs(379);
    outputs(2792) <= not(layer0_outputs(4561));
    outputs(2793) <= not(layer0_outputs(4098)) or (layer0_outputs(5490));
    outputs(2794) <= (layer0_outputs(8851)) xor (layer0_outputs(3475));
    outputs(2795) <= not(layer0_outputs(343)) or (layer0_outputs(2056));
    outputs(2796) <= layer0_outputs(9911);
    outputs(2797) <= not((layer0_outputs(5024)) and (layer0_outputs(8438)));
    outputs(2798) <= layer0_outputs(2988);
    outputs(2799) <= not(layer0_outputs(10161));
    outputs(2800) <= layer0_outputs(8466);
    outputs(2801) <= not(layer0_outputs(3225));
    outputs(2802) <= not(layer0_outputs(5006));
    outputs(2803) <= not((layer0_outputs(9048)) xor (layer0_outputs(8795)));
    outputs(2804) <= not(layer0_outputs(3922)) or (layer0_outputs(4185));
    outputs(2805) <= not(layer0_outputs(7057));
    outputs(2806) <= not((layer0_outputs(8162)) or (layer0_outputs(3349)));
    outputs(2807) <= not((layer0_outputs(10072)) or (layer0_outputs(6889)));
    outputs(2808) <= (layer0_outputs(7380)) xor (layer0_outputs(4295));
    outputs(2809) <= not(layer0_outputs(10198));
    outputs(2810) <= not(layer0_outputs(9345));
    outputs(2811) <= (layer0_outputs(1492)) or (layer0_outputs(8163));
    outputs(2812) <= layer0_outputs(8614);
    outputs(2813) <= not(layer0_outputs(8604));
    outputs(2814) <= not(layer0_outputs(5502));
    outputs(2815) <= (layer0_outputs(6664)) xor (layer0_outputs(1562));
    outputs(2816) <= (layer0_outputs(7889)) and not (layer0_outputs(5066));
    outputs(2817) <= not((layer0_outputs(7864)) and (layer0_outputs(2900)));
    outputs(2818) <= not((layer0_outputs(1785)) xor (layer0_outputs(9544)));
    outputs(2819) <= layer0_outputs(6174);
    outputs(2820) <= not((layer0_outputs(2064)) xor (layer0_outputs(7217)));
    outputs(2821) <= not(layer0_outputs(5514));
    outputs(2822) <= (layer0_outputs(586)) and not (layer0_outputs(5851));
    outputs(2823) <= layer0_outputs(5520);
    outputs(2824) <= not(layer0_outputs(227));
    outputs(2825) <= not((layer0_outputs(343)) and (layer0_outputs(5301)));
    outputs(2826) <= not(layer0_outputs(6332)) or (layer0_outputs(5338));
    outputs(2827) <= not(layer0_outputs(3962));
    outputs(2828) <= layer0_outputs(9971);
    outputs(2829) <= not((layer0_outputs(4875)) xor (layer0_outputs(278)));
    outputs(2830) <= not(layer0_outputs(7132));
    outputs(2831) <= not((layer0_outputs(553)) and (layer0_outputs(4026)));
    outputs(2832) <= (layer0_outputs(1034)) xor (layer0_outputs(1361));
    outputs(2833) <= not(layer0_outputs(1094)) or (layer0_outputs(212));
    outputs(2834) <= (layer0_outputs(9372)) xor (layer0_outputs(6626));
    outputs(2835) <= (layer0_outputs(672)) xor (layer0_outputs(7745));
    outputs(2836) <= not((layer0_outputs(5448)) xor (layer0_outputs(9415)));
    outputs(2837) <= (layer0_outputs(7618)) and not (layer0_outputs(5360));
    outputs(2838) <= layer0_outputs(9325);
    outputs(2839) <= not(layer0_outputs(9891)) or (layer0_outputs(7942));
    outputs(2840) <= not(layer0_outputs(2131));
    outputs(2841) <= (layer0_outputs(624)) and (layer0_outputs(572));
    outputs(2842) <= (layer0_outputs(4634)) and not (layer0_outputs(362));
    outputs(2843) <= (layer0_outputs(8288)) or (layer0_outputs(5267));
    outputs(2844) <= (layer0_outputs(8112)) xor (layer0_outputs(1719));
    outputs(2845) <= not(layer0_outputs(5074));
    outputs(2846) <= (layer0_outputs(9269)) and (layer0_outputs(8864));
    outputs(2847) <= not(layer0_outputs(6880));
    outputs(2848) <= not(layer0_outputs(6000)) or (layer0_outputs(742));
    outputs(2849) <= (layer0_outputs(5303)) and not (layer0_outputs(4544));
    outputs(2850) <= not(layer0_outputs(5806));
    outputs(2851) <= not((layer0_outputs(7483)) xor (layer0_outputs(5699)));
    outputs(2852) <= (layer0_outputs(2247)) xor (layer0_outputs(7292));
    outputs(2853) <= not((layer0_outputs(4459)) or (layer0_outputs(3705)));
    outputs(2854) <= not(layer0_outputs(1455)) or (layer0_outputs(4552));
    outputs(2855) <= not((layer0_outputs(7176)) xor (layer0_outputs(6604)));
    outputs(2856) <= not((layer0_outputs(7237)) or (layer0_outputs(7117)));
    outputs(2857) <= layer0_outputs(5338);
    outputs(2858) <= (layer0_outputs(4226)) and not (layer0_outputs(8343));
    outputs(2859) <= layer0_outputs(1610);
    outputs(2860) <= not(layer0_outputs(3243));
    outputs(2861) <= layer0_outputs(7098);
    outputs(2862) <= (layer0_outputs(8422)) xor (layer0_outputs(1354));
    outputs(2863) <= not(layer0_outputs(8293));
    outputs(2864) <= (layer0_outputs(312)) or (layer0_outputs(9564));
    outputs(2865) <= (layer0_outputs(5251)) and not (layer0_outputs(5773));
    outputs(2866) <= (layer0_outputs(5047)) and not (layer0_outputs(1230));
    outputs(2867) <= not(layer0_outputs(3017));
    outputs(2868) <= not((layer0_outputs(5082)) xor (layer0_outputs(2641)));
    outputs(2869) <= layer0_outputs(9833);
    outputs(2870) <= not((layer0_outputs(6226)) and (layer0_outputs(9335)));
    outputs(2871) <= (layer0_outputs(1938)) xor (layer0_outputs(7941));
    outputs(2872) <= layer0_outputs(7769);
    outputs(2873) <= layer0_outputs(7326);
    outputs(2874) <= not((layer0_outputs(2074)) and (layer0_outputs(9156)));
    outputs(2875) <= layer0_outputs(7665);
    outputs(2876) <= not(layer0_outputs(9178));
    outputs(2877) <= not((layer0_outputs(1076)) and (layer0_outputs(6251)));
    outputs(2878) <= (layer0_outputs(7022)) or (layer0_outputs(6297));
    outputs(2879) <= not((layer0_outputs(1738)) and (layer0_outputs(8675)));
    outputs(2880) <= not(layer0_outputs(815));
    outputs(2881) <= not((layer0_outputs(6088)) or (layer0_outputs(143)));
    outputs(2882) <= layer0_outputs(4221);
    outputs(2883) <= not((layer0_outputs(9630)) or (layer0_outputs(2693)));
    outputs(2884) <= (layer0_outputs(3205)) xor (layer0_outputs(4640));
    outputs(2885) <= layer0_outputs(3677);
    outputs(2886) <= not(layer0_outputs(924));
    outputs(2887) <= (layer0_outputs(7929)) and not (layer0_outputs(4696));
    outputs(2888) <= (layer0_outputs(8523)) xor (layer0_outputs(8587));
    outputs(2889) <= (layer0_outputs(2819)) or (layer0_outputs(4159));
    outputs(2890) <= not((layer0_outputs(5973)) xor (layer0_outputs(213)));
    outputs(2891) <= not(layer0_outputs(1416));
    outputs(2892) <= layer0_outputs(952);
    outputs(2893) <= not((layer0_outputs(7833)) and (layer0_outputs(8593)));
    outputs(2894) <= layer0_outputs(1608);
    outputs(2895) <= (layer0_outputs(5431)) and (layer0_outputs(6521));
    outputs(2896) <= not(layer0_outputs(293));
    outputs(2897) <= (layer0_outputs(7226)) or (layer0_outputs(1591));
    outputs(2898) <= layer0_outputs(2535);
    outputs(2899) <= (layer0_outputs(5394)) and not (layer0_outputs(9143));
    outputs(2900) <= (layer0_outputs(7113)) and not (layer0_outputs(2048));
    outputs(2901) <= not(layer0_outputs(508));
    outputs(2902) <= not(layer0_outputs(2411)) or (layer0_outputs(1595));
    outputs(2903) <= (layer0_outputs(685)) xor (layer0_outputs(1771));
    outputs(2904) <= not((layer0_outputs(8788)) xor (layer0_outputs(1195)));
    outputs(2905) <= (layer0_outputs(2629)) or (layer0_outputs(2775));
    outputs(2906) <= not(layer0_outputs(7580)) or (layer0_outputs(2647));
    outputs(2907) <= (layer0_outputs(6142)) or (layer0_outputs(1261));
    outputs(2908) <= (layer0_outputs(9995)) and not (layer0_outputs(2151));
    outputs(2909) <= not(layer0_outputs(6729));
    outputs(2910) <= layer0_outputs(9377);
    outputs(2911) <= (layer0_outputs(4641)) or (layer0_outputs(455));
    outputs(2912) <= not(layer0_outputs(5420));
    outputs(2913) <= (layer0_outputs(3813)) and (layer0_outputs(2945));
    outputs(2914) <= layer0_outputs(5646);
    outputs(2915) <= not(layer0_outputs(5454)) or (layer0_outputs(1092));
    outputs(2916) <= not((layer0_outputs(1684)) xor (layer0_outputs(603)));
    outputs(2917) <= not(layer0_outputs(5260));
    outputs(2918) <= layer0_outputs(2933);
    outputs(2919) <= layer0_outputs(6445);
    outputs(2920) <= (layer0_outputs(1886)) xor (layer0_outputs(7978));
    outputs(2921) <= not((layer0_outputs(8686)) xor (layer0_outputs(10096)));
    outputs(2922) <= not((layer0_outputs(6189)) xor (layer0_outputs(1820)));
    outputs(2923) <= (layer0_outputs(1583)) xor (layer0_outputs(9129));
    outputs(2924) <= layer0_outputs(9830);
    outputs(2925) <= not(layer0_outputs(1877));
    outputs(2926) <= not((layer0_outputs(6496)) and (layer0_outputs(4467)));
    outputs(2927) <= layer0_outputs(9990);
    outputs(2928) <= not((layer0_outputs(5829)) and (layer0_outputs(5476)));
    outputs(2929) <= (layer0_outputs(8559)) or (layer0_outputs(9621));
    outputs(2930) <= not(layer0_outputs(4602));
    outputs(2931) <= (layer0_outputs(2245)) xor (layer0_outputs(7810));
    outputs(2932) <= layer0_outputs(573);
    outputs(2933) <= not((layer0_outputs(3656)) and (layer0_outputs(2289)));
    outputs(2934) <= layer0_outputs(8315);
    outputs(2935) <= not(layer0_outputs(3177)) or (layer0_outputs(1201));
    outputs(2936) <= not((layer0_outputs(595)) or (layer0_outputs(7282)));
    outputs(2937) <= layer0_outputs(2960);
    outputs(2938) <= not(layer0_outputs(5034));
    outputs(2939) <= layer0_outputs(4996);
    outputs(2940) <= not(layer0_outputs(9315)) or (layer0_outputs(9261));
    outputs(2941) <= layer0_outputs(1904);
    outputs(2942) <= layer0_outputs(9320);
    outputs(2943) <= not(layer0_outputs(2522));
    outputs(2944) <= not((layer0_outputs(9797)) xor (layer0_outputs(3391)));
    outputs(2945) <= not(layer0_outputs(7814));
    outputs(2946) <= not(layer0_outputs(9361)) or (layer0_outputs(9147));
    outputs(2947) <= layer0_outputs(3871);
    outputs(2948) <= layer0_outputs(5500);
    outputs(2949) <= layer0_outputs(8968);
    outputs(2950) <= not((layer0_outputs(3358)) or (layer0_outputs(2913)));
    outputs(2951) <= not(layer0_outputs(9216));
    outputs(2952) <= (layer0_outputs(8402)) xor (layer0_outputs(784));
    outputs(2953) <= (layer0_outputs(3591)) and (layer0_outputs(2925));
    outputs(2954) <= not(layer0_outputs(5783));
    outputs(2955) <= not((layer0_outputs(6739)) or (layer0_outputs(5636)));
    outputs(2956) <= (layer0_outputs(2386)) and (layer0_outputs(3733));
    outputs(2957) <= not((layer0_outputs(9180)) xor (layer0_outputs(4128)));
    outputs(2958) <= not(layer0_outputs(2595)) or (layer0_outputs(5497));
    outputs(2959) <= not(layer0_outputs(9255)) or (layer0_outputs(429));
    outputs(2960) <= layer0_outputs(471);
    outputs(2961) <= not((layer0_outputs(2194)) xor (layer0_outputs(8550)));
    outputs(2962) <= not(layer0_outputs(1086));
    outputs(2963) <= (layer0_outputs(2337)) or (layer0_outputs(10126));
    outputs(2964) <= not(layer0_outputs(9956));
    outputs(2965) <= layer0_outputs(3924);
    outputs(2966) <= not((layer0_outputs(3204)) xor (layer0_outputs(6022)));
    outputs(2967) <= not(layer0_outputs(3020));
    outputs(2968) <= (layer0_outputs(9574)) and not (layer0_outputs(9101));
    outputs(2969) <= layer0_outputs(4829);
    outputs(2970) <= (layer0_outputs(10017)) xor (layer0_outputs(7443));
    outputs(2971) <= (layer0_outputs(4804)) or (layer0_outputs(1816));
    outputs(2972) <= not((layer0_outputs(6618)) or (layer0_outputs(6738)));
    outputs(2973) <= layer0_outputs(10007);
    outputs(2974) <= not(layer0_outputs(8644));
    outputs(2975) <= not((layer0_outputs(4026)) and (layer0_outputs(9285)));
    outputs(2976) <= not((layer0_outputs(570)) xor (layer0_outputs(2163)));
    outputs(2977) <= not(layer0_outputs(6497)) or (layer0_outputs(7573));
    outputs(2978) <= not((layer0_outputs(10098)) xor (layer0_outputs(8554)));
    outputs(2979) <= layer0_outputs(1191);
    outputs(2980) <= not(layer0_outputs(2850)) or (layer0_outputs(3337));
    outputs(2981) <= not((layer0_outputs(9919)) and (layer0_outputs(4974)));
    outputs(2982) <= layer0_outputs(5972);
    outputs(2983) <= not(layer0_outputs(4842));
    outputs(2984) <= not(layer0_outputs(5390));
    outputs(2985) <= not(layer0_outputs(5277));
    outputs(2986) <= not(layer0_outputs(10136));
    outputs(2987) <= layer0_outputs(8105);
    outputs(2988) <= layer0_outputs(7235);
    outputs(2989) <= not((layer0_outputs(7193)) or (layer0_outputs(5639)));
    outputs(2990) <= not(layer0_outputs(346));
    outputs(2991) <= not(layer0_outputs(6923)) or (layer0_outputs(601));
    outputs(2992) <= not((layer0_outputs(730)) xor (layer0_outputs(1071)));
    outputs(2993) <= (layer0_outputs(8482)) xor (layer0_outputs(2986));
    outputs(2994) <= not((layer0_outputs(2284)) and (layer0_outputs(1943)));
    outputs(2995) <= not(layer0_outputs(6969));
    outputs(2996) <= not(layer0_outputs(2670));
    outputs(2997) <= not(layer0_outputs(324));
    outputs(2998) <= not((layer0_outputs(2493)) xor (layer0_outputs(69)));
    outputs(2999) <= not(layer0_outputs(9124));
    outputs(3000) <= not((layer0_outputs(5090)) and (layer0_outputs(1527)));
    outputs(3001) <= not(layer0_outputs(4172)) or (layer0_outputs(2241));
    outputs(3002) <= layer0_outputs(7175);
    outputs(3003) <= not(layer0_outputs(4063)) or (layer0_outputs(6011));
    outputs(3004) <= (layer0_outputs(8015)) xor (layer0_outputs(792));
    outputs(3005) <= layer0_outputs(2596);
    outputs(3006) <= not(layer0_outputs(5657)) or (layer0_outputs(4887));
    outputs(3007) <= layer0_outputs(8756);
    outputs(3008) <= layer0_outputs(2727);
    outputs(3009) <= not(layer0_outputs(8609)) or (layer0_outputs(6509));
    outputs(3010) <= layer0_outputs(9623);
    outputs(3011) <= (layer0_outputs(9437)) or (layer0_outputs(4600));
    outputs(3012) <= (layer0_outputs(6967)) and not (layer0_outputs(3208));
    outputs(3013) <= '1';
    outputs(3014) <= (layer0_outputs(10196)) or (layer0_outputs(6255));
    outputs(3015) <= layer0_outputs(479);
    outputs(3016) <= not(layer0_outputs(1832)) or (layer0_outputs(1379));
    outputs(3017) <= not(layer0_outputs(1768));
    outputs(3018) <= layer0_outputs(669);
    outputs(3019) <= not(layer0_outputs(9303));
    outputs(3020) <= layer0_outputs(7300);
    outputs(3021) <= not((layer0_outputs(6424)) or (layer0_outputs(2460)));
    outputs(3022) <= (layer0_outputs(8054)) and not (layer0_outputs(5639));
    outputs(3023) <= (layer0_outputs(3063)) xor (layer0_outputs(2633));
    outputs(3024) <= layer0_outputs(7609);
    outputs(3025) <= not((layer0_outputs(9583)) and (layer0_outputs(1280)));
    outputs(3026) <= not((layer0_outputs(6465)) or (layer0_outputs(806)));
    outputs(3027) <= (layer0_outputs(7787)) xor (layer0_outputs(3301));
    outputs(3028) <= not((layer0_outputs(2718)) xor (layer0_outputs(4578)));
    outputs(3029) <= not(layer0_outputs(136)) or (layer0_outputs(789));
    outputs(3030) <= layer0_outputs(447);
    outputs(3031) <= layer0_outputs(8149);
    outputs(3032) <= not(layer0_outputs(2747));
    outputs(3033) <= not(layer0_outputs(7876)) or (layer0_outputs(6586));
    outputs(3034) <= not(layer0_outputs(4703));
    outputs(3035) <= layer0_outputs(6230);
    outputs(3036) <= (layer0_outputs(4666)) xor (layer0_outputs(7478));
    outputs(3037) <= not(layer0_outputs(1674));
    outputs(3038) <= not(layer0_outputs(2890));
    outputs(3039) <= not(layer0_outputs(1163));
    outputs(3040) <= not(layer0_outputs(460)) or (layer0_outputs(8601));
    outputs(3041) <= (layer0_outputs(7273)) xor (layer0_outputs(2023));
    outputs(3042) <= (layer0_outputs(8693)) xor (layer0_outputs(6057));
    outputs(3043) <= not(layer0_outputs(4511));
    outputs(3044) <= not((layer0_outputs(1044)) or (layer0_outputs(8957)));
    outputs(3045) <= not((layer0_outputs(5876)) or (layer0_outputs(5661)));
    outputs(3046) <= (layer0_outputs(9784)) xor (layer0_outputs(5118));
    outputs(3047) <= not(layer0_outputs(2246));
    outputs(3048) <= not(layer0_outputs(1674));
    outputs(3049) <= layer0_outputs(1440);
    outputs(3050) <= not(layer0_outputs(3590)) or (layer0_outputs(5792));
    outputs(3051) <= not(layer0_outputs(3635));
    outputs(3052) <= not((layer0_outputs(9826)) or (layer0_outputs(6286)));
    outputs(3053) <= not(layer0_outputs(6579));
    outputs(3054) <= (layer0_outputs(6803)) and (layer0_outputs(524));
    outputs(3055) <= not((layer0_outputs(63)) xor (layer0_outputs(8797)));
    outputs(3056) <= (layer0_outputs(640)) or (layer0_outputs(5254));
    outputs(3057) <= not(layer0_outputs(3419));
    outputs(3058) <= not(layer0_outputs(9976)) or (layer0_outputs(3323));
    outputs(3059) <= layer0_outputs(5490);
    outputs(3060) <= not(layer0_outputs(2611));
    outputs(3061) <= (layer0_outputs(4109)) xor (layer0_outputs(3337));
    outputs(3062) <= not((layer0_outputs(4897)) xor (layer0_outputs(9879)));
    outputs(3063) <= layer0_outputs(9701);
    outputs(3064) <= not(layer0_outputs(5281)) or (layer0_outputs(826));
    outputs(3065) <= layer0_outputs(3953);
    outputs(3066) <= (layer0_outputs(5093)) or (layer0_outputs(1159));
    outputs(3067) <= (layer0_outputs(5823)) xor (layer0_outputs(10154));
    outputs(3068) <= not(layer0_outputs(2961)) or (layer0_outputs(4105));
    outputs(3069) <= not(layer0_outputs(9011));
    outputs(3070) <= not(layer0_outputs(1049));
    outputs(3071) <= not(layer0_outputs(1467));
    outputs(3072) <= not(layer0_outputs(10003));
    outputs(3073) <= layer0_outputs(10056);
    outputs(3074) <= not(layer0_outputs(898));
    outputs(3075) <= not(layer0_outputs(9991));
    outputs(3076) <= layer0_outputs(3371);
    outputs(3077) <= not(layer0_outputs(4615)) or (layer0_outputs(4683));
    outputs(3078) <= layer0_outputs(8203);
    outputs(3079) <= not(layer0_outputs(2208)) or (layer0_outputs(667));
    outputs(3080) <= layer0_outputs(3777);
    outputs(3081) <= not((layer0_outputs(7832)) and (layer0_outputs(769)));
    outputs(3082) <= not((layer0_outputs(9228)) xor (layer0_outputs(9882)));
    outputs(3083) <= not((layer0_outputs(4890)) xor (layer0_outputs(4667)));
    outputs(3084) <= not(layer0_outputs(5571));
    outputs(3085) <= not((layer0_outputs(6611)) xor (layer0_outputs(7319)));
    outputs(3086) <= layer0_outputs(5556);
    outputs(3087) <= layer0_outputs(2206);
    outputs(3088) <= layer0_outputs(3952);
    outputs(3089) <= layer0_outputs(3964);
    outputs(3090) <= (layer0_outputs(7470)) and (layer0_outputs(6233));
    outputs(3091) <= not(layer0_outputs(936)) or (layer0_outputs(5396));
    outputs(3092) <= not((layer0_outputs(1998)) xor (layer0_outputs(3482)));
    outputs(3093) <= not(layer0_outputs(7270));
    outputs(3094) <= not(layer0_outputs(3239));
    outputs(3095) <= (layer0_outputs(1919)) or (layer0_outputs(8532));
    outputs(3096) <= not(layer0_outputs(1897));
    outputs(3097) <= (layer0_outputs(701)) and not (layer0_outputs(2469));
    outputs(3098) <= not(layer0_outputs(7718)) or (layer0_outputs(6063));
    outputs(3099) <= layer0_outputs(7046);
    outputs(3100) <= not(layer0_outputs(1297));
    outputs(3101) <= layer0_outputs(23);
    outputs(3102) <= not((layer0_outputs(5831)) xor (layer0_outputs(4752)));
    outputs(3103) <= not((layer0_outputs(5410)) xor (layer0_outputs(8433)));
    outputs(3104) <= not(layer0_outputs(1764));
    outputs(3105) <= (layer0_outputs(3887)) or (layer0_outputs(9333));
    outputs(3106) <= (layer0_outputs(9735)) xor (layer0_outputs(3074));
    outputs(3107) <= (layer0_outputs(4539)) and not (layer0_outputs(9745));
    outputs(3108) <= (layer0_outputs(5231)) xor (layer0_outputs(8971));
    outputs(3109) <= (layer0_outputs(7700)) and (layer0_outputs(9677));
    outputs(3110) <= (layer0_outputs(970)) xor (layer0_outputs(3416));
    outputs(3111) <= not(layer0_outputs(6049));
    outputs(3112) <= (layer0_outputs(8084)) xor (layer0_outputs(7224));
    outputs(3113) <= (layer0_outputs(2274)) xor (layer0_outputs(3131));
    outputs(3114) <= (layer0_outputs(6278)) or (layer0_outputs(1963));
    outputs(3115) <= not((layer0_outputs(1091)) and (layer0_outputs(6093)));
    outputs(3116) <= (layer0_outputs(1419)) xor (layer0_outputs(9556));
    outputs(3117) <= not(layer0_outputs(5014));
    outputs(3118) <= layer0_outputs(9185);
    outputs(3119) <= not(layer0_outputs(9742)) or (layer0_outputs(3772));
    outputs(3120) <= not((layer0_outputs(4210)) xor (layer0_outputs(9383)));
    outputs(3121) <= not(layer0_outputs(2278)) or (layer0_outputs(5492));
    outputs(3122) <= not(layer0_outputs(7342));
    outputs(3123) <= not(layer0_outputs(9791));
    outputs(3124) <= not(layer0_outputs(3293)) or (layer0_outputs(3390));
    outputs(3125) <= not(layer0_outputs(3694));
    outputs(3126) <= not((layer0_outputs(5214)) and (layer0_outputs(5177)));
    outputs(3127) <= not((layer0_outputs(3870)) xor (layer0_outputs(1667)));
    outputs(3128) <= layer0_outputs(10060);
    outputs(3129) <= not((layer0_outputs(3670)) xor (layer0_outputs(10105)));
    outputs(3130) <= layer0_outputs(5834);
    outputs(3131) <= layer0_outputs(1859);
    outputs(3132) <= not((layer0_outputs(8953)) and (layer0_outputs(6665)));
    outputs(3133) <= layer0_outputs(558);
    outputs(3134) <= layer0_outputs(8883);
    outputs(3135) <= not(layer0_outputs(5501));
    outputs(3136) <= not(layer0_outputs(6323)) or (layer0_outputs(2029));
    outputs(3137) <= layer0_outputs(9243);
    outputs(3138) <= layer0_outputs(5079);
    outputs(3139) <= layer0_outputs(7856);
    outputs(3140) <= '0';
    outputs(3141) <= not(layer0_outputs(5682));
    outputs(3142) <= not((layer0_outputs(8676)) xor (layer0_outputs(9957)));
    outputs(3143) <= not(layer0_outputs(4327));
    outputs(3144) <= not(layer0_outputs(5706));
    outputs(3145) <= (layer0_outputs(8284)) xor (layer0_outputs(5495));
    outputs(3146) <= not((layer0_outputs(9049)) xor (layer0_outputs(9247)));
    outputs(3147) <= layer0_outputs(1461);
    outputs(3148) <= not((layer0_outputs(1977)) and (layer0_outputs(74)));
    outputs(3149) <= layer0_outputs(1256);
    outputs(3150) <= layer0_outputs(8949);
    outputs(3151) <= not((layer0_outputs(6766)) or (layer0_outputs(7406)));
    outputs(3152) <= not(layer0_outputs(1001));
    outputs(3153) <= (layer0_outputs(4072)) and not (layer0_outputs(3598));
    outputs(3154) <= not(layer0_outputs(1540));
    outputs(3155) <= not(layer0_outputs(7211));
    outputs(3156) <= not(layer0_outputs(7749));
    outputs(3157) <= layer0_outputs(7668);
    outputs(3158) <= layer0_outputs(930);
    outputs(3159) <= layer0_outputs(1099);
    outputs(3160) <= layer0_outputs(4913);
    outputs(3161) <= layer0_outputs(6656);
    outputs(3162) <= not(layer0_outputs(1921));
    outputs(3163) <= (layer0_outputs(3881)) xor (layer0_outputs(9940));
    outputs(3164) <= layer0_outputs(2031);
    outputs(3165) <= layer0_outputs(9017);
    outputs(3166) <= not(layer0_outputs(1233)) or (layer0_outputs(994));
    outputs(3167) <= layer0_outputs(1760);
    outputs(3168) <= layer0_outputs(4601);
    outputs(3169) <= not((layer0_outputs(2895)) and (layer0_outputs(8538)));
    outputs(3170) <= not((layer0_outputs(3769)) xor (layer0_outputs(6404)));
    outputs(3171) <= layer0_outputs(8251);
    outputs(3172) <= layer0_outputs(2089);
    outputs(3173) <= not(layer0_outputs(9321)) or (layer0_outputs(9739));
    outputs(3174) <= layer0_outputs(398);
    outputs(3175) <= (layer0_outputs(4555)) xor (layer0_outputs(4149));
    outputs(3176) <= not(layer0_outputs(4094)) or (layer0_outputs(5));
    outputs(3177) <= (layer0_outputs(9042)) xor (layer0_outputs(5903));
    outputs(3178) <= not(layer0_outputs(5989));
    outputs(3179) <= not(layer0_outputs(3216));
    outputs(3180) <= (layer0_outputs(1220)) and not (layer0_outputs(3868));
    outputs(3181) <= (layer0_outputs(624)) xor (layer0_outputs(2656));
    outputs(3182) <= not(layer0_outputs(8465));
    outputs(3183) <= not(layer0_outputs(6489));
    outputs(3184) <= not((layer0_outputs(6365)) and (layer0_outputs(1617)));
    outputs(3185) <= (layer0_outputs(2382)) xor (layer0_outputs(2719));
    outputs(3186) <= (layer0_outputs(521)) xor (layer0_outputs(7232));
    outputs(3187) <= layer0_outputs(8059);
    outputs(3188) <= layer0_outputs(9916);
    outputs(3189) <= (layer0_outputs(6459)) and not (layer0_outputs(1610));
    outputs(3190) <= not(layer0_outputs(1943));
    outputs(3191) <= not(layer0_outputs(229));
    outputs(3192) <= not((layer0_outputs(7294)) xor (layer0_outputs(8232)));
    outputs(3193) <= (layer0_outputs(2936)) xor (layer0_outputs(6539));
    outputs(3194) <= layer0_outputs(10111);
    outputs(3195) <= (layer0_outputs(9202)) and (layer0_outputs(7049));
    outputs(3196) <= not((layer0_outputs(5179)) xor (layer0_outputs(5448)));
    outputs(3197) <= not((layer0_outputs(10203)) xor (layer0_outputs(7026)));
    outputs(3198) <= layer0_outputs(8880);
    outputs(3199) <= not((layer0_outputs(8852)) xor (layer0_outputs(3343)));
    outputs(3200) <= not(layer0_outputs(9309)) or (layer0_outputs(2037));
    outputs(3201) <= not(layer0_outputs(2965));
    outputs(3202) <= not(layer0_outputs(9468));
    outputs(3203) <= (layer0_outputs(10238)) xor (layer0_outputs(8830));
    outputs(3204) <= layer0_outputs(10234);
    outputs(3205) <= not(layer0_outputs(7661)) or (layer0_outputs(6770));
    outputs(3206) <= (layer0_outputs(2221)) xor (layer0_outputs(9596));
    outputs(3207) <= not((layer0_outputs(4163)) xor (layer0_outputs(6326)));
    outputs(3208) <= not((layer0_outputs(4849)) and (layer0_outputs(6479)));
    outputs(3209) <= (layer0_outputs(7164)) and not (layer0_outputs(10162));
    outputs(3210) <= not(layer0_outputs(5088));
    outputs(3211) <= not((layer0_outputs(5152)) xor (layer0_outputs(4734)));
    outputs(3212) <= layer0_outputs(6845);
    outputs(3213) <= not((layer0_outputs(8524)) xor (layer0_outputs(3466)));
    outputs(3214) <= (layer0_outputs(8706)) xor (layer0_outputs(7606));
    outputs(3215) <= not(layer0_outputs(4896));
    outputs(3216) <= layer0_outputs(5561);
    outputs(3217) <= not(layer0_outputs(1129));
    outputs(3218) <= not((layer0_outputs(9047)) xor (layer0_outputs(6734)));
    outputs(3219) <= layer0_outputs(8388);
    outputs(3220) <= (layer0_outputs(2113)) xor (layer0_outputs(654));
    outputs(3221) <= not(layer0_outputs(9959)) or (layer0_outputs(9670));
    outputs(3222) <= not(layer0_outputs(2132));
    outputs(3223) <= not((layer0_outputs(7334)) xor (layer0_outputs(9942)));
    outputs(3224) <= (layer0_outputs(10000)) and not (layer0_outputs(4628));
    outputs(3225) <= (layer0_outputs(3125)) xor (layer0_outputs(6014));
    outputs(3226) <= not((layer0_outputs(696)) xor (layer0_outputs(2374)));
    outputs(3227) <= (layer0_outputs(608)) xor (layer0_outputs(9334));
    outputs(3228) <= not((layer0_outputs(9077)) xor (layer0_outputs(2127)));
    outputs(3229) <= layer0_outputs(70);
    outputs(3230) <= not(layer0_outputs(8759)) or (layer0_outputs(2247));
    outputs(3231) <= not(layer0_outputs(4200));
    outputs(3232) <= layer0_outputs(6361);
    outputs(3233) <= not(layer0_outputs(4041)) or (layer0_outputs(7053));
    outputs(3234) <= (layer0_outputs(3496)) or (layer0_outputs(4822));
    outputs(3235) <= (layer0_outputs(8754)) or (layer0_outputs(5080));
    outputs(3236) <= layer0_outputs(3203);
    outputs(3237) <= layer0_outputs(410);
    outputs(3238) <= layer0_outputs(7171);
    outputs(3239) <= layer0_outputs(1188);
    outputs(3240) <= layer0_outputs(1801);
    outputs(3241) <= not((layer0_outputs(6331)) and (layer0_outputs(7973)));
    outputs(3242) <= not(layer0_outputs(1186));
    outputs(3243) <= not((layer0_outputs(1373)) xor (layer0_outputs(3596)));
    outputs(3244) <= not(layer0_outputs(4041));
    outputs(3245) <= not(layer0_outputs(2553));
    outputs(3246) <= not(layer0_outputs(9445));
    outputs(3247) <= not(layer0_outputs(8491));
    outputs(3248) <= not(layer0_outputs(3404));
    outputs(3249) <= not((layer0_outputs(2976)) xor (layer0_outputs(6657)));
    outputs(3250) <= not(layer0_outputs(6051));
    outputs(3251) <= not(layer0_outputs(524)) or (layer0_outputs(7011));
    outputs(3252) <= not((layer0_outputs(6867)) xor (layer0_outputs(4714)));
    outputs(3253) <= not((layer0_outputs(8189)) xor (layer0_outputs(8711)));
    outputs(3254) <= (layer0_outputs(7137)) xor (layer0_outputs(9673));
    outputs(3255) <= layer0_outputs(725);
    outputs(3256) <= not(layer0_outputs(2720)) or (layer0_outputs(1211));
    outputs(3257) <= (layer0_outputs(4463)) and not (layer0_outputs(7334));
    outputs(3258) <= (layer0_outputs(6959)) xor (layer0_outputs(6360));
    outputs(3259) <= not(layer0_outputs(3085));
    outputs(3260) <= layer0_outputs(7429);
    outputs(3261) <= (layer0_outputs(5475)) and not (layer0_outputs(2055));
    outputs(3262) <= layer0_outputs(854);
    outputs(3263) <= (layer0_outputs(7717)) xor (layer0_outputs(2461));
    outputs(3264) <= (layer0_outputs(4239)) xor (layer0_outputs(5703));
    outputs(3265) <= not((layer0_outputs(5224)) xor (layer0_outputs(7146)));
    outputs(3266) <= (layer0_outputs(7762)) and (layer0_outputs(3163));
    outputs(3267) <= not(layer0_outputs(6507)) or (layer0_outputs(6125));
    outputs(3268) <= layer0_outputs(6311);
    outputs(3269) <= not((layer0_outputs(411)) and (layer0_outputs(6913)));
    outputs(3270) <= layer0_outputs(931);
    outputs(3271) <= not(layer0_outputs(8333));
    outputs(3272) <= (layer0_outputs(363)) or (layer0_outputs(9057));
    outputs(3273) <= (layer0_outputs(6332)) xor (layer0_outputs(6680));
    outputs(3274) <= not((layer0_outputs(2306)) xor (layer0_outputs(247)));
    outputs(3275) <= not(layer0_outputs(8498)) or (layer0_outputs(2705));
    outputs(3276) <= (layer0_outputs(9927)) xor (layer0_outputs(2200));
    outputs(3277) <= not(layer0_outputs(8028));
    outputs(3278) <= not((layer0_outputs(5665)) and (layer0_outputs(9596)));
    outputs(3279) <= layer0_outputs(6714);
    outputs(3280) <= not(layer0_outputs(3025));
    outputs(3281) <= layer0_outputs(3732);
    outputs(3282) <= not(layer0_outputs(2715));
    outputs(3283) <= not(layer0_outputs(8238));
    outputs(3284) <= not(layer0_outputs(5773));
    outputs(3285) <= layer0_outputs(9418);
    outputs(3286) <= (layer0_outputs(5468)) and not (layer0_outputs(6297));
    outputs(3287) <= (layer0_outputs(2043)) xor (layer0_outputs(6237));
    outputs(3288) <= layer0_outputs(8869);
    outputs(3289) <= not(layer0_outputs(7069)) or (layer0_outputs(2532));
    outputs(3290) <= not((layer0_outputs(6064)) xor (layer0_outputs(2927)));
    outputs(3291) <= not((layer0_outputs(2048)) or (layer0_outputs(10023)));
    outputs(3292) <= (layer0_outputs(2816)) or (layer0_outputs(5965));
    outputs(3293) <= (layer0_outputs(8885)) and not (layer0_outputs(9928));
    outputs(3294) <= not(layer0_outputs(3687));
    outputs(3295) <= (layer0_outputs(7964)) and not (layer0_outputs(215));
    outputs(3296) <= (layer0_outputs(5882)) xor (layer0_outputs(3396));
    outputs(3297) <= layer0_outputs(6327);
    outputs(3298) <= (layer0_outputs(556)) and not (layer0_outputs(516));
    outputs(3299) <= not((layer0_outputs(5731)) xor (layer0_outputs(10040)));
    outputs(3300) <= (layer0_outputs(4225)) or (layer0_outputs(5585));
    outputs(3301) <= (layer0_outputs(4936)) and not (layer0_outputs(6557));
    outputs(3302) <= not((layer0_outputs(5530)) xor (layer0_outputs(8756)));
    outputs(3303) <= (layer0_outputs(5984)) and not (layer0_outputs(9780));
    outputs(3304) <= (layer0_outputs(10010)) xor (layer0_outputs(2290));
    outputs(3305) <= not(layer0_outputs(4679)) or (layer0_outputs(9355));
    outputs(3306) <= (layer0_outputs(4875)) and (layer0_outputs(1930));
    outputs(3307) <= layer0_outputs(3300);
    outputs(3308) <= layer0_outputs(8857);
    outputs(3309) <= (layer0_outputs(5325)) xor (layer0_outputs(7807));
    outputs(3310) <= layer0_outputs(4972);
    outputs(3311) <= not((layer0_outputs(8213)) xor (layer0_outputs(148)));
    outputs(3312) <= (layer0_outputs(6401)) xor (layer0_outputs(3674));
    outputs(3313) <= not((layer0_outputs(3035)) xor (layer0_outputs(5723)));
    outputs(3314) <= not((layer0_outputs(2425)) and (layer0_outputs(342)));
    outputs(3315) <= not(layer0_outputs(6257)) or (layer0_outputs(2698));
    outputs(3316) <= layer0_outputs(2697);
    outputs(3317) <= not(layer0_outputs(1528)) or (layer0_outputs(7666));
    outputs(3318) <= not(layer0_outputs(2749));
    outputs(3319) <= not((layer0_outputs(5225)) xor (layer0_outputs(9248)));
    outputs(3320) <= not(layer0_outputs(9198));
    outputs(3321) <= not(layer0_outputs(6649));
    outputs(3322) <= (layer0_outputs(3061)) xor (layer0_outputs(1111));
    outputs(3323) <= not(layer0_outputs(8553));
    outputs(3324) <= (layer0_outputs(5940)) xor (layer0_outputs(1365));
    outputs(3325) <= layer0_outputs(7492);
    outputs(3326) <= not((layer0_outputs(2645)) and (layer0_outputs(9876)));
    outputs(3327) <= not(layer0_outputs(7406)) or (layer0_outputs(3839));
    outputs(3328) <= not(layer0_outputs(5769)) or (layer0_outputs(2217));
    outputs(3329) <= layer0_outputs(1571);
    outputs(3330) <= not((layer0_outputs(5863)) or (layer0_outputs(1405)));
    outputs(3331) <= not((layer0_outputs(4932)) xor (layer0_outputs(5290)));
    outputs(3332) <= layer0_outputs(2627);
    outputs(3333) <= not(layer0_outputs(991));
    outputs(3334) <= (layer0_outputs(820)) or (layer0_outputs(596));
    outputs(3335) <= not(layer0_outputs(7889));
    outputs(3336) <= not(layer0_outputs(9700)) or (layer0_outputs(4952));
    outputs(3337) <= layer0_outputs(1920);
    outputs(3338) <= '1';
    outputs(3339) <= not(layer0_outputs(256));
    outputs(3340) <= not(layer0_outputs(2669));
    outputs(3341) <= layer0_outputs(1969);
    outputs(3342) <= (layer0_outputs(7251)) and not (layer0_outputs(2160));
    outputs(3343) <= not((layer0_outputs(6379)) and (layer0_outputs(9893)));
    outputs(3344) <= not(layer0_outputs(6970)) or (layer0_outputs(3898));
    outputs(3345) <= (layer0_outputs(3406)) and not (layer0_outputs(8167));
    outputs(3346) <= not(layer0_outputs(6005));
    outputs(3347) <= not(layer0_outputs(7497));
    outputs(3348) <= not((layer0_outputs(4859)) and (layer0_outputs(1800)));
    outputs(3349) <= not(layer0_outputs(7179));
    outputs(3350) <= not((layer0_outputs(8286)) xor (layer0_outputs(7640)));
    outputs(3351) <= not(layer0_outputs(3567));
    outputs(3352) <= layer0_outputs(5202);
    outputs(3353) <= (layer0_outputs(1784)) and not (layer0_outputs(7651));
    outputs(3354) <= not(layer0_outputs(3593)) or (layer0_outputs(5921));
    outputs(3355) <= (layer0_outputs(9571)) or (layer0_outputs(7691));
    outputs(3356) <= layer0_outputs(886);
    outputs(3357) <= not((layer0_outputs(135)) xor (layer0_outputs(1264)));
    outputs(3358) <= layer0_outputs(1309);
    outputs(3359) <= layer0_outputs(381);
    outputs(3360) <= not(layer0_outputs(4133)) or (layer0_outputs(4069));
    outputs(3361) <= (layer0_outputs(7664)) xor (layer0_outputs(4396));
    outputs(3362) <= (layer0_outputs(1723)) and (layer0_outputs(4176));
    outputs(3363) <= not(layer0_outputs(3988)) or (layer0_outputs(2622));
    outputs(3364) <= (layer0_outputs(7831)) xor (layer0_outputs(2597));
    outputs(3365) <= (layer0_outputs(7129)) xor (layer0_outputs(509));
    outputs(3366) <= (layer0_outputs(4472)) or (layer0_outputs(6522));
    outputs(3367) <= not((layer0_outputs(6195)) or (layer0_outputs(416)));
    outputs(3368) <= (layer0_outputs(1335)) xor (layer0_outputs(3276));
    outputs(3369) <= not(layer0_outputs(8086));
    outputs(3370) <= not((layer0_outputs(4961)) xor (layer0_outputs(9561)));
    outputs(3371) <= not(layer0_outputs(9665)) or (layer0_outputs(2261));
    outputs(3372) <= layer0_outputs(8993);
    outputs(3373) <= not((layer0_outputs(9640)) and (layer0_outputs(5217)));
    outputs(3374) <= (layer0_outputs(3866)) and not (layer0_outputs(7508));
    outputs(3375) <= not(layer0_outputs(2184));
    outputs(3376) <= (layer0_outputs(7155)) or (layer0_outputs(8190));
    outputs(3377) <= (layer0_outputs(2767)) xor (layer0_outputs(8368));
    outputs(3378) <= not(layer0_outputs(183));
    outputs(3379) <= layer0_outputs(6495);
    outputs(3380) <= layer0_outputs(846);
    outputs(3381) <= layer0_outputs(2701);
    outputs(3382) <= (layer0_outputs(2443)) xor (layer0_outputs(9418));
    outputs(3383) <= (layer0_outputs(7095)) xor (layer0_outputs(3125));
    outputs(3384) <= not((layer0_outputs(3115)) xor (layer0_outputs(4568)));
    outputs(3385) <= (layer0_outputs(2572)) or (layer0_outputs(2577));
    outputs(3386) <= not(layer0_outputs(8070)) or (layer0_outputs(8126));
    outputs(3387) <= not(layer0_outputs(6277));
    outputs(3388) <= not((layer0_outputs(559)) xor (layer0_outputs(4733)));
    outputs(3389) <= (layer0_outputs(2071)) and not (layer0_outputs(2154));
    outputs(3390) <= (layer0_outputs(1048)) xor (layer0_outputs(4710));
    outputs(3391) <= layer0_outputs(2931);
    outputs(3392) <= not(layer0_outputs(2342)) or (layer0_outputs(8783));
    outputs(3393) <= not((layer0_outputs(4841)) and (layer0_outputs(7574)));
    outputs(3394) <= not(layer0_outputs(5597));
    outputs(3395) <= layer0_outputs(1086);
    outputs(3396) <= not(layer0_outputs(3363));
    outputs(3397) <= not((layer0_outputs(9482)) xor (layer0_outputs(7440)));
    outputs(3398) <= not((layer0_outputs(3912)) xor (layer0_outputs(1413)));
    outputs(3399) <= not(layer0_outputs(2170)) or (layer0_outputs(8160));
    outputs(3400) <= (layer0_outputs(2010)) or (layer0_outputs(7358));
    outputs(3401) <= not((layer0_outputs(2737)) and (layer0_outputs(7151)));
    outputs(3402) <= not((layer0_outputs(6755)) xor (layer0_outputs(8685)));
    outputs(3403) <= layer0_outputs(3981);
    outputs(3404) <= (layer0_outputs(990)) xor (layer0_outputs(9496));
    outputs(3405) <= not((layer0_outputs(60)) and (layer0_outputs(5809)));
    outputs(3406) <= not((layer0_outputs(1032)) xor (layer0_outputs(5853)));
    outputs(3407) <= not(layer0_outputs(8430));
    outputs(3408) <= layer0_outputs(1575);
    outputs(3409) <= (layer0_outputs(1334)) and not (layer0_outputs(1097));
    outputs(3410) <= (layer0_outputs(6765)) xor (layer0_outputs(10053));
    outputs(3411) <= not(layer0_outputs(8258));
    outputs(3412) <= (layer0_outputs(24)) xor (layer0_outputs(4492));
    outputs(3413) <= (layer0_outputs(6422)) xor (layer0_outputs(923));
    outputs(3414) <= not(layer0_outputs(6473)) or (layer0_outputs(9062));
    outputs(3415) <= not(layer0_outputs(7192));
    outputs(3416) <= not(layer0_outputs(4355));
    outputs(3417) <= not((layer0_outputs(7423)) and (layer0_outputs(7206)));
    outputs(3418) <= not((layer0_outputs(1064)) xor (layer0_outputs(3918)));
    outputs(3419) <= layer0_outputs(7722);
    outputs(3420) <= not(layer0_outputs(5186)) or (layer0_outputs(2910));
    outputs(3421) <= layer0_outputs(4921);
    outputs(3422) <= not((layer0_outputs(9429)) or (layer0_outputs(5616)));
    outputs(3423) <= (layer0_outputs(5155)) xor (layer0_outputs(9149));
    outputs(3424) <= not((layer0_outputs(8319)) xor (layer0_outputs(5546)));
    outputs(3425) <= layer0_outputs(6407);
    outputs(3426) <= not((layer0_outputs(4365)) xor (layer0_outputs(6081)));
    outputs(3427) <= not(layer0_outputs(8008));
    outputs(3428) <= layer0_outputs(1010);
    outputs(3429) <= (layer0_outputs(3575)) xor (layer0_outputs(8806));
    outputs(3430) <= (layer0_outputs(8100)) xor (layer0_outputs(4263));
    outputs(3431) <= layer0_outputs(584);
    outputs(3432) <= layer0_outputs(6086);
    outputs(3433) <= not(layer0_outputs(3191)) or (layer0_outputs(907));
    outputs(3434) <= layer0_outputs(8296);
    outputs(3435) <= layer0_outputs(4716);
    outputs(3436) <= (layer0_outputs(383)) and not (layer0_outputs(6855));
    outputs(3437) <= layer0_outputs(2081);
    outputs(3438) <= not(layer0_outputs(3819));
    outputs(3439) <= (layer0_outputs(7630)) xor (layer0_outputs(5376));
    outputs(3440) <= layer0_outputs(5962);
    outputs(3441) <= (layer0_outputs(4118)) and (layer0_outputs(4147));
    outputs(3442) <= not(layer0_outputs(3614)) or (layer0_outputs(7213));
    outputs(3443) <= layer0_outputs(3584);
    outputs(3444) <= layer0_outputs(9964);
    outputs(3445) <= '0';
    outputs(3446) <= not(layer0_outputs(8950));
    outputs(3447) <= not((layer0_outputs(7794)) or (layer0_outputs(5571)));
    outputs(3448) <= not((layer0_outputs(1918)) or (layer0_outputs(7026)));
    outputs(3449) <= (layer0_outputs(1403)) xor (layer0_outputs(5649));
    outputs(3450) <= layer0_outputs(7507);
    outputs(3451) <= not((layer0_outputs(9470)) and (layer0_outputs(1293)));
    outputs(3452) <= not((layer0_outputs(9145)) xor (layer0_outputs(7741)));
    outputs(3453) <= (layer0_outputs(7355)) and (layer0_outputs(338));
    outputs(3454) <= layer0_outputs(3315);
    outputs(3455) <= layer0_outputs(4432);
    outputs(3456) <= not((layer0_outputs(4045)) or (layer0_outputs(6433)));
    outputs(3457) <= (layer0_outputs(9091)) xor (layer0_outputs(3380));
    outputs(3458) <= (layer0_outputs(6571)) and (layer0_outputs(8002));
    outputs(3459) <= not(layer0_outputs(2504)) or (layer0_outputs(9328));
    outputs(3460) <= not(layer0_outputs(7517));
    outputs(3461) <= layer0_outputs(6516);
    outputs(3462) <= (layer0_outputs(9090)) and (layer0_outputs(197));
    outputs(3463) <= not((layer0_outputs(4163)) xor (layer0_outputs(2235)));
    outputs(3464) <= not(layer0_outputs(898));
    outputs(3465) <= not(layer0_outputs(3292));
    outputs(3466) <= not(layer0_outputs(376));
    outputs(3467) <= layer0_outputs(9793);
    outputs(3468) <= not((layer0_outputs(2721)) or (layer0_outputs(2610)));
    outputs(3469) <= layer0_outputs(10177);
    outputs(3470) <= not(layer0_outputs(7615));
    outputs(3471) <= (layer0_outputs(2454)) xor (layer0_outputs(7902));
    outputs(3472) <= (layer0_outputs(2617)) xor (layer0_outputs(5002));
    outputs(3473) <= (layer0_outputs(60)) xor (layer0_outputs(1175));
    outputs(3474) <= layer0_outputs(7134);
    outputs(3475) <= (layer0_outputs(5475)) and (layer0_outputs(4268));
    outputs(3476) <= (layer0_outputs(6629)) and (layer0_outputs(678));
    outputs(3477) <= layer0_outputs(5373);
    outputs(3478) <= layer0_outputs(5257);
    outputs(3479) <= not((layer0_outputs(6565)) and (layer0_outputs(9157)));
    outputs(3480) <= not(layer0_outputs(4923));
    outputs(3481) <= not((layer0_outputs(5779)) xor (layer0_outputs(9670)));
    outputs(3482) <= not(layer0_outputs(2687)) or (layer0_outputs(10120));
    outputs(3483) <= not((layer0_outputs(3707)) xor (layer0_outputs(331)));
    outputs(3484) <= not((layer0_outputs(4569)) and (layer0_outputs(7404)));
    outputs(3485) <= layer0_outputs(1562);
    outputs(3486) <= (layer0_outputs(6582)) xor (layer0_outputs(2967));
    outputs(3487) <= (layer0_outputs(340)) and not (layer0_outputs(6667));
    outputs(3488) <= layer0_outputs(287);
    outputs(3489) <= layer0_outputs(4161);
    outputs(3490) <= not((layer0_outputs(6588)) or (layer0_outputs(9592)));
    outputs(3491) <= (layer0_outputs(2118)) and not (layer0_outputs(5327));
    outputs(3492) <= not(layer0_outputs(3335));
    outputs(3493) <= layer0_outputs(4673);
    outputs(3494) <= (layer0_outputs(7619)) xor (layer0_outputs(7781));
    outputs(3495) <= not(layer0_outputs(6737));
    outputs(3496) <= not(layer0_outputs(8606)) or (layer0_outputs(7175));
    outputs(3497) <= layer0_outputs(6050);
    outputs(3498) <= (layer0_outputs(9368)) and (layer0_outputs(1884));
    outputs(3499) <= (layer0_outputs(1278)) and not (layer0_outputs(8017));
    outputs(3500) <= (layer0_outputs(8749)) xor (layer0_outputs(2699));
    outputs(3501) <= not(layer0_outputs(3031));
    outputs(3502) <= not(layer0_outputs(9219)) or (layer0_outputs(1200));
    outputs(3503) <= layer0_outputs(3681);
    outputs(3504) <= layer0_outputs(5187);
    outputs(3505) <= not((layer0_outputs(4680)) and (layer0_outputs(5438)));
    outputs(3506) <= not(layer0_outputs(2147));
    outputs(3507) <= layer0_outputs(4169);
    outputs(3508) <= not(layer0_outputs(6460)) or (layer0_outputs(273));
    outputs(3509) <= not(layer0_outputs(5219));
    outputs(3510) <= (layer0_outputs(5371)) xor (layer0_outputs(65));
    outputs(3511) <= (layer0_outputs(399)) or (layer0_outputs(1250));
    outputs(3512) <= layer0_outputs(405);
    outputs(3513) <= not(layer0_outputs(2670));
    outputs(3514) <= not(layer0_outputs(7467));
    outputs(3515) <= layer0_outputs(5603);
    outputs(3516) <= not(layer0_outputs(9202)) or (layer0_outputs(2249));
    outputs(3517) <= layer0_outputs(3402);
    outputs(3518) <= not(layer0_outputs(5055));
    outputs(3519) <= not((layer0_outputs(6922)) xor (layer0_outputs(2957)));
    outputs(3520) <= not(layer0_outputs(9626));
    outputs(3521) <= layer0_outputs(5041);
    outputs(3522) <= not(layer0_outputs(3011));
    outputs(3523) <= layer0_outputs(626);
    outputs(3524) <= layer0_outputs(7268);
    outputs(3525) <= not(layer0_outputs(3824)) or (layer0_outputs(6399));
    outputs(3526) <= not(layer0_outputs(3109));
    outputs(3527) <= not(layer0_outputs(2317)) or (layer0_outputs(17));
    outputs(3528) <= not((layer0_outputs(5223)) xor (layer0_outputs(9086)));
    outputs(3529) <= not((layer0_outputs(951)) xor (layer0_outputs(9381)));
    outputs(3530) <= layer0_outputs(10194);
    outputs(3531) <= (layer0_outputs(4524)) and not (layer0_outputs(10121));
    outputs(3532) <= not(layer0_outputs(7187));
    outputs(3533) <= (layer0_outputs(5683)) or (layer0_outputs(3329));
    outputs(3534) <= not(layer0_outputs(472));
    outputs(3535) <= not(layer0_outputs(6372)) or (layer0_outputs(7957));
    outputs(3536) <= not((layer0_outputs(8206)) xor (layer0_outputs(10079)));
    outputs(3537) <= (layer0_outputs(6395)) xor (layer0_outputs(6736));
    outputs(3538) <= layer0_outputs(1456);
    outputs(3539) <= not((layer0_outputs(8943)) or (layer0_outputs(2469)));
    outputs(3540) <= (layer0_outputs(5572)) and not (layer0_outputs(2626));
    outputs(3541) <= not((layer0_outputs(1308)) xor (layer0_outputs(2040)));
    outputs(3542) <= layer0_outputs(276);
    outputs(3543) <= not(layer0_outputs(7366));
    outputs(3544) <= not(layer0_outputs(5173));
    outputs(3545) <= not(layer0_outputs(8351));
    outputs(3546) <= not(layer0_outputs(4487));
    outputs(3547) <= layer0_outputs(6594);
    outputs(3548) <= not((layer0_outputs(6832)) and (layer0_outputs(4946)));
    outputs(3549) <= (layer0_outputs(4684)) or (layer0_outputs(5841));
    outputs(3550) <= (layer0_outputs(3386)) xor (layer0_outputs(1817));
    outputs(3551) <= layer0_outputs(5311);
    outputs(3552) <= not(layer0_outputs(2391)) or (layer0_outputs(8695));
    outputs(3553) <= not((layer0_outputs(7383)) xor (layer0_outputs(3830)));
    outputs(3554) <= not((layer0_outputs(9850)) and (layer0_outputs(6341)));
    outputs(3555) <= layer0_outputs(8564);
    outputs(3556) <= layer0_outputs(3792);
    outputs(3557) <= layer0_outputs(4882);
    outputs(3558) <= (layer0_outputs(9153)) xor (layer0_outputs(9757));
    outputs(3559) <= not((layer0_outputs(234)) and (layer0_outputs(8581)));
    outputs(3560) <= not((layer0_outputs(6519)) and (layer0_outputs(574)));
    outputs(3561) <= layer0_outputs(6767);
    outputs(3562) <= not(layer0_outputs(5174)) or (layer0_outputs(3313));
    outputs(3563) <= (layer0_outputs(2081)) and (layer0_outputs(6729));
    outputs(3564) <= not((layer0_outputs(1066)) xor (layer0_outputs(7957)));
    outputs(3565) <= layer0_outputs(4353);
    outputs(3566) <= not(layer0_outputs(8636));
    outputs(3567) <= not(layer0_outputs(6378));
    outputs(3568) <= not((layer0_outputs(4117)) and (layer0_outputs(2446)));
    outputs(3569) <= (layer0_outputs(9598)) or (layer0_outputs(2024));
    outputs(3570) <= not(layer0_outputs(6543)) or (layer0_outputs(7758));
    outputs(3571) <= (layer0_outputs(8399)) xor (layer0_outputs(2995));
    outputs(3572) <= not(layer0_outputs(2190));
    outputs(3573) <= (layer0_outputs(1517)) or (layer0_outputs(1812));
    outputs(3574) <= layer0_outputs(1108);
    outputs(3575) <= not(layer0_outputs(8929)) or (layer0_outputs(1629));
    outputs(3576) <= (layer0_outputs(6208)) and (layer0_outputs(6463));
    outputs(3577) <= not(layer0_outputs(9385));
    outputs(3578) <= not((layer0_outputs(10066)) xor (layer0_outputs(4765)));
    outputs(3579) <= not((layer0_outputs(9040)) xor (layer0_outputs(1707)));
    outputs(3580) <= (layer0_outputs(6302)) xor (layer0_outputs(8583));
    outputs(3581) <= not(layer0_outputs(5154));
    outputs(3582) <= not(layer0_outputs(4719));
    outputs(3583) <= not(layer0_outputs(5430));
    outputs(3584) <= (layer0_outputs(6465)) xor (layer0_outputs(9296));
    outputs(3585) <= (layer0_outputs(2867)) xor (layer0_outputs(431));
    outputs(3586) <= (layer0_outputs(10125)) xor (layer0_outputs(2919));
    outputs(3587) <= not(layer0_outputs(6227));
    outputs(3588) <= not(layer0_outputs(2051));
    outputs(3589) <= (layer0_outputs(1073)) xor (layer0_outputs(5436));
    outputs(3590) <= (layer0_outputs(3316)) xor (layer0_outputs(3165));
    outputs(3591) <= layer0_outputs(5040);
    outputs(3592) <= (layer0_outputs(4846)) xor (layer0_outputs(2125));
    outputs(3593) <= layer0_outputs(7831);
    outputs(3594) <= not(layer0_outputs(3631)) or (layer0_outputs(5369));
    outputs(3595) <= not((layer0_outputs(2973)) xor (layer0_outputs(9271)));
    outputs(3596) <= (layer0_outputs(568)) or (layer0_outputs(40));
    outputs(3597) <= layer0_outputs(6280);
    outputs(3598) <= not(layer0_outputs(1339));
    outputs(3599) <= not((layer0_outputs(3017)) xor (layer0_outputs(5742)));
    outputs(3600) <= layer0_outputs(6700);
    outputs(3601) <= not(layer0_outputs(9313));
    outputs(3602) <= layer0_outputs(3611);
    outputs(3603) <= not(layer0_outputs(8300));
    outputs(3604) <= (layer0_outputs(7097)) xor (layer0_outputs(1948));
    outputs(3605) <= layer0_outputs(2192);
    outputs(3606) <= (layer0_outputs(6177)) xor (layer0_outputs(7448));
    outputs(3607) <= (layer0_outputs(583)) xor (layer0_outputs(1554));
    outputs(3608) <= not(layer0_outputs(10043));
    outputs(3609) <= not(layer0_outputs(738));
    outputs(3610) <= (layer0_outputs(6448)) xor (layer0_outputs(10229));
    outputs(3611) <= layer0_outputs(6342);
    outputs(3612) <= not(layer0_outputs(9085)) or (layer0_outputs(4537));
    outputs(3613) <= not(layer0_outputs(8444));
    outputs(3614) <= not(layer0_outputs(1228));
    outputs(3615) <= not(layer0_outputs(1358));
    outputs(3616) <= (layer0_outputs(6887)) xor (layer0_outputs(9497));
    outputs(3617) <= not((layer0_outputs(7528)) xor (layer0_outputs(6392)));
    outputs(3618) <= not((layer0_outputs(4482)) xor (layer0_outputs(5385)));
    outputs(3619) <= not(layer0_outputs(4656)) or (layer0_outputs(1784));
    outputs(3620) <= not(layer0_outputs(3283)) or (layer0_outputs(6651));
    outputs(3621) <= layer0_outputs(5572);
    outputs(3622) <= layer0_outputs(10109);
    outputs(3623) <= not(layer0_outputs(9226));
    outputs(3624) <= layer0_outputs(897);
    outputs(3625) <= not(layer0_outputs(14)) or (layer0_outputs(8115));
    outputs(3626) <= (layer0_outputs(3853)) or (layer0_outputs(2418));
    outputs(3627) <= layer0_outputs(9581);
    outputs(3628) <= not((layer0_outputs(1104)) and (layer0_outputs(8829)));
    outputs(3629) <= (layer0_outputs(5164)) xor (layer0_outputs(3415));
    outputs(3630) <= not((layer0_outputs(6133)) and (layer0_outputs(2731)));
    outputs(3631) <= layer0_outputs(7872);
    outputs(3632) <= not(layer0_outputs(1741));
    outputs(3633) <= not(layer0_outputs(10147)) or (layer0_outputs(2980));
    outputs(3634) <= not(layer0_outputs(7424));
    outputs(3635) <= not((layer0_outputs(2253)) xor (layer0_outputs(1498)));
    outputs(3636) <= layer0_outputs(3721);
    outputs(3637) <= (layer0_outputs(254)) xor (layer0_outputs(189));
    outputs(3638) <= (layer0_outputs(6919)) or (layer0_outputs(7621));
    outputs(3639) <= not(layer0_outputs(2720));
    outputs(3640) <= (layer0_outputs(3863)) xor (layer0_outputs(502));
    outputs(3641) <= layer0_outputs(5493);
    outputs(3642) <= not(layer0_outputs(9638));
    outputs(3643) <= not(layer0_outputs(2926));
    outputs(3644) <= layer0_outputs(2881);
    outputs(3645) <= (layer0_outputs(10005)) xor (layer0_outputs(9469));
    outputs(3646) <= not(layer0_outputs(4744));
    outputs(3647) <= not(layer0_outputs(2959)) or (layer0_outputs(6161));
    outputs(3648) <= not(layer0_outputs(10019));
    outputs(3649) <= not((layer0_outputs(10097)) and (layer0_outputs(2810)));
    outputs(3650) <= not((layer0_outputs(4600)) xor (layer0_outputs(1991)));
    outputs(3651) <= not(layer0_outputs(954));
    outputs(3652) <= not((layer0_outputs(5310)) and (layer0_outputs(3459)));
    outputs(3653) <= layer0_outputs(6191);
    outputs(3654) <= (layer0_outputs(233)) xor (layer0_outputs(9224));
    outputs(3655) <= (layer0_outputs(5945)) xor (layer0_outputs(1212));
    outputs(3656) <= layer0_outputs(9764);
    outputs(3657) <= not((layer0_outputs(3065)) xor (layer0_outputs(5865)));
    outputs(3658) <= not((layer0_outputs(7858)) xor (layer0_outputs(4758)));
    outputs(3659) <= not((layer0_outputs(1547)) xor (layer0_outputs(1018)));
    outputs(3660) <= not((layer0_outputs(2641)) xor (layer0_outputs(5602)));
    outputs(3661) <= layer0_outputs(8602);
    outputs(3662) <= not(layer0_outputs(1401));
    outputs(3663) <= layer0_outputs(4906);
    outputs(3664) <= (layer0_outputs(42)) and not (layer0_outputs(2528));
    outputs(3665) <= not(layer0_outputs(2649));
    outputs(3666) <= layer0_outputs(1147);
    outputs(3667) <= layer0_outputs(8113);
    outputs(3668) <= layer0_outputs(9071);
    outputs(3669) <= not(layer0_outputs(5638));
    outputs(3670) <= not(layer0_outputs(5713));
    outputs(3671) <= layer0_outputs(5849);
    outputs(3672) <= not(layer0_outputs(3970));
    outputs(3673) <= layer0_outputs(1324);
    outputs(3674) <= not(layer0_outputs(683)) or (layer0_outputs(6777));
    outputs(3675) <= layer0_outputs(6023);
    outputs(3676) <= not(layer0_outputs(4055)) or (layer0_outputs(8905));
    outputs(3677) <= not((layer0_outputs(561)) xor (layer0_outputs(3634)));
    outputs(3678) <= layer0_outputs(9980);
    outputs(3679) <= (layer0_outputs(8413)) xor (layer0_outputs(5035));
    outputs(3680) <= not(layer0_outputs(7092));
    outputs(3681) <= layer0_outputs(2120);
    outputs(3682) <= layer0_outputs(3890);
    outputs(3683) <= (layer0_outputs(9462)) xor (layer0_outputs(9770));
    outputs(3684) <= (layer0_outputs(4050)) xor (layer0_outputs(4519));
    outputs(3685) <= not(layer0_outputs(7243));
    outputs(3686) <= not(layer0_outputs(9638)) or (layer0_outputs(8330));
    outputs(3687) <= not((layer0_outputs(9328)) xor (layer0_outputs(458)));
    outputs(3688) <= layer0_outputs(8737);
    outputs(3689) <= not(layer0_outputs(9258));
    outputs(3690) <= not(layer0_outputs(4361));
    outputs(3691) <= not(layer0_outputs(5395));
    outputs(3692) <= not(layer0_outputs(7445)) or (layer0_outputs(6426));
    outputs(3693) <= layer0_outputs(1910);
    outputs(3694) <= (layer0_outputs(6829)) and (layer0_outputs(3906));
    outputs(3695) <= not(layer0_outputs(4083)) or (layer0_outputs(10021));
    outputs(3696) <= (layer0_outputs(1387)) xor (layer0_outputs(3083));
    outputs(3697) <= (layer0_outputs(6126)) xor (layer0_outputs(173));
    outputs(3698) <= layer0_outputs(3253);
    outputs(3699) <= layer0_outputs(4227);
    outputs(3700) <= not(layer0_outputs(6775));
    outputs(3701) <= (layer0_outputs(4286)) xor (layer0_outputs(109));
    outputs(3702) <= (layer0_outputs(9813)) and not (layer0_outputs(5692));
    outputs(3703) <= (layer0_outputs(7793)) xor (layer0_outputs(9173));
    outputs(3704) <= not(layer0_outputs(2642));
    outputs(3705) <= not(layer0_outputs(2059));
    outputs(3706) <= (layer0_outputs(2501)) xor (layer0_outputs(1501));
    outputs(3707) <= not((layer0_outputs(2473)) xor (layer0_outputs(2602)));
    outputs(3708) <= not(layer0_outputs(8116));
    outputs(3709) <= (layer0_outputs(7746)) and not (layer0_outputs(3914));
    outputs(3710) <= layer0_outputs(5137);
    outputs(3711) <= not(layer0_outputs(1688)) or (layer0_outputs(3451));
    outputs(3712) <= (layer0_outputs(3366)) xor (layer0_outputs(2230));
    outputs(3713) <= layer0_outputs(2003);
    outputs(3714) <= (layer0_outputs(2730)) xor (layer0_outputs(4220));
    outputs(3715) <= (layer0_outputs(4410)) and not (layer0_outputs(5948));
    outputs(3716) <= (layer0_outputs(9800)) xor (layer0_outputs(4287));
    outputs(3717) <= layer0_outputs(3067);
    outputs(3718) <= not((layer0_outputs(1742)) xor (layer0_outputs(6875)));
    outputs(3719) <= not(layer0_outputs(2144));
    outputs(3720) <= layer0_outputs(5017);
    outputs(3721) <= layer0_outputs(6547);
    outputs(3722) <= not(layer0_outputs(8656));
    outputs(3723) <= not(layer0_outputs(9282));
    outputs(3724) <= '1';
    outputs(3725) <= layer0_outputs(7422);
    outputs(3726) <= not(layer0_outputs(19)) or (layer0_outputs(7030));
    outputs(3727) <= not(layer0_outputs(8228));
    outputs(3728) <= not(layer0_outputs(9449)) or (layer0_outputs(9903));
    outputs(3729) <= not(layer0_outputs(6792)) or (layer0_outputs(4263));
    outputs(3730) <= (layer0_outputs(4876)) xor (layer0_outputs(988));
    outputs(3731) <= (layer0_outputs(8069)) and not (layer0_outputs(1694));
    outputs(3732) <= not((layer0_outputs(3833)) xor (layer0_outputs(9148)));
    outputs(3733) <= not((layer0_outputs(8551)) and (layer0_outputs(8173)));
    outputs(3734) <= layer0_outputs(8899);
    outputs(3735) <= not(layer0_outputs(6027));
    outputs(3736) <= (layer0_outputs(936)) and (layer0_outputs(3969));
    outputs(3737) <= (layer0_outputs(673)) and (layer0_outputs(8133));
    outputs(3738) <= (layer0_outputs(2717)) xor (layer0_outputs(6190));
    outputs(3739) <= not((layer0_outputs(1159)) or (layer0_outputs(10044)));
    outputs(3740) <= (layer0_outputs(7712)) xor (layer0_outputs(2688));
    outputs(3741) <= (layer0_outputs(4457)) xor (layer0_outputs(2708));
    outputs(3742) <= layer0_outputs(369);
    outputs(3743) <= not((layer0_outputs(1139)) xor (layer0_outputs(7280)));
    outputs(3744) <= layer0_outputs(6405);
    outputs(3745) <= (layer0_outputs(8557)) xor (layer0_outputs(7365));
    outputs(3746) <= not((layer0_outputs(1369)) xor (layer0_outputs(817)));
    outputs(3747) <= (layer0_outputs(6614)) xor (layer0_outputs(244));
    outputs(3748) <= not((layer0_outputs(2626)) and (layer0_outputs(7734)));
    outputs(3749) <= not((layer0_outputs(2357)) xor (layer0_outputs(5816)));
    outputs(3750) <= not(layer0_outputs(10223)) or (layer0_outputs(8438));
    outputs(3751) <= (layer0_outputs(7394)) xor (layer0_outputs(5798));
    outputs(3752) <= layer0_outputs(4515);
    outputs(3753) <= not(layer0_outputs(883));
    outputs(3754) <= not((layer0_outputs(8473)) xor (layer0_outputs(2612)));
    outputs(3755) <= not((layer0_outputs(1716)) xor (layer0_outputs(4818)));
    outputs(3756) <= not(layer0_outputs(769));
    outputs(3757) <= not((layer0_outputs(7950)) or (layer0_outputs(5847)));
    outputs(3758) <= (layer0_outputs(5636)) xor (layer0_outputs(4993));
    outputs(3759) <= not(layer0_outputs(719)) or (layer0_outputs(2141));
    outputs(3760) <= (layer0_outputs(8174)) or (layer0_outputs(8038));
    outputs(3761) <= layer0_outputs(7261);
    outputs(3762) <= not((layer0_outputs(3246)) xor (layer0_outputs(8035)));
    outputs(3763) <= not((layer0_outputs(7529)) xor (layer0_outputs(1716)));
    outputs(3764) <= not((layer0_outputs(5985)) xor (layer0_outputs(5393)));
    outputs(3765) <= not((layer0_outputs(9096)) xor (layer0_outputs(4122)));
    outputs(3766) <= not(layer0_outputs(7559));
    outputs(3767) <= layer0_outputs(4807);
    outputs(3768) <= not(layer0_outputs(9076)) or (layer0_outputs(6548));
    outputs(3769) <= layer0_outputs(3817);
    outputs(3770) <= (layer0_outputs(2471)) xor (layer0_outputs(9122));
    outputs(3771) <= (layer0_outputs(1836)) xor (layer0_outputs(9289));
    outputs(3772) <= layer0_outputs(454);
    outputs(3773) <= not((layer0_outputs(9953)) xor (layer0_outputs(3139)));
    outputs(3774) <= (layer0_outputs(480)) xor (layer0_outputs(4649));
    outputs(3775) <= not((layer0_outputs(2300)) xor (layer0_outputs(2922)));
    outputs(3776) <= (layer0_outputs(1743)) and (layer0_outputs(3967));
    outputs(3777) <= (layer0_outputs(9696)) or (layer0_outputs(4693));
    outputs(3778) <= (layer0_outputs(6035)) or (layer0_outputs(2685));
    outputs(3779) <= layer0_outputs(996);
    outputs(3780) <= layer0_outputs(5962);
    outputs(3781) <= layer0_outputs(8301);
    outputs(3782) <= not((layer0_outputs(4765)) xor (layer0_outputs(7400)));
    outputs(3783) <= not((layer0_outputs(2512)) or (layer0_outputs(2364)));
    outputs(3784) <= not(layer0_outputs(274));
    outputs(3785) <= not(layer0_outputs(320));
    outputs(3786) <= (layer0_outputs(9031)) and not (layer0_outputs(2890));
    outputs(3787) <= layer0_outputs(3234);
    outputs(3788) <= (layer0_outputs(550)) xor (layer0_outputs(4406));
    outputs(3789) <= not(layer0_outputs(3928)) or (layer0_outputs(3356));
    outputs(3790) <= layer0_outputs(4113);
    outputs(3791) <= layer0_outputs(6430);
    outputs(3792) <= layer0_outputs(9182);
    outputs(3793) <= not((layer0_outputs(4522)) and (layer0_outputs(1355)));
    outputs(3794) <= layer0_outputs(983);
    outputs(3795) <= not(layer0_outputs(3532)) or (layer0_outputs(9899));
    outputs(3796) <= (layer0_outputs(3110)) and not (layer0_outputs(822));
    outputs(3797) <= not(layer0_outputs(10163)) or (layer0_outputs(8572));
    outputs(3798) <= layer0_outputs(8339);
    outputs(3799) <= layer0_outputs(9450);
    outputs(3800) <= (layer0_outputs(3865)) xor (layer0_outputs(952));
    outputs(3801) <= layer0_outputs(9046);
    outputs(3802) <= not(layer0_outputs(10155));
    outputs(3803) <= not((layer0_outputs(3891)) xor (layer0_outputs(8964)));
    outputs(3804) <= layer0_outputs(3140);
    outputs(3805) <= layer0_outputs(9351);
    outputs(3806) <= layer0_outputs(9188);
    outputs(3807) <= not((layer0_outputs(6783)) xor (layer0_outputs(5099)));
    outputs(3808) <= (layer0_outputs(573)) and not (layer0_outputs(4312));
    outputs(3809) <= (layer0_outputs(3893)) xor (layer0_outputs(5749));
    outputs(3810) <= (layer0_outputs(2420)) xor (layer0_outputs(645));
    outputs(3811) <= layer0_outputs(5018);
    outputs(3812) <= not((layer0_outputs(6866)) xor (layer0_outputs(6552)));
    outputs(3813) <= not(layer0_outputs(6060));
    outputs(3814) <= layer0_outputs(3);
    outputs(3815) <= (layer0_outputs(8545)) and not (layer0_outputs(4409));
    outputs(3816) <= not(layer0_outputs(9881));
    outputs(3817) <= not((layer0_outputs(2904)) and (layer0_outputs(2219)));
    outputs(3818) <= not(layer0_outputs(8452));
    outputs(3819) <= not((layer0_outputs(6293)) xor (layer0_outputs(6412)));
    outputs(3820) <= not((layer0_outputs(2151)) or (layer0_outputs(284)));
    outputs(3821) <= (layer0_outputs(7391)) and not (layer0_outputs(5094));
    outputs(3822) <= (layer0_outputs(3603)) xor (layer0_outputs(9303));
    outputs(3823) <= not((layer0_outputs(424)) xor (layer0_outputs(656)));
    outputs(3824) <= (layer0_outputs(7582)) and not (layer0_outputs(9929));
    outputs(3825) <= not(layer0_outputs(4316));
    outputs(3826) <= not(layer0_outputs(2279));
    outputs(3827) <= (layer0_outputs(7540)) xor (layer0_outputs(10051));
    outputs(3828) <= layer0_outputs(7030);
    outputs(3829) <= (layer0_outputs(8624)) and not (layer0_outputs(7107));
    outputs(3830) <= layer0_outputs(861);
    outputs(3831) <= layer0_outputs(7835);
    outputs(3832) <= (layer0_outputs(164)) xor (layer0_outputs(2457));
    outputs(3833) <= (layer0_outputs(9584)) xor (layer0_outputs(1080));
    outputs(3834) <= not(layer0_outputs(2472));
    outputs(3835) <= (layer0_outputs(8017)) xor (layer0_outputs(277));
    outputs(3836) <= not(layer0_outputs(7308));
    outputs(3837) <= layer0_outputs(8106);
    outputs(3838) <= not(layer0_outputs(10038));
    outputs(3839) <= layer0_outputs(9350);
    outputs(3840) <= (layer0_outputs(6500)) xor (layer0_outputs(2841));
    outputs(3841) <= layer0_outputs(1144);
    outputs(3842) <= not(layer0_outputs(2390));
    outputs(3843) <= (layer0_outputs(8680)) xor (layer0_outputs(3875));
    outputs(3844) <= (layer0_outputs(7293)) and not (layer0_outputs(7105));
    outputs(3845) <= layer0_outputs(8096);
    outputs(3846) <= not(layer0_outputs(1385)) or (layer0_outputs(3554));
    outputs(3847) <= not((layer0_outputs(9777)) and (layer0_outputs(906)));
    outputs(3848) <= not((layer0_outputs(571)) and (layer0_outputs(1749)));
    outputs(3849) <= not((layer0_outputs(7586)) xor (layer0_outputs(8317)));
    outputs(3850) <= layer0_outputs(8079);
    outputs(3851) <= not(layer0_outputs(7326));
    outputs(3852) <= not(layer0_outputs(1268));
    outputs(3853) <= not(layer0_outputs(5472)) or (layer0_outputs(3001));
    outputs(3854) <= not(layer0_outputs(3341)) or (layer0_outputs(3432));
    outputs(3855) <= not(layer0_outputs(2955));
    outputs(3856) <= not(layer0_outputs(1080)) or (layer0_outputs(3039));
    outputs(3857) <= not(layer0_outputs(7369)) or (layer0_outputs(8257));
    outputs(3858) <= not(layer0_outputs(10192));
    outputs(3859) <= (layer0_outputs(2369)) and not (layer0_outputs(7172));
    outputs(3860) <= not(layer0_outputs(9791));
    outputs(3861) <= (layer0_outputs(5748)) and not (layer0_outputs(7821));
    outputs(3862) <= not(layer0_outputs(5771));
    outputs(3863) <= not((layer0_outputs(1586)) or (layer0_outputs(33)));
    outputs(3864) <= layer0_outputs(6367);
    outputs(3865) <= layer0_outputs(4413);
    outputs(3866) <= (layer0_outputs(6857)) or (layer0_outputs(3648));
    outputs(3867) <= (layer0_outputs(6625)) xor (layer0_outputs(3881));
    outputs(3868) <= not((layer0_outputs(8391)) xor (layer0_outputs(311)));
    outputs(3869) <= (layer0_outputs(4249)) xor (layer0_outputs(202));
    outputs(3870) <= not(layer0_outputs(3507));
    outputs(3871) <= not(layer0_outputs(361));
    outputs(3872) <= not(layer0_outputs(9421));
    outputs(3873) <= not(layer0_outputs(3000));
    outputs(3874) <= layer0_outputs(2703);
    outputs(3875) <= not(layer0_outputs(2548)) or (layer0_outputs(1541));
    outputs(3876) <= '1';
    outputs(3877) <= (layer0_outputs(3555)) and (layer0_outputs(2985));
    outputs(3878) <= not(layer0_outputs(9127)) or (layer0_outputs(1362));
    outputs(3879) <= not(layer0_outputs(8078));
    outputs(3880) <= layer0_outputs(7909);
    outputs(3881) <= not(layer0_outputs(9187));
    outputs(3882) <= not(layer0_outputs(6432));
    outputs(3883) <= not(layer0_outputs(7093)) or (layer0_outputs(1712));
    outputs(3884) <= not(layer0_outputs(1497));
    outputs(3885) <= not((layer0_outputs(8867)) xor (layer0_outputs(2375)));
    outputs(3886) <= not((layer0_outputs(8367)) xor (layer0_outputs(7101)));
    outputs(3887) <= (layer0_outputs(8664)) or (layer0_outputs(8941));
    outputs(3888) <= not(layer0_outputs(7729));
    outputs(3889) <= not(layer0_outputs(2461)) or (layer0_outputs(7504));
    outputs(3890) <= not(layer0_outputs(6628)) or (layer0_outputs(2358));
    outputs(3891) <= layer0_outputs(2854);
    outputs(3892) <= (layer0_outputs(7287)) and (layer0_outputs(4592));
    outputs(3893) <= layer0_outputs(6762);
    outputs(3894) <= layer0_outputs(7811);
    outputs(3895) <= not(layer0_outputs(7923));
    outputs(3896) <= not(layer0_outputs(6418));
    outputs(3897) <= (layer0_outputs(3604)) and not (layer0_outputs(7906));
    outputs(3898) <= layer0_outputs(5925);
    outputs(3899) <= (layer0_outputs(6179)) xor (layer0_outputs(9632));
    outputs(3900) <= not((layer0_outputs(2551)) xor (layer0_outputs(5198)));
    outputs(3901) <= not(layer0_outputs(9975));
    outputs(3902) <= not(layer0_outputs(1252));
    outputs(3903) <= layer0_outputs(6269);
    outputs(3904) <= not((layer0_outputs(3305)) xor (layer0_outputs(4824)));
    outputs(3905) <= (layer0_outputs(6773)) xor (layer0_outputs(1949));
    outputs(3906) <= not(layer0_outputs(2373));
    outputs(3907) <= layer0_outputs(2753);
    outputs(3908) <= not(layer0_outputs(6578)) or (layer0_outputs(6840));
    outputs(3909) <= layer0_outputs(2426);
    outputs(3910) <= not(layer0_outputs(9817)) or (layer0_outputs(2791));
    outputs(3911) <= not(layer0_outputs(3124));
    outputs(3912) <= not((layer0_outputs(9546)) xor (layer0_outputs(5755)));
    outputs(3913) <= (layer0_outputs(8508)) xor (layer0_outputs(9582));
    outputs(3914) <= (layer0_outputs(4448)) or (layer0_outputs(8840));
    outputs(3915) <= not(layer0_outputs(1876));
    outputs(3916) <= not((layer0_outputs(5426)) xor (layer0_outputs(7983)));
    outputs(3917) <= layer0_outputs(9958);
    outputs(3918) <= not(layer0_outputs(2365)) or (layer0_outputs(7247));
    outputs(3919) <= not(layer0_outputs(4021));
    outputs(3920) <= layer0_outputs(2511);
    outputs(3921) <= not(layer0_outputs(4883));
    outputs(3922) <= (layer0_outputs(1318)) xor (layer0_outputs(6903));
    outputs(3923) <= not(layer0_outputs(4455));
    outputs(3924) <= (layer0_outputs(4699)) or (layer0_outputs(10103));
    outputs(3925) <= layer0_outputs(388);
    outputs(3926) <= not((layer0_outputs(3175)) xor (layer0_outputs(10105)));
    outputs(3927) <= not(layer0_outputs(9257)) or (layer0_outputs(1813));
    outputs(3928) <= not((layer0_outputs(7490)) or (layer0_outputs(1367)));
    outputs(3929) <= (layer0_outputs(373)) and not (layer0_outputs(6871));
    outputs(3930) <= (layer0_outputs(8014)) and not (layer0_outputs(1398));
    outputs(3931) <= not((layer0_outputs(9782)) or (layer0_outputs(6075)));
    outputs(3932) <= layer0_outputs(7988);
    outputs(3933) <= layer0_outputs(8185);
    outputs(3934) <= (layer0_outputs(1702)) or (layer0_outputs(8183));
    outputs(3935) <= not(layer0_outputs(9140));
    outputs(3936) <= not(layer0_outputs(7514));
    outputs(3937) <= '1';
    outputs(3938) <= layer0_outputs(8639);
    outputs(3939) <= not(layer0_outputs(364));
    outputs(3940) <= (layer0_outputs(9041)) and not (layer0_outputs(9594));
    outputs(3941) <= layer0_outputs(1284);
    outputs(3942) <= not(layer0_outputs(7111));
    outputs(3943) <= not(layer0_outputs(5515));
    outputs(3944) <= not(layer0_outputs(7556)) or (layer0_outputs(9111));
    outputs(3945) <= not(layer0_outputs(2825));
    outputs(3946) <= not((layer0_outputs(4253)) xor (layer0_outputs(7725)));
    outputs(3947) <= not(layer0_outputs(8789));
    outputs(3948) <= not(layer0_outputs(3065));
    outputs(3949) <= (layer0_outputs(7568)) or (layer0_outputs(3888));
    outputs(3950) <= not((layer0_outputs(5142)) and (layer0_outputs(5466)));
    outputs(3951) <= not(layer0_outputs(16)) or (layer0_outputs(8226));
    outputs(3952) <= not((layer0_outputs(5122)) or (layer0_outputs(1253)));
    outputs(3953) <= not(layer0_outputs(3944));
    outputs(3954) <= not(layer0_outputs(9043));
    outputs(3955) <= not((layer0_outputs(2180)) xor (layer0_outputs(9481)));
    outputs(3956) <= not(layer0_outputs(285)) or (layer0_outputs(7498));
    outputs(3957) <= layer0_outputs(6895);
    outputs(3958) <= not((layer0_outputs(5983)) xor (layer0_outputs(166)));
    outputs(3959) <= (layer0_outputs(5871)) and not (layer0_outputs(5948));
    outputs(3960) <= not((layer0_outputs(9986)) xor (layer0_outputs(4166)));
    outputs(3961) <= not((layer0_outputs(8136)) xor (layer0_outputs(2966)));
    outputs(3962) <= not(layer0_outputs(4787));
    outputs(3963) <= (layer0_outputs(5943)) xor (layer0_outputs(2768));
    outputs(3964) <= not((layer0_outputs(3904)) xor (layer0_outputs(561)));
    outputs(3965) <= layer0_outputs(6289);
    outputs(3966) <= layer0_outputs(5633);
    outputs(3967) <= not(layer0_outputs(7408));
    outputs(3968) <= (layer0_outputs(9211)) and (layer0_outputs(6987));
    outputs(3969) <= layer0_outputs(668);
    outputs(3970) <= not(layer0_outputs(2834));
    outputs(3971) <= not(layer0_outputs(757)) or (layer0_outputs(7538));
    outputs(3972) <= (layer0_outputs(4073)) xor (layer0_outputs(3375));
    outputs(3973) <= not(layer0_outputs(6096));
    outputs(3974) <= (layer0_outputs(2897)) xor (layer0_outputs(2288));
    outputs(3975) <= layer0_outputs(6082);
    outputs(3976) <= not(layer0_outputs(8827));
    outputs(3977) <= layer0_outputs(2465);
    outputs(3978) <= layer0_outputs(6547);
    outputs(3979) <= (layer0_outputs(1263)) xor (layer0_outputs(7993));
    outputs(3980) <= layer0_outputs(5212);
    outputs(3981) <= not(layer0_outputs(5145));
    outputs(3982) <= not(layer0_outputs(4923));
    outputs(3983) <= (layer0_outputs(3537)) or (layer0_outputs(605));
    outputs(3984) <= not(layer0_outputs(9877));
    outputs(3985) <= not(layer0_outputs(5991)) or (layer0_outputs(6692));
    outputs(3986) <= (layer0_outputs(5898)) xor (layer0_outputs(3865));
    outputs(3987) <= '1';
    outputs(3988) <= not(layer0_outputs(9215));
    outputs(3989) <= (layer0_outputs(8912)) xor (layer0_outputs(1457));
    outputs(3990) <= (layer0_outputs(2703)) and (layer0_outputs(7512));
    outputs(3991) <= not(layer0_outputs(4801));
    outputs(3992) <= layer0_outputs(3651);
    outputs(3993) <= not((layer0_outputs(290)) xor (layer0_outputs(3350)));
    outputs(3994) <= layer0_outputs(4950);
    outputs(3995) <= not(layer0_outputs(6181));
    outputs(3996) <= (layer0_outputs(8256)) xor (layer0_outputs(7500));
    outputs(3997) <= not(layer0_outputs(4278)) or (layer0_outputs(5181));
    outputs(3998) <= (layer0_outputs(6764)) xor (layer0_outputs(811));
    outputs(3999) <= (layer0_outputs(4004)) and (layer0_outputs(6801));
    outputs(4000) <= (layer0_outputs(2447)) xor (layer0_outputs(2348));
    outputs(4001) <= layer0_outputs(1273);
    outputs(4002) <= not(layer0_outputs(2780));
    outputs(4003) <= not(layer0_outputs(8570)) or (layer0_outputs(5849));
    outputs(4004) <= not((layer0_outputs(3330)) or (layer0_outputs(6710)));
    outputs(4005) <= (layer0_outputs(10108)) and not (layer0_outputs(3448));
    outputs(4006) <= (layer0_outputs(8768)) xor (layer0_outputs(10125));
    outputs(4007) <= (layer0_outputs(1372)) xor (layer0_outputs(771));
    outputs(4008) <= not((layer0_outputs(1789)) and (layer0_outputs(7667)));
    outputs(4009) <= (layer0_outputs(2584)) xor (layer0_outputs(7542));
    outputs(4010) <= layer0_outputs(358);
    outputs(4011) <= not(layer0_outputs(2663)) or (layer0_outputs(4846));
    outputs(4012) <= not((layer0_outputs(2883)) xor (layer0_outputs(2001)));
    outputs(4013) <= not(layer0_outputs(7685));
    outputs(4014) <= not(layer0_outputs(529));
    outputs(4015) <= not(layer0_outputs(4399));
    outputs(4016) <= (layer0_outputs(5282)) xor (layer0_outputs(5263));
    outputs(4017) <= layer0_outputs(8590);
    outputs(4018) <= layer0_outputs(2979);
    outputs(4019) <= (layer0_outputs(5827)) xor (layer0_outputs(5710));
    outputs(4020) <= not(layer0_outputs(11)) or (layer0_outputs(4681));
    outputs(4021) <= not(layer0_outputs(10155));
    outputs(4022) <= (layer0_outputs(2104)) or (layer0_outputs(6607));
    outputs(4023) <= not((layer0_outputs(7433)) and (layer0_outputs(3534)));
    outputs(4024) <= layer0_outputs(4335);
    outputs(4025) <= '0';
    outputs(4026) <= layer0_outputs(724);
    outputs(4027) <= (layer0_outputs(8888)) and not (layer0_outputs(9227));
    outputs(4028) <= not((layer0_outputs(5421)) xor (layer0_outputs(2297)));
    outputs(4029) <= not(layer0_outputs(7730));
    outputs(4030) <= (layer0_outputs(6558)) xor (layer0_outputs(6689));
    outputs(4031) <= not(layer0_outputs(3136)) or (layer0_outputs(4407));
    outputs(4032) <= not((layer0_outputs(8092)) xor (layer0_outputs(3364)));
    outputs(4033) <= (layer0_outputs(129)) and not (layer0_outputs(8416));
    outputs(4034) <= not(layer0_outputs(779)) or (layer0_outputs(6749));
    outputs(4035) <= layer0_outputs(7819);
    outputs(4036) <= layer0_outputs(4367);
    outputs(4037) <= not((layer0_outputs(1506)) and (layer0_outputs(6265)));
    outputs(4038) <= not((layer0_outputs(2705)) xor (layer0_outputs(8890)));
    outputs(4039) <= layer0_outputs(9430);
    outputs(4040) <= (layer0_outputs(2396)) or (layer0_outputs(9495));
    outputs(4041) <= layer0_outputs(370);
    outputs(4042) <= (layer0_outputs(3258)) and (layer0_outputs(794));
    outputs(4043) <= not(layer0_outputs(4971)) or (layer0_outputs(6490));
    outputs(4044) <= not((layer0_outputs(376)) or (layer0_outputs(10078)));
    outputs(4045) <= not(layer0_outputs(691));
    outputs(4046) <= not(layer0_outputs(860));
    outputs(4047) <= layer0_outputs(10227);
    outputs(4048) <= not(layer0_outputs(3663)) or (layer0_outputs(5530));
    outputs(4049) <= (layer0_outputs(1903)) and not (layer0_outputs(4647));
    outputs(4050) <= not(layer0_outputs(10134));
    outputs(4051) <= not((layer0_outputs(6772)) or (layer0_outputs(10082)));
    outputs(4052) <= (layer0_outputs(2054)) and (layer0_outputs(2385));
    outputs(4053) <= layer0_outputs(9416);
    outputs(4054) <= (layer0_outputs(119)) xor (layer0_outputs(10108));
    outputs(4055) <= (layer0_outputs(8139)) xor (layer0_outputs(2226));
    outputs(4056) <= not(layer0_outputs(8116));
    outputs(4057) <= not((layer0_outputs(4905)) xor (layer0_outputs(9780)));
    outputs(4058) <= not(layer0_outputs(9778)) or (layer0_outputs(6537));
    outputs(4059) <= (layer0_outputs(2400)) xor (layer0_outputs(5093));
    outputs(4060) <= layer0_outputs(7791);
    outputs(4061) <= layer0_outputs(7748);
    outputs(4062) <= not(layer0_outputs(7078)) or (layer0_outputs(1866));
    outputs(4063) <= (layer0_outputs(6921)) or (layer0_outputs(4175));
    outputs(4064) <= not(layer0_outputs(5697)) or (layer0_outputs(3476));
    outputs(4065) <= (layer0_outputs(8329)) or (layer0_outputs(3949));
    outputs(4066) <= not(layer0_outputs(8901)) or (layer0_outputs(8670));
    outputs(4067) <= not((layer0_outputs(3665)) and (layer0_outputs(2640)));
    outputs(4068) <= layer0_outputs(2595);
    outputs(4069) <= not(layer0_outputs(7490));
    outputs(4070) <= not((layer0_outputs(4651)) xor (layer0_outputs(2765)));
    outputs(4071) <= (layer0_outputs(8966)) xor (layer0_outputs(2543));
    outputs(4072) <= (layer0_outputs(8778)) xor (layer0_outputs(3700));
    outputs(4073) <= (layer0_outputs(7253)) xor (layer0_outputs(5685));
    outputs(4074) <= (layer0_outputs(6010)) and not (layer0_outputs(10164));
    outputs(4075) <= not(layer0_outputs(2438)) or (layer0_outputs(3423));
    outputs(4076) <= layer0_outputs(4572);
    outputs(4077) <= layer0_outputs(2590);
    outputs(4078) <= not(layer0_outputs(10045)) or (layer0_outputs(4168));
    outputs(4079) <= not((layer0_outputs(2592)) and (layer0_outputs(2209)));
    outputs(4080) <= layer0_outputs(8942);
    outputs(4081) <= layer0_outputs(8746);
    outputs(4082) <= not(layer0_outputs(2566));
    outputs(4083) <= not(layer0_outputs(3207));
    outputs(4084) <= not((layer0_outputs(7285)) xor (layer0_outputs(1012)));
    outputs(4085) <= layer0_outputs(9196);
    outputs(4086) <= (layer0_outputs(1591)) or (layer0_outputs(4024));
    outputs(4087) <= layer0_outputs(3581);
    outputs(4088) <= (layer0_outputs(7141)) xor (layer0_outputs(7912));
    outputs(4089) <= not(layer0_outputs(286));
    outputs(4090) <= not((layer0_outputs(9046)) and (layer0_outputs(39)));
    outputs(4091) <= not(layer0_outputs(4881));
    outputs(4092) <= not(layer0_outputs(57)) or (layer0_outputs(6480));
    outputs(4093) <= (layer0_outputs(8338)) xor (layer0_outputs(5419));
    outputs(4094) <= not((layer0_outputs(9291)) xor (layer0_outputs(9827)));
    outputs(4095) <= (layer0_outputs(3808)) and not (layer0_outputs(1316));
    outputs(4096) <= not((layer0_outputs(2867)) or (layer0_outputs(3353)));
    outputs(4097) <= layer0_outputs(935);
    outputs(4098) <= (layer0_outputs(9585)) and not (layer0_outputs(9431));
    outputs(4099) <= (layer0_outputs(6216)) and not (layer0_outputs(4975));
    outputs(4100) <= not((layer0_outputs(6394)) xor (layer0_outputs(8099)));
    outputs(4101) <= layer0_outputs(7902);
    outputs(4102) <= not(layer0_outputs(1338)) or (layer0_outputs(7690));
    outputs(4103) <= not((layer0_outputs(3756)) xor (layer0_outputs(9687)));
    outputs(4104) <= (layer0_outputs(5401)) xor (layer0_outputs(5054));
    outputs(4105) <= not(layer0_outputs(4294));
    outputs(4106) <= (layer0_outputs(1384)) and (layer0_outputs(4740));
    outputs(4107) <= (layer0_outputs(3450)) and not (layer0_outputs(164));
    outputs(4108) <= not((layer0_outputs(5721)) or (layer0_outputs(7919)));
    outputs(4109) <= not(layer0_outputs(3923));
    outputs(4110) <= not((layer0_outputs(7703)) or (layer0_outputs(8308)));
    outputs(4111) <= layer0_outputs(5917);
    outputs(4112) <= not((layer0_outputs(2861)) and (layer0_outputs(1628)));
    outputs(4113) <= layer0_outputs(1876);
    outputs(4114) <= (layer0_outputs(6953)) and (layer0_outputs(2664));
    outputs(4115) <= (layer0_outputs(7663)) xor (layer0_outputs(4218));
    outputs(4116) <= (layer0_outputs(6668)) and not (layer0_outputs(1317));
    outputs(4117) <= (layer0_outputs(3321)) xor (layer0_outputs(3378));
    outputs(4118) <= not(layer0_outputs(2486));
    outputs(4119) <= (layer0_outputs(2445)) and not (layer0_outputs(1517));
    outputs(4120) <= not(layer0_outputs(2907));
    outputs(4121) <= not(layer0_outputs(5431));
    outputs(4122) <= (layer0_outputs(7332)) xor (layer0_outputs(1377));
    outputs(4123) <= not((layer0_outputs(1392)) xor (layer0_outputs(1729)));
    outputs(4124) <= (layer0_outputs(6505)) and not (layer0_outputs(4791));
    outputs(4125) <= not((layer0_outputs(7827)) and (layer0_outputs(3935)));
    outputs(4126) <= (layer0_outputs(2069)) and not (layer0_outputs(6176));
    outputs(4127) <= not(layer0_outputs(7060));
    outputs(4128) <= layer0_outputs(8772);
    outputs(4129) <= not(layer0_outputs(7306));
    outputs(4130) <= not((layer0_outputs(5935)) xor (layer0_outputs(5324)));
    outputs(4131) <= not((layer0_outputs(2233)) or (layer0_outputs(3036)));
    outputs(4132) <= layer0_outputs(5397);
    outputs(4133) <= (layer0_outputs(4390)) xor (layer0_outputs(3652));
    outputs(4134) <= not(layer0_outputs(8045));
    outputs(4135) <= not((layer0_outputs(9034)) and (layer0_outputs(9696)));
    outputs(4136) <= (layer0_outputs(7992)) xor (layer0_outputs(3655));
    outputs(4137) <= not((layer0_outputs(8682)) xor (layer0_outputs(5878)));
    outputs(4138) <= not((layer0_outputs(2466)) or (layer0_outputs(5772)));
    outputs(4139) <= layer0_outputs(1258);
    outputs(4140) <= layer0_outputs(8590);
    outputs(4141) <= not((layer0_outputs(4903)) xor (layer0_outputs(6140)));
    outputs(4142) <= not(layer0_outputs(2052));
    outputs(4143) <= not((layer0_outputs(2301)) xor (layer0_outputs(5550)));
    outputs(4144) <= (layer0_outputs(4325)) and not (layer0_outputs(237));
    outputs(4145) <= not((layer0_outputs(347)) xor (layer0_outputs(9721)));
    outputs(4146) <= not(layer0_outputs(8879));
    outputs(4147) <= (layer0_outputs(3129)) and (layer0_outputs(274));
    outputs(4148) <= layer0_outputs(8242);
    outputs(4149) <= not(layer0_outputs(3781));
    outputs(4150) <= not(layer0_outputs(4223)) or (layer0_outputs(8679));
    outputs(4151) <= not(layer0_outputs(4036));
    outputs(4152) <= layer0_outputs(1186);
    outputs(4153) <= (layer0_outputs(8796)) xor (layer0_outputs(1649));
    outputs(4154) <= layer0_outputs(5846);
    outputs(4155) <= layer0_outputs(1438);
    outputs(4156) <= not(layer0_outputs(7793));
    outputs(4157) <= (layer0_outputs(7075)) and not (layer0_outputs(6037));
    outputs(4158) <= not(layer0_outputs(9650));
    outputs(4159) <= layer0_outputs(2525);
    outputs(4160) <= layer0_outputs(319);
    outputs(4161) <= not((layer0_outputs(6871)) or (layer0_outputs(7879)));
    outputs(4162) <= (layer0_outputs(3155)) xor (layer0_outputs(2120));
    outputs(4163) <= not(layer0_outputs(6238));
    outputs(4164) <= not(layer0_outputs(8108));
    outputs(4165) <= (layer0_outputs(3324)) and (layer0_outputs(6657));
    outputs(4166) <= not(layer0_outputs(404));
    outputs(4167) <= not((layer0_outputs(7878)) or (layer0_outputs(6767)));
    outputs(4168) <= (layer0_outputs(895)) and not (layer0_outputs(7857));
    outputs(4169) <= layer0_outputs(4857);
    outputs(4170) <= (layer0_outputs(146)) and not (layer0_outputs(9800));
    outputs(4171) <= (layer0_outputs(2839)) and not (layer0_outputs(4334));
    outputs(4172) <= not((layer0_outputs(1485)) xor (layer0_outputs(9122)));
    outputs(4173) <= layer0_outputs(10110);
    outputs(4174) <= (layer0_outputs(5304)) xor (layer0_outputs(972));
    outputs(4175) <= not(layer0_outputs(3346));
    outputs(4176) <= layer0_outputs(8385);
    outputs(4177) <= (layer0_outputs(9239)) and not (layer0_outputs(8095));
    outputs(4178) <= (layer0_outputs(5349)) and not (layer0_outputs(2932));
    outputs(4179) <= not(layer0_outputs(4578));
    outputs(4180) <= not(layer0_outputs(4392)) or (layer0_outputs(9686));
    outputs(4181) <= layer0_outputs(2302);
    outputs(4182) <= (layer0_outputs(8786)) and not (layer0_outputs(9979));
    outputs(4183) <= not(layer0_outputs(7290));
    outputs(4184) <= not(layer0_outputs(6702));
    outputs(4185) <= (layer0_outputs(3469)) xor (layer0_outputs(8916));
    outputs(4186) <= not(layer0_outputs(7290)) or (layer0_outputs(9938));
    outputs(4187) <= not((layer0_outputs(10203)) or (layer0_outputs(8275)));
    outputs(4188) <= not((layer0_outputs(9010)) or (layer0_outputs(10071)));
    outputs(4189) <= (layer0_outputs(5109)) xor (layer0_outputs(5881));
    outputs(4190) <= (layer0_outputs(6533)) and not (layer0_outputs(4526));
    outputs(4191) <= not(layer0_outputs(7221));
    outputs(4192) <= layer0_outputs(5345);
    outputs(4193) <= not((layer0_outputs(6149)) xor (layer0_outputs(3496)));
    outputs(4194) <= (layer0_outputs(5938)) xor (layer0_outputs(2715));
    outputs(4195) <= layer0_outputs(4003);
    outputs(4196) <= not((layer0_outputs(3426)) xor (layer0_outputs(8221)));
    outputs(4197) <= layer0_outputs(1368);
    outputs(4198) <= not(layer0_outputs(5167));
    outputs(4199) <= layer0_outputs(5515);
    outputs(4200) <= not((layer0_outputs(4298)) xor (layer0_outputs(4047)));
    outputs(4201) <= (layer0_outputs(2259)) and not (layer0_outputs(4121));
    outputs(4202) <= not(layer0_outputs(116));
    outputs(4203) <= (layer0_outputs(1496)) and not (layer0_outputs(9002));
    outputs(4204) <= layer0_outputs(3834);
    outputs(4205) <= not(layer0_outputs(10041));
    outputs(4206) <= not((layer0_outputs(10074)) and (layer0_outputs(8209)));
    outputs(4207) <= not(layer0_outputs(7841)) or (layer0_outputs(8763));
    outputs(4208) <= layer0_outputs(10166);
    outputs(4209) <= (layer0_outputs(3407)) and (layer0_outputs(506));
    outputs(4210) <= (layer0_outputs(1500)) xor (layer0_outputs(9668));
    outputs(4211) <= (layer0_outputs(7873)) and not (layer0_outputs(7948));
    outputs(4212) <= not((layer0_outputs(7244)) xor (layer0_outputs(6924)));
    outputs(4213) <= layer0_outputs(1785);
    outputs(4214) <= not(layer0_outputs(4082)) or (layer0_outputs(3457));
    outputs(4215) <= (layer0_outputs(4348)) and (layer0_outputs(3219));
    outputs(4216) <= (layer0_outputs(4612)) and not (layer0_outputs(6639));
    outputs(4217) <= (layer0_outputs(8930)) xor (layer0_outputs(5036));
    outputs(4218) <= not(layer0_outputs(3262));
    outputs(4219) <= not((layer0_outputs(2585)) or (layer0_outputs(8862)));
    outputs(4220) <= (layer0_outputs(10098)) and not (layer0_outputs(590));
    outputs(4221) <= not((layer0_outputs(1495)) xor (layer0_outputs(1504)));
    outputs(4222) <= not((layer0_outputs(4434)) or (layer0_outputs(2750)));
    outputs(4223) <= (layer0_outputs(808)) xor (layer0_outputs(8584));
    outputs(4224) <= layer0_outputs(1934);
    outputs(4225) <= (layer0_outputs(7847)) and not (layer0_outputs(6847));
    outputs(4226) <= layer0_outputs(10153);
    outputs(4227) <= not(layer0_outputs(7801));
    outputs(4228) <= not(layer0_outputs(9685));
    outputs(4229) <= (layer0_outputs(4126)) and not (layer0_outputs(9524));
    outputs(4230) <= layer0_outputs(1516);
    outputs(4231) <= not(layer0_outputs(8498));
    outputs(4232) <= not(layer0_outputs(8936));
    outputs(4233) <= (layer0_outputs(1475)) or (layer0_outputs(1105));
    outputs(4234) <= layer0_outputs(2982);
    outputs(4235) <= not(layer0_outputs(1955)) or (layer0_outputs(6946));
    outputs(4236) <= (layer0_outputs(1681)) and (layer0_outputs(7750));
    outputs(4237) <= layer0_outputs(3748);
    outputs(4238) <= not(layer0_outputs(7642));
    outputs(4239) <= (layer0_outputs(7388)) xor (layer0_outputs(7071));
    outputs(4240) <= (layer0_outputs(5178)) xor (layer0_outputs(4224));
    outputs(4241) <= not(layer0_outputs(1619));
    outputs(4242) <= not((layer0_outputs(5200)) xor (layer0_outputs(999)));
    outputs(4243) <= not((layer0_outputs(4107)) xor (layer0_outputs(9234)));
    outputs(4244) <= (layer0_outputs(5491)) and not (layer0_outputs(9612));
    outputs(4245) <= (layer0_outputs(2790)) and not (layer0_outputs(4032));
    outputs(4246) <= not((layer0_outputs(36)) xor (layer0_outputs(3005)));
    outputs(4247) <= layer0_outputs(7533);
    outputs(4248) <= layer0_outputs(861);
    outputs(4249) <= not((layer0_outputs(3280)) xor (layer0_outputs(1972)));
    outputs(4250) <= layer0_outputs(4706);
    outputs(4251) <= (layer0_outputs(6352)) and not (layer0_outputs(7766));
    outputs(4252) <= not(layer0_outputs(3935));
    outputs(4253) <= '0';
    outputs(4254) <= layer0_outputs(4573);
    outputs(4255) <= layer0_outputs(8712);
    outputs(4256) <= (layer0_outputs(9516)) xor (layer0_outputs(4998));
    outputs(4257) <= '0';
    outputs(4258) <= (layer0_outputs(3388)) and not (layer0_outputs(3241));
    outputs(4259) <= layer0_outputs(3261);
    outputs(4260) <= layer0_outputs(8876);
    outputs(4261) <= (layer0_outputs(3072)) xor (layer0_outputs(5170));
    outputs(4262) <= not(layer0_outputs(4462)) or (layer0_outputs(2167));
    outputs(4263) <= (layer0_outputs(1100)) and not (layer0_outputs(3138));
    outputs(4264) <= not((layer0_outputs(9016)) xor (layer0_outputs(1284)));
    outputs(4265) <= not(layer0_outputs(1760));
    outputs(4266) <= not(layer0_outputs(5566));
    outputs(4267) <= (layer0_outputs(10173)) xor (layer0_outputs(8363));
    outputs(4268) <= not(layer0_outputs(2667));
    outputs(4269) <= (layer0_outputs(8327)) and not (layer0_outputs(4691));
    outputs(4270) <= not(layer0_outputs(9627));
    outputs(4271) <= layer0_outputs(4524);
    outputs(4272) <= layer0_outputs(5897);
    outputs(4273) <= layer0_outputs(3158);
    outputs(4274) <= not(layer0_outputs(9037)) or (layer0_outputs(650));
    outputs(4275) <= layer0_outputs(6545);
    outputs(4276) <= not((layer0_outputs(6006)) xor (layer0_outputs(5777)));
    outputs(4277) <= not((layer0_outputs(8502)) or (layer0_outputs(9998)));
    outputs(4278) <= (layer0_outputs(7698)) and not (layer0_outputs(8266));
    outputs(4279) <= (layer0_outputs(3558)) and not (layer0_outputs(3016));
    outputs(4280) <= layer0_outputs(1389);
    outputs(4281) <= (layer0_outputs(7167)) and not (layer0_outputs(5345));
    outputs(4282) <= '0';
    outputs(4283) <= not((layer0_outputs(9143)) xor (layer0_outputs(5150)));
    outputs(4284) <= (layer0_outputs(2871)) xor (layer0_outputs(7411));
    outputs(4285) <= (layer0_outputs(5730)) and not (layer0_outputs(7140));
    outputs(4286) <= not((layer0_outputs(2485)) or (layer0_outputs(3919)));
    outputs(4287) <= not((layer0_outputs(1189)) xor (layer0_outputs(9937)));
    outputs(4288) <= not((layer0_outputs(5166)) xor (layer0_outputs(3046)));
    outputs(4289) <= not(layer0_outputs(5620));
    outputs(4290) <= layer0_outputs(8858);
    outputs(4291) <= (layer0_outputs(162)) and not (layer0_outputs(3184));
    outputs(4292) <= (layer0_outputs(6967)) xor (layer0_outputs(2182));
    outputs(4293) <= (layer0_outputs(3839)) xor (layer0_outputs(1960));
    outputs(4294) <= not((layer0_outputs(2235)) xor (layer0_outputs(2826)));
    outputs(4295) <= layer0_outputs(7577);
    outputs(4296) <= not((layer0_outputs(5188)) and (layer0_outputs(5877)));
    outputs(4297) <= not(layer0_outputs(6683)) or (layer0_outputs(1396));
    outputs(4298) <= (layer0_outputs(632)) and not (layer0_outputs(482));
    outputs(4299) <= layer0_outputs(2487);
    outputs(4300) <= layer0_outputs(857);
    outputs(4301) <= not((layer0_outputs(7805)) xor (layer0_outputs(7314)));
    outputs(4302) <= not(layer0_outputs(3556));
    outputs(4303) <= layer0_outputs(4934);
    outputs(4304) <= '1';
    outputs(4305) <= not(layer0_outputs(6662));
    outputs(4306) <= not((layer0_outputs(1043)) xor (layer0_outputs(7102)));
    outputs(4307) <= (layer0_outputs(9744)) and not (layer0_outputs(332));
    outputs(4308) <= (layer0_outputs(5160)) and (layer0_outputs(6717));
    outputs(4309) <= (layer0_outputs(5819)) xor (layer0_outputs(5411));
    outputs(4310) <= not((layer0_outputs(10085)) or (layer0_outputs(8619)));
    outputs(4311) <= not((layer0_outputs(5615)) xor (layer0_outputs(7857)));
    outputs(4312) <= (layer0_outputs(7121)) xor (layer0_outputs(4839));
    outputs(4313) <= layer0_outputs(1985);
    outputs(4314) <= not((layer0_outputs(8839)) or (layer0_outputs(4582)));
    outputs(4315) <= (layer0_outputs(7095)) xor (layer0_outputs(982));
    outputs(4316) <= (layer0_outputs(3621)) xor (layer0_outputs(1423));
    outputs(4317) <= not(layer0_outputs(4848));
    outputs(4318) <= (layer0_outputs(5666)) and not (layer0_outputs(2832));
    outputs(4319) <= (layer0_outputs(2243)) xor (layer0_outputs(8294));
    outputs(4320) <= (layer0_outputs(5626)) and (layer0_outputs(675));
    outputs(4321) <= layer0_outputs(8000);
    outputs(4322) <= not(layer0_outputs(3110)) or (layer0_outputs(5585));
    outputs(4323) <= not((layer0_outputs(1243)) or (layer0_outputs(6691)));
    outputs(4324) <= (layer0_outputs(1027)) and not (layer0_outputs(9259));
    outputs(4325) <= (layer0_outputs(18)) and not (layer0_outputs(8991));
    outputs(4326) <= layer0_outputs(5857);
    outputs(4327) <= not(layer0_outputs(9619));
    outputs(4328) <= (layer0_outputs(7727)) xor (layer0_outputs(308));
    outputs(4329) <= (layer0_outputs(2591)) xor (layer0_outputs(4494));
    outputs(4330) <= not((layer0_outputs(833)) xor (layer0_outputs(7413)));
    outputs(4331) <= layer0_outputs(10015);
    outputs(4332) <= (layer0_outputs(3486)) and not (layer0_outputs(5937));
    outputs(4333) <= (layer0_outputs(9577)) xor (layer0_outputs(1614));
    outputs(4334) <= layer0_outputs(4560);
    outputs(4335) <= layer0_outputs(9932);
    outputs(4336) <= not(layer0_outputs(8342));
    outputs(4337) <= layer0_outputs(7228);
    outputs(4338) <= (layer0_outputs(10114)) and not (layer0_outputs(874));
    outputs(4339) <= not(layer0_outputs(7656)) or (layer0_outputs(4313));
    outputs(4340) <= (layer0_outputs(1632)) and (layer0_outputs(9982));
    outputs(4341) <= (layer0_outputs(5829)) and not (layer0_outputs(8269));
    outputs(4342) <= not(layer0_outputs(325));
    outputs(4343) <= not((layer0_outputs(5900)) xor (layer0_outputs(5863)));
    outputs(4344) <= (layer0_outputs(8810)) and not (layer0_outputs(2207));
    outputs(4345) <= not((layer0_outputs(4261)) xor (layer0_outputs(5482)));
    outputs(4346) <= not(layer0_outputs(2108)) or (layer0_outputs(5586));
    outputs(4347) <= not((layer0_outputs(9908)) xor (layer0_outputs(1518)));
    outputs(4348) <= layer0_outputs(5803);
    outputs(4349) <= not(layer0_outputs(5613)) or (layer0_outputs(9501));
    outputs(4350) <= not(layer0_outputs(4104));
    outputs(4351) <= not(layer0_outputs(7538));
    outputs(4352) <= layer0_outputs(1641);
    outputs(4353) <= not(layer0_outputs(3851));
    outputs(4354) <= (layer0_outputs(5244)) xor (layer0_outputs(7094));
    outputs(4355) <= (layer0_outputs(7472)) and not (layer0_outputs(5826));
    outputs(4356) <= (layer0_outputs(4907)) and not (layer0_outputs(4934));
    outputs(4357) <= not(layer0_outputs(4260));
    outputs(4358) <= not(layer0_outputs(2419));
    outputs(4359) <= not((layer0_outputs(4930)) xor (layer0_outputs(1668)));
    outputs(4360) <= (layer0_outputs(6644)) xor (layer0_outputs(9233));
    outputs(4361) <= (layer0_outputs(7501)) xor (layer0_outputs(4260));
    outputs(4362) <= (layer0_outputs(9726)) and not (layer0_outputs(778));
    outputs(4363) <= (layer0_outputs(3232)) and not (layer0_outputs(1348));
    outputs(4364) <= (layer0_outputs(4229)) xor (layer0_outputs(1085));
    outputs(4365) <= (layer0_outputs(4949)) and not (layer0_outputs(2401));
    outputs(4366) <= layer0_outputs(6711);
    outputs(4367) <= not(layer0_outputs(8989));
    outputs(4368) <= (layer0_outputs(10096)) and (layer0_outputs(3798));
    outputs(4369) <= layer0_outputs(6864);
    outputs(4370) <= (layer0_outputs(1312)) xor (layer0_outputs(6040));
    outputs(4371) <= not(layer0_outputs(7293));
    outputs(4372) <= not((layer0_outputs(5197)) or (layer0_outputs(6230)));
    outputs(4373) <= (layer0_outputs(6359)) and (layer0_outputs(8411));
    outputs(4374) <= not((layer0_outputs(913)) or (layer0_outputs(8577)));
    outputs(4375) <= not(layer0_outputs(6622));
    outputs(4376) <= layer0_outputs(1468);
    outputs(4377) <= layer0_outputs(4265);
    outputs(4378) <= not((layer0_outputs(8148)) or (layer0_outputs(5727)));
    outputs(4379) <= not((layer0_outputs(3119)) or (layer0_outputs(7738)));
    outputs(4380) <= (layer0_outputs(1096)) and (layer0_outputs(6079));
    outputs(4381) <= not((layer0_outputs(4303)) and (layer0_outputs(6728)));
    outputs(4382) <= not(layer0_outputs(7887));
    outputs(4383) <= layer0_outputs(6047);
    outputs(4384) <= (layer0_outputs(8328)) and (layer0_outputs(803));
    outputs(4385) <= layer0_outputs(1380);
    outputs(4386) <= (layer0_outputs(5939)) xor (layer0_outputs(8120));
    outputs(4387) <= (layer0_outputs(4480)) xor (layer0_outputs(6396));
    outputs(4388) <= layer0_outputs(2836);
    outputs(4389) <= (layer0_outputs(544)) and not (layer0_outputs(6599));
    outputs(4390) <= layer0_outputs(9952);
    outputs(4391) <= (layer0_outputs(2894)) and (layer0_outputs(4792));
    outputs(4392) <= not(layer0_outputs(2747));
    outputs(4393) <= not((layer0_outputs(7137)) and (layer0_outputs(4954)));
    outputs(4394) <= not(layer0_outputs(8142));
    outputs(4395) <= layer0_outputs(5634);
    outputs(4396) <= (layer0_outputs(10078)) and (layer0_outputs(5548));
    outputs(4397) <= not((layer0_outputs(6811)) or (layer0_outputs(9587)));
    outputs(4398) <= not((layer0_outputs(1281)) or (layer0_outputs(5980)));
    outputs(4399) <= (layer0_outputs(6981)) and not (layer0_outputs(5292));
    outputs(4400) <= layer0_outputs(8372);
    outputs(4401) <= not(layer0_outputs(8093)) or (layer0_outputs(3548));
    outputs(4402) <= '0';
    outputs(4403) <= not((layer0_outputs(6303)) or (layer0_outputs(4143)));
    outputs(4404) <= not(layer0_outputs(10037));
    outputs(4405) <= (layer0_outputs(6165)) and not (layer0_outputs(1872));
    outputs(4406) <= (layer0_outputs(8873)) and (layer0_outputs(8934));
    outputs(4407) <= (layer0_outputs(3947)) and (layer0_outputs(122));
    outputs(4408) <= (layer0_outputs(6440)) xor (layer0_outputs(4472));
    outputs(4409) <= not(layer0_outputs(301));
    outputs(4410) <= not(layer0_outputs(8480));
    outputs(4411) <= not((layer0_outputs(8834)) xor (layer0_outputs(5513)));
    outputs(4412) <= (layer0_outputs(3270)) and not (layer0_outputs(2162));
    outputs(4413) <= (layer0_outputs(702)) and not (layer0_outputs(5591));
    outputs(4414) <= (layer0_outputs(8264)) xor (layer0_outputs(7572));
    outputs(4415) <= not((layer0_outputs(7676)) or (layer0_outputs(5196)));
    outputs(4416) <= '0';
    outputs(4417) <= layer0_outputs(9278);
    outputs(4418) <= not(layer0_outputs(1003)) or (layer0_outputs(1459));
    outputs(4419) <= layer0_outputs(6272);
    outputs(4420) <= not(layer0_outputs(9051)) or (layer0_outputs(5976));
    outputs(4421) <= (layer0_outputs(6303)) xor (layer0_outputs(619));
    outputs(4422) <= not(layer0_outputs(1733)) or (layer0_outputs(8447));
    outputs(4423) <= not(layer0_outputs(4252));
    outputs(4424) <= layer0_outputs(8957);
    outputs(4425) <= not((layer0_outputs(3522)) xor (layer0_outputs(2173)));
    outputs(4426) <= not((layer0_outputs(5485)) xor (layer0_outputs(5523)));
    outputs(4427) <= (layer0_outputs(3566)) xor (layer0_outputs(7096));
    outputs(4428) <= layer0_outputs(7169);
    outputs(4429) <= layer0_outputs(1364);
    outputs(4430) <= (layer0_outputs(4328)) and not (layer0_outputs(1144));
    outputs(4431) <= (layer0_outputs(6132)) and (layer0_outputs(3056));
    outputs(4432) <= not((layer0_outputs(5149)) or (layer0_outputs(7202)));
    outputs(4433) <= not(layer0_outputs(3201));
    outputs(4434) <= layer0_outputs(4199);
    outputs(4435) <= (layer0_outputs(2283)) and (layer0_outputs(2014));
    outputs(4436) <= not(layer0_outputs(2707));
    outputs(4437) <= layer0_outputs(3523);
    outputs(4438) <= not((layer0_outputs(6028)) xor (layer0_outputs(3310)));
    outputs(4439) <= not((layer0_outputs(1331)) or (layer0_outputs(5689)));
    outputs(4440) <= layer0_outputs(3720);
    outputs(4441) <= not(layer0_outputs(7359));
    outputs(4442) <= not(layer0_outputs(8859));
    outputs(4443) <= not((layer0_outputs(9537)) xor (layer0_outputs(8744)));
    outputs(4444) <= layer0_outputs(3102);
    outputs(4445) <= layer0_outputs(5923);
    outputs(4446) <= (layer0_outputs(5131)) and not (layer0_outputs(3015));
    outputs(4447) <= not(layer0_outputs(5734));
    outputs(4448) <= not(layer0_outputs(1136));
    outputs(4449) <= not(layer0_outputs(8523));
    outputs(4450) <= (layer0_outputs(5372)) and not (layer0_outputs(9172));
    outputs(4451) <= (layer0_outputs(8470)) or (layer0_outputs(3434));
    outputs(4452) <= (layer0_outputs(7389)) xor (layer0_outputs(2911));
    outputs(4453) <= (layer0_outputs(9210)) xor (layer0_outputs(8546));
    outputs(4454) <= not((layer0_outputs(1700)) xor (layer0_outputs(3652)));
    outputs(4455) <= not(layer0_outputs(8764));
    outputs(4456) <= not(layer0_outputs(6616)) or (layer0_outputs(7397));
    outputs(4457) <= not((layer0_outputs(9008)) or (layer0_outputs(6495)));
    outputs(4458) <= (layer0_outputs(7688)) and (layer0_outputs(3900));
    outputs(4459) <= not(layer0_outputs(6101));
    outputs(4460) <= layer0_outputs(8134);
    outputs(4461) <= not(layer0_outputs(1971));
    outputs(4462) <= not((layer0_outputs(7979)) or (layer0_outputs(9389)));
    outputs(4463) <= (layer0_outputs(7961)) and not (layer0_outputs(6046));
    outputs(4464) <= not((layer0_outputs(4277)) xor (layer0_outputs(9914)));
    outputs(4465) <= layer0_outputs(10073);
    outputs(4466) <= layer0_outputs(5926);
    outputs(4467) <= not(layer0_outputs(9565));
    outputs(4468) <= not(layer0_outputs(8775));
    outputs(4469) <= not(layer0_outputs(9955)) or (layer0_outputs(1134));
    outputs(4470) <= not(layer0_outputs(4505));
    outputs(4471) <= not(layer0_outputs(49));
    outputs(4472) <= layer0_outputs(5446);
    outputs(4473) <= not((layer0_outputs(8196)) or (layer0_outputs(7067)));
    outputs(4474) <= not((layer0_outputs(2410)) xor (layer0_outputs(443)));
    outputs(4475) <= (layer0_outputs(6557)) and (layer0_outputs(3650));
    outputs(4476) <= not((layer0_outputs(6818)) xor (layer0_outputs(4763)));
    outputs(4477) <= not((layer0_outputs(5558)) xor (layer0_outputs(3461)));
    outputs(4478) <= not(layer0_outputs(3312));
    outputs(4479) <= (layer0_outputs(8263)) and not (layer0_outputs(4585));
    outputs(4480) <= not(layer0_outputs(877));
    outputs(4481) <= not(layer0_outputs(8348));
    outputs(4482) <= not((layer0_outputs(2526)) xor (layer0_outputs(8016)));
    outputs(4483) <= (layer0_outputs(9060)) xor (layer0_outputs(8703));
    outputs(4484) <= not((layer0_outputs(10149)) xor (layer0_outputs(9734)));
    outputs(4485) <= not((layer0_outputs(231)) xor (layer0_outputs(3939)));
    outputs(4486) <= (layer0_outputs(8928)) xor (layer0_outputs(2078));
    outputs(4487) <= not(layer0_outputs(3605));
    outputs(4488) <= layer0_outputs(2685);
    outputs(4489) <= not((layer0_outputs(565)) xor (layer0_outputs(6956)));
    outputs(4490) <= (layer0_outputs(2935)) xor (layer0_outputs(5970));
    outputs(4491) <= (layer0_outputs(9591)) or (layer0_outputs(10003));
    outputs(4492) <= (layer0_outputs(4791)) or (layer0_outputs(837));
    outputs(4493) <= not(layer0_outputs(5212));
    outputs(4494) <= layer0_outputs(9890);
    outputs(4495) <= layer0_outputs(1294);
    outputs(4496) <= not(layer0_outputs(4802)) or (layer0_outputs(4864));
    outputs(4497) <= (layer0_outputs(2688)) and not (layer0_outputs(2637));
    outputs(4498) <= (layer0_outputs(503)) xor (layer0_outputs(8431));
    outputs(4499) <= not(layer0_outputs(4397));
    outputs(4500) <= (layer0_outputs(5048)) and (layer0_outputs(5717));
    outputs(4501) <= not(layer0_outputs(4));
    outputs(4502) <= (layer0_outputs(2255)) xor (layer0_outputs(9376));
    outputs(4503) <= layer0_outputs(1255);
    outputs(4504) <= (layer0_outputs(8307)) xor (layer0_outputs(5971));
    outputs(4505) <= not(layer0_outputs(1477));
    outputs(4506) <= (layer0_outputs(115)) xor (layer0_outputs(1922));
    outputs(4507) <= (layer0_outputs(3030)) and not (layer0_outputs(6902));
    outputs(4508) <= layer0_outputs(1397);
    outputs(4509) <= layer0_outputs(8058);
    outputs(4510) <= not((layer0_outputs(3565)) xor (layer0_outputs(6989)));
    outputs(4511) <= not((layer0_outputs(6528)) xor (layer0_outputs(6122)));
    outputs(4512) <= not(layer0_outputs(640));
    outputs(4513) <= '0';
    outputs(4514) <= not(layer0_outputs(8776));
    outputs(4515) <= layer0_outputs(6814);
    outputs(4516) <= (layer0_outputs(6684)) xor (layer0_outputs(9164));
    outputs(4517) <= not(layer0_outputs(7672));
    outputs(4518) <= not(layer0_outputs(1544));
    outputs(4519) <= not((layer0_outputs(4125)) xor (layer0_outputs(283)));
    outputs(4520) <= not(layer0_outputs(9634));
    outputs(4521) <= not(layer0_outputs(9073));
    outputs(4522) <= layer0_outputs(4348);
    outputs(4523) <= layer0_outputs(3512);
    outputs(4524) <= (layer0_outputs(8318)) xor (layer0_outputs(5175));
    outputs(4525) <= layer0_outputs(7157);
    outputs(4526) <= layer0_outputs(3281);
    outputs(4527) <= (layer0_outputs(1110)) xor (layer0_outputs(6132));
    outputs(4528) <= (layer0_outputs(3555)) and (layer0_outputs(513));
    outputs(4529) <= layer0_outputs(3212);
    outputs(4530) <= not((layer0_outputs(3315)) and (layer0_outputs(1589)));
    outputs(4531) <= not(layer0_outputs(9715));
    outputs(4532) <= (layer0_outputs(607)) xor (layer0_outputs(1665));
    outputs(4533) <= not((layer0_outputs(1931)) xor (layer0_outputs(849)));
    outputs(4534) <= layer0_outputs(3320);
    outputs(4535) <= (layer0_outputs(3878)) and not (layer0_outputs(7623));
    outputs(4536) <= not(layer0_outputs(7438));
    outputs(4537) <= (layer0_outputs(4827)) and (layer0_outputs(6318));
    outputs(4538) <= (layer0_outputs(7768)) or (layer0_outputs(7925));
    outputs(4539) <= not(layer0_outputs(3903));
    outputs(4540) <= not((layer0_outputs(4939)) xor (layer0_outputs(8304)));
    outputs(4541) <= not(layer0_outputs(3175));
    outputs(4542) <= layer0_outputs(7911);
    outputs(4543) <= not(layer0_outputs(4581));
    outputs(4544) <= layer0_outputs(7627);
    outputs(4545) <= (layer0_outputs(250)) and (layer0_outputs(367));
    outputs(4546) <= not(layer0_outputs(9716));
    outputs(4547) <= (layer0_outputs(2404)) and not (layer0_outputs(2366));
    outputs(4548) <= not(layer0_outputs(1247)) or (layer0_outputs(5339));
    outputs(4549) <= (layer0_outputs(2759)) and (layer0_outputs(3237));
    outputs(4550) <= not((layer0_outputs(6290)) or (layer0_outputs(1944)));
    outputs(4551) <= (layer0_outputs(1831)) and not (layer0_outputs(3565));
    outputs(4552) <= layer0_outputs(4400);
    outputs(4553) <= not(layer0_outputs(1301));
    outputs(4554) <= not(layer0_outputs(5893));
    outputs(4555) <= (layer0_outputs(3716)) and (layer0_outputs(6466));
    outputs(4556) <= layer0_outputs(9048);
    outputs(4557) <= not(layer0_outputs(9423));
    outputs(4558) <= (layer0_outputs(2686)) xor (layer0_outputs(9632));
    outputs(4559) <= (layer0_outputs(1082)) and not (layer0_outputs(4032));
    outputs(4560) <= (layer0_outputs(8069)) xor (layer0_outputs(8320));
    outputs(4561) <= (layer0_outputs(7639)) and (layer0_outputs(6890));
    outputs(4562) <= not(layer0_outputs(3026));
    outputs(4563) <= not((layer0_outputs(4294)) or (layer0_outputs(3528)));
    outputs(4564) <= (layer0_outputs(7609)) and not (layer0_outputs(8833));
    outputs(4565) <= not((layer0_outputs(4998)) or (layer0_outputs(4197)));
    outputs(4566) <= not(layer0_outputs(3991));
    outputs(4567) <= (layer0_outputs(6019)) and (layer0_outputs(7907));
    outputs(4568) <= not((layer0_outputs(8241)) and (layer0_outputs(5371)));
    outputs(4569) <= (layer0_outputs(218)) and not (layer0_outputs(5851));
    outputs(4570) <= not(layer0_outputs(2038));
    outputs(4571) <= layer0_outputs(7956);
    outputs(4572) <= layer0_outputs(9533);
    outputs(4573) <= not(layer0_outputs(3094));
    outputs(4574) <= not(layer0_outputs(3938)) or (layer0_outputs(3544));
    outputs(4575) <= not((layer0_outputs(412)) or (layer0_outputs(2028)));
    outputs(4576) <= layer0_outputs(4736);
    outputs(4577) <= layer0_outputs(8236);
    outputs(4578) <= layer0_outputs(7003);
    outputs(4579) <= layer0_outputs(3682);
    outputs(4580) <= not(layer0_outputs(3990)) or (layer0_outputs(8563));
    outputs(4581) <= layer0_outputs(1543);
    outputs(4582) <= layer0_outputs(7884);
    outputs(4583) <= layer0_outputs(4325);
    outputs(4584) <= not(layer0_outputs(2738));
    outputs(4585) <= not((layer0_outputs(9749)) or (layer0_outputs(29)));
    outputs(4586) <= layer0_outputs(3114);
    outputs(4587) <= not((layer0_outputs(8666)) xor (layer0_outputs(9329)));
    outputs(4588) <= not(layer0_outputs(2571));
    outputs(4589) <= layer0_outputs(651);
    outputs(4590) <= not((layer0_outputs(713)) xor (layer0_outputs(9531)));
    outputs(4591) <= layer0_outputs(9170);
    outputs(4592) <= (layer0_outputs(7441)) or (layer0_outputs(6048));
    outputs(4593) <= layer0_outputs(8799);
    outputs(4594) <= (layer0_outputs(3621)) xor (layer0_outputs(9796));
    outputs(4595) <= (layer0_outputs(4228)) and not (layer0_outputs(3328));
    outputs(4596) <= not((layer0_outputs(4182)) or (layer0_outputs(8255)));
    outputs(4597) <= '0';
    outputs(4598) <= (layer0_outputs(1888)) and (layer0_outputs(9157));
    outputs(4599) <= not(layer0_outputs(7160));
    outputs(4600) <= (layer0_outputs(4180)) xor (layer0_outputs(4880));
    outputs(4601) <= layer0_outputs(1460);
    outputs(4602) <= not(layer0_outputs(841));
    outputs(4603) <= not((layer0_outputs(2712)) xor (layer0_outputs(7136)));
    outputs(4604) <= '0';
    outputs(4605) <= layer0_outputs(2027);
    outputs(4606) <= not(layer0_outputs(9576)) or (layer0_outputs(5875));
    outputs(4607) <= not(layer0_outputs(7809));
    outputs(4608) <= (layer0_outputs(9708)) and not (layer0_outputs(3617));
    outputs(4609) <= (layer0_outputs(2712)) xor (layer0_outputs(9984));
    outputs(4610) <= not(layer0_outputs(605));
    outputs(4611) <= not((layer0_outputs(7697)) xor (layer0_outputs(5426)));
    outputs(4612) <= layer0_outputs(4385);
    outputs(4613) <= layer0_outputs(4202);
    outputs(4614) <= not((layer0_outputs(5452)) xor (layer0_outputs(6346)));
    outputs(4615) <= (layer0_outputs(4363)) or (layer0_outputs(6556));
    outputs(4616) <= (layer0_outputs(2291)) xor (layer0_outputs(5203));
    outputs(4617) <= (layer0_outputs(7511)) and not (layer0_outputs(6109));
    outputs(4618) <= (layer0_outputs(3448)) xor (layer0_outputs(8032));
    outputs(4619) <= layer0_outputs(10052);
    outputs(4620) <= (layer0_outputs(7014)) xor (layer0_outputs(1926));
    outputs(4621) <= (layer0_outputs(4155)) and not (layer0_outputs(2718));
    outputs(4622) <= not(layer0_outputs(3919)) or (layer0_outputs(6229));
    outputs(4623) <= not(layer0_outputs(48));
    outputs(4624) <= not((layer0_outputs(9131)) or (layer0_outputs(3663)));
    outputs(4625) <= (layer0_outputs(8641)) and not (layer0_outputs(8334));
    outputs(4626) <= (layer0_outputs(4206)) and not (layer0_outputs(2064));
    outputs(4627) <= layer0_outputs(4272);
    outputs(4628) <= not(layer0_outputs(10010)) or (layer0_outputs(9689));
    outputs(4629) <= layer0_outputs(7452);
    outputs(4630) <= (layer0_outputs(5314)) xor (layer0_outputs(612));
    outputs(4631) <= not(layer0_outputs(9354));
    outputs(4632) <= (layer0_outputs(7801)) xor (layer0_outputs(3847));
    outputs(4633) <= layer0_outputs(8847);
    outputs(4634) <= not(layer0_outputs(1063));
    outputs(4635) <= not((layer0_outputs(4683)) or (layer0_outputs(41)));
    outputs(4636) <= not((layer0_outputs(7131)) or (layer0_outputs(7162)));
    outputs(4637) <= not(layer0_outputs(2206));
    outputs(4638) <= (layer0_outputs(9362)) and not (layer0_outputs(5592));
    outputs(4639) <= layer0_outputs(2539);
    outputs(4640) <= layer0_outputs(65);
    outputs(4641) <= not((layer0_outputs(9921)) xor (layer0_outputs(4701)));
    outputs(4642) <= not(layer0_outputs(6600));
    outputs(4643) <= not(layer0_outputs(7655));
    outputs(4644) <= layer0_outputs(4235);
    outputs(4645) <= not(layer0_outputs(4085));
    outputs(4646) <= not((layer0_outputs(2697)) or (layer0_outputs(8849)));
    outputs(4647) <= not((layer0_outputs(6931)) xor (layer0_outputs(5828)));
    outputs(4648) <= layer0_outputs(10099);
    outputs(4649) <= (layer0_outputs(1208)) and not (layer0_outputs(3757));
    outputs(4650) <= (layer0_outputs(4318)) xor (layer0_outputs(6546));
    outputs(4651) <= not(layer0_outputs(6124)) or (layer0_outputs(7690));
    outputs(4652) <= not(layer0_outputs(6063));
    outputs(4653) <= (layer0_outputs(2785)) and not (layer0_outputs(6138));
    outputs(4654) <= (layer0_outputs(245)) and not (layer0_outputs(1617));
    outputs(4655) <= (layer0_outputs(3463)) and (layer0_outputs(9944));
    outputs(4656) <= layer0_outputs(2123);
    outputs(4657) <= (layer0_outputs(10039)) and (layer0_outputs(7627));
    outputs(4658) <= not((layer0_outputs(2154)) xor (layer0_outputs(8407)));
    outputs(4659) <= (layer0_outputs(6675)) and not (layer0_outputs(3829));
    outputs(4660) <= not((layer0_outputs(2076)) or (layer0_outputs(456)));
    outputs(4661) <= (layer0_outputs(5098)) and not (layer0_outputs(5886));
    outputs(4662) <= not((layer0_outputs(389)) or (layer0_outputs(7358)));
    outputs(4663) <= not(layer0_outputs(5011)) or (layer0_outputs(888));
    outputs(4664) <= (layer0_outputs(2340)) and not (layer0_outputs(6347));
    outputs(4665) <= (layer0_outputs(3528)) xor (layer0_outputs(9275));
    outputs(4666) <= not((layer0_outputs(1830)) xor (layer0_outputs(4350)));
    outputs(4667) <= not((layer0_outputs(8936)) or (layer0_outputs(7473)));
    outputs(4668) <= layer0_outputs(1659);
    outputs(4669) <= layer0_outputs(9603);
    outputs(4670) <= not(layer0_outputs(7805));
    outputs(4671) <= (layer0_outputs(1306)) xor (layer0_outputs(9076));
    outputs(4672) <= not(layer0_outputs(9201));
    outputs(4673) <= not((layer0_outputs(5721)) xor (layer0_outputs(3348)));
    outputs(4674) <= (layer0_outputs(174)) and (layer0_outputs(5473));
    outputs(4675) <= layer0_outputs(4193);
    outputs(4676) <= layer0_outputs(4913);
    outputs(4677) <= not((layer0_outputs(2824)) or (layer0_outputs(7074)));
    outputs(4678) <= (layer0_outputs(9580)) and not (layer0_outputs(5091));
    outputs(4679) <= (layer0_outputs(830)) and not (layer0_outputs(1974));
    outputs(4680) <= (layer0_outputs(2809)) and not (layer0_outputs(2140));
    outputs(4681) <= (layer0_outputs(630)) and (layer0_outputs(3441));
    outputs(4682) <= (layer0_outputs(8355)) and (layer0_outputs(2080));
    outputs(4683) <= not((layer0_outputs(8222)) and (layer0_outputs(8018)));
    outputs(4684) <= layer0_outputs(1593);
    outputs(4685) <= layer0_outputs(6947);
    outputs(4686) <= not(layer0_outputs(5747));
    outputs(4687) <= not((layer0_outputs(10035)) and (layer0_outputs(7817)));
    outputs(4688) <= not((layer0_outputs(1410)) or (layer0_outputs(453)));
    outputs(4689) <= not((layer0_outputs(3342)) xor (layer0_outputs(477)));
    outputs(4690) <= not((layer0_outputs(3698)) xor (layer0_outputs(1824)));
    outputs(4691) <= (layer0_outputs(1503)) and not (layer0_outputs(3763));
    outputs(4692) <= not(layer0_outputs(456));
    outputs(4693) <= layer0_outputs(349);
    outputs(4694) <= not((layer0_outputs(4344)) xor (layer0_outputs(2411)));
    outputs(4695) <= (layer0_outputs(9798)) and not (layer0_outputs(6865));
    outputs(4696) <= (layer0_outputs(9250)) xor (layer0_outputs(9085));
    outputs(4697) <= not((layer0_outputs(7241)) xor (layer0_outputs(4571)));
    outputs(4698) <= (layer0_outputs(1770)) and not (layer0_outputs(7420));
    outputs(4699) <= layer0_outputs(5429);
    outputs(4700) <= not((layer0_outputs(3800)) or (layer0_outputs(5764)));
    outputs(4701) <= (layer0_outputs(118)) xor (layer0_outputs(4458));
    outputs(4702) <= not((layer0_outputs(8125)) xor (layer0_outputs(2751)));
    outputs(4703) <= not(layer0_outputs(691));
    outputs(4704) <= layer0_outputs(3815);
    outputs(4705) <= not(layer0_outputs(8731));
    outputs(4706) <= not(layer0_outputs(1513));
    outputs(4707) <= not(layer0_outputs(7583));
    outputs(4708) <= not(layer0_outputs(10106));
    outputs(4709) <= not(layer0_outputs(2117));
    outputs(4710) <= not((layer0_outputs(9223)) or (layer0_outputs(5498)));
    outputs(4711) <= not((layer0_outputs(5768)) or (layer0_outputs(8534)));
    outputs(4712) <= layer0_outputs(3889);
    outputs(4713) <= not(layer0_outputs(3096));
    outputs(4714) <= not(layer0_outputs(2458));
    outputs(4715) <= not(layer0_outputs(6929));
    outputs(4716) <= not(layer0_outputs(3651));
    outputs(4717) <= (layer0_outputs(1878)) and not (layer0_outputs(9650));
    outputs(4718) <= (layer0_outputs(1963)) xor (layer0_outputs(583));
    outputs(4719) <= not(layer0_outputs(1752));
    outputs(4720) <= not((layer0_outputs(9950)) xor (layer0_outputs(6809)));
    outputs(4721) <= layer0_outputs(3058);
    outputs(4722) <= layer0_outputs(6240);
    outputs(4723) <= (layer0_outputs(4880)) and not (layer0_outputs(9225));
    outputs(4724) <= (layer0_outputs(7371)) and (layer0_outputs(6948));
    outputs(4725) <= (layer0_outputs(879)) and not (layer0_outputs(5982));
    outputs(4726) <= '0';
    outputs(4727) <= (layer0_outputs(8391)) and (layer0_outputs(9427));
    outputs(4728) <= not((layer0_outputs(1340)) or (layer0_outputs(1866)));
    outputs(4729) <= (layer0_outputs(3234)) and not (layer0_outputs(4035));
    outputs(4730) <= (layer0_outputs(8902)) and not (layer0_outputs(3993));
    outputs(4731) <= not(layer0_outputs(598));
    outputs(4732) <= not((layer0_outputs(1759)) xor (layer0_outputs(3155)));
    outputs(4733) <= not(layer0_outputs(2920));
    outputs(4734) <= (layer0_outputs(4191)) and (layer0_outputs(1569));
    outputs(4735) <= not((layer0_outputs(715)) xor (layer0_outputs(4990)));
    outputs(4736) <= (layer0_outputs(270)) xor (layer0_outputs(5981));
    outputs(4737) <= not((layer0_outputs(4891)) xor (layer0_outputs(5852)));
    outputs(4738) <= not((layer0_outputs(3325)) and (layer0_outputs(6971)));
    outputs(4739) <= not(layer0_outputs(4192));
    outputs(4740) <= not((layer0_outputs(7020)) xor (layer0_outputs(7210)));
    outputs(4741) <= not(layer0_outputs(288));
    outputs(4742) <= not((layer0_outputs(1383)) and (layer0_outputs(3808)));
    outputs(4743) <= layer0_outputs(3887);
    outputs(4744) <= layer0_outputs(2646);
    outputs(4745) <= (layer0_outputs(6903)) and not (layer0_outputs(4412));
    outputs(4746) <= (layer0_outputs(3547)) and not (layer0_outputs(5532));
    outputs(4747) <= layer0_outputs(5535);
    outputs(4748) <= (layer0_outputs(6931)) and not (layer0_outputs(8903));
    outputs(4749) <= layer0_outputs(516);
    outputs(4750) <= (layer0_outputs(6366)) and not (layer0_outputs(8096));
    outputs(4751) <= (layer0_outputs(1659)) xor (layer0_outputs(9193));
    outputs(4752) <= not(layer0_outputs(6405));
    outputs(4753) <= (layer0_outputs(463)) and not (layer0_outputs(9652));
    outputs(4754) <= not(layer0_outputs(7085));
    outputs(4755) <= (layer0_outputs(7001)) and not (layer0_outputs(5761));
    outputs(4756) <= not((layer0_outputs(6852)) or (layer0_outputs(9466)));
    outputs(4757) <= (layer0_outputs(1476)) and (layer0_outputs(9900));
    outputs(4758) <= not(layer0_outputs(853));
    outputs(4759) <= (layer0_outputs(1952)) and not (layer0_outputs(6593));
    outputs(4760) <= (layer0_outputs(8675)) and not (layer0_outputs(3762));
    outputs(4761) <= not(layer0_outputs(9851));
    outputs(4762) <= (layer0_outputs(3034)) and (layer0_outputs(7010));
    outputs(4763) <= (layer0_outputs(5842)) xor (layer0_outputs(3594));
    outputs(4764) <= (layer0_outputs(5995)) and not (layer0_outputs(9591));
    outputs(4765) <= not((layer0_outputs(5243)) xor (layer0_outputs(2744)));
    outputs(4766) <= not((layer0_outputs(5577)) or (layer0_outputs(9175)));
    outputs(4767) <= layer0_outputs(7845);
    outputs(4768) <= not(layer0_outputs(3859));
    outputs(4769) <= (layer0_outputs(8986)) and not (layer0_outputs(9343));
    outputs(4770) <= layer0_outputs(9245);
    outputs(4771) <= layer0_outputs(2226);
    outputs(4772) <= (layer0_outputs(4633)) or (layer0_outputs(5462));
    outputs(4773) <= not(layer0_outputs(8555));
    outputs(4774) <= not(layer0_outputs(2608));
    outputs(4775) <= (layer0_outputs(2187)) and not (layer0_outputs(2601));
    outputs(4776) <= layer0_outputs(9145);
    outputs(4777) <= not((layer0_outputs(2316)) xor (layer0_outputs(4358)));
    outputs(4778) <= (layer0_outputs(9323)) xor (layer0_outputs(67));
    outputs(4779) <= layer0_outputs(1615);
    outputs(4780) <= layer0_outputs(8536);
    outputs(4781) <= (layer0_outputs(177)) xor (layer0_outputs(4625));
    outputs(4782) <= not(layer0_outputs(4894)) or (layer0_outputs(1354));
    outputs(4783) <= (layer0_outputs(1274)) and not (layer0_outputs(788));
    outputs(4784) <= not(layer0_outputs(2269));
    outputs(4785) <= not(layer0_outputs(8380));
    outputs(4786) <= (layer0_outputs(4584)) and (layer0_outputs(8848));
    outputs(4787) <= not((layer0_outputs(5466)) or (layer0_outputs(8696)));
    outputs(4788) <= layer0_outputs(2265);
    outputs(4789) <= (layer0_outputs(7461)) and not (layer0_outputs(4247));
    outputs(4790) <= (layer0_outputs(7990)) and not (layer0_outputs(7924));
    outputs(4791) <= (layer0_outputs(9994)) xor (layer0_outputs(9593));
    outputs(4792) <= (layer0_outputs(2852)) and not (layer0_outputs(717));
    outputs(4793) <= (layer0_outputs(9892)) or (layer0_outputs(8706));
    outputs(4794) <= not(layer0_outputs(8309));
    outputs(4795) <= layer0_outputs(4861);
    outputs(4796) <= not(layer0_outputs(5748));
    outputs(4797) <= not((layer0_outputs(2427)) xor (layer0_outputs(2393)));
    outputs(4798) <= not(layer0_outputs(7846));
    outputs(4799) <= (layer0_outputs(2368)) or (layer0_outputs(3440));
    outputs(4800) <= (layer0_outputs(7472)) and not (layer0_outputs(10226));
    outputs(4801) <= layer0_outputs(3645);
    outputs(4802) <= (layer0_outputs(6904)) and not (layer0_outputs(3166));
    outputs(4803) <= (layer0_outputs(9216)) xor (layer0_outputs(8164));
    outputs(4804) <= not((layer0_outputs(9518)) xor (layer0_outputs(6584)));
    outputs(4805) <= layer0_outputs(3518);
    outputs(4806) <= layer0_outputs(4114);
    outputs(4807) <= not((layer0_outputs(3246)) xor (layer0_outputs(8298)));
    outputs(4808) <= not(layer0_outputs(5602));
    outputs(4809) <= not(layer0_outputs(3966));
    outputs(4810) <= (layer0_outputs(8047)) and (layer0_outputs(2173));
    outputs(4811) <= (layer0_outputs(8779)) and (layer0_outputs(1497));
    outputs(4812) <= layer0_outputs(2478);
    outputs(4813) <= (layer0_outputs(2234)) and (layer0_outputs(3294));
    outputs(4814) <= (layer0_outputs(393)) and not (layer0_outputs(4565));
    outputs(4815) <= not(layer0_outputs(4113));
    outputs(4816) <= (layer0_outputs(2733)) xor (layer0_outputs(6646));
    outputs(4817) <= not((layer0_outputs(3176)) and (layer0_outputs(7204)));
    outputs(4818) <= '0';
    outputs(4819) <= not(layer0_outputs(6077));
    outputs(4820) <= layer0_outputs(3500);
    outputs(4821) <= layer0_outputs(3352);
    outputs(4822) <= not(layer0_outputs(9324)) or (layer0_outputs(6159));
    outputs(4823) <= (layer0_outputs(4174)) and (layer0_outputs(752));
    outputs(4824) <= not((layer0_outputs(418)) xor (layer0_outputs(6750)));
    outputs(4825) <= (layer0_outputs(3853)) xor (layer0_outputs(4955));
    outputs(4826) <= layer0_outputs(3639);
    outputs(4827) <= not(layer0_outputs(4527));
    outputs(4828) <= layer0_outputs(6998);
    outputs(4829) <= layer0_outputs(10085);
    outputs(4830) <= not((layer0_outputs(7036)) and (layer0_outputs(5719)));
    outputs(4831) <= not(layer0_outputs(3676));
    outputs(4832) <= not((layer0_outputs(3372)) xor (layer0_outputs(875)));
    outputs(4833) <= (layer0_outputs(3037)) and not (layer0_outputs(5715));
    outputs(4834) <= not((layer0_outputs(6781)) xor (layer0_outputs(6554)));
    outputs(4835) <= not((layer0_outputs(7273)) xor (layer0_outputs(8532)));
    outputs(4836) <= not((layer0_outputs(947)) or (layer0_outputs(7144)));
    outputs(4837) <= (layer0_outputs(1153)) xor (layer0_outputs(1070));
    outputs(4838) <= (layer0_outputs(4019)) and not (layer0_outputs(8387));
    outputs(4839) <= not((layer0_outputs(496)) xor (layer0_outputs(5070)));
    outputs(4840) <= (layer0_outputs(7005)) and (layer0_outputs(6965));
    outputs(4841) <= not(layer0_outputs(8015));
    outputs(4842) <= (layer0_outputs(26)) xor (layer0_outputs(3728));
    outputs(4843) <= layer0_outputs(3243);
    outputs(4844) <= (layer0_outputs(9001)) xor (layer0_outputs(8387));
    outputs(4845) <= (layer0_outputs(7190)) and not (layer0_outputs(6109));
    outputs(4846) <= (layer0_outputs(9969)) and not (layer0_outputs(4708));
    outputs(4847) <= not(layer0_outputs(968));
    outputs(4848) <= (layer0_outputs(9554)) and (layer0_outputs(2203));
    outputs(4849) <= layer0_outputs(4873);
    outputs(4850) <= not((layer0_outputs(10032)) xor (layer0_outputs(8709)));
    outputs(4851) <= not(layer0_outputs(4330));
    outputs(4852) <= not((layer0_outputs(1925)) xor (layer0_outputs(5576)));
    outputs(4853) <= not((layer0_outputs(8576)) or (layer0_outputs(7619)));
    outputs(4854) <= not(layer0_outputs(3864));
    outputs(4855) <= layer0_outputs(4795);
    outputs(4856) <= not(layer0_outputs(7971)) or (layer0_outputs(6786));
    outputs(4857) <= not(layer0_outputs(8090));
    outputs(4858) <= (layer0_outputs(6510)) and not (layer0_outputs(9204));
    outputs(4859) <= layer0_outputs(3363);
    outputs(4860) <= not((layer0_outputs(6126)) or (layer0_outputs(8208)));
    outputs(4861) <= not((layer0_outputs(6234)) or (layer0_outputs(80)));
    outputs(4862) <= (layer0_outputs(2901)) and not (layer0_outputs(425));
    outputs(4863) <= not(layer0_outputs(6704));
    outputs(4864) <= layer0_outputs(8273);
    outputs(4865) <= not(layer0_outputs(2740));
    outputs(4866) <= (layer0_outputs(161)) and not (layer0_outputs(1224));
    outputs(4867) <= layer0_outputs(9722);
    outputs(4868) <= not(layer0_outputs(9298)) or (layer0_outputs(3924));
    outputs(4869) <= (layer0_outputs(844)) and not (layer0_outputs(8396));
    outputs(4870) <= layer0_outputs(705);
    outputs(4871) <= (layer0_outputs(3756)) and (layer0_outputs(8263));
    outputs(4872) <= layer0_outputs(349);
    outputs(4873) <= (layer0_outputs(8771)) and not (layer0_outputs(5255));
    outputs(4874) <= (layer0_outputs(6511)) and not (layer0_outputs(3846));
    outputs(4875) <= layer0_outputs(435);
    outputs(4876) <= not(layer0_outputs(4967));
    outputs(4877) <= (layer0_outputs(7087)) and (layer0_outputs(4728));
    outputs(4878) <= not(layer0_outputs(5433));
    outputs(4879) <= (layer0_outputs(4658)) and not (layer0_outputs(6593));
    outputs(4880) <= (layer0_outputs(6645)) xor (layer0_outputs(6071));
    outputs(4881) <= (layer0_outputs(2422)) xor (layer0_outputs(5852));
    outputs(4882) <= (layer0_outputs(1802)) xor (layer0_outputs(9712));
    outputs(4883) <= not((layer0_outputs(8843)) xor (layer0_outputs(8194)));
    outputs(4884) <= layer0_outputs(9493);
    outputs(4885) <= (layer0_outputs(8039)) and (layer0_outputs(8287));
    outputs(4886) <= (layer0_outputs(7272)) and not (layer0_outputs(5985));
    outputs(4887) <= (layer0_outputs(4153)) xor (layer0_outputs(9976));
    outputs(4888) <= (layer0_outputs(3244)) and (layer0_outputs(6388));
    outputs(4889) <= (layer0_outputs(1770)) xor (layer0_outputs(2946));
    outputs(4890) <= (layer0_outputs(5594)) and not (layer0_outputs(6963));
    outputs(4891) <= not(layer0_outputs(2502)) or (layer0_outputs(8186));
    outputs(4892) <= (layer0_outputs(3818)) and (layer0_outputs(759));
    outputs(4893) <= not((layer0_outputs(7297)) and (layer0_outputs(7861)));
    outputs(4894) <= not((layer0_outputs(538)) or (layer0_outputs(7588)));
    outputs(4895) <= layer0_outputs(1683);
    outputs(4896) <= not(layer0_outputs(5424));
    outputs(4897) <= (layer0_outputs(2135)) and not (layer0_outputs(7333));
    outputs(4898) <= (layer0_outputs(9832)) and (layer0_outputs(5716));
    outputs(4899) <= (layer0_outputs(7642)) xor (layer0_outputs(8525));
    outputs(4900) <= not((layer0_outputs(8657)) xor (layer0_outputs(2464)));
    outputs(4901) <= (layer0_outputs(2556)) xor (layer0_outputs(4087));
    outputs(4902) <= (layer0_outputs(10042)) xor (layer0_outputs(2530));
    outputs(4903) <= not(layer0_outputs(2134));
    outputs(4904) <= not(layer0_outputs(9462)) or (layer0_outputs(3391));
    outputs(4905) <= not(layer0_outputs(9876));
    outputs(4906) <= not((layer0_outputs(1152)) xor (layer0_outputs(1246)));
    outputs(4907) <= layer0_outputs(6814);
    outputs(4908) <= (layer0_outputs(6320)) and not (layer0_outputs(6651));
    outputs(4909) <= (layer0_outputs(1918)) and not (layer0_outputs(8884));
    outputs(4910) <= (layer0_outputs(4555)) and not (layer0_outputs(2476));
    outputs(4911) <= (layer0_outputs(10030)) xor (layer0_outputs(2542));
    outputs(4912) <= (layer0_outputs(4886)) xor (layer0_outputs(3799));
    outputs(4913) <= not((layer0_outputs(7223)) xor (layer0_outputs(1299)));
    outputs(4914) <= (layer0_outputs(9349)) xor (layer0_outputs(292));
    outputs(4915) <= layer0_outputs(5356);
    outputs(4916) <= not((layer0_outputs(7248)) or (layer0_outputs(9536)));
    outputs(4917) <= layer0_outputs(604);
    outputs(4918) <= layer0_outputs(5089);
    outputs(4919) <= not(layer0_outputs(7279));
    outputs(4920) <= not(layer0_outputs(5487));
    outputs(4921) <= (layer0_outputs(7456)) and not (layer0_outputs(9206));
    outputs(4922) <= not(layer0_outputs(80));
    outputs(4923) <= (layer0_outputs(2335)) and (layer0_outputs(8483));
    outputs(4924) <= not((layer0_outputs(8732)) or (layer0_outputs(6380)));
    outputs(4925) <= not((layer0_outputs(306)) or (layer0_outputs(1289)));
    outputs(4926) <= not(layer0_outputs(1792));
    outputs(4927) <= not(layer0_outputs(3754));
    outputs(4928) <= (layer0_outputs(4205)) and not (layer0_outputs(9471));
    outputs(4929) <= layer0_outputs(3376);
    outputs(4930) <= (layer0_outputs(2958)) and (layer0_outputs(5335));
    outputs(4931) <= not(layer0_outputs(848)) or (layer0_outputs(4843));
    outputs(4932) <= not((layer0_outputs(7143)) xor (layer0_outputs(4554)));
    outputs(4933) <= (layer0_outputs(8484)) and not (layer0_outputs(8854));
    outputs(4934) <= layer0_outputs(2065);
    outputs(4935) <= (layer0_outputs(6966)) and not (layer0_outputs(5104));
    outputs(4936) <= (layer0_outputs(3659)) or (layer0_outputs(5340));
    outputs(4937) <= not((layer0_outputs(7581)) xor (layer0_outputs(1533)));
    outputs(4938) <= not((layer0_outputs(2621)) or (layer0_outputs(6822)));
    outputs(4939) <= layer0_outputs(7972);
    outputs(4940) <= not(layer0_outputs(6805));
    outputs(4941) <= not((layer0_outputs(76)) xor (layer0_outputs(639)));
    outputs(4942) <= not(layer0_outputs(2128));
    outputs(4943) <= not(layer0_outputs(679));
    outputs(4944) <= (layer0_outputs(20)) and not (layer0_outputs(5504));
    outputs(4945) <= (layer0_outputs(9973)) or (layer0_outputs(1400));
    outputs(4946) <= not((layer0_outputs(405)) xor (layer0_outputs(8507)));
    outputs(4947) <= not(layer0_outputs(4941));
    outputs(4948) <= '0';
    outputs(4949) <= not((layer0_outputs(4676)) or (layer0_outputs(6436)));
    outputs(4950) <= (layer0_outputs(158)) xor (layer0_outputs(3558));
    outputs(4951) <= (layer0_outputs(9137)) and not (layer0_outputs(647));
    outputs(4952) <= layer0_outputs(4624);
    outputs(4953) <= not(layer0_outputs(8076));
    outputs(4954) <= layer0_outputs(1074);
    outputs(4955) <= not(layer0_outputs(5072));
    outputs(4956) <= not((layer0_outputs(2265)) xor (layer0_outputs(2421)));
    outputs(4957) <= layer0_outputs(986);
    outputs(4958) <= not(layer0_outputs(4476));
    outputs(4959) <= not((layer0_outputs(4556)) xor (layer0_outputs(523)));
    outputs(4960) <= (layer0_outputs(2442)) and (layer0_outputs(7735));
    outputs(4961) <= not(layer0_outputs(2736));
    outputs(4962) <= not(layer0_outputs(10139));
    outputs(4963) <= not((layer0_outputs(6377)) xor (layer0_outputs(8638)));
    outputs(4964) <= (layer0_outputs(5972)) and not (layer0_outputs(9325));
    outputs(4965) <= (layer0_outputs(8299)) xor (layer0_outputs(7691));
    outputs(4966) <= (layer0_outputs(9504)) xor (layer0_outputs(3584));
    outputs(4967) <= (layer0_outputs(5650)) xor (layer0_outputs(4696));
    outputs(4968) <= layer0_outputs(8753);
    outputs(4969) <= not(layer0_outputs(7552));
    outputs(4970) <= (layer0_outputs(1860)) xor (layer0_outputs(4686));
    outputs(4971) <= not(layer0_outputs(7759));
    outputs(4972) <= not((layer0_outputs(3910)) xor (layer0_outputs(5161)));
    outputs(4973) <= not((layer0_outputs(7707)) or (layer0_outputs(5818)));
    outputs(4974) <= not((layer0_outputs(814)) or (layer0_outputs(305)));
    outputs(4975) <= (layer0_outputs(9331)) xor (layer0_outputs(4929));
    outputs(4976) <= not(layer0_outputs(1120));
    outputs(4977) <= not((layer0_outputs(2090)) or (layer0_outputs(2845)));
    outputs(4978) <= layer0_outputs(7630);
    outputs(4979) <= (layer0_outputs(6595)) and not (layer0_outputs(6636));
    outputs(4980) <= not(layer0_outputs(50)) or (layer0_outputs(5897));
    outputs(4981) <= (layer0_outputs(3432)) and not (layer0_outputs(5125));
    outputs(4982) <= (layer0_outputs(8191)) and (layer0_outputs(10064));
    outputs(4983) <= layer0_outputs(694);
    outputs(4984) <= not((layer0_outputs(5489)) or (layer0_outputs(4343)));
    outputs(4985) <= not(layer0_outputs(247));
    outputs(4986) <= not(layer0_outputs(5083));
    outputs(4987) <= layer0_outputs(2844);
    outputs(4988) <= not(layer0_outputs(4767));
    outputs(4989) <= layer0_outputs(8330);
    outputs(4990) <= (layer0_outputs(1936)) and not (layer0_outputs(6270));
    outputs(4991) <= (layer0_outputs(333)) xor (layer0_outputs(428));
    outputs(4992) <= layer0_outputs(10144);
    outputs(4993) <= layer0_outputs(10236);
    outputs(4994) <= not((layer0_outputs(3894)) xor (layer0_outputs(981)));
    outputs(4995) <= layer0_outputs(4901);
    outputs(4996) <= layer0_outputs(2378);
    outputs(4997) <= not((layer0_outputs(3536)) and (layer0_outputs(4040)));
    outputs(4998) <= layer0_outputs(6640);
    outputs(4999) <= not((layer0_outputs(1412)) xor (layer0_outputs(3042)));
    outputs(5000) <= (layer0_outputs(10180)) and not (layer0_outputs(7240));
    outputs(5001) <= not((layer0_outputs(2524)) xor (layer0_outputs(7577)));
    outputs(5002) <= not(layer0_outputs(3752)) or (layer0_outputs(6484));
    outputs(5003) <= (layer0_outputs(1933)) and not (layer0_outputs(181));
    outputs(5004) <= (layer0_outputs(2433)) and not (layer0_outputs(3034));
    outputs(5005) <= not((layer0_outputs(8259)) xor (layer0_outputs(9007)));
    outputs(5006) <= (layer0_outputs(7285)) xor (layer0_outputs(2413));
    outputs(5007) <= (layer0_outputs(4936)) and not (layer0_outputs(193));
    outputs(5008) <= not(layer0_outputs(3658));
    outputs(5009) <= (layer0_outputs(6288)) and not (layer0_outputs(8463));
    outputs(5010) <= layer0_outputs(871);
    outputs(5011) <= not((layer0_outputs(2510)) xor (layer0_outputs(6858)));
    outputs(5012) <= (layer0_outputs(2392)) and (layer0_outputs(1855));
    outputs(5013) <= not((layer0_outputs(7645)) and (layer0_outputs(10103)));
    outputs(5014) <= (layer0_outputs(4816)) and not (layer0_outputs(5567));
    outputs(5015) <= not((layer0_outputs(6206)) or (layer0_outputs(2653)));
    outputs(5016) <= not((layer0_outputs(9537)) xor (layer0_outputs(6760)));
    outputs(5017) <= not(layer0_outputs(8510));
    outputs(5018) <= layer0_outputs(4751);
    outputs(5019) <= layer0_outputs(4444);
    outputs(5020) <= not((layer0_outputs(8028)) or (layer0_outputs(3795)));
    outputs(5021) <= (layer0_outputs(4053)) or (layer0_outputs(7852));
    outputs(5022) <= (layer0_outputs(9029)) xor (layer0_outputs(9622));
    outputs(5023) <= (layer0_outputs(4619)) xor (layer0_outputs(9341));
    outputs(5024) <= layer0_outputs(1913);
    outputs(5025) <= layer0_outputs(6014);
    outputs(5026) <= (layer0_outputs(3726)) and (layer0_outputs(8676));
    outputs(5027) <= not((layer0_outputs(7233)) xor (layer0_outputs(5784)));
    outputs(5028) <= not(layer0_outputs(7758));
    outputs(5029) <= not(layer0_outputs(2963)) or (layer0_outputs(299));
    outputs(5030) <= (layer0_outputs(6201)) xor (layer0_outputs(6099));
    outputs(5031) <= not(layer0_outputs(9304));
    outputs(5032) <= (layer0_outputs(9177)) and (layer0_outputs(7404));
    outputs(5033) <= not(layer0_outputs(7659));
    outputs(5034) <= (layer0_outputs(876)) and (layer0_outputs(6934));
    outputs(5035) <= (layer0_outputs(8774)) xor (layer0_outputs(8596));
    outputs(5036) <= not(layer0_outputs(3197));
    outputs(5037) <= layer0_outputs(8801);
    outputs(5038) <= (layer0_outputs(4627)) xor (layer0_outputs(5901));
    outputs(5039) <= (layer0_outputs(6778)) and not (layer0_outputs(9459));
    outputs(5040) <= (layer0_outputs(8000)) and not (layer0_outputs(1253));
    outputs(5041) <= not(layer0_outputs(2883));
    outputs(5042) <= not(layer0_outputs(1790));
    outputs(5043) <= not((layer0_outputs(4315)) or (layer0_outputs(8567)));
    outputs(5044) <= (layer0_outputs(977)) and not (layer0_outputs(8533));
    outputs(5045) <= not(layer0_outputs(3142));
    outputs(5046) <= layer0_outputs(6224);
    outputs(5047) <= not(layer0_outputs(1126));
    outputs(5048) <= not(layer0_outputs(4504));
    outputs(5049) <= (layer0_outputs(9396)) xor (layer0_outputs(3832));
    outputs(5050) <= (layer0_outputs(5318)) and not (layer0_outputs(9446));
    outputs(5051) <= (layer0_outputs(7466)) and not (layer0_outputs(8192));
    outputs(5052) <= (layer0_outputs(845)) and (layer0_outputs(8599));
    outputs(5053) <= (layer0_outputs(6036)) and not (layer0_outputs(3829));
    outputs(5054) <= (layer0_outputs(3446)) and not (layer0_outputs(7891));
    outputs(5055) <= (layer0_outputs(7056)) xor (layer0_outputs(2614));
    outputs(5056) <= not((layer0_outputs(7950)) or (layer0_outputs(8213)));
    outputs(5057) <= not((layer0_outputs(736)) xor (layer0_outputs(3921)));
    outputs(5058) <= layer0_outputs(6131);
    outputs(5059) <= not(layer0_outputs(3004));
    outputs(5060) <= not(layer0_outputs(5600));
    outputs(5061) <= not(layer0_outputs(7281));
    outputs(5062) <= not(layer0_outputs(6739)) or (layer0_outputs(7197));
    outputs(5063) <= layer0_outputs(459);
    outputs(5064) <= layer0_outputs(6893);
    outputs(5065) <= not(layer0_outputs(645));
    outputs(5066) <= layer0_outputs(9930);
    outputs(5067) <= not((layer0_outputs(4783)) xor (layer0_outputs(686)));
    outputs(5068) <= not(layer0_outputs(2061));
    outputs(5069) <= (layer0_outputs(6731)) and not (layer0_outputs(7127));
    outputs(5070) <= (layer0_outputs(2038)) xor (layer0_outputs(3698));
    outputs(5071) <= (layer0_outputs(614)) and (layer0_outputs(7589));
    outputs(5072) <= not((layer0_outputs(4111)) or (layer0_outputs(7813)));
    outputs(5073) <= (layer0_outputs(3984)) and not (layer0_outputs(438));
    outputs(5074) <= (layer0_outputs(684)) and not (layer0_outputs(2212));
    outputs(5075) <= not((layer0_outputs(2971)) xor (layer0_outputs(6271)));
    outputs(5076) <= (layer0_outputs(1267)) and (layer0_outputs(880));
    outputs(5077) <= not(layer0_outputs(10158));
    outputs(5078) <= layer0_outputs(5008);
    outputs(5079) <= (layer0_outputs(1409)) xor (layer0_outputs(1976));
    outputs(5080) <= not(layer0_outputs(775));
    outputs(5081) <= (layer0_outputs(8197)) and not (layer0_outputs(10094));
    outputs(5082) <= (layer0_outputs(2983)) and (layer0_outputs(2741));
    outputs(5083) <= not(layer0_outputs(2240));
    outputs(5084) <= layer0_outputs(7557);
    outputs(5085) <= (layer0_outputs(2314)) and not (layer0_outputs(8364));
    outputs(5086) <= not(layer0_outputs(5458));
    outputs(5087) <= (layer0_outputs(2230)) and (layer0_outputs(648));
    outputs(5088) <= not((layer0_outputs(1382)) or (layer0_outputs(1930)));
    outputs(5089) <= not(layer0_outputs(7435));
    outputs(5090) <= layer0_outputs(2693);
    outputs(5091) <= not((layer0_outputs(4393)) or (layer0_outputs(3427)));
    outputs(5092) <= layer0_outputs(1022);
    outputs(5093) <= not(layer0_outputs(2519)) or (layer0_outputs(5279));
    outputs(5094) <= (layer0_outputs(10221)) and (layer0_outputs(4152));
    outputs(5095) <= not((layer0_outputs(8504)) or (layer0_outputs(7528)));
    outputs(5096) <= not(layer0_outputs(10131));
    outputs(5097) <= (layer0_outputs(3032)) xor (layer0_outputs(195));
    outputs(5098) <= layer0_outputs(5709);
    outputs(5099) <= (layer0_outputs(4209)) and (layer0_outputs(9407));
    outputs(5100) <= layer0_outputs(5368);
    outputs(5101) <= not(layer0_outputs(8927));
    outputs(5102) <= layer0_outputs(160);
    outputs(5103) <= not((layer0_outputs(8612)) and (layer0_outputs(8888)));
    outputs(5104) <= layer0_outputs(993);
    outputs(5105) <= (layer0_outputs(1688)) xor (layer0_outputs(637));
    outputs(5106) <= layer0_outputs(248);
    outputs(5107) <= not((layer0_outputs(2281)) or (layer0_outputs(1141)));
    outputs(5108) <= not(layer0_outputs(2503));
    outputs(5109) <= not(layer0_outputs(2974));
    outputs(5110) <= layer0_outputs(5609);
    outputs(5111) <= layer0_outputs(4389);
    outputs(5112) <= layer0_outputs(792);
    outputs(5113) <= not(layer0_outputs(1483));
    outputs(5114) <= not(layer0_outputs(5266));
    outputs(5115) <= (layer0_outputs(802)) or (layer0_outputs(2992));
    outputs(5116) <= (layer0_outputs(3583)) and (layer0_outputs(6069));
    outputs(5117) <= layer0_outputs(1870);
    outputs(5118) <= (layer0_outputs(3928)) and not (layer0_outputs(4083));
    outputs(5119) <= (layer0_outputs(8336)) xor (layer0_outputs(5791));
    outputs(5120) <= (layer0_outputs(9605)) and not (layer0_outputs(2706));
    outputs(5121) <= layer0_outputs(3754);
    outputs(5122) <= layer0_outputs(7421);
    outputs(5123) <= (layer0_outputs(1819)) xor (layer0_outputs(517));
    outputs(5124) <= (layer0_outputs(5037)) and (layer0_outputs(4079));
    outputs(5125) <= (layer0_outputs(5519)) and not (layer0_outputs(3913));
    outputs(5126) <= not(layer0_outputs(7318));
    outputs(5127) <= layer0_outputs(5830);
    outputs(5128) <= not(layer0_outputs(4202));
    outputs(5129) <= not((layer0_outputs(5347)) xor (layer0_outputs(9485)));
    outputs(5130) <= not((layer0_outputs(132)) xor (layer0_outputs(3377)));
    outputs(5131) <= layer0_outputs(9115);
    outputs(5132) <= not(layer0_outputs(4926)) or (layer0_outputs(3929));
    outputs(5133) <= (layer0_outputs(7812)) xor (layer0_outputs(2115));
    outputs(5134) <= not(layer0_outputs(3683));
    outputs(5135) <= (layer0_outputs(4466)) or (layer0_outputs(7662));
    outputs(5136) <= not((layer0_outputs(5930)) and (layer0_outputs(1910)));
    outputs(5137) <= not(layer0_outputs(615));
    outputs(5138) <= (layer0_outputs(7772)) and (layer0_outputs(5260));
    outputs(5139) <= layer0_outputs(8325);
    outputs(5140) <= (layer0_outputs(9823)) xor (layer0_outputs(3394));
    outputs(5141) <= (layer0_outputs(8686)) and not (layer0_outputs(8053));
    outputs(5142) <= (layer0_outputs(6640)) xor (layer0_outputs(4866));
    outputs(5143) <= not(layer0_outputs(3589));
    outputs(5144) <= not(layer0_outputs(159));
    outputs(5145) <= layer0_outputs(1701);
    outputs(5146) <= not(layer0_outputs(2866));
    outputs(5147) <= not(layer0_outputs(9270));
    outputs(5148) <= not(layer0_outputs(1062)) or (layer0_outputs(8283));
    outputs(5149) <= not(layer0_outputs(2419));
    outputs(5150) <= not((layer0_outputs(239)) or (layer0_outputs(4241)));
    outputs(5151) <= (layer0_outputs(708)) xor (layer0_outputs(9913));
    outputs(5152) <= not(layer0_outputs(1673));
    outputs(5153) <= layer0_outputs(6271);
    outputs(5154) <= (layer0_outputs(6024)) xor (layer0_outputs(2795));
    outputs(5155) <= not((layer0_outputs(9843)) xor (layer0_outputs(8274)));
    outputs(5156) <= not((layer0_outputs(9032)) xor (layer0_outputs(1675)));
    outputs(5157) <= not((layer0_outputs(672)) xor (layer0_outputs(6453)));
    outputs(5158) <= layer0_outputs(10076);
    outputs(5159) <= (layer0_outputs(627)) or (layer0_outputs(63));
    outputs(5160) <= (layer0_outputs(282)) xor (layer0_outputs(1603));
    outputs(5161) <= not((layer0_outputs(3230)) xor (layer0_outputs(7385)));
    outputs(5162) <= (layer0_outputs(2820)) xor (layer0_outputs(218));
    outputs(5163) <= not(layer0_outputs(335));
    outputs(5164) <= layer0_outputs(1983);
    outputs(5165) <= not(layer0_outputs(4622));
    outputs(5166) <= (layer0_outputs(9043)) xor (layer0_outputs(3525));
    outputs(5167) <= not(layer0_outputs(4368));
    outputs(5168) <= (layer0_outputs(8592)) xor (layer0_outputs(8664));
    outputs(5169) <= not(layer0_outputs(1875));
    outputs(5170) <= layer0_outputs(3307);
    outputs(5171) <= not(layer0_outputs(8097));
    outputs(5172) <= (layer0_outputs(5033)) and not (layer0_outputs(4309));
    outputs(5173) <= not((layer0_outputs(5526)) xor (layer0_outputs(5554)));
    outputs(5174) <= (layer0_outputs(66)) xor (layer0_outputs(7946));
    outputs(5175) <= not((layer0_outputs(3783)) or (layer0_outputs(1529)));
    outputs(5176) <= layer0_outputs(168);
    outputs(5177) <= not(layer0_outputs(7102));
    outputs(5178) <= layer0_outputs(6929);
    outputs(5179) <= not((layer0_outputs(6450)) xor (layer0_outputs(6660)));
    outputs(5180) <= not((layer0_outputs(9660)) xor (layer0_outputs(7632)));
    outputs(5181) <= layer0_outputs(7254);
    outputs(5182) <= not((layer0_outputs(1653)) xor (layer0_outputs(762)));
    outputs(5183) <= not(layer0_outputs(10168));
    outputs(5184) <= not((layer0_outputs(9472)) and (layer0_outputs(2623)));
    outputs(5185) <= layer0_outputs(1337);
    outputs(5186) <= not(layer0_outputs(398));
    outputs(5187) <= (layer0_outputs(3943)) or (layer0_outputs(9266));
    outputs(5188) <= (layer0_outputs(3240)) xor (layer0_outputs(246));
    outputs(5189) <= (layer0_outputs(4548)) or (layer0_outputs(201));
    outputs(5190) <= (layer0_outputs(9322)) or (layer0_outputs(6432));
    outputs(5191) <= not(layer0_outputs(4921));
    outputs(5192) <= not((layer0_outputs(484)) and (layer0_outputs(8497)));
    outputs(5193) <= layer0_outputs(6103);
    outputs(5194) <= (layer0_outputs(6452)) and not (layer0_outputs(2367));
    outputs(5195) <= not((layer0_outputs(3411)) xor (layer0_outputs(3824)));
    outputs(5196) <= (layer0_outputs(6820)) xor (layer0_outputs(2460));
    outputs(5197) <= layer0_outputs(6098);
    outputs(5198) <= not(layer0_outputs(668));
    outputs(5199) <= not(layer0_outputs(5117));
    outputs(5200) <= not(layer0_outputs(6881)) or (layer0_outputs(6290));
    outputs(5201) <= (layer0_outputs(2127)) xor (layer0_outputs(2036));
    outputs(5202) <= (layer0_outputs(5357)) xor (layer0_outputs(7658));
    outputs(5203) <= not((layer0_outputs(4566)) xor (layer0_outputs(4451)));
    outputs(5204) <= (layer0_outputs(3608)) xor (layer0_outputs(5385));
    outputs(5205) <= not((layer0_outputs(10211)) and (layer0_outputs(2114)));
    outputs(5206) <= (layer0_outputs(2228)) xor (layer0_outputs(4477));
    outputs(5207) <= not((layer0_outputs(5023)) xor (layer0_outputs(7790)));
    outputs(5208) <= not((layer0_outputs(2556)) and (layer0_outputs(4317)));
    outputs(5209) <= not(layer0_outputs(3777));
    outputs(5210) <= not((layer0_outputs(8352)) or (layer0_outputs(67)));
    outputs(5211) <= (layer0_outputs(6030)) and (layer0_outputs(4425));
    outputs(5212) <= not((layer0_outputs(7004)) or (layer0_outputs(3279)));
    outputs(5213) <= (layer0_outputs(8944)) and not (layer0_outputs(1754));
    outputs(5214) <= not((layer0_outputs(4300)) xor (layer0_outputs(4442)));
    outputs(5215) <= layer0_outputs(8734);
    outputs(5216) <= (layer0_outputs(6020)) xor (layer0_outputs(4103));
    outputs(5217) <= (layer0_outputs(8895)) xor (layer0_outputs(95));
    outputs(5218) <= not((layer0_outputs(3247)) or (layer0_outputs(5802)));
    outputs(5219) <= (layer0_outputs(52)) xor (layer0_outputs(6242));
    outputs(5220) <= layer0_outputs(7648);
    outputs(5221) <= (layer0_outputs(6452)) and (layer0_outputs(9417));
    outputs(5222) <= (layer0_outputs(5370)) or (layer0_outputs(1530));
    outputs(5223) <= not((layer0_outputs(289)) or (layer0_outputs(7032)));
    outputs(5224) <= not(layer0_outputs(3815));
    outputs(5225) <= not(layer0_outputs(7874)) or (layer0_outputs(2844));
    outputs(5226) <= (layer0_outputs(4994)) xor (layer0_outputs(959));
    outputs(5227) <= not(layer0_outputs(8380)) or (layer0_outputs(950));
    outputs(5228) <= (layer0_outputs(6151)) and not (layer0_outputs(6390));
    outputs(5229) <= not((layer0_outputs(1415)) xor (layer0_outputs(5331)));
    outputs(5230) <= (layer0_outputs(317)) xor (layer0_outputs(1915));
    outputs(5231) <= not(layer0_outputs(10067));
    outputs(5232) <= (layer0_outputs(8602)) and not (layer0_outputs(8219));
    outputs(5233) <= not((layer0_outputs(7347)) xor (layer0_outputs(8030)));
    outputs(5234) <= (layer0_outputs(4023)) xor (layer0_outputs(2267));
    outputs(5235) <= (layer0_outputs(7426)) and not (layer0_outputs(7414));
    outputs(5236) <= not((layer0_outputs(8009)) or (layer0_outputs(90)));
    outputs(5237) <= layer0_outputs(7539);
    outputs(5238) <= layer0_outputs(3296);
    outputs(5239) <= not((layer0_outputs(5015)) and (layer0_outputs(756)));
    outputs(5240) <= (layer0_outputs(1980)) xor (layer0_outputs(5388));
    outputs(5241) <= layer0_outputs(3169);
    outputs(5242) <= not(layer0_outputs(3399));
    outputs(5243) <= not(layer0_outputs(7493));
    outputs(5244) <= (layer0_outputs(4431)) xor (layer0_outputs(6127));
    outputs(5245) <= (layer0_outputs(7752)) xor (layer0_outputs(4490));
    outputs(5246) <= not(layer0_outputs(9249));
    outputs(5247) <= (layer0_outputs(9963)) and not (layer0_outputs(7119));
    outputs(5248) <= (layer0_outputs(8004)) xor (layer0_outputs(441));
    outputs(5249) <= not((layer0_outputs(5779)) or (layer0_outputs(5845)));
    outputs(5250) <= layer0_outputs(6233);
    outputs(5251) <= (layer0_outputs(61)) and not (layer0_outputs(4546));
    outputs(5252) <= (layer0_outputs(10152)) xor (layer0_outputs(4511));
    outputs(5253) <= not(layer0_outputs(2698)) or (layer0_outputs(3208));
    outputs(5254) <= not(layer0_outputs(6510)) or (layer0_outputs(1390));
    outputs(5255) <= not(layer0_outputs(7225)) or (layer0_outputs(4981));
    outputs(5256) <= not(layer0_outputs(5893));
    outputs(5257) <= not((layer0_outputs(8635)) and (layer0_outputs(5000)));
    outputs(5258) <= not(layer0_outputs(5825));
    outputs(5259) <= not((layer0_outputs(1914)) and (layer0_outputs(8025)));
    outputs(5260) <= (layer0_outputs(8218)) or (layer0_outputs(4411));
    outputs(5261) <= not(layer0_outputs(1429));
    outputs(5262) <= not((layer0_outputs(8138)) xor (layer0_outputs(9965)));
    outputs(5263) <= not(layer0_outputs(1304));
    outputs(5264) <= not(layer0_outputs(202)) or (layer0_outputs(4579));
    outputs(5265) <= not(layer0_outputs(3979));
    outputs(5266) <= (layer0_outputs(1333)) and not (layer0_outputs(6677));
    outputs(5267) <= not(layer0_outputs(6538));
    outputs(5268) <= not(layer0_outputs(5811));
    outputs(5269) <= not(layer0_outputs(6389));
    outputs(5270) <= not(layer0_outputs(4703));
    outputs(5271) <= (layer0_outputs(122)) xor (layer0_outputs(899));
    outputs(5272) <= (layer0_outputs(3463)) and not (layer0_outputs(9858));
    outputs(5273) <= not(layer0_outputs(9526));
    outputs(5274) <= not(layer0_outputs(10179)) or (layer0_outputs(9087));
    outputs(5275) <= (layer0_outputs(2371)) or (layer0_outputs(2420));
    outputs(5276) <= not(layer0_outputs(8371)) or (layer0_outputs(5930));
    outputs(5277) <= not(layer0_outputs(646)) or (layer0_outputs(1630));
    outputs(5278) <= (layer0_outputs(1361)) and (layer0_outputs(2339));
    outputs(5279) <= not(layer0_outputs(8245)) or (layer0_outputs(8193));
    outputs(5280) <= (layer0_outputs(2925)) and not (layer0_outputs(9892));
    outputs(5281) <= (layer0_outputs(3681)) and not (layer0_outputs(3051));
    outputs(5282) <= not((layer0_outputs(83)) xor (layer0_outputs(8350)));
    outputs(5283) <= not((layer0_outputs(8531)) or (layer0_outputs(7873)));
    outputs(5284) <= (layer0_outputs(2232)) and not (layer0_outputs(533));
    outputs(5285) <= (layer0_outputs(1572)) xor (layer0_outputs(3351));
    outputs(5286) <= (layer0_outputs(6958)) and not (layer0_outputs(8131));
    outputs(5287) <= layer0_outputs(5437);
    outputs(5288) <= layer0_outputs(7055);
    outputs(5289) <= layer0_outputs(5766);
    outputs(5290) <= (layer0_outputs(7773)) or (layer0_outputs(4430));
    outputs(5291) <= (layer0_outputs(4013)) xor (layer0_outputs(690));
    outputs(5292) <= layer0_outputs(6647);
    outputs(5293) <= (layer0_outputs(1990)) xor (layer0_outputs(7712));
    outputs(5294) <= (layer0_outputs(3836)) xor (layer0_outputs(7114));
    outputs(5295) <= not((layer0_outputs(470)) or (layer0_outputs(7451)));
    outputs(5296) <= not((layer0_outputs(2790)) and (layer0_outputs(313)));
    outputs(5297) <= not((layer0_outputs(3534)) xor (layer0_outputs(4916)));
    outputs(5298) <= layer0_outputs(629);
    outputs(5299) <= layer0_outputs(2662);
    outputs(5300) <= not((layer0_outputs(10230)) and (layer0_outputs(1822)));
    outputs(5301) <= not((layer0_outputs(5996)) xor (layer0_outputs(9058)));
    outputs(5302) <= (layer0_outputs(9294)) and not (layer0_outputs(4449));
    outputs(5303) <= not((layer0_outputs(8822)) and (layer0_outputs(2152)));
    outputs(5304) <= not(layer0_outputs(6523)) or (layer0_outputs(1828));
    outputs(5305) <= layer0_outputs(8184);
    outputs(5306) <= layer0_outputs(8223);
    outputs(5307) <= (layer0_outputs(256)) and not (layer0_outputs(3386));
    outputs(5308) <= not(layer0_outputs(8711)) or (layer0_outputs(9945));
    outputs(5309) <= layer0_outputs(8208);
    outputs(5310) <= not(layer0_outputs(491)) or (layer0_outputs(8671));
    outputs(5311) <= (layer0_outputs(1139)) xor (layer0_outputs(3936));
    outputs(5312) <= layer0_outputs(793);
    outputs(5313) <= (layer0_outputs(8364)) xor (layer0_outputs(1362));
    outputs(5314) <= not((layer0_outputs(2567)) or (layer0_outputs(6553)));
    outputs(5315) <= not(layer0_outputs(5583));
    outputs(5316) <= (layer0_outputs(7487)) and not (layer0_outputs(4945));
    outputs(5317) <= (layer0_outputs(6481)) xor (layer0_outputs(6532));
    outputs(5318) <= (layer0_outputs(2882)) xor (layer0_outputs(2070));
    outputs(5319) <= layer0_outputs(1463);
    outputs(5320) <= not(layer0_outputs(2916)) or (layer0_outputs(4464));
    outputs(5321) <= (layer0_outputs(10080)) xor (layer0_outputs(1466));
    outputs(5322) <= layer0_outputs(1882);
    outputs(5323) <= layer0_outputs(7453);
    outputs(5324) <= '1';
    outputs(5325) <= layer0_outputs(5403);
    outputs(5326) <= (layer0_outputs(7434)) xor (layer0_outputs(8095));
    outputs(5327) <= (layer0_outputs(3003)) xor (layer0_outputs(5384));
    outputs(5328) <= layer0_outputs(4420);
    outputs(5329) <= not(layer0_outputs(8767));
    outputs(5330) <= not((layer0_outputs(850)) and (layer0_outputs(1339)));
    outputs(5331) <= not((layer0_outputs(1845)) xor (layer0_outputs(9573)));
    outputs(5332) <= not(layer0_outputs(6054));
    outputs(5333) <= layer0_outputs(4850);
    outputs(5334) <= not(layer0_outputs(8323));
    outputs(5335) <= not(layer0_outputs(3509));
    outputs(5336) <= (layer0_outputs(6609)) or (layer0_outputs(697));
    outputs(5337) <= (layer0_outputs(1939)) and not (layer0_outputs(3615));
    outputs(5338) <= not(layer0_outputs(2042));
    outputs(5339) <= not(layer0_outputs(7479));
    outputs(5340) <= layer0_outputs(7975);
    outputs(5341) <= (layer0_outputs(5343)) and not (layer0_outputs(1727));
    outputs(5342) <= not(layer0_outputs(5222));
    outputs(5343) <= not((layer0_outputs(1650)) xor (layer0_outputs(658)));
    outputs(5344) <= layer0_outputs(1481);
    outputs(5345) <= (layer0_outputs(6255)) and (layer0_outputs(9825));
    outputs(5346) <= layer0_outputs(3602);
    outputs(5347) <= layer0_outputs(9002);
    outputs(5348) <= layer0_outputs(2654);
    outputs(5349) <= (layer0_outputs(1135)) and not (layer0_outputs(1028));
    outputs(5350) <= not((layer0_outputs(8280)) xor (layer0_outputs(5988)));
    outputs(5351) <= not((layer0_outputs(1686)) xor (layer0_outputs(5980)));
    outputs(5352) <= not(layer0_outputs(7346)) or (layer0_outputs(6317));
    outputs(5353) <= not((layer0_outputs(10087)) xor (layer0_outputs(7182)));
    outputs(5354) <= not((layer0_outputs(6757)) xor (layer0_outputs(7457)));
    outputs(5355) <= layer0_outputs(3405);
    outputs(5356) <= not(layer0_outputs(9736)) or (layer0_outputs(847));
    outputs(5357) <= not(layer0_outputs(2962));
    outputs(5358) <= not(layer0_outputs(1951)) or (layer0_outputs(1239));
    outputs(5359) <= (layer0_outputs(6661)) xor (layer0_outputs(3784));
    outputs(5360) <= not(layer0_outputs(9869)) or (layer0_outputs(8928));
    outputs(5361) <= not(layer0_outputs(6743));
    outputs(5362) <= layer0_outputs(5231);
    outputs(5363) <= not((layer0_outputs(7788)) and (layer0_outputs(10109)));
    outputs(5364) <= not(layer0_outputs(5726));
    outputs(5365) <= (layer0_outputs(5095)) or (layer0_outputs(4847));
    outputs(5366) <= layer0_outputs(3867);
    outputs(5367) <= not((layer0_outputs(9023)) xor (layer0_outputs(9314)));
    outputs(5368) <= not((layer0_outputs(579)) or (layer0_outputs(7930)));
    outputs(5369) <= not(layer0_outputs(890));
    outputs(5370) <= (layer0_outputs(3992)) and not (layer0_outputs(1810));
    outputs(5371) <= (layer0_outputs(9378)) xor (layer0_outputs(2793));
    outputs(5372) <= not((layer0_outputs(8348)) and (layer0_outputs(279)));
    outputs(5373) <= (layer0_outputs(9801)) and (layer0_outputs(9674));
    outputs(5374) <= not(layer0_outputs(10073)) or (layer0_outputs(739));
    outputs(5375) <= not(layer0_outputs(8535)) or (layer0_outputs(7321));
    outputs(5376) <= not(layer0_outputs(2996)) or (layer0_outputs(8863));
    outputs(5377) <= not((layer0_outputs(9455)) and (layer0_outputs(8994)));
    outputs(5378) <= not(layer0_outputs(8506));
    outputs(5379) <= layer0_outputs(5138);
    outputs(5380) <= layer0_outputs(9606);
    outputs(5381) <= (layer0_outputs(4843)) xor (layer0_outputs(6129));
    outputs(5382) <= not((layer0_outputs(766)) xor (layer0_outputs(9022)));
    outputs(5383) <= (layer0_outputs(3219)) xor (layer0_outputs(7724));
    outputs(5384) <= not(layer0_outputs(495));
    outputs(5385) <= not(layer0_outputs(4590));
    outputs(5386) <= layer0_outputs(3640);
    outputs(5387) <= not(layer0_outputs(1028));
    outputs(5388) <= (layer0_outputs(1864)) xor (layer0_outputs(8574));
    outputs(5389) <= not((layer0_outputs(3285)) xor (layer0_outputs(1332)));
    outputs(5390) <= (layer0_outputs(3719)) or (layer0_outputs(3347));
    outputs(5391) <= not(layer0_outputs(8339));
    outputs(5392) <= not(layer0_outputs(9390));
    outputs(5393) <= not(layer0_outputs(4499)) or (layer0_outputs(3233));
    outputs(5394) <= (layer0_outputs(5643)) or (layer0_outputs(3506));
    outputs(5395) <= not(layer0_outputs(493));
    outputs(5396) <= not(layer0_outputs(4862));
    outputs(5397) <= (layer0_outputs(3929)) or (layer0_outputs(9979));
    outputs(5398) <= not(layer0_outputs(6263));
    outputs(5399) <= layer0_outputs(3959);
    outputs(5400) <= not((layer0_outputs(2696)) xor (layer0_outputs(6324)));
    outputs(5401) <= (layer0_outputs(2618)) or (layer0_outputs(7974));
    outputs(5402) <= not(layer0_outputs(7181));
    outputs(5403) <= not((layer0_outputs(4737)) xor (layer0_outputs(8358)));
    outputs(5404) <= not(layer0_outputs(3011));
    outputs(5405) <= layer0_outputs(3498);
    outputs(5406) <= not((layer0_outputs(1499)) xor (layer0_outputs(8397)));
    outputs(5407) <= not((layer0_outputs(1156)) xor (layer0_outputs(6535)));
    outputs(5408) <= (layer0_outputs(696)) xor (layer0_outputs(3107));
    outputs(5409) <= not(layer0_outputs(9448));
    outputs(5410) <= (layer0_outputs(3038)) xor (layer0_outputs(6753));
    outputs(5411) <= (layer0_outputs(5182)) or (layer0_outputs(1701));
    outputs(5412) <= layer0_outputs(8130);
    outputs(5413) <= not(layer0_outputs(1927));
    outputs(5414) <= (layer0_outputs(5103)) and not (layer0_outputs(8850));
    outputs(5415) <= (layer0_outputs(481)) or (layer0_outputs(5424));
    outputs(5416) <= (layer0_outputs(1372)) xor (layer0_outputs(8514));
    outputs(5417) <= not(layer0_outputs(121));
    outputs(5418) <= not(layer0_outputs(7502));
    outputs(5419) <= not(layer0_outputs(2311)) or (layer0_outputs(5057));
    outputs(5420) <= (layer0_outputs(4810)) or (layer0_outputs(6530));
    outputs(5421) <= not(layer0_outputs(4483));
    outputs(5422) <= (layer0_outputs(450)) xor (layer0_outputs(10097));
    outputs(5423) <= not((layer0_outputs(10204)) xor (layer0_outputs(3955)));
    outputs(5424) <= layer0_outputs(4244);
    outputs(5425) <= (layer0_outputs(9621)) and not (layer0_outputs(9025));
    outputs(5426) <= not(layer0_outputs(9655));
    outputs(5427) <= layer0_outputs(6249);
    outputs(5428) <= not(layer0_outputs(2987)) or (layer0_outputs(8757));
    outputs(5429) <= not(layer0_outputs(4560));
    outputs(5430) <= not((layer0_outputs(6990)) or (layer0_outputs(4785)));
    outputs(5431) <= (layer0_outputs(1093)) and not (layer0_outputs(2535));
    outputs(5432) <= not((layer0_outputs(4522)) and (layer0_outputs(903)));
    outputs(5433) <= layer0_outputs(9787);
    outputs(5434) <= not(layer0_outputs(8087));
    outputs(5435) <= not(layer0_outputs(3227));
    outputs(5436) <= (layer0_outputs(1435)) xor (layer0_outputs(7220));
    outputs(5437) <= (layer0_outputs(4782)) and not (layer0_outputs(7896));
    outputs(5438) <= not(layer0_outputs(8717));
    outputs(5439) <= layer0_outputs(3542);
    outputs(5440) <= layer0_outputs(3767);
    outputs(5441) <= (layer0_outputs(8585)) and not (layer0_outputs(7510));
    outputs(5442) <= not(layer0_outputs(123)) or (layer0_outputs(9863));
    outputs(5443) <= not(layer0_outputs(4311));
    outputs(5444) <= (layer0_outputs(1402)) xor (layer0_outputs(5979));
    outputs(5445) <= not((layer0_outputs(9011)) xor (layer0_outputs(7648)));
    outputs(5446) <= layer0_outputs(7919);
    outputs(5447) <= not(layer0_outputs(927));
    outputs(5448) <= not(layer0_outputs(3057));
    outputs(5449) <= not(layer0_outputs(1328));
    outputs(5450) <= (layer0_outputs(8752)) or (layer0_outputs(7837));
    outputs(5451) <= (layer0_outputs(3348)) and not (layer0_outputs(2726));
    outputs(5452) <= not(layer0_outputs(2292));
    outputs(5453) <= layer0_outputs(8041);
    outputs(5454) <= not((layer0_outputs(363)) or (layer0_outputs(6615)));
    outputs(5455) <= layer0_outputs(8001);
    outputs(5456) <= not((layer0_outputs(6650)) or (layer0_outputs(2651)));
    outputs(5457) <= layer0_outputs(9306);
    outputs(5458) <= layer0_outputs(813);
    outputs(5459) <= (layer0_outputs(1025)) xor (layer0_outputs(4024));
    outputs(5460) <= not(layer0_outputs(7894));
    outputs(5461) <= (layer0_outputs(6839)) and (layer0_outputs(4668));
    outputs(5462) <= not((layer0_outputs(2191)) xor (layer0_outputs(2794)));
    outputs(5463) <= layer0_outputs(545);
    outputs(5464) <= not((layer0_outputs(4304)) or (layer0_outputs(723)));
    outputs(5465) <= (layer0_outputs(4789)) and not (layer0_outputs(3665));
    outputs(5466) <= layer0_outputs(5415);
    outputs(5467) <= not(layer0_outputs(7742)) or (layer0_outputs(9010));
    outputs(5468) <= not((layer0_outputs(7135)) xor (layer0_outputs(1670)));
    outputs(5469) <= (layer0_outputs(2096)) xor (layer0_outputs(6594));
    outputs(5470) <= not((layer0_outputs(6585)) xor (layer0_outputs(4440)));
    outputs(5471) <= not(layer0_outputs(4108));
    outputs(5472) <= not((layer0_outputs(2059)) or (layer0_outputs(8098)));
    outputs(5473) <= layer0_outputs(4038);
    outputs(5474) <= not(layer0_outputs(9725)) or (layer0_outputs(8070));
    outputs(5475) <= (layer0_outputs(4495)) xor (layer0_outputs(4326));
    outputs(5476) <= layer0_outputs(5527);
    outputs(5477) <= not(layer0_outputs(1702));
    outputs(5478) <= not(layer0_outputs(6922));
    outputs(5479) <= not((layer0_outputs(3388)) xor (layer0_outputs(3581)));
    outputs(5480) <= not(layer0_outputs(3940));
    outputs(5481) <= not(layer0_outputs(2455));
    outputs(5482) <= layer0_outputs(6373);
    outputs(5483) <= not(layer0_outputs(6671));
    outputs(5484) <= not((layer0_outputs(5765)) xor (layer0_outputs(3974)));
    outputs(5485) <= layer0_outputs(1846);
    outputs(5486) <= not((layer0_outputs(7986)) xor (layer0_outputs(5763)));
    outputs(5487) <= (layer0_outputs(1322)) or (layer0_outputs(1121));
    outputs(5488) <= not(layer0_outputs(890));
    outputs(5489) <= not((layer0_outputs(8804)) and (layer0_outputs(6909)));
    outputs(5490) <= (layer0_outputs(5941)) and not (layer0_outputs(7333));
    outputs(5491) <= not(layer0_outputs(8982));
    outputs(5492) <= (layer0_outputs(8215)) xor (layer0_outputs(2020));
    outputs(5493) <= (layer0_outputs(6883)) and not (layer0_outputs(5764));
    outputs(5494) <= (layer0_outputs(7418)) and not (layer0_outputs(6685));
    outputs(5495) <= layer0_outputs(9825);
    outputs(5496) <= not((layer0_outputs(4001)) or (layer0_outputs(4860)));
    outputs(5497) <= not((layer0_outputs(7450)) and (layer0_outputs(8418)));
    outputs(5498) <= not(layer0_outputs(6588));
    outputs(5499) <= not(layer0_outputs(563)) or (layer0_outputs(3311));
    outputs(5500) <= not(layer0_outputs(6634)) or (layer0_outputs(2508));
    outputs(5501) <= not(layer0_outputs(2973)) or (layer0_outputs(5606));
    outputs(5502) <= (layer0_outputs(7920)) xor (layer0_outputs(9860));
    outputs(5503) <= not(layer0_outputs(6401));
    outputs(5504) <= layer0_outputs(9724);
    outputs(5505) <= layer0_outputs(1531);
    outputs(5506) <= (layer0_outputs(5610)) xor (layer0_outputs(2462));
    outputs(5507) <= not((layer0_outputs(753)) xor (layer0_outputs(2144)));
    outputs(5508) <= (layer0_outputs(1614)) xor (layer0_outputs(8074));
    outputs(5509) <= layer0_outputs(9993);
    outputs(5510) <= layer0_outputs(1956);
    outputs(5511) <= layer0_outputs(4563);
    outputs(5512) <= (layer0_outputs(6238)) and not (layer0_outputs(8601));
    outputs(5513) <= not(layer0_outputs(7432));
    outputs(5514) <= (layer0_outputs(2889)) xor (layer0_outputs(4343));
    outputs(5515) <= not(layer0_outputs(6502)) or (layer0_outputs(1123));
    outputs(5516) <= layer0_outputs(8522);
    outputs(5517) <= (layer0_outputs(702)) and (layer0_outputs(7830));
    outputs(5518) <= not(layer0_outputs(9453));
    outputs(5519) <= not(layer0_outputs(5667)) or (layer0_outputs(1380));
    outputs(5520) <= (layer0_outputs(5299)) xor (layer0_outputs(1013));
    outputs(5521) <= (layer0_outputs(8571)) xor (layer0_outputs(10102));
    outputs(5522) <= not((layer0_outputs(3100)) xor (layer0_outputs(2559)));
    outputs(5523) <= (layer0_outputs(4395)) xor (layer0_outputs(2335));
    outputs(5524) <= (layer0_outputs(7575)) and (layer0_outputs(3193));
    outputs(5525) <= (layer0_outputs(4752)) xor (layer0_outputs(1906));
    outputs(5526) <= (layer0_outputs(4919)) or (layer0_outputs(1832));
    outputs(5527) <= not((layer0_outputs(7337)) xor (layer0_outputs(7588)));
    outputs(5528) <= not(layer0_outputs(8837)) or (layer0_outputs(1977));
    outputs(5529) <= layer0_outputs(8742);
    outputs(5530) <= not(layer0_outputs(7467));
    outputs(5531) <= not(layer0_outputs(9533)) or (layer0_outputs(9682));
    outputs(5532) <= not(layer0_outputs(9928));
    outputs(5533) <= not((layer0_outputs(4826)) xor (layer0_outputs(10231)));
    outputs(5534) <= not(layer0_outputs(8324)) or (layer0_outputs(2099));
    outputs(5535) <= (layer0_outputs(1251)) and not (layer0_outputs(9614));
    outputs(5536) <= (layer0_outputs(3492)) xor (layer0_outputs(1706));
    outputs(5537) <= (layer0_outputs(3755)) xor (layer0_outputs(3568));
    outputs(5538) <= (layer0_outputs(1616)) and (layer0_outputs(8345));
    outputs(5539) <= (layer0_outputs(8342)) xor (layer0_outputs(3835));
    outputs(5540) <= '1';
    outputs(5541) <= (layer0_outputs(8660)) and (layer0_outputs(1965));
    outputs(5542) <= layer0_outputs(6321);
    outputs(5543) <= not((layer0_outputs(697)) xor (layer0_outputs(4014)));
    outputs(5544) <= (layer0_outputs(5815)) and (layer0_outputs(5634));
    outputs(5545) <= (layer0_outputs(7886)) xor (layer0_outputs(6019));
    outputs(5546) <= (layer0_outputs(7884)) xor (layer0_outputs(25));
    outputs(5547) <= not(layer0_outputs(675));
    outputs(5548) <= not(layer0_outputs(3159));
    outputs(5549) <= not((layer0_outputs(3532)) xor (layer0_outputs(7678)));
    outputs(5550) <= layer0_outputs(3989);
    outputs(5551) <= not(layer0_outputs(2634));
    outputs(5552) <= not((layer0_outputs(9972)) xor (layer0_outputs(235)));
    outputs(5553) <= layer0_outputs(4240);
    outputs(5554) <= layer0_outputs(9802);
    outputs(5555) <= not(layer0_outputs(6193));
    outputs(5556) <= not((layer0_outputs(10234)) or (layer0_outputs(8101)));
    outputs(5557) <= not((layer0_outputs(881)) xor (layer0_outputs(4040)));
    outputs(5558) <= (layer0_outputs(7616)) and not (layer0_outputs(893));
    outputs(5559) <= layer0_outputs(3901);
    outputs(5560) <= not(layer0_outputs(4309));
    outputs(5561) <= (layer0_outputs(6610)) and not (layer0_outputs(4862));
    outputs(5562) <= (layer0_outputs(3789)) xor (layer0_outputs(8728));
    outputs(5563) <= layer0_outputs(6932);
    outputs(5564) <= not(layer0_outputs(7479));
    outputs(5565) <= not(layer0_outputs(8240));
    outputs(5566) <= not(layer0_outputs(7961));
    outputs(5567) <= not((layer0_outputs(9183)) xor (layer0_outputs(6797)));
    outputs(5568) <= not(layer0_outputs(5656));
    outputs(5569) <= layer0_outputs(6312);
    outputs(5570) <= not((layer0_outputs(3514)) and (layer0_outputs(3668)));
    outputs(5571) <= layer0_outputs(1834);
    outputs(5572) <= (layer0_outputs(4047)) or (layer0_outputs(5722));
    outputs(5573) <= (layer0_outputs(6843)) xor (layer0_outputs(3983));
    outputs(5574) <= not(layer0_outputs(32));
    outputs(5575) <= not(layer0_outputs(7532));
    outputs(5576) <= (layer0_outputs(8089)) or (layer0_outputs(5158));
    outputs(5577) <= not(layer0_outputs(8033));
    outputs(5578) <= not((layer0_outputs(3896)) and (layer0_outputs(302)));
    outputs(5579) <= (layer0_outputs(296)) or (layer0_outputs(3249));
    outputs(5580) <= (layer0_outputs(4533)) and not (layer0_outputs(8921));
    outputs(5581) <= not(layer0_outputs(4164)) or (layer0_outputs(5903));
    outputs(5582) <= not((layer0_outputs(3920)) xor (layer0_outputs(2094)));
    outputs(5583) <= not(layer0_outputs(3896)) or (layer0_outputs(9136));
    outputs(5584) <= layer0_outputs(5195);
    outputs(5585) <= (layer0_outputs(1841)) or (layer0_outputs(5919));
    outputs(5586) <= not((layer0_outputs(4488)) xor (layer0_outputs(6354)));
    outputs(5587) <= layer0_outputs(9894);
    outputs(5588) <= layer0_outputs(1711);
    outputs(5589) <= not((layer0_outputs(3841)) or (layer0_outputs(10236)));
    outputs(5590) <= not((layer0_outputs(4275)) xor (layer0_outputs(6155)));
    outputs(5591) <= (layer0_outputs(4362)) xor (layer0_outputs(3055));
    outputs(5592) <= (layer0_outputs(3480)) xor (layer0_outputs(9478));
    outputs(5593) <= not(layer0_outputs(8157));
    outputs(5594) <= not(layer0_outputs(2652)) or (layer0_outputs(5651));
    outputs(5595) <= not(layer0_outputs(4812));
    outputs(5596) <= not((layer0_outputs(6598)) or (layer0_outputs(4189)));
    outputs(5597) <= layer0_outputs(5266);
    outputs(5598) <= (layer0_outputs(1620)) xor (layer0_outputs(5509));
    outputs(5599) <= not(layer0_outputs(9999));
    outputs(5600) <= (layer0_outputs(8044)) or (layer0_outputs(1957));
    outputs(5601) <= layer0_outputs(908);
    outputs(5602) <= (layer0_outputs(43)) and not (layer0_outputs(9467));
    outputs(5603) <= (layer0_outputs(5164)) and not (layer0_outputs(9786));
    outputs(5604) <= not((layer0_outputs(2077)) xor (layer0_outputs(1132)));
    outputs(5605) <= layer0_outputs(1273);
    outputs(5606) <= (layer0_outputs(4246)) xor (layer0_outputs(6199));
    outputs(5607) <= not((layer0_outputs(2482)) xor (layer0_outputs(9575)));
    outputs(5608) <= not(layer0_outputs(3861)) or (layer0_outputs(4930));
    outputs(5609) <= not((layer0_outputs(3060)) or (layer0_outputs(7054)));
    outputs(5610) <= (layer0_outputs(8579)) xor (layer0_outputs(3332));
    outputs(5611) <= layer0_outputs(8571);
    outputs(5612) <= (layer0_outputs(2102)) and (layer0_outputs(5071));
    outputs(5613) <= (layer0_outputs(2683)) xor (layer0_outputs(5635));
    outputs(5614) <= layer0_outputs(8475);
    outputs(5615) <= layer0_outputs(158);
    outputs(5616) <= not(layer0_outputs(3516));
    outputs(5617) <= not(layer0_outputs(3686));
    outputs(5618) <= (layer0_outputs(4129)) xor (layer0_outputs(7771));
    outputs(5619) <= not(layer0_outputs(5276));
    outputs(5620) <= not(layer0_outputs(8818)) or (layer0_outputs(7756));
    outputs(5621) <= (layer0_outputs(6483)) xor (layer0_outputs(9916));
    outputs(5622) <= not(layer0_outputs(1959));
    outputs(5623) <= not(layer0_outputs(4829)) or (layer0_outputs(5024));
    outputs(5624) <= not(layer0_outputs(10032));
    outputs(5625) <= layer0_outputs(6134);
    outputs(5626) <= not((layer0_outputs(5358)) xor (layer0_outputs(6609)));
    outputs(5627) <= layer0_outputs(781);
    outputs(5628) <= (layer0_outputs(8075)) and not (layer0_outputs(7584));
    outputs(5629) <= not((layer0_outputs(3773)) xor (layer0_outputs(1084)));
    outputs(5630) <= (layer0_outputs(2426)) or (layer0_outputs(7542));
    outputs(5631) <= (layer0_outputs(10235)) and not (layer0_outputs(5101));
    outputs(5632) <= not(layer0_outputs(4346));
    outputs(5633) <= not((layer0_outputs(1277)) xor (layer0_outputs(5281)));
    outputs(5634) <= not(layer0_outputs(7073)) or (layer0_outputs(6222));
    outputs(5635) <= (layer0_outputs(6907)) xor (layer0_outputs(4516));
    outputs(5636) <= not((layer0_outputs(7898)) xor (layer0_outputs(8534)));
    outputs(5637) <= not(layer0_outputs(6829));
    outputs(5638) <= (layer0_outputs(8761)) or (layer0_outputs(7620));
    outputs(5639) <= not(layer0_outputs(2940));
    outputs(5640) <= layer0_outputs(4762);
    outputs(5641) <= (layer0_outputs(6178)) xor (layer0_outputs(7338));
    outputs(5642) <= not(layer0_outputs(1762));
    outputs(5643) <= (layer0_outputs(7393)) xor (layer0_outputs(6468));
    outputs(5644) <= not(layer0_outputs(4812)) or (layer0_outputs(3350));
    outputs(5645) <= layer0_outputs(814);
    outputs(5646) <= not(layer0_outputs(4190));
    outputs(5647) <= not((layer0_outputs(5810)) xor (layer0_outputs(5328)));
    outputs(5648) <= (layer0_outputs(6308)) xor (layer0_outputs(5358));
    outputs(5649) <= not((layer0_outputs(2190)) or (layer0_outputs(857)));
    outputs(5650) <= (layer0_outputs(2348)) xor (layer0_outputs(8214));
    outputs(5651) <= layer0_outputs(4624);
    outputs(5652) <= not((layer0_outputs(22)) xor (layer0_outputs(7081)));
    outputs(5653) <= (layer0_outputs(5374)) xor (layer0_outputs(7491));
    outputs(5654) <= (layer0_outputs(5344)) or (layer0_outputs(9257));
    outputs(5655) <= layer0_outputs(6524);
    outputs(5656) <= not(layer0_outputs(2954)) or (layer0_outputs(6224));
    outputs(5657) <= not(layer0_outputs(2994));
    outputs(5658) <= not((layer0_outputs(6306)) xor (layer0_outputs(7771)));
    outputs(5659) <= (layer0_outputs(6225)) and not (layer0_outputs(6745));
    outputs(5660) <= (layer0_outputs(4545)) and not (layer0_outputs(6447));
    outputs(5661) <= (layer0_outputs(7397)) and not (layer0_outputs(2761));
    outputs(5662) <= not(layer0_outputs(4646));
    outputs(5663) <= (layer0_outputs(5551)) xor (layer0_outputs(6335));
    outputs(5664) <= not((layer0_outputs(8481)) xor (layer0_outputs(8848)));
    outputs(5665) <= not((layer0_outputs(9768)) xor (layer0_outputs(8305)));
    outputs(5666) <= layer0_outputs(4515);
    outputs(5667) <= (layer0_outputs(5955)) or (layer0_outputs(7348));
    outputs(5668) <= layer0_outputs(7264);
    outputs(5669) <= not((layer0_outputs(1563)) and (layer0_outputs(6632)));
    outputs(5670) <= not((layer0_outputs(2849)) xor (layer0_outputs(598)));
    outputs(5671) <= layer0_outputs(3689);
    outputs(5672) <= (layer0_outputs(9985)) and (layer0_outputs(7778));
    outputs(5673) <= not((layer0_outputs(8735)) xor (layer0_outputs(3501)));
    outputs(5674) <= layer0_outputs(4229);
    outputs(5675) <= (layer0_outputs(1295)) xor (layer0_outputs(2813));
    outputs(5676) <= layer0_outputs(4196);
    outputs(5677) <= (layer0_outputs(171)) or (layer0_outputs(8115));
    outputs(5678) <= not(layer0_outputs(8399));
    outputs(5679) <= not(layer0_outputs(4999));
    outputs(5680) <= not(layer0_outputs(1993)) or (layer0_outputs(1968));
    outputs(5681) <= not(layer0_outputs(37));
    outputs(5682) <= not(layer0_outputs(327));
    outputs(5683) <= not(layer0_outputs(4120)) or (layer0_outputs(5967));
    outputs(5684) <= not(layer0_outputs(6672)) or (layer0_outputs(8554));
    outputs(5685) <= not(layer0_outputs(6139));
    outputs(5686) <= not(layer0_outputs(6928));
    outputs(5687) <= layer0_outputs(9553);
    outputs(5688) <= (layer0_outputs(3945)) or (layer0_outputs(9762));
    outputs(5689) <= (layer0_outputs(4690)) xor (layer0_outputs(8574));
    outputs(5690) <= not(layer0_outputs(4379));
    outputs(5691) <= not(layer0_outputs(2913));
    outputs(5692) <= not((layer0_outputs(2527)) or (layer0_outputs(8618)));
    outputs(5693) <= not((layer0_outputs(8779)) and (layer0_outputs(3255)));
    outputs(5694) <= (layer0_outputs(1602)) or (layer0_outputs(6652));
    outputs(5695) <= (layer0_outputs(4589)) and not (layer0_outputs(593));
    outputs(5696) <= '1';
    outputs(5697) <= (layer0_outputs(3934)) and not (layer0_outputs(6152));
    outputs(5698) <= not(layer0_outputs(9555));
    outputs(5699) <= layer0_outputs(9189);
    outputs(5700) <= not(layer0_outputs(8012)) or (layer0_outputs(1287));
    outputs(5701) <= (layer0_outputs(875)) xor (layer0_outputs(4461));
    outputs(5702) <= not(layer0_outputs(7499));
    outputs(5703) <= layer0_outputs(6551);
    outputs(5704) <= (layer0_outputs(3260)) xor (layer0_outputs(3458));
    outputs(5705) <= (layer0_outputs(4115)) or (layer0_outputs(9994));
    outputs(5706) <= not((layer0_outputs(5450)) and (layer0_outputs(113)));
    outputs(5707) <= not((layer0_outputs(5462)) xor (layer0_outputs(2276)));
    outputs(5708) <= layer0_outputs(5390);
    outputs(5709) <= layer0_outputs(2618);
    outputs(5710) <= not(layer0_outputs(5905)) or (layer0_outputs(8910));
    outputs(5711) <= layer0_outputs(2389);
    outputs(5712) <= not((layer0_outputs(6236)) xor (layer0_outputs(9103)));
    outputs(5713) <= not(layer0_outputs(3794));
    outputs(5714) <= not((layer0_outputs(7591)) and (layer0_outputs(5814)));
    outputs(5715) <= layer0_outputs(6319);
    outputs(5716) <= not(layer0_outputs(5806));
    outputs(5717) <= not(layer0_outputs(10224));
    outputs(5718) <= layer0_outputs(4316);
    outputs(5719) <= not((layer0_outputs(498)) and (layer0_outputs(9812)));
    outputs(5720) <= (layer0_outputs(1781)) or (layer0_outputs(7224));
    outputs(5721) <= (layer0_outputs(470)) xor (layer0_outputs(40));
    outputs(5722) <= (layer0_outputs(4607)) xor (layer0_outputs(3159));
    outputs(5723) <= not(layer0_outputs(7604));
    outputs(5724) <= not(layer0_outputs(8777)) or (layer0_outputs(733));
    outputs(5725) <= not(layer0_outputs(9106)) or (layer0_outputs(1627));
    outputs(5726) <= (layer0_outputs(7380)) and not (layer0_outputs(8233));
    outputs(5727) <= not(layer0_outputs(5925)) or (layer0_outputs(8905));
    outputs(5728) <= layer0_outputs(3855);
    outputs(5729) <= not((layer0_outputs(9053)) and (layer0_outputs(9626)));
    outputs(5730) <= not(layer0_outputs(490)) or (layer0_outputs(8694));
    outputs(5731) <= not((layer0_outputs(3095)) and (layer0_outputs(1729)));
    outputs(5732) <= (layer0_outputs(1734)) and not (layer0_outputs(2075));
    outputs(5733) <= (layer0_outputs(8166)) xor (layer0_outputs(7665));
    outputs(5734) <= not(layer0_outputs(7742)) or (layer0_outputs(3974));
    outputs(5735) <= not(layer0_outputs(1996)) or (layer0_outputs(9466));
    outputs(5736) <= not(layer0_outputs(2100));
    outputs(5737) <= '0';
    outputs(5738) <= not(layer0_outputs(8451));
    outputs(5739) <= not((layer0_outputs(3471)) and (layer0_outputs(1493)));
    outputs(5740) <= (layer0_outputs(3002)) xor (layer0_outputs(3725));
    outputs(5741) <= (layer0_outputs(2183)) xor (layer0_outputs(6195));
    outputs(5742) <= layer0_outputs(3204);
    outputs(5743) <= layer0_outputs(9618);
    outputs(5744) <= (layer0_outputs(2879)) and not (layer0_outputs(1666));
    outputs(5745) <= (layer0_outputs(9409)) or (layer0_outputs(3688));
    outputs(5746) <= (layer0_outputs(8356)) xor (layer0_outputs(4086));
    outputs(5747) <= (layer0_outputs(800)) or (layer0_outputs(3772));
    outputs(5748) <= (layer0_outputs(144)) xor (layer0_outputs(5581));
    outputs(5749) <= not((layer0_outputs(2338)) and (layer0_outputs(3094)));
    outputs(5750) <= not((layer0_outputs(7940)) xor (layer0_outputs(395)));
    outputs(5751) <= not(layer0_outputs(9105));
    outputs(5752) <= not(layer0_outputs(1567)) or (layer0_outputs(2734));
    outputs(5753) <= (layer0_outputs(9149)) xor (layer0_outputs(9558));
    outputs(5754) <= not(layer0_outputs(2901)) or (layer0_outputs(536));
    outputs(5755) <= not((layer0_outputs(8369)) and (layer0_outputs(3456)));
    outputs(5756) <= (layer0_outputs(8547)) xor (layer0_outputs(4631));
    outputs(5757) <= not(layer0_outputs(2257)) or (layer0_outputs(2997));
    outputs(5758) <= not(layer0_outputs(7018)) or (layer0_outputs(7394));
    outputs(5759) <= (layer0_outputs(4320)) and not (layer0_outputs(6975));
    outputs(5760) <= (layer0_outputs(8862)) and not (layer0_outputs(1374));
    outputs(5761) <= (layer0_outputs(3601)) xor (layer0_outputs(7531));
    outputs(5762) <= (layer0_outputs(1671)) and (layer0_outputs(4107));
    outputs(5763) <= not(layer0_outputs(5782)) or (layer0_outputs(9954));
    outputs(5764) <= (layer0_outputs(9196)) and not (layer0_outputs(6410));
    outputs(5765) <= not(layer0_outputs(4449));
    outputs(5766) <= layer0_outputs(3271);
    outputs(5767) <= (layer0_outputs(8044)) and (layer0_outputs(4485));
    outputs(5768) <= not((layer0_outputs(671)) and (layer0_outputs(7754)));
    outputs(5769) <= not((layer0_outputs(925)) xor (layer0_outputs(226)));
    outputs(5770) <= layer0_outputs(1693);
    outputs(5771) <= layer0_outputs(7830);
    outputs(5772) <= (layer0_outputs(8758)) or (layer0_outputs(2550));
    outputs(5773) <= not((layer0_outputs(4131)) or (layer0_outputs(298)));
    outputs(5774) <= (layer0_outputs(780)) and not (layer0_outputs(5120));
    outputs(5775) <= (layer0_outputs(4065)) and not (layer0_outputs(2885));
    outputs(5776) <= layer0_outputs(2650);
    outputs(5777) <= layer0_outputs(8511);
    outputs(5778) <= not(layer0_outputs(2977));
    outputs(5779) <= (layer0_outputs(2748)) and (layer0_outputs(1042));
    outputs(5780) <= not((layer0_outputs(9541)) and (layer0_outputs(82)));
    outputs(5781) <= not(layer0_outputs(7569));
    outputs(5782) <= (layer0_outputs(6182)) xor (layer0_outputs(2807));
    outputs(5783) <= not((layer0_outputs(7594)) or (layer0_outputs(8247)));
    outputs(5784) <= not(layer0_outputs(5225)) or (layer0_outputs(3104));
    outputs(5785) <= not((layer0_outputs(8629)) xor (layer0_outputs(417)));
    outputs(5786) <= (layer0_outputs(6421)) and not (layer0_outputs(4988));
    outputs(5787) <= not(layer0_outputs(254));
    outputs(5788) <= not(layer0_outputs(2227)) or (layer0_outputs(7080));
    outputs(5789) <= (layer0_outputs(5356)) xor (layer0_outputs(3814));
    outputs(5790) <= (layer0_outputs(7370)) xor (layer0_outputs(7154));
    outputs(5791) <= layer0_outputs(8539);
    outputs(5792) <= not(layer0_outputs(8073));
    outputs(5793) <= layer0_outputs(2406);
    outputs(5794) <= (layer0_outputs(7574)) or (layer0_outputs(6043));
    outputs(5795) <= (layer0_outputs(6477)) and not (layer0_outputs(4346));
    outputs(5796) <= not(layer0_outputs(1022));
    outputs(5797) <= (layer0_outputs(7311)) or (layer0_outputs(4951));
    outputs(5798) <= not(layer0_outputs(6654));
    outputs(5799) <= (layer0_outputs(5932)) xor (layer0_outputs(344));
    outputs(5800) <= not(layer0_outputs(7138)) or (layer0_outputs(3472));
    outputs(5801) <= not(layer0_outputs(9448)) or (layer0_outputs(8987));
    outputs(5802) <= not(layer0_outputs(2891)) or (layer0_outputs(2466));
    outputs(5803) <= (layer0_outputs(9919)) and not (layer0_outputs(5276));
    outputs(5804) <= (layer0_outputs(5088)) xor (layer0_outputs(3594));
    outputs(5805) <= (layer0_outputs(9290)) and (layer0_outputs(916));
    outputs(5806) <= layer0_outputs(5658);
    outputs(5807) <= not((layer0_outputs(5766)) xor (layer0_outputs(2849)));
    outputs(5808) <= not((layer0_outputs(7453)) xor (layer0_outputs(4016)));
    outputs(5809) <= layer0_outputs(4491);
    outputs(5810) <= layer0_outputs(3658);
    outputs(5811) <= not((layer0_outputs(5329)) and (layer0_outputs(9200)));
    outputs(5812) <= layer0_outputs(6583);
    outputs(5813) <= not((layer0_outputs(6489)) xor (layer0_outputs(6460)));
    outputs(5814) <= not(layer0_outputs(5833));
    outputs(5815) <= layer0_outputs(3926);
    outputs(5816) <= (layer0_outputs(1070)) and not (layer0_outputs(2143));
    outputs(5817) <= not(layer0_outputs(8578));
    outputs(5818) <= (layer0_outputs(1288)) and (layer0_outputs(1672));
    outputs(5819) <= (layer0_outputs(8800)) xor (layer0_outputs(8736));
    outputs(5820) <= not(layer0_outputs(7085));
    outputs(5821) <= not(layer0_outputs(7790));
    outputs(5822) <= not((layer0_outputs(8849)) or (layer0_outputs(6402)));
    outputs(5823) <= not((layer0_outputs(3615)) xor (layer0_outputs(6728)));
    outputs(5824) <= not(layer0_outputs(7121));
    outputs(5825) <= (layer0_outputs(7819)) and (layer0_outputs(91));
    outputs(5826) <= not(layer0_outputs(1148)) or (layer0_outputs(6526));
    outputs(5827) <= not((layer0_outputs(5590)) xor (layer0_outputs(4158)));
    outputs(5828) <= (layer0_outputs(9335)) xor (layer0_outputs(5889));
    outputs(5829) <= layer0_outputs(1024);
    outputs(5830) <= (layer0_outputs(6118)) and not (layer0_outputs(6799));
    outputs(5831) <= (layer0_outputs(3858)) and not (layer0_outputs(7106));
    outputs(5832) <= not((layer0_outputs(5362)) xor (layer0_outputs(8998)));
    outputs(5833) <= (layer0_outputs(1331)) xor (layer0_outputs(2965));
    outputs(5834) <= not(layer0_outputs(2381)) or (layer0_outputs(1581));
    outputs(5835) <= (layer0_outputs(9731)) and not (layer0_outputs(7115));
    outputs(5836) <= (layer0_outputs(2565)) xor (layer0_outputs(819));
    outputs(5837) <= not(layer0_outputs(205)) or (layer0_outputs(3620));
    outputs(5838) <= '1';
    outputs(5839) <= not((layer0_outputs(1048)) and (layer0_outputs(1409)));
    outputs(5840) <= (layer0_outputs(7786)) and (layer0_outputs(1717));
    outputs(5841) <= not(layer0_outputs(4048));
    outputs(5842) <= layer0_outputs(6259);
    outputs(5843) <= not(layer0_outputs(8982));
    outputs(5844) <= (layer0_outputs(1772)) and not (layer0_outputs(2273));
    outputs(5845) <= not(layer0_outputs(9756)) or (layer0_outputs(8813));
    outputs(5846) <= not((layer0_outputs(3114)) or (layer0_outputs(448)));
    outputs(5847) <= layer0_outputs(8372);
    outputs(5848) <= layer0_outputs(2133);
    outputs(5849) <= (layer0_outputs(6359)) xor (layer0_outputs(5914));
    outputs(5850) <= not(layer0_outputs(7711));
    outputs(5851) <= layer0_outputs(3743);
    outputs(5852) <= not(layer0_outputs(6329)) or (layer0_outputs(9252));
    outputs(5853) <= not((layer0_outputs(3050)) xor (layer0_outputs(8316)));
    outputs(5854) <= layer0_outputs(884);
    outputs(5855) <= not((layer0_outputs(420)) xor (layer0_outputs(6261)));
    outputs(5856) <= (layer0_outputs(7396)) and not (layer0_outputs(4718));
    outputs(5857) <= (layer0_outputs(8737)) xor (layer0_outputs(1993));
    outputs(5858) <= layer0_outputs(1533);
    outputs(5859) <= not(layer0_outputs(1874));
    outputs(5860) <= not(layer0_outputs(2007));
    outputs(5861) <= not((layer0_outputs(8897)) and (layer0_outputs(1773)));
    outputs(5862) <= (layer0_outputs(8332)) xor (layer0_outputs(9770));
    outputs(5863) <= not(layer0_outputs(9181));
    outputs(5864) <= not(layer0_outputs(5743)) or (layer0_outputs(7694));
    outputs(5865) <= not((layer0_outputs(3060)) and (layer0_outputs(5245)));
    outputs(5866) <= not((layer0_outputs(3303)) and (layer0_outputs(7791)));
    outputs(5867) <= not(layer0_outputs(4279)) or (layer0_outputs(5447));
    outputs(5868) <= not(layer0_outputs(1783));
    outputs(5869) <= not(layer0_outputs(331));
    outputs(5870) <= (layer0_outputs(5744)) and not (layer0_outputs(4532));
    outputs(5871) <= layer0_outputs(4567);
    outputs(5872) <= layer0_outputs(8816);
    outputs(5873) <= not(layer0_outputs(4345));
    outputs(5874) <= layer0_outputs(8212);
    outputs(5875) <= layer0_outputs(9322);
    outputs(5876) <= (layer0_outputs(2417)) xor (layer0_outputs(6942));
    outputs(5877) <= not(layer0_outputs(2845)) or (layer0_outputs(44));
    outputs(5878) <= not(layer0_outputs(2160));
    outputs(5879) <= not(layer0_outputs(2588));
    outputs(5880) <= (layer0_outputs(4425)) and (layer0_outputs(1488));
    outputs(5881) <= layer0_outputs(6347);
    outputs(5882) <= (layer0_outputs(2313)) or (layer0_outputs(5628));
    outputs(5883) <= layer0_outputs(4283);
    outputs(5884) <= (layer0_outputs(1724)) and not (layer0_outputs(1596));
    outputs(5885) <= (layer0_outputs(10026)) xor (layer0_outputs(4454));
    outputs(5886) <= (layer0_outputs(9278)) and not (layer0_outputs(8918));
    outputs(5887) <= (layer0_outputs(1328)) xor (layer0_outputs(9820));
    outputs(5888) <= not((layer0_outputs(4264)) xor (layer0_outputs(5816)));
    outputs(5889) <= not(layer0_outputs(3611)) or (layer0_outputs(7998));
    outputs(5890) <= layer0_outputs(307);
    outputs(5891) <= not(layer0_outputs(7064));
    outputs(5892) <= not(layer0_outputs(5209));
    outputs(5893) <= layer0_outputs(6945);
    outputs(5894) <= not(layer0_outputs(2539));
    outputs(5895) <= not((layer0_outputs(3115)) xor (layer0_outputs(3637)));
    outputs(5896) <= layer0_outputs(7173);
    outputs(5897) <= not(layer0_outputs(4310));
    outputs(5898) <= layer0_outputs(4650);
    outputs(5899) <= not(layer0_outputs(3437)) or (layer0_outputs(9959));
    outputs(5900) <= (layer0_outputs(2237)) or (layer0_outputs(8374));
    outputs(5901) <= (layer0_outputs(6994)) and not (layer0_outputs(242));
    outputs(5902) <= layer0_outputs(8029);
    outputs(5903) <= not(layer0_outputs(5522));
    outputs(5904) <= not(layer0_outputs(3538)) or (layer0_outputs(8719));
    outputs(5905) <= layer0_outputs(6617);
    outputs(5906) <= layer0_outputs(3187);
    outputs(5907) <= (layer0_outputs(923)) and not (layer0_outputs(681));
    outputs(5908) <= not(layer0_outputs(9095));
    outputs(5909) <= not(layer0_outputs(276));
    outputs(5910) <= layer0_outputs(8526);
    outputs(5911) <= not(layer0_outputs(8034)) or (layer0_outputs(6914));
    outputs(5912) <= (layer0_outputs(8873)) and (layer0_outputs(4067));
    outputs(5913) <= not(layer0_outputs(4221));
    outputs(5914) <= not(layer0_outputs(6527)) or (layer0_outputs(9336));
    outputs(5915) <= layer0_outputs(4338);
    outputs(5916) <= not(layer0_outputs(6834));
    outputs(5917) <= not(layer0_outputs(6994)) or (layer0_outputs(2893));
    outputs(5918) <= not(layer0_outputs(8671));
    outputs(5919) <= not(layer0_outputs(6859));
    outputs(5920) <= layer0_outputs(7183);
    outputs(5921) <= (layer0_outputs(5626)) and not (layer0_outputs(407));
    outputs(5922) <= not(layer0_outputs(6291));
    outputs(5923) <= layer0_outputs(6314);
    outputs(5924) <= not(layer0_outputs(9082)) or (layer0_outputs(3092));
    outputs(5925) <= layer0_outputs(5879);
    outputs(5926) <= not(layer0_outputs(7496));
    outputs(5927) <= not((layer0_outputs(8998)) or (layer0_outputs(3730)));
    outputs(5928) <= (layer0_outputs(6633)) and not (layer0_outputs(6349));
    outputs(5929) <= (layer0_outputs(8812)) or (layer0_outputs(9205));
    outputs(5930) <= not(layer0_outputs(1003));
    outputs(5931) <= not(layer0_outputs(7562));
    outputs(5932) <= not(layer0_outputs(8804)) or (layer0_outputs(9558));
    outputs(5933) <= not(layer0_outputs(8544)) or (layer0_outputs(9098));
    outputs(5934) <= (layer0_outputs(3182)) or (layer0_outputs(9567));
    outputs(5935) <= (layer0_outputs(7595)) and not (layer0_outputs(8677));
    outputs(5936) <= (layer0_outputs(5619)) xor (layer0_outputs(908));
    outputs(5937) <= not(layer0_outputs(9503));
    outputs(5938) <= not(layer0_outputs(280));
    outputs(5939) <= (layer0_outputs(2605)) and not (layer0_outputs(2458));
    outputs(5940) <= layer0_outputs(704);
    outputs(5941) <= layer0_outputs(4793);
    outputs(5942) <= not(layer0_outputs(7892));
    outputs(5943) <= not((layer0_outputs(9142)) xor (layer0_outputs(3153)));
    outputs(5944) <= (layer0_outputs(1221)) and (layer0_outputs(1251));
    outputs(5945) <= not((layer0_outputs(3530)) xor (layer0_outputs(4856)));
    outputs(5946) <= not((layer0_outputs(9765)) xor (layer0_outputs(1112)));
    outputs(5947) <= not((layer0_outputs(4603)) and (layer0_outputs(3539)));
    outputs(5948) <= layer0_outputs(7539);
    outputs(5949) <= layer0_outputs(299);
    outputs(5950) <= layer0_outputs(3606);
    outputs(5951) <= (layer0_outputs(9583)) or (layer0_outputs(4509));
    outputs(5952) <= (layer0_outputs(1494)) or (layer0_outputs(2499));
    outputs(5953) <= layer0_outputs(1534);
    outputs(5954) <= not((layer0_outputs(2587)) and (layer0_outputs(8785)));
    outputs(5955) <= (layer0_outputs(2884)) and (layer0_outputs(9566));
    outputs(5956) <= not((layer0_outputs(8668)) xor (layer0_outputs(3417)));
    outputs(5957) <= (layer0_outputs(4722)) or (layer0_outputs(7107));
    outputs(5958) <= (layer0_outputs(1962)) xor (layer0_outputs(9396));
    outputs(5959) <= not((layer0_outputs(3864)) and (layer0_outputs(1989)));
    outputs(5960) <= (layer0_outputs(2543)) or (layer0_outputs(5033));
    outputs(5961) <= not((layer0_outputs(7181)) or (layer0_outputs(3753)));
    outputs(5962) <= not((layer0_outputs(4953)) xor (layer0_outputs(8988)));
    outputs(5963) <= (layer0_outputs(939)) or (layer0_outputs(6324));
    outputs(5964) <= not(layer0_outputs(3403));
    outputs(5965) <= layer0_outputs(7926);
    outputs(5966) <= not((layer0_outputs(8893)) and (layer0_outputs(9874)));
    outputs(5967) <= not((layer0_outputs(4080)) and (layer0_outputs(941)));
    outputs(5968) <= (layer0_outputs(4713)) xor (layer0_outputs(9934));
    outputs(5969) <= not(layer0_outputs(659));
    outputs(5970) <= not((layer0_outputs(3797)) xor (layer0_outputs(5917)));
    outputs(5971) <= (layer0_outputs(7862)) xor (layer0_outputs(3317));
    outputs(5972) <= not(layer0_outputs(8558));
    outputs(5973) <= layer0_outputs(6232);
    outputs(5974) <= not(layer0_outputs(6919));
    outputs(5975) <= not(layer0_outputs(2384));
    outputs(5976) <= (layer0_outputs(6550)) and (layer0_outputs(4977));
    outputs(5977) <= (layer0_outputs(5022)) xor (layer0_outputs(3991));
    outputs(5978) <= layer0_outputs(5517);
    outputs(5979) <= (layer0_outputs(9087)) xor (layer0_outputs(7161));
    outputs(5980) <= not(layer0_outputs(6603));
    outputs(5981) <= layer0_outputs(7170);
    outputs(5982) <= not(layer0_outputs(5947));
    outputs(5983) <= not(layer0_outputs(610));
    outputs(5984) <= not((layer0_outputs(5215)) and (layer0_outputs(9669)));
    outputs(5985) <= not(layer0_outputs(2310)) or (layer0_outputs(2514));
    outputs(5986) <= not(layer0_outputs(3711)) or (layer0_outputs(614));
    outputs(5987) <= not((layer0_outputs(6164)) or (layer0_outputs(6808)));
    outputs(5988) <= layer0_outputs(2018);
    outputs(5989) <= (layer0_outputs(9472)) and not (layer0_outputs(6414));
    outputs(5990) <= not((layer0_outputs(596)) xor (layer0_outputs(2939)));
    outputs(5991) <= not(layer0_outputs(4332));
    outputs(5992) <= (layer0_outputs(910)) and not (layer0_outputs(6509));
    outputs(5993) <= not(layer0_outputs(2763)) or (layer0_outputs(1351));
    outputs(5994) <= layer0_outputs(519);
    outputs(5995) <= not((layer0_outputs(6148)) or (layer0_outputs(8791)));
    outputs(5996) <= not(layer0_outputs(1229)) or (layer0_outputs(9656));
    outputs(5997) <= not((layer0_outputs(3336)) or (layer0_outputs(9836)));
    outputs(5998) <= (layer0_outputs(3186)) xor (layer0_outputs(9413));
    outputs(5999) <= not((layer0_outputs(3418)) xor (layer0_outputs(357)));
    outputs(6000) <= not((layer0_outputs(2401)) xor (layer0_outputs(5579)));
    outputs(6001) <= (layer0_outputs(337)) xor (layer0_outputs(5814));
    outputs(6002) <= not(layer0_outputs(9611));
    outputs(6003) <= not(layer0_outputs(2957)) or (layer0_outputs(300));
    outputs(6004) <= not(layer0_outputs(6872));
    outputs(6005) <= not(layer0_outputs(137));
    outputs(6006) <= (layer0_outputs(3455)) or (layer0_outputs(1805));
    outputs(6007) <= not(layer0_outputs(6051));
    outputs(6008) <= not(layer0_outputs(8045));
    outputs(6009) <= not((layer0_outputs(6301)) xor (layer0_outputs(3544)));
    outputs(6010) <= not((layer0_outputs(956)) and (layer0_outputs(1138)));
    outputs(6011) <= not((layer0_outputs(172)) and (layer0_outputs(1055)));
    outputs(6012) <= not((layer0_outputs(5443)) xor (layer0_outputs(5494)));
    outputs(6013) <= not(layer0_outputs(2850));
    outputs(6014) <= (layer0_outputs(2371)) xor (layer0_outputs(7643));
    outputs(6015) <= layer0_outputs(1422);
    outputs(6016) <= not((layer0_outputs(4820)) xor (layer0_outputs(1550)));
    outputs(6017) <= not(layer0_outputs(5505)) or (layer0_outputs(1221));
    outputs(6018) <= layer0_outputs(501);
    outputs(6019) <= (layer0_outputs(1787)) and not (layer0_outputs(6186));
    outputs(6020) <= not(layer0_outputs(9730)) or (layer0_outputs(6715));
    outputs(6021) <= (layer0_outputs(1175)) xor (layer0_outputs(2546));
    outputs(6022) <= not(layer0_outputs(2914));
    outputs(6023) <= '1';
    outputs(6024) <= not(layer0_outputs(6813)) or (layer0_outputs(1098));
    outputs(6025) <= layer0_outputs(9538);
    outputs(6026) <= (layer0_outputs(7154)) xor (layer0_outputs(4042));
    outputs(6027) <= not((layer0_outputs(5846)) and (layer0_outputs(9781)));
    outputs(6028) <= not(layer0_outputs(7492));
    outputs(6029) <= layer0_outputs(7164);
    outputs(6030) <= (layer0_outputs(92)) xor (layer0_outputs(1260));
    outputs(6031) <= not(layer0_outputs(2263));
    outputs(6032) <= layer0_outputs(6938);
    outputs(6033) <= not((layer0_outputs(9265)) xor (layer0_outputs(9067)));
    outputs(6034) <= not((layer0_outputs(6954)) xor (layer0_outputs(7658)));
    outputs(6035) <= not(layer0_outputs(4395));
    outputs(6036) <= not((layer0_outputs(1595)) xor (layer0_outputs(2325)));
    outputs(6037) <= (layer0_outputs(7462)) xor (layer0_outputs(6010));
    outputs(6038) <= (layer0_outputs(4002)) and (layer0_outputs(3890));
    outputs(6039) <= (layer0_outputs(9648)) and not (layer0_outputs(4275));
    outputs(6040) <= (layer0_outputs(4711)) xor (layer0_outputs(5406));
    outputs(6041) <= layer0_outputs(584);
    outputs(6042) <= not((layer0_outputs(7826)) xor (layer0_outputs(3684)));
    outputs(6043) <= not((layer0_outputs(8042)) and (layer0_outputs(3218)));
    outputs(6044) <= not((layer0_outputs(8046)) xor (layer0_outputs(673)));
    outputs(6045) <= (layer0_outputs(5668)) and not (layer0_outputs(618));
    outputs(6046) <= not(layer0_outputs(6969)) or (layer0_outputs(2606));
    outputs(6047) <= (layer0_outputs(9408)) xor (layer0_outputs(6755));
    outputs(6048) <= (layer0_outputs(1587)) and not (layer0_outputs(2080));
    outputs(6049) <= (layer0_outputs(8461)) and (layer0_outputs(1114));
    outputs(6050) <= not(layer0_outputs(1152)) or (layer0_outputs(2150));
    outputs(6051) <= not(layer0_outputs(2923)) or (layer0_outputs(8204));
    outputs(6052) <= (layer0_outputs(7908)) or (layer0_outputs(3849));
    outputs(6053) <= layer0_outputs(4654);
    outputs(6054) <= (layer0_outputs(8295)) and not (layer0_outputs(1823));
    outputs(6055) <= not((layer0_outputs(1239)) xor (layer0_outputs(412)));
    outputs(6056) <= layer0_outputs(3393);
    outputs(6057) <= layer0_outputs(2244);
    outputs(6058) <= '0';
    outputs(6059) <= not(layer0_outputs(5720));
    outputs(6060) <= (layer0_outputs(2301)) xor (layer0_outputs(5046));
    outputs(6061) <= (layer0_outputs(3529)) and not (layer0_outputs(5727));
    outputs(6062) <= (layer0_outputs(2277)) and not (layer0_outputs(6544));
    outputs(6063) <= (layer0_outputs(2139)) xor (layer0_outputs(6261));
    outputs(6064) <= layer0_outputs(5870);
    outputs(6065) <= not(layer0_outputs(1311));
    outputs(6066) <= not(layer0_outputs(7976)) or (layer0_outputs(2499));
    outputs(6067) <= layer0_outputs(2650);
    outputs(6068) <= not((layer0_outputs(3770)) xor (layer0_outputs(2016)));
    outputs(6069) <= not(layer0_outputs(1838)) or (layer0_outputs(7133));
    outputs(6070) <= not((layer0_outputs(5400)) xor (layer0_outputs(9386)));
    outputs(6071) <= layer0_outputs(2878);
    outputs(6072) <= not((layer0_outputs(8322)) xor (layer0_outputs(9592)));
    outputs(6073) <= not((layer0_outputs(5679)) xor (layer0_outputs(9436)));
    outputs(6074) <= not((layer0_outputs(1662)) and (layer0_outputs(9080)));
    outputs(6075) <= (layer0_outputs(2908)) xor (layer0_outputs(7739));
    outputs(6076) <= (layer0_outputs(6587)) and (layer0_outputs(3071));
    outputs(6077) <= not((layer0_outputs(3340)) xor (layer0_outputs(3677)));
    outputs(6078) <= not(layer0_outputs(4201));
    outputs(6079) <= not((layer0_outputs(6843)) xor (layer0_outputs(7814)));
    outputs(6080) <= (layer0_outputs(2678)) and (layer0_outputs(3883));
    outputs(6081) <= (layer0_outputs(6399)) xor (layer0_outputs(5412));
    outputs(6082) <= not(layer0_outputs(1718));
    outputs(6083) <= layer0_outputs(5768);
    outputs(6084) <= (layer0_outputs(8410)) or (layer0_outputs(560));
    outputs(6085) <= (layer0_outputs(5087)) and not (layer0_outputs(8102));
    outputs(6086) <= not(layer0_outputs(1058)) or (layer0_outputs(9101));
    outputs(6087) <= not(layer0_outputs(2105));
    outputs(6088) <= not((layer0_outputs(1209)) or (layer0_outputs(5919)));
    outputs(6089) <= layer0_outputs(2760);
    outputs(6090) <= not(layer0_outputs(585)) or (layer0_outputs(2554));
    outputs(6091) <= (layer0_outputs(5151)) and (layer0_outputs(4333));
    outputs(6092) <= not(layer0_outputs(1231)) or (layer0_outputs(6158));
    outputs(6093) <= not(layer0_outputs(845)) or (layer0_outputs(8839));
    outputs(6094) <= not((layer0_outputs(8291)) xor (layer0_outputs(6511)));
    outputs(6095) <= (layer0_outputs(1265)) xor (layer0_outputs(7935));
    outputs(6096) <= not(layer0_outputs(4736));
    outputs(6097) <= (layer0_outputs(2662)) or (layer0_outputs(8101));
    outputs(6098) <= layer0_outputs(5670);
    outputs(6099) <= (layer0_outputs(7991)) and not (layer0_outputs(2347));
    outputs(6100) <= (layer0_outputs(7057)) or (layer0_outputs(6813));
    outputs(6101) <= (layer0_outputs(3731)) and (layer0_outputs(7323));
    outputs(6102) <= (layer0_outputs(5288)) xor (layer0_outputs(2433));
    outputs(6103) <= not(layer0_outputs(9595)) or (layer0_outputs(4261));
    outputs(6104) <= not(layer0_outputs(8436));
    outputs(6105) <= not(layer0_outputs(1967));
    outputs(6106) <= layer0_outputs(4652);
    outputs(6107) <= (layer0_outputs(819)) xor (layer0_outputs(2551));
    outputs(6108) <= (layer0_outputs(6231)) and (layer0_outputs(1755));
    outputs(6109) <= not(layer0_outputs(3482)) or (layer0_outputs(404));
    outputs(6110) <= (layer0_outputs(5969)) and not (layer0_outputs(850));
    outputs(6111) <= layer0_outputs(6912);
    outputs(6112) <= layer0_outputs(562);
    outputs(6113) <= not(layer0_outputs(9829)) or (layer0_outputs(2298));
    outputs(6114) <= not((layer0_outputs(1599)) xor (layer0_outputs(7882)));
    outputs(6115) <= not((layer0_outputs(2057)) xor (layer0_outputs(3062)));
    outputs(6116) <= layer0_outputs(277);
    outputs(6117) <= layer0_outputs(6240);
    outputs(6118) <= not(layer0_outputs(4091));
    outputs(6119) <= layer0_outputs(1241);
    outputs(6120) <= layer0_outputs(6103);
    outputs(6121) <= not(layer0_outputs(9728));
    outputs(6122) <= not((layer0_outputs(6741)) xor (layer0_outputs(3477)));
    outputs(6123) <= (layer0_outputs(2019)) and not (layer0_outputs(1435));
    outputs(6124) <= not(layer0_outputs(7330));
    outputs(6125) <= not((layer0_outputs(155)) xor (layer0_outputs(661)));
    outputs(6126) <= not((layer0_outputs(3740)) or (layer0_outputs(394)));
    outputs(6127) <= (layer0_outputs(1684)) xor (layer0_outputs(835));
    outputs(6128) <= not((layer0_outputs(4780)) or (layer0_outputs(5111)));
    outputs(6129) <= layer0_outputs(2653);
    outputs(6130) <= (layer0_outputs(48)) and not (layer0_outputs(10));
    outputs(6131) <= not(layer0_outputs(8634));
    outputs(6132) <= not((layer0_outputs(2725)) xor (layer0_outputs(9000)));
    outputs(6133) <= (layer0_outputs(567)) or (layer0_outputs(7726));
    outputs(6134) <= not((layer0_outputs(1378)) xor (layer0_outputs(2776)));
    outputs(6135) <= not(layer0_outputs(9308)) or (layer0_outputs(8983));
    outputs(6136) <= not((layer0_outputs(5725)) xor (layer0_outputs(9045)));
    outputs(6137) <= layer0_outputs(904);
    outputs(6138) <= not(layer0_outputs(9516));
    outputs(6139) <= layer0_outputs(3676);
    outputs(6140) <= (layer0_outputs(5516)) and not (layer0_outputs(1448));
    outputs(6141) <= (layer0_outputs(1954)) and not (layer0_outputs(3111));
    outputs(6142) <= (layer0_outputs(10212)) or (layer0_outputs(5580));
    outputs(6143) <= layer0_outputs(2180);
    outputs(6144) <= layer0_outputs(7163);
    outputs(6145) <= not(layer0_outputs(2087));
    outputs(6146) <= (layer0_outputs(6186)) xor (layer0_outputs(6715));
    outputs(6147) <= not((layer0_outputs(4606)) xor (layer0_outputs(4737)));
    outputs(6148) <= layer0_outputs(8795);
    outputs(6149) <= not(layer0_outputs(8642));
    outputs(6150) <= not(layer0_outputs(4251));
    outputs(6151) <= layer0_outputs(3322);
    outputs(6152) <= not((layer0_outputs(10176)) and (layer0_outputs(4871)));
    outputs(6153) <= not(layer0_outputs(3472));
    outputs(6154) <= not(layer0_outputs(1631));
    outputs(6155) <= layer0_outputs(288);
    outputs(6156) <= not(layer0_outputs(139));
    outputs(6157) <= '0';
    outputs(6158) <= (layer0_outputs(4416)) and not (layer0_outputs(2169));
    outputs(6159) <= layer0_outputs(9270);
    outputs(6160) <= (layer0_outputs(4636)) and (layer0_outputs(1811));
    outputs(6161) <= layer0_outputs(3223);
    outputs(6162) <= not(layer0_outputs(9512));
    outputs(6163) <= (layer0_outputs(3770)) xor (layer0_outputs(6122));
    outputs(6164) <= (layer0_outputs(6731)) xor (layer0_outputs(1071));
    outputs(6165) <= not((layer0_outputs(128)) and (layer0_outputs(8815)));
    outputs(6166) <= (layer0_outputs(3147)) xor (layer0_outputs(1853));
    outputs(6167) <= (layer0_outputs(4997)) and not (layer0_outputs(5083));
    outputs(6168) <= not(layer0_outputs(6417));
    outputs(6169) <= not((layer0_outputs(4143)) or (layer0_outputs(1002)));
    outputs(6170) <= (layer0_outputs(8168)) xor (layer0_outputs(7145));
    outputs(6171) <= not(layer0_outputs(7755)) or (layer0_outputs(4111));
    outputs(6172) <= (layer0_outputs(9930)) or (layer0_outputs(2766));
    outputs(6173) <= not((layer0_outputs(3298)) xor (layer0_outputs(9064)));
    outputs(6174) <= layer0_outputs(8499);
    outputs(6175) <= not((layer0_outputs(9212)) xor (layer0_outputs(1471)));
    outputs(6176) <= not(layer0_outputs(2166)) or (layer0_outputs(7208));
    outputs(6177) <= not(layer0_outputs(2714));
    outputs(6178) <= not((layer0_outputs(8455)) xor (layer0_outputs(8382)));
    outputs(6179) <= layer0_outputs(2306);
    outputs(6180) <= not((layer0_outputs(7596)) and (layer0_outputs(3778)));
    outputs(6181) <= (layer0_outputs(2147)) xor (layer0_outputs(8433));
    outputs(6182) <= layer0_outputs(4724);
    outputs(6183) <= not(layer0_outputs(5332)) or (layer0_outputs(9585));
    outputs(6184) <= (layer0_outputs(7199)) xor (layer0_outputs(9499));
    outputs(6185) <= (layer0_outputs(5978)) xor (layer0_outputs(9717));
    outputs(6186) <= layer0_outputs(10124);
    outputs(6187) <= (layer0_outputs(6284)) and not (layer0_outputs(558));
    outputs(6188) <= not(layer0_outputs(946));
    outputs(6189) <= (layer0_outputs(5922)) and (layer0_outputs(582));
    outputs(6190) <= layer0_outputs(608);
    outputs(6191) <= not(layer0_outputs(3627));
    outputs(6192) <= not(layer0_outputs(4571));
    outputs(6193) <= layer0_outputs(152);
    outputs(6194) <= (layer0_outputs(6123)) xor (layer0_outputs(5826));
    outputs(6195) <= not((layer0_outputs(1594)) xor (layer0_outputs(9624)));
    outputs(6196) <= not(layer0_outputs(5063));
    outputs(6197) <= layer0_outputs(3209);
    outputs(6198) <= not(layer0_outputs(6458));
    outputs(6199) <= not(layer0_outputs(4458));
    outputs(6200) <= not(layer0_outputs(15));
    outputs(6201) <= layer0_outputs(963);
    outputs(6202) <= (layer0_outputs(5736)) xor (layer0_outputs(6558));
    outputs(6203) <= layer0_outputs(4250);
    outputs(6204) <= layer0_outputs(1690);
    outputs(6205) <= layer0_outputs(7291);
    outputs(6206) <= (layer0_outputs(4384)) xor (layer0_outputs(1652));
    outputs(6207) <= not(layer0_outputs(2205));
    outputs(6208) <= not(layer0_outputs(8780));
    outputs(6209) <= not(layer0_outputs(9862));
    outputs(6210) <= layer0_outputs(3666);
    outputs(6211) <= (layer0_outputs(2067)) xor (layer0_outputs(8802));
    outputs(6212) <= not(layer0_outputs(3812));
    outputs(6213) <= not(layer0_outputs(3768));
    outputs(6214) <= (layer0_outputs(6241)) xor (layer0_outputs(3746));
    outputs(6215) <= layer0_outputs(896);
    outputs(6216) <= not(layer0_outputs(9463));
    outputs(6217) <= not(layer0_outputs(6930));
    outputs(6218) <= (layer0_outputs(1725)) or (layer0_outputs(9280));
    outputs(6219) <= (layer0_outputs(7449)) or (layer0_outputs(5778));
    outputs(6220) <= layer0_outputs(2538);
    outputs(6221) <= (layer0_outputs(8189)) and not (layer0_outputs(4140));
    outputs(6222) <= not(layer0_outputs(1798));
    outputs(6223) <= (layer0_outputs(7233)) and not (layer0_outputs(3035));
    outputs(6224) <= layer0_outputs(2599);
    outputs(6225) <= not((layer0_outputs(3007)) xor (layer0_outputs(4068)));
    outputs(6226) <= (layer0_outputs(8282)) and not (layer0_outputs(6017));
    outputs(6227) <= not((layer0_outputs(2222)) or (layer0_outputs(1557)));
    outputs(6228) <= not((layer0_outputs(3750)) xor (layer0_outputs(2610)));
    outputs(6229) <= (layer0_outputs(3080)) xor (layer0_outputs(6528));
    outputs(6230) <= not((layer0_outputs(3414)) and (layer0_outputs(6131)));
    outputs(6231) <= not(layer0_outputs(6458));
    outputs(6232) <= layer0_outputs(3927);
    outputs(6233) <= layer0_outputs(3925);
    outputs(6234) <= not(layer0_outputs(1598));
    outputs(6235) <= not((layer0_outputs(2836)) and (layer0_outputs(5815)));
    outputs(6236) <= not(layer0_outputs(3743));
    outputs(6237) <= not((layer0_outputs(9902)) xor (layer0_outputs(3228)));
    outputs(6238) <= (layer0_outputs(7125)) and (layer0_outputs(88));
    outputs(6239) <= (layer0_outputs(4669)) and not (layer0_outputs(344));
    outputs(6240) <= (layer0_outputs(606)) and (layer0_outputs(7779));
    outputs(6241) <= not(layer0_outputs(4096));
    outputs(6242) <= layer0_outputs(7923);
    outputs(6243) <= not(layer0_outputs(772));
    outputs(6244) <= layer0_outputs(1755);
    outputs(6245) <= not(layer0_outputs(6444));
    outputs(6246) <= (layer0_outputs(9954)) xor (layer0_outputs(2691));
    outputs(6247) <= layer0_outputs(6435);
    outputs(6248) <= not((layer0_outputs(1718)) or (layer0_outputs(6158)));
    outputs(6249) <= layer0_outputs(8628);
    outputs(6250) <= not((layer0_outputs(2529)) xor (layer0_outputs(2098)));
    outputs(6251) <= not(layer0_outputs(2043));
    outputs(6252) <= (layer0_outputs(5119)) and not (layer0_outputs(6260));
    outputs(6253) <= not((layer0_outputs(385)) or (layer0_outputs(5421)));
    outputs(6254) <= layer0_outputs(9256);
    outputs(6255) <= not((layer0_outputs(8340)) or (layer0_outputs(2021)));
    outputs(6256) <= not((layer0_outputs(7972)) or (layer0_outputs(9811)));
    outputs(6257) <= layer0_outputs(815);
    outputs(6258) <= layer0_outputs(5273);
    outputs(6259) <= '0';
    outputs(6260) <= (layer0_outputs(3230)) and not (layer0_outputs(3310));
    outputs(6261) <= layer0_outputs(9481);
    outputs(6262) <= (layer0_outputs(9299)) or (layer0_outputs(3263));
    outputs(6263) <= (layer0_outputs(7869)) xor (layer0_outputs(5896));
    outputs(6264) <= (layer0_outputs(7521)) xor (layer0_outputs(1621));
    outputs(6265) <= not(layer0_outputs(978));
    outputs(6266) <= (layer0_outputs(5573)) xor (layer0_outputs(8401));
    outputs(6267) <= not((layer0_outputs(8420)) xor (layer0_outputs(8072)));
    outputs(6268) <= not(layer0_outputs(8919));
    outputs(6269) <= not((layer0_outputs(8791)) or (layer0_outputs(6513)));
    outputs(6270) <= not((layer0_outputs(620)) xor (layer0_outputs(4183)));
    outputs(6271) <= not(layer0_outputs(4347)) or (layer0_outputs(5075));
    outputs(6272) <= (layer0_outputs(2286)) and (layer0_outputs(2628));
    outputs(6273) <= not(layer0_outputs(2827));
    outputs(6274) <= not(layer0_outputs(9741));
    outputs(6275) <= not(layer0_outputs(8925));
    outputs(6276) <= not(layer0_outputs(6850));
    outputs(6277) <= (layer0_outputs(7622)) xor (layer0_outputs(1600));
    outputs(6278) <= layer0_outputs(9476);
    outputs(6279) <= not(layer0_outputs(5625)) or (layer0_outputs(361));
    outputs(6280) <= not(layer0_outputs(9238)) or (layer0_outputs(4498));
    outputs(6281) <= not(layer0_outputs(2735)) or (layer0_outputs(9337));
    outputs(6282) <= not((layer0_outputs(4990)) xor (layer0_outputs(4710)));
    outputs(6283) <= not(layer0_outputs(3002));
    outputs(6284) <= (layer0_outputs(4401)) and not (layer0_outputs(3757));
    outputs(6285) <= not(layer0_outputs(10028));
    outputs(6286) <= not(layer0_outputs(2374)) or (layer0_outputs(8287));
    outputs(6287) <= (layer0_outputs(476)) xor (layer0_outputs(2525));
    outputs(6288) <= not(layer0_outputs(8907));
    outputs(6289) <= not((layer0_outputs(2435)) or (layer0_outputs(6210)));
    outputs(6290) <= (layer0_outputs(4744)) xor (layer0_outputs(4104));
    outputs(6291) <= layer0_outputs(6936);
    outputs(6292) <= not(layer0_outputs(6363));
    outputs(6293) <= (layer0_outputs(8501)) and not (layer0_outputs(7398));
    outputs(6294) <= not((layer0_outputs(2298)) xor (layer0_outputs(7870)));
    outputs(6295) <= layer0_outputs(3822);
    outputs(6296) <= not((layer0_outputs(5141)) or (layer0_outputs(6639)));
    outputs(6297) <= not(layer0_outputs(7316));
    outputs(6298) <= layer0_outputs(2707);
    outputs(6299) <= (layer0_outputs(1243)) or (layer0_outputs(579));
    outputs(6300) <= (layer0_outputs(10101)) and (layer0_outputs(7535));
    outputs(6301) <= (layer0_outputs(9461)) and (layer0_outputs(3058));
    outputs(6302) <= not(layer0_outputs(6336)) or (layer0_outputs(1520));
    outputs(6303) <= not(layer0_outputs(7778));
    outputs(6304) <= layer0_outputs(6326);
    outputs(6305) <= not(layer0_outputs(2349));
    outputs(6306) <= (layer0_outputs(8762)) xor (layer0_outputs(9588));
    outputs(6307) <= not(layer0_outputs(4830));
    outputs(6308) <= layer0_outputs(9139);
    outputs(6309) <= not(layer0_outputs(4527));
    outputs(6310) <= not(layer0_outputs(764));
    outputs(6311) <= not(layer0_outputs(5106));
    outputs(6312) <= layer0_outputs(8699);
    outputs(6313) <= (layer0_outputs(1601)) xor (layer0_outputs(1363));
    outputs(6314) <= (layer0_outputs(5163)) or (layer0_outputs(2079));
    outputs(6315) <= not(layer0_outputs(1259));
    outputs(6316) <= (layer0_outputs(530)) xor (layer0_outputs(242));
    outputs(6317) <= (layer0_outputs(4211)) xor (layer0_outputs(6574));
    outputs(6318) <= layer0_outputs(2410);
    outputs(6319) <= not(layer0_outputs(3506));
    outputs(6320) <= not(layer0_outputs(1618)) or (layer0_outputs(6555));
    outputs(6321) <= layer0_outputs(9310);
    outputs(6322) <= not((layer0_outputs(1303)) or (layer0_outputs(8713)));
    outputs(6323) <= not(layer0_outputs(575));
    outputs(6324) <= not(layer0_outputs(1663));
    outputs(6325) <= not(layer0_outputs(872));
    outputs(6326) <= not((layer0_outputs(5062)) or (layer0_outputs(6870)));
    outputs(6327) <= layer0_outputs(901);
    outputs(6328) <= not((layer0_outputs(9260)) xor (layer0_outputs(7773)));
    outputs(6329) <= layer0_outputs(7186);
    outputs(6330) <= layer0_outputs(6833);
    outputs(6331) <= (layer0_outputs(7881)) xor (layer0_outputs(9576));
    outputs(6332) <= not(layer0_outputs(9939));
    outputs(6333) <= (layer0_outputs(9246)) and not (layer0_outputs(6600));
    outputs(6334) <= layer0_outputs(3085);
    outputs(6335) <= not((layer0_outputs(6569)) or (layer0_outputs(2205)));
    outputs(6336) <= not(layer0_outputs(2386)) or (layer0_outputs(9327));
    outputs(6337) <= (layer0_outputs(2011)) or (layer0_outputs(8046));
    outputs(6338) <= (layer0_outputs(9829)) xor (layer0_outputs(2322));
    outputs(6339) <= not((layer0_outputs(10209)) xor (layer0_outputs(7578)));
    outputs(6340) <= layer0_outputs(5719);
    outputs(6341) <= (layer0_outputs(4554)) or (layer0_outputs(10212));
    outputs(6342) <= not(layer0_outputs(5649));
    outputs(6343) <= (layer0_outputs(3773)) xor (layer0_outputs(2801));
    outputs(6344) <= (layer0_outputs(8221)) xor (layer0_outputs(5236));
    outputs(6345) <= (layer0_outputs(4537)) xor (layer0_outputs(4337));
    outputs(6346) <= not(layer0_outputs(1336));
    outputs(6347) <= not((layer0_outputs(4356)) xor (layer0_outputs(43)));
    outputs(6348) <= (layer0_outputs(711)) and (layer0_outputs(9305));
    outputs(6349) <= (layer0_outputs(97)) and (layer0_outputs(4423));
    outputs(6350) <= not(layer0_outputs(1740));
    outputs(6351) <= layer0_outputs(7207);
    outputs(6352) <= (layer0_outputs(2899)) or (layer0_outputs(4006));
    outputs(6353) <= not(layer0_outputs(9073));
    outputs(6354) <= not(layer0_outputs(5416));
    outputs(6355) <= (layer0_outputs(2579)) and not (layer0_outputs(8160));
    outputs(6356) <= (layer0_outputs(6624)) and not (layer0_outputs(85));
    outputs(6357) <= not(layer0_outputs(5504));
    outputs(6358) <= (layer0_outputs(7039)) and (layer0_outputs(708));
    outputs(6359) <= not(layer0_outputs(300));
    outputs(6360) <= layer0_outputs(5417);
    outputs(6361) <= (layer0_outputs(7419)) xor (layer0_outputs(7323));
    outputs(6362) <= (layer0_outputs(6358)) and not (layer0_outputs(8172));
    outputs(6363) <= (layer0_outputs(2873)) and not (layer0_outputs(3194));
    outputs(6364) <= layer0_outputs(8149);
    outputs(6365) <= layer0_outputs(1077);
    outputs(6366) <= (layer0_outputs(2020)) and not (layer0_outputs(100));
    outputs(6367) <= not(layer0_outputs(5540));
    outputs(6368) <= not((layer0_outputs(2624)) xor (layer0_outputs(2806)));
    outputs(6369) <= not(layer0_outputs(6042));
    outputs(6370) <= (layer0_outputs(406)) or (layer0_outputs(3153));
    outputs(6371) <= (layer0_outputs(7403)) and not (layer0_outputs(2781));
    outputs(6372) <= not(layer0_outputs(5286));
    outputs(6373) <= not((layer0_outputs(4557)) xor (layer0_outputs(10049)));
    outputs(6374) <= (layer0_outputs(5731)) and (layer0_outputs(3504));
    outputs(6375) <= not((layer0_outputs(1523)) xor (layer0_outputs(4662)));
    outputs(6376) <= not(layer0_outputs(5728));
    outputs(6377) <= (layer0_outputs(9108)) and (layer0_outputs(9226));
    outputs(6378) <= layer0_outputs(8271);
    outputs(6379) <= (layer0_outputs(7836)) xor (layer0_outputs(9613));
    outputs(6380) <= (layer0_outputs(1061)) xor (layer0_outputs(5275));
    outputs(6381) <= not((layer0_outputs(4419)) xor (layer0_outputs(8608)));
    outputs(6382) <= (layer0_outputs(1476)) and (layer0_outputs(2072));
    outputs(6383) <= (layer0_outputs(4371)) xor (layer0_outputs(3216));
    outputs(6384) <= not(layer0_outputs(3284));
    outputs(6385) <= layer0_outputs(10068);
    outputs(6386) <= not((layer0_outputs(7464)) xor (layer0_outputs(2178)));
    outputs(6387) <= not(layer0_outputs(7331));
    outputs(6388) <= not(layer0_outputs(3416));
    outputs(6389) <= (layer0_outputs(7730)) and not (layer0_outputs(1631));
    outputs(6390) <= layer0_outputs(7887);
    outputs(6391) <= not(layer0_outputs(9981));
    outputs(6392) <= not(layer0_outputs(5250));
    outputs(6393) <= not((layer0_outputs(4520)) or (layer0_outputs(8543)));
    outputs(6394) <= (layer0_outputs(3425)) or (layer0_outputs(4429));
    outputs(6395) <= not(layer0_outputs(10029));
    outputs(6396) <= not((layer0_outputs(4486)) or (layer0_outputs(6367)));
    outputs(6397) <= not(layer0_outputs(1798));
    outputs(6398) <= not((layer0_outputs(3965)) or (layer0_outputs(6159)));
    outputs(6399) <= (layer0_outputs(7705)) or (layer0_outputs(2174));
    outputs(6400) <= not((layer0_outputs(7262)) xor (layer0_outputs(8648)));
    outputs(6401) <= not(layer0_outputs(3852));
    outputs(6402) <= (layer0_outputs(1471)) or (layer0_outputs(5778));
    outputs(6403) <= not((layer0_outputs(8404)) or (layer0_outputs(6322)));
    outputs(6404) <= not(layer0_outputs(9821));
    outputs(6405) <= (layer0_outputs(630)) and not (layer0_outputs(7611));
    outputs(6406) <= (layer0_outputs(6790)) and (layer0_outputs(5933));
    outputs(6407) <= (layer0_outputs(5137)) xor (layer0_outputs(8082));
    outputs(6408) <= not(layer0_outputs(7335)) or (layer0_outputs(3063));
    outputs(6409) <= not(layer0_outputs(10036));
    outputs(6410) <= (layer0_outputs(683)) and (layer0_outputs(6029));
    outputs(6411) <= (layer0_outputs(5705)) and not (layer0_outputs(4811));
    outputs(6412) <= layer0_outputs(3097);
    outputs(6413) <= (layer0_outputs(5970)) xor (layer0_outputs(5804));
    outputs(6414) <= not(layer0_outputs(1633));
    outputs(6415) <= not(layer0_outputs(5967));
    outputs(6416) <= not(layer0_outputs(7706));
    outputs(6417) <= layer0_outputs(7932);
    outputs(6418) <= (layer0_outputs(8933)) and not (layer0_outputs(2495));
    outputs(6419) <= not(layer0_outputs(9283)) or (layer0_outputs(927));
    outputs(6420) <= (layer0_outputs(5193)) xor (layer0_outputs(2558));
    outputs(6421) <= not((layer0_outputs(149)) or (layer0_outputs(4300)));
    outputs(6422) <= '1';
    outputs(6423) <= (layer0_outputs(7853)) and not (layer0_outputs(423));
    outputs(6424) <= not(layer0_outputs(4548));
    outputs(6425) <= (layer0_outputs(5145)) and not (layer0_outputs(7368));
    outputs(6426) <= (layer0_outputs(7188)) or (layer0_outputs(3520));
    outputs(6427) <= layer0_outputs(8451);
    outputs(6428) <= layer0_outputs(1974);
    outputs(6429) <= not((layer0_outputs(8588)) or (layer0_outputs(4373)));
    outputs(6430) <= not((layer0_outputs(3116)) xor (layer0_outputs(6690)));
    outputs(6431) <= not(layer0_outputs(5958));
    outputs(6432) <= not((layer0_outputs(5162)) or (layer0_outputs(1176)));
    outputs(6433) <= not((layer0_outputs(9307)) or (layer0_outputs(8207)));
    outputs(6434) <= (layer0_outputs(2508)) or (layer0_outputs(1727));
    outputs(6435) <= not((layer0_outputs(4922)) and (layer0_outputs(4618)));
    outputs(6436) <= (layer0_outputs(5963)) xor (layer0_outputs(580));
    outputs(6437) <= not((layer0_outputs(9938)) xor (layer0_outputs(4756)));
    outputs(6438) <= layer0_outputs(10053);
    outputs(6439) <= (layer0_outputs(3277)) and (layer0_outputs(7343));
    outputs(6440) <= not((layer0_outputs(9842)) or (layer0_outputs(1887)));
    outputs(6441) <= not(layer0_outputs(7871));
    outputs(6442) <= (layer0_outputs(9577)) and not (layer0_outputs(3569));
    outputs(6443) <= not(layer0_outputs(2673));
    outputs(6444) <= not(layer0_outputs(1265)) or (layer0_outputs(5961));
    outputs(6445) <= not((layer0_outputs(6985)) xor (layer0_outputs(4085)));
    outputs(6446) <= not(layer0_outputs(106)) or (layer0_outputs(1173));
    outputs(6447) <= (layer0_outputs(1545)) or (layer0_outputs(4323));
    outputs(6448) <= not(layer0_outputs(4010));
    outputs(6449) <= not(layer0_outputs(3368)) or (layer0_outputs(5384));
    outputs(6450) <= layer0_outputs(1757);
    outputs(6451) <= (layer0_outputs(1604)) xor (layer0_outputs(9664));
    outputs(6452) <= not(layer0_outputs(5459));
    outputs(6453) <= layer0_outputs(7042);
    outputs(6454) <= not((layer0_outputs(9019)) xor (layer0_outputs(5817)));
    outputs(6455) <= not((layer0_outputs(359)) xor (layer0_outputs(5352)));
    outputs(6456) <= layer0_outputs(2224);
    outputs(6457) <= not(layer0_outputs(6916));
    outputs(6458) <= (layer0_outputs(4048)) or (layer0_outputs(5287));
    outputs(6459) <= not((layer0_outputs(8729)) or (layer0_outputs(2764)));
    outputs(6460) <= (layer0_outputs(5974)) xor (layer0_outputs(1995));
    outputs(6461) <= (layer0_outputs(8817)) xor (layer0_outputs(1464));
    outputs(6462) <= layer0_outputs(9844);
    outputs(6463) <= (layer0_outputs(3497)) xor (layer0_outputs(8754));
    outputs(6464) <= not((layer0_outputs(7689)) and (layer0_outputs(5048)));
    outputs(6465) <= (layer0_outputs(3447)) xor (layer0_outputs(4639));
    outputs(6466) <= (layer0_outputs(1883)) and not (layer0_outputs(2679));
    outputs(6467) <= (layer0_outputs(5799)) and not (layer0_outputs(7901));
    outputs(6468) <= (layer0_outputs(2445)) xor (layer0_outputs(4991));
    outputs(6469) <= (layer0_outputs(1077)) and (layer0_outputs(582));
    outputs(6470) <= not(layer0_outputs(1898)) or (layer0_outputs(2829));
    outputs(6471) <= (layer0_outputs(7021)) and not (layer0_outputs(8843));
    outputs(6472) <= not(layer0_outputs(271)) or (layer0_outputs(1736));
    outputs(6473) <= layer0_outputs(1376);
    outputs(6474) <= not(layer0_outputs(1005));
    outputs(6475) <= not((layer0_outputs(2683)) xor (layer0_outputs(4588)));
    outputs(6476) <= (layer0_outputs(5138)) and not (layer0_outputs(8373));
    outputs(6477) <= (layer0_outputs(9392)) xor (layer0_outputs(6774));
    outputs(6478) <= layer0_outputs(3794);
    outputs(6479) <= layer0_outputs(3750);
    outputs(6480) <= layer0_outputs(5032);
    outputs(6481) <= not(layer0_outputs(8552)) or (layer0_outputs(4288));
    outputs(6482) <= (layer0_outputs(5612)) xor (layer0_outputs(7903));
    outputs(6483) <= (layer0_outputs(3026)) and (layer0_outputs(374));
    outputs(6484) <= layer0_outputs(114);
    outputs(6485) <= not((layer0_outputs(8550)) or (layer0_outputs(2402)));
    outputs(6486) <= not(layer0_outputs(1877));
    outputs(6487) <= not((layer0_outputs(5872)) and (layer0_outputs(1375)));
    outputs(6488) <= not(layer0_outputs(1294));
    outputs(6489) <= layer0_outputs(9565);
    outputs(6490) <= layer0_outputs(6419);
    outputs(6491) <= not(layer0_outputs(3508));
    outputs(6492) <= (layer0_outputs(1985)) xor (layer0_outputs(4132));
    outputs(6493) <= not((layer0_outputs(9937)) or (layer0_outputs(9152)));
    outputs(6494) <= (layer0_outputs(3031)) and (layer0_outputs(5877));
    outputs(6495) <= (layer0_outputs(4541)) and not (layer0_outputs(5477));
    outputs(6496) <= not((layer0_outputs(7718)) xor (layer0_outputs(3937)));
    outputs(6497) <= not(layer0_outputs(4899));
    outputs(6498) <= (layer0_outputs(2018)) and (layer0_outputs(2117));
    outputs(6499) <= (layer0_outputs(10080)) xor (layer0_outputs(4501));
    outputs(6500) <= (layer0_outputs(7916)) and not (layer0_outputs(10199));
    outputs(6501) <= not(layer0_outputs(1598));
    outputs(6502) <= layer0_outputs(9641);
    outputs(6503) <= layer0_outputs(2575);
    outputs(6504) <= layer0_outputs(5509);
    outputs(6505) <= (layer0_outputs(5001)) and (layer0_outputs(9806));
    outputs(6506) <= not((layer0_outputs(3657)) and (layer0_outputs(3994)));
    outputs(6507) <= not(layer0_outputs(6768));
    outputs(6508) <= (layer0_outputs(6178)) and (layer0_outputs(9754));
    outputs(6509) <= (layer0_outputs(5947)) xor (layer0_outputs(407));
    outputs(6510) <= not(layer0_outputs(9167));
    outputs(6511) <= not((layer0_outputs(8129)) or (layer0_outputs(7402)));
    outputs(6512) <= (layer0_outputs(8872)) xor (layer0_outputs(5644));
    outputs(6513) <= not((layer0_outputs(1853)) xor (layer0_outputs(7503)));
    outputs(6514) <= not(layer0_outputs(3211));
    outputs(6515) <= layer0_outputs(7527);
    outputs(6516) <= not(layer0_outputs(7274));
    outputs(6517) <= (layer0_outputs(2172)) or (layer0_outputs(8194));
    outputs(6518) <= (layer0_outputs(1164)) and not (layer0_outputs(4978));
    outputs(6519) <= not(layer0_outputs(1417));
    outputs(6520) <= not(layer0_outputs(7112));
    outputs(6521) <= layer0_outputs(1382);
    outputs(6522) <= (layer0_outputs(2811)) xor (layer0_outputs(3875));
    outputs(6523) <= not((layer0_outputs(5278)) xor (layer0_outputs(2121)));
    outputs(6524) <= (layer0_outputs(2490)) xor (layer0_outputs(7523));
    outputs(6525) <= not(layer0_outputs(6288)) or (layer0_outputs(2352));
    outputs(6526) <= layer0_outputs(3096);
    outputs(6527) <= (layer0_outputs(6602)) and not (layer0_outputs(10090));
    outputs(6528) <= not(layer0_outputs(5438));
    outputs(6529) <= not(layer0_outputs(670));
    outputs(6530) <= layer0_outputs(3831);
    outputs(6531) <= not((layer0_outputs(9851)) or (layer0_outputs(75)));
    outputs(6532) <= not(layer0_outputs(8464));
    outputs(6533) <= (layer0_outputs(8696)) xor (layer0_outputs(8674));
    outputs(6534) <= layer0_outputs(2175);
    outputs(6535) <= '0';
    outputs(6536) <= not(layer0_outputs(9704));
    outputs(6537) <= not(layer0_outputs(2489));
    outputs(6538) <= not((layer0_outputs(4217)) or (layer0_outputs(9905)));
    outputs(6539) <= not(layer0_outputs(228));
    outputs(6540) <= layer0_outputs(5774);
    outputs(6541) <= not(layer0_outputs(9375));
    outputs(6542) <= not((layer0_outputs(6029)) xor (layer0_outputs(6650)));
    outputs(6543) <= not(layer0_outputs(6371));
    outputs(6544) <= (layer0_outputs(8227)) xor (layer0_outputs(6350));
    outputs(6545) <= not((layer0_outputs(8150)) xor (layer0_outputs(9485)));
    outputs(6546) <= not((layer0_outputs(7459)) xor (layer0_outputs(4564)));
    outputs(6547) <= (layer0_outputs(4568)) xor (layer0_outputs(946));
    outputs(6548) <= (layer0_outputs(1728)) and (layer0_outputs(3917));
    outputs(6549) <= not((layer0_outputs(7968)) and (layer0_outputs(4823)));
    outputs(6550) <= not((layer0_outputs(1452)) xor (layer0_outputs(6643)));
    outputs(6551) <= layer0_outputs(5661);
    outputs(6552) <= layer0_outputs(2364);
    outputs(6553) <= (layer0_outputs(3302)) xor (layer0_outputs(4178));
    outputs(6554) <= layer0_outputs(4360);
    outputs(6555) <= not(layer0_outputs(604));
    outputs(6556) <= not(layer0_outputs(5830)) or (layer0_outputs(2084));
    outputs(6557) <= layer0_outputs(2366);
    outputs(6558) <= not(layer0_outputs(7518));
    outputs(6559) <= layer0_outputs(5280);
    outputs(6560) <= (layer0_outputs(2360)) and not (layer0_outputs(5295));
    outputs(6561) <= (layer0_outputs(5687)) and (layer0_outputs(629));
    outputs(6562) <= not(layer0_outputs(3817));
    outputs(6563) <= not((layer0_outputs(2001)) xor (layer0_outputs(10128)));
    outputs(6564) <= not(layer0_outputs(9248)) or (layer0_outputs(2802));
    outputs(6565) <= (layer0_outputs(7981)) or (layer0_outputs(4234));
    outputs(6566) <= not((layer0_outputs(3554)) or (layer0_outputs(6837)));
    outputs(6567) <= (layer0_outputs(180)) xor (layer0_outputs(2800));
    outputs(6568) <= (layer0_outputs(8740)) xor (layer0_outputs(6560));
    outputs(6569) <= (layer0_outputs(9492)) xor (layer0_outputs(9412));
    outputs(6570) <= layer0_outputs(5107);
    outputs(6571) <= layer0_outputs(1228);
    outputs(6572) <= layer0_outputs(1313);
    outputs(6573) <= not(layer0_outputs(2165));
    outputs(6574) <= (layer0_outputs(9316)) and (layer0_outputs(5632));
    outputs(6575) <= layer0_outputs(4250);
    outputs(6576) <= not(layer0_outputs(8010));
    outputs(6577) <= not(layer0_outputs(3478));
    outputs(6578) <= layer0_outputs(2303);
    outputs(6579) <= (layer0_outputs(6027)) xor (layer0_outputs(5020));
    outputs(6580) <= layer0_outputs(2125);
    outputs(6581) <= not((layer0_outputs(986)) xor (layer0_outputs(3550)));
    outputs(6582) <= layer0_outputs(9234);
    outputs(6583) <= not(layer0_outputs(8940));
    outputs(6584) <= (layer0_outputs(6085)) and (layer0_outputs(2657));
    outputs(6585) <= not(layer0_outputs(7738));
    outputs(6586) <= not((layer0_outputs(4759)) and (layer0_outputs(5946)));
    outputs(6587) <= not(layer0_outputs(656)) or (layer0_outputs(3708));
    outputs(6588) <= not(layer0_outputs(2760));
    outputs(6589) <= (layer0_outputs(8816)) xor (layer0_outputs(862));
    outputs(6590) <= not(layer0_outputs(1166)) or (layer0_outputs(777));
    outputs(6591) <= not((layer0_outputs(314)) xor (layer0_outputs(9192)));
    outputs(6592) <= not((layer0_outputs(4274)) xor (layer0_outputs(7613)));
    outputs(6593) <= not(layer0_outputs(8375));
    outputs(6594) <= layer0_outputs(6733);
    outputs(6595) <= '0';
    outputs(6596) <= (layer0_outputs(5809)) or (layer0_outputs(6740));
    outputs(6597) <= (layer0_outputs(9564)) xor (layer0_outputs(8494));
    outputs(6598) <= layer0_outputs(8347);
    outputs(6599) <= not((layer0_outputs(6961)) or (layer0_outputs(5471)));
    outputs(6600) <= layer0_outputs(9515);
    outputs(6601) <= not(layer0_outputs(6151));
    outputs(6602) <= (layer0_outputs(7978)) and not (layer0_outputs(6254));
    outputs(6603) <= layer0_outputs(7679);
    outputs(6604) <= layer0_outputs(5132);
    outputs(6605) <= layer0_outputs(3737);
    outputs(6606) <= not(layer0_outputs(3561));
    outputs(6607) <= not(layer0_outputs(8667));
    outputs(6608) <= (layer0_outputs(8886)) and not (layer0_outputs(7960));
    outputs(6609) <= not(layer0_outputs(35)) or (layer0_outputs(2162));
    outputs(6610) <= (layer0_outputs(7687)) or (layer0_outputs(8154));
    outputs(6611) <= not((layer0_outputs(4900)) xor (layer0_outputs(540)));
    outputs(6612) <= (layer0_outputs(1094)) xor (layer0_outputs(7270));
    outputs(6613) <= not(layer0_outputs(2799));
    outputs(6614) <= not(layer0_outputs(6125));
    outputs(6615) <= layer0_outputs(3921);
    outputs(6616) <= not(layer0_outputs(6467)) or (layer0_outputs(721));
    outputs(6617) <= not(layer0_outputs(2821));
    outputs(6618) <= not(layer0_outputs(1348));
    outputs(6619) <= layer0_outputs(2412);
    outputs(6620) <= (layer0_outputs(105)) and (layer0_outputs(910));
    outputs(6621) <= not((layer0_outputs(9507)) xor (layer0_outputs(4794)));
    outputs(6622) <= (layer0_outputs(6487)) and not (layer0_outputs(6661));
    outputs(6623) <= layer0_outputs(5818);
    outputs(6624) <= not(layer0_outputs(1475));
    outputs(6625) <= (layer0_outputs(905)) and (layer0_outputs(1753));
    outputs(6626) <= layer0_outputs(7958);
    outputs(6627) <= (layer0_outputs(5405)) xor (layer0_outputs(3917));
    outputs(6628) <= not((layer0_outputs(4969)) xor (layer0_outputs(8695)));
    outputs(6629) <= (layer0_outputs(4738)) or (layer0_outputs(681));
    outputs(6630) <= not((layer0_outputs(5653)) xor (layer0_outputs(7798)));
    outputs(6631) <= not(layer0_outputs(8589)) or (layer0_outputs(679));
    outputs(6632) <= layer0_outputs(5679);
    outputs(6633) <= (layer0_outputs(3664)) xor (layer0_outputs(3441));
    outputs(6634) <= layer0_outputs(7760);
    outputs(6635) <= layer0_outputs(2752);
    outputs(6636) <= (layer0_outputs(8019)) and (layer0_outputs(6141));
    outputs(6637) <= not((layer0_outputs(7374)) xor (layer0_outputs(2804)));
    outputs(6638) <= layer0_outputs(2058);
    outputs(6639) <= (layer0_outputs(20)) and (layer0_outputs(1862));
    outputs(6640) <= not(layer0_outputs(8383)) or (layer0_outputs(5968));
    outputs(6641) <= layer0_outputs(9911);
    outputs(6642) <= (layer0_outputs(9675)) xor (layer0_outputs(2972));
    outputs(6643) <= not(layer0_outputs(1053));
    outputs(6644) <= not(layer0_outputs(6491));
    outputs(6645) <= (layer0_outputs(4124)) xor (layer0_outputs(5298));
    outputs(6646) <= layer0_outputs(6031);
    outputs(6647) <= (layer0_outputs(5781)) and not (layer0_outputs(1053));
    outputs(6648) <= not(layer0_outputs(1989));
    outputs(6649) <= (layer0_outputs(10057)) and not (layer0_outputs(222));
    outputs(6650) <= not(layer0_outputs(9078));
    outputs(6651) <= not(layer0_outputs(3513));
    outputs(6652) <= not(layer0_outputs(4944));
    outputs(6653) <= layer0_outputs(9684);
    outputs(6654) <= not(layer0_outputs(3713));
    outputs(6655) <= not(layer0_outputs(5495)) or (layer0_outputs(3702));
    outputs(6656) <= layer0_outputs(1874);
    outputs(6657) <= '1';
    outputs(6658) <= not((layer0_outputs(8616)) xor (layer0_outputs(9881)));
    outputs(6659) <= layer0_outputs(3748);
    outputs(6660) <= not((layer0_outputs(1546)) or (layer0_outputs(2403)));
    outputs(6661) <= (layer0_outputs(5265)) and not (layer0_outputs(4157));
    outputs(6662) <= layer0_outputs(2608);
    outputs(6663) <= (layer0_outputs(130)) and (layer0_outputs(8134));
    outputs(6664) <= not((layer0_outputs(2299)) or (layer0_outputs(7118)));
    outputs(6665) <= not((layer0_outputs(8889)) xor (layer0_outputs(6305)));
    outputs(6666) <= (layer0_outputs(5918)) xor (layer0_outputs(9123));
    outputs(6667) <= not(layer0_outputs(7228));
    outputs(6668) <= not(layer0_outputs(7483));
    outputs(6669) <= not(layer0_outputs(6216));
    outputs(6670) <= layer0_outputs(6873);
    outputs(6671) <= (layer0_outputs(8630)) and (layer0_outputs(8560));
    outputs(6672) <= (layer0_outputs(8268)) xor (layer0_outputs(2679));
    outputs(6673) <= (layer0_outputs(1925)) and (layer0_outputs(6683));
    outputs(6674) <= (layer0_outputs(1034)) and not (layer0_outputs(2708));
    outputs(6675) <= (layer0_outputs(3951)) xor (layer0_outputs(8886));
    outputs(6676) <= not(layer0_outputs(6899));
    outputs(6677) <= layer0_outputs(8310);
    outputs(6678) <= not(layer0_outputs(7700)) or (layer0_outputs(1868));
    outputs(6679) <= not(layer0_outputs(1247));
    outputs(6680) <= layer0_outputs(1122);
    outputs(6681) <= not((layer0_outputs(4693)) or (layer0_outputs(154)));
    outputs(6682) <= (layer0_outputs(894)) and (layer0_outputs(6895));
    outputs(6683) <= not(layer0_outputs(9188));
    outputs(6684) <= layer0_outputs(3474);
    outputs(6685) <= layer0_outputs(9022);
    outputs(6686) <= (layer0_outputs(7347)) and not (layer0_outputs(7232));
    outputs(6687) <= layer0_outputs(4806);
    outputs(6688) <= (layer0_outputs(8477)) and not (layer0_outputs(449));
    outputs(6689) <= layer0_outputs(537);
    outputs(6690) <= not(layer0_outputs(1594)) or (layer0_outputs(4663));
    outputs(6691) <= (layer0_outputs(7272)) or (layer0_outputs(45));
    outputs(6692) <= layer0_outputs(1615);
    outputs(6693) <= (layer0_outputs(6515)) and not (layer0_outputs(9384));
    outputs(6694) <= not(layer0_outputs(4469));
    outputs(6695) <= (layer0_outputs(59)) xor (layer0_outputs(4357));
    outputs(6696) <= (layer0_outputs(7084)) xor (layer0_outputs(4542));
    outputs(6697) <= (layer0_outputs(2204)) and not (layer0_outputs(8645));
    outputs(6698) <= layer0_outputs(7599);
    outputs(6699) <= not(layer0_outputs(2644));
    outputs(6700) <= (layer0_outputs(4185)) xor (layer0_outputs(4566));
    outputs(6701) <= (layer0_outputs(6832)) and not (layer0_outputs(5537));
    outputs(6702) <= layer0_outputs(6627);
    outputs(6703) <= not((layer0_outputs(5975)) or (layer0_outputs(732)));
    outputs(6704) <= (layer0_outputs(5184)) and not (layer0_outputs(9200));
    outputs(6705) <= not((layer0_outputs(7274)) or (layer0_outputs(9912)));
    outputs(6706) <= layer0_outputs(8276);
    outputs(6707) <= not(layer0_outputs(3689));
    outputs(6708) <= not((layer0_outputs(6985)) xor (layer0_outputs(8241)));
    outputs(6709) <= not(layer0_outputs(2833));
    outputs(6710) <= layer0_outputs(783);
    outputs(6711) <= not(layer0_outputs(8072));
    outputs(6712) <= layer0_outputs(1121);
    outputs(6713) <= not(layer0_outputs(5951));
    outputs(6714) <= layer0_outputs(9983);
    outputs(6715) <= layer0_outputs(9991);
    outputs(6716) <= (layer0_outputs(2763)) xor (layer0_outputs(6707));
    outputs(6717) <= not(layer0_outputs(10055));
    outputs(6718) <= layer0_outputs(5110);
    outputs(6719) <= (layer0_outputs(9341)) xor (layer0_outputs(9155));
    outputs(6720) <= '0';
    outputs(6721) <= layer0_outputs(4292);
    outputs(6722) <= (layer0_outputs(4622)) xor (layer0_outputs(1177));
    outputs(6723) <= layer0_outputs(1794);
    outputs(6724) <= layer0_outputs(5687);
    outputs(6725) <= not(layer0_outputs(4668));
    outputs(6726) <= not((layer0_outputs(410)) or (layer0_outputs(7743)));
    outputs(6727) <= (layer0_outputs(1530)) xor (layer0_outputs(1519));
    outputs(6728) <= (layer0_outputs(8457)) xor (layer0_outputs(3575));
    outputs(6729) <= (layer0_outputs(482)) and (layer0_outputs(2545));
    outputs(6730) <= not(layer0_outputs(6047)) or (layer0_outputs(8553));
    outputs(6731) <= (layer0_outputs(9440)) and not (layer0_outputs(3256));
    outputs(6732) <= layer0_outputs(8341);
    outputs(6733) <= not((layer0_outputs(321)) xor (layer0_outputs(1374)));
    outputs(6734) <= layer0_outputs(8938);
    outputs(6735) <= (layer0_outputs(5010)) xor (layer0_outputs(9740));
    outputs(6736) <= layer0_outputs(1917);
    outputs(6737) <= (layer0_outputs(1911)) and (layer0_outputs(2384));
    outputs(6738) <= layer0_outputs(9428);
    outputs(6739) <= layer0_outputs(2538);
    outputs(6740) <= not((layer0_outputs(7865)) or (layer0_outputs(1271)));
    outputs(6741) <= not(layer0_outputs(2989));
    outputs(6742) <= (layer0_outputs(5653)) and not (layer0_outputs(6080));
    outputs(6743) <= not(layer0_outputs(5416));
    outputs(6744) <= layer0_outputs(9886);
    outputs(6745) <= not(layer0_outputs(5808)) or (layer0_outputs(1658));
    outputs(6746) <= layer0_outputs(5430);
    outputs(6747) <= layer0_outputs(9798);
    outputs(6748) <= layer0_outputs(4603);
    outputs(6749) <= (layer0_outputs(4139)) or (layer0_outputs(9505));
    outputs(6750) <= (layer0_outputs(5069)) and (layer0_outputs(7422));
    outputs(6751) <= (layer0_outputs(4870)) and not (layer0_outputs(2495));
    outputs(6752) <= not((layer0_outputs(6772)) xor (layer0_outputs(9161)));
    outputs(6753) <= not((layer0_outputs(10210)) or (layer0_outputs(14)));
    outputs(6754) <= (layer0_outputs(6716)) and not (layer0_outputs(1988));
    outputs(6755) <= not((layer0_outputs(2399)) and (layer0_outputs(4901)));
    outputs(6756) <= not(layer0_outputs(461));
    outputs(6757) <= not(layer0_outputs(8346)) or (layer0_outputs(8112));
    outputs(6758) <= not((layer0_outputs(6633)) or (layer0_outputs(3479)));
    outputs(6759) <= (layer0_outputs(5050)) and (layer0_outputs(6936));
    outputs(6760) <= (layer0_outputs(3428)) or (layer0_outputs(5795));
    outputs(6761) <= layer0_outputs(7506);
    outputs(6762) <= not((layer0_outputs(9642)) xor (layer0_outputs(6941)));
    outputs(6763) <= layer0_outputs(2336);
    outputs(6764) <= layer0_outputs(9317);
    outputs(6765) <= not((layer0_outputs(6631)) xor (layer0_outputs(2168)));
    outputs(6766) <= not((layer0_outputs(8907)) xor (layer0_outputs(4856)));
    outputs(6767) <= layer0_outputs(8135);
    outputs(6768) <= (layer0_outputs(603)) and (layer0_outputs(1656));
    outputs(6769) <= not((layer0_outputs(3736)) and (layer0_outputs(5483)));
    outputs(6770) <= not(layer0_outputs(2239));
    outputs(6771) <= layer0_outputs(8693);
    outputs(6772) <= not((layer0_outputs(4099)) and (layer0_outputs(2031)));
    outputs(6773) <= layer0_outputs(3874);
    outputs(6774) <= layer0_outputs(6362);
    outputs(6775) <= not(layer0_outputs(1765));
    outputs(6776) <= (layer0_outputs(6861)) and not (layer0_outputs(226));
    outputs(6777) <= (layer0_outputs(1436)) and not (layer0_outputs(5255));
    outputs(6778) <= not(layer0_outputs(1316));
    outputs(6779) <= not(layer0_outputs(8661));
    outputs(6780) <= not(layer0_outputs(1323));
    outputs(6781) <= (layer0_outputs(1421)) xor (layer0_outputs(1031));
    outputs(6782) <= not(layer0_outputs(2387));
    outputs(6783) <= not(layer0_outputs(1076));
    outputs(6784) <= (layer0_outputs(1539)) and not (layer0_outputs(9021));
    outputs(6785) <= layer0_outputs(4327);
    outputs(6786) <= not(layer0_outputs(6634));
    outputs(6787) <= layer0_outputs(9395);
    outputs(6788) <= (layer0_outputs(5742)) and not (layer0_outputs(6888));
    outputs(6789) <= (layer0_outputs(1236)) xor (layer0_outputs(1983));
    outputs(6790) <= (layer0_outputs(638)) and (layer0_outputs(6976));
    outputs(6791) <= layer0_outputs(7054);
    outputs(6792) <= not((layer0_outputs(5896)) xor (layer0_outputs(3149)));
    outputs(6793) <= not((layer0_outputs(4892)) xor (layer0_outputs(9602)));
    outputs(6794) <= not(layer0_outputs(587));
    outputs(6795) <= (layer0_outputs(7605)) xor (layer0_outputs(4148));
    outputs(6796) <= layer0_outputs(4997);
    outputs(6797) <= not((layer0_outputs(7360)) and (layer0_outputs(329)));
    outputs(6798) <= not((layer0_outputs(2328)) xor (layer0_outputs(5982)));
    outputs(6799) <= not(layer0_outputs(9898)) or (layer0_outputs(4417));
    outputs(6800) <= not((layer0_outputs(9028)) or (layer0_outputs(7931)));
    outputs(6801) <= not((layer0_outputs(9529)) xor (layer0_outputs(1237)));
    outputs(6802) <= (layer0_outputs(9831)) and not (layer0_outputs(1606));
    outputs(6803) <= not(layer0_outputs(7637));
    outputs(6804) <= (layer0_outputs(10083)) xor (layer0_outputs(3693));
    outputs(6805) <= not(layer0_outputs(3033)) or (layer0_outputs(9865));
    outputs(6806) <= layer0_outputs(1826);
    outputs(6807) <= layer0_outputs(6121);
    outputs(6808) <= not((layer0_outputs(5946)) xor (layer0_outputs(5173)));
    outputs(6809) <= (layer0_outputs(1079)) and not (layer0_outputs(10159));
    outputs(6810) <= (layer0_outputs(2331)) and (layer0_outputs(2017));
    outputs(6811) <= not((layer0_outputs(3820)) xor (layer0_outputs(9220)));
    outputs(6812) <= layer0_outputs(9982);
    outputs(6813) <= (layer0_outputs(7448)) xor (layer0_outputs(3056));
    outputs(6814) <= layer0_outputs(7237);
    outputs(6815) <= (layer0_outputs(6232)) xor (layer0_outputs(6642));
    outputs(6816) <= not(layer0_outputs(6835)) or (layer0_outputs(3259));
    outputs(6817) <= layer0_outputs(87);
    outputs(6818) <= not(layer0_outputs(6798)) or (layer0_outputs(9715));
    outputs(6819) <= layer0_outputs(2620);
    outputs(6820) <= (layer0_outputs(8633)) or (layer0_outputs(842));
    outputs(6821) <= not(layer0_outputs(5026)) or (layer0_outputs(8834));
    outputs(6822) <= layer0_outputs(5363);
    outputs(6823) <= not((layer0_outputs(9403)) and (layer0_outputs(400)));
    outputs(6824) <= not(layer0_outputs(1212)) or (layer0_outputs(8036));
    outputs(6825) <= layer0_outputs(9218);
    outputs(6826) <= not((layer0_outputs(6567)) xor (layer0_outputs(7576)));
    outputs(6827) <= not(layer0_outputs(884));
    outputs(6828) <= layer0_outputs(3334);
    outputs(6829) <= layer0_outputs(1090);
    outputs(6830) <= layer0_outputs(1585);
    outputs(6831) <= not(layer0_outputs(9657));
    outputs(6832) <= not((layer0_outputs(3309)) xor (layer0_outputs(2327)));
    outputs(6833) <= not(layer0_outputs(7239));
    outputs(6834) <= layer0_outputs(8327);
    outputs(6835) <= not(layer0_outputs(7989));
    outputs(6836) <= not(layer0_outputs(403));
    outputs(6837) <= layer0_outputs(7551);
    outputs(6838) <= (layer0_outputs(9755)) xor (layer0_outputs(2015));
    outputs(6839) <= not(layer0_outputs(4750));
    outputs(6840) <= (layer0_outputs(6110)) and not (layer0_outputs(8778));
    outputs(6841) <= not(layer0_outputs(5351));
    outputs(6842) <= (layer0_outputs(445)) and not (layer0_outputs(7988));
    outputs(6843) <= not(layer0_outputs(5051));
    outputs(6844) <= not(layer0_outputs(3873));
    outputs(6845) <= (layer0_outputs(6249)) xor (layer0_outputs(156));
    outputs(6846) <= not(layer0_outputs(1625));
    outputs(6847) <= (layer0_outputs(6448)) xor (layer0_outputs(2489));
    outputs(6848) <= not((layer0_outputs(8485)) and (layer0_outputs(9399)));
    outputs(6849) <= layer0_outputs(8377);
    outputs(6850) <= layer0_outputs(4691);
    outputs(6851) <= (layer0_outputs(3686)) and (layer0_outputs(5417));
    outputs(6852) <= (layer0_outputs(3744)) or (layer0_outputs(5123));
    outputs(6853) <= not(layer0_outputs(3513)) or (layer0_outputs(9420));
    outputs(6854) <= not(layer0_outputs(5836));
    outputs(6855) <= not(layer0_outputs(3546));
    outputs(6856) <= (layer0_outputs(4144)) and not (layer0_outputs(7720));
    outputs(6857) <= not((layer0_outputs(4916)) xor (layer0_outputs(5346)));
    outputs(6858) <= (layer0_outputs(8254)) and not (layer0_outputs(3431));
    outputs(6859) <= (layer0_outputs(9238)) xor (layer0_outputs(6493));
    outputs(6860) <= layer0_outputs(6040);
    outputs(6861) <= (layer0_outputs(8345)) and not (layer0_outputs(6115));
    outputs(6862) <= not(layer0_outputs(1155));
    outputs(6863) <= layer0_outputs(795);
    outputs(6864) <= not((layer0_outputs(6921)) xor (layer0_outputs(8716)));
    outputs(6865) <= not(layer0_outputs(2673)) or (layer0_outputs(504));
    outputs(6866) <= not(layer0_outputs(7149));
    outputs(6867) <= not((layer0_outputs(4397)) xor (layer0_outputs(1157)));
    outputs(6868) <= layer0_outputs(6481);
    outputs(6869) <= (layer0_outputs(3012)) and (layer0_outputs(1088));
    outputs(6870) <= not(layer0_outputs(6319));
    outputs(6871) <= not(layer0_outputs(5114));
    outputs(6872) <= not(layer0_outputs(2350));
    outputs(6873) <= (layer0_outputs(8486)) xor (layer0_outputs(9988));
    outputs(6874) <= layer0_outputs(5547);
    outputs(6875) <= layer0_outputs(7760);
    outputs(6876) <= not((layer0_outputs(10116)) and (layer0_outputs(4326)));
    outputs(6877) <= (layer0_outputs(6779)) xor (layer0_outputs(5461));
    outputs(6878) <= layer0_outputs(1185);
    outputs(6879) <= (layer0_outputs(1444)) xor (layer0_outputs(3286));
    outputs(6880) <= (layer0_outputs(2928)) xor (layer0_outputs(4158));
    outputs(6881) <= (layer0_outputs(4917)) xor (layer0_outputs(5642));
    outputs(6882) <= not((layer0_outputs(5678)) xor (layer0_outputs(3958)));
    outputs(6883) <= not((layer0_outputs(7774)) and (layer0_outputs(1154)));
    outputs(6884) <= layer0_outputs(7587);
    outputs(6885) <= not(layer0_outputs(3473)) or (layer0_outputs(6982));
    outputs(6886) <= layer0_outputs(409);
    outputs(6887) <= layer0_outputs(4285);
    outputs(6888) <= (layer0_outputs(2559)) and not (layer0_outputs(5327));
    outputs(6889) <= layer0_outputs(5442);
    outputs(6890) <= not(layer0_outputs(1244));
    outputs(6891) <= not(layer0_outputs(1038));
    outputs(6892) <= layer0_outputs(4376);
    outputs(6893) <= not((layer0_outputs(9861)) xor (layer0_outputs(9623)));
    outputs(6894) <= not((layer0_outputs(7584)) xor (layer0_outputs(6220)));
    outputs(6895) <= (layer0_outputs(2259)) xor (layer0_outputs(5712));
    outputs(6896) <= layer0_outputs(5890);
    outputs(6897) <= not(layer0_outputs(4704));
    outputs(6898) <= layer0_outputs(3963);
    outputs(6899) <= layer0_outputs(1721);
    outputs(6900) <= not(layer0_outputs(8955));
    outputs(6901) <= not((layer0_outputs(891)) xor (layer0_outputs(1292)));
    outputs(6902) <= (layer0_outputs(3977)) and (layer0_outputs(5467));
    outputs(6903) <= not(layer0_outputs(4010));
    outputs(6904) <= layer0_outputs(0);
    outputs(6905) <= not((layer0_outputs(3539)) xor (layer0_outputs(4816)));
    outputs(6906) <= not(layer0_outputs(2403));
    outputs(6907) <= not(layer0_outputs(7880));
    outputs(6908) <= not(layer0_outputs(5309)) or (layer0_outputs(1908));
    outputs(6909) <= not((layer0_outputs(6421)) and (layer0_outputs(4538)));
    outputs(6910) <= not((layer0_outputs(2505)) xor (layer0_outputs(5279)));
    outputs(6911) <= not(layer0_outputs(5414));
    outputs(6912) <= not((layer0_outputs(9549)) xor (layer0_outputs(3087)));
    outputs(6913) <= layer0_outputs(8021);
    outputs(6914) <= not(layer0_outputs(6822));
    outputs(6915) <= layer0_outputs(6252);
    outputs(6916) <= layer0_outputs(1912);
    outputs(6917) <= not(layer0_outputs(6485)) or (layer0_outputs(3937));
    outputs(6918) <= not(layer0_outputs(9249));
    outputs(6919) <= not((layer0_outputs(1548)) or (layer0_outputs(2998)));
    outputs(6920) <= not(layer0_outputs(1509));
    outputs(6921) <= (layer0_outputs(5789)) and not (layer0_outputs(6697));
    outputs(6922) <= not((layer0_outputs(98)) xor (layer0_outputs(7286)));
    outputs(6923) <= layer0_outputs(2107);
    outputs(6924) <= layer0_outputs(6163);
    outputs(6925) <= not((layer0_outputs(8205)) or (layer0_outputs(7810)));
    outputs(6926) <= not((layer0_outputs(4101)) or (layer0_outputs(13)));
    outputs(6927) <= not(layer0_outputs(5348));
    outputs(6928) <= not((layer0_outputs(4051)) xor (layer0_outputs(4073)));
    outputs(6929) <= (layer0_outputs(9374)) xor (layer0_outputs(7621));
    outputs(6930) <= (layer0_outputs(2397)) xor (layer0_outputs(2155));
    outputs(6931) <= (layer0_outputs(9998)) and (layer0_outputs(9873));
    outputs(6932) <= layer0_outputs(5284);
    outputs(6933) <= not((layer0_outputs(2097)) and (layer0_outputs(3429)));
    outputs(6934) <= not((layer0_outputs(8638)) and (layer0_outputs(3790)));
    outputs(6935) <= not(layer0_outputs(7478));
    outputs(6936) <= layer0_outputs(7022);
    outputs(6937) <= not(layer0_outputs(2812));
    outputs(6938) <= (layer0_outputs(6636)) xor (layer0_outputs(2303));
    outputs(6939) <= not(layer0_outputs(4947));
    outputs(6940) <= layer0_outputs(8976);
    outputs(6941) <= (layer0_outputs(1297)) and not (layer0_outputs(7895));
    outputs(6942) <= not(layer0_outputs(2907));
    outputs(6943) <= not((layer0_outputs(693)) or (layer0_outputs(2355)));
    outputs(6944) <= not(layer0_outputs(8284));
    outputs(6945) <= not((layer0_outputs(7855)) xor (layer0_outputs(7196)));
    outputs(6946) <= not(layer0_outputs(5171)) or (layer0_outputs(4911));
    outputs(6947) <= not((layer0_outputs(8639)) xor (layer0_outputs(5960)));
    outputs(6948) <= layer0_outputs(2079);
    outputs(6949) <= not((layer0_outputs(2888)) xor (layer0_outputs(7386)));
    outputs(6950) <= (layer0_outputs(7729)) and not (layer0_outputs(5468));
    outputs(6951) <= not(layer0_outputs(5825)) or (layer0_outputs(5069));
    outputs(6952) <= not((layer0_outputs(6664)) xor (layer0_outputs(1776)));
    outputs(6953) <= layer0_outputs(2449);
    outputs(6954) <= layer0_outputs(4259);
    outputs(6955) <= not(layer0_outputs(9699));
    outputs(6956) <= not(layer0_outputs(6859));
    outputs(6957) <= not(layer0_outputs(2574)) or (layer0_outputs(2084));
    outputs(6958) <= (layer0_outputs(7881)) and not (layer0_outputs(2129));
    outputs(6959) <= (layer0_outputs(4746)) xor (layer0_outputs(8446));
    outputs(6960) <= not(layer0_outputs(3607));
    outputs(6961) <= not((layer0_outputs(2772)) or (layer0_outputs(7931)));
    outputs(6962) <= (layer0_outputs(7572)) and (layer0_outputs(1508));
    outputs(6963) <= not(layer0_outputs(8939));
    outputs(6964) <= layer0_outputs(5365);
    outputs(6965) <= not(layer0_outputs(5064));
    outputs(6966) <= layer0_outputs(9805);
    outputs(6967) <= not((layer0_outputs(921)) xor (layer0_outputs(1833)));
    outputs(6968) <= (layer0_outputs(6106)) and (layer0_outputs(8127));
    outputs(6969) <= layer0_outputs(1386);
    outputs(6970) <= layer0_outputs(8469);
    outputs(6971) <= not(layer0_outputs(9386));
    outputs(6972) <= not(layer0_outputs(2383));
    outputs(6973) <= layer0_outputs(1906);
    outputs(6974) <= (layer0_outputs(2136)) and (layer0_outputs(5230));
    outputs(6975) <= not(layer0_outputs(9866));
    outputs(6976) <= (layer0_outputs(1103)) xor (layer0_outputs(6305));
    outputs(6977) <= not((layer0_outputs(511)) xor (layer0_outputs(4707)));
    outputs(6978) <= (layer0_outputs(8114)) and not (layer0_outputs(3805));
    outputs(6979) <= not((layer0_outputs(7732)) or (layer0_outputs(3766)));
    outputs(6980) <= not(layer0_outputs(1041)) or (layer0_outputs(268));
    outputs(6981) <= (layer0_outputs(2428)) and not (layer0_outputs(2793));
    outputs(6982) <= not((layer0_outputs(7628)) xor (layer0_outputs(268)));
    outputs(6983) <= not((layer0_outputs(3361)) or (layer0_outputs(3669)));
    outputs(6984) <= not((layer0_outputs(3786)) xor (layer0_outputs(3705)));
    outputs(6985) <= not((layer0_outputs(2290)) xor (layer0_outputs(3646)));
    outputs(6986) <= not(layer0_outputs(1370));
    outputs(6987) <= not((layer0_outputs(2370)) xor (layer0_outputs(3307)));
    outputs(6988) <= not(layer0_outputs(9187));
    outputs(6989) <= not(layer0_outputs(9931));
    outputs(6990) <= layer0_outputs(902);
    outputs(6991) <= (layer0_outputs(2138)) and (layer0_outputs(711));
    outputs(6992) <= not((layer0_outputs(6512)) xor (layer0_outputs(7345)));
    outputs(6993) <= not(layer0_outputs(724)) or (layer0_outputs(3619));
    outputs(6994) <= (layer0_outputs(2515)) and not (layer0_outputs(8748));
    outputs(6995) <= layer0_outputs(6219);
    outputs(6996) <= layer0_outputs(3893);
    outputs(6997) <= layer0_outputs(5565);
    outputs(6998) <= (layer0_outputs(9769)) xor (layer0_outputs(255));
    outputs(6999) <= not(layer0_outputs(4219)) or (layer0_outputs(3577));
    outputs(7000) <= (layer0_outputs(9633)) xor (layer0_outputs(10102));
    outputs(7001) <= not(layer0_outputs(7327));
    outputs(7002) <= not(layer0_outputs(8068));
    outputs(7003) <= layer0_outputs(4022);
    outputs(7004) <= (layer0_outputs(9769)) xor (layer0_outputs(8812));
    outputs(7005) <= layer0_outputs(2914);
    outputs(7006) <= not((layer0_outputs(7772)) and (layer0_outputs(395)));
    outputs(7007) <= (layer0_outputs(5171)) and (layer0_outputs(9227));
    outputs(7008) <= layer0_outputs(6265);
    outputs(7009) <= not((layer0_outputs(9176)) xor (layer0_outputs(1663)));
    outputs(7010) <= (layer0_outputs(9218)) and (layer0_outputs(4502));
    outputs(7011) <= (layer0_outputs(6984)) and not (layer0_outputs(4732));
    outputs(7012) <= (layer0_outputs(4285)) and not (layer0_outputs(592));
    outputs(7013) <= not(layer0_outputs(3003));
    outputs(7014) <= layer0_outputs(4985);
    outputs(7015) <= (layer0_outputs(4591)) xor (layer0_outputs(5895));
    outputs(7016) <= not((layer0_outputs(945)) xor (layer0_outputs(4256)));
    outputs(7017) <= (layer0_outputs(5158)) xor (layer0_outputs(7795));
    outputs(7018) <= layer0_outputs(4340);
    outputs(7019) <= (layer0_outputs(9553)) xor (layer0_outputs(4747));
    outputs(7020) <= (layer0_outputs(1523)) xor (layer0_outputs(6395));
    outputs(7021) <= layer0_outputs(8475);
    outputs(7022) <= not(layer0_outputs(3442));
    outputs(7023) <= (layer0_outputs(3895)) and not (layer0_outputs(8898));
    outputs(7024) <= not(layer0_outputs(5520));
    outputs(7025) <= not((layer0_outputs(8969)) xor (layer0_outputs(7762)));
    outputs(7026) <= (layer0_outputs(7269)) and not (layer0_outputs(9627));
    outputs(7027) <= not(layer0_outputs(250));
    outputs(7028) <= not(layer0_outputs(6306));
    outputs(7029) <= not(layer0_outputs(2724));
    outputs(7030) <= not(layer0_outputs(3997));
    outputs(7031) <= (layer0_outputs(917)) and not (layer0_outputs(2285));
    outputs(7032) <= not(layer0_outputs(1596));
    outputs(7033) <= (layer0_outputs(1635)) xor (layer0_outputs(54));
    outputs(7034) <= (layer0_outputs(6860)) and not (layer0_outputs(6955));
    outputs(7035) <= not((layer0_outputs(175)) and (layer0_outputs(5928)));
    outputs(7036) <= not(layer0_outputs(2220));
    outputs(7037) <= (layer0_outputs(4769)) and not (layer0_outputs(1190));
    outputs(7038) <= layer0_outputs(1640);
    outputs(7039) <= layer0_outputs(1731);
    outputs(7040) <= not(layer0_outputs(4060)) or (layer0_outputs(5162));
    outputs(7041) <= layer0_outputs(8687);
    outputs(7042) <= layer0_outputs(8414);
    outputs(7043) <= (layer0_outputs(10191)) and not (layer0_outputs(4314));
    outputs(7044) <= (layer0_outputs(8427)) xor (layer0_outputs(4210));
    outputs(7045) <= not(layer0_outputs(5334));
    outputs(7046) <= not((layer0_outputs(1137)) and (layer0_outputs(7571)));
    outputs(7047) <= not(layer0_outputs(234));
    outputs(7048) <= not((layer0_outputs(7979)) xor (layer0_outputs(3629)));
    outputs(7049) <= (layer0_outputs(8354)) xor (layer0_outputs(8672));
    outputs(7050) <= (layer0_outputs(8906)) or (layer0_outputs(7945));
    outputs(7051) <= (layer0_outputs(2518)) xor (layer0_outputs(41));
    outputs(7052) <= (layer0_outputs(8688)) and not (layer0_outputs(4572));
    outputs(7053) <= not((layer0_outputs(4424)) xor (layer0_outputs(9510)));
    outputs(7054) <= not((layer0_outputs(3880)) xor (layer0_outputs(6619)));
    outputs(7055) <= not(layer0_outputs(5126)) or (layer0_outputs(1057));
    outputs(7056) <= not((layer0_outputs(334)) xor (layer0_outputs(321)));
    outputs(7057) <= (layer0_outputs(2575)) and not (layer0_outputs(3869));
    outputs(7058) <= layer0_outputs(2940);
    outputs(7059) <= not(layer0_outputs(4650));
    outputs(7060) <= not((layer0_outputs(6071)) xor (layer0_outputs(8075)));
    outputs(7061) <= layer0_outputs(680);
    outputs(7062) <= not(layer0_outputs(3982));
    outputs(7063) <= (layer0_outputs(8085)) and (layer0_outputs(10079));
    outputs(7064) <= (layer0_outputs(919)) and not (layer0_outputs(1842));
    outputs(7065) <= layer0_outputs(3564);
    outputs(7066) <= not(layer0_outputs(6166)) or (layer0_outputs(1849));
    outputs(7067) <= layer0_outputs(5623);
    outputs(7068) <= layer0_outputs(5413);
    outputs(7069) <= not(layer0_outputs(1588));
    outputs(7070) <= layer0_outputs(3409);
    outputs(7071) <= not(layer0_outputs(6430));
    outputs(7072) <= (layer0_outputs(6957)) xor (layer0_outputs(3489));
    outputs(7073) <= (layer0_outputs(6482)) xor (layer0_outputs(5258));
    outputs(7074) <= layer0_outputs(8248);
    outputs(7075) <= not(layer0_outputs(3776));
    outputs(7076) <= layer0_outputs(8566);
    outputs(7077) <= not((layer0_outputs(3852)) xor (layer0_outputs(8625)));
    outputs(7078) <= layer0_outputs(6420);
    outputs(7079) <= layer0_outputs(3523);
    outputs(7080) <= layer0_outputs(7059);
    outputs(7081) <= (layer0_outputs(4404)) xor (layer0_outputs(2050));
    outputs(7082) <= (layer0_outputs(5229)) and not (layer0_outputs(1467));
    outputs(7083) <= (layer0_outputs(8723)) and not (layer0_outputs(4677));
    outputs(7084) <= (layer0_outputs(8441)) xor (layer0_outputs(5963));
    outputs(7085) <= not(layer0_outputs(6837)) or (layer0_outputs(4044));
    outputs(7086) <= not(layer0_outputs(5235)) or (layer0_outputs(9072));
    outputs(7087) <= (layer0_outputs(4904)) and not (layer0_outputs(9532));
    outputs(7088) <= not((layer0_outputs(8760)) or (layer0_outputs(4160)));
    outputs(7089) <= not(layer0_outputs(139));
    outputs(7090) <= not(layer0_outputs(5062)) or (layer0_outputs(4007));
    outputs(7091) <= (layer0_outputs(4339)) xor (layer0_outputs(2188));
    outputs(7092) <= (layer0_outputs(3551)) and (layer0_outputs(6795));
    outputs(7093) <= (layer0_outputs(4544)) xor (layer0_outputs(6214));
    outputs(7094) <= layer0_outputs(284);
    outputs(7095) <= not(layer0_outputs(3510));
    outputs(7096) <= not(layer0_outputs(4642));
    outputs(7097) <= layer0_outputs(8043);
    outputs(7098) <= layer0_outputs(3166);
    outputs(7099) <= (layer0_outputs(2887)) and not (layer0_outputs(8051));
    outputs(7100) <= layer0_outputs(6638);
    outputs(7101) <= not(layer0_outputs(6569));
    outputs(7102) <= (layer0_outputs(9839)) and (layer0_outputs(6708));
    outputs(7103) <= not(layer0_outputs(1804));
    outputs(7104) <= layer0_outputs(3383);
    outputs(7105) <= not((layer0_outputs(9284)) xor (layer0_outputs(7524)));
    outputs(7106) <= (layer0_outputs(1122)) xor (layer0_outputs(7722));
    outputs(7107) <= (layer0_outputs(6000)) and not (layer0_outputs(9186));
    outputs(7108) <= (layer0_outputs(3259)) xor (layer0_outputs(8176));
    outputs(7109) <= (layer0_outputs(2815)) and (layer0_outputs(2888));
    outputs(7110) <= not(layer0_outputs(5478));
    outputs(7111) <= not(layer0_outputs(8874));
    outputs(7112) <= not((layer0_outputs(3278)) xor (layer0_outputs(1327)));
    outputs(7113) <= not(layer0_outputs(5037));
    outputs(7114) <= (layer0_outputs(6045)) xor (layer0_outputs(5435));
    outputs(7115) <= (layer0_outputs(9189)) xor (layer0_outputs(9604));
    outputs(7116) <= not((layer0_outputs(5270)) and (layer0_outputs(7220)));
    outputs(7117) <= (layer0_outputs(804)) xor (layer0_outputs(5733));
    outputs(7118) <= not(layer0_outputs(9009));
    outputs(7119) <= not(layer0_outputs(9958));
    outputs(7120) <= (layer0_outputs(8654)) xor (layer0_outputs(4919));
    outputs(7121) <= layer0_outputs(6008);
    outputs(7122) <= not(layer0_outputs(7255));
    outputs(7123) <= not(layer0_outputs(1093));
    outputs(7124) <= not(layer0_outputs(7898));
    outputs(7125) <= (layer0_outputs(7543)) or (layer0_outputs(8279));
    outputs(7126) <= not((layer0_outputs(2520)) xor (layer0_outputs(8426)));
    outputs(7127) <= (layer0_outputs(7900)) xor (layer0_outputs(1414));
    outputs(7128) <= not(layer0_outputs(5387)) or (layer0_outputs(6621));
    outputs(7129) <= not((layer0_outputs(6827)) xor (layer0_outputs(787)));
    outputs(7130) <= (layer0_outputs(3816)) xor (layer0_outputs(7167));
    outputs(7131) <= not(layer0_outputs(2034));
    outputs(7132) <= (layer0_outputs(9519)) xor (layer0_outputs(10052));
    outputs(7133) <= not(layer0_outputs(2531));
    outputs(7134) <= (layer0_outputs(7875)) and (layer0_outputs(4808));
    outputs(7135) <= not(layer0_outputs(9373));
    outputs(7136) <= not(layer0_outputs(2483));
    outputs(7137) <= (layer0_outputs(2770)) or (layer0_outputs(6171));
    outputs(7138) <= (layer0_outputs(1634)) or (layer0_outputs(2243));
    outputs(7139) <= (layer0_outputs(5214)) xor (layer0_outputs(6732));
    outputs(7140) <= not(layer0_outputs(5949));
    outputs(7141) <= not(layer0_outputs(352));
    outputs(7142) <= (layer0_outputs(5460)) and (layer0_outputs(7124));
    outputs(7143) <= layer0_outputs(546);
    outputs(7144) <= (layer0_outputs(2581)) and not (layer0_outputs(8951));
    outputs(7145) <= layer0_outputs(7945);
    outputs(7146) <= not(layer0_outputs(4077));
    outputs(7147) <= (layer0_outputs(7362)) xor (layer0_outputs(7861));
    outputs(7148) <= not((layer0_outputs(7)) or (layer0_outputs(1367)));
    outputs(7149) <= not((layer0_outputs(4054)) or (layer0_outputs(3164)));
    outputs(7150) <= layer0_outputs(1692);
    outputs(7151) <= not(layer0_outputs(1343));
    outputs(7152) <= not(layer0_outputs(9042));
    outputs(7153) <= not((layer0_outputs(4087)) xor (layer0_outputs(2358)));
    outputs(7154) <= not((layer0_outputs(1837)) xor (layer0_outputs(9667)));
    outputs(7155) <= not((layer0_outputs(1639)) xor (layer0_outputs(4338)));
    outputs(7156) <= (layer0_outputs(5783)) and not (layer0_outputs(8620));
    outputs(7157) <= layer0_outputs(8924);
    outputs(7158) <= layer0_outputs(3511);
    outputs(7159) <= (layer0_outputs(8397)) xor (layer0_outputs(7277));
    outputs(7160) <= layer0_outputs(9490);
    outputs(7161) <= layer0_outputs(2373);
    outputs(7162) <= not((layer0_outputs(7680)) xor (layer0_outputs(4422)));
    outputs(7163) <= layer0_outputs(6149);
    outputs(7164) <= (layer0_outputs(10115)) xor (layer0_outputs(8246));
    outputs(7165) <= layer0_outputs(1150);
    outputs(7166) <= (layer0_outputs(5043)) and not (layer0_outputs(4473));
    outputs(7167) <= not((layer0_outputs(8230)) xor (layer0_outputs(9137)));
    outputs(7168) <= not((layer0_outputs(623)) xor (layer0_outputs(9285)));
    outputs(7169) <= (layer0_outputs(4687)) xor (layer0_outputs(1456));
    outputs(7170) <= (layer0_outputs(1590)) and not (layer0_outputs(3086));
    outputs(7171) <= (layer0_outputs(1510)) and not (layer0_outputs(9886));
    outputs(7172) <= (layer0_outputs(6274)) xor (layer0_outputs(6351));
    outputs(7173) <= (layer0_outputs(1945)) and (layer0_outputs(1978));
    outputs(7174) <= not((layer0_outputs(3093)) xor (layer0_outputs(3679)));
    outputs(7175) <= not((layer0_outputs(1507)) xor (layer0_outputs(3699)));
    outputs(7176) <= (layer0_outputs(1588)) xor (layer0_outputs(6765));
    outputs(7177) <= (layer0_outputs(9153)) and not (layer0_outputs(4357));
    outputs(7178) <= not(layer0_outputs(4460));
    outputs(7179) <= layer0_outputs(2857);
    outputs(7180) <= not(layer0_outputs(7303)) or (layer0_outputs(5931));
    outputs(7181) <= not((layer0_outputs(6568)) xor (layer0_outputs(2999)));
    outputs(7182) <= (layer0_outputs(8408)) and (layer0_outputs(5001));
    outputs(7183) <= layer0_outputs(13);
    outputs(7184) <= not(layer0_outputs(3206));
    outputs(7185) <= not(layer0_outputs(7451));
    outputs(7186) <= not((layer0_outputs(262)) xor (layer0_outputs(6884)));
    outputs(7187) <= (layer0_outputs(1193)) and not (layer0_outputs(8279));
    outputs(7188) <= (layer0_outputs(7012)) and not (layer0_outputs(1498));
    outputs(7189) <= (layer0_outputs(5923)) xor (layer0_outputs(5867));
    outputs(7190) <= not(layer0_outputs(7545)) or (layer0_outputs(9772));
    outputs(7191) <= (layer0_outputs(978)) and (layer0_outputs(2413));
    outputs(7192) <= not(layer0_outputs(10184));
    outputs(7193) <= not((layer0_outputs(7947)) and (layer0_outputs(2272)));
    outputs(7194) <= layer0_outputs(7838);
    outputs(7195) <= not(layer0_outputs(3792));
    outputs(7196) <= not(layer0_outputs(4337));
    outputs(7197) <= layer0_outputs(1190);
    outputs(7198) <= not(layer0_outputs(8487));
    outputs(7199) <= layer0_outputs(2488);
    outputs(7200) <= not((layer0_outputs(8933)) xor (layer0_outputs(4847)));
    outputs(7201) <= not(layer0_outputs(1196));
    outputs(7202) <= not(layer0_outputs(6189));
    outputs(7203) <= (layer0_outputs(1791)) and not (layer0_outputs(5910));
    outputs(7204) <= not(layer0_outputs(796));
    outputs(7205) <= layer0_outputs(1686);
    outputs(7206) <= layer0_outputs(3570);
    outputs(7207) <= (layer0_outputs(1428)) xor (layer0_outputs(1218));
    outputs(7208) <= '1';
    outputs(7209) <= not(layer0_outputs(5473));
    outputs(7210) <= (layer0_outputs(134)) xor (layer0_outputs(4898));
    outputs(7211) <= (layer0_outputs(8519)) xor (layer0_outputs(2083));
    outputs(7212) <= (layer0_outputs(2112)) or (layer0_outputs(8319));
    outputs(7213) <= not((layer0_outputs(444)) or (layer0_outputs(7960)));
    outputs(7214) <= not(layer0_outputs(1696));
    outputs(7215) <= not((layer0_outputs(7222)) xor (layer0_outputs(4148)));
    outputs(7216) <= not((layer0_outputs(5800)) xor (layer0_outputs(4479)));
    outputs(7217) <= not((layer0_outputs(7215)) or (layer0_outputs(4450)));
    outputs(7218) <= layer0_outputs(1);
    outputs(7219) <= not(layer0_outputs(9074));
    outputs(7220) <= not(layer0_outputs(6554)) or (layer0_outputs(4980));
    outputs(7221) <= not(layer0_outputs(4821));
    outputs(7222) <= not(layer0_outputs(3070)) or (layer0_outputs(578));
    outputs(7223) <= not((layer0_outputs(6580)) or (layer0_outputs(8131)));
    outputs(7224) <= not((layer0_outputs(4823)) xor (layer0_outputs(1416)));
    outputs(7225) <= (layer0_outputs(3538)) and not (layer0_outputs(1115));
    outputs(7226) <= (layer0_outputs(6723)) xor (layer0_outputs(4437));
    outputs(7227) <= (layer0_outputs(9050)) xor (layer0_outputs(10031));
    outputs(7228) <= not((layer0_outputs(2795)) xor (layer0_outputs(7759)));
    outputs(7229) <= not(layer0_outputs(5737));
    outputs(7230) <= layer0_outputs(906);
    outputs(7231) <= not(layer0_outputs(1214)) or (layer0_outputs(2505));
    outputs(7232) <= not(layer0_outputs(5019));
    outputs(7233) <= (layer0_outputs(9039)) or (layer0_outputs(59));
    outputs(7234) <= not(layer0_outputs(4167));
    outputs(7235) <= not((layer0_outputs(9657)) xor (layer0_outputs(2475)));
    outputs(7236) <= not(layer0_outputs(4948));
    outputs(7237) <= (layer0_outputs(9209)) xor (layer0_outputs(4859));
    outputs(7238) <= not(layer0_outputs(5676));
    outputs(7239) <= layer0_outputs(4526);
    outputs(7240) <= not(layer0_outputs(5249));
    outputs(7241) <= not(layer0_outputs(6444));
    outputs(7242) <= (layer0_outputs(2057)) and not (layer0_outputs(6339));
    outputs(7243) <= not(layer0_outputs(8975));
    outputs(7244) <= not((layer0_outputs(9608)) or (layer0_outputs(8865)));
    outputs(7245) <= (layer0_outputs(5150)) or (layer0_outputs(4742));
    outputs(7246) <= not((layer0_outputs(1138)) or (layer0_outputs(9848)));
    outputs(7247) <= not(layer0_outputs(5621));
    outputs(7248) <= layer0_outputs(1317);
    outputs(7249) <= not((layer0_outputs(8273)) or (layer0_outputs(1404)));
    outputs(7250) <= layer0_outputs(4503);
    outputs(7251) <= layer0_outputs(8883);
    outputs(7252) <= (layer0_outputs(9207)) xor (layer0_outputs(7114));
    outputs(7253) <= (layer0_outputs(8378)) and not (layer0_outputs(1315));
    outputs(7254) <= not(layer0_outputs(3041));
    outputs(7255) <= layer0_outputs(2005);
    outputs(7256) <= not(layer0_outputs(5820));
    outputs(7257) <= not(layer0_outputs(4170));
    outputs(7258) <= not(layer0_outputs(8458));
    outputs(7259) <= (layer0_outputs(4084)) and not (layer0_outputs(5718));
    outputs(7260) <= layer0_outputs(1358);
    outputs(7261) <= not(layer0_outputs(2133));
    outputs(7262) <= not((layer0_outputs(7242)) xor (layer0_outputs(10022)));
    outputs(7263) <= not((layer0_outputs(433)) or (layer0_outputs(5190)));
    outputs(7264) <= not((layer0_outputs(9166)) or (layer0_outputs(8111)));
    outputs(7265) <= not((layer0_outputs(5312)) xor (layer0_outputs(7768)));
    outputs(7266) <= not((layer0_outputs(2305)) xor (layer0_outputs(8361)));
    outputs(7267) <= layer0_outputs(8860);
    outputs(7268) <= (layer0_outputs(6431)) xor (layer0_outputs(7485));
    outputs(7269) <= not(layer0_outputs(1757));
    outputs(7270) <= not(layer0_outputs(1827)) or (layer0_outputs(156));
    outputs(7271) <= not((layer0_outputs(5854)) xor (layer0_outputs(9158)));
    outputs(7272) <= layer0_outputs(9054);
    outputs(7273) <= (layer0_outputs(3458)) and not (layer0_outputs(5737));
    outputs(7274) <= not(layer0_outputs(3605));
    outputs(7275) <= not(layer0_outputs(2701));
    outputs(7276) <= layer0_outputs(7317);
    outputs(7277) <= (layer0_outputs(8285)) xor (layer0_outputs(6906));
    outputs(7278) <= not((layer0_outputs(3171)) or (layer0_outputs(2517)));
    outputs(7279) <= not(layer0_outputs(2010));
    outputs(7280) <= not((layer0_outputs(9913)) xor (layer0_outputs(720)));
    outputs(7281) <= not((layer0_outputs(6873)) xor (layer0_outputs(9229)));
    outputs(7282) <= (layer0_outputs(9675)) xor (layer0_outputs(7751));
    outputs(7283) <= not((layer0_outputs(9295)) xor (layer0_outputs(6574)));
    outputs(7284) <= not(layer0_outputs(1771)) or (layer0_outputs(8984));
    outputs(7285) <= not(layer0_outputs(9435));
    outputs(7286) <= not(layer0_outputs(9393)) or (layer0_outputs(7032));
    outputs(7287) <= (layer0_outputs(6486)) and not (layer0_outputs(29));
    outputs(7288) <= (layer0_outputs(384)) and not (layer0_outputs(58));
    outputs(7289) <= (layer0_outputs(6437)) and not (layer0_outputs(985));
    outputs(7290) <= not(layer0_outputs(6865));
    outputs(7291) <= not((layer0_outputs(5560)) xor (layer0_outputs(1752)));
    outputs(7292) <= layer0_outputs(7043);
    outputs(7293) <= (layer0_outputs(4238)) and (layer0_outputs(9348));
    outputs(7294) <= layer0_outputs(2327);
    outputs(7295) <= (layer0_outputs(3662)) xor (layer0_outputs(6809));
    outputs(7296) <= layer0_outputs(1021);
    outputs(7297) <= (layer0_outputs(2809)) and not (layer0_outputs(8137));
    outputs(7298) <= (layer0_outputs(4570)) or (layer0_outputs(3105));
    outputs(7299) <= layer0_outputs(8684);
    outputs(7300) <= not(layer0_outputs(5107));
    outputs(7301) <= not((layer0_outputs(4731)) or (layer0_outputs(5993)));
    outputs(7302) <= layer0_outputs(6694);
    outputs(7303) <= not(layer0_outputs(7977)) or (layer0_outputs(634));
    outputs(7304) <= layer0_outputs(1955);
    outputs(7305) <= not(layer0_outputs(8707));
    outputs(7306) <= layer0_outputs(529);
    outputs(7307) <= (layer0_outputs(8819)) and (layer0_outputs(1680));
    outputs(7308) <= not(layer0_outputs(8658));
    outputs(7309) <= not((layer0_outputs(5929)) xor (layer0_outputs(4160)));
    outputs(7310) <= layer0_outputs(160);
    outputs(7311) <= layer0_outputs(4886);
    outputs(7312) <= not((layer0_outputs(7894)) xor (layer0_outputs(7028)));
    outputs(7313) <= (layer0_outputs(7905)) and not (layer0_outputs(5248));
    outputs(7314) <= layer0_outputs(6507);
    outputs(7315) <= layer0_outputs(10074);
    outputs(7316) <= not(layer0_outputs(5716)) or (layer0_outputs(3825));
    outputs(7317) <= (layer0_outputs(5378)) xor (layer0_outputs(8876));
    outputs(7318) <= not((layer0_outputs(6074)) xor (layer0_outputs(1909)));
    outputs(7319) <= not((layer0_outputs(10168)) xor (layer0_outputs(5298)));
    outputs(7320) <= (layer0_outputs(7294)) or (layer0_outputs(4714));
    outputs(7321) <= (layer0_outputs(1744)) xor (layer0_outputs(9179));
    outputs(7322) <= (layer0_outputs(7327)) and not (layer0_outputs(2063));
    outputs(7323) <= not(layer0_outputs(6039));
    outputs(7324) <= (layer0_outputs(6145)) xor (layer0_outputs(6194));
    outputs(7325) <= not(layer0_outputs(889));
    outputs(7326) <= not((layer0_outputs(2856)) or (layer0_outputs(4393)));
    outputs(7327) <= not((layer0_outputs(2268)) or (layer0_outputs(9259)));
    outputs(7328) <= (layer0_outputs(8735)) and not (layer0_outputs(4989));
    outputs(7329) <= layer0_outputs(9176);
    outputs(7330) <= not((layer0_outputs(9109)) xor (layer0_outputs(4340)));
    outputs(7331) <= layer0_outputs(8024);
    outputs(7332) <= (layer0_outputs(4489)) xor (layer0_outputs(8492));
    outputs(7333) <= not(layer0_outputs(7488));
    outputs(7334) <= not((layer0_outputs(1777)) or (layer0_outputs(9163)));
    outputs(7335) <= not(layer0_outputs(737)) or (layer0_outputs(6128));
    outputs(7336) <= not(layer0_outputs(4103));
    outputs(7337) <= (layer0_outputs(89)) and not (layer0_outputs(4203));
    outputs(7338) <= not(layer0_outputs(6992)) or (layer0_outputs(4106));
    outputs(7339) <= (layer0_outputs(6052)) and (layer0_outputs(5673));
    outputs(7340) <= (layer0_outputs(5367)) xor (layer0_outputs(8138));
    outputs(7341) <= (layer0_outputs(5249)) xor (layer0_outputs(7513));
    outputs(7342) <= (layer0_outputs(5429)) and (layer0_outputs(2903));
    outputs(7343) <= not((layer0_outputs(2631)) xor (layer0_outputs(5106)));
    outputs(7344) <= layer0_outputs(757);
    outputs(7345) <= layer0_outputs(1811);
    outputs(7346) <= layer0_outputs(189);
    outputs(7347) <= (layer0_outputs(592)) and not (layer0_outputs(2256));
    outputs(7348) <= layer0_outputs(8448);
    outputs(7349) <= (layer0_outputs(1884)) and not (layer0_outputs(6599));
    outputs(7350) <= not(layer0_outputs(8146));
    outputs(7351) <= not((layer0_outputs(3936)) xor (layer0_outputs(9563)));
    outputs(7352) <= layer0_outputs(9616);
    outputs(7353) <= (layer0_outputs(9890)) and not (layer0_outputs(8090));
    outputs(7354) <= (layer0_outputs(3052)) xor (layer0_outputs(2255));
    outputs(7355) <= not((layer0_outputs(9063)) or (layer0_outputs(1078)));
    outputs(7356) <= not((layer0_outputs(3020)) or (layer0_outputs(2221)));
    outputs(7357) <= (layer0_outputs(1842)) xor (layer0_outputs(2164));
    outputs(7358) <= not((layer0_outputs(340)) xor (layer0_outputs(1973)));
    outputs(7359) <= not((layer0_outputs(3006)) xor (layer0_outputs(2590)));
    outputs(7360) <= not(layer0_outputs(3813));
    outputs(7361) <= not((layer0_outputs(3775)) or (layer0_outputs(9269)));
    outputs(7362) <= (layer0_outputs(3306)) xor (layer0_outputs(3769));
    outputs(7363) <= layer0_outputs(9353);
    outputs(7364) <= layer0_outputs(759);
    outputs(7365) <= (layer0_outputs(8300)) xor (layer0_outputs(1051));
    outputs(7366) <= not((layer0_outputs(125)) xor (layer0_outputs(5043)));
    outputs(7367) <= (layer0_outputs(6213)) and not (layer0_outputs(8137));
    outputs(7368) <= not(layer0_outputs(9125));
    outputs(7369) <= not(layer0_outputs(3151)) or (layer0_outputs(6927));
    outputs(7370) <= not((layer0_outputs(8618)) xor (layer0_outputs(998)));
    outputs(7371) <= (layer0_outputs(7746)) and not (layer0_outputs(1980));
    outputs(7372) <= not(layer0_outputs(2926));
    outputs(7373) <= not(layer0_outputs(6314)) or (layer0_outputs(1422));
    outputs(7374) <= (layer0_outputs(8165)) xor (layer0_outputs(7457));
    outputs(7375) <= (layer0_outputs(979)) and not (layer0_outputs(5297));
    outputs(7376) <= (layer0_outputs(2337)) xor (layer0_outputs(7600));
    outputs(7377) <= (layer0_outputs(9367)) and not (layer0_outputs(6916));
    outputs(7378) <= (layer0_outputs(4507)) and (layer0_outputs(1679));
    outputs(7379) <= not((layer0_outputs(5570)) or (layer0_outputs(6280)));
    outputs(7380) <= not((layer0_outputs(4767)) xor (layer0_outputs(1429)));
    outputs(7381) <= not(layer0_outputs(6498));
    outputs(7382) <= layer0_outputs(3071);
    outputs(7383) <= (layer0_outputs(8689)) and not (layer0_outputs(7229));
    outputs(7384) <= layer0_outputs(9706);
    outputs(7385) <= (layer0_outputs(5502)) and not (layer0_outputs(6746));
    outputs(7386) <= not(layer0_outputs(7266)) or (layer0_outputs(10214));
    outputs(7387) <= not(layer0_outputs(6466));
    outputs(7388) <= not(layer0_outputs(2223));
    outputs(7389) <= (layer0_outputs(9845)) and (layer0_outputs(5383));
    outputs(7390) <= (layer0_outputs(7816)) xor (layer0_outputs(1689));
    outputs(7391) <= (layer0_outputs(2308)) xor (layer0_outputs(6701));
    outputs(7392) <= layer0_outputs(8422);
    outputs(7393) <= not(layer0_outputs(7916));
    outputs(7394) <= layer0_outputs(9379);
    outputs(7395) <= layer0_outputs(4495);
    outputs(7396) <= not((layer0_outputs(5860)) or (layer0_outputs(2710)));
    outputs(7397) <= not(layer0_outputs(5656)) or (layer0_outputs(6532));
    outputs(7398) <= not((layer0_outputs(5130)) xor (layer0_outputs(3439)));
    outputs(7399) <= (layer0_outputs(5574)) xor (layer0_outputs(6358));
    outputs(7400) <= not((layer0_outputs(10091)) xor (layer0_outputs(7128)));
    outputs(7401) <= layer0_outputs(5476);
    outputs(7402) <= not(layer0_outputs(9319));
    outputs(7403) <= not((layer0_outputs(7469)) or (layer0_outputs(5256)));
    outputs(7404) <= not(layer0_outputs(9124)) or (layer0_outputs(3828));
    outputs(7405) <= not(layer0_outputs(2357));
    outputs(7406) <= not(layer0_outputs(5481));
    outputs(7407) <= not(layer0_outputs(3226));
    outputs(7408) <= layer0_outputs(1458);
    outputs(7409) <= (layer0_outputs(6998)) xor (layer0_outputs(1177));
    outputs(7410) <= (layer0_outputs(8947)) and not (layer0_outputs(710));
    outputs(7411) <= not(layer0_outputs(3759));
    outputs(7412) <= not((layer0_outputs(1007)) xor (layer0_outputs(6935)));
    outputs(7413) <= layer0_outputs(931);
    outputs(7414) <= not((layer0_outputs(5538)) xor (layer0_outputs(7133)));
    outputs(7415) <= (layer0_outputs(8916)) and not (layer0_outputs(8895));
    outputs(7416) <= (layer0_outputs(3047)) and not (layer0_outputs(2826));
    outputs(7417) <= (layer0_outputs(1483)) xor (layer0_outputs(5102));
    outputs(7418) <= not(layer0_outputs(8909)) or (layer0_outputs(4839));
    outputs(7419) <= (layer0_outputs(1352)) xor (layer0_outputs(8353));
    outputs(7420) <= (layer0_outputs(9873)) and (layer0_outputs(6828));
    outputs(7421) <= layer0_outputs(6020);
    outputs(7422) <= layer0_outputs(1462);
    outputs(7423) <= not(layer0_outputs(1125)) or (layer0_outputs(7876));
    outputs(7424) <= (layer0_outputs(1895)) and not (layer0_outputs(4457));
    outputs(7425) <= not((layer0_outputs(4688)) xor (layer0_outputs(9651)));
    outputs(7426) <= (layer0_outputs(8733)) xor (layer0_outputs(126));
    outputs(7427) <= not((layer0_outputs(6854)) xor (layer0_outputs(120)));
    outputs(7428) <= '0';
    outputs(7429) <= layer0_outputs(8889);
    outputs(7430) <= not((layer0_outputs(8408)) or (layer0_outputs(6234)));
    outputs(7431) <= layer0_outputs(1706);
    outputs(7432) <= not((layer0_outputs(2937)) xor (layer0_outputs(8809)));
    outputs(7433) <= layer0_outputs(5617);
    outputs(7434) <= (layer0_outputs(7982)) and (layer0_outputs(6821));
    outputs(7435) <= not(layer0_outputs(8239));
    outputs(7436) <= not((layer0_outputs(9701)) xor (layer0_outputs(3385)));
    outputs(7437) <= not((layer0_outputs(5847)) xor (layer0_outputs(5673)));
    outputs(7438) <= not(layer0_outputs(2182));
    outputs(7439) <= layer0_outputs(528);
    outputs(7440) <= not(layer0_outputs(7942));
    outputs(7441) <= not((layer0_outputs(4213)) xor (layer0_outputs(6561)));
    outputs(7442) <= layer0_outputs(9722);
    outputs(7443) <= not((layer0_outputs(6)) or (layer0_outputs(2256)));
    outputs(7444) <= not(layer0_outputs(1564));
    outputs(7445) <= layer0_outputs(9405);
    outputs(7446) <= not((layer0_outputs(9097)) xor (layer0_outputs(478)));
    outputs(7447) <= not((layer0_outputs(9415)) or (layer0_outputs(9434)));
    outputs(7448) <= not((layer0_outputs(4970)) xor (layer0_outputs(8249)));
    outputs(7449) <= not((layer0_outputs(2997)) xor (layer0_outputs(3468)));
    outputs(7450) <= layer0_outputs(2308);
    outputs(7451) <= (layer0_outputs(511)) or (layer0_outputs(6229));
    outputs(7452) <= not(layer0_outputs(1871)) or (layer0_outputs(4017));
    outputs(7453) <= layer0_outputs(6492);
    outputs(7454) <= not(layer0_outputs(3241));
    outputs(7455) <= (layer0_outputs(1941)) and (layer0_outputs(701));
    outputs(7456) <= '0';
    outputs(7457) <= not(layer0_outputs(8503));
    outputs(7458) <= (layer0_outputs(4643)) and not (layer0_outputs(5532));
    outputs(7459) <= layer0_outputs(5455);
    outputs(7460) <= not(layer0_outputs(9261));
    outputs(7461) <= layer0_outputs(6366);
    outputs(7462) <= not(layer0_outputs(8978));
    outputs(7463) <= not(layer0_outputs(1871));
    outputs(7464) <= layer0_outputs(1852);
    outputs(7465) <= (layer0_outputs(5887)) and not (layer0_outputs(1414));
    outputs(7466) <= not((layer0_outputs(5622)) xor (layer0_outputs(619)));
    outputs(7467) <= (layer0_outputs(5796)) xor (layer0_outputs(5655));
    outputs(7468) <= not((layer0_outputs(2277)) or (layer0_outputs(5447)));
    outputs(7469) <= layer0_outputs(1039);
    outputs(7470) <= not(layer0_outputs(6894));
    outputs(7471) <= layer0_outputs(4046);
    outputs(7472) <= not(layer0_outputs(4841)) or (layer0_outputs(6973));
    outputs(7473) <= not(layer0_outputs(2709)) or (layer0_outputs(6977));
    outputs(7474) <= not(layer0_outputs(9986));
    outputs(7475) <= not((layer0_outputs(8445)) or (layer0_outputs(9629)));
    outputs(7476) <= not(layer0_outputs(426));
    outputs(7477) <= (layer0_outputs(4454)) and (layer0_outputs(873));
    outputs(7478) <= not((layer0_outputs(1124)) or (layer0_outputs(2462)));
    outputs(7479) <= (layer0_outputs(9795)) and not (layer0_outputs(4418));
    outputs(7480) <= (layer0_outputs(1040)) and (layer0_outputs(8055));
    outputs(7481) <= (layer0_outputs(6668)) xor (layer0_outputs(8504));
    outputs(7482) <= not((layer0_outputs(6218)) or (layer0_outputs(1624)));
    outputs(7483) <= not(layer0_outputs(6397));
    outputs(7484) <= not(layer0_outputs(5886));
    outputs(7485) <= layer0_outputs(2839);
    outputs(7486) <= layer0_outputs(7017);
    outputs(7487) <= (layer0_outputs(4721)) xor (layer0_outputs(9428));
    outputs(7488) <= not((layer0_outputs(5608)) xor (layer0_outputs(4794)));
    outputs(7489) <= (layer0_outputs(7353)) and not (layer0_outputs(1140));
    outputs(7490) <= layer0_outputs(4190);
    outputs(7491) <= layer0_outputs(7511);
    outputs(7492) <= layer0_outputs(5574);
    outputs(7493) <= (layer0_outputs(2756)) and not (layer0_outputs(377));
    outputs(7494) <= (layer0_outputs(8092)) xor (layer0_outputs(1803));
    outputs(7495) <= (layer0_outputs(5568)) xor (layer0_outputs(8429));
    outputs(7496) <= layer0_outputs(9117);
    outputs(7497) <= (layer0_outputs(4563)) and not (layer0_outputs(6517));
    outputs(7498) <= layer0_outputs(9904);
    outputs(7499) <= (layer0_outputs(7429)) or (layer0_outputs(9653));
    outputs(7500) <= (layer0_outputs(9363)) and (layer0_outputs(551));
    outputs(7501) <= not((layer0_outputs(113)) xor (layer0_outputs(4761)));
    outputs(7502) <= (layer0_outputs(1957)) and not (layer0_outputs(1797));
    outputs(7503) <= layer0_outputs(338);
    outputs(7504) <= layer0_outputs(1746);
    outputs(7505) <= (layer0_outputs(7620)) or (layer0_outputs(3356));
    outputs(7506) <= not((layer0_outputs(527)) xor (layer0_outputs(7156)));
    outputs(7507) <= not((layer0_outputs(3180)) or (layer0_outputs(4745)));
    outputs(7508) <= (layer0_outputs(4133)) and not (layer0_outputs(3671));
    outputs(7509) <= not(layer0_outputs(4768));
    outputs(7510) <= (layer0_outputs(1485)) and not (layer0_outputs(3242));
    outputs(7511) <= (layer0_outputs(3837)) xor (layer0_outputs(10235));
    outputs(7512) <= (layer0_outputs(4115)) and not (layer0_outputs(179));
    outputs(7513) <= not(layer0_outputs(8011)) or (layer0_outputs(4402));
    outputs(7514) <= layer0_outputs(1613);
    outputs(7515) <= (layer0_outputs(7061)) and (layer0_outputs(3221));
    outputs(7516) <= not(layer0_outputs(7520)) or (layer0_outputs(5977));
    outputs(7517) <= not((layer0_outputs(6975)) xor (layer0_outputs(2803)));
    outputs(7518) <= (layer0_outputs(3931)) and not (layer0_outputs(1602));
    outputs(7519) <= (layer0_outputs(785)) xor (layer0_outputs(8200));
    outputs(7520) <= not((layer0_outputs(7948)) xor (layer0_outputs(7169)));
    outputs(7521) <= not((layer0_outputs(9633)) or (layer0_outputs(9659)));
    outputs(7522) <= layer0_outputs(3479);
    outputs(7523) <= not((layer0_outputs(3339)) xor (layer0_outputs(2740)));
    outputs(7524) <= layer0_outputs(9838);
    outputs(7525) <= (layer0_outputs(6810)) xor (layer0_outputs(6383));
    outputs(7526) <= not(layer0_outputs(8122));
    outputs(7527) <= not((layer0_outputs(2116)) xor (layer0_outputs(7999)));
    outputs(7528) <= layer0_outputs(770);
    outputs(7529) <= layer0_outputs(4789);
    outputs(7530) <= not(layer0_outputs(801));
    outputs(7531) <= not((layer0_outputs(9063)) xor (layer0_outputs(8821)));
    outputs(7532) <= layer0_outputs(7689);
    outputs(7533) <= not((layer0_outputs(5990)) or (layer0_outputs(713)));
    outputs(7534) <= (layer0_outputs(7529)) and (layer0_outputs(3254));
    outputs(7535) <= (layer0_outputs(4508)) xor (layer0_outputs(7201));
    outputs(7536) <= not(layer0_outputs(1794));
    outputs(7537) <= (layer0_outputs(4723)) and not (layer0_outputs(10026));
    outputs(7538) <= (layer0_outputs(7653)) xor (layer0_outputs(8631));
    outputs(7539) <= not((layer0_outputs(6789)) xor (layer0_outputs(4271)));
    outputs(7540) <= layer0_outputs(9524);
    outputs(7541) <= not(layer0_outputs(1825)) or (layer0_outputs(178));
    outputs(7542) <= not(layer0_outputs(4797));
    outputs(7543) <= (layer0_outputs(3438)) and not (layer0_outputs(6779));
    outputs(7544) <= not(layer0_outputs(3296));
    outputs(7545) <= not(layer0_outputs(9683));
    outputs(7546) <= not(layer0_outputs(6706));
    outputs(7547) <= (layer0_outputs(4381)) xor (layer0_outputs(7736));
    outputs(7548) <= not(layer0_outputs(2947)) or (layer0_outputs(7899));
    outputs(7549) <= layer0_outputs(520);
    outputs(7550) <= (layer0_outputs(6812)) and not (layer0_outputs(581));
    outputs(7551) <= layer0_outputs(90);
    outputs(7552) <= layer0_outputs(990);
    outputs(7553) <= (layer0_outputs(523)) xor (layer0_outputs(6009));
    outputs(7554) <= layer0_outputs(1735);
    outputs(7555) <= not(layer0_outputs(2884));
    outputs(7556) <= layer0_outputs(9197);
    outputs(7557) <= not((layer0_outputs(6455)) xor (layer0_outputs(3260)));
    outputs(7558) <= not(layer0_outputs(10128));
    outputs(7559) <= not((layer0_outputs(9971)) or (layer0_outputs(9880)));
    outputs(7560) <= not(layer0_outputs(8347));
    outputs(7561) <= not(layer0_outputs(7104)) or (layer0_outputs(4124));
    outputs(7562) <= layer0_outputs(4615);
    outputs(7563) <= not((layer0_outputs(4433)) xor (layer0_outputs(1310)));
    outputs(7564) <= layer0_outputs(7258);
    outputs(7565) <= not(layer0_outputs(8793));
    outputs(7566) <= layer0_outputs(4675);
    outputs(7567) <= not(layer0_outputs(6533));
    outputs(7568) <= (layer0_outputs(6207)) or (layer0_outputs(4559));
    outputs(7569) <= (layer0_outputs(1084)) xor (layer0_outputs(10034));
    outputs(7570) <= not(layer0_outputs(9806));
    outputs(7571) <= not(layer0_outputs(7382));
    outputs(7572) <= not((layer0_outputs(2248)) or (layer0_outputs(7301)));
    outputs(7573) <= (layer0_outputs(4341)) and not (layer0_outputs(1262));
    outputs(7574) <= (layer0_outputs(3976)) and (layer0_outputs(9013));
    outputs(7575) <= layer0_outputs(2805);
    outputs(7576) <= layer0_outputs(1920);
    outputs(7577) <= not((layer0_outputs(2334)) xor (layer0_outputs(3672)));
    outputs(7578) <= (layer0_outputs(6091)) and not (layer0_outputs(2405));
    outputs(7579) <= (layer0_outputs(5702)) or (layer0_outputs(7510));
    outputs(7580) <= layer0_outputs(851);
    outputs(7581) <= layer0_outputs(5455);
    outputs(7582) <= (layer0_outputs(8782)) or (layer0_outputs(9401));
    outputs(7583) <= not(layer0_outputs(1163));
    outputs(7584) <= not((layer0_outputs(4173)) or (layer0_outputs(184)));
    outputs(7585) <= not((layer0_outputs(4699)) xor (layer0_outputs(3603)));
    outputs(7586) <= not((layer0_outputs(7431)) or (layer0_outputs(7328)));
    outputs(7587) <= not(layer0_outputs(1826));
    outputs(7588) <= layer0_outputs(8529);
    outputs(7589) <= not(layer0_outputs(8576));
    outputs(7590) <= layer0_outputs(1902);
    outputs(7591) <= layer0_outputs(1213);
    outputs(7592) <= not((layer0_outputs(7882)) xor (layer0_outputs(2450)));
    outputs(7593) <= not(layer0_outputs(5790));
    outputs(7594) <= (layer0_outputs(473)) xor (layer0_outputs(670));
    outputs(7595) <= (layer0_outputs(4863)) xor (layer0_outputs(1738));
    outputs(7596) <= not(layer0_outputs(9966)) or (layer0_outputs(4102));
    outputs(7597) <= not(layer0_outputs(791));
    outputs(7598) <= not(layer0_outputs(4776)) or (layer0_outputs(8371));
    outputs(7599) <= (layer0_outputs(2439)) and not (layer0_outputs(375));
    outputs(7600) <= (layer0_outputs(2023)) and not (layer0_outputs(10092));
    outputs(7601) <= layer0_outputs(2770);
    outputs(7602) <= (layer0_outputs(3745)) or (layer0_outputs(8992));
    outputs(7603) <= not((layer0_outputs(2130)) xor (layer0_outputs(9643)));
    outputs(7604) <= not((layer0_outputs(8533)) xor (layer0_outputs(504)));
    outputs(7605) <= (layer0_outputs(1856)) and not (layer0_outputs(459));
    outputs(7606) <= not((layer0_outputs(3922)) xor (layer0_outputs(5820)));
    outputs(7607) <= layer0_outputs(4612);
    outputs(7608) <= not(layer0_outputs(116));
    outputs(7609) <= not((layer0_outputs(7439)) xor (layer0_outputs(2695)));
    outputs(7610) <= (layer0_outputs(2863)) xor (layer0_outputs(8830));
    outputs(7611) <= layer0_outputs(8962);
    outputs(7612) <= not(layer0_outputs(5597));
    outputs(7613) <= not((layer0_outputs(2569)) or (layer0_outputs(2851)));
    outputs(7614) <= not(layer0_outputs(9936));
    outputs(7615) <= layer0_outputs(682);
    outputs(7616) <= (layer0_outputs(258)) xor (layer0_outputs(3909));
    outputs(7617) <= not((layer0_outputs(5641)) xor (layer0_outputs(5151)));
    outputs(7618) <= not(layer0_outputs(3899));
    outputs(7619) <= not(layer0_outputs(1917));
    outputs(7620) <= (layer0_outputs(3390)) xor (layer0_outputs(10101));
    outputs(7621) <= not(layer0_outputs(1818));
    outputs(7622) <= not(layer0_outputs(2272)) or (layer0_outputs(7937));
    outputs(7623) <= layer0_outputs(8489);
    outputs(7624) <= (layer0_outputs(4000)) and (layer0_outputs(10061));
    outputs(7625) <= not((layer0_outputs(7685)) and (layer0_outputs(4976)));
    outputs(7626) <= (layer0_outputs(7849)) and (layer0_outputs(4233));
    outputs(7627) <= (layer0_outputs(1401)) and (layer0_outputs(4070));
    outputs(7628) <= not((layer0_outputs(7048)) xor (layer0_outputs(7470)));
    outputs(7629) <= not(layer0_outputs(467));
    outputs(7630) <= not(layer0_outputs(7824));
    outputs(7631) <= layer0_outputs(7554);
    outputs(7632) <= not(layer0_outputs(4567)) or (layer0_outputs(8701));
    outputs(7633) <= layer0_outputs(6720);
    outputs(7634) <= (layer0_outputs(3054)) xor (layer0_outputs(3460));
    outputs(7635) <= not(layer0_outputs(3977)) or (layer0_outputs(4860));
    outputs(7636) <= not((layer0_outputs(4697)) and (layer0_outputs(8500)));
    outputs(7637) <= not(layer0_outputs(5599));
    outputs(7638) <= not(layer0_outputs(8170));
    outputs(7639) <= (layer0_outputs(9887)) and not (layer0_outputs(8193));
    outputs(7640) <= not(layer0_outputs(9398));
    outputs(7641) <= '0';
    outputs(7642) <= (layer0_outputs(5253)) xor (layer0_outputs(2930));
    outputs(7643) <= layer0_outputs(1023);
    outputs(7644) <= (layer0_outputs(1981)) and not (layer0_outputs(7202));
    outputs(7645) <= layer0_outputs(6563);
    outputs(7646) <= (layer0_outputs(1111)) xor (layer0_outputs(8289));
    outputs(7647) <= not((layer0_outputs(7541)) or (layer0_outputs(10181)));
    outputs(7648) <= layer0_outputs(8884);
    outputs(7649) <= (layer0_outputs(2309)) xor (layer0_outputs(3678));
    outputs(7650) <= layer0_outputs(3511);
    outputs(7651) <= not((layer0_outputs(6315)) xor (layer0_outputs(7033)));
    outputs(7652) <= (layer0_outputs(1334)) xor (layer0_outputs(3533));
    outputs(7653) <= not((layer0_outputs(176)) xor (layer0_outputs(6130)));
    outputs(7654) <= not(layer0_outputs(9775));
    outputs(7655) <= layer0_outputs(4844);
    outputs(7656) <= not(layer0_outputs(9284)) or (layer0_outputs(7537));
    outputs(7657) <= (layer0_outputs(935)) and not (layer0_outputs(4854));
    outputs(7658) <= not((layer0_outputs(289)) or (layer0_outputs(2066)));
    outputs(7659) <= not(layer0_outputs(6154));
    outputs(7660) <= (layer0_outputs(8152)) and (layer0_outputs(6304));
    outputs(7661) <= not(layer0_outputs(5563));
    outputs(7662) <= layer0_outputs(5960);
    outputs(7663) <= layer0_outputs(3738);
    outputs(7664) <= layer0_outputs(1267);
    outputs(7665) <= (layer0_outputs(4467)) and not (layer0_outputs(2736));
    outputs(7666) <= (layer0_outputs(2372)) or (layer0_outputs(5953));
    outputs(7667) <= not(layer0_outputs(2101));
    outputs(7668) <= (layer0_outputs(9557)) and (layer0_outputs(7965));
    outputs(7669) <= not(layer0_outputs(1546));
    outputs(7670) <= (layer0_outputs(2009)) and (layer0_outputs(9098));
    outputs(7671) <= layer0_outputs(2156);
    outputs(7672) <= not(layer0_outputs(5824));
    outputs(7673) <= layer0_outputs(722);
    outputs(7674) <= layer0_outputs(6505);
    outputs(7675) <= layer0_outputs(5453);
    outputs(7676) <= (layer0_outputs(1921)) xor (layer0_outputs(2586));
    outputs(7677) <= layer0_outputs(914);
    outputs(7678) <= (layer0_outputs(4793)) xor (layer0_outputs(6015));
    outputs(7679) <= not(layer0_outputs(9209)) or (layer0_outputs(9402));
    outputs(7680) <= layer0_outputs(3628);
    outputs(7681) <= not((layer0_outputs(1973)) and (layer0_outputs(216)));
    outputs(7682) <= not(layer0_outputs(3943));
    outputs(7683) <= layer0_outputs(2297);
    outputs(7684) <= (layer0_outputs(4973)) xor (layer0_outputs(506));
    outputs(7685) <= not(layer0_outputs(8425));
    outputs(7686) <= (layer0_outputs(836)) and not (layer0_outputs(1697));
    outputs(7687) <= (layer0_outputs(6572)) and not (layer0_outputs(2834));
    outputs(7688) <= (layer0_outputs(2119)) or (layer0_outputs(4928));
    outputs(7689) <= (layer0_outputs(2733)) and not (layer0_outputs(1500));
    outputs(7690) <= (layer0_outputs(760)) and not (layer0_outputs(3334));
    outputs(7691) <= layer0_outputs(7900);
    outputs(7692) <= not(layer0_outputs(4481));
    outputs(7693) <= layer0_outputs(3286);
    outputs(7694) <= not((layer0_outputs(2454)) xor (layer0_outputs(1903)));
    outputs(7695) <= not((layer0_outputs(8924)) and (layer0_outputs(1681)));
    outputs(7696) <= not(layer0_outputs(9362));
    outputs(7697) <= layer0_outputs(5523);
    outputs(7698) <= not((layer0_outputs(4394)) or (layer0_outputs(7869)));
    outputs(7699) <= not(layer0_outputs(8023));
    outputs(7700) <= (layer0_outputs(5155)) and not (layer0_outputs(8896));
    outputs(7701) <= (layer0_outputs(6874)) xor (layer0_outputs(3519));
    outputs(7702) <= layer0_outputs(1568);
    outputs(7703) <= (layer0_outputs(8225)) and (layer0_outputs(3442));
    outputs(7704) <= '0';
    outputs(7705) <= not(layer0_outputs(9717));
    outputs(7706) <= not(layer0_outputs(9152));
    outputs(7707) <= not(layer0_outputs(2369));
    outputs(7708) <= not((layer0_outputs(6)) or (layer0_outputs(669)));
    outputs(7709) <= '0';
    outputs(7710) <= not(layer0_outputs(4611));
    outputs(7711) <= (layer0_outputs(2879)) xor (layer0_outputs(3564));
    outputs(7712) <= (layer0_outputs(3547)) or (layer0_outputs(4902));
    outputs(7713) <= not((layer0_outputs(4238)) xor (layer0_outputs(7260)));
    outputs(7714) <= (layer0_outputs(6167)) and not (layer0_outputs(826));
    outputs(7715) <= not(layer0_outputs(8568)) or (layer0_outputs(9915));
    outputs(7716) <= not(layer0_outputs(555));
    outputs(7717) <= layer0_outputs(6480);
    outputs(7718) <= not(layer0_outputs(3625));
    outputs(7719) <= (layer0_outputs(127)) and not (layer0_outputs(7184));
    outputs(7720) <= layer0_outputs(4016);
    outputs(7721) <= layer0_outputs(7211);
    outputs(7722) <= (layer0_outputs(2376)) or (layer0_outputs(10031));
    outputs(7723) <= not(layer0_outputs(7303));
    outputs(7724) <= (layer0_outputs(4181)) and (layer0_outputs(2456));
    outputs(7725) <= layer0_outputs(442);
    outputs(7726) <= (layer0_outputs(4345)) xor (layer0_outputs(5064));
    outputs(7727) <= (layer0_outputs(1894)) and (layer0_outputs(9884));
    outputs(7728) <= (layer0_outputs(6174)) xor (layer0_outputs(3180));
    outputs(7729) <= layer0_outputs(649);
    outputs(7730) <= not(layer0_outputs(1633)) or (layer0_outputs(2376));
    outputs(7731) <= not(layer0_outputs(2876));
    outputs(7732) <= not(layer0_outputs(5139));
    outputs(7733) <= not(layer0_outputs(1045));
    outputs(7734) <= not((layer0_outputs(5425)) and (layer0_outputs(2936)));
    outputs(7735) <= not(layer0_outputs(3847)) or (layer0_outputs(3516));
    outputs(7736) <= layer0_outputs(1987);
    outputs(7737) <= not((layer0_outputs(3475)) or (layer0_outputs(7666)));
    outputs(7738) <= layer0_outputs(8853);
    outputs(7739) <= not(layer0_outputs(8836));
    outputs(7740) <= not((layer0_outputs(10150)) and (layer0_outputs(589)));
    outputs(7741) <= layer0_outputs(5418);
    outputs(7742) <= not((layer0_outputs(2012)) xor (layer0_outputs(9105)));
    outputs(7743) <= (layer0_outputs(1558)) xor (layer0_outputs(1878));
    outputs(7744) <= not((layer0_outputs(8518)) or (layer0_outputs(631)));
    outputs(7745) <= (layer0_outputs(1012)) xor (layer0_outputs(8286));
    outputs(7746) <= layer0_outputs(4716);
    outputs(7747) <= not((layer0_outputs(9664)) xor (layer0_outputs(864)));
    outputs(7748) <= (layer0_outputs(7915)) xor (layer0_outputs(808));
    outputs(7749) <= layer0_outputs(378);
    outputs(7750) <= (layer0_outputs(3860)) and not (layer0_outputs(8996));
    outputs(7751) <= not(layer0_outputs(1488));
    outputs(7752) <= not((layer0_outputs(4834)) or (layer0_outputs(4879)));
    outputs(7753) <= layer0_outputs(8770);
    outputs(7754) <= not(layer0_outputs(9763)) or (layer0_outputs(7709));
    outputs(7755) <= (layer0_outputs(5659)) and (layer0_outputs(6800));
    outputs(7756) <= (layer0_outputs(6596)) and not (layer0_outputs(4506));
    outputs(7757) <= (layer0_outputs(9699)) xor (layer0_outputs(7767));
    outputs(7758) <= not(layer0_outputs(6852));
    outputs(7759) <= not(layer0_outputs(9064)) or (layer0_outputs(8797));
    outputs(7760) <= not(layer0_outputs(5237));
    outputs(7761) <= not(layer0_outputs(5755)) or (layer0_outputs(3465));
    outputs(7762) <= (layer0_outputs(4627)) and not (layer0_outputs(2555));
    outputs(7763) <= (layer0_outputs(1567)) and not (layer0_outputs(9828));
    outputs(7764) <= not(layer0_outputs(4410));
    outputs(7765) <= not(layer0_outputs(1499));
    outputs(7766) <= (layer0_outputs(7853)) and not (layer0_outputs(3268));
    outputs(7767) <= (layer0_outputs(676)) and (layer0_outputs(5418));
    outputs(7768) <= layer0_outputs(3167);
    outputs(7769) <= layer0_outputs(9104);
    outputs(7770) <= layer0_outputs(12);
    outputs(7771) <= not(layer0_outputs(2181));
    outputs(7772) <= (layer0_outputs(2935)) and not (layer0_outputs(9279));
    outputs(7773) <= layer0_outputs(1703);
    outputs(7774) <= not((layer0_outputs(5326)) xor (layer0_outputs(8079)));
    outputs(7775) <= not((layer0_outputs(7328)) or (layer0_outputs(7387)));
    outputs(7776) <= not(layer0_outputs(2613));
    outputs(7777) <= not((layer0_outputs(9868)) xor (layer0_outputs(2948)));
    outputs(7778) <= not((layer0_outputs(2724)) xor (layer0_outputs(4222)));
    outputs(7779) <= not(layer0_outputs(4850));
    outputs(7780) <= (layer0_outputs(1679)) and not (layer0_outputs(1490));
    outputs(7781) <= layer0_outputs(1882);
    outputs(7782) <= (layer0_outputs(396)) and not (layer0_outputs(4959));
    outputs(7783) <= not((layer0_outputs(9482)) xor (layer0_outputs(9433)));
    outputs(7784) <= (layer0_outputs(7086)) and not (layer0_outputs(5075));
    outputs(7785) <= not((layer0_outputs(2681)) xor (layer0_outputs(6274)));
    outputs(7786) <= not(layer0_outputs(9480));
    outputs(7787) <= not(layer0_outputs(6802));
    outputs(7788) <= layer0_outputs(9450);
    outputs(7789) <= not(layer0_outputs(2749));
    outputs(7790) <= not((layer0_outputs(1109)) xor (layer0_outputs(9819)));
    outputs(7791) <= (layer0_outputs(7512)) and not (layer0_outputs(2078));
    outputs(7792) <= (layer0_outputs(9605)) and not (layer0_outputs(1730));
    outputs(7793) <= not(layer0_outputs(6622));
    outputs(7794) <= (layer0_outputs(8720)) and not (layer0_outputs(4396));
    outputs(7795) <= (layer0_outputs(2501)) xor (layer0_outputs(3719));
    outputs(7796) <= (layer0_outputs(597)) and not (layer0_outputs(2184));
    outputs(7797) <= not((layer0_outputs(3517)) xor (layer0_outputs(7782)));
    outputs(7798) <= (layer0_outputs(7246)) and not (layer0_outputs(6228));
    outputs(7799) <= (layer0_outputs(4274)) xor (layer0_outputs(5702));
    outputs(7800) <= not((layer0_outputs(8769)) xor (layer0_outputs(3764)));
    outputs(7801) <= (layer0_outputs(3654)) and not (layer0_outputs(10037));
    outputs(7802) <= layer0_outputs(8108);
    outputs(7803) <= (layer0_outputs(8219)) or (layer0_outputs(4));
    outputs(7804) <= not((layer0_outputs(892)) xor (layer0_outputs(3080)));
    outputs(7805) <= not(layer0_outputs(9121));
    outputs(7806) <= layer0_outputs(10227);
    outputs(7807) <= not((layer0_outputs(6135)) xor (layer0_outputs(4479)));
    outputs(7808) <= layer0_outputs(6318);
    outputs(7809) <= not((layer0_outputs(9977)) and (layer0_outputs(7796)));
    outputs(7810) <= (layer0_outputs(3673)) xor (layer0_outputs(91));
    outputs(7811) <= (layer0_outputs(471)) and (layer0_outputs(8786));
    outputs(7812) <= not(layer0_outputs(4154));
    outputs(7813) <= not((layer0_outputs(4062)) or (layer0_outputs(3780)));
    outputs(7814) <= not((layer0_outputs(544)) xor (layer0_outputs(5246)));
    outputs(7815) <= (layer0_outputs(903)) and (layer0_outputs(3783));
    outputs(7816) <= layer0_outputs(6578);
    outputs(7817) <= (layer0_outputs(5932)) xor (layer0_outputs(8392));
    outputs(7818) <= layer0_outputs(802);
    outputs(7819) <= (layer0_outputs(10018)) xor (layer0_outputs(10056));
    outputs(7820) <= not(layer0_outputs(6889));
    outputs(7821) <= layer0_outputs(4060);
    outputs(7822) <= not(layer0_outputs(1205)) or (layer0_outputs(969));
    outputs(7823) <= not((layer0_outputs(1009)) xor (layer0_outputs(6016)));
    outputs(7824) <= (layer0_outputs(7284)) and (layer0_outputs(10238));
    outputs(7825) <= not(layer0_outputs(9024));
    outputs(7826) <= layer0_outputs(5965);
    outputs(7827) <= (layer0_outputs(5996)) xor (layer0_outputs(4322));
    outputs(7828) <= (layer0_outputs(1584)) and not (layer0_outputs(797));
    outputs(7829) <= not(layer0_outputs(8718));
    outputs(7830) <= not((layer0_outputs(9313)) xor (layer0_outputs(2356)));
    outputs(7831) <= not(layer0_outputs(9317));
    outputs(7832) <= not((layer0_outputs(1929)) xor (layer0_outputs(8640)));
    outputs(7833) <= layer0_outputs(5053);
    outputs(7834) <= not((layer0_outputs(7362)) or (layer0_outputs(6591)));
    outputs(7835) <= (layer0_outputs(52)) xor (layer0_outputs(5868));
    outputs(7836) <= (layer0_outputs(5434)) xor (layer0_outputs(4319));
    outputs(7837) <= not(layer0_outputs(7575));
    outputs(7838) <= layer0_outputs(6108);
    outputs(7839) <= not(layer0_outputs(730));
    outputs(7840) <= not(layer0_outputs(6226)) or (layer0_outputs(8145));
    outputs(7841) <= not(layer0_outputs(8946));
    outputs(7842) <= layer0_outputs(8269);
    outputs(7843) <= layer0_outputs(4095);
    outputs(7844) <= (layer0_outputs(7480)) xor (layer0_outputs(3344));
    outputs(7845) <= (layer0_outputs(9382)) or (layer0_outputs(9357));
    outputs(7846) <= not(layer0_outputs(6708)) or (layer0_outputs(9655));
    outputs(7847) <= not((layer0_outputs(10211)) xor (layer0_outputs(6107)));
    outputs(7848) <= layer0_outputs(4031);
    outputs(7849) <= (layer0_outputs(896)) xor (layer0_outputs(6191));
    outputs(7850) <= (layer0_outputs(4465)) xor (layer0_outputs(7594));
    outputs(7851) <= (layer0_outputs(6243)) and (layer0_outputs(8898));
    outputs(7852) <= (layer0_outputs(4398)) and not (layer0_outputs(5131));
    outputs(7853) <= not((layer0_outputs(8454)) xor (layer0_outputs(8362)));
    outputs(7854) <= not((layer0_outputs(4943)) xor (layer0_outputs(7485)));
    outputs(7855) <= layer0_outputs(4505);
    outputs(7856) <= (layer0_outputs(6696)) and not (layer0_outputs(6789));
    outputs(7857) <= not((layer0_outputs(5933)) xor (layer0_outputs(4362)));
    outputs(7858) <= not(layer0_outputs(4186));
    outputs(7859) <= (layer0_outputs(8157)) and not (layer0_outputs(6033));
    outputs(7860) <= (layer0_outputs(9579)) and not (layer0_outputs(3981));
    outputs(7861) <= not((layer0_outputs(8048)) xor (layer0_outputs(3248)));
    outputs(7862) <= not(layer0_outputs(3191));
    outputs(7863) <= not(layer0_outputs(5427));
    outputs(7864) <= (layer0_outputs(5006)) and not (layer0_outputs(7035));
    outputs(7865) <= (layer0_outputs(6905)) and not (layer0_outputs(9214));
    outputs(7866) <= not((layer0_outputs(4276)) xor (layer0_outputs(8369)));
    outputs(7867) <= layer0_outputs(753);
    outputs(7868) <= not(layer0_outputs(2578)) or (layer0_outputs(7939));
    outputs(7869) <= not(layer0_outputs(10197));
    outputs(7870) <= (layer0_outputs(4517)) and not (layer0_outputs(3638));
    outputs(7871) <= not(layer0_outputs(3021)) or (layer0_outputs(1459));
    outputs(7872) <= not(layer0_outputs(1307));
    outputs(7873) <= (layer0_outputs(4130)) and (layer0_outputs(9315));
    outputs(7874) <= (layer0_outputs(5834)) and (layer0_outputs(4779));
    outputs(7875) <= not(layer0_outputs(6680)) or (layer0_outputs(5756));
    outputs(7876) <= not(layer0_outputs(6181));
    outputs(7877) <= (layer0_outputs(7459)) and (layer0_outputs(7015));
    outputs(7878) <= (layer0_outputs(6754)) and not (layer0_outputs(4551));
    outputs(7879) <= (layer0_outputs(5310)) and not (layer0_outputs(4430));
    outputs(7880) <= not(layer0_outputs(5269));
    outputs(7881) <= (layer0_outputs(7068)) and (layer0_outputs(8617));
    outputs(7882) <= not((layer0_outputs(8007)) or (layer0_outputs(8863)));
    outputs(7883) <= layer0_outputs(10119);
    outputs(7884) <= (layer0_outputs(5594)) xor (layer0_outputs(7038));
    outputs(7885) <= layer0_outputs(5954);
    outputs(7886) <= layer0_outputs(7905);
    outputs(7887) <= '1';
    outputs(7888) <= layer0_outputs(7363);
    outputs(7889) <= not((layer0_outputs(4366)) or (layer0_outputs(9737)));
    outputs(7890) <= layer0_outputs(2005);
    outputs(7891) <= layer0_outputs(2837);
    outputs(7892) <= layer0_outputs(10001);
    outputs(7893) <= not(layer0_outputs(1774));
    outputs(7894) <= (layer0_outputs(8217)) xor (layer0_outputs(4631));
    outputs(7895) <= not(layer0_outputs(8561));
    outputs(7896) <= not((layer0_outputs(5373)) xor (layer0_outputs(10071)));
    outputs(7897) <= (layer0_outputs(5663)) or (layer0_outputs(1687));
    outputs(7898) <= layer0_outputs(8913);
    outputs(7899) <= not(layer0_outputs(6482));
    outputs(7900) <= layer0_outputs(9859);
    outputs(7901) <= (layer0_outputs(5328)) xor (layer0_outputs(633));
    outputs(7902) <= not((layer0_outputs(7859)) xor (layer0_outputs(7918)));
    outputs(7903) <= (layer0_outputs(9444)) and not (layer0_outputs(1896));
    outputs(7904) <= (layer0_outputs(7438)) xor (layer0_outputs(394));
    outputs(7905) <= not((layer0_outputs(9371)) xor (layer0_outputs(291)));
    outputs(7906) <= not((layer0_outputs(7953)) xor (layer0_outputs(3995)));
    outputs(7907) <= not(layer0_outputs(4171));
    outputs(7908) <= not(layer0_outputs(9020));
    outputs(7909) <= not((layer0_outputs(9451)) xor (layer0_outputs(3273)));
    outputs(7910) <= (layer0_outputs(2500)) xor (layer0_outputs(7527));
    outputs(7911) <= (layer0_outputs(5293)) and (layer0_outputs(3672));
    outputs(7912) <= (layer0_outputs(3059)) and (layer0_outputs(7535));
    outputs(7913) <= layer0_outputs(134);
    outputs(7914) <= (layer0_outputs(9366)) and not (layer0_outputs(9134));
    outputs(7915) <= layer0_outputs(2193);
    outputs(7916) <= (layer0_outputs(47)) or (layer0_outputs(641));
    outputs(7917) <= layer0_outputs(8606);
    outputs(7918) <= not((layer0_outputs(9811)) xor (layer0_outputs(2428)));
    outputs(7919) <= (layer0_outputs(746)) xor (layer0_outputs(411));
    outputs(7920) <= (layer0_outputs(957)) and not (layer0_outputs(1875));
    outputs(7921) <= layer0_outputs(9142);
    outputs(7922) <= (layer0_outputs(1940)) and (layer0_outputs(4760));
    outputs(7923) <= not(layer0_outputs(8652));
    outputs(7924) <= layer0_outputs(8340);
    outputs(7925) <= layer0_outputs(5976);
    outputs(7926) <= not(layer0_outputs(9781)) or (layer0_outputs(2407));
    outputs(7927) <= (layer0_outputs(5801)) or (layer0_outputs(6184));
    outputs(7928) <= not(layer0_outputs(9166));
    outputs(7929) <= not(layer0_outputs(8908));
    outputs(7930) <= layer0_outputs(8062);
    outputs(7931) <= (layer0_outputs(9712)) xor (layer0_outputs(3541));
    outputs(7932) <= (layer0_outputs(9645)) and (layer0_outputs(488));
    outputs(7933) <= not((layer0_outputs(1451)) xor (layer0_outputs(2873)));
    outputs(7934) <= layer0_outputs(1433);
    outputs(7935) <= (layer0_outputs(3998)) and not (layer0_outputs(10084));
    outputs(7936) <= not((layer0_outputs(7463)) xor (layer0_outputs(912)));
    outputs(7937) <= (layer0_outputs(6988)) xor (layer0_outputs(8026));
    outputs(7938) <= layer0_outputs(7259);
    outputs(7939) <= (layer0_outputs(9754)) and (layer0_outputs(7155));
    outputs(7940) <= not((layer0_outputs(9761)) or (layer0_outputs(6498)));
    outputs(7941) <= not(layer0_outputs(8472));
    outputs(7942) <= layer0_outputs(7296);
    outputs(7943) <= not((layer0_outputs(4900)) or (layer0_outputs(4105)));
    outputs(7944) <= layer0_outputs(6744);
    outputs(7945) <= layer0_outputs(9542);
    outputs(7946) <= (layer0_outputs(8560)) and (layer0_outputs(9968));
    outputs(7947) <= not((layer0_outputs(2069)) and (layer0_outputs(6258)));
    outputs(7948) <= layer0_outputs(3168);
    outputs(7949) <= layer0_outputs(432);
    outputs(7950) <= layer0_outputs(1732);
    outputs(7951) <= not(layer0_outputs(1999));
    outputs(7952) <= not(layer0_outputs(1609)) or (layer0_outputs(6291));
    outputs(7953) <= (layer0_outputs(5934)) xor (layer0_outputs(238));
    outputs(7954) <= (layer0_outputs(6576)) xor (layer0_outputs(3325));
    outputs(7955) <= not(layer0_outputs(4176));
    outputs(7956) <= layer0_outputs(7699);
    outputs(7957) <= not((layer0_outputs(6734)) xor (layer0_outputs(6699)));
    outputs(7958) <= not(layer0_outputs(3933));
    outputs(7959) <= (layer0_outputs(6486)) and not (layer0_outputs(4116));
    outputs(7960) <= (layer0_outputs(4280)) xor (layer0_outputs(4570));
    outputs(7961) <= (layer0_outputs(7071)) xor (layer0_outputs(4471));
    outputs(7962) <= (layer0_outputs(8250)) or (layer0_outputs(1225));
    outputs(7963) <= not((layer0_outputs(3938)) and (layer0_outputs(688)));
    outputs(7964) <= not(layer0_outputs(7629));
    outputs(7965) <= (layer0_outputs(6677)) and not (layer0_outputs(4138));
    outputs(7966) <= not(layer0_outputs(8049));
    outputs(7967) <= (layer0_outputs(6076)) or (layer0_outputs(4255));
    outputs(7968) <= layer0_outputs(10075);
    outputs(7969) <= not(layer0_outputs(2315));
    outputs(7970) <= not(layer0_outputs(5969));
    outputs(7971) <= not(layer0_outputs(2696));
    outputs(7972) <= not(layer0_outputs(2175));
    outputs(7973) <= (layer0_outputs(469)) xor (layer0_outputs(8110));
    outputs(7974) <= layer0_outputs(832);
    outputs(7975) <= not((layer0_outputs(6643)) xor (layer0_outputs(21)));
    outputs(7976) <= (layer0_outputs(8962)) and (layer0_outputs(10048));
    outputs(7977) <= layer0_outputs(2307);
    outputs(7978) <= not(layer0_outputs(5587));
    outputs(7979) <= (layer0_outputs(7544)) and not (layer0_outputs(554));
    outputs(7980) <= (layer0_outputs(9361)) and (layer0_outputs(1101));
    outputs(7981) <= layer0_outputs(6827);
    outputs(7982) <= not((layer0_outputs(5793)) xor (layer0_outputs(9008)));
    outputs(7983) <= not(layer0_outputs(5760));
    outputs(7984) <= (layer0_outputs(8272)) xor (layer0_outputs(4889));
    outputs(7985) <= not(layer0_outputs(1300));
    outputs(7986) <= (layer0_outputs(5148)) and not (layer0_outputs(9113));
    outputs(7987) <= (layer0_outputs(4296)) and not (layer0_outputs(6055));
    outputs(7988) <= (layer0_outputs(6808)) and not (layer0_outputs(5319));
    outputs(7989) <= not((layer0_outputs(1322)) or (layer0_outputs(6963)));
    outputs(7990) <= not((layer0_outputs(10046)) and (layer0_outputs(9459)));
    outputs(7991) <= not(layer0_outputs(9788));
    outputs(7992) <= not(layer0_outputs(6621));
    outputs(7993) <= (layer0_outputs(8632)) and not (layer0_outputs(9089));
    outputs(7994) <= (layer0_outputs(5296)) and not (layer0_outputs(5201));
    outputs(7995) <= (layer0_outputs(6404)) and (layer0_outputs(1480));
    outputs(7996) <= (layer0_outputs(2984)) and not (layer0_outputs(8956));
    outputs(7997) <= not((layer0_outputs(5592)) xor (layer0_outputs(4575)));
    outputs(7998) <= not((layer0_outputs(4166)) xor (layer0_outputs(414)));
    outputs(7999) <= (layer0_outputs(3187)) and not (layer0_outputs(4116));
    outputs(8000) <= (layer0_outputs(232)) xor (layer0_outputs(9669));
    outputs(8001) <= not((layer0_outputs(5077)) xor (layer0_outputs(7807)));
    outputs(8002) <= not(layer0_outputs(5353));
    outputs(8003) <= layer0_outputs(1245);
    outputs(8004) <= (layer0_outputs(8874)) and not (layer0_outputs(159));
    outputs(8005) <= not((layer0_outputs(3205)) or (layer0_outputs(125)));
    outputs(8006) <= not((layer0_outputs(4162)) xor (layer0_outputs(1495)));
    outputs(8007) <= not(layer0_outputs(7726));
    outputs(8008) <= not((layer0_outputs(4552)) xor (layer0_outputs(3521)));
    outputs(8009) <= (layer0_outputs(3947)) and not (layer0_outputs(217));
    outputs(8010) <= not((layer0_outputs(7840)) or (layer0_outputs(7843)));
    outputs(8011) <= (layer0_outputs(2097)) and not (layer0_outputs(2317));
    outputs(8012) <= not((layer0_outputs(4049)) xor (layer0_outputs(1207)));
    outputs(8013) <= (layer0_outputs(7890)) xor (layer0_outputs(7638));
    outputs(8014) <= (layer0_outputs(6877)) xor (layer0_outputs(5966));
    outputs(8015) <= layer0_outputs(9706);
    outputs(8016) <= not(layer0_outputs(3193));
    outputs(8017) <= layer0_outputs(8729);
    outputs(8018) <= not(layer0_outputs(611));
    outputs(8019) <= not(layer0_outputs(3362));
    outputs(8020) <= not(layer0_outputs(5988)) or (layer0_outputs(3942));
    outputs(8021) <= (layer0_outputs(3281)) and (layer0_outputs(1000));
    outputs(8022) <= (layer0_outputs(5350)) and not (layer0_outputs(7381));
    outputs(8023) <= (layer0_outputs(3029)) and not (layer0_outputs(4021));
    outputs(8024) <= not(layer0_outputs(8432));
    outputs(8025) <= not(layer0_outputs(7692));
    outputs(8026) <= not((layer0_outputs(9880)) or (layer0_outputs(1848)));
    outputs(8027) <= layer0_outputs(2167);
    outputs(8028) <= not((layer0_outputs(4634)) xor (layer0_outputs(2993)));
    outputs(8029) <= not(layer0_outputs(4029));
    outputs(8030) <= not(layer0_outputs(7021));
    outputs(8031) <= not((layer0_outputs(6309)) xor (layer0_outputs(6939)));
    outputs(8032) <= not((layer0_outputs(2208)) xor (layer0_outputs(400)));
    outputs(8033) <= (layer0_outputs(8145)) or (layer0_outputs(9342));
    outputs(8034) <= not((layer0_outputs(7136)) xor (layer0_outputs(1291)));
    outputs(8035) <= not((layer0_outputs(7372)) xor (layer0_outputs(8056)));
    outputs(8036) <= (layer0_outputs(7304)) xor (layer0_outputs(1928));
    outputs(8037) <= layer0_outputs(553);
    outputs(8038) <= not(layer0_outputs(2545));
    outputs(8039) <= (layer0_outputs(6376)) and not (layer0_outputs(2481));
    outputs(8040) <= not(layer0_outputs(1855));
    outputs(8041) <= layer0_outputs(10165);
    outputs(8042) <= not(layer0_outputs(7142));
    outputs(8043) <= layer0_outputs(1552);
    outputs(8044) <= not((layer0_outputs(8291)) xor (layer0_outputs(5868)));
    outputs(8045) <= not(layer0_outputs(8836));
    outputs(8046) <= not(layer0_outputs(6801)) or (layer0_outputs(2114));
    outputs(8047) <= not(layer0_outputs(4709));
    outputs(8048) <= not(layer0_outputs(4226));
    outputs(8049) <= layer0_outputs(543);
    outputs(8050) <= not(layer0_outputs(3502));
    outputs(8051) <= not((layer0_outputs(9760)) xor (layer0_outputs(3319)));
    outputs(8052) <= not((layer0_outputs(5242)) xor (layer0_outputs(5021)));
    outputs(8053) <= (layer0_outputs(5329)) xor (layer0_outputs(3018));
    outputs(8054) <= not(layer0_outputs(2939));
    outputs(8055) <= layer0_outputs(996);
    outputs(8056) <= (layer0_outputs(8726)) xor (layer0_outputs(2947));
    outputs(8057) <= (layer0_outputs(735)) xor (layer0_outputs(1444));
    outputs(8058) <= not(layer0_outputs(6175));
    outputs(8059) <= not(layer0_outputs(1477));
    outputs(8060) <= not(layer0_outputs(9693));
    outputs(8061) <= (layer0_outputs(7115)) xor (layer0_outputs(1269));
    outputs(8062) <= not(layer0_outputs(3124));
    outputs(8063) <= layer0_outputs(8666);
    outputs(8064) <= layer0_outputs(5915);
    outputs(8065) <= layer0_outputs(4543);
    outputs(8066) <= not(layer0_outputs(5148)) or (layer0_outputs(390));
    outputs(8067) <= (layer0_outputs(6356)) xor (layer0_outputs(6272));
    outputs(8068) <= not((layer0_outputs(9645)) xor (layer0_outputs(5568)));
    outputs(8069) <= not((layer0_outputs(8239)) xor (layer0_outputs(1737)));
    outputs(8070) <= layer0_outputs(303);
    outputs(8071) <= not((layer0_outputs(1491)) xor (layer0_outputs(3961)));
    outputs(8072) <= layer0_outputs(5535);
    outputs(8073) <= not((layer0_outputs(409)) xor (layer0_outputs(5747)));
    outputs(8074) <= not(layer0_outputs(4932));
    outputs(8075) <= (layer0_outputs(3107)) xor (layer0_outputs(8513));
    outputs(8076) <= (layer0_outputs(6273)) and not (layer0_outputs(4697));
    outputs(8077) <= (layer0_outputs(9635)) xor (layer0_outputs(3960));
    outputs(8078) <= layer0_outputs(1286);
    outputs(8079) <= not(layer0_outputs(6799));
    outputs(8080) <= (layer0_outputs(5939)) or (layer0_outputs(2513));
    outputs(8081) <= (layer0_outputs(2211)) xor (layer0_outputs(1204));
    outputs(8082) <= not(layer0_outputs(2299));
    outputs(8083) <= (layer0_outputs(7034)) or (layer0_outputs(5892));
    outputs(8084) <= layer0_outputs(3048);
    outputs(8085) <= not(layer0_outputs(327));
    outputs(8086) <= not(layer0_outputs(4056));
    outputs(8087) <= not(layer0_outputs(8846)) or (layer0_outputs(5439));
    outputs(8088) <= layer0_outputs(6313);
    outputs(8089) <= (layer0_outputs(948)) xor (layer0_outputs(2484));
    outputs(8090) <= layer0_outputs(9671);
    outputs(8091) <= not(layer0_outputs(2994));
    outputs(8092) <= not((layer0_outputs(136)) xor (layer0_outputs(5805)));
    outputs(8093) <= (layer0_outputs(9530)) and (layer0_outputs(8216));
    outputs(8094) <= layer0_outputs(3889);
    outputs(8095) <= (layer0_outputs(206)) and not (layer0_outputs(2659));
    outputs(8096) <= (layer0_outputs(7938)) xor (layer0_outputs(2671));
    outputs(8097) <= layer0_outputs(1547);
    outputs(8098) <= not(layer0_outputs(3194));
    outputs(8099) <= (layer0_outputs(1553)) xor (layer0_outputs(9118));
    outputs(8100) <= not((layer0_outputs(7072)) or (layer0_outputs(5016)));
    outputs(8101) <= layer0_outputs(8156);
    outputs(8102) <= not((layer0_outputs(4220)) xor (layer0_outputs(5883)));
    outputs(8103) <= not(layer0_outputs(1465));
    outputs(8104) <= not((layer0_outputs(4408)) xor (layer0_outputs(3288)));
    outputs(8105) <= not(layer0_outputs(2181));
    outputs(8106) <= layer0_outputs(9168);
    outputs(8107) <= not((layer0_outputs(3381)) xor (layer0_outputs(7880)));
    outputs(8108) <= layer0_outputs(1705);
    outputs(8109) <= layer0_outputs(10077);
    outputs(8110) <= layer0_outputs(2791);
    outputs(8111) <= not(layer0_outputs(4558)) or (layer0_outputs(3338));
    outputs(8112) <= not((layer0_outputs(6328)) xor (layer0_outputs(960)));
    outputs(8113) <= (layer0_outputs(4547)) xor (layer0_outputs(4531));
    outputs(8114) <= (layer0_outputs(6451)) and (layer0_outputs(2232));
    outputs(8115) <= layer0_outputs(2009);
    outputs(8116) <= (layer0_outputs(638)) and (layer0_outputs(4922));
    outputs(8117) <= layer0_outputs(1552);
    outputs(8118) <= not(layer0_outputs(774)) or (layer0_outputs(6556));
    outputs(8119) <= not(layer0_outputs(2598));
    outputs(8120) <= not(layer0_outputs(4247));
    outputs(8121) <= (layer0_outputs(1823)) or (layer0_outputs(9817));
    outputs(8122) <= not((layer0_outputs(271)) or (layer0_outputs(3710)));
    outputs(8123) <= not(layer0_outputs(9167));
    outputs(8124) <= (layer0_outputs(8939)) xor (layer0_outputs(7138));
    outputs(8125) <= not(layer0_outputs(333)) or (layer0_outputs(1419));
    outputs(8126) <= (layer0_outputs(10213)) xor (layer0_outputs(853));
    outputs(8127) <= (layer0_outputs(4006)) xor (layer0_outputs(9293));
    outputs(8128) <= layer0_outputs(3353);
    outputs(8129) <= (layer0_outputs(4188)) and not (layer0_outputs(6747));
    outputs(8130) <= not(layer0_outputs(3327));
    outputs(8131) <= not(layer0_outputs(3446));
    outputs(8132) <= not((layer0_outputs(7951)) xor (layer0_outputs(1109)));
    outputs(8133) <= layer0_outputs(9009);
    outputs(8134) <= (layer0_outputs(6004)) and not (layer0_outputs(2165));
    outputs(8135) <= layer0_outputs(9403);
    outputs(8136) <= layer0_outputs(7236);
    outputs(8137) <= not((layer0_outputs(7442)) xor (layer0_outputs(1426)));
    outputs(8138) <= (layer0_outputs(5704)) and not (layer0_outputs(4203));
    outputs(8139) <= (layer0_outputs(8598)) and (layer0_outputs(5866));
    outputs(8140) <= (layer0_outputs(5704)) xor (layer0_outputs(3078));
    outputs(8141) <= not(layer0_outputs(9199)) or (layer0_outputs(4473));
    outputs(8142) <= layer0_outputs(5752);
    outputs(8143) <= not(layer0_outputs(5621));
    outputs(8144) <= not((layer0_outputs(9790)) xor (layer0_outputs(4441)));
    outputs(8145) <= (layer0_outputs(6831)) and (layer0_outputs(4705));
    outputs(8146) <= not((layer0_outputs(5596)) xor (layer0_outputs(8817)));
    outputs(8147) <= not((layer0_outputs(1288)) xor (layer0_outputs(8018)));
    outputs(8148) <= not((layer0_outputs(1438)) or (layer0_outputs(6252)));
    outputs(8149) <= (layer0_outputs(6197)) or (layer0_outputs(1405));
    outputs(8150) <= not((layer0_outputs(9175)) xor (layer0_outputs(9672)));
    outputs(8151) <= layer0_outputs(7299);
    outputs(8152) <= not((layer0_outputs(3323)) xor (layer0_outputs(4435)));
    outputs(8153) <= (layer0_outputs(9843)) and (layer0_outputs(473));
    outputs(8154) <= (layer0_outputs(3305)) xor (layer0_outputs(5997));
    outputs(8155) <= layer0_outputs(6623);
    outputs(8156) <= not(layer0_outputs(1635));
    outputs(8157) <= not(layer0_outputs(6185)) or (layer0_outputs(5875));
    outputs(8158) <= (layer0_outputs(220)) and not (layer0_outputs(7802));
    outputs(8159) <= not(layer0_outputs(4713));
    outputs(8160) <= not((layer0_outputs(8651)) or (layer0_outputs(8958)));
    outputs(8161) <= (layer0_outputs(7976)) or (layer0_outputs(4150));
    outputs(8162) <= layer0_outputs(8211);
    outputs(8163) <= not(layer0_outputs(3972));
    outputs(8164) <= (layer0_outputs(8198)) xor (layer0_outputs(809));
    outputs(8165) <= (layer0_outputs(6974)) xor (layer0_outputs(9560));
    outputs(8166) <= not(layer0_outputs(8418));
    outputs(8167) <= not(layer0_outputs(1516));
    outputs(8168) <= (layer0_outputs(6168)) and not (layer0_outputs(8726));
    outputs(8169) <= layer0_outputs(4332);
    outputs(8170) <= not(layer0_outputs(963));
    outputs(8171) <= not(layer0_outputs(7713));
    outputs(8172) <= not((layer0_outputs(8333)) xor (layer0_outputs(10229)));
    outputs(8173) <= not(layer0_outputs(2004));
    outputs(8174) <= not(layer0_outputs(8206));
    outputs(8175) <= not(layer0_outputs(4194)) or (layer0_outputs(6365));
    outputs(8176) <= layer0_outputs(4844);
    outputs(8177) <= (layer0_outputs(7178)) and not (layer0_outputs(275));
    outputs(8178) <= (layer0_outputs(6787)) xor (layer0_outputs(10001));
    outputs(8179) <= (layer0_outputs(5078)) xor (layer0_outputs(4878));
    outputs(8180) <= (layer0_outputs(8727)) xor (layer0_outputs(740));
    outputs(8181) <= not((layer0_outputs(6874)) xor (layer0_outputs(1225)));
    outputs(8182) <= layer0_outputs(9061);
    outputs(8183) <= layer0_outputs(6425);
    outputs(8184) <= (layer0_outputs(2061)) xor (layer0_outputs(7728));
    outputs(8185) <= (layer0_outputs(353)) xor (layer0_outputs(2095));
    outputs(8186) <= not((layer0_outputs(7268)) xor (layer0_outputs(7586)));
    outputs(8187) <= not(layer0_outputs(2548));
    outputs(8188) <= not(layer0_outputs(5927));
    outputs(8189) <= not(layer0_outputs(1775)) or (layer0_outputs(4017));
    outputs(8190) <= (layer0_outputs(1651)) and not (layer0_outputs(6002));
    outputs(8191) <= layer0_outputs(8447);
    outputs(8192) <= (layer0_outputs(6146)) and (layer0_outputs(6345));
    outputs(8193) <= not(layer0_outputs(454));
    outputs(8194) <= not(layer0_outputs(4272));
    outputs(8195) <= not((layer0_outputs(8632)) xor (layer0_outputs(3267)));
    outputs(8196) <= not(layer0_outputs(1835));
    outputs(8197) <= not((layer0_outputs(1901)) xor (layer0_outputs(5536)));
    outputs(8198) <= not(layer0_outputs(6201)) or (layer0_outputs(152));
    outputs(8199) <= (layer0_outputs(934)) xor (layer0_outputs(9609));
    outputs(8200) <= (layer0_outputs(4682)) xor (layer0_outputs(4012));
    outputs(8201) <= (layer0_outputs(2783)) xor (layer0_outputs(8443));
    outputs(8202) <= (layer0_outputs(2142)) and not (layer0_outputs(5437));
    outputs(8203) <= not(layer0_outputs(4598)) or (layer0_outputs(6673));
    outputs(8204) <= (layer0_outputs(5313)) or (layer0_outputs(5233));
    outputs(8205) <= (layer0_outputs(5223)) or (layer0_outputs(1833));
    outputs(8206) <= (layer0_outputs(10087)) xor (layer0_outputs(5013));
    outputs(8207) <= not((layer0_outputs(974)) and (layer0_outputs(4216)));
    outputs(8208) <= layer0_outputs(7364);
    outputs(8209) <= (layer0_outputs(5216)) xor (layer0_outputs(7158));
    outputs(8210) <= not(layer0_outputs(315)) or (layer0_outputs(1470));
    outputs(8211) <= not((layer0_outputs(7864)) and (layer0_outputs(4444)));
    outputs(8212) <= (layer0_outputs(8482)) xor (layer0_outputs(828));
    outputs(8213) <= not(layer0_outputs(3045));
    outputs(8214) <= not((layer0_outputs(715)) and (layer0_outputs(3683)));
    outputs(8215) <= not((layer0_outputs(86)) xor (layer0_outputs(3541)));
    outputs(8216) <= not((layer0_outputs(7534)) and (layer0_outputs(9864)));
    outputs(8217) <= not((layer0_outputs(5786)) xor (layer0_outputs(7139)));
    outputs(8218) <= layer0_outputs(1165);
    outputs(8219) <= not((layer0_outputs(1470)) and (layer0_outputs(5686)));
    outputs(8220) <= not(layer0_outputs(77));
    outputs(8221) <= (layer0_outputs(7089)) and not (layer0_outputs(4957));
    outputs(8222) <= not(layer0_outputs(1113)) or (layer0_outputs(9918));
    outputs(8223) <= not((layer0_outputs(3993)) xor (layer0_outputs(8961)));
    outputs(8224) <= (layer0_outputs(5613)) xor (layer0_outputs(9562));
    outputs(8225) <= not(layer0_outputs(5025));
    outputs(8226) <= (layer0_outputs(6529)) xor (layer0_outputs(9084));
    outputs(8227) <= not(layer0_outputs(8088));
    outputs(8228) <= not((layer0_outputs(10143)) or (layer0_outputs(3503)));
    outputs(8229) <= not(layer0_outputs(10151)) or (layer0_outputs(8481));
    outputs(8230) <= not(layer0_outputs(4657)) or (layer0_outputs(7731));
    outputs(8231) <= not(layer0_outputs(5518));
    outputs(8232) <= not((layer0_outputs(3494)) xor (layer0_outputs(4405)));
    outputs(8233) <= not(layer0_outputs(1625)) or (layer0_outputs(3073));
    outputs(8234) <= '0';
    outputs(8235) <= not((layer0_outputs(9467)) xor (layer0_outputs(1780)));
    outputs(8236) <= (layer0_outputs(5192)) and not (layer0_outputs(5525));
    outputs(8237) <= not((layer0_outputs(2874)) xor (layer0_outputs(1388)));
    outputs(8238) <= not((layer0_outputs(8366)) or (layer0_outputs(2692)));
    outputs(8239) <= not((layer0_outputs(3247)) or (layer0_outputs(5254)));
    outputs(8240) <= layer0_outputs(3505);
    outputs(8241) <= layer0_outputs(5676);
    outputs(8242) <= layer0_outputs(4538);
    outputs(8243) <= layer0_outputs(3848);
    outputs(8244) <= not((layer0_outputs(4662)) xor (layer0_outputs(4958)));
    outputs(8245) <= (layer0_outputs(10134)) xor (layer0_outputs(10008));
    outputs(8246) <= not((layer0_outputs(8235)) xor (layer0_outputs(5110)));
    outputs(8247) <= layer0_outputs(6703);
    outputs(8248) <= not((layer0_outputs(10223)) xor (layer0_outputs(6606)));
    outputs(8249) <= not(layer0_outputs(4550));
    outputs(8250) <= (layer0_outputs(9931)) and (layer0_outputs(6077));
    outputs(8251) <= not(layer0_outputs(6750));
    outputs(8252) <= layer0_outputs(7360);
    outputs(8253) <= layer0_outputs(58);
    outputs(8254) <= layer0_outputs(9062);
    outputs(8255) <= (layer0_outputs(7486)) xor (layer0_outputs(6428));
    outputs(8256) <= (layer0_outputs(507)) and (layer0_outputs(9573));
    outputs(8257) <= not((layer0_outputs(7025)) and (layer0_outputs(2316)));
    outputs(8258) <= not((layer0_outputs(9508)) xor (layer0_outputs(5215)));
    outputs(8259) <= not((layer0_outputs(5030)) xor (layer0_outputs(9345)));
    outputs(8260) <= layer0_outputs(5481);
    outputs(8261) <= layer0_outputs(1415);
    outputs(8262) <= not((layer0_outputs(9247)) xor (layer0_outputs(9100)));
    outputs(8263) <= (layer0_outputs(6072)) and not (layer0_outputs(10092));
    outputs(8264) <= '1';
    outputs(8265) <= (layer0_outputs(5510)) xor (layer0_outputs(3914));
    outputs(8266) <= not(layer0_outputs(2777)) or (layer0_outputs(4610));
    outputs(8267) <= (layer0_outputs(230)) xor (layer0_outputs(4751));
    outputs(8268) <= (layer0_outputs(9720)) and not (layer0_outputs(5305));
    outputs(8269) <= not((layer0_outputs(3968)) and (layer0_outputs(2943)));
    outputs(8270) <= not(layer0_outputs(9094)) or (layer0_outputs(5330));
    outputs(8271) <= layer0_outputs(3915);
    outputs(8272) <= not(layer0_outputs(1263));
    outputs(8273) <= not(layer0_outputs(2191));
    outputs(8274) <= not(layer0_outputs(10206));
    outputs(8275) <= not((layer0_outputs(7602)) xor (layer0_outputs(5675)));
    outputs(8276) <= not(layer0_outputs(3758));
    outputs(8277) <= (layer0_outputs(8121)) xor (layer0_outputs(3642));
    outputs(8278) <= layer0_outputs(4982);
    outputs(8279) <= (layer0_outputs(9123)) or (layer0_outputs(1208));
    outputs(8280) <= layer0_outputs(3880);
    outputs(8281) <= (layer0_outputs(8952)) xor (layer0_outputs(8132));
    outputs(8282) <= not(layer0_outputs(360));
    outputs(8283) <= (layer0_outputs(10069)) or (layer0_outputs(8462));
    outputs(8284) <= (layer0_outputs(2072)) or (layer0_outputs(6933));
    outputs(8285) <= not((layer0_outputs(3145)) and (layer0_outputs(3283)));
    outputs(8286) <= not((layer0_outputs(5317)) xor (layer0_outputs(1051)));
    outputs(8287) <= not(layer0_outputs(4280));
    outputs(8288) <= layer0_outputs(6879);
    outputs(8289) <= not((layer0_outputs(5604)) or (layer0_outputs(590)));
    outputs(8290) <= not(layer0_outputs(6056));
    outputs(8291) <= not((layer0_outputs(510)) xor (layer0_outputs(689)));
    outputs(8292) <= '1';
    outputs(8293) <= (layer0_outputs(9992)) xor (layer0_outputs(3226));
    outputs(8294) <= not(layer0_outputs(7433));
    outputs(8295) <= layer0_outputs(5708);
    outputs(8296) <= not((layer0_outputs(2432)) or (layer0_outputs(3223)));
    outputs(8297) <= not(layer0_outputs(4754));
    outputs(8298) <= (layer0_outputs(6670)) or (layer0_outputs(119));
    outputs(8299) <= not(layer0_outputs(6292));
    outputs(8300) <= (layer0_outputs(7632)) or (layer0_outputs(5821));
    outputs(8301) <= layer0_outputs(3490);
    outputs(8302) <= layer0_outputs(719);
    outputs(8303) <= layer0_outputs(3860);
    outputs(8304) <= (layer0_outputs(6298)) xor (layer0_outputs(2946));
    outputs(8305) <= layer0_outputs(1560);
    outputs(8306) <= (layer0_outputs(3116)) xor (layer0_outputs(1352));
    outputs(8307) <= not(layer0_outputs(9686));
    outputs(8308) <= not((layer0_outputs(2323)) xor (layer0_outputs(317)));
    outputs(8309) <= not((layer0_outputs(3066)) and (layer0_outputs(6992)));
    outputs(8310) <= (layer0_outputs(5348)) or (layer0_outputs(4605));
    outputs(8311) <= layer0_outputs(10189);
    outputs(8312) <= not(layer0_outputs(526));
    outputs(8313) <= (layer0_outputs(987)) and not (layer0_outputs(1764));
    outputs(8314) <= not(layer0_outputs(8177));
    outputs(8315) <= (layer0_outputs(178)) xor (layer0_outputs(3332));
    outputs(8316) <= not((layer0_outputs(1532)) and (layer0_outputs(1753)));
    outputs(8317) <= layer0_outputs(6120);
    outputs(8318) <= layer0_outputs(9451);
    outputs(8319) <= (layer0_outputs(245)) and (layer0_outputs(5789));
    outputs(8320) <= not(layer0_outputs(9231));
    outputs(8321) <= not(layer0_outputs(6525)) or (layer0_outputs(10127));
    outputs(8322) <= not(layer0_outputs(4825));
    outputs(8323) <= not(layer0_outputs(5934));
    outputs(8324) <= (layer0_outputs(502)) xor (layer0_outputs(4597));
    outputs(8325) <= not(layer0_outputs(8153));
    outputs(8326) <= not(layer0_outputs(1108));
    outputs(8327) <= (layer0_outputs(955)) or (layer0_outputs(3054));
    outputs(8328) <= layer0_outputs(6762);
    outputs(8329) <= (layer0_outputs(1565)) and not (layer0_outputs(3956));
    outputs(8330) <= (layer0_outputs(3238)) and not (layer0_outputs(8932));
    outputs(8331) <= not(layer0_outputs(2452)) or (layer0_outputs(1541));
    outputs(8332) <= not(layer0_outputs(4518));
    outputs(8333) <= not((layer0_outputs(7850)) xor (layer0_outputs(2661)));
    outputs(8334) <= (layer0_outputs(4058)) xor (layer0_outputs(9914));
    outputs(8335) <= not((layer0_outputs(8956)) xor (layer0_outputs(3033)));
    outputs(8336) <= not((layer0_outputs(8479)) xor (layer0_outputs(3552)));
    outputs(8337) <= layer0_outputs(2329);
    outputs(8338) <= layer0_outputs(5019);
    outputs(8339) <= (layer0_outputs(7427)) and (layer0_outputs(7357));
    outputs(8340) <= not((layer0_outputs(10002)) xor (layer0_outputs(7369)));
    outputs(8341) <= not((layer0_outputs(9302)) xor (layer0_outputs(3248)));
    outputs(8342) <= not((layer0_outputs(5419)) xor (layer0_outputs(7302)));
    outputs(8343) <= not(layer0_outputs(8731));
    outputs(8344) <= (layer0_outputs(4307)) or (layer0_outputs(428));
    outputs(8345) <= not(layer0_outputs(562));
    outputs(8346) <= not((layer0_outputs(10196)) or (layer0_outputs(4436)));
    outputs(8347) <= not((layer0_outputs(4755)) xor (layer0_outputs(1446)));
    outputs(8348) <= layer0_outputs(9375);
    outputs(8349) <= not(layer0_outputs(7561));
    outputs(8350) <= not((layer0_outputs(6462)) or (layer0_outputs(1240)));
    outputs(8351) <= not(layer0_outputs(8891)) or (layer0_outputs(2818));
    outputs(8352) <= not((layer0_outputs(5101)) xor (layer0_outputs(2579)));
    outputs(8353) <= (layer0_outputs(3791)) xor (layer0_outputs(7304));
    outputs(8354) <= (layer0_outputs(2216)) xor (layer0_outputs(2885));
    outputs(8355) <= not(layer0_outputs(3401));
    outputs(8356) <= (layer0_outputs(1118)) or (layer0_outputs(2821));
    outputs(8357) <= layer0_outputs(7558);
    outputs(8358) <= not((layer0_outputs(243)) xor (layer0_outputs(5500)));
    outputs(8359) <= layer0_outputs(9586);
    outputs(8360) <= (layer0_outputs(576)) and (layer0_outputs(3983));
    outputs(8361) <= (layer0_outputs(2758)) and not (layer0_outputs(5901));
    outputs(8362) <= layer0_outputs(5788);
    outputs(8363) <= (layer0_outputs(9312)) xor (layer0_outputs(3364));
    outputs(8364) <= not((layer0_outputs(5770)) and (layer0_outputs(5525)));
    outputs(8365) <= not((layer0_outputs(8396)) or (layer0_outputs(748)));
    outputs(8366) <= not((layer0_outputs(6048)) or (layer0_outputs(1016)));
    outputs(8367) <= layer0_outputs(4912);
    outputs(8368) <= not(layer0_outputs(10202));
    outputs(8369) <= layer0_outputs(4370);
    outputs(8370) <= layer0_outputs(9509);
    outputs(8371) <= layer0_outputs(6035);
    outputs(8372) <= not((layer0_outputs(3295)) or (layer0_outputs(3905)));
    outputs(8373) <= layer0_outputs(8708);
    outputs(8374) <= not(layer0_outputs(3771));
    outputs(8375) <= not((layer0_outputs(2302)) xor (layer0_outputs(4331)));
    outputs(8376) <= not(layer0_outputs(8757));
    outputs(8377) <= (layer0_outputs(1742)) and not (layer0_outputs(937));
    outputs(8378) <= (layer0_outputs(2648)) and not (layer0_outputs(2960));
    outputs(8379) <= layer0_outputs(8580);
    outputs(8380) <= not(layer0_outputs(10230));
    outputs(8381) <= (layer0_outputs(1189)) or (layer0_outputs(2408));
    outputs(8382) <= not(layer0_outputs(4438));
    outputs(8383) <= not(layer0_outputs(8468));
    outputs(8384) <= layer0_outputs(3933);
    outputs(8385) <= not((layer0_outputs(2424)) or (layer0_outputs(1469)));
    outputs(8386) <= not(layer0_outputs(1535)) or (layer0_outputs(6912));
    outputs(8387) <= not((layer0_outputs(2278)) or (layer0_outputs(806)));
    outputs(8388) <= layer0_outputs(7284);
    outputs(8389) <= not((layer0_outputs(9241)) xor (layer0_outputs(6073)));
    outputs(8390) <= not((layer0_outputs(9514)) xor (layer0_outputs(4959)));
    outputs(8391) <= not(layer0_outputs(9031));
    outputs(8392) <= layer0_outputs(5459);
    outputs(8393) <= not(layer0_outputs(2126));
    outputs(8394) <= not((layer0_outputs(8376)) xor (layer0_outputs(9856)));
    outputs(8395) <= (layer0_outputs(8841)) and not (layer0_outputs(1831));
    outputs(8396) <= not(layer0_outputs(2280));
    outputs(8397) <= (layer0_outputs(10175)) xor (layer0_outputs(2775));
    outputs(8398) <= not((layer0_outputs(223)) xor (layer0_outputs(4771)));
    outputs(8399) <= not((layer0_outputs(4466)) xor (layer0_outputs(1999)));
    outputs(8400) <= not(layer0_outputs(2619));
    outputs(8401) <= not(layer0_outputs(9191));
    outputs(8402) <= not(layer0_outputs(5283)) or (layer0_outputs(4826));
    outputs(8403) <= not(layer0_outputs(6712));
    outputs(8404) <= not((layer0_outputs(5351)) xor (layer0_outputs(1576)));
    outputs(8405) <= (layer0_outputs(9146)) or (layer0_outputs(5677));
    outputs(8406) <= layer0_outputs(1090);
    outputs(8407) <= (layer0_outputs(4291)) xor (layer0_outputs(8450));
    outputs(8408) <= (layer0_outputs(648)) xor (layer0_outputs(2321));
    outputs(8409) <= (layer0_outputs(2324)) xor (layer0_outputs(7610));
    outputs(8410) <= (layer0_outputs(1793)) xor (layer0_outputs(1697));
    outputs(8411) <= not(layer0_outputs(9853));
    outputs(8412) <= not(layer0_outputs(8414));
    outputs(8413) <= not((layer0_outputs(6300)) xor (layer0_outputs(1290)));
    outputs(8414) <= not(layer0_outputs(2632));
    outputs(8415) <= not((layer0_outputs(920)) xor (layer0_outputs(6277)));
    outputs(8416) <= layer0_outputs(4535);
    outputs(8417) <= not(layer0_outputs(1639)) or (layer0_outputs(9004));
    outputs(8418) <= layer0_outputs(9162);
    outputs(8419) <= (layer0_outputs(9477)) xor (layer0_outputs(75));
    outputs(8420) <= not(layer0_outputs(7827));
    outputs(8421) <= not(layer0_outputs(197)) or (layer0_outputs(7465));
    outputs(8422) <= not(layer0_outputs(2024));
    outputs(8423) <= (layer0_outputs(8064)) and not (layer0_outputs(8633));
    outputs(8424) <= layer0_outputs(5321);
    outputs(8425) <= (layer0_outputs(10138)) and not (layer0_outputs(6385));
    outputs(8426) <= not((layer0_outputs(1191)) and (layer0_outputs(9195)));
    outputs(8427) <= (layer0_outputs(7816)) and not (layer0_outputs(6313));
    outputs(8428) <= (layer0_outputs(5715)) xor (layer0_outputs(2491));
    outputs(8429) <= layer0_outputs(4498);
    outputs(8430) <= not(layer0_outputs(2912));
    outputs(8431) <= layer0_outputs(9363);
    outputs(8432) <= (layer0_outputs(798)) xor (layer0_outputs(911));
    outputs(8433) <= (layer0_outputs(6783)) xor (layer0_outputs(642));
    outputs(8434) <= not(layer0_outputs(4550));
    outputs(8435) <= layer0_outputs(7837);
    outputs(8436) <= layer0_outputs(9709);
    outputs(8437) <= layer0_outputs(9772);
    outputs(8438) <= (layer0_outputs(53)) or (layer0_outputs(3636));
    outputs(8439) <= layer0_outputs(9785);
    outputs(8440) <= (layer0_outputs(7636)) xor (layer0_outputs(569));
    outputs(8441) <= not((layer0_outputs(6693)) and (layer0_outputs(3842)));
    outputs(8442) <= (layer0_outputs(204)) and (layer0_outputs(5499));
    outputs(8443) <= (layer0_outputs(851)) and not (layer0_outputs(7784));
    outputs(8444) <= (layer0_outputs(9114)) xor (layer0_outputs(7205));
    outputs(8445) <= not(layer0_outputs(591));
    outputs(8446) <= not(layer0_outputs(2999));
    outputs(8447) <= (layer0_outputs(7593)) and not (layer0_outputs(7546));
    outputs(8448) <= (layer0_outputs(311)) or (layer0_outputs(5192));
    outputs(8449) <= not(layer0_outputs(9687)) or (layer0_outputs(5071));
    outputs(8450) <= not(layer0_outputs(9972));
    outputs(8451) <= not(layer0_outputs(2841));
    outputs(8452) <= (layer0_outputs(2509)) xor (layer0_outputs(751));
    outputs(8453) <= not(layer0_outputs(223)) or (layer0_outputs(7376));
    outputs(8454) <= '1';
    outputs(8455) <= not(layer0_outputs(8234));
    outputs(8456) <= not(layer0_outputs(6084));
    outputs(8457) <= (layer0_outputs(4981)) and not (layer0_outputs(4970));
    outputs(8458) <= layer0_outputs(8412);
    outputs(8459) <= not((layer0_outputs(6996)) and (layer0_outputs(4095)));
    outputs(8460) <= (layer0_outputs(6884)) xor (layer0_outputs(7234));
    outputs(8461) <= layer0_outputs(6617);
    outputs(8462) <= not(layer0_outputs(9061));
    outputs(8463) <= (layer0_outputs(71)) and not (layer0_outputs(2313));
    outputs(8464) <= not(layer0_outputs(6751));
    outputs(8465) <= (layer0_outputs(9727)) and (layer0_outputs(8252));
    outputs(8466) <= not(layer0_outputs(5781)) or (layer0_outputs(5837));
    outputs(8467) <= (layer0_outputs(1959)) or (layer0_outputs(8767));
    outputs(8468) <= not((layer0_outputs(1888)) or (layer0_outputs(4629)));
    outputs(8469) <= not(layer0_outputs(3411)) or (layer0_outputs(7436));
    outputs(8470) <= (layer0_outputs(3978)) xor (layer0_outputs(5953));
    outputs(8471) <= not(layer0_outputs(2842)) or (layer0_outputs(8626));
    outputs(8472) <= not((layer0_outputs(5066)) or (layer0_outputs(9093)));
    outputs(8473) <= not((layer0_outputs(933)) or (layer0_outputs(5522)));
    outputs(8474) <= layer0_outputs(9804);
    outputs(8475) <= (layer0_outputs(811)) xor (layer0_outputs(3417));
    outputs(8476) <= layer0_outputs(2329);
    outputs(8477) <= not(layer0_outputs(8973));
    outputs(8478) <= (layer0_outputs(3944)) and not (layer0_outputs(5555));
    outputs(8479) <= not(layer0_outputs(3973)) or (layer0_outputs(2738));
    outputs(8480) <= (layer0_outputs(9367)) and (layer0_outputs(7112));
    outputs(8481) <= not((layer0_outputs(2434)) or (layer0_outputs(38)));
    outputs(8482) <= (layer0_outputs(9151)) xor (layer0_outputs(8150));
    outputs(8483) <= not((layer0_outputs(9812)) xor (layer0_outputs(4364)));
    outputs(8484) <= layer0_outputs(6522);
    outputs(8485) <= not(layer0_outputs(4869));
    outputs(8486) <= (layer0_outputs(8292)) xor (layer0_outputs(3220));
    outputs(8487) <= layer0_outputs(7536);
    outputs(8488) <= not(layer0_outputs(1942)) or (layer0_outputs(6018));
    outputs(8489) <= layer0_outputs(6242);
    outputs(8490) <= layer0_outputs(767);
    outputs(8491) <= not(layer0_outputs(7879));
    outputs(8492) <= not((layer0_outputs(4540)) xor (layer0_outputs(5172)));
    outputs(8493) <= layer0_outputs(9321);
    outputs(8494) <= (layer0_outputs(8001)) and (layer0_outputs(2405));
    outputs(8495) <= layer0_outputs(827);
    outputs(8496) <= not((layer0_outputs(625)) xor (layer0_outputs(2731)));
    outputs(8497) <= not((layer0_outputs(1241)) or (layer0_outputs(348)));
    outputs(8498) <= not(layer0_outputs(9522));
    outputs(8499) <= not(layer0_outputs(2864));
    outputs(8500) <= '1';
    outputs(8501) <= layer0_outputs(10172);
    outputs(8502) <= layer0_outputs(799);
    outputs(8503) <= not((layer0_outputs(4632)) xor (layer0_outputs(253)));
    outputs(8504) <= (layer0_outputs(5318)) xor (layer0_outputs(7455));
    outputs(8505) <= (layer0_outputs(8592)) and not (layer0_outputs(6454));
    outputs(8506) <= not(layer0_outputs(8897));
    outputs(8507) <= not((layer0_outputs(9455)) and (layer0_outputs(9492)));
    outputs(8508) <= (layer0_outputs(6984)) xor (layer0_outputs(5099));
    outputs(8509) <= (layer0_outputs(423)) xor (layer0_outputs(8997));
    outputs(8510) <= (layer0_outputs(2318)) xor (layer0_outputs(6618));
    outputs(8511) <= (layer0_outputs(4164)) and (layer0_outputs(7785));
    outputs(8512) <= (layer0_outputs(4635)) xor (layer0_outputs(8918));
    outputs(8513) <= not(layer0_outputs(4037));
    outputs(8514) <= (layer0_outputs(6391)) xor (layer0_outputs(4137));
    outputs(8515) <= not((layer0_outputs(6100)) xor (layer0_outputs(2087)));
    outputs(8516) <= layer0_outputs(4432);
    outputs(8517) <= (layer0_outputs(4035)) xor (layer0_outputs(8135));
    outputs(8518) <= not((layer0_outputs(341)) xor (layer0_outputs(4140)));
    outputs(8519) <= (layer0_outputs(6872)) or (layer0_outputs(6743));
    outputs(8520) <= (layer0_outputs(8623)) and not (layer0_outputs(6463));
    outputs(8521) <= not((layer0_outputs(7723)) xor (layer0_outputs(6389)));
    outputs(8522) <= (layer0_outputs(5264)) xor (layer0_outputs(5856));
    outputs(8523) <= not((layer0_outputs(8637)) xor (layer0_outputs(9526)));
    outputs(8524) <= (layer0_outputs(9288)) xor (layer0_outputs(147));
    outputs(8525) <= not((layer0_outputs(9353)) or (layer0_outputs(5140)));
    outputs(8526) <= not(layer0_outputs(6425));
    outputs(8527) <= layer0_outputs(4965);
    outputs(8528) <= not(layer0_outputs(8739));
    outputs(8529) <= layer0_outputs(9032);
    outputs(8530) <= not(layer0_outputs(758)) or (layer0_outputs(5363));
    outputs(8531) <= not(layer0_outputs(2578));
    outputs(8532) <= not(layer0_outputs(2746));
    outputs(8533) <= not(layer0_outputs(4764));
    outputs(8534) <= not(layer0_outputs(1505)) or (layer0_outputs(2049));
    outputs(8535) <= not(layer0_outputs(1394)) or (layer0_outputs(3978));
    outputs(8536) <= not(layer0_outputs(4831));
    outputs(8537) <= not(layer0_outputs(5402));
    outputs(8538) <= not((layer0_outputs(2091)) xor (layer0_outputs(5183)));
    outputs(8539) <= not((layer0_outputs(8832)) xor (layer0_outputs(5652)));
    outputs(8540) <= not((layer0_outputs(10012)) and (layer0_outputs(7249)));
    outputs(8541) <= layer0_outputs(264);
    outputs(8542) <= not((layer0_outputs(9120)) xor (layer0_outputs(2820)));
    outputs(8543) <= not(layer0_outputs(2694)) or (layer0_outputs(62));
    outputs(8544) <= (layer0_outputs(8999)) xor (layer0_outputs(7456));
    outputs(8545) <= (layer0_outputs(5712)) xor (layer0_outputs(3137));
    outputs(8546) <= not(layer0_outputs(9199)) or (layer0_outputs(7116));
    outputs(8547) <= not(layer0_outputs(8484));
    outputs(8548) <= (layer0_outputs(6144)) xor (layer0_outputs(940));
    outputs(8549) <= (layer0_outputs(1818)) xor (layer0_outputs(6325));
    outputs(8550) <= not(layer0_outputs(1658));
    outputs(8551) <= (layer0_outputs(7888)) xor (layer0_outputs(7865));
    outputs(8552) <= not((layer0_outputs(4302)) xor (layer0_outputs(5247)));
    outputs(8553) <= not(layer0_outputs(4352)) or (layer0_outputs(10043));
    outputs(8554) <= (layer0_outputs(7551)) xor (layer0_outputs(6635));
    outputs(8555) <= not(layer0_outputs(2264));
    outputs(8556) <= '1';
    outputs(8557) <= not((layer0_outputs(8665)) xor (layer0_outputs(10028)));
    outputs(8558) <= (layer0_outputs(5090)) and not (layer0_outputs(4408));
    outputs(8559) <= not(layer0_outputs(6003));
    outputs(8560) <= not((layer0_outputs(9447)) xor (layer0_outputs(9253)));
    outputs(8561) <= (layer0_outputs(5118)) xor (layer0_outputs(10106));
    outputs(8562) <= not(layer0_outputs(4637));
    outputs(8563) <= (layer0_outputs(1193)) xor (layer0_outputs(4698));
    outputs(8564) <= (layer0_outputs(1950)) or (layer0_outputs(266));
    outputs(8565) <= layer0_outputs(4985);
    outputs(8566) <= not(layer0_outputs(3657)) or (layer0_outputs(9782));
    outputs(8567) <= not(layer0_outputs(2604)) or (layer0_outputs(64));
    outputs(8568) <= not((layer0_outputs(1116)) xor (layer0_outputs(6563)));
    outputs(8569) <= (layer0_outputs(6241)) and (layer0_outputs(7590));
    outputs(8570) <= (layer0_outputs(3009)) xor (layer0_outputs(7877));
    outputs(8571) <= not(layer0_outputs(9607)) or (layer0_outputs(655));
    outputs(8572) <= (layer0_outputs(4265)) and not (layer0_outputs(4991));
    outputs(8573) <= (layer0_outputs(5234)) xor (layer0_outputs(7182));
    outputs(8574) <= layer0_outputs(6656);
    outputs(8575) <= (layer0_outputs(4225)) or (layer0_outputs(1559));
    outputs(8576) <= not(layer0_outputs(3160)) or (layer0_outputs(8130));
    outputs(8577) <= (layer0_outputs(3560)) xor (layer0_outputs(5519));
    outputs(8578) <= layer0_outputs(10190);
    outputs(8579) <= layer0_outputs(4593);
    outputs(8580) <= layer0_outputs(8747);
    outputs(8581) <= layer0_outputs(5315);
    outputs(8582) <= not((layer0_outputs(2952)) and (layer0_outputs(9412)));
    outputs(8583) <= layer0_outputs(8539);
    outputs(8584) <= layer0_outputs(9901);
    outputs(8585) <= layer0_outputs(9774);
    outputs(8586) <= (layer0_outputs(5042)) xor (layer0_outputs(6043));
    outputs(8587) <= (layer0_outputs(2039)) xor (layer0_outputs(8497));
    outputs(8588) <= not(layer0_outputs(7571));
    outputs(8589) <= layer0_outputs(2909);
    outputs(8590) <= not(layer0_outputs(895));
    outputs(8591) <= not(layer0_outputs(2312)) or (layer0_outputs(8743));
    outputs(8592) <= not((layer0_outputs(7765)) or (layer0_outputs(771)));
    outputs(8593) <= not((layer0_outputs(2573)) xor (layer0_outputs(6059)));
    outputs(8594) <= (layer0_outputs(8805)) and not (layer0_outputs(3975));
    outputs(8595) <= not((layer0_outputs(8446)) xor (layer0_outputs(1869)));
    outputs(8596) <= not((layer0_outputs(5228)) xor (layer0_outputs(9005)));
    outputs(8597) <= not((layer0_outputs(2130)) xor (layer0_outputs(776)));
    outputs(8598) <= (layer0_outputs(1260)) and (layer0_outputs(1937));
    outputs(8599) <= (layer0_outputs(358)) xor (layer0_outputs(6202));
    outputs(8600) <= (layer0_outputs(7694)) xor (layer0_outputs(5038));
    outputs(8601) <= not(layer0_outputs(6069));
    outputs(8602) <= (layer0_outputs(6926)) and (layer0_outputs(3009));
    outputs(8603) <= not((layer0_outputs(9513)) xor (layer0_outputs(1819)));
    outputs(8604) <= layer0_outputs(9952);
    outputs(8605) <= (layer0_outputs(1325)) and not (layer0_outputs(6403));
    outputs(8606) <= (layer0_outputs(6958)) and (layer0_outputs(2783));
    outputs(8607) <= not(layer0_outputs(194));
    outputs(8608) <= not((layer0_outputs(3015)) and (layer0_outputs(6566)));
    outputs(8609) <= not((layer0_outputs(5964)) xor (layer0_outputs(2969)));
    outputs(8610) <= not(layer0_outputs(5817)) or (layer0_outputs(7411));
    outputs(8611) <= not(layer0_outputs(2307)) or (layer0_outputs(5819));
    outputs(8612) <= (layer0_outputs(4204)) xor (layer0_outputs(1368));
    outputs(8613) <= not((layer0_outputs(328)) or (layer0_outputs(9947)));
    outputs(8614) <= not((layer0_outputs(7505)) and (layer0_outputs(6424)));
    outputs(8615) <= not(layer0_outputs(2363)) or (layer0_outputs(5788));
    outputs(8616) <= not((layer0_outputs(525)) xor (layer0_outputs(7829)));
    outputs(8617) <= layer0_outputs(586);
    outputs(8618) <= not(layer0_outputs(9515));
    outputs(8619) <= not((layer0_outputs(509)) xor (layer0_outputs(5776)));
    outputs(8620) <= not(layer0_outputs(7076));
    outputs(8621) <= not((layer0_outputs(270)) xor (layer0_outputs(7834)));
    outputs(8622) <= (layer0_outputs(7890)) or (layer0_outputs(6331));
    outputs(8623) <= not((layer0_outputs(6712)) or (layer0_outputs(1447)));
    outputs(8624) <= layer0_outputs(2906);
    outputs(8625) <= not(layer0_outputs(8705));
    outputs(8626) <= not((layer0_outputs(8232)) xor (layer0_outputs(4307)));
    outputs(8627) <= not(layer0_outputs(7863));
    outputs(8628) <= not(layer0_outputs(7626));
    outputs(8629) <= (layer0_outputs(3549)) and not (layer0_outputs(3626));
    outputs(8630) <= (layer0_outputs(7893)) xor (layer0_outputs(3075));
    outputs(8631) <= (layer0_outputs(3738)) or (layer0_outputs(942));
    outputs(8632) <= (layer0_outputs(1936)) xor (layer0_outputs(3568));
    outputs(8633) <= not(layer0_outputs(123)) or (layer0_outputs(1997));
    outputs(8634) <= not(layer0_outputs(6888));
    outputs(8635) <= layer0_outputs(720);
    outputs(8636) <= not((layer0_outputs(7385)) xor (layer0_outputs(8537)));
    outputs(8637) <= not((layer0_outputs(3655)) or (layer0_outputs(8118)));
    outputs(8638) <= (layer0_outputs(4004)) or (layer0_outputs(1577));
    outputs(8639) <= not((layer0_outputs(741)) xor (layer0_outputs(489)));
    outputs(8640) <= not(layer0_outputs(7622));
    outputs(8641) <= (layer0_outputs(4771)) or (layer0_outputs(183));
    outputs(8642) <= not(layer0_outputs(1450)) or (layer0_outputs(9203));
    outputs(8643) <= (layer0_outputs(8508)) and not (layer0_outputs(3143));
    outputs(8644) <= not(layer0_outputs(6761)) or (layer0_outputs(2455));
    outputs(8645) <= not(layer0_outputs(1324));
    outputs(8646) <= (layer0_outputs(4788)) xor (layer0_outputs(9824));
    outputs(8647) <= not(layer0_outputs(6105)) or (layer0_outputs(9330));
    outputs(8648) <= not((layer0_outputs(5141)) or (layer0_outputs(5732)));
    outputs(8649) <= not((layer0_outputs(1275)) xor (layer0_outputs(3374)));
    outputs(8650) <= not(layer0_outputs(7482)) or (layer0_outputs(594));
    outputs(8651) <= not(layer0_outputs(7458));
    outputs(8652) <= not(layer0_outputs(2854));
    outputs(8653) <= not((layer0_outputs(1399)) xor (layer0_outputs(9323)));
    outputs(8654) <= not(layer0_outputs(1015));
    outputs(8655) <= (layer0_outputs(3715)) and not (layer0_outputs(6403));
    outputs(8656) <= (layer0_outputs(8835)) or (layer0_outputs(7088));
    outputs(8657) <= layer0_outputs(5355);
    outputs(8658) <= not((layer0_outputs(4582)) and (layer0_outputs(192)));
    outputs(8659) <= not(layer0_outputs(3098)) or (layer0_outputs(1947));
    outputs(8660) <= not((layer0_outputs(5312)) or (layer0_outputs(1412)));
    outputs(8661) <= not((layer0_outputs(6953)) xor (layer0_outputs(6711)));
    outputs(8662) <= (layer0_outputs(8616)) or (layer0_outputs(2577));
    outputs(8663) <= (layer0_outputs(6606)) and not (layer0_outputs(141));
    outputs(8664) <= (layer0_outputs(8337)) xor (layer0_outputs(2434));
    outputs(8665) <= not(layer0_outputs(1487));
    outputs(8666) <= not((layer0_outputs(10012)) xor (layer0_outputs(2924)));
    outputs(8667) <= not(layer0_outputs(9266));
    outputs(8668) <= (layer0_outputs(8914)) or (layer0_outputs(7344));
    outputs(8669) <= (layer0_outputs(3925)) and (layer0_outputs(3293));
    outputs(8670) <= not(layer0_outputs(9872));
    outputs(8671) <= (layer0_outputs(6471)) xor (layer0_outputs(2700));
    outputs(8672) <= (layer0_outputs(4192)) and not (layer0_outputs(5294));
    outputs(8673) <= layer0_outputs(969);
    outputs(8674) <= (layer0_outputs(671)) and (layer0_outputs(5854));
    outputs(8675) <= not(layer0_outputs(2655));
    outputs(8676) <= not((layer0_outputs(10177)) xor (layer0_outputs(3897)));
    outputs(8677) <= not((layer0_outputs(6521)) xor (layer0_outputs(7187)));
    outputs(8678) <= not((layer0_outputs(1229)) or (layer0_outputs(3960)));
    outputs(8679) <= (layer0_outputs(5920)) or (layer0_outputs(9752));
    outputs(8680) <= not((layer0_outputs(5646)) xor (layer0_outputs(3179)));
    outputs(8681) <= not((layer0_outputs(7567)) xor (layer0_outputs(1732)));
    outputs(8682) <= not(layer0_outputs(10059)) or (layer0_outputs(1128));
    outputs(8683) <= (layer0_outputs(7989)) xor (layer0_outputs(2468));
    outputs(8684) <= (layer0_outputs(4558)) xor (layer0_outputs(9366));
    outputs(8685) <= not(layer0_outputs(9730)) or (layer0_outputs(6575));
    outputs(8686) <= not(layer0_outputs(3131)) or (layer0_outputs(3377));
    outputs(8687) <= layer0_outputs(4760);
    outputs(8688) <= (layer0_outputs(9595)) xor (layer0_outputs(945));
    outputs(8689) <= not((layer0_outputs(1555)) xor (layer0_outputs(7449)));
    outputs(8690) <= layer0_outputs(5787);
    outputs(8691) <= layer0_outputs(1937);
    outputs(8692) <= layer0_outputs(9620);
    outputs(8693) <= not(layer0_outputs(1981));
    outputs(8694) <= not(layer0_outputs(6239)) or (layer0_outputs(9867));
    outputs(8695) <= (layer0_outputs(9821)) and not (layer0_outputs(8030));
    outputs(8696) <= not((layer0_outputs(5263)) xor (layer0_outputs(4761)));
    outputs(8697) <= not((layer0_outputs(6682)) xor (layer0_outputs(9302)));
    outputs(8698) <= (layer0_outputs(2085)) and not (layer0_outputs(2158));
    outputs(8699) <= layer0_outputs(4514);
    outputs(8700) <= layer0_outputs(6821);
    outputs(8701) <= not(layer0_outputs(9505));
    outputs(8702) <= (layer0_outputs(6846)) and not (layer0_outputs(4292));
    outputs(8703) <= not((layer0_outputs(723)) xor (layer0_outputs(5908)));
    outputs(8704) <= (layer0_outputs(7078)) and not (layer0_outputs(6577));
    outputs(8705) <= (layer0_outputs(7091)) xor (layer0_outputs(8537));
    outputs(8706) <= (layer0_outputs(9713)) and not (layer0_outputs(141));
    outputs(8707) <= not((layer0_outputs(3866)) xor (layer0_outputs(261)));
    outputs(8708) <= not(layer0_outputs(8251));
    outputs(8709) <= layer0_outputs(8078);
    outputs(8710) <= not((layer0_outputs(1715)) or (layer0_outputs(6152)));
    outputs(8711) <= (layer0_outputs(9135)) xor (layer0_outputs(36));
    outputs(8712) <= not(layer0_outputs(2963));
    outputs(8713) <= not(layer0_outputs(5670)) or (layer0_outputs(31));
    outputs(8714) <= layer0_outputs(9523);
    outputs(8715) <= not((layer0_outputs(8055)) and (layer0_outputs(9946)));
    outputs(8716) <= not(layer0_outputs(2424));
    outputs(8717) <= layer0_outputs(2394);
    outputs(8718) <= layer0_outputs(547);
    outputs(8719) <= not((layer0_outputs(1726)) and (layer0_outputs(7885)));
    outputs(8720) <= not((layer0_outputs(7481)) xor (layer0_outputs(9815)));
    outputs(8721) <= '1';
    outputs(8722) <= (layer0_outputs(3666)) and not (layer0_outputs(7886));
    outputs(8723) <= not((layer0_outputs(5968)) or (layer0_outputs(8973)));
    outputs(8724) <= layer0_outputs(4894);
    outputs(8725) <= not(layer0_outputs(7461)) or (layer0_outputs(7914));
    outputs(8726) <= (layer0_outputs(9365)) xor (layer0_outputs(3057));
    outputs(8727) <= not((layer0_outputs(2521)) and (layer0_outputs(4849)));
    outputs(8728) <= not((layer0_outputs(8282)) or (layer0_outputs(7775)));
    outputs(8729) <= not(layer0_outputs(3764));
    outputs(8730) <= not((layer0_outputs(1807)) xor (layer0_outputs(6781)));
    outputs(8731) <= not((layer0_outputs(10219)) or (layer0_outputs(7212)));
    outputs(8732) <= not((layer0_outputs(9222)) xor (layer0_outputs(3995)));
    outputs(8733) <= (layer0_outputs(8587)) or (layer0_outputs(9483));
    outputs(8734) <= not((layer0_outputs(9347)) xor (layer0_outputs(822)));
    outputs(8735) <= not((layer0_outputs(4033)) and (layer0_outputs(4061)));
    outputs(8736) <= layer0_outputs(8176);
    outputs(8737) <= (layer0_outputs(10019)) and not (layer0_outputs(2743));
    outputs(8738) <= (layer0_outputs(5726)) xor (layer0_outputs(7798));
    outputs(8739) <= (layer0_outputs(4383)) xor (layer0_outputs(2523));
    outputs(8740) <= layer0_outputs(597);
    outputs(8741) <= '1';
    outputs(8742) <= not(layer0_outputs(6210));
    outputs(8743) <= not(layer0_outputs(1669));
    outputs(8744) <= not((layer0_outputs(3423)) xor (layer0_outputs(7073)));
    outputs(8745) <= layer0_outputs(5812);
    outputs(8746) <= not(layer0_outputs(5503)) or (layer0_outputs(8600));
    outputs(8747) <= not((layer0_outputs(8524)) and (layer0_outputs(6735)));
    outputs(8748) <= not((layer0_outputs(1648)) or (layer0_outputs(77)));
    outputs(8749) <= not((layer0_outputs(2254)) xor (layer0_outputs(7705)));
    outputs(8750) <= not(layer0_outputs(3474));
    outputs(8751) <= not(layer0_outputs(3990));
    outputs(8752) <= layer0_outputs(9479);
    outputs(8753) <= layer0_outputs(6950);
    outputs(8754) <= layer0_outputs(6387);
    outputs(8755) <= (layer0_outputs(9360)) and (layer0_outputs(4023));
    outputs(8756) <= not((layer0_outputs(3706)) xor (layer0_outputs(552)));
    outputs(8757) <= not((layer0_outputs(2497)) xor (layer0_outputs(9975)));
    outputs(8758) <= not(layer0_outputs(3299));
    outputs(8759) <= (layer0_outputs(5308)) or (layer0_outputs(6564));
    outputs(8760) <= layer0_outputs(9587);
    outputs(8761) <= layer0_outputs(5797);
    outputs(8762) <= layer0_outputs(2201);
    outputs(8763) <= not((layer0_outputs(3622)) xor (layer0_outputs(7815)));
    outputs(8764) <= not(layer0_outputs(9262));
    outputs(8765) <= (layer0_outputs(8931)) xor (layer0_outputs(515));
    outputs(8766) <= layer0_outputs(8968);
    outputs(8767) <= layer0_outputs(5758);
    outputs(8768) <= (layer0_outputs(10107)) xor (layer0_outputs(7981));
    outputs(8769) <= layer0_outputs(1892);
    outputs(8770) <= not((layer0_outputs(8006)) xor (layer0_outputs(4657)));
    outputs(8771) <= (layer0_outputs(4686)) xor (layer0_outputs(4863));
    outputs(8772) <= not(layer0_outputs(7260));
    outputs(8773) <= (layer0_outputs(6317)) and not (layer0_outputs(5220));
    outputs(8774) <= not((layer0_outputs(4675)) xor (layer0_outputs(9828)));
    outputs(8775) <= (layer0_outputs(3857)) and (layer0_outputs(5987));
    outputs(8776) <= not((layer0_outputs(7074)) xor (layer0_outputs(9079)));
    outputs(8777) <= not(layer0_outputs(4529));
    outputs(8778) <= not((layer0_outputs(4739)) and (layer0_outputs(2351)));
    outputs(8779) <= not(layer0_outputs(4754));
    outputs(8780) <= (layer0_outputs(458)) or (layer0_outputs(6104));
    outputs(8781) <= not((layer0_outputs(4906)) xor (layer0_outputs(8436)));
    outputs(8782) <= (layer0_outputs(8041)) xor (layer0_outputs(9661));
    outputs(8783) <= (layer0_outputs(4706)) and not (layer0_outputs(4898));
    outputs(8784) <= not((layer0_outputs(5147)) xor (layer0_outputs(8321)));
    outputs(8785) <= not((layer0_outputs(3609)) and (layer0_outputs(8683)));
    outputs(8786) <= (layer0_outputs(5115)) xor (layer0_outputs(1970));
    outputs(8787) <= not(layer0_outputs(774)) or (layer0_outputs(7753));
    outputs(8788) <= not((layer0_outputs(3724)) and (layer0_outputs(7545)));
    outputs(8789) <= not((layer0_outputs(341)) xor (layer0_outputs(7065)));
    outputs(8790) <= (layer0_outputs(2870)) and not (layer0_outputs(1640));
    outputs(8791) <= not((layer0_outputs(3563)) xor (layer0_outputs(9088)));
    outputs(8792) <= not((layer0_outputs(6908)) and (layer0_outputs(2728)));
    outputs(8793) <= (layer0_outputs(3415)) xor (layer0_outputs(2573));
    outputs(8794) <= layer0_outputs(6113);
    outputs(8795) <= (layer0_outputs(4127)) xor (layer0_outputs(2287));
    outputs(8796) <= layer0_outputs(8763);
    outputs(8797) <= not(layer0_outputs(8103)) or (layer0_outputs(6136));
    outputs(8798) <= (layer0_outputs(5503)) or (layer0_outputs(6620));
    outputs(8799) <= not((layer0_outputs(4025)) xor (layer0_outputs(5945)));
    outputs(8800) <= not(layer0_outputs(5238));
    outputs(8801) <= not(layer0_outputs(2876));
    outputs(8802) <= (layer0_outputs(128)) xor (layer0_outputs(9110));
    outputs(8803) <= (layer0_outputs(8867)) xor (layer0_outputs(8226));
    outputs(8804) <= (layer0_outputs(2732)) xor (layer0_outputs(7402));
    outputs(8805) <= not(layer0_outputs(2444));
    outputs(8806) <= not(layer0_outputs(1199));
    outputs(8807) <= not(layer0_outputs(2805));
    outputs(8808) <= not((layer0_outputs(9893)) and (layer0_outputs(7386)));
    outputs(8809) <= layer0_outputs(1772);
    outputs(8810) <= (layer0_outputs(8807)) or (layer0_outputs(6745));
    outputs(8811) <= layer0_outputs(7526);
    outputs(8812) <= not(layer0_outputs(2792));
    outputs(8813) <= not(layer0_outputs(3562));
    outputs(8814) <= layer0_outputs(1394);
    outputs(8815) <= (layer0_outputs(4809)) and not (layer0_outputs(750));
    outputs(8816) <= (layer0_outputs(5909)) or (layer0_outputs(92));
    outputs(8817) <= not(layer0_outputs(6479)) or (layer0_outputs(4942));
    outputs(8818) <= (layer0_outputs(10069)) xor (layer0_outputs(510));
    outputs(8819) <= not((layer0_outputs(4242)) xor (layer0_outputs(8439)));
    outputs(8820) <= not(layer0_outputs(4964));
    outputs(8821) <= (layer0_outputs(9155)) xor (layer0_outputs(3559));
    outputs(8822) <= '1';
    outputs(8823) <= (layer0_outputs(8773)) and not (layer0_outputs(1065));
    outputs(8824) <= (layer0_outputs(6258)) and not (layer0_outputs(2056));
    outputs(8825) <= not((layer0_outputs(8276)) xor (layer0_outputs(1377)));
    outputs(8826) <= (layer0_outputs(8202)) xor (layer0_outputs(1033));
    outputs(8827) <= (layer0_outputs(2448)) xor (layer0_outputs(9680));
    outputs(8828) <= layer0_outputs(5044);
    outputs(8829) <= (layer0_outputs(6294)) and not (layer0_outputs(5791));
    outputs(8830) <= not((layer0_outputs(4987)) xor (layer0_outputs(2822)));
    outputs(8831) <= not((layer0_outputs(7982)) xor (layer0_outputs(6536)));
    outputs(8832) <= not(layer0_outputs(4130));
    outputs(8833) <= not((layer0_outputs(5227)) xor (layer0_outputs(2882)));
    outputs(8834) <= (layer0_outputs(2554)) xor (layer0_outputs(9174));
    outputs(8835) <= (layer0_outputs(8917)) xor (layer0_outputs(2624));
    outputs(8836) <= layer0_outputs(4039);
    outputs(8837) <= not(layer0_outputs(6133));
    outputs(8838) <= (layer0_outputs(1059)) and (layer0_outputs(5247));
    outputs(8839) <= layer0_outputs(970);
    outputs(8840) <= layer0_outputs(5482);
    outputs(8841) <= layer0_outputs(3803);
    outputs(8842) <= layer0_outputs(8691);
    outputs(8843) <= (layer0_outputs(3256)) or (layer0_outputs(1863));
    outputs(8844) <= not(layer0_outputs(2481)) or (layer0_outputs(3294));
    outputs(8845) <= not((layer0_outputs(2493)) xor (layer0_outputs(3872)));
    outputs(8846) <= not((layer0_outputs(9525)) xor (layer0_outputs(7185)));
    outputs(8847) <= not(layer0_outputs(8980)) or (layer0_outputs(6267));
    outputs(8848) <= (layer0_outputs(3920)) or (layer0_outputs(3667));
    outputs(8849) <= not(layer0_outputs(2846)) or (layer0_outputs(9070));
    outputs(8850) <= (layer0_outputs(7037)) and not (layer0_outputs(6500));
    outputs(8851) <= not((layer0_outputs(441)) or (layer0_outputs(8203)));
    outputs(8852) <= (layer0_outputs(5078)) xor (layer0_outputs(7192));
    outputs(8853) <= (layer0_outputs(9735)) or (layer0_outputs(8223));
    outputs(8854) <= not((layer0_outputs(163)) and (layer0_outputs(6006)));
    outputs(8855) <= not((layer0_outputs(1536)) xor (layer0_outputs(716)));
    outputs(8856) <= not(layer0_outputs(2238));
    outputs(8857) <= (layer0_outputs(2945)) and (layer0_outputs(2128));
    outputs(8858) <= (layer0_outputs(1789)) xor (layer0_outputs(6053));
    outputs(8859) <= not((layer0_outputs(9490)) xor (layer0_outputs(2903)));
    outputs(8860) <= (layer0_outputs(6707)) or (layer0_outputs(7587));
    outputs(8861) <= (layer0_outputs(447)) and not (layer0_outputs(5470));
    outputs(8862) <= layer0_outputs(9599);
    outputs(8863) <= layer0_outputs(616);
    outputs(8864) <= not((layer0_outputs(3466)) xor (layer0_outputs(3643)));
    outputs(8865) <= not((layer0_outputs(5908)) xor (layer0_outputs(5297)));
    outputs(8866) <= (layer0_outputs(5668)) and not (layer0_outputs(5688));
    outputs(8867) <= layer0_outputs(4196);
    outputs(8868) <= (layer0_outputs(5452)) or (layer0_outputs(6383));
    outputs(8869) <= (layer0_outputs(3957)) xor (layer0_outputs(2042));
    outputs(8870) <= not(layer0_outputs(6941));
    outputs(8871) <= layer0_outputs(7471);
    outputs(8872) <= not((layer0_outputs(3228)) xor (layer0_outputs(891)));
    outputs(8873) <= layer0_outputs(6022);
    outputs(8874) <= not((layer0_outputs(9219)) xor (layer0_outputs(7980)));
    outputs(8875) <= (layer0_outputs(6907)) xor (layer0_outputs(117));
    outputs(8876) <= not((layer0_outputs(962)) xor (layer0_outputs(375)));
    outputs(8877) <= (layer0_outputs(9456)) and not (layer0_outputs(3793));
    outputs(8878) <= (layer0_outputs(7927)) xor (layer0_outputs(3291));
    outputs(8879) <= layer0_outputs(5631);
    outputs(8880) <= not(layer0_outputs(8039)) or (layer0_outputs(3636));
    outputs(8881) <= not((layer0_outputs(3842)) and (layer0_outputs(8526)));
    outputs(8882) <= (layer0_outputs(5133)) and not (layer0_outputs(17));
    outputs(8883) <= not(layer0_outputs(6150));
    outputs(8884) <= not((layer0_outputs(4786)) xor (layer0_outputs(2938)));
    outputs(8885) <= layer0_outputs(926);
    outputs(8886) <= (layer0_outputs(9290)) xor (layer0_outputs(5971));
    outputs(8887) <= not(layer0_outputs(10067)) or (layer0_outputs(6644));
    outputs(8888) <= not((layer0_outputs(7344)) xor (layer0_outputs(5191)));
    outputs(8889) <= '1';
    outputs(8890) <= layer0_outputs(4606);
    outputs(8891) <= layer0_outputs(9016);
    outputs(8892) <= (layer0_outputs(5514)) xor (layer0_outputs(4659));
    outputs(8893) <= not((layer0_outputs(7367)) or (layer0_outputs(314)));
    outputs(8894) <= layer0_outputs(3886);
    outputs(8895) <= (layer0_outputs(3822)) xor (layer0_outputs(3520));
    outputs(8896) <= (layer0_outputs(6630)) and (layer0_outputs(6771));
    outputs(8897) <= not(layer0_outputs(3782));
    outputs(8898) <= not(layer0_outputs(10081));
    outputs(8899) <= not(layer0_outputs(8080));
    outputs(8900) <= not(layer0_outputs(5746)) or (layer0_outputs(7066));
    outputs(8901) <= (layer0_outputs(9534)) xor (layer0_outputs(3162));
    outputs(8902) <= layer0_outputs(6803);
    outputs(8903) <= not((layer0_outputs(4728)) xor (layer0_outputs(4364)));
    outputs(8904) <= layer0_outputs(5888);
    outputs(8905) <= (layer0_outputs(6753)) or (layer0_outputs(4861));
    outputs(8906) <= (layer0_outputs(5601)) or (layer0_outputs(9169));
    outputs(8907) <= (layer0_outputs(2975)) and not (layer0_outputs(7205));
    outputs(8908) <= (layer0_outputs(7580)) or (layer0_outputs(2132));
    outputs(8909) <= layer0_outputs(8052);
    outputs(8910) <= (layer0_outputs(10139)) and not (layer0_outputs(10058));
    outputs(8911) <= not(layer0_outputs(4214)) or (layer0_outputs(9138));
    outputs(8912) <= (layer0_outputs(5608)) xor (layer0_outputs(6078));
    outputs(8913) <= layer0_outputs(3287);
    outputs(8914) <= (layer0_outputs(2620)) or (layer0_outputs(4009));
    outputs(8915) <= not(layer0_outputs(1899)) or (layer0_outputs(7991));
    outputs(8916) <= not(layer0_outputs(5204));
    outputs(8917) <= not(layer0_outputs(1194)) or (layer0_outputs(6802));
    outputs(8918) <= layer0_outputs(188);
    outputs(8919) <= not(layer0_outputs(4311));
    outputs(8920) <= not((layer0_outputs(1408)) xor (layer0_outputs(10194)));
    outputs(8921) <= layer0_outputs(9454);
    outputs(8922) <= not(layer0_outputs(8536)) or (layer0_outputs(1161));
    outputs(8923) <= not((layer0_outputs(5073)) or (layer0_outputs(330)));
    outputs(8924) <= not((layer0_outputs(653)) and (layer0_outputs(1905)));
    outputs(8925) <= layer0_outputs(2886);
    outputs(8926) <= not((layer0_outputs(5143)) or (layer0_outputs(6139)));
    outputs(8927) <= (layer0_outputs(6416)) xor (layer0_outputs(7062));
    outputs(8928) <= (layer0_outputs(3717)) xor (layer0_outputs(1713));
    outputs(8929) <= not((layer0_outputs(1171)) xor (layer0_outputs(977)));
    outputs(8930) <= not((layer0_outputs(489)) xor (layer0_outputs(821)));
    outputs(8931) <= not(layer0_outputs(8942));
    outputs(8932) <= (layer0_outputs(1814)) or (layer0_outputs(7214));
    outputs(8933) <= not(layer0_outputs(229));
    outputs(8934) <= layer0_outputs(377);
    outputs(8935) <= not((layer0_outputs(4534)) xor (layer0_outputs(7937)));
    outputs(8936) <= layer0_outputs(7170);
    outputs(8937) <= not((layer0_outputs(1285)) xor (layer0_outputs(4217)));
    outputs(8938) <= (layer0_outputs(7416)) and not (layer0_outputs(747));
    outputs(8939) <= not(layer0_outputs(8801));
    outputs(8940) <= (layer0_outputs(1035)) or (layer0_outputs(9997));
    outputs(8941) <= not(layer0_outputs(2829));
    outputs(8942) <= not(layer0_outputs(4382)) or (layer0_outputs(7547));
    outputs(8943) <= (layer0_outputs(6279)) xor (layer0_outputs(172));
    outputs(8944) <= layer0_outputs(4535);
    outputs(8945) <= not(layer0_outputs(6788));
    outputs(8946) <= not(layer0_outputs(7650));
    outputs(8947) <= (layer0_outputs(7415)) and (layer0_outputs(24));
    outputs(8948) <= (layer0_outputs(1796)) xor (layer0_outputs(6137));
    outputs(8949) <= layer0_outputs(4593);
    outputs(8950) <= not((layer0_outputs(3207)) and (layer0_outputs(4388)));
    outputs(8951) <= not(layer0_outputs(1650)) or (layer0_outputs(7500));
    outputs(8952) <= not((layer0_outputs(8597)) and (layer0_outputs(3394)));
    outputs(8953) <= not((layer0_outputs(2294)) xor (layer0_outputs(2334)));
    outputs(8954) <= not(layer0_outputs(443)) or (layer0_outputs(1050));
    outputs(8955) <= not(layer0_outputs(5185));
    outputs(8956) <= not(layer0_outputs(493)) or (layer0_outputs(3379));
    outputs(8957) <= not((layer0_outputs(1496)) and (layer0_outputs(6945)));
    outputs(8958) <= (layer0_outputs(6719)) xor (layer0_outputs(1518));
    outputs(8959) <= layer0_outputs(2847);
    outputs(8960) <= not((layer0_outputs(2138)) xor (layer0_outputs(3147)));
    outputs(8961) <= (layer0_outputs(7331)) and (layer0_outputs(1306));
    outputs(8962) <= not(layer0_outputs(8866)) or (layer0_outputs(3422));
    outputs(8963) <= not(layer0_outputs(2728));
    outputs(8964) <= not((layer0_outputs(9255)) and (layer0_outputs(8668)));
    outputs(8965) <= not((layer0_outputs(6435)) and (layer0_outputs(328)));
    outputs(8966) <= not((layer0_outputs(165)) xor (layer0_outputs(9312)));
    outputs(8967) <= not((layer0_outputs(303)) and (layer0_outputs(7359)));
    outputs(8968) <= not((layer0_outputs(8564)) and (layer0_outputs(2103)));
    outputs(8969) <= (layer0_outputs(9889)) xor (layer0_outputs(2630));
    outputs(8970) <= not((layer0_outputs(4915)) xor (layer0_outputs(1822)));
    outputs(8971) <= (layer0_outputs(5050)) and (layer0_outputs(1788));
    outputs(8972) <= not(layer0_outputs(4179));
    outputs(8973) <= layer0_outputs(7944);
    outputs(8974) <= (layer0_outputs(6066)) xor (layer0_outputs(3831));
    outputs(8975) <= (layer0_outputs(3099)) and not (layer0_outputs(4336));
    outputs(8976) <= not((layer0_outputs(7390)) and (layer0_outputs(4626)));
    outputs(8977) <= not(layer0_outputs(5582)) or (layer0_outputs(5607));
    outputs(8978) <= (layer0_outputs(7933)) and not (layer0_outputs(888));
    outputs(8979) <= not(layer0_outputs(10136));
    outputs(8980) <= (layer0_outputs(951)) xor (layer0_outputs(275));
    outputs(8981) <= layer0_outputs(9473);
    outputs(8982) <= not(layer0_outputs(2694));
    outputs(8983) <= (layer0_outputs(4604)) and not (layer0_outputs(5112));
    outputs(8984) <= layer0_outputs(8562);
    outputs(8985) <= (layer0_outputs(4352)) xor (layer0_outputs(6513));
    outputs(8986) <= not((layer0_outputs(1677)) xor (layer0_outputs(9570)));
    outputs(8987) <= not((layer0_outputs(3793)) xor (layer0_outputs(5711)));
    outputs(8988) <= not(layer0_outputs(9878)) or (layer0_outputs(10112));
    outputs(8989) <= layer0_outputs(100);
    outputs(8990) <= not((layer0_outputs(10192)) xor (layer0_outputs(3787)));
    outputs(8991) <= layer0_outputs(4817);
    outputs(8992) <= (layer0_outputs(3400)) xor (layer0_outputs(3526));
    outputs(8993) <= not(layer0_outputs(512)) or (layer0_outputs(3154));
    outputs(8994) <= not(layer0_outputs(8967)) or (layer0_outputs(552));
    outputs(8995) <= (layer0_outputs(157)) and not (layer0_outputs(3680));
    outputs(8996) <= not(layer0_outputs(1896));
    outputs(8997) <= not(layer0_outputs(1000));
    outputs(8998) <= (layer0_outputs(3901)) xor (layer0_outputs(4701));
    outputs(8999) <= layer0_outputs(6384);
    outputs(9000) <= not(layer0_outputs(8993));
    outputs(9001) <= not(layer0_outputs(6157)) or (layer0_outputs(3640));
    outputs(9002) <= (layer0_outputs(7975)) and not (layer0_outputs(3951));
    outputs(9003) <= not(layer0_outputs(350)) or (layer0_outputs(9509));
    outputs(9004) <= (layer0_outputs(9138)) xor (layer0_outputs(7113));
    outputs(9005) <= not((layer0_outputs(9726)) xor (layer0_outputs(2773)));
    outputs(9006) <= (layer0_outputs(3610)) and not (layer0_outputs(6160));
    outputs(9007) <= layer0_outputs(2856);
    outputs(9008) <= not(layer0_outputs(6751));
    outputs(9009) <= (layer0_outputs(623)) or (layer0_outputs(6183));
    outputs(9010) <= (layer0_outputs(2661)) and not (layer0_outputs(8421));
    outputs(9011) <= (layer0_outputs(7125)) xor (layer0_outputs(9507));
    outputs(9012) <= (layer0_outputs(3174)) and (layer0_outputs(5699));
    outputs(9013) <= (layer0_outputs(3037)) or (layer0_outputs(776));
    outputs(9014) <= layer0_outputs(1018);
    outputs(9015) <= (layer0_outputs(2919)) xor (layer0_outputs(6162));
    outputs(9016) <= not(layer0_outputs(6952)) or (layer0_outputs(9909));
    outputs(9017) <= layer0_outputs(9038);
    outputs(9018) <= not(layer0_outputs(7070)) or (layer0_outputs(5694));
    outputs(9019) <= not(layer0_outputs(1758));
    outputs(9020) <= (layer0_outputs(3703)) xor (layer0_outputs(9545));
    outputs(9021) <= layer0_outputs(1902);
    outputs(9022) <= not(layer0_outputs(7430)) or (layer0_outputs(3326));
    outputs(9023) <= (layer0_outputs(816)) xor (layer0_outputs(3710));
    outputs(9024) <= (layer0_outputs(9693)) and not (layer0_outputs(7913));
    outputs(9025) <= (layer0_outputs(6378)) xor (layer0_outputs(5058));
    outputs(9026) <= layer0_outputs(6663);
    outputs(9027) <= (layer0_outputs(3354)) and not (layer0_outputs(928));
    outputs(9028) <= not((layer0_outputs(8267)) xor (layer0_outputs(3224)));
    outputs(9029) <= not((layer0_outputs(1252)) xor (layer0_outputs(4525)));
    outputs(9030) <= not((layer0_outputs(4118)) xor (layer0_outputs(5689)));
    outputs(9031) <= not(layer0_outputs(10156));
    outputs(9032) <= (layer0_outputs(9243)) xor (layer0_outputs(9019));
    outputs(9033) <= not(layer0_outputs(1129));
    outputs(9034) <= (layer0_outputs(9307)) xor (layer0_outputs(8398));
    outputs(9035) <= not(layer0_outputs(7954));
    outputs(9036) <= (layer0_outputs(4223)) and (layer0_outputs(6906));
    outputs(9037) <= (layer0_outputs(7024)) xor (layer0_outputs(9432));
    outputs(9038) <= (layer0_outputs(3290)) and not (layer0_outputs(1529));
    outputs(9039) <= not(layer0_outputs(3245));
    outputs(9040) <= not((layer0_outputs(8019)) and (layer0_outputs(5844)));
    outputs(9041) <= not((layer0_outputs(1040)) xor (layer0_outputs(9788)));
    outputs(9042) <= not((layer0_outputs(7549)) or (layer0_outputs(8824)));
    outputs(9043) <= not((layer0_outputs(818)) xor (layer0_outputs(3873)));
    outputs(9044) <= not((layer0_outputs(8856)) xor (layer0_outputs(9794)));
    outputs(9045) <= layer0_outputs(5952);
    outputs(9046) <= not(layer0_outputs(9691));
    outputs(9047) <= (layer0_outputs(3779)) and not (layer0_outputs(167));
    outputs(9048) <= not(layer0_outputs(422));
    outputs(9049) <= not(layer0_outputs(7355));
    outputs(9050) <= (layer0_outputs(1612)) or (layer0_outputs(8444));
    outputs(9051) <= not((layer0_outputs(8790)) xor (layer0_outputs(3134)));
    outputs(9052) <= not((layer0_outputs(9426)) xor (layer0_outputs(7152)));
    outputs(9053) <= not(layer0_outputs(5484)) or (layer0_outputs(3635));
    outputs(9054) <= not((layer0_outputs(4825)) or (layer0_outputs(3401)));
    outputs(9055) <= layer0_outputs(9933);
    outputs(9056) <= (layer0_outputs(3587)) xor (layer0_outputs(6804));
    outputs(9057) <= (layer0_outputs(6185)) and (layer0_outputs(3613));
    outputs(9058) <= not((layer0_outputs(7242)) and (layer0_outputs(1119)));
    outputs(9059) <= not(layer0_outputs(8500)) or (layer0_outputs(4594));
    outputs(9060) <= not(layer0_outputs(8938));
    outputs(9061) <= '1';
    outputs(9062) <= layer0_outputs(4950);
    outputs(9063) <= (layer0_outputs(4665)) or (layer0_outputs(9385));
    outputs(9064) <= layer0_outputs(7335);
    outputs(9065) <= (layer0_outputs(9235)) xor (layer0_outputs(3196));
    outputs(9066) <= not(layer0_outputs(9745));
    outputs(9067) <= layer0_outputs(2349);
    outputs(9068) <= (layer0_outputs(9923)) and (layer0_outputs(6340));
    outputs(9069) <= not((layer0_outputs(7707)) and (layer0_outputs(2321)));
    outputs(9070) <= not(layer0_outputs(457));
    outputs(9071) <= layer0_outputs(9708);
    outputs(9072) <= not(layer0_outputs(5305));
    outputs(9073) <= not((layer0_outputs(8425)) or (layer0_outputs(3143)));
    outputs(9074) <= (layer0_outputs(6548)) or (layer0_outputs(5370));
    outputs(9075) <= not(layer0_outputs(9208));
    outputs(9076) <= layer0_outputs(1641);
    outputs(9077) <= not((layer0_outputs(10024)) xor (layer0_outputs(1692)));
    outputs(9078) <= not((layer0_outputs(6213)) xor (layer0_outputs(4414)));
    outputs(9079) <= not((layer0_outputs(5588)) xor (layer0_outputs(1750)));
    outputs(9080) <= (layer0_outputs(804)) xor (layer0_outputs(5027));
    outputs(9081) <= layer0_outputs(9033);
    outputs(9082) <= (layer0_outputs(4207)) xor (layer0_outputs(7351));
    outputs(9083) <= not(layer0_outputs(3739)) or (layer0_outputs(1091));
    outputs(9084) <= (layer0_outputs(7256)) or (layer0_outputs(5850));
    outputs(9085) <= not((layer0_outputs(9208)) or (layer0_outputs(6695)));
    outputs(9086) <= not((layer0_outputs(1257)) xor (layer0_outputs(2711)));
    outputs(9087) <= not((layer0_outputs(6362)) xor (layer0_outputs(27)));
    outputs(9088) <= (layer0_outputs(3701)) xor (layer0_outputs(6867));
    outputs(9089) <= (layer0_outputs(7583)) xor (layer0_outputs(2345));
    outputs(9090) <= not(layer0_outputs(124)) or (layer0_outputs(1460));
    outputs(9091) <= not(layer0_outputs(7517)) or (layer0_outputs(3826));
    outputs(9092) <= (layer0_outputs(5471)) xor (layer0_outputs(9924));
    outputs(9093) <= not((layer0_outputs(3445)) xor (layer0_outputs(9025)));
    outputs(9094) <= (layer0_outputs(8140)) xor (layer0_outputs(1311));
    outputs(9095) <= layer0_outputs(8169);
    outputs(9096) <= not(layer0_outputs(2258));
    outputs(9097) <= not(layer0_outputs(8113)) or (layer0_outputs(5797));
    outputs(9098) <= not((layer0_outputs(4126)) or (layer0_outputs(9107)));
    outputs(9099) <= not(layer0_outputs(8358)) or (layer0_outputs(9021));
    outputs(9100) <= (layer0_outputs(8773)) and not (layer0_outputs(5038));
    outputs(9101) <= not((layer0_outputs(1148)) xor (layer0_outputs(565)));
    outputs(9102) <= not(layer0_outputs(1407));
    outputs(9103) <= (layer0_outputs(5994)) xor (layer0_outputs(9486));
    outputs(9104) <= not((layer0_outputs(9235)) and (layer0_outputs(810)));
    outputs(9105) <= (layer0_outputs(5157)) xor (layer0_outputs(1691));
    outputs(9106) <= layer0_outputs(10015);
    outputs(9107) <= not((layer0_outputs(2840)) xor (layer0_outputs(3270)));
    outputs(9108) <= not(layer0_outputs(3926));
    outputs(9109) <= layer0_outputs(6754);
    outputs(9110) <= '1';
    outputs(9111) <= (layer0_outputs(1192)) or (layer0_outputs(1424));
    outputs(9112) <= not((layer0_outputs(7231)) xor (layer0_outputs(9920)));
    outputs(9113) <= not((layer0_outputs(5369)) xor (layer0_outputs(3987)));
    outputs(9114) <= (layer0_outputs(6388)) xor (layer0_outputs(262));
    outputs(9115) <= not((layer0_outputs(7616)) and (layer0_outputs(6079)));
    outputs(9116) <= layer0_outputs(613);
    outputs(9117) <= not(layer0_outputs(5630));
    outputs(9118) <= (layer0_outputs(2772)) xor (layer0_outputs(1059));
    outputs(9119) <= not((layer0_outputs(3690)) xor (layer0_outputs(1934)));
    outputs(9120) <= not((layer0_outputs(6918)) and (layer0_outputs(4808)));
    outputs(9121) <= layer0_outputs(8766);
    outputs(9122) <= layer0_outputs(7591);
    outputs(9123) <= layer0_outputs(7711);
    outputs(9124) <= not((layer0_outputs(709)) xor (layer0_outputs(1528)));
    outputs(9125) <= (layer0_outputs(2467)) and not (layer0_outputs(7684));
    outputs(9126) <= not((layer0_outputs(9037)) xor (layer0_outputs(5647)));
    outputs(9127) <= not(layer0_outputs(9380)) or (layer0_outputs(9081));
    outputs(9128) <= layer0_outputs(4177);
    outputs(9129) <= not(layer0_outputs(1486)) or (layer0_outputs(7704));
    outputs(9130) <= not(layer0_outputs(2155));
    outputs(9131) <= (layer0_outputs(9344)) xor (layer0_outputs(2634));
    outputs(9132) <= not((layer0_outputs(5604)) xor (layer0_outputs(2003)));
    outputs(9133) <= (layer0_outputs(4468)) xor (layer0_outputs(8720));
    outputs(9134) <= (layer0_outputs(5559)) xor (layer0_outputs(3215));
    outputs(9135) <= not((layer0_outputs(9126)) xor (layer0_outputs(4446)));
    outputs(9136) <= (layer0_outputs(5717)) xor (layer0_outputs(3869));
    outputs(9137) <= not((layer0_outputs(2293)) or (layer0_outputs(2189)));
    outputs(9138) <= (layer0_outputs(5644)) and (layer0_outputs(7645));
    outputs(9139) <= not((layer0_outputs(6530)) and (layer0_outputs(8212)));
    outputs(9140) <= (layer0_outputs(2613)) and not (layer0_outputs(8692));
    outputs(9141) <= layer0_outputs(3381);
    outputs(9142) <= layer0_outputs(9517);
    outputs(9143) <= not(layer0_outputs(3843)) or (layer0_outputs(3588));
    outputs(9144) <= not(layer0_outputs(10181));
    outputs(9145) <= not((layer0_outputs(7671)) xor (layer0_outputs(4135)));
    outputs(9146) <= (layer0_outputs(1011)) xor (layer0_outputs(4730));
    outputs(9147) <= not(layer0_outputs(9374)) or (layer0_outputs(10182));
    outputs(9148) <= layer0_outputs(883);
    outputs(9149) <= not(layer0_outputs(4723));
    outputs(9150) <= (layer0_outputs(5395)) or (layer0_outputs(5487));
    outputs(9151) <= not((layer0_outputs(4730)) xor (layer0_outputs(6933)));
    outputs(9152) <= (layer0_outputs(9663)) and not (layer0_outputs(4763));
    outputs(9153) <= not(layer0_outputs(5021));
    outputs(9154) <= not(layer0_outputs(1230));
    outputs(9155) <= layer0_outputs(8755);
    outputs(9156) <= (layer0_outputs(7076)) xor (layer0_outputs(72));
    outputs(9157) <= (layer0_outputs(2516)) and not (layer0_outputs(9165));
    outputs(9158) <= (layer0_outputs(3202)) xor (layer0_outputs(481));
    outputs(9159) <= not(layer0_outputs(5052));
    outputs(9160) <= layer0_outputs(6806);
    outputs(9161) <= not((layer0_outputs(10185)) or (layer0_outputs(3170)));
    outputs(9162) <= not(layer0_outputs(7012));
    outputs(9163) <= not(layer0_outputs(464));
    outputs(9164) <= not((layer0_outputs(2916)) xor (layer0_outputs(2025)));
    outputs(9165) <= (layer0_outputs(6467)) or (layer0_outputs(5984));
    outputs(9166) <= not((layer0_outputs(932)) or (layer0_outputs(6138)));
    outputs(9167) <= not(layer0_outputs(2193));
    outputs(9168) <= layer0_outputs(1020);
    outputs(9169) <= layer0_outputs(1573);
    outputs(9170) <= not((layer0_outputs(9835)) and (layer0_outputs(882)));
    outputs(9171) <= not((layer0_outputs(5341)) and (layer0_outputs(350)));
    outputs(9172) <= (layer0_outputs(9120)) xor (layer0_outputs(7007));
    outputs(9173) <= not(layer0_outputs(1180));
    outputs(9174) <= (layer0_outputs(6119)) and (layer0_outputs(8491));
    outputs(9175) <= '1';
    outputs(9176) <= (layer0_outputs(4857)) and not (layer0_outputs(6408));
    outputs(9177) <= layer0_outputs(956);
    outputs(9178) <= not(layer0_outputs(1480));
    outputs(9179) <= not(layer0_outputs(8540)) or (layer0_outputs(1198));
    outputs(9180) <= (layer0_outputs(9154)) xor (layer0_outputs(4866));
    outputs(9181) <= (layer0_outputs(7585)) and not (layer0_outputs(8179));
    outputs(9182) <= not(layer0_outputs(8202));
    outputs(9183) <= (layer0_outputs(4853)) xor (layer0_outputs(1717));
    outputs(9184) <= not((layer0_outputs(7727)) and (layer0_outputs(3040)));
    outputs(9185) <= (layer0_outputs(6199)) and not (layer0_outputs(1023));
    outputs(9186) <= not(layer0_outputs(3966));
    outputs(9187) <= not(layer0_outputs(1088));
    outputs(9188) <= layer0_outputs(4817);
    outputs(9189) <= not(layer0_outputs(7468));
    outputs(9190) <= not((layer0_outputs(1741)) xor (layer0_outputs(6730)));
    outputs(9191) <= not(layer0_outputs(2014));
    outputs(9192) <= not((layer0_outputs(2629)) and (layer0_outputs(2615)));
    outputs(9193) <= '0';
    outputs(9194) <= layer0_outputs(1642);
    outputs(9195) <= not(layer0_outputs(8173)) or (layer0_outputs(9630));
    outputs(9196) <= not((layer0_outputs(9082)) or (layer0_outputs(3885)));
    outputs(9197) <= not(layer0_outputs(4182)) or (layer0_outputs(1804));
    outputs(9198) <= layer0_outputs(10023);
    outputs(9199) <= not((layer0_outputs(9443)) xor (layer0_outputs(7617)));
    outputs(9200) <= not(layer0_outputs(4468));
    outputs(9201) <= (layer0_outputs(9797)) or (layer0_outputs(6786));
    outputs(9202) <= layer0_outputs(4254);
    outputs(9203) <= layer0_outputs(3962);
    outputs(9204) <= layer0_outputs(2689);
    outputs(9205) <= (layer0_outputs(4895)) and not (layer0_outputs(2287));
    outputs(9206) <= not((layer0_outputs(5028)) xor (layer0_outputs(3282)));
    outputs(9207) <= (layer0_outputs(2691)) and not (layer0_outputs(627));
    outputs(9208) <= not(layer0_outputs(2746));
    outputs(9209) <= layer0_outputs(6091);
    outputs(9210) <= layer0_outputs(4635);
    outputs(9211) <= layer0_outputs(4688);
    outputs(9212) <= layer0_outputs(5188);
    outputs(9213) <= not((layer0_outputs(7610)) xor (layer0_outputs(1014)));
    outputs(9214) <= layer0_outputs(2905);
    outputs(9215) <= (layer0_outputs(6470)) and not (layer0_outputs(4310));
    outputs(9216) <= not(layer0_outputs(1654)) or (layer0_outputs(6170));
    outputs(9217) <= layer0_outputs(2417);
    outputs(9218) <= (layer0_outputs(3480)) xor (layer0_outputs(7922));
    outputs(9219) <= (layer0_outputs(4787)) and not (layer0_outputs(5470));
    outputs(9220) <= not((layer0_outputs(2474)) or (layer0_outputs(4540)));
    outputs(9221) <= (layer0_outputs(9579)) and not (layer0_outputs(6730));
    outputs(9222) <= (layer0_outputs(1514)) xor (layer0_outputs(6141));
    outputs(9223) <= (layer0_outputs(2819)) and (layer0_outputs(4273));
    outputs(9224) <= layer0_outputs(5998);
    outputs(9225) <= not((layer0_outputs(5025)) xor (layer0_outputs(2723)));
    outputs(9226) <= not(layer0_outputs(6612)) or (layer0_outputs(3690));
    outputs(9227) <= not(layer0_outputs(2392));
    outputs(9228) <= not(layer0_outputs(9212)) or (layer0_outputs(3907));
    outputs(9229) <= (layer0_outputs(7122)) xor (layer0_outputs(700));
    outputs(9230) <= layer0_outputs(7109);
    outputs(9231) <= not((layer0_outputs(2083)) xor (layer0_outputs(7555)));
    outputs(9232) <= (layer0_outputs(8714)) xor (layer0_outputs(1830));
    outputs(9233) <= not((layer0_outputs(500)) xor (layer0_outputs(2992)));
    outputs(9234) <= not((layer0_outputs(7426)) xor (layer0_outputs(10126)));
    outputs(9235) <= '1';
    outputs(9236) <= layer0_outputs(6083);
    outputs(9237) <= (layer0_outputs(8615)) and (layer0_outputs(9557));
    outputs(9238) <= (layer0_outputs(8557)) and (layer0_outputs(8021));
    outputs(9239) <= not(layer0_outputs(1611));
    outputs(9240) <= (layer0_outputs(4964)) and not (layer0_outputs(3543));
    outputs(9241) <= not(layer0_outputs(944));
    outputs(9242) <= (layer0_outputs(10239)) and not (layer0_outputs(10119));
    outputs(9243) <= layer0_outputs(9721);
    outputs(9244) <= not(layer0_outputs(9479));
    outputs(9245) <= layer0_outputs(7866);
    outputs(9246) <= (layer0_outputs(7148)) xor (layer0_outputs(5337));
    outputs(9247) <= not(layer0_outputs(602));
    outputs(9248) <= (layer0_outputs(6478)) xor (layer0_outputs(6243));
    outputs(9249) <= (layer0_outputs(4594)) and (layer0_outputs(7612));
    outputs(9250) <= not((layer0_outputs(9694)) xor (layer0_outputs(9300)));
    outputs(9251) <= not((layer0_outputs(7239)) xor (layer0_outputs(6819)));
    outputs(9252) <= not((layer0_outputs(8260)) xor (layer0_outputs(8227)));
    outputs(9253) <= not(layer0_outputs(1628));
    outputs(9254) <= (layer0_outputs(346)) and (layer0_outputs(4324));
    outputs(9255) <= not((layer0_outputs(8463)) or (layer0_outputs(2521)));
    outputs(9256) <= not(layer0_outputs(10062)) or (layer0_outputs(7803));
    outputs(9257) <= (layer0_outputs(9371)) and not (layer0_outputs(4219));
    outputs(9258) <= not((layer0_outputs(4610)) xor (layer0_outputs(3553)));
    outputs(9259) <= (layer0_outputs(3010)) xor (layer0_outputs(9090));
    outputs(9260) <= layer0_outputs(1695);
    outputs(9261) <= (layer0_outputs(8518)) xor (layer0_outputs(6446));
    outputs(9262) <= not((layer0_outputs(4546)) or (layer0_outputs(5889)));
    outputs(9263) <= (layer0_outputs(5759)) and not (layer0_outputs(2092));
    outputs(9264) <= not(layer0_outputs(5927));
    outputs(9265) <= (layer0_outputs(355)) and not (layer0_outputs(3449));
    outputs(9266) <= not((layer0_outputs(4790)) or (layer0_outputs(8357)));
    outputs(9267) <= layer0_outputs(5521);
    outputs(9268) <= not((layer0_outputs(9733)) or (layer0_outputs(6784)));
    outputs(9269) <= (layer0_outputs(8483)) xor (layer0_outputs(5975));
    outputs(9270) <= (layer0_outputs(5765)) or (layer0_outputs(2486));
    outputs(9271) <= (layer0_outputs(5073)) and not (layer0_outputs(3797));
    outputs(9272) <= not((layer0_outputs(8911)) xor (layer0_outputs(9488)));
    outputs(9273) <= not((layer0_outputs(655)) or (layer0_outputs(928)));
    outputs(9274) <= layer0_outputs(5910);
    outputs(9275) <= not(layer0_outputs(1932));
    outputs(9276) <= not((layer0_outputs(1276)) or (layer0_outputs(4493)));
    outputs(9277) <= (layer0_outputs(652)) and not (layer0_outputs(7525));
    outputs(9278) <= layer0_outputs(5289);
    outputs(9279) <= (layer0_outputs(7822)) and not (layer0_outputs(7770));
    outputs(9280) <= not((layer0_outputs(5845)) or (layer0_outputs(7684)));
    outputs(9281) <= (layer0_outputs(5245)) xor (layer0_outputs(6517));
    outputs(9282) <= not(layer0_outputs(1809));
    outputs(9283) <= layer0_outputs(2592);
    outputs(9284) <= '0';
    outputs(9285) <= not(layer0_outputs(465));
    outputs(9286) <= not(layer0_outputs(8595));
    outputs(9287) <= (layer0_outputs(8893)) and not (layer0_outputs(7959));
    outputs(9288) <= not((layer0_outputs(8068)) xor (layer0_outputs(9559)));
    outputs(9289) <= layer0_outputs(1551);
    outputs(9290) <= '0';
    outputs(9291) <= not(layer0_outputs(7158));
    outputs(9292) <= not((layer0_outputs(354)) xor (layer0_outputs(6542)));
    outputs(9293) <= layer0_outputs(3437);
    outputs(9294) <= layer0_outputs(4236);
    outputs(9295) <= not((layer0_outputs(4306)) and (layer0_outputs(7686)));
    outputs(9296) <= not(layer0_outputs(4313)) or (layer0_outputs(1986));
    outputs(9297) <= not(layer0_outputs(8690));
    outputs(9298) <= (layer0_outputs(1916)) and not (layer0_outputs(9133));
    outputs(9299) <= layer0_outputs(2988);
    outputs(9300) <= (layer0_outputs(5272)) and (layer0_outputs(4447));
    outputs(9301) <= '0';
    outputs(9302) <= not((layer0_outputs(6346)) xor (layer0_outputs(8598)));
    outputs(9303) <= layer0_outputs(714);
    outputs(9304) <= layer0_outputs(5642);
    outputs(9305) <= (layer0_outputs(3081)) and not (layer0_outputs(5650));
    outputs(9306) <= not(layer0_outputs(430));
    outputs(9307) <= (layer0_outputs(9102)) xor (layer0_outputs(5420));
    outputs(9308) <= (layer0_outputs(5840)) xor (layer0_outputs(7834));
    outputs(9309) <= (layer0_outputs(2961)) and (layer0_outputs(6815));
    outputs(9310) <= not(layer0_outputs(3008));
    outputs(9311) <= (layer0_outputs(1997)) xor (layer0_outputs(836));
    outputs(9312) <= not(layer0_outputs(5311));
    outputs(9313) <= (layer0_outputs(7818)) xor (layer0_outputs(4828));
    outputs(9314) <= (layer0_outputs(7566)) xor (layer0_outputs(2974));
    outputs(9315) <= (layer0_outputs(2250)) and not (layer0_outputs(1619));
    outputs(9316) <= (layer0_outputs(10183)) and (layer0_outputs(4324));
    outputs(9317) <= (layer0_outputs(6198)) and (layer0_outputs(3700));
    outputs(9318) <= (layer0_outputs(8528)) xor (layer0_outputs(5978));
    outputs(9319) <= not(layer0_outputs(5156));
    outputs(9320) <= (layer0_outputs(1302)) and not (layer0_outputs(8493));
    outputs(9321) <= not((layer0_outputs(1427)) xor (layer0_outputs(3774)));
    outputs(9322) <= (layer0_outputs(3090)) and not (layer0_outputs(2644));
    outputs(9323) <= not((layer0_outputs(3712)) or (layer0_outputs(399)));
    outputs(9324) <= not((layer0_outputs(6641)) or (layer0_outputs(4074)));
    outputs(9325) <= (layer0_outputs(7614)) xor (layer0_outputs(1458));
    outputs(9326) <= (layer0_outputs(4109)) and not (layer0_outputs(2769));
    outputs(9327) <= (layer0_outputs(9871)) and not (layer0_outputs(8509));
    outputs(9328) <= not(layer0_outputs(5008));
    outputs(9329) <= not((layer0_outputs(1852)) xor (layer0_outputs(9584)));
    outputs(9330) <= not(layer0_outputs(1511));
    outputs(9331) <= not((layer0_outputs(1214)) xor (layer0_outputs(4390)));
    outputs(9332) <= not((layer0_outputs(2263)) xor (layer0_outputs(6892)));
    outputs(9333) <= not((layer0_outputs(5550)) xor (layer0_outputs(3370)));
    outputs(9334) <= not(layer0_outputs(7039)) or (layer0_outputs(8123));
    outputs(9335) <= not(layer0_outputs(4461));
    outputs(9336) <= layer0_outputs(3804);
    outputs(9337) <= (layer0_outputs(3237)) xor (layer0_outputs(4982));
    outputs(9338) <= (layer0_outputs(8798)) or (layer0_outputs(2179));
    outputs(9339) <= not((layer0_outputs(4491)) or (layer0_outputs(9186)));
    outputs(9340) <= not((layer0_outputs(1327)) or (layer0_outputs(7904)));
    outputs(9341) <= layer0_outputs(7564);
    outputs(9342) <= layer0_outputs(1187);
    outputs(9343) <= (layer0_outputs(2459)) and (layer0_outputs(4401));
    outputs(9344) <= (layer0_outputs(4264)) xor (layer0_outputs(8566));
    outputs(9345) <= (layer0_outputs(8759)) and not (layer0_outputs(6830));
    outputs(9346) <= layer0_outputs(989);
    outputs(9347) <= not(layer0_outputs(8409));
    outputs(9348) <= (layer0_outputs(9600)) and not (layer0_outputs(5533));
    outputs(9349) <= (layer0_outputs(9611)) and not (layer0_outputs(4781));
    outputs(9350) <= (layer0_outputs(5218)) and (layer0_outputs(403));
    outputs(9351) <= (layer0_outputs(6925)) and not (layer0_outputs(9619));
    outputs(9352) <= layer0_outputs(6205);
    outputs(9353) <= layer0_outputs(4868);
    outputs(9354) <= layer0_outputs(1713);
    outputs(9355) <= (layer0_outputs(4628)) or (layer0_outputs(1384));
    outputs(9356) <= (layer0_outputs(8093)) xor (layer0_outputs(2106));
    outputs(9357) <= not(layer0_outputs(5280)) or (layer0_outputs(1492));
    outputs(9358) <= layer0_outputs(9846);
    outputs(9359) <= (layer0_outputs(9055)) and not (layer0_outputs(6112));
    outputs(9360) <= not((layer0_outputs(2560)) or (layer0_outputs(8721)));
    outputs(9361) <= not((layer0_outputs(9617)) xor (layer0_outputs(149)));
    outputs(9362) <= layer0_outputs(9228);
    outputs(9363) <= layer0_outputs(9613);
    outputs(9364) <= (layer0_outputs(3616)) xor (layer0_outputs(3727));
    outputs(9365) <= not((layer0_outputs(9646)) xor (layer0_outputs(186)));
    outputs(9366) <= (layer0_outputs(6018)) xor (layer0_outputs(3249));
    outputs(9367) <= not(layer0_outputs(5858));
    outputs(9368) <= (layer0_outputs(356)) xor (layer0_outputs(5593));
    outputs(9369) <= not((layer0_outputs(9056)) or (layer0_outputs(6499)));
    outputs(9370) <= not((layer0_outputs(3952)) xor (layer0_outputs(3127)));
    outputs(9371) <= not(layer0_outputs(3557)) or (layer0_outputs(5387));
    outputs(9372) <= (layer0_outputs(8972)) xor (layer0_outputs(8636));
    outputs(9373) <= layer0_outputs(2512);
    outputs(9374) <= not(layer0_outputs(8585));
    outputs(9375) <= (layer0_outputs(5762)) xor (layer0_outputs(9517));
    outputs(9376) <= (layer0_outputs(9018)) and not (layer0_outputs(6539));
    outputs(9377) <= layer0_outputs(2431);
    outputs(9378) <= not(layer0_outputs(3504));
    outputs(9379) <= layer0_outputs(2602);
    outputs(9380) <= not(layer0_outputs(1244));
    outputs(9381) <= not(layer0_outputs(6386));
    outputs(9382) <= not(layer0_outputs(9026));
    outputs(9383) <= (layer0_outputs(8738)) or (layer0_outputs(6810));
    outputs(9384) <= (layer0_outputs(8435)) xor (layer0_outputs(2183));
    outputs(9385) <= layer0_outputs(1894);
    outputs(9386) <= not((layer0_outputs(790)) or (layer0_outputs(2496)));
    outputs(9387) <= not(layer0_outputs(1867));
    outputs(9388) <= (layer0_outputs(3957)) and not (layer0_outputs(9698));
    outputs(9389) <= not(layer0_outputs(1184)) or (layer0_outputs(6173));
    outputs(9390) <= (layer0_outputs(2372)) xor (layer0_outputs(434));
    outputs(9391) <= not(layer0_outputs(6329));
    outputs(9392) <= not(layer0_outputs(3308));
    outputs(9393) <= not((layer0_outputs(4110)) xor (layer0_outputs(9503)));
    outputs(9394) <= not((layer0_outputs(1624)) xor (layer0_outputs(9531)));
    outputs(9395) <= (layer0_outputs(1200)) and not (layer0_outputs(8266));
    outputs(9396) <= not(layer0_outputs(8390)) or (layer0_outputs(831));
    outputs(9397) <= layer0_outputs(3507);
    outputs(9398) <= layer0_outputs(305);
    outputs(9399) <= not((layer0_outputs(4084)) xor (layer0_outputs(1982)));
    outputs(9400) <= layer0_outputs(1870);
    outputs(9401) <= layer0_outputs(8772);
    outputs(9402) <= layer0_outputs(5744);
    outputs(9403) <= (layer0_outputs(6937)) xor (layer0_outputs(1995));
    outputs(9404) <= not(layer0_outputs(9346));
    outputs(9405) <= (layer0_outputs(8031)) xor (layer0_outputs(7400));
    outputs(9406) <= layer0_outputs(2492);
    outputs(9407) <= not(layer0_outputs(4520)) or (layer0_outputs(10006));
    outputs(9408) <= (layer0_outputs(8758)) or (layer0_outputs(4496));
    outputs(9409) <= not(layer0_outputs(9301));
    outputs(9410) <= layer0_outputs(9692);
    outputs(9411) <= layer0_outputs(3396);
    outputs(9412) <= not((layer0_outputs(397)) or (layer0_outputs(1549)));
    outputs(9413) <= (layer0_outputs(5498)) xor (layer0_outputs(2848));
    outputs(9414) <= layer0_outputs(3941);
    outputs(9415) <= not((layer0_outputs(5201)) or (layer0_outputs(8516)));
    outputs(9416) <= not(layer0_outputs(2047));
    outputs(9417) <= (layer0_outputs(5184)) and not (layer0_outputs(2189));
    outputs(9418) <= (layer0_outputs(486)) and (layer0_outputs(5745));
    outputs(9419) <= not(layer0_outputs(2628));
    outputs(9420) <= not((layer0_outputs(4516)) xor (layer0_outputs(9059)));
    outputs(9421) <= not((layer0_outputs(5302)) xor (layer0_outputs(8765)));
    outputs(9422) <= layer0_outputs(280);
    outputs(9423) <= (layer0_outputs(3562)) and not (layer0_outputs(8));
    outputs(9424) <= not(layer0_outputs(4822));
    outputs(9425) <= not(layer0_outputs(329));
    outputs(9426) <= layer0_outputs(2942);
    outputs(9427) <= not(layer0_outputs(1440));
    outputs(9428) <= not(layer0_outputs(5730));
    outputs(9429) <= (layer0_outputs(6214)) or (layer0_outputs(2557));
    outputs(9430) <= (layer0_outputs(3181)) and not (layer0_outputs(2177));
    outputs(9431) <= not((layer0_outputs(7564)) xor (layer0_outputs(2704)));
    outputs(9432) <= (layer0_outputs(10021)) xor (layer0_outputs(9917));
    outputs(9433) <= not(layer0_outputs(8941));
    outputs(9434) <= (layer0_outputs(5413)) and not (layer0_outputs(3004));
    outputs(9435) <= layer0_outputs(7715);
    outputs(9436) <= (layer0_outputs(2312)) xor (layer0_outputs(7663));
    outputs(9437) <= (layer0_outputs(4877)) and not (layer0_outputs(3723));
    outputs(9438) <= not(layer0_outputs(388));
    outputs(9439) <= layer0_outputs(8712);
    outputs(9440) <= not(layer0_outputs(5593)) or (layer0_outputs(1381));
    outputs(9441) <= layer0_outputs(3585);
    outputs(9442) <= not((layer0_outputs(4891)) xor (layer0_outputs(5552)));
    outputs(9443) <= (layer0_outputs(4477)) xor (layer0_outputs(8930));
    outputs(9444) <= (layer0_outputs(5457)) xor (layer0_outputs(1131));
    outputs(9445) <= not(layer0_outputs(2107));
    outputs(9446) <= layer0_outputs(8850);
    outputs(9447) <= (layer0_outputs(9978)) and not (layer0_outputs(1050));
    outputs(9448) <= not((layer0_outputs(9165)) xor (layer0_outputs(9933)));
    outputs(9449) <= layer0_outputs(5876);
    outputs(9450) <= '0';
    outputs(9451) <= not((layer0_outputs(4644)) xor (layer0_outputs(3758)));
    outputs(9452) <= layer0_outputs(5262);
    outputs(9453) <= (layer0_outputs(6250)) xor (layer0_outputs(9695));
    outputs(9454) <= (layer0_outputs(9967)) and not (layer0_outputs(6246));
    outputs(9455) <= (layer0_outputs(2123)) and (layer0_outputs(5291));
    outputs(9456) <= layer0_outputs(4629);
    outputs(9457) <= not(layer0_outputs(7787)) or (layer0_outputs(281));
    outputs(9458) <= not(layer0_outputs(6457)) or (layer0_outputs(6710));
    outputs(9459) <= (layer0_outputs(3106)) and not (layer0_outputs(8896));
    outputs(9460) <= (layer0_outputs(6469)) xor (layer0_outputs(9446));
    outputs(9461) <= not(layer0_outputs(842));
    outputs(9462) <= (layer0_outputs(1032)) xor (layer0_outputs(5924));
    outputs(9463) <= layer0_outputs(7019);
    outputs(9464) <= layer0_outputs(5128);
    outputs(9465) <= layer0_outputs(320);
    outputs(9466) <= not(layer0_outputs(9694));
    outputs(9467) <= not((layer0_outputs(9539)) xor (layer0_outputs(5028)));
    outputs(9468) <= not(layer0_outputs(1181));
    outputs(9469) <= (layer0_outputs(9773)) or (layer0_outputs(962));
    outputs(9470) <= not(layer0_outputs(3076));
    outputs(9471) <= not(layer0_outputs(9110)) or (layer0_outputs(8460));
    outputs(9472) <= (layer0_outputs(9178)) xor (layer0_outputs(5964));
    outputs(9473) <= not(layer0_outputs(5632));
    outputs(9474) <= layer0_outputs(3821);
    outputs(9475) <= (layer0_outputs(3044)) and not (layer0_outputs(8375));
    outputs(9476) <= not(layer0_outputs(5372));
    outputs(9477) <= (layer0_outputs(1373)) xor (layer0_outputs(2870));
    outputs(9478) <= (layer0_outputs(1778)) xor (layer0_outputs(6287));
    outputs(9479) <= not((layer0_outputs(5693)) xor (layer0_outputs(7518)));
    outputs(9480) <= (layer0_outputs(7672)) and not (layer0_outputs(7674));
    outputs(9481) <= not((layer0_outputs(9789)) xor (layer0_outputs(6119)));
    outputs(9482) <= (layer0_outputs(71)) and (layer0_outputs(8960));
    outputs(9483) <= (layer0_outputs(9944)) and not (layer0_outputs(10033));
    outputs(9484) <= (layer0_outputs(7662)) xor (layer0_outputs(7494));
    outputs(9485) <= not((layer0_outputs(1657)) or (layer0_outputs(4620)));
    outputs(9486) <= not(layer0_outputs(5880));
    outputs(9487) <= not(layer0_outputs(4038));
    outputs(9488) <= not(layer0_outputs(1170));
    outputs(9489) <= layer0_outputs(830);
    outputs(9490) <= not(layer0_outputs(8838));
    outputs(9491) <= (layer0_outputs(6943)) and not (layer0_outputs(2073));
    outputs(9492) <= (layer0_outputs(1425)) xor (layer0_outputs(6072));
    outputs(9493) <= (layer0_outputs(5586)) and not (layer0_outputs(3453));
    outputs(9494) <= (layer0_outputs(8022)) and not (layer0_outputs(8612));
    outputs(9495) <= not(layer0_outputs(2818));
    outputs(9496) <= not(layer0_outputs(591));
    outputs(9497) <= not((layer0_outputs(2008)) xor (layer0_outputs(8594)));
    outputs(9498) <= (layer0_outputs(2640)) and not (layer0_outputs(2552));
    outputs(9499) <= not(layer0_outputs(8158)) or (layer0_outputs(10051));
    outputs(9500) <= layer0_outputs(705);
    outputs(9501) <= (layer0_outputs(7638)) xor (layer0_outputs(4996));
    outputs(9502) <= not(layer0_outputs(1378));
    outputs(9503) <= (layer0_outputs(8777)) and (layer0_outputs(1996));
    outputs(9504) <= not((layer0_outputs(494)) xor (layer0_outputs(7792)));
    outputs(9505) <= (layer0_outputs(4810)) xor (layer0_outputs(8496));
    outputs(9506) <= not(layer0_outputs(3108));
    outputs(9507) <= not(layer0_outputs(5444)) or (layer0_outputs(7282));
    outputs(9508) <= not((layer0_outputs(2725)) and (layer0_outputs(6756)));
    outputs(9509) <= (layer0_outputs(476)) xor (layer0_outputs(8495));
    outputs(9510) <= not((layer0_outputs(480)) xor (layer0_outputs(131)));
    outputs(9511) <= not((layer0_outputs(6427)) xor (layer0_outputs(4720)));
    outputs(9512) <= not(layer0_outputs(2468)) or (layer0_outputs(9845));
    outputs(9513) <= (layer0_outputs(8823)) and not (layer0_outputs(6805));
    outputs(9514) <= (layer0_outputs(3097)) xor (layer0_outputs(5784));
    outputs(9515) <= layer0_outputs(3398);
    outputs(9516) <= not(layer0_outputs(893));
    outputs(9517) <= not((layer0_outputs(5241)) or (layer0_outputs(6426)));
    outputs(9518) <= (layer0_outputs(7754)) and (layer0_outputs(9298));
    outputs(9519) <= not((layer0_outputs(7108)) or (layer0_outputs(3264)));
    outputs(9520) <= (layer0_outputs(4156)) and (layer0_outputs(4845));
    outputs(9521) <= not(layer0_outputs(8136));
    outputs(9522) <= layer0_outputs(4000);
    outputs(9523) <= not(layer0_outputs(3620));
    outputs(9524) <= (layer0_outputs(1893)) and not (layer0_outputs(1967));
    outputs(9525) <= not((layer0_outputs(6671)) xor (layer0_outputs(4881)));
    outputs(9526) <= not(layer0_outputs(3238));
    outputs(9527) <= not((layer0_outputs(3313)) xor (layer0_outputs(7802)));
    outputs(9528) <= (layer0_outputs(2896)) or (layer0_outputs(9594));
    outputs(9529) <= (layer0_outputs(7949)) xor (layer0_outputs(1061));
    outputs(9530) <= layer0_outputs(1843);
    outputs(9531) <= layer0_outputs(6205);
    outputs(9532) <= (layer0_outputs(2046)) and not (layer0_outputs(1512));
    outputs(9533) <= (layer0_outputs(4433)) and not (layer0_outputs(7659));
    outputs(9534) <= not(layer0_outputs(3030));
    outputs(9535) <= '0';
    outputs(9536) <= layer0_outputs(9453);
    outputs(9537) <= (layer0_outputs(2332)) xor (layer0_outputs(150));
    outputs(9538) <= layer0_outputs(542);
    outputs(9539) <= (layer0_outputs(61)) and not (layer0_outputs(503));
    outputs(9540) <= not(layer0_outputs(3626));
    outputs(9541) <= (layer0_outputs(9171)) and (layer0_outputs(1929));
    outputs(9542) <= not(layer0_outputs(1673));
    outputs(9543) <= layer0_outputs(1411);
    outputs(9544) <= not((layer0_outputs(3023)) xor (layer0_outputs(7045)));
    outputs(9545) <= (layer0_outputs(4591)) or (layer0_outputs(5526));
    outputs(9546) <= layer0_outputs(3706);
    outputs(9547) <= not(layer0_outputs(5032));
    outputs(9548) <= layer0_outputs(636);
    outputs(9549) <= (layer0_outputs(4883)) and not (layer0_outputs(9857));
    outputs(9550) <= not((layer0_outputs(6988)) xor (layer0_outputs(3971)));
    outputs(9551) <= (layer0_outputs(2874)) and not (layer0_outputs(1366));
    outputs(9552) <= not((layer0_outputs(8880)) and (layer0_outputs(1441)));
    outputs(9553) <= (layer0_outputs(3435)) xor (layer0_outputs(2868));
    outputs(9554) <= not(layer0_outputs(7086));
    outputs(9555) <= not(layer0_outputs(9547));
    outputs(9556) <= layer0_outputs(3375);
    outputs(9557) <= not((layer0_outputs(6866)) xor (layer0_outputs(5640)));
    outputs(9558) <= layer0_outputs(8088);
    outputs(9559) <= not((layer0_outputs(1232)) xor (layer0_outputs(5914)));
    outputs(9560) <= layer0_outputs(547);
    outputs(9561) <= not(layer0_outputs(9258));
    outputs(9562) <= (layer0_outputs(7309)) and not (layer0_outputs(1145));
    outputs(9563) <= (layer0_outputs(3265)) and (layer0_outputs(1856));
    outputs(9564) <= layer0_outputs(370);
    outputs(9565) <= (layer0_outputs(2547)) xor (layer0_outputs(4938));
    outputs(9566) <= not(layer0_outputs(10093));
    outputs(9567) <= layer0_outputs(9883);
    outputs(9568) <= (layer0_outputs(3103)) and not (layer0_outputs(5512));
    outputs(9569) <= (layer0_outputs(8977)) xor (layer0_outputs(2032));
    outputs(9570) <= layer0_outputs(2288);
    outputs(9571) <= (layer0_outputs(2135)) and not (layer0_outputs(9071));
    outputs(9572) <= layer0_outputs(5992);
    outputs(9573) <= not(layer0_outputs(6718));
    outputs(9574) <= layer0_outputs(8242);
    outputs(9575) <= not(layer0_outputs(5324));
    outputs(9576) <= (layer0_outputs(8416)) or (layer0_outputs(4082));
    outputs(9577) <= (layer0_outputs(3326)) and not (layer0_outputs(5627));
    outputs(9578) <= not((layer0_outputs(8265)) xor (layer0_outputs(7401)));
    outputs(9579) <= (layer0_outputs(7502)) and not (layer0_outputs(7655));
    outputs(9580) <= not((layer0_outputs(129)) and (layer0_outputs(6225)));
    outputs(9581) <= (layer0_outputs(2831)) xor (layer0_outputs(3333));
    outputs(9582) <= (layer0_outputs(4551)) or (layer0_outputs(949));
    outputs(9583) <= (layer0_outputs(8525)) and (layer0_outputs(3563));
    outputs(9584) <= (layer0_outputs(4379)) xor (layer0_outputs(10189));
    outputs(9585) <= (layer0_outputs(5992)) and not (layer0_outputs(4925));
    outputs(9586) <= layer0_outputs(8023);
    outputs(9587) <= not(layer0_outputs(8466));
    outputs(9588) <= not((layer0_outputs(2220)) or (layer0_outputs(9511)));
    outputs(9589) <= (layer0_outputs(1507)) and not (layer0_outputs(380));
    outputs(9590) <= not(layer0_outputs(1522));
    outputs(9591) <= (layer0_outputs(2249)) xor (layer0_outputs(7573));
    outputs(9592) <= not(layer0_outputs(10045)) or (layer0_outputs(1991));
    outputs(9593) <= not(layer0_outputs(3328));
    outputs(9594) <= layer0_outputs(6130);
    outputs(9595) <= not(layer0_outputs(5472));
    outputs(9596) <= (layer0_outputs(5211)) or (layer0_outputs(869));
    outputs(9597) <= not((layer0_outputs(5906)) xor (layer0_outputs(7854)));
    outputs(9598) <= layer0_outputs(4621);
    outputs(9599) <= layer0_outputs(3083);
    outputs(9600) <= layer0_outputs(7523);
    outputs(9601) <= (layer0_outputs(1393)) and not (layer0_outputs(5009));
    outputs(9602) <= not(layer0_outputs(5323));
    outputs(9603) <= not((layer0_outputs(6203)) xor (layer0_outputs(1550)));
    outputs(9604) <= (layer0_outputs(2488)) and not (layer0_outputs(6835));
    outputs(9605) <= not((layer0_outputs(2808)) xor (layer0_outputs(5287)));
    outputs(9606) <= (layer0_outputs(9006)) and not (layer0_outputs(7279));
    outputs(9607) <= not(layer0_outputs(8775));
    outputs(9608) <= layer0_outputs(8442);
    outputs(9609) <= not(layer0_outputs(6423));
    outputs(9610) <= (layer0_outputs(3645)) xor (layer0_outputs(196));
    outputs(9611) <= not(layer0_outputs(3470)) or (layer0_outputs(62));
    outputs(9612) <= layer0_outputs(4243);
    outputs(9613) <= layer0_outputs(7353);
    outputs(9614) <= (layer0_outputs(1815)) and not (layer0_outputs(32));
    outputs(9615) <= not(layer0_outputs(2174));
    outputs(9616) <= layer0_outputs(2452);
    outputs(9617) <= layer0_outputs(8738);
    outputs(9618) <= (layer0_outputs(3122)) xor (layer0_outputs(9840));
    outputs(9619) <= not((layer0_outputs(8031)) or (layer0_outputs(968)));
    outputs(9620) <= not((layer0_outputs(3685)) xor (layer0_outputs(5790)));
    outputs(9621) <= (layer0_outputs(2159)) and (layer0_outputs(9981));
    outputs(9622) <= (layer0_outputs(4146)) or (layer0_outputs(421));
    outputs(9623) <= not((layer0_outputs(9614)) xor (layer0_outputs(2330)));
    outputs(9624) <= not((layer0_outputs(7134)) or (layer0_outputs(863)));
    outputs(9625) <= not((layer0_outputs(4755)) or (layer0_outputs(4944)));
    outputs(9626) <= not((layer0_outputs(8478)) xor (layer0_outputs(9681)));
    outputs(9627) <= (layer0_outputs(5389)) xor (layer0_outputs(6239));
    outputs(9628) <= not((layer0_outputs(1493)) xor (layer0_outputs(8979)));
    outputs(9629) <= not(layer0_outputs(658));
    outputs(9630) <= layer0_outputs(2900);
    outputs(9631) <= layer0_outputs(6534);
    outputs(9632) <= not(layer0_outputs(8793));
    outputs(9633) <= not((layer0_outputs(1128)) and (layer0_outputs(9040)));
    outputs(9634) <= not((layer0_outputs(4297)) or (layer0_outputs(7835)));
    outputs(9635) <= not((layer0_outputs(3612)) xor (layer0_outputs(1188)));
    outputs(9636) <= layer0_outputs(5692);
    outputs(9637) <= (layer0_outputs(5397)) and not (layer0_outputs(107));
    outputs(9638) <= (layer0_outputs(3172)) xor (layer0_outputs(726));
    outputs(9639) <= (layer0_outputs(761)) or (layer0_outputs(6955));
    outputs(9640) <= layer0_outputs(9224);
    outputs(9641) <= (layer0_outputs(9921)) xor (layer0_outputs(1911));
    outputs(9642) <= layer0_outputs(862);
    outputs(9643) <= not((layer0_outputs(2237)) or (layer0_outputs(6299)));
    outputs(9644) <= (layer0_outputs(7635)) and (layer0_outputs(5178));
    outputs(9645) <= layer0_outputs(6269);
    outputs(9646) <= (layer0_outputs(5873)) and (layer0_outputs(1895));
    outputs(9647) <= not((layer0_outputs(2979)) or (layer0_outputs(3162)));
    outputs(9648) <= (layer0_outputs(1572)) and not (layer0_outputs(9240));
    outputs(9649) <= not(layer0_outputs(6847));
    outputs(9650) <= not((layer0_outputs(4939)) xor (layer0_outputs(2379)));
    outputs(9651) <= not(layer0_outputs(2121));
    outputs(9652) <= layer0_outputs(2616);
    outputs(9653) <= not(layer0_outputs(2955));
    outputs(9654) <= not(layer0_outputs(2052));
    outputs(9655) <= (layer0_outputs(6503)) and not (layer0_outputs(4354));
    outputs(9656) <= not((layer0_outputs(7832)) and (layer0_outputs(4439)));
    outputs(9657) <= layer0_outputs(7949);
    outputs(9658) <= (layer0_outputs(5662)) and not (layer0_outputs(3911));
    outputs(9659) <= (layer0_outputs(2381)) xor (layer0_outputs(34));
    outputs(9660) <= (layer0_outputs(8355)) and not (layer0_outputs(5762));
    outputs(9661) <= (layer0_outputs(4497)) and (layer0_outputs(9347));
    outputs(9662) <= not((layer0_outputs(9949)) xor (layer0_outputs(1695)));
    outputs(9663) <= not((layer0_outputs(9838)) xor (layer0_outputs(1582)));
    outputs(9664) <= (layer0_outputs(4453)) and (layer0_outputs(8635));
    outputs(9665) <= not(layer0_outputs(6387));
    outputs(9666) <= not(layer0_outputs(739));
    outputs(9667) <= (layer0_outputs(7680)) and not (layer0_outputs(211));
    outputs(9668) <= layer0_outputs(6939);
    outputs(9669) <= not(layer0_outputs(916));
    outputs(9670) <= layer0_outputs(5567);
    outputs(9671) <= layer0_outputs(1606);
    outputs(9672) <= (layer0_outputs(8470)) xor (layer0_outputs(45));
    outputs(9673) <= layer0_outputs(6356);
    outputs(9674) <= layer0_outputs(70);
    outputs(9675) <= not((layer0_outputs(7935)) xor (layer0_outputs(6973)));
    outputs(9676) <= (layer0_outputs(4828)) xor (layer0_outputs(1762));
    outputs(9677) <= layer0_outputs(7757);
    outputs(9678) <= layer0_outputs(1926);
    outputs(9679) <= (layer0_outputs(1231)) and not (layer0_outputs(8894));
    outputs(9680) <= (layer0_outputs(8379)) and (layer0_outputs(5379));
    outputs(9681) <= not(layer0_outputs(5561));
    outputs(9682) <= not((layer0_outputs(8471)) xor (layer0_outputs(2339)));
    outputs(9683) <= (layer0_outputs(1720)) or (layer0_outputs(8906));
    outputs(9684) <= not(layer0_outputs(6499));
    outputs(9685) <= not((layer0_outputs(2507)) or (layer0_outputs(7341)));
    outputs(9686) <= (layer0_outputs(4644)) xor (layer0_outputs(4694));
    outputs(9687) <= not(layer0_outputs(2036));
    outputs(9688) <= not(layer0_outputs(9044));
    outputs(9689) <= not((layer0_outputs(6320)) and (layer0_outputs(7437)));
    outputs(9690) <= not(layer0_outputs(6862));
    outputs(9691) <= not((layer0_outputs(3081)) and (layer0_outputs(7867)));
    outputs(9692) <= not((layer0_outputs(587)) xor (layer0_outputs(3217)));
    outputs(9693) <= not((layer0_outputs(5537)) or (layer0_outputs(3642)));
    outputs(9694) <= (layer0_outputs(1576)) and not (layer0_outputs(9447));
    outputs(9695) <= (layer0_outputs(7710)) and not (layer0_outputs(2743));
    outputs(9696) <= layer0_outputs(4885);
    outputs(9697) <= (layer0_outputs(4077)) and (layer0_outputs(8011));
    outputs(9698) <= not(layer0_outputs(1837));
    outputs(9699) <= '1';
    outputs(9700) <= layer0_outputs(1849);
    outputs(9701) <= (layer0_outputs(4386)) or (layer0_outputs(9704));
    outputs(9702) <= layer0_outputs(1258);
    outputs(9703) <= not(layer0_outputs(6289));
    outputs(9704) <= (layer0_outputs(2442)) and (layer0_outputs(1274));
    outputs(9705) <= not(layer0_outputs(7863));
    outputs(9706) <= not(layer0_outputs(1652));
    outputs(9707) <= not(layer0_outputs(4617));
    outputs(9708) <= not(layer0_outputs(4800));
    outputs(9709) <= not(layer0_outputs(9299)) or (layer0_outputs(5584));
    outputs(9710) <= not((layer0_outputs(4589)) and (layer0_outputs(5357)));
    outputs(9711) <= (layer0_outputs(450)) or (layer0_outputs(6097));
    outputs(9712) <= not((layer0_outputs(9232)) xor (layer0_outputs(5800)));
    outputs(9713) <= layer0_outputs(432);
    outputs(9714) <= (layer0_outputs(9915)) xor (layer0_outputs(1223));
    outputs(9715) <= layer0_outputs(10137);
    outputs(9716) <= (layer0_outputs(5060)) xor (layer0_outputs(674));
    outputs(9717) <= not(layer0_outputs(918)) or (layer0_outputs(7731));
    outputs(9718) <= not(layer0_outputs(3498));
    outputs(9719) <= (layer0_outputs(4553)) and not (layer0_outputs(2633));
    outputs(9720) <= not(layer0_outputs(1304));
    outputs(9721) <= (layer0_outputs(6869)) and (layer0_outputs(4422));
    outputs(9722) <= (layer0_outputs(5843)) xor (layer0_outputs(8195));
    outputs(9723) <= layer0_outputs(7203);
    outputs(9724) <= (layer0_outputs(7299)) xor (layer0_outputs(2622));
    outputs(9725) <= not(layer0_outputs(6938));
    outputs(9726) <= (layer0_outputs(2778)) and not (layer0_outputs(2006));
    outputs(9727) <= (layer0_outputs(8597)) xor (layer0_outputs(5706));
    outputs(9728) <= not(layer0_outputs(8790));
    outputs(9729) <= (layer0_outputs(6679)) and (layer0_outputs(4605));
    outputs(9730) <= layer0_outputs(1687);
    outputs(9731) <= (layer0_outputs(2812)) and (layer0_outputs(829));
    outputs(9732) <= (layer0_outputs(5261)) xor (layer0_outputs(4726));
    outputs(9733) <= layer0_outputs(7106);
    outputs(9734) <= (layer0_outputs(6568)) xor (layer0_outputs(9141));
    outputs(9735) <= (layer0_outputs(2808)) xor (layer0_outputs(4749));
    outputs(9736) <= (layer0_outputs(3271)) xor (layer0_outputs(219));
    outputs(9737) <= layer0_outputs(6194);
    outputs(9738) <= (layer0_outputs(6099)) or (layer0_outputs(5611));
    outputs(9739) <= layer0_outputs(4543);
    outputs(9740) <= not((layer0_outputs(2643)) xor (layer0_outputs(3882)));
    outputs(9741) <= (layer0_outputs(10020)) xor (layer0_outputs(9339));
    outputs(9742) <= (layer0_outputs(6266)) xor (layer0_outputs(4780));
    outputs(9743) <= '0';
    outputs(9744) <= layer0_outputs(222);
    outputs(9745) <= not(layer0_outputs(3408));
    outputs(9746) <= not(layer0_outputs(7221));
    outputs(9747) <= (layer0_outputs(7130)) xor (layer0_outputs(8443));
    outputs(9748) <= (layer0_outputs(3930)) xor (layer0_outputs(9955));
    outputs(9749) <= (layer0_outputs(8175)) xor (layer0_outputs(387));
    outputs(9750) <= (layer0_outputs(2473)) xor (layer0_outputs(1089));
    outputs(9751) <= not((layer0_outputs(8593)) or (layer0_outputs(1207)));
    outputs(9752) <= layer0_outputs(1360);
    outputs(9753) <= (layer0_outputs(4957)) and (layer0_outputs(1708));
    outputs(9754) <= (layer0_outputs(1964)) xor (layer0_outputs(5121));
    outputs(9755) <= not((layer0_outputs(2871)) or (layer0_outputs(2594)));
    outputs(9756) <= layer0_outputs(4028);
    outputs(9757) <= layer0_outputs(8730);
    outputs(9758) <= (layer0_outputs(7180)) xor (layer0_outputs(4905));
    outputs(9759) <= (layer0_outputs(7661)) and not (layer0_outputs(4966));
    outputs(9760) <= (layer0_outputs(2544)) and (layer0_outputs(9779));
    outputs(9761) <= not((layer0_outputs(2902)) xor (layer0_outputs(7389)));
    outputs(9762) <= (layer0_outputs(490)) and not (layer0_outputs(4545));
    outputs(9763) <= not(layer0_outputs(5316));
    outputs(9764) <= not((layer0_outputs(9014)) xor (layer0_outputs(6807)));
    outputs(9765) <= not((layer0_outputs(2968)) xor (layer0_outputs(1434)));
    outputs(9766) <= not(layer0_outputs(4879)) or (layer0_outputs(635));
    outputs(9767) <= (layer0_outputs(4595)) and not (layer0_outputs(5423));
    outputs(9768) <= (layer0_outputs(5936)) or (layer0_outputs(295));
    outputs(9769) <= (layer0_outputs(10210)) xor (layer0_outputs(829));
    outputs(9770) <= not(layer0_outputs(3436));
    outputs(9771) <= layer0_outputs(5549);
    outputs(9772) <= not(layer0_outputs(976));
    outputs(9773) <= not(layer0_outputs(7218));
    outputs(9774) <= not(layer0_outputs(1736)) or (layer0_outputs(6949));
    outputs(9775) <= (layer0_outputs(3113)) xor (layer0_outputs(8304));
    outputs(9776) <= not(layer0_outputs(5758));
    outputs(9777) <= not((layer0_outputs(1305)) or (layer0_outputs(260)));
    outputs(9778) <= (layer0_outputs(6442)) xor (layer0_outputs(1646));
    outputs(9779) <= (layer0_outputs(1634)) xor (layer0_outputs(3373));
    outputs(9780) <= not((layer0_outputs(7639)) xor (layer0_outputs(1058)));
    outputs(9781) <= (layer0_outputs(7501)) and not (layer0_outputs(5149));
    outputs(9782) <= layer0_outputs(5496);
    outputs(9783) <= not(layer0_outputs(8513));
    outputs(9784) <= layer0_outputs(7288);
    outputs(9785) <= (layer0_outputs(6694)) xor (layer0_outputs(55));
    outputs(9786) <= (layer0_outputs(664)) or (layer0_outputs(9834));
    outputs(9787) <= (layer0_outputs(8915)) and not (layer0_outputs(646));
    outputs(9788) <= layer0_outputs(2397);
    outputs(9789) <= not(layer0_outputs(617)) or (layer0_outputs(7751));
    outputs(9790) <= (layer0_outputs(7180)) xor (layer0_outputs(9012));
    outputs(9791) <= (layer0_outputs(3327)) xor (layer0_outputs(8406));
    outputs(9792) <= not((layer0_outputs(6559)) and (layer0_outputs(10006)));
    outputs(9793) <= not(layer0_outputs(3536)) or (layer0_outputs(7213));
    outputs(9794) <= (layer0_outputs(10218)) xor (layer0_outputs(9007));
    outputs(9795) <= not(layer0_outputs(644));
    outputs(9796) <= not(layer0_outputs(3126));
    outputs(9797) <= (layer0_outputs(4902)) and (layer0_outputs(8037));
    outputs(9798) <= layer0_outputs(8892);
    outputs(9799) <= layer0_outputs(659);
    outputs(9800) <= (layer0_outputs(6908)) xor (layer0_outputs(4359));
    outputs(9801) <= (layer0_outputs(6581)) xor (layer0_outputs(8439));
    outputs(9802) <= not((layer0_outputs(28)) or (layer0_outputs(278)));
    outputs(9803) <= layer0_outputs(2649);
    outputs(9804) <= layer0_outputs(7140);
    outputs(9805) <= not(layer0_outputs(8611));
    outputs(9806) <= (layer0_outputs(4596)) and not (layer0_outputs(9271));
    outputs(9807) <= not(layer0_outputs(8181));
    outputs(9808) <= not((layer0_outputs(3359)) xor (layer0_outputs(266)));
    outputs(9809) <= not((layer0_outputs(118)) xor (layer0_outputs(7858)));
    outputs(9810) <= not((layer0_outputs(5671)) xor (layer0_outputs(1618)));
    outputs(9811) <= not((layer0_outputs(6722)) xor (layer0_outputs(2606)));
    outputs(9812) <= (layer0_outputs(6220)) and (layer0_outputs(4649));
    outputs(9813) <= not((layer0_outputs(7311)) xor (layer0_outputs(1778)));
    outputs(9814) <= (layer0_outputs(7860)) xor (layer0_outputs(7513));
    outputs(9815) <= not(layer0_outputs(2090)) or (layer0_outputs(1445));
    outputs(9816) <= (layer0_outputs(1156)) xor (layer0_outputs(4813));
    outputs(9817) <= (layer0_outputs(7716)) xor (layer0_outputs(4233));
    outputs(9818) <= not((layer0_outputs(2787)) xor (layer0_outputs(1689)));
    outputs(9819) <= not(layer0_outputs(5242));
    outputs(9820) <= not(layer0_outputs(4512));
    outputs(9821) <= not((layer0_outputs(8605)) xor (layer0_outputs(434)));
    outputs(9822) <= layer0_outputs(3397);
    outputs(9823) <= (layer0_outputs(4764)) and (layer0_outputs(7984));
    outputs(9824) <= (layer0_outputs(6247)) and not (layer0_outputs(7693));
    outputs(9825) <= not(layer0_outputs(3133));
    outputs(9826) <= layer0_outputs(7);
    outputs(9827) <= not((layer0_outputs(1162)) and (layer0_outputs(8215)));
    outputs(9828) <= (layer0_outputs(764)) and not (layer0_outputs(4821));
    outputs(9829) <= not((layer0_outputs(1402)) xor (layer0_outputs(2687)));
    outputs(9830) <= not(layer0_outputs(8974));
    outputs(9831) <= (layer0_outputs(8709)) and (layer0_outputs(7027));
    outputs(9832) <= layer0_outputs(2202);
    outputs(9833) <= not((layer0_outputs(7654)) or (layer0_outputs(6116)));
    outputs(9834) <= (layer0_outputs(7670)) and not (layer0_outputs(8781));
    outputs(9835) <= layer0_outputs(9422);
    outputs(9836) <= layer0_outputs(2776);
    outputs(9837) <= layer0_outputs(8403);
    outputs(9838) <= not((layer0_outputs(2638)) or (layer0_outputs(3872)));
    outputs(9839) <= not(layer0_outputs(1226));
    outputs(9840) <= not((layer0_outputs(3593)) or (layer0_outputs(6627)));
    outputs(9841) <= not((layer0_outputs(5361)) or (layer0_outputs(38)));
    outputs(9842) <= not((layer0_outputs(993)) or (layer0_outputs(637)));
    outputs(9843) <= not(layer0_outputs(4989));
    outputs(9844) <= (layer0_outputs(1047)) and (layer0_outputs(1766));
    outputs(9845) <= (layer0_outputs(7081)) xor (layer0_outputs(4141));
    outputs(9846) <= not(layer0_outputs(1883)) or (layer0_outputs(6075));
    outputs(9847) <= (layer0_outputs(7493)) and not (layer0_outputs(4573));
    outputs(9848) <= not(layer0_outputs(1464));
    outputs(9849) <= not(layer0_outputs(8881));
    outputs(9850) <= not((layer0_outputs(5042)) xor (layer0_outputs(3344)));
    outputs(9851) <= not(layer0_outputs(4157));
    outputs(9852) <= (layer0_outputs(3948)) and (layer0_outputs(3464));
    outputs(9853) <= not(layer0_outputs(7229));
    outputs(9854) <= not(layer0_outputs(6153));
    outputs(9855) <= not((layer0_outputs(7383)) xor (layer0_outputs(7992)));
    outputs(9856) <= not(layer0_outputs(93));
    outputs(9857) <= layer0_outputs(8617);
    outputs(9858) <= layer0_outputs(2365);
    outputs(9859) <= not(layer0_outputs(1520));
    outputs(9860) <= not(layer0_outputs(4531)) or (layer0_outputs(5193));
    outputs(9861) <= (layer0_outputs(3624)) and not (layer0_outputs(2157));
    outputs(9862) <= layer0_outputs(2784);
    outputs(9863) <= not(layer0_outputs(8622));
    outputs(9864) <= layer0_outputs(413);
    outputs(9865) <= layer0_outputs(2129);
    outputs(9866) <= not(layer0_outputs(3156));
    outputs(9867) <= (layer0_outputs(3714)) xor (layer0_outputs(1197));
    outputs(9868) <= (layer0_outputs(7696)) and not (layer0_outputs(3361));
    outputs(9869) <= not((layer0_outputs(6343)) xor (layer0_outputs(5091)));
    outputs(9870) <= layer0_outputs(744);
    outputs(9871) <= not(layer0_outputs(4711));
    outputs(9872) <= (layer0_outputs(4464)) or (layer0_outputs(485));
    outputs(9873) <= not((layer0_outputs(8914)) or (layer0_outputs(6184)));
    outputs(9874) <= not(layer0_outputs(3112));
    outputs(9875) <= not((layer0_outputs(8169)) xor (layer0_outputs(354)));
    outputs(9876) <= layer0_outputs(3257);
    outputs(9877) <= (layer0_outputs(2924)) and not (layer0_outputs(8721));
    outputs(9878) <= (layer0_outputs(7177)) and (layer0_outputs(8417));
    outputs(9879) <= not((layer0_outputs(4424)) xor (layer0_outputs(3362)));
    outputs(9880) <= not((layer0_outputs(5782)) or (layer0_outputs(2414)));
    outputs(9881) <= (layer0_outputs(664)) and not (layer0_outputs(2178));
    outputs(9882) <= layer0_outputs(9856);
    outputs(9883) <= (layer0_outputs(2409)) xor (layer0_outputs(3644));
    outputs(9884) <= layer0_outputs(589);
    outputs(9885) <= (layer0_outputs(6747)) xor (layer0_outputs(7851));
    outputs(9886) <= not(layer0_outputs(9409));
    outputs(9887) <= (layer0_outputs(8062)) xor (layer0_outputs(6064));
    outputs(9888) <= layer0_outputs(616);
    outputs(9889) <= not((layer0_outputs(7227)) xor (layer0_outputs(3245)));
    outputs(9890) <= not(layer0_outputs(4199));
    outputs(9891) <= (layer0_outputs(3545)) xor (layer0_outputs(4485));
    outputs(9892) <= not((layer0_outputs(8029)) xor (layer0_outputs(4663)));
    outputs(9893) <= layer0_outputs(2899);
    outputs(9894) <= layer0_outputs(4065);
    outputs(9895) <= not((layer0_outputs(734)) xor (layer0_outputs(4893)));
    outputs(9896) <= (layer0_outputs(4501)) xor (layer0_outputs(8875));
    outputs(9897) <= layer0_outputs(6472);
    outputs(9898) <= (layer0_outputs(9690)) and not (layer0_outputs(813));
    outputs(9899) <= not((layer0_outputs(4018)) xor (layer0_outputs(85)));
    outputs(9900) <= (layer0_outputs(3801)) and (layer0_outputs(9359));
    outputs(9901) <= (layer0_outputs(8792)) and (layer0_outputs(973));
    outputs(9902) <= (layer0_outputs(8384)) and not (layer0_outputs(686));
    outputs(9903) <= layer0_outputs(1862);
    outputs(9904) <= (layer0_outputs(7126)) xor (layer0_outputs(9464));
    outputs(9905) <= not((layer0_outputs(4165)) xor (layer0_outputs(941)));
    outputs(9906) <= (layer0_outputs(1019)) xor (layer0_outputs(3357));
    outputs(9907) <= not(layer0_outputs(7964));
    outputs(9908) <= not((layer0_outputs(2217)) or (layer0_outputs(3461)));
    outputs(9909) <= not((layer0_outputs(6589)) and (layer0_outputs(4094)));
    outputs(9910) <= (layer0_outputs(7092)) xor (layer0_outputs(7428));
    outputs(9911) <= layer0_outputs(5207);
    outputs(9912) <= layer0_outputs(8780);
    outputs(9913) <= not(layer0_outputs(4814)) or (layer0_outputs(3410));
    outputs(9914) <= (layer0_outputs(1582)) or (layer0_outputs(1506));
    outputs(9915) <= (layer0_outputs(606)) and not (layer0_outputs(8181));
    outputs(9916) <= not((layer0_outputs(4947)) xor (layer0_outputs(4781)));
    outputs(9917) <= not((layer0_outputs(4734)) xor (layer0_outputs(10055)));
    outputs(9918) <= not(layer0_outputs(297));
    outputs(9919) <= not(layer0_outputs(7458));
    outputs(9920) <= not(layer0_outputs(3493));
    outputs(9921) <= (layer0_outputs(1443)) xor (layer0_outputs(210));
    outputs(9922) <= (layer0_outputs(4376)) and not (layer0_outputs(6840));
    outputs(9923) <= layer0_outputs(4681);
    outputs(9924) <= layer0_outputs(3297);
    outputs(9925) <= (layer0_outputs(8792)) and not (layer0_outputs(3741));
    outputs(9926) <= (layer0_outputs(174)) and not (layer0_outputs(9233));
    outputs(9927) <= '0';
    outputs(9928) <= not((layer0_outputs(8944)) or (layer0_outputs(9369)));
    outputs(9929) <= not(layer0_outputs(4512));
    outputs(9930) <= layer0_outputs(7994);
    outputs(9931) <= (layer0_outputs(2941)) and not (layer0_outputs(1743));
    outputs(9932) <= not((layer0_outputs(3989)) xor (layer0_outputs(201)));
    outputs(9933) <= not((layer0_outputs(9475)) xor (layer0_outputs(7634)));
    outputs(9934) <= not((layer0_outputs(2950)) xor (layer0_outputs(3771)));
    outputs(9935) <= layer0_outputs(9667);
    outputs(9936) <= not(layer0_outputs(8377));
    outputs(9937) <= (layer0_outputs(1935)) and (layer0_outputs(252));
    outputs(9938) <= not((layer0_outputs(5528)) or (layer0_outputs(3604)));
    outputs(9939) <= not(layer0_outputs(3130));
    outputs(9940) <= not((layer0_outputs(0)) xor (layer0_outputs(5767)));
    outputs(9941) <= '0';
    outputs(9942) <= not(layer0_outputs(7245));
    outputs(9943) <= layer0_outputs(6083);
    outputs(9944) <= (layer0_outputs(9719)) xor (layer0_outputs(5479));
    outputs(9945) <= not((layer0_outputs(4837)) or (layer0_outputs(5172)));
    outputs(9946) <= (layer0_outputs(7009)) and (layer0_outputs(2477));
    outputs(9947) <= (layer0_outputs(9946)) and not (layer0_outputs(3384));
    outputs(9948) <= not((layer0_outputs(1914)) xor (layer0_outputs(9411)));
    outputs(9949) <= (layer0_outputs(8424)) and (layer0_outputs(7829));
    outputs(9950) <= not(layer0_outputs(3573));
    outputs(9951) <= not(layer0_outputs(3704));
    outputs(9952) <= (layer0_outputs(8071)) and not (layer0_outputs(7150));
    outputs(9953) <= not(layer0_outputs(6824));
    outputs(9954) <= not((layer0_outputs(3346)) and (layer0_outputs(1233)));
    outputs(9955) <= (layer0_outputs(9837)) xor (layer0_outputs(7629));
    outputs(9956) <= (layer0_outputs(4553)) and not (layer0_outputs(2092));
    outputs(9957) <= (layer0_outputs(295)) xor (layer0_outputs(7849));
    outputs(9958) <= (layer0_outputs(4834)) and (layer0_outputs(8806));
    outputs(9959) <= (layer0_outputs(8256)) and (layer0_outputs(532));
    outputs(9960) <= not((layer0_outputs(449)) xor (layer0_outputs(6296)));
    outputs(9961) <= layer0_outputs(1543);
    outputs(9962) <= (layer0_outputs(6117)) or (layer0_outputs(1972));
    outputs(9963) <= not(layer0_outputs(4638));
    outputs(9964) <= not(layer0_outputs(5580));
    outputs(9965) <= not(layer0_outputs(7859));
    outputs(9966) <= not((layer0_outputs(5181)) xor (layer0_outputs(5510)));
    outputs(9967) <= layer0_outputs(214);
    outputs(9968) <= (layer0_outputs(7444)) xor (layer0_outputs(3195));
    outputs(9969) <= not((layer0_outputs(2077)) xor (layer0_outputs(5709)));
    outputs(9970) <= (layer0_outputs(7152)) and not (layer0_outputs(3812));
    outputs(9971) <= (layer0_outputs(5874)) xor (layer0_outputs(6784));
    outputs(9972) <= not(layer0_outputs(5282));
    outputs(9973) <= not(layer0_outputs(7415));
    outputs(9974) <= not((layer0_outputs(1067)) xor (layer0_outputs(5105)));
    outputs(9975) <= (layer0_outputs(3476)) or (layer0_outputs(5160));
    outputs(9976) <= not((layer0_outputs(4798)) or (layer0_outputs(4803)));
    outputs(9977) <= (layer0_outputs(4666)) xor (layer0_outputs(8989));
    outputs(9978) <= not((layer0_outputs(3687)) xor (layer0_outputs(2261)));
    outputs(9979) <= not(layer0_outputs(10226)) or (layer0_outputs(9156));
    outputs(9980) <= not(layer0_outputs(244));
    outputs(9981) <= not(layer0_outputs(7325));
    outputs(9982) <= not((layer0_outputs(9732)) xor (layer0_outputs(4419)));
    outputs(9983) <= not((layer0_outputs(2664)) xor (layer0_outputs(215)));
    outputs(9984) <= not(layer0_outputs(330));
    outputs(9985) <= (layer0_outputs(6164)) xor (layer0_outputs(8492));
    outputs(9986) <= not((layer0_outputs(7061)) xor (layer0_outputs(1014)));
    outputs(9987) <= (layer0_outputs(3571)) and not (layer0_outputs(10178));
    outputs(9988) <= layer0_outputs(199);
    outputs(9989) <= not(layer0_outputs(9170));
    outputs(9990) <= not(layer0_outputs(7430));
    outputs(9991) <= not(layer0_outputs(9842));
    outputs(9992) <= not((layer0_outputs(4437)) and (layer0_outputs(9658)));
    outputs(9993) <= (layer0_outputs(2609)) and (layer0_outputs(1026));
    outputs(9994) <= not(layer0_outputs(1537));
    outputs(9995) <= (layer0_outputs(323)) or (layer0_outputs(9918));
    outputs(9996) <= (layer0_outputs(337)) and not (layer0_outputs(9493));
    outputs(9997) <= layer0_outputs(439);
    outputs(9998) <= not(layer0_outputs(3213));
    outputs(9999) <= not((layer0_outputs(9498)) xor (layer0_outputs(975)));
    outputs(10000) <= not((layer0_outputs(1756)) xor (layer0_outputs(9024)));
    outputs(10001) <= not(layer0_outputs(5518)) or (layer0_outputs(1421));
    outputs(10002) <= not(layer0_outputs(3113));
    outputs(10003) <= not((layer0_outputs(10086)) xor (layer0_outputs(7058)));
    outputs(10004) <= layer0_outputs(3451);
    outputs(10005) <= layer0_outputs(316);
    outputs(10006) <= (layer0_outputs(7340)) and (layer0_outputs(4917));
    outputs(10007) <= not((layer0_outputs(9483)) or (layer0_outputs(9047)));
    outputs(10008) <= not(layer0_outputs(2086));
    outputs(10009) <= not(layer0_outputs(4689));
    outputs(10010) <= (layer0_outputs(2583)) xor (layer0_outputs(5244));
    outputs(10011) <= layer0_outputs(8680);
    outputs(10012) <= not((layer0_outputs(3389)) and (layer0_outputs(2853)));
    outputs(10013) <= (layer0_outputs(709)) and not (layer0_outputs(1211));
    outputs(10014) <= layer0_outputs(68);
    outputs(10015) <= not((layer0_outputs(8803)) or (layer0_outputs(1277)));
    outputs(10016) <= (layer0_outputs(4360)) xor (layer0_outputs(8541));
    outputs(10017) <= (layer0_outputs(1442)) or (layer0_outputs(9568));
    outputs(10018) <= layer0_outputs(2689);
    outputs(10019) <= layer0_outputs(5777);
    outputs(10020) <= not(layer0_outputs(6352));
    outputs(10021) <= (layer0_outputs(2319)) xor (layer0_outputs(6372));
    outputs(10022) <= (layer0_outputs(4370)) and (layer0_outputs(10077));
    outputs(10023) <= (layer0_outputs(10201)) and not (layer0_outputs(6914));
    outputs(10024) <= (layer0_outputs(1174)) and (layer0_outputs(9639));
    outputs(10025) <= not((layer0_outputs(2588)) xor (layer0_outputs(7559)));
    outputs(10026) <= (layer0_outputs(5116)) xor (layer0_outputs(1270));
    outputs(10027) <= (layer0_outputs(2682)) xor (layer0_outputs(8268));
    outputs(10028) <= not(layer0_outputs(2815));
    outputs(10029) <= (layer0_outputs(4252)) and not (layer0_outputs(6861));
    outputs(10030) <= (layer0_outputs(1232)) and not (layer0_outputs(5320));
    outputs(10031) <= not(layer0_outputs(2583)) or (layer0_outputs(8209));
    outputs(10032) <= not((layer0_outputs(1806)) or (layer0_outputs(2075)));
    outputs(10033) <= not((layer0_outputs(4549)) xor (layer0_outputs(3566)));
    outputs(10034) <= not(layer0_outputs(3082)) or (layer0_outputs(1540));
    outputs(10035) <= not(layer0_outputs(3964));
    outputs(10036) <= (layer0_outputs(4909)) and not (layer0_outputs(840));
    outputs(10037) <= not((layer0_outputs(8155)) xor (layer0_outputs(3444)));
    outputs(10038) <= (layer0_outputs(6212)) and (layer0_outputs(3830));
    outputs(10039) <= (layer0_outputs(758)) and not (layer0_outputs(9339));
    outputs(10040) <= (layer0_outputs(5620)) and (layer0_outputs(9006));
    outputs(10041) <= not(layer0_outputs(7806));
    outputs(10042) <= not(layer0_outputs(7002));
    outputs(10043) <= not(layer0_outputs(7996));
    outputs(10044) <= (layer0_outputs(6817)) xor (layer0_outputs(9688));
    outputs(10045) <= layer0_outputs(2993);
    outputs(10046) <= not((layer0_outputs(5190)) xor (layer0_outputs(4001)));
    outputs(10047) <= (layer0_outputs(8631)) or (layer0_outputs(7197));
    outputs(10048) <= not((layer0_outputs(9929)) or (layer0_outputs(2506)));
    outputs(10049) <= (layer0_outputs(6058)) or (layer0_outputs(7109));
    outputs(10050) <= (layer0_outputs(7911)) xor (layer0_outputs(6515));
    outputs(10051) <= (layer0_outputs(9406)) and (layer0_outputs(6304));
    outputs(10052) <= (layer0_outputs(4892)) and not (layer0_outputs(5700));
    outputs(10053) <= not((layer0_outputs(6669)) and (layer0_outputs(9671)));
    outputs(10054) <= layer0_outputs(1948);
    outputs(10055) <= (layer0_outputs(1984)) and (layer0_outputs(984));
    outputs(10056) <= layer0_outputs(9);
    outputs(10057) <= not(layer0_outputs(4830)) or (layer0_outputs(3522));
    outputs(10058) <= (layer0_outputs(8623)) or (layer0_outputs(1548));
    outputs(10059) <= not(layer0_outputs(6737));
    outputs(10060) <= not(layer0_outputs(7841)) or (layer0_outputs(9520));
    outputs(10061) <= (layer0_outputs(6760)) and not (layer0_outputs(6105));
    outputs(10062) <= layer0_outputs(8948);
    outputs(10063) <= not((layer0_outputs(2260)) xor (layer0_outputs(2643)));
    outputs(10064) <= not(layer0_outputs(3404));
    outputs(10065) <= (layer0_outputs(3836)) and (layer0_outputs(7954));
    outputs(10066) <= not(layer0_outputs(4878));
    outputs(10067) <= not((layer0_outputs(9681)) xor (layer0_outputs(899)));
    outputs(10068) <= not((layer0_outputs(8575)) xor (layer0_outputs(1869)));
    outputs(10069) <= (layer0_outputs(5785)) xor (layer0_outputs(4855));
    outputs(10070) <= (layer0_outputs(3904)) and not (layer0_outputs(859));
    outputs(10071) <= not((layer0_outputs(1246)) or (layer0_outputs(2103)));
    outputs(10072) <= not((layer0_outputs(9879)) xor (layer0_outputs(2467)));
    outputs(10073) <= not((layer0_outputs(4428)) xor (layer0_outputs(8253)));
    outputs(10074) <= not((layer0_outputs(8978)) xor (layer0_outputs(9723)));
    outputs(10075) <= not(layer0_outputs(1323)) or (layer0_outputs(7637));
    outputs(10076) <= layer0_outputs(7361);
    outputs(10077) <= (layer0_outputs(2472)) and (layer0_outputs(6742));
    outputs(10078) <= (layer0_outputs(2250)) or (layer0_outputs(865));
    outputs(10079) <= layer0_outputs(7015);
    outputs(10080) <= layer0_outputs(3660);
    outputs(10081) <= (layer0_outputs(950)) and not (layer0_outputs(106));
    outputs(10082) <= layer0_outputs(1315);
    outputs(10083) <= (layer0_outputs(8725)) and (layer0_outputs(6780));
    outputs(10084) <= layer0_outputs(10193);
    outputs(10085) <= layer0_outputs(920);
    outputs(10086) <= layer0_outputs(2440);
    outputs(10087) <= not((layer0_outputs(5322)) and (layer0_outputs(9807)));
    outputs(10088) <= (layer0_outputs(8609)) and not (layer0_outputs(3157));
    outputs(10089) <= '1';
    outputs(10090) <= not(layer0_outputs(8931));
    outputs(10091) <= not(layer0_outputs(6620)) or (layer0_outputs(9753));
    outputs(10092) <= not((layer0_outputs(9419)) or (layer0_outputs(2587)));
    outputs(10093) <= not((layer0_outputs(4915)) xor (layer0_outputs(8547)));
    outputs(10094) <= not((layer0_outputs(3946)) xor (layer0_outputs(4377)));
    outputs(10095) <= not(layer0_outputs(1292)) or (layer0_outputs(3430));
    outputs(10096) <= (layer0_outputs(7083)) and not (layer0_outputs(5867));
    outputs(10097) <= (layer0_outputs(4523)) and not (layer0_outputs(7997));
    outputs(10098) <= not((layer0_outputs(5474)) xor (layer0_outputs(1938)));
    outputs(10099) <= not(layer0_outputs(9058));
    outputs(10100) <= (layer0_outputs(8810)) and not (layer0_outputs(8142));
    outputs(10101) <= layer0_outputs(1913);
    outputs(10102) <= not(layer0_outputs(9121));
    outputs(10103) <= not((layer0_outputs(1395)) xor (layer0_outputs(2213)));
    outputs(10104) <= (layer0_outputs(7147)) or (layer0_outputs(10038));
    outputs(10105) <= not(layer0_outputs(1123)) or (layer0_outputs(301));
    outputs(10106) <= (layer0_outputs(8222)) and not (layer0_outputs(9571));
    outputs(10107) <= (layer0_outputs(7579)) xor (layer0_outputs(2904));
    outputs(10108) <= layer0_outputs(413);
    outputs(10109) <= not(layer0_outputs(10089));
    outputs(10110) <= not(layer0_outputs(9643));
    outputs(10111) <= layer0_outputs(9003);
    outputs(10112) <= '0';
    outputs(10113) <= not(layer0_outputs(7382));
    outputs(10114) <= (layer0_outputs(1418)) and not (layer0_outputs(8833));
    outputs(10115) <= not((layer0_outputs(4813)) or (layer0_outputs(4051)));
    outputs(10116) <= (layer0_outputs(6610)) and not (layer0_outputs(7582));
    outputs(10117) <= not((layer0_outputs(8649)) xor (layer0_outputs(8511)));
    outputs(10118) <= not((layer0_outputs(6595)) xor (layer0_outputs(5848)));
    outputs(10119) <= layer0_outputs(3735);
    outputs(10120) <= (layer0_outputs(6590)) and not (layer0_outputs(940));
    outputs(10121) <= (layer0_outputs(2479)) and (layer0_outputs(8794));
    outputs(10122) <= not((layer0_outputs(9818)) or (layer0_outputs(4299)));
    outputs(10123) <= not((layer0_outputs(4994)) or (layer0_outputs(10233)));
    outputs(10124) <= (layer0_outputs(2185)) and (layer0_outputs(3863));
    outputs(10125) <= (layer0_outputs(381)) and not (layer0_outputs(5361));
    outputs(10126) <= layer0_outputs(7203);
    outputs(10127) <= layer0_outputs(3200);
    outputs(10128) <= (layer0_outputs(6675)) and not (layer0_outputs(9737));
    outputs(10129) <= layer0_outputs(832);
    outputs(10130) <= not(layer0_outputs(3129)) or (layer0_outputs(5331));
    outputs(10131) <= not((layer0_outputs(2833)) xor (layer0_outputs(9948)));
    outputs(10132) <= not((layer0_outputs(8270)) and (layer0_outputs(8736)));
    outputs(10133) <= not(layer0_outputs(4067));
    outputs(10134) <= not(layer0_outputs(7320));
    outputs(10135) <= not(layer0_outputs(2296)) or (layer0_outputs(8684));
    outputs(10136) <= (layer0_outputs(7984)) xor (layer0_outputs(7006));
    outputs(10137) <= (layer0_outputs(7506)) xor (layer0_outputs(6278));
    outputs(10138) <= layer0_outputs(8236);
    outputs(10139) <= layer0_outputs(4792);
    outputs(10140) <= not(layer0_outputs(3133)) or (layer0_outputs(9660));
    outputs(10141) <= not((layer0_outputs(5595)) xor (layer0_outputs(3953)));
    outputs(10142) <= layer0_outputs(8710);
    outputs(10143) <= not(layer0_outputs(4598));
    outputs(10144) <= not(layer0_outputs(6087));
    outputs(10145) <= layer0_outputs(7519);
    outputs(10146) <= not((layer0_outputs(5890)) xor (layer0_outputs(4777)));
    outputs(10147) <= layer0_outputs(3530);
    outputs(10148) <= not((layer0_outputs(7354)) or (layer0_outputs(9397)));
    outputs(10149) <= not((layer0_outputs(2838)) or (layer0_outputs(2444)));
    outputs(10150) <= (layer0_outputs(6400)) and (layer0_outputs(1513));
    outputs(10151) <= layer0_outputs(1106);
    outputs(10152) <= not(layer0_outputs(6283));
    outputs(10153) <= not(layer0_outputs(7142)) or (layer0_outputs(7082));
    outputs(10154) <= not((layer0_outputs(8495)) xor (layer0_outputs(4903)));
    outputs(10155) <= not(layer0_outputs(6978));
    outputs(10156) <= layer0_outputs(9398);
    outputs(10157) <= not(layer0_outputs(10151));
    outputs(10158) <= (layer0_outputs(4328)) and not (layer0_outputs(3093));
    outputs(10159) <= not((layer0_outputs(1765)) xor (layer0_outputs(10215)));
    outputs(10160) <= (layer0_outputs(6217)) and not (layer0_outputs(8178));
    outputs(10161) <= layer0_outputs(2229);
    outputs(10162) <= (layer0_outputs(3903)) and not (layer0_outputs(9206));
    outputs(10163) <= (layer0_outputs(9132)) and not (layer0_outputs(7193));
    outputs(10164) <= (layer0_outputs(6264)) xor (layer0_outputs(6864));
    outputs(10165) <= layer0_outputs(559);
    outputs(10166) <= (layer0_outputs(8489)) and (layer0_outputs(6351));
    outputs(10167) <= not(layer0_outputs(7844));
    outputs(10168) <= (layer0_outputs(5394)) and not (layer0_outputs(841));
    outputs(10169) <= layer0_outputs(5895);
    outputs(10170) <= layer0_outputs(8211);
    outputs(10171) <= layer0_outputs(1089);
    outputs(10172) <= not(layer0_outputs(5203));
    outputs(10173) <= (layer0_outputs(5757)) and (layer0_outputs(9732));
    outputs(10174) <= layer0_outputs(3810);
    outputs(10175) <= not(layer0_outputs(7123));
    outputs(10176) <= not(layer0_outputs(5912));
    outputs(10177) <= layer0_outputs(2862);
    outputs(10178) <= not((layer0_outputs(4014)) xor (layer0_outputs(3389)));
    outputs(10179) <= (layer0_outputs(7536)) and not (layer0_outputs(323));
    outputs(10180) <= (layer0_outputs(5986)) and not (layer0_outputs(10179));
    outputs(10181) <= not(layer0_outputs(6263));
    outputs(10182) <= layer0_outputs(10183);
    outputs(10183) <= layer0_outputs(4770);
    outputs(10184) <= not(layer0_outputs(5631)) or (layer0_outputs(199));
    outputs(10185) <= (layer0_outputs(4406)) and (layer0_outputs(5086));
    outputs(10186) <= (layer0_outputs(8538)) and (layer0_outputs(6573));
    outputs(10187) <= not(layer0_outputs(5606)) or (layer0_outputs(7111));
    outputs(10188) <= layer0_outputs(8452);
    outputs(10189) <= not((layer0_outputs(9799)) or (layer0_outputs(9534)));
    outputs(10190) <= not((layer0_outputs(5506)) xor (layer0_outputs(9872)));
    outputs(10191) <= not(layer0_outputs(8334));
    outputs(10192) <= not(layer0_outputs(2008));
    outputs(10193) <= layer0_outputs(1469);
    outputs(10194) <= not((layer0_outputs(7590)) xor (layer0_outputs(6106)));
    outputs(10195) <= not(layer0_outputs(5541)) or (layer0_outputs(10004));
    outputs(10196) <= not(layer0_outputs(2990)) or (layer0_outputs(4735));
    outputs(10197) <= (layer0_outputs(10095)) and not (layer0_outputs(740));
    outputs(10198) <= (layer0_outputs(5380)) and not (layer0_outputs(551));
    outputs(10199) <= not(layer0_outputs(9649));
    outputs(10200) <= not((layer0_outputs(3128)) xor (layer0_outputs(4207)));
    outputs(10201) <= (layer0_outputs(2224)) xor (layer0_outputs(6586));
    outputs(10202) <= not((layer0_outputs(3785)) xor (layer0_outputs(783)));
    outputs(10203) <= layer0_outputs(4496);
    outputs(10204) <= not(layer0_outputs(6997));
    outputs(10205) <= (layer0_outputs(6180)) xor (layer0_outputs(6991));
    outputs(10206) <= (layer0_outputs(114)) and (layer0_outputs(5750));
    outputs(10207) <= not((layer0_outputs(2264)) xor (layer0_outputs(332)));
    outputs(10208) <= not(layer0_outputs(3908));
    outputs(10209) <= (layer0_outputs(7049)) and not (layer0_outputs(6740));
    outputs(10210) <= not(layer0_outputs(9964));
    outputs(10211) <= (layer0_outputs(9902)) xor (layer0_outputs(9000));
    outputs(10212) <= not(layer0_outputs(10061));
    outputs(10213) <= not(layer0_outputs(9456));
    outputs(10214) <= not(layer0_outputs(9232));
    outputs(10215) <= layer0_outputs(6292);
    outputs(10216) <= not((layer0_outputs(9230)) xor (layer0_outputs(2013)));
    outputs(10217) <= not((layer0_outputs(9747)) xor (layer0_outputs(3492)));
    outputs(10218) <= (layer0_outputs(620)) xor (layer0_outputs(5859));
    outputs(10219) <= not(layer0_outputs(4884)) or (layer0_outputs(7034));
    outputs(10220) <= (layer0_outputs(1551)) xor (layer0_outputs(9300));
    outputs(10221) <= not(layer0_outputs(834)) or (layer0_outputs(7372));
    outputs(10222) <= not(layer0_outputs(8477)) or (layer0_outputs(2561));
    outputs(10223) <= (layer0_outputs(9365)) and not (layer0_outputs(1808));
    outputs(10224) <= (layer0_outputs(8128)) xor (layer0_outputs(8356));
    outputs(10225) <= (layer0_outputs(6501)) and (layer0_outputs(2019));
    outputs(10226) <= not(layer0_outputs(4914)) or (layer0_outputs(6794));
    outputs(10227) <= (layer0_outputs(7250)) and not (layer0_outputs(3499));
    outputs(10228) <= layer0_outputs(1653);
    outputs(10229) <= (layer0_outputs(2030)) xor (layer0_outputs(8814));
    outputs(10230) <= not(layer0_outputs(5135));
    outputs(10231) <= not(layer0_outputs(2589));
    outputs(10232) <= layer0_outputs(3602);
    outputs(10233) <= (layer0_outputs(2742)) and not (layer0_outputs(6603));
    outputs(10234) <= (layer0_outputs(7560)) and not (layer0_outputs(1482));
    outputs(10235) <= layer0_outputs(3001);
    outputs(10236) <= (layer0_outputs(9542)) xor (layer0_outputs(9552));
    outputs(10237) <= not(layer0_outputs(7971));
    outputs(10238) <= not((layer0_outputs(5862)) xor (layer0_outputs(3578)));
    outputs(10239) <= (layer0_outputs(5979)) xor (layer0_outputs(5004));

end Behavioral;
