library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs : in std_logic_vector(255 downto 0);
        outputs : out std_logic_vector(7679 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs : std_logic_vector(7679 downto 0);

begin

    layer0_outputs(0) <= not(inputs(139)) or (inputs(41));
    layer0_outputs(1) <= not(inputs(50));
    layer0_outputs(2) <= (inputs(42)) or (inputs(33));
    layer0_outputs(3) <= (inputs(45)) xor (inputs(30));
    layer0_outputs(4) <= inputs(195);
    layer0_outputs(5) <= not((inputs(255)) xor (inputs(96)));
    layer0_outputs(6) <= not((inputs(248)) or (inputs(215)));
    layer0_outputs(7) <= not((inputs(94)) or (inputs(6)));
    layer0_outputs(8) <= (inputs(45)) or (inputs(29));
    layer0_outputs(9) <= not(inputs(44));
    layer0_outputs(10) <= (inputs(4)) or (inputs(227));
    layer0_outputs(11) <= (inputs(204)) and not (inputs(112));
    layer0_outputs(12) <= not(inputs(74));
    layer0_outputs(13) <= not(inputs(247)) or (inputs(123));
    layer0_outputs(14) <= (inputs(160)) and not (inputs(147));
    layer0_outputs(15) <= (inputs(39)) and not (inputs(221));
    layer0_outputs(16) <= inputs(204);
    layer0_outputs(17) <= inputs(58);
    layer0_outputs(18) <= not(inputs(168)) or (inputs(79));
    layer0_outputs(19) <= not(inputs(209));
    layer0_outputs(20) <= not(inputs(18));
    layer0_outputs(21) <= not((inputs(97)) or (inputs(104)));
    layer0_outputs(22) <= (inputs(185)) and not (inputs(235));
    layer0_outputs(23) <= inputs(88);
    layer0_outputs(24) <= not(inputs(193));
    layer0_outputs(25) <= not((inputs(38)) or (inputs(47)));
    layer0_outputs(26) <= not(inputs(208)) or (inputs(234));
    layer0_outputs(27) <= not((inputs(163)) or (inputs(251)));
    layer0_outputs(28) <= not(inputs(183));
    layer0_outputs(29) <= (inputs(37)) or (inputs(46));
    layer0_outputs(30) <= inputs(185);
    layer0_outputs(31) <= inputs(145);
    layer0_outputs(32) <= (inputs(54)) and not (inputs(105));
    layer0_outputs(33) <= not((inputs(193)) or (inputs(176)));
    layer0_outputs(34) <= not((inputs(80)) or (inputs(53)));
    layer0_outputs(35) <= not((inputs(83)) or (inputs(65)));
    layer0_outputs(36) <= (inputs(24)) xor (inputs(55));
    layer0_outputs(37) <= not((inputs(81)) or (inputs(156)));
    layer0_outputs(38) <= not(inputs(76));
    layer0_outputs(39) <= not(inputs(31));
    layer0_outputs(40) <= '1';
    layer0_outputs(41) <= not((inputs(9)) and (inputs(161)));
    layer0_outputs(42) <= (inputs(179)) or (inputs(175));
    layer0_outputs(43) <= not(inputs(139));
    layer0_outputs(44) <= not(inputs(77));
    layer0_outputs(45) <= not(inputs(205)) or (inputs(107));
    layer0_outputs(46) <= (inputs(46)) or (inputs(101));
    layer0_outputs(47) <= (inputs(122)) xor (inputs(134));
    layer0_outputs(48) <= not(inputs(13));
    layer0_outputs(49) <= (inputs(164)) and not (inputs(94));
    layer0_outputs(50) <= not(inputs(234));
    layer0_outputs(51) <= (inputs(52)) or (inputs(6));
    layer0_outputs(52) <= not(inputs(53));
    layer0_outputs(53) <= not((inputs(10)) xor (inputs(106)));
    layer0_outputs(54) <= inputs(22);
    layer0_outputs(55) <= not(inputs(22));
    layer0_outputs(56) <= not(inputs(230));
    layer0_outputs(57) <= inputs(201);
    layer0_outputs(58) <= not(inputs(26));
    layer0_outputs(59) <= not(inputs(214));
    layer0_outputs(60) <= (inputs(184)) and not (inputs(111));
    layer0_outputs(61) <= (inputs(112)) or (inputs(131));
    layer0_outputs(62) <= (inputs(230)) or (inputs(254));
    layer0_outputs(63) <= not((inputs(83)) or (inputs(46)));
    layer0_outputs(64) <= (inputs(212)) and not (inputs(19));
    layer0_outputs(65) <= not(inputs(0)) or (inputs(237));
    layer0_outputs(66) <= not(inputs(19));
    layer0_outputs(67) <= (inputs(202)) xor (inputs(38));
    layer0_outputs(68) <= (inputs(104)) and (inputs(26));
    layer0_outputs(69) <= not((inputs(142)) or (inputs(32)));
    layer0_outputs(70) <= not(inputs(42));
    layer0_outputs(71) <= inputs(175);
    layer0_outputs(72) <= '0';
    layer0_outputs(73) <= not((inputs(163)) or (inputs(195)));
    layer0_outputs(74) <= (inputs(194)) or (inputs(222));
    layer0_outputs(75) <= (inputs(179)) or (inputs(64));
    layer0_outputs(76) <= not((inputs(96)) or (inputs(252)));
    layer0_outputs(77) <= not((inputs(21)) or (inputs(30)));
    layer0_outputs(78) <= not(inputs(229));
    layer0_outputs(79) <= not(inputs(179)) or (inputs(95));
    layer0_outputs(80) <= (inputs(156)) or (inputs(172));
    layer0_outputs(81) <= not((inputs(102)) or (inputs(47)));
    layer0_outputs(82) <= inputs(249);
    layer0_outputs(83) <= not((inputs(221)) and (inputs(114)));
    layer0_outputs(84) <= (inputs(8)) and not (inputs(162));
    layer0_outputs(85) <= (inputs(189)) or (inputs(3));
    layer0_outputs(86) <= (inputs(38)) and not (inputs(109));
    layer0_outputs(87) <= (inputs(157)) and not (inputs(45));
    layer0_outputs(88) <= not(inputs(88));
    layer0_outputs(89) <= not(inputs(50));
    layer0_outputs(90) <= (inputs(166)) and not (inputs(238));
    layer0_outputs(91) <= (inputs(194)) xor (inputs(198));
    layer0_outputs(92) <= (inputs(203)) and not (inputs(32));
    layer0_outputs(93) <= not(inputs(93));
    layer0_outputs(94) <= (inputs(216)) or (inputs(176));
    layer0_outputs(95) <= not((inputs(22)) xor (inputs(177)));
    layer0_outputs(96) <= (inputs(106)) and not (inputs(149));
    layer0_outputs(97) <= not(inputs(136)) or (inputs(57));
    layer0_outputs(98) <= '0';
    layer0_outputs(99) <= (inputs(28)) or (inputs(15));
    layer0_outputs(100) <= inputs(100);
    layer0_outputs(101) <= inputs(42);
    layer0_outputs(102) <= inputs(156);
    layer0_outputs(103) <= (inputs(146)) xor (inputs(12));
    layer0_outputs(104) <= (inputs(225)) or (inputs(193));
    layer0_outputs(105) <= inputs(35);
    layer0_outputs(106) <= not(inputs(134));
    layer0_outputs(107) <= inputs(23);
    layer0_outputs(108) <= not(inputs(153));
    layer0_outputs(109) <= not(inputs(104));
    layer0_outputs(110) <= (inputs(122)) and not (inputs(44));
    layer0_outputs(111) <= not(inputs(128));
    layer0_outputs(112) <= not(inputs(125)) or (inputs(250));
    layer0_outputs(113) <= not(inputs(2));
    layer0_outputs(114) <= (inputs(122)) and not (inputs(214));
    layer0_outputs(115) <= not((inputs(126)) or (inputs(8)));
    layer0_outputs(116) <= (inputs(140)) or (inputs(59));
    layer0_outputs(117) <= not(inputs(199)) or (inputs(25));
    layer0_outputs(118) <= not((inputs(170)) and (inputs(251)));
    layer0_outputs(119) <= not((inputs(223)) xor (inputs(140)));
    layer0_outputs(120) <= (inputs(108)) xor (inputs(89));
    layer0_outputs(121) <= (inputs(103)) xor (inputs(173));
    layer0_outputs(122) <= not((inputs(37)) or (inputs(221)));
    layer0_outputs(123) <= inputs(129);
    layer0_outputs(124) <= (inputs(169)) or (inputs(3));
    layer0_outputs(125) <= (inputs(121)) and (inputs(69));
    layer0_outputs(126) <= inputs(212);
    layer0_outputs(127) <= (inputs(212)) and not (inputs(52));
    layer0_outputs(128) <= not(inputs(233)) or (inputs(43));
    layer0_outputs(129) <= (inputs(0)) or (inputs(216));
    layer0_outputs(130) <= (inputs(195)) and not (inputs(125));
    layer0_outputs(131) <= not((inputs(59)) xor (inputs(107)));
    layer0_outputs(132) <= not((inputs(213)) or (inputs(108)));
    layer0_outputs(133) <= (inputs(141)) and not (inputs(19));
    layer0_outputs(134) <= not(inputs(161));
    layer0_outputs(135) <= (inputs(38)) and not (inputs(109));
    layer0_outputs(136) <= (inputs(113)) and not (inputs(57));
    layer0_outputs(137) <= inputs(231);
    layer0_outputs(138) <= not(inputs(167)) or (inputs(158));
    layer0_outputs(139) <= (inputs(248)) or (inputs(143));
    layer0_outputs(140) <= (inputs(253)) and not (inputs(207));
    layer0_outputs(141) <= not(inputs(50));
    layer0_outputs(142) <= inputs(236);
    layer0_outputs(143) <= not(inputs(197));
    layer0_outputs(144) <= inputs(38);
    layer0_outputs(145) <= not((inputs(60)) xor (inputs(113)));
    layer0_outputs(146) <= not((inputs(193)) or (inputs(167)));
    layer0_outputs(147) <= (inputs(220)) or (inputs(222));
    layer0_outputs(148) <= (inputs(196)) and not (inputs(221));
    layer0_outputs(149) <= not((inputs(111)) or (inputs(138)));
    layer0_outputs(150) <= not(inputs(196)) or (inputs(17));
    layer0_outputs(151) <= not((inputs(42)) or (inputs(206)));
    layer0_outputs(152) <= not(inputs(96));
    layer0_outputs(153) <= not((inputs(7)) or (inputs(92)));
    layer0_outputs(154) <= not(inputs(202));
    layer0_outputs(155) <= inputs(221);
    layer0_outputs(156) <= not((inputs(46)) xor (inputs(60)));
    layer0_outputs(157) <= not(inputs(62));
    layer0_outputs(158) <= not((inputs(34)) xor (inputs(242)));
    layer0_outputs(159) <= not(inputs(137));
    layer0_outputs(160) <= inputs(101);
    layer0_outputs(161) <= not(inputs(105));
    layer0_outputs(162) <= (inputs(6)) and not (inputs(239));
    layer0_outputs(163) <= (inputs(39)) xor (inputs(161));
    layer0_outputs(164) <= not(inputs(244)) or (inputs(181));
    layer0_outputs(165) <= (inputs(154)) and not (inputs(14));
    layer0_outputs(166) <= not(inputs(60)) or (inputs(33));
    layer0_outputs(167) <= not(inputs(99));
    layer0_outputs(168) <= not(inputs(194)) or (inputs(128));
    layer0_outputs(169) <= inputs(164);
    layer0_outputs(170) <= not((inputs(38)) or (inputs(15)));
    layer0_outputs(171) <= inputs(84);
    layer0_outputs(172) <= not((inputs(248)) xor (inputs(14)));
    layer0_outputs(173) <= not((inputs(180)) and (inputs(180)));
    layer0_outputs(174) <= not(inputs(86));
    layer0_outputs(175) <= (inputs(231)) and not (inputs(123));
    layer0_outputs(176) <= (inputs(35)) or (inputs(108));
    layer0_outputs(177) <= not((inputs(20)) or (inputs(162)));
    layer0_outputs(178) <= not((inputs(203)) or (inputs(72)));
    layer0_outputs(179) <= not((inputs(169)) or (inputs(126)));
    layer0_outputs(180) <= (inputs(28)) or (inputs(162));
    layer0_outputs(181) <= (inputs(187)) or (inputs(97));
    layer0_outputs(182) <= (inputs(183)) xor (inputs(186));
    layer0_outputs(183) <= not(inputs(219)) or (inputs(6));
    layer0_outputs(184) <= (inputs(120)) and not (inputs(180));
    layer0_outputs(185) <= (inputs(68)) or (inputs(128));
    layer0_outputs(186) <= (inputs(123)) xor (inputs(145));
    layer0_outputs(187) <= (inputs(99)) and (inputs(189));
    layer0_outputs(188) <= not(inputs(210));
    layer0_outputs(189) <= not((inputs(249)) or (inputs(247)));
    layer0_outputs(190) <= inputs(8);
    layer0_outputs(191) <= (inputs(189)) or (inputs(196));
    layer0_outputs(192) <= not(inputs(57)) or (inputs(101));
    layer0_outputs(193) <= inputs(103);
    layer0_outputs(194) <= not(inputs(19));
    layer0_outputs(195) <= inputs(135);
    layer0_outputs(196) <= (inputs(211)) xor (inputs(100));
    layer0_outputs(197) <= not(inputs(179));
    layer0_outputs(198) <= inputs(142);
    layer0_outputs(199) <= inputs(213);
    layer0_outputs(200) <= (inputs(239)) xor (inputs(123));
    layer0_outputs(201) <= not((inputs(6)) xor (inputs(190)));
    layer0_outputs(202) <= '1';
    layer0_outputs(203) <= (inputs(20)) or (inputs(163));
    layer0_outputs(204) <= (inputs(113)) or (inputs(51));
    layer0_outputs(205) <= not((inputs(110)) and (inputs(87)));
    layer0_outputs(206) <= not((inputs(62)) xor (inputs(248)));
    layer0_outputs(207) <= not((inputs(72)) or (inputs(140)));
    layer0_outputs(208) <= (inputs(122)) and not (inputs(203));
    layer0_outputs(209) <= inputs(174);
    layer0_outputs(210) <= not((inputs(140)) xor (inputs(66)));
    layer0_outputs(211) <= not(inputs(86)) or (inputs(90));
    layer0_outputs(212) <= not((inputs(70)) or (inputs(132)));
    layer0_outputs(213) <= not(inputs(136));
    layer0_outputs(214) <= not((inputs(168)) xor (inputs(246)));
    layer0_outputs(215) <= inputs(229);
    layer0_outputs(216) <= not(inputs(211));
    layer0_outputs(217) <= not((inputs(232)) xor (inputs(168)));
    layer0_outputs(218) <= not((inputs(26)) or (inputs(74)));
    layer0_outputs(219) <= inputs(145);
    layer0_outputs(220) <= not(inputs(25));
    layer0_outputs(221) <= not((inputs(202)) xor (inputs(80)));
    layer0_outputs(222) <= (inputs(200)) and (inputs(16));
    layer0_outputs(223) <= not(inputs(78));
    layer0_outputs(224) <= not(inputs(41));
    layer0_outputs(225) <= not(inputs(131));
    layer0_outputs(226) <= not((inputs(94)) or (inputs(95)));
    layer0_outputs(227) <= inputs(103);
    layer0_outputs(228) <= not(inputs(252));
    layer0_outputs(229) <= not((inputs(99)) or (inputs(80)));
    layer0_outputs(230) <= not((inputs(110)) or (inputs(115)));
    layer0_outputs(231) <= not(inputs(234));
    layer0_outputs(232) <= (inputs(41)) and not (inputs(164));
    layer0_outputs(233) <= not(inputs(119));
    layer0_outputs(234) <= (inputs(179)) or (inputs(63));
    layer0_outputs(235) <= not(inputs(60)) or (inputs(118));
    layer0_outputs(236) <= inputs(26);
    layer0_outputs(237) <= not(inputs(136));
    layer0_outputs(238) <= not((inputs(11)) or (inputs(20)));
    layer0_outputs(239) <= not((inputs(157)) xor (inputs(108)));
    layer0_outputs(240) <= not(inputs(2)) or (inputs(112));
    layer0_outputs(241) <= inputs(54);
    layer0_outputs(242) <= not((inputs(80)) or (inputs(46)));
    layer0_outputs(243) <= (inputs(238)) and (inputs(111));
    layer0_outputs(244) <= inputs(164);
    layer0_outputs(245) <= not(inputs(150));
    layer0_outputs(246) <= (inputs(195)) and not (inputs(170));
    layer0_outputs(247) <= (inputs(177)) or (inputs(161));
    layer0_outputs(248) <= not((inputs(115)) or (inputs(11)));
    layer0_outputs(249) <= inputs(148);
    layer0_outputs(250) <= not((inputs(7)) or (inputs(53)));
    layer0_outputs(251) <= not((inputs(225)) or (inputs(106)));
    layer0_outputs(252) <= (inputs(245)) or (inputs(4));
    layer0_outputs(253) <= inputs(167);
    layer0_outputs(254) <= not((inputs(16)) or (inputs(17)));
    layer0_outputs(255) <= (inputs(169)) xor (inputs(44));
    layer0_outputs(256) <= (inputs(155)) or (inputs(45));
    layer0_outputs(257) <= not(inputs(58)) or (inputs(193));
    layer0_outputs(258) <= (inputs(80)) or (inputs(229));
    layer0_outputs(259) <= not(inputs(226));
    layer0_outputs(260) <= inputs(102);
    layer0_outputs(261) <= inputs(91);
    layer0_outputs(262) <= not((inputs(236)) xor (inputs(135)));
    layer0_outputs(263) <= inputs(212);
    layer0_outputs(264) <= not(inputs(233)) or (inputs(95));
    layer0_outputs(265) <= (inputs(74)) or (inputs(60));
    layer0_outputs(266) <= not(inputs(44));
    layer0_outputs(267) <= (inputs(57)) or (inputs(46));
    layer0_outputs(268) <= (inputs(251)) or (inputs(209));
    layer0_outputs(269) <= not(inputs(114));
    layer0_outputs(270) <= (inputs(99)) and not (inputs(126));
    layer0_outputs(271) <= not((inputs(39)) xor (inputs(85)));
    layer0_outputs(272) <= not((inputs(146)) xor (inputs(116)));
    layer0_outputs(273) <= not((inputs(183)) xor (inputs(191)));
    layer0_outputs(274) <= inputs(86);
    layer0_outputs(275) <= not(inputs(188));
    layer0_outputs(276) <= not((inputs(169)) or (inputs(82)));
    layer0_outputs(277) <= (inputs(138)) xor (inputs(223));
    layer0_outputs(278) <= inputs(192);
    layer0_outputs(279) <= not(inputs(1));
    layer0_outputs(280) <= (inputs(146)) or (inputs(65));
    layer0_outputs(281) <= not(inputs(198));
    layer0_outputs(282) <= (inputs(184)) or (inputs(252));
    layer0_outputs(283) <= not(inputs(81)) or (inputs(255));
    layer0_outputs(284) <= not(inputs(121)) or (inputs(99));
    layer0_outputs(285) <= not(inputs(6));
    layer0_outputs(286) <= not(inputs(20));
    layer0_outputs(287) <= (inputs(160)) and (inputs(102));
    layer0_outputs(288) <= not((inputs(109)) and (inputs(227)));
    layer0_outputs(289) <= not((inputs(146)) xor (inputs(133)));
    layer0_outputs(290) <= inputs(106);
    layer0_outputs(291) <= (inputs(201)) and not (inputs(51));
    layer0_outputs(292) <= not(inputs(125));
    layer0_outputs(293) <= (inputs(4)) and (inputs(81));
    layer0_outputs(294) <= '1';
    layer0_outputs(295) <= inputs(144);
    layer0_outputs(296) <= not(inputs(155)) or (inputs(89));
    layer0_outputs(297) <= not((inputs(229)) xor (inputs(145)));
    layer0_outputs(298) <= (inputs(67)) and not (inputs(151));
    layer0_outputs(299) <= not((inputs(178)) xor (inputs(181)));
    layer0_outputs(300) <= not(inputs(22));
    layer0_outputs(301) <= inputs(201);
    layer0_outputs(302) <= (inputs(173)) xor (inputs(51));
    layer0_outputs(303) <= not(inputs(228));
    layer0_outputs(304) <= not(inputs(233)) or (inputs(111));
    layer0_outputs(305) <= (inputs(126)) and not (inputs(112));
    layer0_outputs(306) <= not(inputs(63));
    layer0_outputs(307) <= not(inputs(194));
    layer0_outputs(308) <= not(inputs(183));
    layer0_outputs(309) <= not(inputs(248));
    layer0_outputs(310) <= inputs(120);
    layer0_outputs(311) <= not((inputs(45)) xor (inputs(223)));
    layer0_outputs(312) <= not(inputs(234));
    layer0_outputs(313) <= not(inputs(165));
    layer0_outputs(314) <= not((inputs(154)) xor (inputs(249)));
    layer0_outputs(315) <= not((inputs(61)) xor (inputs(150)));
    layer0_outputs(316) <= not(inputs(60));
    layer0_outputs(317) <= not((inputs(255)) or (inputs(147)));
    layer0_outputs(318) <= '1';
    layer0_outputs(319) <= (inputs(187)) and not (inputs(70));
    layer0_outputs(320) <= (inputs(233)) and not (inputs(191));
    layer0_outputs(321) <= inputs(26);
    layer0_outputs(322) <= not((inputs(179)) or (inputs(219)));
    layer0_outputs(323) <= not(inputs(233)) or (inputs(216));
    layer0_outputs(324) <= (inputs(67)) and not (inputs(108));
    layer0_outputs(325) <= (inputs(54)) or (inputs(102));
    layer0_outputs(326) <= not(inputs(84));
    layer0_outputs(327) <= (inputs(234)) or (inputs(149));
    layer0_outputs(328) <= not(inputs(227)) or (inputs(253));
    layer0_outputs(329) <= (inputs(192)) and not (inputs(8));
    layer0_outputs(330) <= (inputs(223)) and not (inputs(1));
    layer0_outputs(331) <= not((inputs(196)) or (inputs(227)));
    layer0_outputs(332) <= inputs(108);
    layer0_outputs(333) <= not(inputs(210));
    layer0_outputs(334) <= '1';
    layer0_outputs(335) <= (inputs(118)) and (inputs(86));
    layer0_outputs(336) <= inputs(208);
    layer0_outputs(337) <= (inputs(197)) or (inputs(11));
    layer0_outputs(338) <= not((inputs(84)) and (inputs(142)));
    layer0_outputs(339) <= (inputs(37)) xor (inputs(87));
    layer0_outputs(340) <= not((inputs(27)) xor (inputs(50)));
    layer0_outputs(341) <= inputs(178);
    layer0_outputs(342) <= (inputs(159)) xor (inputs(54));
    layer0_outputs(343) <= not(inputs(18));
    layer0_outputs(344) <= not((inputs(5)) xor (inputs(101)));
    layer0_outputs(345) <= (inputs(12)) and not (inputs(243));
    layer0_outputs(346) <= inputs(178);
    layer0_outputs(347) <= inputs(224);
    layer0_outputs(348) <= inputs(147);
    layer0_outputs(349) <= (inputs(248)) and (inputs(138));
    layer0_outputs(350) <= inputs(124);
    layer0_outputs(351) <= inputs(212);
    layer0_outputs(352) <= not(inputs(134)) or (inputs(139));
    layer0_outputs(353) <= (inputs(53)) xor (inputs(203));
    layer0_outputs(354) <= inputs(193);
    layer0_outputs(355) <= inputs(162);
    layer0_outputs(356) <= not(inputs(58)) or (inputs(183));
    layer0_outputs(357) <= not(inputs(168));
    layer0_outputs(358) <= not((inputs(8)) or (inputs(94)));
    layer0_outputs(359) <= not((inputs(112)) or (inputs(114)));
    layer0_outputs(360) <= (inputs(17)) or (inputs(19));
    layer0_outputs(361) <= not(inputs(10));
    layer0_outputs(362) <= not((inputs(164)) or (inputs(71)));
    layer0_outputs(363) <= inputs(236);
    layer0_outputs(364) <= '1';
    layer0_outputs(365) <= (inputs(14)) or (inputs(190));
    layer0_outputs(366) <= not((inputs(11)) xor (inputs(10)));
    layer0_outputs(367) <= not(inputs(160));
    layer0_outputs(368) <= (inputs(13)) and not (inputs(47));
    layer0_outputs(369) <= not((inputs(77)) or (inputs(24)));
    layer0_outputs(370) <= inputs(158);
    layer0_outputs(371) <= not(inputs(166)) or (inputs(118));
    layer0_outputs(372) <= not((inputs(185)) xor (inputs(163)));
    layer0_outputs(373) <= not(inputs(246));
    layer0_outputs(374) <= not(inputs(152)) or (inputs(219));
    layer0_outputs(375) <= inputs(20);
    layer0_outputs(376) <= not(inputs(230));
    layer0_outputs(377) <= not((inputs(22)) or (inputs(51)));
    layer0_outputs(378) <= not(inputs(157)) or (inputs(160));
    layer0_outputs(379) <= (inputs(143)) xor (inputs(62));
    layer0_outputs(380) <= not(inputs(41));
    layer0_outputs(381) <= inputs(168);
    layer0_outputs(382) <= not(inputs(110));
    layer0_outputs(383) <= (inputs(4)) xor (inputs(91));
    layer0_outputs(384) <= (inputs(188)) and not (inputs(83));
    layer0_outputs(385) <= inputs(43);
    layer0_outputs(386) <= not(inputs(174));
    layer0_outputs(387) <= (inputs(95)) xor (inputs(91));
    layer0_outputs(388) <= (inputs(73)) xor (inputs(208));
    layer0_outputs(389) <= not(inputs(168));
    layer0_outputs(390) <= not(inputs(212)) or (inputs(239));
    layer0_outputs(391) <= not(inputs(26));
    layer0_outputs(392) <= not((inputs(176)) xor (inputs(63)));
    layer0_outputs(393) <= not(inputs(112)) or (inputs(235));
    layer0_outputs(394) <= not(inputs(80));
    layer0_outputs(395) <= (inputs(57)) or (inputs(136));
    layer0_outputs(396) <= not((inputs(94)) or (inputs(103)));
    layer0_outputs(397) <= not(inputs(105));
    layer0_outputs(398) <= (inputs(170)) and not (inputs(5));
    layer0_outputs(399) <= (inputs(184)) and not (inputs(191));
    layer0_outputs(400) <= not(inputs(85)) or (inputs(16));
    layer0_outputs(401) <= inputs(125);
    layer0_outputs(402) <= inputs(183);
    layer0_outputs(403) <= not((inputs(77)) or (inputs(24)));
    layer0_outputs(404) <= (inputs(136)) and not (inputs(168));
    layer0_outputs(405) <= inputs(203);
    layer0_outputs(406) <= not(inputs(21));
    layer0_outputs(407) <= (inputs(207)) and not (inputs(97));
    layer0_outputs(408) <= not((inputs(223)) or (inputs(211)));
    layer0_outputs(409) <= not(inputs(211)) or (inputs(125));
    layer0_outputs(410) <= (inputs(91)) xor (inputs(18));
    layer0_outputs(411) <= (inputs(169)) xor (inputs(138));
    layer0_outputs(412) <= not((inputs(228)) or (inputs(127)));
    layer0_outputs(413) <= not(inputs(44)) or (inputs(205));
    layer0_outputs(414) <= '1';
    layer0_outputs(415) <= not((inputs(82)) or (inputs(121)));
    layer0_outputs(416) <= inputs(167);
    layer0_outputs(417) <= not(inputs(38));
    layer0_outputs(418) <= inputs(186);
    layer0_outputs(419) <= not(inputs(215)) or (inputs(31));
    layer0_outputs(420) <= inputs(167);
    layer0_outputs(421) <= not(inputs(150)) or (inputs(60));
    layer0_outputs(422) <= (inputs(182)) or (inputs(89));
    layer0_outputs(423) <= (inputs(77)) xor (inputs(71));
    layer0_outputs(424) <= inputs(19);
    layer0_outputs(425) <= (inputs(254)) or (inputs(131));
    layer0_outputs(426) <= not(inputs(18)) or (inputs(80));
    layer0_outputs(427) <= not((inputs(65)) xor (inputs(199)));
    layer0_outputs(428) <= (inputs(214)) and not (inputs(152));
    layer0_outputs(429) <= not((inputs(174)) or (inputs(183)));
    layer0_outputs(430) <= not(inputs(213));
    layer0_outputs(431) <= not(inputs(226)) or (inputs(94));
    layer0_outputs(432) <= not((inputs(8)) or (inputs(33)));
    layer0_outputs(433) <= inputs(14);
    layer0_outputs(434) <= not((inputs(221)) or (inputs(42)));
    layer0_outputs(435) <= (inputs(19)) or (inputs(74));
    layer0_outputs(436) <= (inputs(180)) and not (inputs(166));
    layer0_outputs(437) <= not((inputs(188)) or (inputs(79)));
    layer0_outputs(438) <= (inputs(141)) and not (inputs(214));
    layer0_outputs(439) <= not(inputs(134)) or (inputs(57));
    layer0_outputs(440) <= '0';
    layer0_outputs(441) <= inputs(194);
    layer0_outputs(442) <= inputs(165);
    layer0_outputs(443) <= inputs(251);
    layer0_outputs(444) <= not(inputs(83));
    layer0_outputs(445) <= not((inputs(40)) and (inputs(27)));
    layer0_outputs(446) <= not(inputs(148));
    layer0_outputs(447) <= not(inputs(144));
    layer0_outputs(448) <= (inputs(97)) or (inputs(90));
    layer0_outputs(449) <= not(inputs(223));
    layer0_outputs(450) <= not((inputs(29)) or (inputs(6)));
    layer0_outputs(451) <= (inputs(100)) and not (inputs(188));
    layer0_outputs(452) <= (inputs(231)) or (inputs(99));
    layer0_outputs(453) <= not(inputs(5)) or (inputs(49));
    layer0_outputs(454) <= (inputs(109)) and (inputs(255));
    layer0_outputs(455) <= (inputs(158)) and not (inputs(118));
    layer0_outputs(456) <= (inputs(210)) xor (inputs(67));
    layer0_outputs(457) <= not(inputs(11)) or (inputs(23));
    layer0_outputs(458) <= (inputs(167)) and not (inputs(82));
    layer0_outputs(459) <= not(inputs(18)) or (inputs(80));
    layer0_outputs(460) <= (inputs(62)) xor (inputs(249));
    layer0_outputs(461) <= not(inputs(134)) or (inputs(66));
    layer0_outputs(462) <= inputs(90);
    layer0_outputs(463) <= not(inputs(44)) or (inputs(80));
    layer0_outputs(464) <= not(inputs(142));
    layer0_outputs(465) <= not(inputs(162));
    layer0_outputs(466) <= (inputs(94)) and (inputs(96));
    layer0_outputs(467) <= inputs(228);
    layer0_outputs(468) <= (inputs(33)) or (inputs(25));
    layer0_outputs(469) <= not(inputs(232));
    layer0_outputs(470) <= not((inputs(84)) or (inputs(65)));
    layer0_outputs(471) <= not((inputs(25)) or (inputs(9)));
    layer0_outputs(472) <= inputs(99);
    layer0_outputs(473) <= inputs(182);
    layer0_outputs(474) <= inputs(75);
    layer0_outputs(475) <= (inputs(0)) and not (inputs(240));
    layer0_outputs(476) <= not(inputs(207));
    layer0_outputs(477) <= not((inputs(108)) xor (inputs(190)));
    layer0_outputs(478) <= (inputs(133)) and (inputs(149));
    layer0_outputs(479) <= not((inputs(113)) xor (inputs(172)));
    layer0_outputs(480) <= inputs(9);
    layer0_outputs(481) <= (inputs(210)) and not (inputs(185));
    layer0_outputs(482) <= not(inputs(66));
    layer0_outputs(483) <= not(inputs(86));
    layer0_outputs(484) <= inputs(21);
    layer0_outputs(485) <= (inputs(208)) or (inputs(211));
    layer0_outputs(486) <= (inputs(218)) or (inputs(67));
    layer0_outputs(487) <= inputs(54);
    layer0_outputs(488) <= not((inputs(37)) or (inputs(219)));
    layer0_outputs(489) <= '1';
    layer0_outputs(490) <= (inputs(207)) xor (inputs(173));
    layer0_outputs(491) <= not((inputs(35)) or (inputs(29)));
    layer0_outputs(492) <= (inputs(117)) or (inputs(132));
    layer0_outputs(493) <= not(inputs(7)) or (inputs(179));
    layer0_outputs(494) <= inputs(159);
    layer0_outputs(495) <= not((inputs(12)) and (inputs(50)));
    layer0_outputs(496) <= (inputs(102)) or (inputs(64));
    layer0_outputs(497) <= not(inputs(39)) or (inputs(161));
    layer0_outputs(498) <= (inputs(28)) and not (inputs(130));
    layer0_outputs(499) <= not((inputs(193)) xor (inputs(189)));
    layer0_outputs(500) <= inputs(7);
    layer0_outputs(501) <= (inputs(65)) xor (inputs(192));
    layer0_outputs(502) <= (inputs(189)) or (inputs(158));
    layer0_outputs(503) <= inputs(163);
    layer0_outputs(504) <= inputs(61);
    layer0_outputs(505) <= not((inputs(92)) or (inputs(88)));
    layer0_outputs(506) <= (inputs(111)) or (inputs(4));
    layer0_outputs(507) <= not(inputs(27));
    layer0_outputs(508) <= not((inputs(49)) xor (inputs(2)));
    layer0_outputs(509) <= not(inputs(245));
    layer0_outputs(510) <= (inputs(144)) xor (inputs(230));
    layer0_outputs(511) <= inputs(25);
    layer0_outputs(512) <= not(inputs(234));
    layer0_outputs(513) <= inputs(196);
    layer0_outputs(514) <= not((inputs(187)) or (inputs(52)));
    layer0_outputs(515) <= (inputs(23)) or (inputs(216));
    layer0_outputs(516) <= (inputs(211)) and not (inputs(98));
    layer0_outputs(517) <= inputs(222);
    layer0_outputs(518) <= inputs(162);
    layer0_outputs(519) <= inputs(102);
    layer0_outputs(520) <= inputs(236);
    layer0_outputs(521) <= not(inputs(103));
    layer0_outputs(522) <= not(inputs(153)) or (inputs(66));
    layer0_outputs(523) <= (inputs(139)) or (inputs(237));
    layer0_outputs(524) <= inputs(118);
    layer0_outputs(525) <= not(inputs(34));
    layer0_outputs(526) <= not(inputs(205)) or (inputs(125));
    layer0_outputs(527) <= not((inputs(89)) xor (inputs(185)));
    layer0_outputs(528) <= (inputs(248)) or (inputs(134));
    layer0_outputs(529) <= (inputs(10)) and not (inputs(86));
    layer0_outputs(530) <= not(inputs(26)) or (inputs(193));
    layer0_outputs(531) <= not(inputs(168)) or (inputs(243));
    layer0_outputs(532) <= not((inputs(204)) xor (inputs(195)));
    layer0_outputs(533) <= (inputs(215)) and (inputs(196));
    layer0_outputs(534) <= (inputs(217)) xor (inputs(134));
    layer0_outputs(535) <= not((inputs(245)) or (inputs(219)));
    layer0_outputs(536) <= (inputs(42)) or (inputs(178));
    layer0_outputs(537) <= not(inputs(27)) or (inputs(206));
    layer0_outputs(538) <= (inputs(21)) or (inputs(94));
    layer0_outputs(539) <= inputs(10);
    layer0_outputs(540) <= inputs(247);
    layer0_outputs(541) <= not(inputs(174)) or (inputs(231));
    layer0_outputs(542) <= inputs(200);
    layer0_outputs(543) <= inputs(234);
    layer0_outputs(544) <= not(inputs(11)) or (inputs(81));
    layer0_outputs(545) <= not(inputs(169));
    layer0_outputs(546) <= (inputs(131)) xor (inputs(65));
    layer0_outputs(547) <= not(inputs(21));
    layer0_outputs(548) <= (inputs(165)) or (inputs(80));
    layer0_outputs(549) <= not((inputs(134)) xor (inputs(107)));
    layer0_outputs(550) <= (inputs(39)) or (inputs(76));
    layer0_outputs(551) <= (inputs(27)) xor (inputs(9));
    layer0_outputs(552) <= not((inputs(34)) or (inputs(226)));
    layer0_outputs(553) <= (inputs(223)) or (inputs(103));
    layer0_outputs(554) <= inputs(76);
    layer0_outputs(555) <= not(inputs(27));
    layer0_outputs(556) <= not(inputs(6)) or (inputs(232));
    layer0_outputs(557) <= (inputs(181)) or (inputs(195));
    layer0_outputs(558) <= inputs(152);
    layer0_outputs(559) <= not(inputs(116));
    layer0_outputs(560) <= (inputs(15)) or (inputs(245));
    layer0_outputs(561) <= (inputs(114)) or (inputs(121));
    layer0_outputs(562) <= not((inputs(95)) or (inputs(181)));
    layer0_outputs(563) <= not((inputs(110)) xor (inputs(35)));
    layer0_outputs(564) <= (inputs(42)) and not (inputs(130));
    layer0_outputs(565) <= (inputs(99)) and not (inputs(0));
    layer0_outputs(566) <= not(inputs(41));
    layer0_outputs(567) <= (inputs(68)) and not (inputs(206));
    layer0_outputs(568) <= not(inputs(211)) or (inputs(97));
    layer0_outputs(569) <= '0';
    layer0_outputs(570) <= not(inputs(181));
    layer0_outputs(571) <= inputs(110);
    layer0_outputs(572) <= (inputs(214)) or (inputs(196));
    layer0_outputs(573) <= not(inputs(193)) or (inputs(4));
    layer0_outputs(574) <= (inputs(215)) or (inputs(1));
    layer0_outputs(575) <= not(inputs(92)) or (inputs(242));
    layer0_outputs(576) <= (inputs(194)) or (inputs(168));
    layer0_outputs(577) <= (inputs(16)) xor (inputs(252));
    layer0_outputs(578) <= '1';
    layer0_outputs(579) <= not((inputs(120)) xor (inputs(88)));
    layer0_outputs(580) <= not(inputs(77)) or (inputs(82));
    layer0_outputs(581) <= inputs(136);
    layer0_outputs(582) <= (inputs(190)) or (inputs(15));
    layer0_outputs(583) <= not(inputs(140));
    layer0_outputs(584) <= not(inputs(69)) or (inputs(79));
    layer0_outputs(585) <= not((inputs(36)) xor (inputs(174)));
    layer0_outputs(586) <= not((inputs(249)) or (inputs(206)));
    layer0_outputs(587) <= not(inputs(66));
    layer0_outputs(588) <= not((inputs(114)) or (inputs(97)));
    layer0_outputs(589) <= not(inputs(91)) or (inputs(144));
    layer0_outputs(590) <= not(inputs(83)) or (inputs(253));
    layer0_outputs(591) <= (inputs(52)) or (inputs(235));
    layer0_outputs(592) <= (inputs(220)) and not (inputs(14));
    layer0_outputs(593) <= not(inputs(90)) or (inputs(111));
    layer0_outputs(594) <= not(inputs(213)) or (inputs(87));
    layer0_outputs(595) <= not(inputs(198)) or (inputs(1));
    layer0_outputs(596) <= inputs(58);
    layer0_outputs(597) <= (inputs(20)) or (inputs(59));
    layer0_outputs(598) <= inputs(16);
    layer0_outputs(599) <= inputs(23);
    layer0_outputs(600) <= not(inputs(248));
    layer0_outputs(601) <= not((inputs(43)) and (inputs(124)));
    layer0_outputs(602) <= (inputs(1)) and (inputs(78));
    layer0_outputs(603) <= (inputs(228)) and not (inputs(34));
    layer0_outputs(604) <= (inputs(96)) xor (inputs(176));
    layer0_outputs(605) <= not(inputs(59));
    layer0_outputs(606) <= inputs(162);
    layer0_outputs(607) <= (inputs(189)) and not (inputs(15));
    layer0_outputs(608) <= (inputs(186)) or (inputs(103));
    layer0_outputs(609) <= (inputs(18)) and not (inputs(61));
    layer0_outputs(610) <= (inputs(163)) and not (inputs(143));
    layer0_outputs(611) <= not(inputs(169)) or (inputs(245));
    layer0_outputs(612) <= not(inputs(101)) or (inputs(145));
    layer0_outputs(613) <= not((inputs(229)) and (inputs(36)));
    layer0_outputs(614) <= inputs(115);
    layer0_outputs(615) <= not(inputs(162));
    layer0_outputs(616) <= not((inputs(205)) or (inputs(148)));
    layer0_outputs(617) <= not((inputs(98)) or (inputs(100)));
    layer0_outputs(618) <= '0';
    layer0_outputs(619) <= not((inputs(243)) xor (inputs(230)));
    layer0_outputs(620) <= not((inputs(239)) or (inputs(244)));
    layer0_outputs(621) <= not((inputs(110)) xor (inputs(49)));
    layer0_outputs(622) <= inputs(226);
    layer0_outputs(623) <= not((inputs(242)) and (inputs(162)));
    layer0_outputs(624) <= not(inputs(167)) or (inputs(51));
    layer0_outputs(625) <= inputs(47);
    layer0_outputs(626) <= inputs(179);
    layer0_outputs(627) <= inputs(116);
    layer0_outputs(628) <= not((inputs(167)) or (inputs(34)));
    layer0_outputs(629) <= not((inputs(9)) or (inputs(1)));
    layer0_outputs(630) <= inputs(70);
    layer0_outputs(631) <= (inputs(16)) or (inputs(192));
    layer0_outputs(632) <= (inputs(203)) xor (inputs(183));
    layer0_outputs(633) <= not((inputs(230)) or (inputs(195)));
    layer0_outputs(634) <= not(inputs(122)) or (inputs(1));
    layer0_outputs(635) <= (inputs(161)) or (inputs(74));
    layer0_outputs(636) <= inputs(33);
    layer0_outputs(637) <= not((inputs(79)) and (inputs(216)));
    layer0_outputs(638) <= not((inputs(229)) xor (inputs(163)));
    layer0_outputs(639) <= not(inputs(38));
    layer0_outputs(640) <= not((inputs(125)) xor (inputs(176)));
    layer0_outputs(641) <= not(inputs(148));
    layer0_outputs(642) <= (inputs(122)) or (inputs(96));
    layer0_outputs(643) <= (inputs(133)) or (inputs(212));
    layer0_outputs(644) <= inputs(60);
    layer0_outputs(645) <= not((inputs(88)) and (inputs(199)));
    layer0_outputs(646) <= not((inputs(151)) or (inputs(14)));
    layer0_outputs(647) <= (inputs(141)) and not (inputs(80));
    layer0_outputs(648) <= (inputs(81)) and not (inputs(224));
    layer0_outputs(649) <= inputs(247);
    layer0_outputs(650) <= not(inputs(27)) or (inputs(220));
    layer0_outputs(651) <= not((inputs(103)) or (inputs(237)));
    layer0_outputs(652) <= not((inputs(98)) or (inputs(182)));
    layer0_outputs(653) <= not(inputs(98));
    layer0_outputs(654) <= not((inputs(247)) or (inputs(230)));
    layer0_outputs(655) <= (inputs(185)) and not (inputs(222));
    layer0_outputs(656) <= not((inputs(199)) or (inputs(171)));
    layer0_outputs(657) <= not((inputs(87)) or (inputs(136)));
    layer0_outputs(658) <= inputs(245);
    layer0_outputs(659) <= inputs(185);
    layer0_outputs(660) <= inputs(25);
    layer0_outputs(661) <= not(inputs(224));
    layer0_outputs(662) <= not(inputs(46));
    layer0_outputs(663) <= inputs(82);
    layer0_outputs(664) <= not(inputs(7));
    layer0_outputs(665) <= (inputs(245)) xor (inputs(97));
    layer0_outputs(666) <= not((inputs(68)) or (inputs(5)));
    layer0_outputs(667) <= inputs(100);
    layer0_outputs(668) <= (inputs(149)) xor (inputs(50));
    layer0_outputs(669) <= inputs(60);
    layer0_outputs(670) <= (inputs(143)) or (inputs(33));
    layer0_outputs(671) <= (inputs(205)) xor (inputs(144));
    layer0_outputs(672) <= (inputs(181)) and not (inputs(96));
    layer0_outputs(673) <= (inputs(92)) or (inputs(242));
    layer0_outputs(674) <= not(inputs(98)) or (inputs(49));
    layer0_outputs(675) <= not((inputs(168)) or (inputs(255)));
    layer0_outputs(676) <= not(inputs(126)) or (inputs(225));
    layer0_outputs(677) <= inputs(158);
    layer0_outputs(678) <= not(inputs(214)) or (inputs(34));
    layer0_outputs(679) <= not((inputs(132)) and (inputs(154)));
    layer0_outputs(680) <= (inputs(168)) and not (inputs(47));
    layer0_outputs(681) <= inputs(106);
    layer0_outputs(682) <= not(inputs(115));
    layer0_outputs(683) <= (inputs(191)) or (inputs(201));
    layer0_outputs(684) <= not((inputs(160)) or (inputs(243)));
    layer0_outputs(685) <= not(inputs(75)) or (inputs(222));
    layer0_outputs(686) <= inputs(193);
    layer0_outputs(687) <= (inputs(43)) or (inputs(138));
    layer0_outputs(688) <= not((inputs(139)) xor (inputs(79)));
    layer0_outputs(689) <= '1';
    layer0_outputs(690) <= (inputs(68)) or (inputs(97));
    layer0_outputs(691) <= (inputs(4)) xor (inputs(141));
    layer0_outputs(692) <= not((inputs(55)) or (inputs(22)));
    layer0_outputs(693) <= (inputs(17)) or (inputs(163));
    layer0_outputs(694) <= inputs(82);
    layer0_outputs(695) <= (inputs(10)) xor (inputs(22));
    layer0_outputs(696) <= (inputs(243)) or (inputs(240));
    layer0_outputs(697) <= not(inputs(75));
    layer0_outputs(698) <= (inputs(153)) or (inputs(205));
    layer0_outputs(699) <= (inputs(100)) and not (inputs(20));
    layer0_outputs(700) <= inputs(174);
    layer0_outputs(701) <= (inputs(36)) or (inputs(91));
    layer0_outputs(702) <= not(inputs(150));
    layer0_outputs(703) <= not(inputs(68));
    layer0_outputs(704) <= not(inputs(29));
    layer0_outputs(705) <= not(inputs(129));
    layer0_outputs(706) <= (inputs(24)) or (inputs(39));
    layer0_outputs(707) <= (inputs(192)) and not (inputs(142));
    layer0_outputs(708) <= not(inputs(104)) or (inputs(16));
    layer0_outputs(709) <= inputs(41);
    layer0_outputs(710) <= (inputs(132)) or (inputs(15));
    layer0_outputs(711) <= (inputs(2)) or (inputs(31));
    layer0_outputs(712) <= not(inputs(117)) or (inputs(62));
    layer0_outputs(713) <= (inputs(28)) xor (inputs(192));
    layer0_outputs(714) <= (inputs(42)) or (inputs(7));
    layer0_outputs(715) <= '0';
    layer0_outputs(716) <= (inputs(105)) and (inputs(26));
    layer0_outputs(717) <= (inputs(122)) and not (inputs(96));
    layer0_outputs(718) <= inputs(187);
    layer0_outputs(719) <= not(inputs(65));
    layer0_outputs(720) <= not((inputs(239)) or (inputs(255)));
    layer0_outputs(721) <= (inputs(203)) and (inputs(111));
    layer0_outputs(722) <= inputs(184);
    layer0_outputs(723) <= (inputs(39)) and not (inputs(33));
    layer0_outputs(724) <= not(inputs(61)) or (inputs(69));
    layer0_outputs(725) <= not(inputs(216));
    layer0_outputs(726) <= not(inputs(228));
    layer0_outputs(727) <= (inputs(84)) and not (inputs(91));
    layer0_outputs(728) <= not(inputs(84));
    layer0_outputs(729) <= not(inputs(228)) or (inputs(89));
    layer0_outputs(730) <= (inputs(204)) or (inputs(205));
    layer0_outputs(731) <= not(inputs(63));
    layer0_outputs(732) <= not((inputs(75)) or (inputs(112)));
    layer0_outputs(733) <= (inputs(38)) and not (inputs(156));
    layer0_outputs(734) <= not(inputs(87));
    layer0_outputs(735) <= (inputs(107)) and (inputs(123));
    layer0_outputs(736) <= not(inputs(199));
    layer0_outputs(737) <= (inputs(30)) and (inputs(87));
    layer0_outputs(738) <= not(inputs(63)) or (inputs(38));
    layer0_outputs(739) <= (inputs(173)) xor (inputs(232));
    layer0_outputs(740) <= (inputs(134)) and not (inputs(109));
    layer0_outputs(741) <= not((inputs(91)) or (inputs(104)));
    layer0_outputs(742) <= not((inputs(179)) xor (inputs(209)));
    layer0_outputs(743) <= (inputs(146)) or (inputs(39));
    layer0_outputs(744) <= inputs(173);
    layer0_outputs(745) <= (inputs(240)) and (inputs(81));
    layer0_outputs(746) <= inputs(130);
    layer0_outputs(747) <= (inputs(203)) and (inputs(75));
    layer0_outputs(748) <= (inputs(133)) and not (inputs(189));
    layer0_outputs(749) <= (inputs(240)) or (inputs(24));
    layer0_outputs(750) <= (inputs(25)) or (inputs(105));
    layer0_outputs(751) <= not((inputs(233)) or (inputs(51)));
    layer0_outputs(752) <= not(inputs(146)) or (inputs(71));
    layer0_outputs(753) <= inputs(23);
    layer0_outputs(754) <= inputs(162);
    layer0_outputs(755) <= not(inputs(39));
    layer0_outputs(756) <= not((inputs(165)) xor (inputs(203)));
    layer0_outputs(757) <= inputs(66);
    layer0_outputs(758) <= not((inputs(161)) xor (inputs(25)));
    layer0_outputs(759) <= not(inputs(164));
    layer0_outputs(760) <= (inputs(255)) or (inputs(38));
    layer0_outputs(761) <= not(inputs(199)) or (inputs(192));
    layer0_outputs(762) <= inputs(246);
    layer0_outputs(763) <= (inputs(119)) and (inputs(43));
    layer0_outputs(764) <= not(inputs(28));
    layer0_outputs(765) <= not(inputs(229));
    layer0_outputs(766) <= inputs(59);
    layer0_outputs(767) <= not((inputs(154)) and (inputs(182)));
    layer0_outputs(768) <= (inputs(205)) or (inputs(221));
    layer0_outputs(769) <= not((inputs(53)) xor (inputs(36)));
    layer0_outputs(770) <= not(inputs(162));
    layer0_outputs(771) <= inputs(66);
    layer0_outputs(772) <= (inputs(65)) xor (inputs(83));
    layer0_outputs(773) <= (inputs(241)) or (inputs(120));
    layer0_outputs(774) <= not((inputs(16)) xor (inputs(174)));
    layer0_outputs(775) <= (inputs(149)) xor (inputs(224));
    layer0_outputs(776) <= (inputs(39)) xor (inputs(248));
    layer0_outputs(777) <= not(inputs(179));
    layer0_outputs(778) <= '1';
    layer0_outputs(779) <= not(inputs(51));
    layer0_outputs(780) <= not((inputs(54)) and (inputs(72)));
    layer0_outputs(781) <= not((inputs(250)) xor (inputs(242)));
    layer0_outputs(782) <= not(inputs(216)) or (inputs(49));
    layer0_outputs(783) <= inputs(197);
    layer0_outputs(784) <= inputs(181);
    layer0_outputs(785) <= not(inputs(98));
    layer0_outputs(786) <= inputs(230);
    layer0_outputs(787) <= inputs(94);
    layer0_outputs(788) <= not(inputs(67));
    layer0_outputs(789) <= not(inputs(187));
    layer0_outputs(790) <= inputs(163);
    layer0_outputs(791) <= inputs(245);
    layer0_outputs(792) <= (inputs(175)) or (inputs(195));
    layer0_outputs(793) <= (inputs(210)) or (inputs(197));
    layer0_outputs(794) <= not(inputs(146));
    layer0_outputs(795) <= (inputs(121)) and not (inputs(194));
    layer0_outputs(796) <= not((inputs(40)) and (inputs(31)));
    layer0_outputs(797) <= (inputs(68)) and not (inputs(196));
    layer0_outputs(798) <= not(inputs(183)) or (inputs(46));
    layer0_outputs(799) <= (inputs(78)) or (inputs(90));
    layer0_outputs(800) <= (inputs(153)) and not (inputs(0));
    layer0_outputs(801) <= not(inputs(124));
    layer0_outputs(802) <= (inputs(230)) and not (inputs(96));
    layer0_outputs(803) <= not((inputs(89)) xor (inputs(10)));
    layer0_outputs(804) <= (inputs(92)) xor (inputs(48));
    layer0_outputs(805) <= not((inputs(227)) or (inputs(56)));
    layer0_outputs(806) <= inputs(230);
    layer0_outputs(807) <= (inputs(74)) xor (inputs(60));
    layer0_outputs(808) <= (inputs(229)) xor (inputs(235));
    layer0_outputs(809) <= not(inputs(52));
    layer0_outputs(810) <= not(inputs(196));
    layer0_outputs(811) <= (inputs(219)) or (inputs(172));
    layer0_outputs(812) <= not((inputs(236)) xor (inputs(156)));
    layer0_outputs(813) <= not((inputs(129)) or (inputs(52)));
    layer0_outputs(814) <= (inputs(75)) and not (inputs(109));
    layer0_outputs(815) <= (inputs(169)) or (inputs(172));
    layer0_outputs(816) <= not((inputs(7)) or (inputs(138)));
    layer0_outputs(817) <= (inputs(188)) and not (inputs(254));
    layer0_outputs(818) <= not(inputs(231)) or (inputs(67));
    layer0_outputs(819) <= (inputs(69)) or (inputs(31));
    layer0_outputs(820) <= not((inputs(160)) or (inputs(21)));
    layer0_outputs(821) <= (inputs(152)) or (inputs(105));
    layer0_outputs(822) <= not((inputs(206)) or (inputs(64)));
    layer0_outputs(823) <= (inputs(71)) and (inputs(172));
    layer0_outputs(824) <= not((inputs(100)) or (inputs(132)));
    layer0_outputs(825) <= inputs(232);
    layer0_outputs(826) <= (inputs(7)) or (inputs(156));
    layer0_outputs(827) <= (inputs(89)) and not (inputs(0));
    layer0_outputs(828) <= not(inputs(86));
    layer0_outputs(829) <= not((inputs(13)) or (inputs(213)));
    layer0_outputs(830) <= (inputs(33)) and not (inputs(54));
    layer0_outputs(831) <= not(inputs(145)) or (inputs(240));
    layer0_outputs(832) <= not((inputs(172)) or (inputs(171)));
    layer0_outputs(833) <= not(inputs(150));
    layer0_outputs(834) <= not(inputs(255));
    layer0_outputs(835) <= inputs(210);
    layer0_outputs(836) <= not((inputs(84)) or (inputs(125)));
    layer0_outputs(837) <= not((inputs(222)) or (inputs(14)));
    layer0_outputs(838) <= not(inputs(106));
    layer0_outputs(839) <= inputs(71);
    layer0_outputs(840) <= (inputs(153)) or (inputs(242));
    layer0_outputs(841) <= (inputs(148)) and not (inputs(17));
    layer0_outputs(842) <= inputs(227);
    layer0_outputs(843) <= inputs(36);
    layer0_outputs(844) <= (inputs(92)) or (inputs(123));
    layer0_outputs(845) <= (inputs(217)) and not (inputs(137));
    layer0_outputs(846) <= not(inputs(135));
    layer0_outputs(847) <= not((inputs(63)) or (inputs(78)));
    layer0_outputs(848) <= (inputs(91)) and not (inputs(15));
    layer0_outputs(849) <= not(inputs(125));
    layer0_outputs(850) <= (inputs(240)) or (inputs(80));
    layer0_outputs(851) <= inputs(60);
    layer0_outputs(852) <= not(inputs(99));
    layer0_outputs(853) <= (inputs(37)) xor (inputs(103));
    layer0_outputs(854) <= not(inputs(193));
    layer0_outputs(855) <= not(inputs(227));
    layer0_outputs(856) <= (inputs(85)) and not (inputs(72));
    layer0_outputs(857) <= (inputs(231)) xor (inputs(192));
    layer0_outputs(858) <= not(inputs(176)) or (inputs(206));
    layer0_outputs(859) <= not(inputs(66)) or (inputs(48));
    layer0_outputs(860) <= inputs(217);
    layer0_outputs(861) <= not(inputs(72));
    layer0_outputs(862) <= (inputs(241)) and not (inputs(169));
    layer0_outputs(863) <= (inputs(160)) and not (inputs(95));
    layer0_outputs(864) <= (inputs(120)) and not (inputs(160));
    layer0_outputs(865) <= inputs(170);
    layer0_outputs(866) <= not((inputs(172)) or (inputs(98)));
    layer0_outputs(867) <= inputs(141);
    layer0_outputs(868) <= not((inputs(249)) or (inputs(149)));
    layer0_outputs(869) <= not((inputs(96)) or (inputs(108)));
    layer0_outputs(870) <= not((inputs(38)) xor (inputs(8)));
    layer0_outputs(871) <= (inputs(115)) and not (inputs(80));
    layer0_outputs(872) <= not(inputs(63));
    layer0_outputs(873) <= inputs(123);
    layer0_outputs(874) <= (inputs(5)) or (inputs(207));
    layer0_outputs(875) <= not((inputs(101)) xor (inputs(223)));
    layer0_outputs(876) <= not(inputs(130)) or (inputs(36));
    layer0_outputs(877) <= not((inputs(139)) and (inputs(200)));
    layer0_outputs(878) <= not(inputs(141));
    layer0_outputs(879) <= not(inputs(85)) or (inputs(2));
    layer0_outputs(880) <= not((inputs(213)) or (inputs(116)));
    layer0_outputs(881) <= (inputs(77)) xor (inputs(203));
    layer0_outputs(882) <= (inputs(126)) and not (inputs(32));
    layer0_outputs(883) <= not((inputs(94)) and (inputs(126)));
    layer0_outputs(884) <= (inputs(166)) or (inputs(35));
    layer0_outputs(885) <= inputs(78);
    layer0_outputs(886) <= (inputs(81)) and (inputs(110));
    layer0_outputs(887) <= (inputs(174)) or (inputs(150));
    layer0_outputs(888) <= (inputs(6)) or (inputs(108));
    layer0_outputs(889) <= (inputs(55)) xor (inputs(29));
    layer0_outputs(890) <= (inputs(8)) and not (inputs(58));
    layer0_outputs(891) <= not(inputs(64));
    layer0_outputs(892) <= not((inputs(200)) or (inputs(237)));
    layer0_outputs(893) <= not(inputs(201));
    layer0_outputs(894) <= not((inputs(239)) or (inputs(50)));
    layer0_outputs(895) <= (inputs(117)) xor (inputs(73));
    layer0_outputs(896) <= not(inputs(196)) or (inputs(140));
    layer0_outputs(897) <= not(inputs(105));
    layer0_outputs(898) <= not((inputs(3)) xor (inputs(144)));
    layer0_outputs(899) <= not(inputs(155));
    layer0_outputs(900) <= (inputs(43)) and not (inputs(146));
    layer0_outputs(901) <= inputs(93);
    layer0_outputs(902) <= (inputs(136)) or (inputs(153));
    layer0_outputs(903) <= not(inputs(69));
    layer0_outputs(904) <= inputs(58);
    layer0_outputs(905) <= not((inputs(88)) and (inputs(186)));
    layer0_outputs(906) <= not(inputs(229));
    layer0_outputs(907) <= not((inputs(138)) xor (inputs(169)));
    layer0_outputs(908) <= (inputs(73)) and not (inputs(175));
    layer0_outputs(909) <= not(inputs(202)) or (inputs(248));
    layer0_outputs(910) <= not(inputs(185));
    layer0_outputs(911) <= (inputs(34)) xor (inputs(92));
    layer0_outputs(912) <= (inputs(213)) or (inputs(229));
    layer0_outputs(913) <= inputs(228);
    layer0_outputs(914) <= not((inputs(86)) or (inputs(193)));
    layer0_outputs(915) <= not(inputs(76));
    layer0_outputs(916) <= (inputs(111)) or (inputs(253));
    layer0_outputs(917) <= not((inputs(9)) and (inputs(100)));
    layer0_outputs(918) <= inputs(95);
    layer0_outputs(919) <= inputs(51);
    layer0_outputs(920) <= not(inputs(132)) or (inputs(35));
    layer0_outputs(921) <= not(inputs(222)) or (inputs(240));
    layer0_outputs(922) <= (inputs(203)) xor (inputs(138));
    layer0_outputs(923) <= inputs(188);
    layer0_outputs(924) <= inputs(90);
    layer0_outputs(925) <= (inputs(61)) or (inputs(121));
    layer0_outputs(926) <= inputs(172);
    layer0_outputs(927) <= (inputs(78)) xor (inputs(191));
    layer0_outputs(928) <= (inputs(86)) and not (inputs(212));
    layer0_outputs(929) <= not((inputs(80)) or (inputs(114)));
    layer0_outputs(930) <= inputs(76);
    layer0_outputs(931) <= (inputs(147)) and not (inputs(138));
    layer0_outputs(932) <= not((inputs(206)) xor (inputs(140)));
    layer0_outputs(933) <= '0';
    layer0_outputs(934) <= not(inputs(104));
    layer0_outputs(935) <= inputs(169);
    layer0_outputs(936) <= (inputs(47)) and not (inputs(124));
    layer0_outputs(937) <= '1';
    layer0_outputs(938) <= (inputs(5)) or (inputs(36));
    layer0_outputs(939) <= (inputs(165)) or (inputs(254));
    layer0_outputs(940) <= inputs(27);
    layer0_outputs(941) <= (inputs(235)) xor (inputs(171));
    layer0_outputs(942) <= (inputs(175)) xor (inputs(20));
    layer0_outputs(943) <= (inputs(62)) xor (inputs(207));
    layer0_outputs(944) <= (inputs(177)) and (inputs(160));
    layer0_outputs(945) <= not(inputs(197)) or (inputs(222));
    layer0_outputs(946) <= not((inputs(239)) or (inputs(94)));
    layer0_outputs(947) <= not((inputs(45)) and (inputs(91)));
    layer0_outputs(948) <= not((inputs(16)) or (inputs(38)));
    layer0_outputs(949) <= (inputs(194)) and (inputs(77));
    layer0_outputs(950) <= inputs(164);
    layer0_outputs(951) <= inputs(171);
    layer0_outputs(952) <= not(inputs(243));
    layer0_outputs(953) <= not(inputs(116)) or (inputs(150));
    layer0_outputs(954) <= (inputs(222)) or (inputs(24));
    layer0_outputs(955) <= (inputs(73)) and not (inputs(0));
    layer0_outputs(956) <= not(inputs(41));
    layer0_outputs(957) <= not(inputs(110)) or (inputs(94));
    layer0_outputs(958) <= not((inputs(163)) or (inputs(79)));
    layer0_outputs(959) <= not(inputs(188));
    layer0_outputs(960) <= (inputs(232)) and not (inputs(51));
    layer0_outputs(961) <= (inputs(44)) xor (inputs(253));
    layer0_outputs(962) <= not(inputs(9));
    layer0_outputs(963) <= not((inputs(112)) or (inputs(69)));
    layer0_outputs(964) <= not((inputs(193)) or (inputs(46)));
    layer0_outputs(965) <= (inputs(147)) xor (inputs(240));
    layer0_outputs(966) <= not(inputs(231));
    layer0_outputs(967) <= (inputs(76)) or (inputs(6));
    layer0_outputs(968) <= inputs(213);
    layer0_outputs(969) <= not(inputs(202));
    layer0_outputs(970) <= (inputs(165)) or (inputs(19));
    layer0_outputs(971) <= (inputs(144)) xor (inputs(52));
    layer0_outputs(972) <= (inputs(64)) or (inputs(38));
    layer0_outputs(973) <= not((inputs(78)) and (inputs(220)));
    layer0_outputs(974) <= (inputs(45)) and (inputs(35));
    layer0_outputs(975) <= not(inputs(72)) or (inputs(157));
    layer0_outputs(976) <= (inputs(105)) and not (inputs(237));
    layer0_outputs(977) <= inputs(75);
    layer0_outputs(978) <= not(inputs(115)) or (inputs(223));
    layer0_outputs(979) <= not((inputs(160)) xor (inputs(252)));
    layer0_outputs(980) <= inputs(136);
    layer0_outputs(981) <= (inputs(218)) and not (inputs(248));
    layer0_outputs(982) <= inputs(203);
    layer0_outputs(983) <= not((inputs(164)) xor (inputs(129)));
    layer0_outputs(984) <= not((inputs(57)) and (inputs(123)));
    layer0_outputs(985) <= not((inputs(188)) or (inputs(180)));
    layer0_outputs(986) <= (inputs(51)) and not (inputs(98));
    layer0_outputs(987) <= inputs(104);
    layer0_outputs(988) <= inputs(197);
    layer0_outputs(989) <= (inputs(7)) and not (inputs(66));
    layer0_outputs(990) <= not((inputs(129)) or (inputs(215)));
    layer0_outputs(991) <= '1';
    layer0_outputs(992) <= not((inputs(84)) xor (inputs(97)));
    layer0_outputs(993) <= inputs(244);
    layer0_outputs(994) <= not((inputs(164)) xor (inputs(117)));
    layer0_outputs(995) <= inputs(40);
    layer0_outputs(996) <= (inputs(27)) and not (inputs(175));
    layer0_outputs(997) <= not(inputs(146));
    layer0_outputs(998) <= (inputs(11)) and not (inputs(190));
    layer0_outputs(999) <= inputs(150);
    layer0_outputs(1000) <= inputs(81);
    layer0_outputs(1001) <= not(inputs(245));
    layer0_outputs(1002) <= not(inputs(43)) or (inputs(65));
    layer0_outputs(1003) <= not((inputs(84)) xor (inputs(172)));
    layer0_outputs(1004) <= not((inputs(136)) or (inputs(32)));
    layer0_outputs(1005) <= not(inputs(70)) or (inputs(250));
    layer0_outputs(1006) <= (inputs(134)) or (inputs(132));
    layer0_outputs(1007) <= (inputs(226)) or (inputs(110));
    layer0_outputs(1008) <= inputs(20);
    layer0_outputs(1009) <= not((inputs(126)) or (inputs(164)));
    layer0_outputs(1010) <= inputs(84);
    layer0_outputs(1011) <= not(inputs(204));
    layer0_outputs(1012) <= (inputs(215)) xor (inputs(184));
    layer0_outputs(1013) <= not((inputs(60)) or (inputs(212)));
    layer0_outputs(1014) <= inputs(217);
    layer0_outputs(1015) <= (inputs(46)) and (inputs(88));
    layer0_outputs(1016) <= inputs(133);
    layer0_outputs(1017) <= inputs(195);
    layer0_outputs(1018) <= (inputs(188)) or (inputs(2));
    layer0_outputs(1019) <= not(inputs(44)) or (inputs(209));
    layer0_outputs(1020) <= inputs(173);
    layer0_outputs(1021) <= not((inputs(220)) or (inputs(4)));
    layer0_outputs(1022) <= inputs(216);
    layer0_outputs(1023) <= (inputs(107)) and not (inputs(167));
    layer0_outputs(1024) <= not(inputs(124)) or (inputs(247));
    layer0_outputs(1025) <= (inputs(55)) and not (inputs(66));
    layer0_outputs(1026) <= (inputs(234)) and not (inputs(163));
    layer0_outputs(1027) <= not((inputs(83)) or (inputs(46)));
    layer0_outputs(1028) <= not(inputs(24));
    layer0_outputs(1029) <= not((inputs(126)) xor (inputs(82)));
    layer0_outputs(1030) <= not(inputs(214));
    layer0_outputs(1031) <= (inputs(243)) or (inputs(36));
    layer0_outputs(1032) <= not((inputs(227)) xor (inputs(182)));
    layer0_outputs(1033) <= not(inputs(118));
    layer0_outputs(1034) <= (inputs(158)) xor (inputs(85));
    layer0_outputs(1035) <= (inputs(51)) and not (inputs(145));
    layer0_outputs(1036) <= not(inputs(169));
    layer0_outputs(1037) <= not((inputs(42)) xor (inputs(38)));
    layer0_outputs(1038) <= not(inputs(42)) or (inputs(3));
    layer0_outputs(1039) <= not(inputs(151)) or (inputs(88));
    layer0_outputs(1040) <= not((inputs(141)) xor (inputs(191)));
    layer0_outputs(1041) <= (inputs(5)) xor (inputs(221));
    layer0_outputs(1042) <= (inputs(133)) xor (inputs(151));
    layer0_outputs(1043) <= (inputs(28)) and not (inputs(80));
    layer0_outputs(1044) <= not(inputs(180)) or (inputs(124));
    layer0_outputs(1045) <= not(inputs(109));
    layer0_outputs(1046) <= not(inputs(234)) or (inputs(41));
    layer0_outputs(1047) <= not(inputs(100));
    layer0_outputs(1048) <= '0';
    layer0_outputs(1049) <= not((inputs(150)) or (inputs(177)));
    layer0_outputs(1050) <= not(inputs(74));
    layer0_outputs(1051) <= (inputs(118)) or (inputs(153));
    layer0_outputs(1052) <= not(inputs(248));
    layer0_outputs(1053) <= not(inputs(237));
    layer0_outputs(1054) <= not(inputs(65));
    layer0_outputs(1055) <= not(inputs(121)) or (inputs(213));
    layer0_outputs(1056) <= (inputs(202)) and not (inputs(78));
    layer0_outputs(1057) <= '1';
    layer0_outputs(1058) <= not((inputs(201)) xor (inputs(71)));
    layer0_outputs(1059) <= inputs(126);
    layer0_outputs(1060) <= not((inputs(172)) or (inputs(149)));
    layer0_outputs(1061) <= (inputs(10)) and not (inputs(130));
    layer0_outputs(1062) <= (inputs(92)) and not (inputs(254));
    layer0_outputs(1063) <= inputs(214);
    layer0_outputs(1064) <= (inputs(235)) xor (inputs(196));
    layer0_outputs(1065) <= not((inputs(248)) or (inputs(49)));
    layer0_outputs(1066) <= (inputs(156)) and (inputs(55));
    layer0_outputs(1067) <= inputs(102);
    layer0_outputs(1068) <= (inputs(166)) and not (inputs(2));
    layer0_outputs(1069) <= inputs(203);
    layer0_outputs(1070) <= not(inputs(163)) or (inputs(11));
    layer0_outputs(1071) <= not((inputs(5)) and (inputs(148)));
    layer0_outputs(1072) <= (inputs(94)) or (inputs(222));
    layer0_outputs(1073) <= not(inputs(129));
    layer0_outputs(1074) <= (inputs(211)) xor (inputs(44));
    layer0_outputs(1075) <= not(inputs(106)) or (inputs(70));
    layer0_outputs(1076) <= not((inputs(205)) or (inputs(80)));
    layer0_outputs(1077) <= inputs(28);
    layer0_outputs(1078) <= not(inputs(53));
    layer0_outputs(1079) <= inputs(82);
    layer0_outputs(1080) <= not((inputs(235)) xor (inputs(46)));
    layer0_outputs(1081) <= (inputs(48)) xor (inputs(237));
    layer0_outputs(1082) <= (inputs(106)) or (inputs(253));
    layer0_outputs(1083) <= not((inputs(60)) xor (inputs(4)));
    layer0_outputs(1084) <= inputs(144);
    layer0_outputs(1085) <= inputs(251);
    layer0_outputs(1086) <= not((inputs(119)) xor (inputs(211)));
    layer0_outputs(1087) <= not(inputs(83));
    layer0_outputs(1088) <= (inputs(116)) or (inputs(96));
    layer0_outputs(1089) <= inputs(234);
    layer0_outputs(1090) <= not((inputs(192)) xor (inputs(234)));
    layer0_outputs(1091) <= (inputs(204)) and not (inputs(163));
    layer0_outputs(1092) <= (inputs(213)) or (inputs(150));
    layer0_outputs(1093) <= inputs(98);
    layer0_outputs(1094) <= not(inputs(72));
    layer0_outputs(1095) <= not((inputs(29)) xor (inputs(103)));
    layer0_outputs(1096) <= (inputs(78)) or (inputs(202));
    layer0_outputs(1097) <= inputs(10);
    layer0_outputs(1098) <= (inputs(154)) and not (inputs(38));
    layer0_outputs(1099) <= not((inputs(21)) xor (inputs(78)));
    layer0_outputs(1100) <= (inputs(79)) or (inputs(207));
    layer0_outputs(1101) <= not(inputs(204)) or (inputs(241));
    layer0_outputs(1102) <= not((inputs(15)) and (inputs(29)));
    layer0_outputs(1103) <= '1';
    layer0_outputs(1104) <= '1';
    layer0_outputs(1105) <= (inputs(36)) and not (inputs(125));
    layer0_outputs(1106) <= (inputs(70)) xor (inputs(136));
    layer0_outputs(1107) <= not(inputs(24));
    layer0_outputs(1108) <= not(inputs(136)) or (inputs(14));
    layer0_outputs(1109) <= (inputs(196)) and not (inputs(157));
    layer0_outputs(1110) <= not((inputs(174)) or (inputs(157)));
    layer0_outputs(1111) <= not((inputs(188)) or (inputs(210)));
    layer0_outputs(1112) <= not((inputs(25)) and (inputs(132)));
    layer0_outputs(1113) <= (inputs(59)) and not (inputs(188));
    layer0_outputs(1114) <= (inputs(37)) and not (inputs(178));
    layer0_outputs(1115) <= (inputs(244)) and not (inputs(49));
    layer0_outputs(1116) <= (inputs(176)) and not (inputs(66));
    layer0_outputs(1117) <= not(inputs(230));
    layer0_outputs(1118) <= (inputs(5)) or (inputs(211));
    layer0_outputs(1119) <= not((inputs(233)) or (inputs(187)));
    layer0_outputs(1120) <= (inputs(178)) and not (inputs(78));
    layer0_outputs(1121) <= inputs(24);
    layer0_outputs(1122) <= not(inputs(121)) or (inputs(13));
    layer0_outputs(1123) <= (inputs(11)) xor (inputs(143));
    layer0_outputs(1124) <= not((inputs(133)) or (inputs(224)));
    layer0_outputs(1125) <= (inputs(135)) xor (inputs(103));
    layer0_outputs(1126) <= (inputs(164)) xor (inputs(194));
    layer0_outputs(1127) <= inputs(41);
    layer0_outputs(1128) <= not(inputs(252));
    layer0_outputs(1129) <= inputs(217);
    layer0_outputs(1130) <= not(inputs(215));
    layer0_outputs(1131) <= not(inputs(42));
    layer0_outputs(1132) <= (inputs(101)) xor (inputs(144));
    layer0_outputs(1133) <= not(inputs(61)) or (inputs(240));
    layer0_outputs(1134) <= not((inputs(253)) or (inputs(43)));
    layer0_outputs(1135) <= not(inputs(76));
    layer0_outputs(1136) <= not((inputs(84)) and (inputs(120)));
    layer0_outputs(1137) <= inputs(89);
    layer0_outputs(1138) <= not((inputs(158)) and (inputs(113)));
    layer0_outputs(1139) <= (inputs(140)) xor (inputs(90));
    layer0_outputs(1140) <= inputs(83);
    layer0_outputs(1141) <= (inputs(73)) xor (inputs(47));
    layer0_outputs(1142) <= inputs(62);
    layer0_outputs(1143) <= inputs(123);
    layer0_outputs(1144) <= (inputs(150)) and not (inputs(43));
    layer0_outputs(1145) <= (inputs(119)) and (inputs(107));
    layer0_outputs(1146) <= not((inputs(241)) or (inputs(192)));
    layer0_outputs(1147) <= inputs(84);
    layer0_outputs(1148) <= (inputs(35)) and not (inputs(82));
    layer0_outputs(1149) <= inputs(141);
    layer0_outputs(1150) <= '0';
    layer0_outputs(1151) <= not(inputs(180)) or (inputs(45));
    layer0_outputs(1152) <= not(inputs(162));
    layer0_outputs(1153) <= (inputs(70)) and not (inputs(57));
    layer0_outputs(1154) <= not(inputs(113));
    layer0_outputs(1155) <= (inputs(226)) or (inputs(98));
    layer0_outputs(1156) <= not(inputs(51));
    layer0_outputs(1157) <= not(inputs(245));
    layer0_outputs(1158) <= inputs(101);
    layer0_outputs(1159) <= '0';
    layer0_outputs(1160) <= not(inputs(170)) or (inputs(132));
    layer0_outputs(1161) <= (inputs(63)) or (inputs(158));
    layer0_outputs(1162) <= not(inputs(27)) or (inputs(252));
    layer0_outputs(1163) <= (inputs(241)) or (inputs(145));
    layer0_outputs(1164) <= not((inputs(218)) and (inputs(168)));
    layer0_outputs(1165) <= not((inputs(160)) xor (inputs(148)));
    layer0_outputs(1166) <= (inputs(34)) or (inputs(193));
    layer0_outputs(1167) <= (inputs(186)) and not (inputs(39));
    layer0_outputs(1168) <= (inputs(218)) or (inputs(94));
    layer0_outputs(1169) <= inputs(132);
    layer0_outputs(1170) <= (inputs(147)) xor (inputs(110));
    layer0_outputs(1171) <= (inputs(222)) xor (inputs(24));
    layer0_outputs(1172) <= (inputs(109)) xor (inputs(137));
    layer0_outputs(1173) <= not(inputs(246)) or (inputs(254));
    layer0_outputs(1174) <= not((inputs(131)) or (inputs(145)));
    layer0_outputs(1175) <= (inputs(166)) or (inputs(198));
    layer0_outputs(1176) <= not(inputs(86));
    layer0_outputs(1177) <= (inputs(50)) xor (inputs(22));
    layer0_outputs(1178) <= inputs(120);
    layer0_outputs(1179) <= not((inputs(106)) xor (inputs(137)));
    layer0_outputs(1180) <= not(inputs(131));
    layer0_outputs(1181) <= inputs(151);
    layer0_outputs(1182) <= (inputs(38)) and not (inputs(2));
    layer0_outputs(1183) <= (inputs(96)) xor (inputs(227));
    layer0_outputs(1184) <= (inputs(214)) or (inputs(229));
    layer0_outputs(1185) <= not(inputs(78));
    layer0_outputs(1186) <= (inputs(2)) or (inputs(175));
    layer0_outputs(1187) <= not(inputs(82)) or (inputs(191));
    layer0_outputs(1188) <= inputs(227);
    layer0_outputs(1189) <= (inputs(180)) or (inputs(18));
    layer0_outputs(1190) <= inputs(189);
    layer0_outputs(1191) <= inputs(58);
    layer0_outputs(1192) <= inputs(178);
    layer0_outputs(1193) <= not(inputs(26)) or (inputs(241));
    layer0_outputs(1194) <= not(inputs(89)) or (inputs(143));
    layer0_outputs(1195) <= (inputs(142)) and (inputs(145));
    layer0_outputs(1196) <= not((inputs(47)) xor (inputs(6)));
    layer0_outputs(1197) <= not(inputs(90));
    layer0_outputs(1198) <= (inputs(148)) and not (inputs(0));
    layer0_outputs(1199) <= (inputs(80)) and not (inputs(13));
    layer0_outputs(1200) <= not(inputs(45));
    layer0_outputs(1201) <= not(inputs(113));
    layer0_outputs(1202) <= not(inputs(230)) or (inputs(106));
    layer0_outputs(1203) <= inputs(19);
    layer0_outputs(1204) <= not(inputs(162));
    layer0_outputs(1205) <= not((inputs(232)) or (inputs(211)));
    layer0_outputs(1206) <= (inputs(87)) and not (inputs(88));
    layer0_outputs(1207) <= (inputs(166)) and not (inputs(208));
    layer0_outputs(1208) <= not(inputs(196)) or (inputs(132));
    layer0_outputs(1209) <= not((inputs(156)) or (inputs(118)));
    layer0_outputs(1210) <= inputs(150);
    layer0_outputs(1211) <= not((inputs(113)) or (inputs(208)));
    layer0_outputs(1212) <= not(inputs(91)) or (inputs(196));
    layer0_outputs(1213) <= not((inputs(89)) xor (inputs(37)));
    layer0_outputs(1214) <= (inputs(66)) and not (inputs(2));
    layer0_outputs(1215) <= (inputs(105)) xor (inputs(126));
    layer0_outputs(1216) <= not((inputs(130)) and (inputs(167)));
    layer0_outputs(1217) <= inputs(152);
    layer0_outputs(1218) <= inputs(121);
    layer0_outputs(1219) <= not(inputs(101));
    layer0_outputs(1220) <= inputs(230);
    layer0_outputs(1221) <= not((inputs(170)) xor (inputs(217)));
    layer0_outputs(1222) <= not(inputs(218)) or (inputs(202));
    layer0_outputs(1223) <= not(inputs(101));
    layer0_outputs(1224) <= not((inputs(40)) or (inputs(243)));
    layer0_outputs(1225) <= (inputs(5)) or (inputs(145));
    layer0_outputs(1226) <= inputs(231);
    layer0_outputs(1227) <= not(inputs(194));
    layer0_outputs(1228) <= (inputs(76)) and (inputs(146));
    layer0_outputs(1229) <= not((inputs(15)) or (inputs(83)));
    layer0_outputs(1230) <= inputs(4);
    layer0_outputs(1231) <= not((inputs(205)) and (inputs(185)));
    layer0_outputs(1232) <= (inputs(250)) or (inputs(217));
    layer0_outputs(1233) <= inputs(194);
    layer0_outputs(1234) <= '1';
    layer0_outputs(1235) <= not(inputs(115)) or (inputs(209));
    layer0_outputs(1236) <= (inputs(184)) or (inputs(161));
    layer0_outputs(1237) <= not(inputs(117)) or (inputs(75));
    layer0_outputs(1238) <= not(inputs(131));
    layer0_outputs(1239) <= inputs(62);
    layer0_outputs(1240) <= inputs(149);
    layer0_outputs(1241) <= inputs(112);
    layer0_outputs(1242) <= not(inputs(168));
    layer0_outputs(1243) <= (inputs(245)) or (inputs(160));
    layer0_outputs(1244) <= (inputs(211)) and not (inputs(90));
    layer0_outputs(1245) <= (inputs(183)) and not (inputs(27));
    layer0_outputs(1246) <= not((inputs(202)) or (inputs(127)));
    layer0_outputs(1247) <= (inputs(110)) or (inputs(213));
    layer0_outputs(1248) <= inputs(48);
    layer0_outputs(1249) <= inputs(228);
    layer0_outputs(1250) <= not((inputs(0)) and (inputs(67)));
    layer0_outputs(1251) <= (inputs(206)) xor (inputs(224));
    layer0_outputs(1252) <= (inputs(83)) and not (inputs(43));
    layer0_outputs(1253) <= not(inputs(121));
    layer0_outputs(1254) <= (inputs(161)) or (inputs(160));
    layer0_outputs(1255) <= not((inputs(79)) and (inputs(170)));
    layer0_outputs(1256) <= (inputs(26)) or (inputs(238));
    layer0_outputs(1257) <= (inputs(2)) or (inputs(178));
    layer0_outputs(1258) <= (inputs(19)) or (inputs(211));
    layer0_outputs(1259) <= not(inputs(182));
    layer0_outputs(1260) <= (inputs(250)) and (inputs(37));
    layer0_outputs(1261) <= (inputs(80)) or (inputs(208));
    layer0_outputs(1262) <= not((inputs(41)) xor (inputs(29)));
    layer0_outputs(1263) <= not(inputs(220));
    layer0_outputs(1264) <= not(inputs(3));
    layer0_outputs(1265) <= (inputs(1)) xor (inputs(193));
    layer0_outputs(1266) <= inputs(157);
    layer0_outputs(1267) <= (inputs(118)) and not (inputs(222));
    layer0_outputs(1268) <= (inputs(22)) and (inputs(230));
    layer0_outputs(1269) <= not((inputs(128)) or (inputs(85)));
    layer0_outputs(1270) <= inputs(227);
    layer0_outputs(1271) <= not((inputs(91)) xor (inputs(116)));
    layer0_outputs(1272) <= not(inputs(234)) or (inputs(239));
    layer0_outputs(1273) <= (inputs(226)) or (inputs(159));
    layer0_outputs(1274) <= inputs(121);
    layer0_outputs(1275) <= (inputs(90)) and not (inputs(198));
    layer0_outputs(1276) <= inputs(223);
    layer0_outputs(1277) <= not(inputs(252)) or (inputs(103));
    layer0_outputs(1278) <= not(inputs(119));
    layer0_outputs(1279) <= not(inputs(9));
    layer0_outputs(1280) <= (inputs(196)) and not (inputs(182));
    layer0_outputs(1281) <= (inputs(26)) and not (inputs(199));
    layer0_outputs(1282) <= (inputs(207)) xor (inputs(70));
    layer0_outputs(1283) <= not((inputs(218)) xor (inputs(145)));
    layer0_outputs(1284) <= (inputs(78)) or (inputs(2));
    layer0_outputs(1285) <= inputs(115);
    layer0_outputs(1286) <= (inputs(185)) or (inputs(130));
    layer0_outputs(1287) <= not(inputs(26));
    layer0_outputs(1288) <= inputs(248);
    layer0_outputs(1289) <= not((inputs(123)) or (inputs(5)));
    layer0_outputs(1290) <= (inputs(49)) and not (inputs(37));
    layer0_outputs(1291) <= inputs(83);
    layer0_outputs(1292) <= not(inputs(24)) or (inputs(147));
    layer0_outputs(1293) <= inputs(153);
    layer0_outputs(1294) <= (inputs(182)) or (inputs(172));
    layer0_outputs(1295) <= '1';
    layer0_outputs(1296) <= not(inputs(45));
    layer0_outputs(1297) <= not((inputs(227)) xor (inputs(233)));
    layer0_outputs(1298) <= (inputs(55)) and not (inputs(207));
    layer0_outputs(1299) <= (inputs(38)) xor (inputs(244));
    layer0_outputs(1300) <= (inputs(217)) and not (inputs(18));
    layer0_outputs(1301) <= inputs(112);
    layer0_outputs(1302) <= (inputs(118)) xor (inputs(146));
    layer0_outputs(1303) <= not((inputs(46)) or (inputs(69)));
    layer0_outputs(1304) <= inputs(2);
    layer0_outputs(1305) <= not(inputs(212));
    layer0_outputs(1306) <= (inputs(209)) or (inputs(182));
    layer0_outputs(1307) <= not((inputs(175)) xor (inputs(247)));
    layer0_outputs(1308) <= inputs(121);
    layer0_outputs(1309) <= (inputs(124)) and not (inputs(216));
    layer0_outputs(1310) <= not((inputs(68)) or (inputs(179)));
    layer0_outputs(1311) <= not(inputs(228)) or (inputs(225));
    layer0_outputs(1312) <= not(inputs(121)) or (inputs(41));
    layer0_outputs(1313) <= not((inputs(127)) or (inputs(181)));
    layer0_outputs(1314) <= not(inputs(59));
    layer0_outputs(1315) <= (inputs(222)) and not (inputs(136));
    layer0_outputs(1316) <= (inputs(171)) xor (inputs(109));
    layer0_outputs(1317) <= (inputs(140)) and not (inputs(201));
    layer0_outputs(1318) <= not((inputs(143)) xor (inputs(11)));
    layer0_outputs(1319) <= (inputs(206)) or (inputs(15));
    layer0_outputs(1320) <= (inputs(207)) and not (inputs(161));
    layer0_outputs(1321) <= not((inputs(156)) xor (inputs(6)));
    layer0_outputs(1322) <= not((inputs(55)) or (inputs(96)));
    layer0_outputs(1323) <= (inputs(229)) or (inputs(189));
    layer0_outputs(1324) <= not(inputs(250)) or (inputs(142));
    layer0_outputs(1325) <= inputs(42);
    layer0_outputs(1326) <= not((inputs(158)) xor (inputs(207)));
    layer0_outputs(1327) <= not((inputs(135)) xor (inputs(164)));
    layer0_outputs(1328) <= inputs(228);
    layer0_outputs(1329) <= not((inputs(117)) or (inputs(78)));
    layer0_outputs(1330) <= not((inputs(148)) or (inputs(94)));
    layer0_outputs(1331) <= inputs(129);
    layer0_outputs(1332) <= not((inputs(94)) or (inputs(196)));
    layer0_outputs(1333) <= (inputs(186)) or (inputs(27));
    layer0_outputs(1334) <= inputs(245);
    layer0_outputs(1335) <= not(inputs(40));
    layer0_outputs(1336) <= (inputs(238)) and (inputs(235));
    layer0_outputs(1337) <= not((inputs(43)) or (inputs(207)));
    layer0_outputs(1338) <= not((inputs(254)) xor (inputs(176)));
    layer0_outputs(1339) <= inputs(39);
    layer0_outputs(1340) <= (inputs(80)) or (inputs(108));
    layer0_outputs(1341) <= (inputs(233)) or (inputs(212));
    layer0_outputs(1342) <= (inputs(132)) xor (inputs(128));
    layer0_outputs(1343) <= not(inputs(21)) or (inputs(82));
    layer0_outputs(1344) <= inputs(184);
    layer0_outputs(1345) <= inputs(91);
    layer0_outputs(1346) <= not(inputs(168));
    layer0_outputs(1347) <= inputs(5);
    layer0_outputs(1348) <= (inputs(209)) xor (inputs(177));
    layer0_outputs(1349) <= not(inputs(85)) or (inputs(176));
    layer0_outputs(1350) <= not(inputs(76));
    layer0_outputs(1351) <= (inputs(248)) and not (inputs(245));
    layer0_outputs(1352) <= not(inputs(214));
    layer0_outputs(1353) <= (inputs(73)) xor (inputs(155));
    layer0_outputs(1354) <= not(inputs(12)) or (inputs(168));
    layer0_outputs(1355) <= not(inputs(115));
    layer0_outputs(1356) <= not(inputs(101)) or (inputs(18));
    layer0_outputs(1357) <= not((inputs(217)) or (inputs(238)));
    layer0_outputs(1358) <= not((inputs(35)) or (inputs(160)));
    layer0_outputs(1359) <= not((inputs(255)) or (inputs(219)));
    layer0_outputs(1360) <= not((inputs(48)) or (inputs(188)));
    layer0_outputs(1361) <= inputs(5);
    layer0_outputs(1362) <= not((inputs(199)) xor (inputs(161)));
    layer0_outputs(1363) <= (inputs(74)) or (inputs(61));
    layer0_outputs(1364) <= (inputs(172)) xor (inputs(161));
    layer0_outputs(1365) <= '1';
    layer0_outputs(1366) <= (inputs(251)) xor (inputs(190));
    layer0_outputs(1367) <= (inputs(180)) xor (inputs(155));
    layer0_outputs(1368) <= inputs(220);
    layer0_outputs(1369) <= (inputs(48)) or (inputs(213));
    layer0_outputs(1370) <= not(inputs(67));
    layer0_outputs(1371) <= '1';
    layer0_outputs(1372) <= not((inputs(52)) and (inputs(38)));
    layer0_outputs(1373) <= not(inputs(132)) or (inputs(12));
    layer0_outputs(1374) <= not(inputs(59));
    layer0_outputs(1375) <= not((inputs(23)) or (inputs(225)));
    layer0_outputs(1376) <= (inputs(27)) and not (inputs(206));
    layer0_outputs(1377) <= (inputs(243)) or (inputs(156));
    layer0_outputs(1378) <= not(inputs(69));
    layer0_outputs(1379) <= (inputs(244)) and (inputs(28));
    layer0_outputs(1380) <= not(inputs(37)) or (inputs(191));
    layer0_outputs(1381) <= not((inputs(86)) or (inputs(127)));
    layer0_outputs(1382) <= (inputs(100)) and (inputs(44));
    layer0_outputs(1383) <= (inputs(107)) xor (inputs(1));
    layer0_outputs(1384) <= inputs(111);
    layer0_outputs(1385) <= not(inputs(51));
    layer0_outputs(1386) <= not(inputs(107)) or (inputs(40));
    layer0_outputs(1387) <= (inputs(122)) and not (inputs(73));
    layer0_outputs(1388) <= not((inputs(238)) and (inputs(5)));
    layer0_outputs(1389) <= not(inputs(53)) or (inputs(155));
    layer0_outputs(1390) <= (inputs(116)) and not (inputs(242));
    layer0_outputs(1391) <= (inputs(29)) or (inputs(93));
    layer0_outputs(1392) <= (inputs(42)) xor (inputs(38));
    layer0_outputs(1393) <= '1';
    layer0_outputs(1394) <= inputs(25);
    layer0_outputs(1395) <= (inputs(111)) xor (inputs(65));
    layer0_outputs(1396) <= not(inputs(54));
    layer0_outputs(1397) <= (inputs(196)) and not (inputs(249));
    layer0_outputs(1398) <= not(inputs(144));
    layer0_outputs(1399) <= (inputs(202)) or (inputs(238));
    layer0_outputs(1400) <= not(inputs(176)) or (inputs(139));
    layer0_outputs(1401) <= (inputs(38)) and not (inputs(173));
    layer0_outputs(1402) <= '0';
    layer0_outputs(1403) <= not((inputs(81)) xor (inputs(85)));
    layer0_outputs(1404) <= not(inputs(188)) or (inputs(12));
    layer0_outputs(1405) <= (inputs(147)) and not (inputs(36));
    layer0_outputs(1406) <= inputs(91);
    layer0_outputs(1407) <= inputs(165);
    layer0_outputs(1408) <= inputs(138);
    layer0_outputs(1409) <= (inputs(0)) xor (inputs(229));
    layer0_outputs(1410) <= not((inputs(30)) or (inputs(48)));
    layer0_outputs(1411) <= not(inputs(133)) or (inputs(21));
    layer0_outputs(1412) <= not(inputs(75)) or (inputs(20));
    layer0_outputs(1413) <= not(inputs(130));
    layer0_outputs(1414) <= (inputs(26)) or (inputs(40));
    layer0_outputs(1415) <= (inputs(91)) or (inputs(146));
    layer0_outputs(1416) <= (inputs(187)) xor (inputs(21));
    layer0_outputs(1417) <= not((inputs(90)) or (inputs(2)));
    layer0_outputs(1418) <= inputs(202);
    layer0_outputs(1419) <= inputs(190);
    layer0_outputs(1420) <= inputs(147);
    layer0_outputs(1421) <= not((inputs(250)) xor (inputs(54)));
    layer0_outputs(1422) <= (inputs(118)) xor (inputs(188));
    layer0_outputs(1423) <= (inputs(122)) and not (inputs(1));
    layer0_outputs(1424) <= inputs(118);
    layer0_outputs(1425) <= not(inputs(206));
    layer0_outputs(1426) <= not(inputs(73));
    layer0_outputs(1427) <= not((inputs(89)) or (inputs(223)));
    layer0_outputs(1428) <= (inputs(74)) and not (inputs(208));
    layer0_outputs(1429) <= inputs(9);
    layer0_outputs(1430) <= not(inputs(102));
    layer0_outputs(1431) <= (inputs(92)) or (inputs(47));
    layer0_outputs(1432) <= (inputs(104)) xor (inputs(53));
    layer0_outputs(1433) <= inputs(56);
    layer0_outputs(1434) <= (inputs(118)) and not (inputs(116));
    layer0_outputs(1435) <= inputs(169);
    layer0_outputs(1436) <= (inputs(149)) and (inputs(196));
    layer0_outputs(1437) <= inputs(68);
    layer0_outputs(1438) <= (inputs(59)) or (inputs(111));
    layer0_outputs(1439) <= (inputs(163)) or (inputs(236));
    layer0_outputs(1440) <= not(inputs(226)) or (inputs(159));
    layer0_outputs(1441) <= not((inputs(17)) xor (inputs(73)));
    layer0_outputs(1442) <= (inputs(94)) xor (inputs(142));
    layer0_outputs(1443) <= not((inputs(60)) xor (inputs(30)));
    layer0_outputs(1444) <= not(inputs(85)) or (inputs(252));
    layer0_outputs(1445) <= not((inputs(218)) and (inputs(22)));
    layer0_outputs(1446) <= not((inputs(229)) or (inputs(230)));
    layer0_outputs(1447) <= (inputs(107)) or (inputs(16));
    layer0_outputs(1448) <= not(inputs(90));
    layer0_outputs(1449) <= not((inputs(184)) or (inputs(91)));
    layer0_outputs(1450) <= (inputs(61)) or (inputs(73));
    layer0_outputs(1451) <= not(inputs(9));
    layer0_outputs(1452) <= not(inputs(219)) or (inputs(30));
    layer0_outputs(1453) <= (inputs(213)) and not (inputs(26));
    layer0_outputs(1454) <= not((inputs(177)) or (inputs(86)));
    layer0_outputs(1455) <= not((inputs(44)) xor (inputs(210)));
    layer0_outputs(1456) <= (inputs(31)) and not (inputs(35));
    layer0_outputs(1457) <= not((inputs(85)) xor (inputs(65)));
    layer0_outputs(1458) <= inputs(87);
    layer0_outputs(1459) <= (inputs(2)) xor (inputs(174));
    layer0_outputs(1460) <= not(inputs(31));
    layer0_outputs(1461) <= not((inputs(154)) or (inputs(20)));
    layer0_outputs(1462) <= (inputs(249)) xor (inputs(159));
    layer0_outputs(1463) <= (inputs(166)) and not (inputs(98));
    layer0_outputs(1464) <= '0';
    layer0_outputs(1465) <= (inputs(169)) and not (inputs(63));
    layer0_outputs(1466) <= not((inputs(135)) or (inputs(252)));
    layer0_outputs(1467) <= not(inputs(177));
    layer0_outputs(1468) <= (inputs(77)) and not (inputs(255));
    layer0_outputs(1469) <= (inputs(153)) and not (inputs(188));
    layer0_outputs(1470) <= not((inputs(112)) xor (inputs(232)));
    layer0_outputs(1471) <= (inputs(211)) or (inputs(233));
    layer0_outputs(1472) <= (inputs(167)) and not (inputs(87));
    layer0_outputs(1473) <= not((inputs(76)) xor (inputs(20)));
    layer0_outputs(1474) <= not(inputs(22));
    layer0_outputs(1475) <= not(inputs(137)) or (inputs(239));
    layer0_outputs(1476) <= not(inputs(127));
    layer0_outputs(1477) <= not(inputs(75));
    layer0_outputs(1478) <= inputs(199);
    layer0_outputs(1479) <= (inputs(201)) and not (inputs(214));
    layer0_outputs(1480) <= inputs(120);
    layer0_outputs(1481) <= inputs(52);
    layer0_outputs(1482) <= (inputs(133)) and (inputs(139));
    layer0_outputs(1483) <= not(inputs(137));
    layer0_outputs(1484) <= inputs(204);
    layer0_outputs(1485) <= not(inputs(228));
    layer0_outputs(1486) <= not(inputs(99));
    layer0_outputs(1487) <= not(inputs(67)) or (inputs(114));
    layer0_outputs(1488) <= inputs(3);
    layer0_outputs(1489) <= (inputs(41)) or (inputs(0));
    layer0_outputs(1490) <= inputs(247);
    layer0_outputs(1491) <= (inputs(121)) xor (inputs(150));
    layer0_outputs(1492) <= not((inputs(219)) or (inputs(11)));
    layer0_outputs(1493) <= (inputs(157)) xor (inputs(140));
    layer0_outputs(1494) <= (inputs(1)) or (inputs(179));
    layer0_outputs(1495) <= inputs(74);
    layer0_outputs(1496) <= inputs(72);
    layer0_outputs(1497) <= not((inputs(8)) or (inputs(29)));
    layer0_outputs(1498) <= not((inputs(131)) or (inputs(216)));
    layer0_outputs(1499) <= (inputs(228)) xor (inputs(119));
    layer0_outputs(1500) <= (inputs(179)) and not (inputs(63));
    layer0_outputs(1501) <= not(inputs(107));
    layer0_outputs(1502) <= not((inputs(21)) xor (inputs(54)));
    layer0_outputs(1503) <= (inputs(118)) and not (inputs(5));
    layer0_outputs(1504) <= not(inputs(98)) or (inputs(193));
    layer0_outputs(1505) <= not((inputs(178)) xor (inputs(192)));
    layer0_outputs(1506) <= (inputs(100)) xor (inputs(222));
    layer0_outputs(1507) <= (inputs(76)) or (inputs(141));
    layer0_outputs(1508) <= (inputs(228)) or (inputs(82));
    layer0_outputs(1509) <= inputs(42);
    layer0_outputs(1510) <= not(inputs(130)) or (inputs(49));
    layer0_outputs(1511) <= not((inputs(203)) or (inputs(143)));
    layer0_outputs(1512) <= not(inputs(212));
    layer0_outputs(1513) <= inputs(150);
    layer0_outputs(1514) <= (inputs(244)) and not (inputs(21));
    layer0_outputs(1515) <= not(inputs(97)) or (inputs(30));
    layer0_outputs(1516) <= (inputs(191)) or (inputs(65));
    layer0_outputs(1517) <= not(inputs(122));
    layer0_outputs(1518) <= inputs(152);
    layer0_outputs(1519) <= not((inputs(221)) xor (inputs(219)));
    layer0_outputs(1520) <= not(inputs(90));
    layer0_outputs(1521) <= (inputs(92)) and not (inputs(162));
    layer0_outputs(1522) <= not(inputs(113));
    layer0_outputs(1523) <= (inputs(248)) xor (inputs(239));
    layer0_outputs(1524) <= (inputs(87)) and not (inputs(34));
    layer0_outputs(1525) <= inputs(214);
    layer0_outputs(1526) <= (inputs(218)) or (inputs(141));
    layer0_outputs(1527) <= not((inputs(188)) or (inputs(82)));
    layer0_outputs(1528) <= inputs(57);
    layer0_outputs(1529) <= (inputs(25)) and not (inputs(147));
    layer0_outputs(1530) <= (inputs(219)) or (inputs(81));
    layer0_outputs(1531) <= not((inputs(155)) or (inputs(217)));
    layer0_outputs(1532) <= inputs(55);
    layer0_outputs(1533) <= not(inputs(231));
    layer0_outputs(1534) <= not(inputs(151));
    layer0_outputs(1535) <= (inputs(215)) and not (inputs(106));
    layer0_outputs(1536) <= (inputs(33)) or (inputs(224));
    layer0_outputs(1537) <= not((inputs(249)) xor (inputs(16)));
    layer0_outputs(1538) <= not(inputs(145));
    layer0_outputs(1539) <= inputs(19);
    layer0_outputs(1540) <= '1';
    layer0_outputs(1541) <= not((inputs(105)) or (inputs(6)));
    layer0_outputs(1542) <= not(inputs(233)) or (inputs(107));
    layer0_outputs(1543) <= (inputs(82)) or (inputs(65));
    layer0_outputs(1544) <= inputs(163);
    layer0_outputs(1545) <= not(inputs(242));
    layer0_outputs(1546) <= (inputs(196)) and not (inputs(255));
    layer0_outputs(1547) <= inputs(189);
    layer0_outputs(1548) <= not(inputs(74)) or (inputs(96));
    layer0_outputs(1549) <= not(inputs(20));
    layer0_outputs(1550) <= not(inputs(196)) or (inputs(40));
    layer0_outputs(1551) <= not((inputs(62)) or (inputs(155)));
    layer0_outputs(1552) <= (inputs(129)) or (inputs(130));
    layer0_outputs(1553) <= inputs(41);
    layer0_outputs(1554) <= not(inputs(170)) or (inputs(46));
    layer0_outputs(1555) <= not(inputs(73));
    layer0_outputs(1556) <= (inputs(26)) and not (inputs(172));
    layer0_outputs(1557) <= not(inputs(250));
    layer0_outputs(1558) <= inputs(51);
    layer0_outputs(1559) <= (inputs(192)) and not (inputs(242));
    layer0_outputs(1560) <= not(inputs(59));
    layer0_outputs(1561) <= (inputs(249)) and not (inputs(64));
    layer0_outputs(1562) <= not(inputs(6)) or (inputs(190));
    layer0_outputs(1563) <= not((inputs(24)) or (inputs(192)));
    layer0_outputs(1564) <= not(inputs(152)) or (inputs(144));
    layer0_outputs(1565) <= (inputs(60)) or (inputs(151));
    layer0_outputs(1566) <= not(inputs(211));
    layer0_outputs(1567) <= not(inputs(80));
    layer0_outputs(1568) <= not((inputs(106)) xor (inputs(254)));
    layer0_outputs(1569) <= not(inputs(247)) or (inputs(42));
    layer0_outputs(1570) <= inputs(231);
    layer0_outputs(1571) <= inputs(18);
    layer0_outputs(1572) <= not(inputs(105));
    layer0_outputs(1573) <= not((inputs(15)) or (inputs(134)));
    layer0_outputs(1574) <= (inputs(74)) and not (inputs(243));
    layer0_outputs(1575) <= not(inputs(218)) or (inputs(184));
    layer0_outputs(1576) <= '1';
    layer0_outputs(1577) <= inputs(55);
    layer0_outputs(1578) <= (inputs(118)) and not (inputs(111));
    layer0_outputs(1579) <= (inputs(187)) and not (inputs(99));
    layer0_outputs(1580) <= (inputs(209)) or (inputs(184));
    layer0_outputs(1581) <= not(inputs(181));
    layer0_outputs(1582) <= inputs(147);
    layer0_outputs(1583) <= not((inputs(103)) xor (inputs(182)));
    layer0_outputs(1584) <= not(inputs(189)) or (inputs(46));
    layer0_outputs(1585) <= not((inputs(191)) or (inputs(195)));
    layer0_outputs(1586) <= not(inputs(45)) or (inputs(34));
    layer0_outputs(1587) <= not((inputs(97)) or (inputs(29)));
    layer0_outputs(1588) <= inputs(183);
    layer0_outputs(1589) <= not(inputs(9));
    layer0_outputs(1590) <= not(inputs(41));
    layer0_outputs(1591) <= not((inputs(210)) or (inputs(143)));
    layer0_outputs(1592) <= (inputs(144)) or (inputs(253));
    layer0_outputs(1593) <= not(inputs(207)) or (inputs(162));
    layer0_outputs(1594) <= (inputs(25)) and not (inputs(237));
    layer0_outputs(1595) <= (inputs(35)) or (inputs(42));
    layer0_outputs(1596) <= (inputs(200)) and (inputs(157));
    layer0_outputs(1597) <= not(inputs(229));
    layer0_outputs(1598) <= '1';
    layer0_outputs(1599) <= (inputs(220)) or (inputs(200));
    layer0_outputs(1600) <= not(inputs(11)) or (inputs(218));
    layer0_outputs(1601) <= (inputs(55)) or (inputs(112));
    layer0_outputs(1602) <= inputs(136);
    layer0_outputs(1603) <= inputs(213);
    layer0_outputs(1604) <= not((inputs(188)) or (inputs(245)));
    layer0_outputs(1605) <= '1';
    layer0_outputs(1606) <= not((inputs(75)) or (inputs(177)));
    layer0_outputs(1607) <= (inputs(172)) or (inputs(216));
    layer0_outputs(1608) <= (inputs(134)) and not (inputs(40));
    layer0_outputs(1609) <= (inputs(137)) and not (inputs(224));
    layer0_outputs(1610) <= inputs(22);
    layer0_outputs(1611) <= not(inputs(215));
    layer0_outputs(1612) <= (inputs(119)) and not (inputs(101));
    layer0_outputs(1613) <= not((inputs(22)) and (inputs(23)));
    layer0_outputs(1614) <= not((inputs(158)) or (inputs(115)));
    layer0_outputs(1615) <= not((inputs(218)) xor (inputs(155)));
    layer0_outputs(1616) <= not(inputs(208)) or (inputs(156));
    layer0_outputs(1617) <= not(inputs(21)) or (inputs(115));
    layer0_outputs(1618) <= not(inputs(245)) or (inputs(55));
    layer0_outputs(1619) <= (inputs(73)) or (inputs(45));
    layer0_outputs(1620) <= (inputs(32)) or (inputs(22));
    layer0_outputs(1621) <= '1';
    layer0_outputs(1622) <= inputs(59);
    layer0_outputs(1623) <= not((inputs(242)) xor (inputs(34)));
    layer0_outputs(1624) <= not(inputs(91)) or (inputs(162));
    layer0_outputs(1625) <= not((inputs(234)) or (inputs(15)));
    layer0_outputs(1626) <= not((inputs(197)) or (inputs(146)));
    layer0_outputs(1627) <= (inputs(54)) and not (inputs(225));
    layer0_outputs(1628) <= not((inputs(242)) or (inputs(95)));
    layer0_outputs(1629) <= not(inputs(48)) or (inputs(80));
    layer0_outputs(1630) <= (inputs(136)) xor (inputs(255));
    layer0_outputs(1631) <= not(inputs(103));
    layer0_outputs(1632) <= (inputs(237)) and (inputs(182));
    layer0_outputs(1633) <= not(inputs(134)) or (inputs(177));
    layer0_outputs(1634) <= inputs(25);
    layer0_outputs(1635) <= (inputs(40)) or (inputs(253));
    layer0_outputs(1636) <= (inputs(121)) xor (inputs(150));
    layer0_outputs(1637) <= not(inputs(93));
    layer0_outputs(1638) <= inputs(140);
    layer0_outputs(1639) <= (inputs(12)) xor (inputs(168));
    layer0_outputs(1640) <= not((inputs(13)) xor (inputs(51)));
    layer0_outputs(1641) <= inputs(23);
    layer0_outputs(1642) <= (inputs(229)) and not (inputs(79));
    layer0_outputs(1643) <= not((inputs(65)) or (inputs(83)));
    layer0_outputs(1644) <= not((inputs(179)) or (inputs(80)));
    layer0_outputs(1645) <= (inputs(187)) xor (inputs(62));
    layer0_outputs(1646) <= inputs(195);
    layer0_outputs(1647) <= not(inputs(96));
    layer0_outputs(1648) <= not(inputs(85));
    layer0_outputs(1649) <= (inputs(163)) or (inputs(168));
    layer0_outputs(1650) <= (inputs(52)) and not (inputs(17));
    layer0_outputs(1651) <= not(inputs(165));
    layer0_outputs(1652) <= not(inputs(113));
    layer0_outputs(1653) <= not(inputs(127));
    layer0_outputs(1654) <= (inputs(84)) xor (inputs(54));
    layer0_outputs(1655) <= not((inputs(161)) or (inputs(18)));
    layer0_outputs(1656) <= not((inputs(206)) or (inputs(242)));
    layer0_outputs(1657) <= (inputs(13)) or (inputs(237));
    layer0_outputs(1658) <= (inputs(173)) xor (inputs(209));
    layer0_outputs(1659) <= inputs(99);
    layer0_outputs(1660) <= not(inputs(43));
    layer0_outputs(1661) <= not((inputs(8)) xor (inputs(33)));
    layer0_outputs(1662) <= not((inputs(174)) or (inputs(125)));
    layer0_outputs(1663) <= (inputs(44)) xor (inputs(245));
    layer0_outputs(1664) <= not((inputs(131)) or (inputs(102)));
    layer0_outputs(1665) <= (inputs(177)) or (inputs(166));
    layer0_outputs(1666) <= inputs(116);
    layer0_outputs(1667) <= not(inputs(236)) or (inputs(112));
    layer0_outputs(1668) <= (inputs(79)) or (inputs(1));
    layer0_outputs(1669) <= not((inputs(53)) xor (inputs(121)));
    layer0_outputs(1670) <= (inputs(29)) xor (inputs(75));
    layer0_outputs(1671) <= not(inputs(201));
    layer0_outputs(1672) <= inputs(156);
    layer0_outputs(1673) <= not((inputs(244)) xor (inputs(32)));
    layer0_outputs(1674) <= not((inputs(37)) or (inputs(63)));
    layer0_outputs(1675) <= (inputs(1)) xor (inputs(6));
    layer0_outputs(1676) <= not((inputs(10)) and (inputs(178)));
    layer0_outputs(1677) <= not((inputs(183)) or (inputs(19)));
    layer0_outputs(1678) <= not((inputs(11)) or (inputs(83)));
    layer0_outputs(1679) <= not(inputs(131));
    layer0_outputs(1680) <= (inputs(101)) or (inputs(178));
    layer0_outputs(1681) <= inputs(136);
    layer0_outputs(1682) <= (inputs(160)) xor (inputs(5));
    layer0_outputs(1683) <= inputs(56);
    layer0_outputs(1684) <= not(inputs(67));
    layer0_outputs(1685) <= not((inputs(99)) or (inputs(98)));
    layer0_outputs(1686) <= not((inputs(145)) or (inputs(214)));
    layer0_outputs(1687) <= not(inputs(113));
    layer0_outputs(1688) <= not(inputs(248));
    layer0_outputs(1689) <= (inputs(173)) or (inputs(34));
    layer0_outputs(1690) <= (inputs(157)) or (inputs(130));
    layer0_outputs(1691) <= not(inputs(4));
    layer0_outputs(1692) <= (inputs(84)) or (inputs(48));
    layer0_outputs(1693) <= not(inputs(237));
    layer0_outputs(1694) <= (inputs(38)) xor (inputs(208));
    layer0_outputs(1695) <= not(inputs(165));
    layer0_outputs(1696) <= inputs(180);
    layer0_outputs(1697) <= not((inputs(171)) xor (inputs(121)));
    layer0_outputs(1698) <= not((inputs(236)) or (inputs(133)));
    layer0_outputs(1699) <= not(inputs(43));
    layer0_outputs(1700) <= not((inputs(16)) and (inputs(182)));
    layer0_outputs(1701) <= not(inputs(229));
    layer0_outputs(1702) <= (inputs(71)) and not (inputs(139));
    layer0_outputs(1703) <= not(inputs(234)) or (inputs(26));
    layer0_outputs(1704) <= inputs(136);
    layer0_outputs(1705) <= not(inputs(223));
    layer0_outputs(1706) <= (inputs(221)) xor (inputs(27));
    layer0_outputs(1707) <= not((inputs(231)) xor (inputs(155)));
    layer0_outputs(1708) <= (inputs(209)) or (inputs(245));
    layer0_outputs(1709) <= (inputs(17)) xor (inputs(137));
    layer0_outputs(1710) <= not(inputs(89)) or (inputs(191));
    layer0_outputs(1711) <= not(inputs(165));
    layer0_outputs(1712) <= not(inputs(217));
    layer0_outputs(1713) <= inputs(230);
    layer0_outputs(1714) <= (inputs(90)) or (inputs(59));
    layer0_outputs(1715) <= (inputs(209)) and (inputs(224));
    layer0_outputs(1716) <= (inputs(221)) and not (inputs(206));
    layer0_outputs(1717) <= inputs(43);
    layer0_outputs(1718) <= not(inputs(183));
    layer0_outputs(1719) <= (inputs(120)) xor (inputs(49));
    layer0_outputs(1720) <= not((inputs(237)) or (inputs(232)));
    layer0_outputs(1721) <= not((inputs(111)) or (inputs(19)));
    layer0_outputs(1722) <= not(inputs(21));
    layer0_outputs(1723) <= (inputs(244)) and (inputs(216));
    layer0_outputs(1724) <= (inputs(25)) or (inputs(96));
    layer0_outputs(1725) <= (inputs(3)) xor (inputs(70));
    layer0_outputs(1726) <= (inputs(231)) xor (inputs(203));
    layer0_outputs(1727) <= inputs(10);
    layer0_outputs(1728) <= not((inputs(15)) or (inputs(101)));
    layer0_outputs(1729) <= not((inputs(143)) xor (inputs(99)));
    layer0_outputs(1730) <= inputs(106);
    layer0_outputs(1731) <= (inputs(181)) and not (inputs(144));
    layer0_outputs(1732) <= inputs(59);
    layer0_outputs(1733) <= (inputs(30)) and not (inputs(160));
    layer0_outputs(1734) <= not(inputs(118)) or (inputs(218));
    layer0_outputs(1735) <= not(inputs(66)) or (inputs(72));
    layer0_outputs(1736) <= '1';
    layer0_outputs(1737) <= (inputs(38)) and not (inputs(182));
    layer0_outputs(1738) <= not((inputs(102)) or (inputs(142)));
    layer0_outputs(1739) <= not(inputs(119)) or (inputs(128));
    layer0_outputs(1740) <= (inputs(158)) xor (inputs(144));
    layer0_outputs(1741) <= not(inputs(98));
    layer0_outputs(1742) <= inputs(174);
    layer0_outputs(1743) <= not((inputs(42)) or (inputs(99)));
    layer0_outputs(1744) <= not(inputs(234));
    layer0_outputs(1745) <= not((inputs(116)) or (inputs(114)));
    layer0_outputs(1746) <= not(inputs(179)) or (inputs(112));
    layer0_outputs(1747) <= not((inputs(252)) xor (inputs(179)));
    layer0_outputs(1748) <= not(inputs(121)) or (inputs(141));
    layer0_outputs(1749) <= not((inputs(108)) xor (inputs(190)));
    layer0_outputs(1750) <= not(inputs(67)) or (inputs(64));
    layer0_outputs(1751) <= not((inputs(2)) or (inputs(43)));
    layer0_outputs(1752) <= inputs(106);
    layer0_outputs(1753) <= (inputs(87)) xor (inputs(143));
    layer0_outputs(1754) <= not(inputs(68));
    layer0_outputs(1755) <= inputs(26);
    layer0_outputs(1756) <= (inputs(211)) or (inputs(41));
    layer0_outputs(1757) <= not(inputs(207)) or (inputs(195));
    layer0_outputs(1758) <= inputs(103);
    layer0_outputs(1759) <= (inputs(1)) xor (inputs(94));
    layer0_outputs(1760) <= not(inputs(152)) or (inputs(57));
    layer0_outputs(1761) <= not((inputs(226)) or (inputs(246)));
    layer0_outputs(1762) <= (inputs(217)) and not (inputs(64));
    layer0_outputs(1763) <= not(inputs(131));
    layer0_outputs(1764) <= (inputs(218)) xor (inputs(249));
    layer0_outputs(1765) <= inputs(108);
    layer0_outputs(1766) <= '1';
    layer0_outputs(1767) <= '1';
    layer0_outputs(1768) <= '1';
    layer0_outputs(1769) <= not(inputs(81));
    layer0_outputs(1770) <= not(inputs(200)) or (inputs(193));
    layer0_outputs(1771) <= not(inputs(103)) or (inputs(111));
    layer0_outputs(1772) <= not((inputs(239)) or (inputs(27)));
    layer0_outputs(1773) <= not((inputs(5)) xor (inputs(18)));
    layer0_outputs(1774) <= inputs(248);
    layer0_outputs(1775) <= (inputs(120)) xor (inputs(151));
    layer0_outputs(1776) <= inputs(90);
    layer0_outputs(1777) <= not(inputs(36)) or (inputs(160));
    layer0_outputs(1778) <= '0';
    layer0_outputs(1779) <= (inputs(197)) and not (inputs(219));
    layer0_outputs(1780) <= not((inputs(42)) or (inputs(170)));
    layer0_outputs(1781) <= inputs(237);
    layer0_outputs(1782) <= not((inputs(90)) or (inputs(238)));
    layer0_outputs(1783) <= not((inputs(221)) and (inputs(4)));
    layer0_outputs(1784) <= not(inputs(32)) or (inputs(199));
    layer0_outputs(1785) <= not(inputs(0));
    layer0_outputs(1786) <= not(inputs(35)) or (inputs(139));
    layer0_outputs(1787) <= inputs(154);
    layer0_outputs(1788) <= not(inputs(6));
    layer0_outputs(1789) <= not(inputs(101)) or (inputs(225));
    layer0_outputs(1790) <= (inputs(60)) and not (inputs(165));
    layer0_outputs(1791) <= (inputs(31)) or (inputs(171));
    layer0_outputs(1792) <= (inputs(0)) xor (inputs(224));
    layer0_outputs(1793) <= not(inputs(22));
    layer0_outputs(1794) <= not(inputs(102));
    layer0_outputs(1795) <= (inputs(160)) or (inputs(178));
    layer0_outputs(1796) <= (inputs(212)) or (inputs(173));
    layer0_outputs(1797) <= '0';
    layer0_outputs(1798) <= not((inputs(40)) or (inputs(141)));
    layer0_outputs(1799) <= not(inputs(78)) or (inputs(239));
    layer0_outputs(1800) <= not(inputs(79)) or (inputs(13));
    layer0_outputs(1801) <= (inputs(237)) or (inputs(74));
    layer0_outputs(1802) <= inputs(92);
    layer0_outputs(1803) <= inputs(164);
    layer0_outputs(1804) <= (inputs(95)) or (inputs(99));
    layer0_outputs(1805) <= (inputs(11)) and (inputs(223));
    layer0_outputs(1806) <= (inputs(167)) and not (inputs(96));
    layer0_outputs(1807) <= not((inputs(37)) or (inputs(142)));
    layer0_outputs(1808) <= inputs(162);
    layer0_outputs(1809) <= (inputs(173)) and not (inputs(24));
    layer0_outputs(1810) <= not((inputs(221)) or (inputs(231)));
    layer0_outputs(1811) <= not((inputs(97)) xor (inputs(140)));
    layer0_outputs(1812) <= (inputs(180)) and not (inputs(2));
    layer0_outputs(1813) <= (inputs(27)) or (inputs(172));
    layer0_outputs(1814) <= not(inputs(45));
    layer0_outputs(1815) <= not(inputs(8));
    layer0_outputs(1816) <= (inputs(28)) xor (inputs(62));
    layer0_outputs(1817) <= inputs(165);
    layer0_outputs(1818) <= (inputs(80)) or (inputs(144));
    layer0_outputs(1819) <= (inputs(155)) xor (inputs(199));
    layer0_outputs(1820) <= inputs(229);
    layer0_outputs(1821) <= (inputs(231)) xor (inputs(255));
    layer0_outputs(1822) <= (inputs(123)) xor (inputs(166));
    layer0_outputs(1823) <= not((inputs(33)) or (inputs(214)));
    layer0_outputs(1824) <= not(inputs(106));
    layer0_outputs(1825) <= (inputs(244)) xor (inputs(226));
    layer0_outputs(1826) <= not(inputs(22));
    layer0_outputs(1827) <= inputs(189);
    layer0_outputs(1828) <= not(inputs(213)) or (inputs(152));
    layer0_outputs(1829) <= (inputs(174)) or (inputs(137));
    layer0_outputs(1830) <= not((inputs(116)) or (inputs(130)));
    layer0_outputs(1831) <= not((inputs(160)) xor (inputs(74)));
    layer0_outputs(1832) <= not(inputs(186));
    layer0_outputs(1833) <= not(inputs(239)) or (inputs(109));
    layer0_outputs(1834) <= (inputs(92)) and not (inputs(81));
    layer0_outputs(1835) <= not(inputs(41));
    layer0_outputs(1836) <= inputs(108);
    layer0_outputs(1837) <= not(inputs(35)) or (inputs(145));
    layer0_outputs(1838) <= not((inputs(135)) xor (inputs(1)));
    layer0_outputs(1839) <= inputs(102);
    layer0_outputs(1840) <= not(inputs(195)) or (inputs(222));
    layer0_outputs(1841) <= (inputs(84)) or (inputs(100));
    layer0_outputs(1842) <= (inputs(119)) xor (inputs(201));
    layer0_outputs(1843) <= not((inputs(52)) or (inputs(65)));
    layer0_outputs(1844) <= not((inputs(205)) xor (inputs(165)));
    layer0_outputs(1845) <= (inputs(108)) and not (inputs(188));
    layer0_outputs(1846) <= not((inputs(139)) xor (inputs(113)));
    layer0_outputs(1847) <= not(inputs(90)) or (inputs(206));
    layer0_outputs(1848) <= (inputs(85)) or (inputs(96));
    layer0_outputs(1849) <= not(inputs(180)) or (inputs(113));
    layer0_outputs(1850) <= (inputs(109)) and not (inputs(255));
    layer0_outputs(1851) <= (inputs(54)) and not (inputs(239));
    layer0_outputs(1852) <= not((inputs(155)) or (inputs(28)));
    layer0_outputs(1853) <= not((inputs(144)) xor (inputs(182)));
    layer0_outputs(1854) <= not(inputs(91));
    layer0_outputs(1855) <= (inputs(58)) or (inputs(6));
    layer0_outputs(1856) <= inputs(194);
    layer0_outputs(1857) <= inputs(40);
    layer0_outputs(1858) <= (inputs(182)) or (inputs(85));
    layer0_outputs(1859) <= inputs(158);
    layer0_outputs(1860) <= not((inputs(229)) or (inputs(95)));
    layer0_outputs(1861) <= not((inputs(148)) xor (inputs(117)));
    layer0_outputs(1862) <= (inputs(231)) xor (inputs(16));
    layer0_outputs(1863) <= (inputs(36)) and not (inputs(55));
    layer0_outputs(1864) <= not(inputs(163));
    layer0_outputs(1865) <= (inputs(195)) xor (inputs(194));
    layer0_outputs(1866) <= not(inputs(51));
    layer0_outputs(1867) <= not((inputs(12)) or (inputs(15)));
    layer0_outputs(1868) <= inputs(139);
    layer0_outputs(1869) <= not(inputs(74));
    layer0_outputs(1870) <= (inputs(234)) or (inputs(65));
    layer0_outputs(1871) <= not((inputs(140)) or (inputs(23)));
    layer0_outputs(1872) <= (inputs(192)) or (inputs(237));
    layer0_outputs(1873) <= inputs(231);
    layer0_outputs(1874) <= not((inputs(0)) or (inputs(184)));
    layer0_outputs(1875) <= inputs(149);
    layer0_outputs(1876) <= not((inputs(226)) or (inputs(202)));
    layer0_outputs(1877) <= (inputs(216)) or (inputs(224));
    layer0_outputs(1878) <= not(inputs(198));
    layer0_outputs(1879) <= inputs(9);
    layer0_outputs(1880) <= (inputs(39)) and not (inputs(208));
    layer0_outputs(1881) <= (inputs(195)) and not (inputs(202));
    layer0_outputs(1882) <= inputs(163);
    layer0_outputs(1883) <= not((inputs(0)) or (inputs(171)));
    layer0_outputs(1884) <= inputs(47);
    layer0_outputs(1885) <= not((inputs(118)) xor (inputs(235)));
    layer0_outputs(1886) <= not((inputs(168)) or (inputs(120)));
    layer0_outputs(1887) <= not(inputs(248));
    layer0_outputs(1888) <= inputs(60);
    layer0_outputs(1889) <= inputs(227);
    layer0_outputs(1890) <= not(inputs(118));
    layer0_outputs(1891) <= (inputs(244)) xor (inputs(24));
    layer0_outputs(1892) <= not((inputs(1)) or (inputs(220)));
    layer0_outputs(1893) <= (inputs(29)) xor (inputs(190));
    layer0_outputs(1894) <= inputs(104);
    layer0_outputs(1895) <= (inputs(36)) and not (inputs(124));
    layer0_outputs(1896) <= '1';
    layer0_outputs(1897) <= (inputs(18)) and not (inputs(251));
    layer0_outputs(1898) <= (inputs(228)) and not (inputs(205));
    layer0_outputs(1899) <= not((inputs(38)) xor (inputs(128)));
    layer0_outputs(1900) <= not(inputs(232));
    layer0_outputs(1901) <= not((inputs(214)) or (inputs(191)));
    layer0_outputs(1902) <= not(inputs(169));
    layer0_outputs(1903) <= inputs(195);
    layer0_outputs(1904) <= not(inputs(42));
    layer0_outputs(1905) <= not(inputs(136));
    layer0_outputs(1906) <= not(inputs(38));
    layer0_outputs(1907) <= not(inputs(104)) or (inputs(34));
    layer0_outputs(1908) <= not(inputs(246)) or (inputs(252));
    layer0_outputs(1909) <= inputs(8);
    layer0_outputs(1910) <= (inputs(66)) or (inputs(137));
    layer0_outputs(1911) <= not(inputs(162));
    layer0_outputs(1912) <= (inputs(171)) xor (inputs(112));
    layer0_outputs(1913) <= (inputs(2)) or (inputs(6));
    layer0_outputs(1914) <= (inputs(89)) and not (inputs(232));
    layer0_outputs(1915) <= (inputs(115)) and not (inputs(254));
    layer0_outputs(1916) <= (inputs(213)) and (inputs(216));
    layer0_outputs(1917) <= (inputs(117)) and not (inputs(17));
    layer0_outputs(1918) <= (inputs(2)) or (inputs(51));
    layer0_outputs(1919) <= not((inputs(243)) or (inputs(201)));
    layer0_outputs(1920) <= inputs(175);
    layer0_outputs(1921) <= (inputs(233)) or (inputs(206));
    layer0_outputs(1922) <= (inputs(124)) and not (inputs(84));
    layer0_outputs(1923) <= inputs(65);
    layer0_outputs(1924) <= not(inputs(228));
    layer0_outputs(1925) <= not(inputs(27)) or (inputs(108));
    layer0_outputs(1926) <= not(inputs(202)) or (inputs(111));
    layer0_outputs(1927) <= inputs(183);
    layer0_outputs(1928) <= not((inputs(77)) or (inputs(215)));
    layer0_outputs(1929) <= not((inputs(246)) or (inputs(111)));
    layer0_outputs(1930) <= not((inputs(220)) xor (inputs(237)));
    layer0_outputs(1931) <= not((inputs(157)) and (inputs(37)));
    layer0_outputs(1932) <= not(inputs(208)) or (inputs(45));
    layer0_outputs(1933) <= inputs(7);
    layer0_outputs(1934) <= inputs(67);
    layer0_outputs(1935) <= not(inputs(73)) or (inputs(224));
    layer0_outputs(1936) <= not(inputs(178)) or (inputs(205));
    layer0_outputs(1937) <= (inputs(150)) and not (inputs(96));
    layer0_outputs(1938) <= (inputs(177)) or (inputs(191));
    layer0_outputs(1939) <= inputs(78);
    layer0_outputs(1940) <= inputs(58);
    layer0_outputs(1941) <= not(inputs(149));
    layer0_outputs(1942) <= inputs(166);
    layer0_outputs(1943) <= not((inputs(144)) or (inputs(70)));
    layer0_outputs(1944) <= not((inputs(235)) or (inputs(251)));
    layer0_outputs(1945) <= not((inputs(222)) and (inputs(193)));
    layer0_outputs(1946) <= not((inputs(142)) xor (inputs(129)));
    layer0_outputs(1947) <= (inputs(192)) and not (inputs(97));
    layer0_outputs(1948) <= (inputs(62)) or (inputs(205));
    layer0_outputs(1949) <= (inputs(128)) and not (inputs(224));
    layer0_outputs(1950) <= inputs(105);
    layer0_outputs(1951) <= inputs(247);
    layer0_outputs(1952) <= not(inputs(92));
    layer0_outputs(1953) <= inputs(249);
    layer0_outputs(1954) <= (inputs(113)) or (inputs(212));
    layer0_outputs(1955) <= inputs(24);
    layer0_outputs(1956) <= inputs(88);
    layer0_outputs(1957) <= not(inputs(171)) or (inputs(20));
    layer0_outputs(1958) <= not(inputs(84));
    layer0_outputs(1959) <= not(inputs(190));
    layer0_outputs(1960) <= (inputs(63)) or (inputs(134));
    layer0_outputs(1961) <= not(inputs(25));
    layer0_outputs(1962) <= not((inputs(19)) xor (inputs(100)));
    layer0_outputs(1963) <= (inputs(243)) xor (inputs(211));
    layer0_outputs(1964) <= (inputs(0)) or (inputs(181));
    layer0_outputs(1965) <= inputs(115);
    layer0_outputs(1966) <= not(inputs(232)) or (inputs(123));
    layer0_outputs(1967) <= inputs(155);
    layer0_outputs(1968) <= (inputs(49)) or (inputs(245));
    layer0_outputs(1969) <= '1';
    layer0_outputs(1970) <= (inputs(10)) and not (inputs(33));
    layer0_outputs(1971) <= (inputs(105)) or (inputs(19));
    layer0_outputs(1972) <= not(inputs(215));
    layer0_outputs(1973) <= not(inputs(59)) or (inputs(158));
    layer0_outputs(1974) <= not((inputs(109)) xor (inputs(188)));
    layer0_outputs(1975) <= not(inputs(164));
    layer0_outputs(1976) <= not(inputs(99));
    layer0_outputs(1977) <= not(inputs(162));
    layer0_outputs(1978) <= not(inputs(71));
    layer0_outputs(1979) <= not((inputs(185)) xor (inputs(181)));
    layer0_outputs(1980) <= not((inputs(198)) xor (inputs(60)));
    layer0_outputs(1981) <= '0';
    layer0_outputs(1982) <= inputs(98);
    layer0_outputs(1983) <= (inputs(218)) or (inputs(134));
    layer0_outputs(1984) <= not(inputs(136)) or (inputs(191));
    layer0_outputs(1985) <= (inputs(47)) or (inputs(230));
    layer0_outputs(1986) <= not(inputs(119)) or (inputs(129));
    layer0_outputs(1987) <= inputs(8);
    layer0_outputs(1988) <= not((inputs(173)) and (inputs(218)));
    layer0_outputs(1989) <= not((inputs(255)) or (inputs(101)));
    layer0_outputs(1990) <= (inputs(236)) xor (inputs(138));
    layer0_outputs(1991) <= inputs(122);
    layer0_outputs(1992) <= not(inputs(193));
    layer0_outputs(1993) <= (inputs(35)) xor (inputs(120));
    layer0_outputs(1994) <= (inputs(87)) xor (inputs(31));
    layer0_outputs(1995) <= not((inputs(173)) xor (inputs(219)));
    layer0_outputs(1996) <= (inputs(124)) and not (inputs(150));
    layer0_outputs(1997) <= not(inputs(232));
    layer0_outputs(1998) <= (inputs(249)) or (inputs(147));
    layer0_outputs(1999) <= inputs(91);
    layer0_outputs(2000) <= not(inputs(190));
    layer0_outputs(2001) <= not((inputs(40)) and (inputs(232)));
    layer0_outputs(2002) <= (inputs(71)) and (inputs(245));
    layer0_outputs(2003) <= not(inputs(161));
    layer0_outputs(2004) <= not((inputs(50)) or (inputs(117)));
    layer0_outputs(2005) <= inputs(108);
    layer0_outputs(2006) <= not((inputs(81)) xor (inputs(69)));
    layer0_outputs(2007) <= not(inputs(51)) or (inputs(244));
    layer0_outputs(2008) <= inputs(204);
    layer0_outputs(2009) <= (inputs(155)) and not (inputs(95));
    layer0_outputs(2010) <= not(inputs(54));
    layer0_outputs(2011) <= (inputs(167)) and not (inputs(56));
    layer0_outputs(2012) <= (inputs(156)) xor (inputs(22));
    layer0_outputs(2013) <= (inputs(6)) and not (inputs(157));
    layer0_outputs(2014) <= inputs(233);
    layer0_outputs(2015) <= inputs(58);
    layer0_outputs(2016) <= (inputs(107)) and (inputs(28));
    layer0_outputs(2017) <= (inputs(150)) or (inputs(129));
    layer0_outputs(2018) <= (inputs(203)) and not (inputs(240));
    layer0_outputs(2019) <= (inputs(5)) or (inputs(191));
    layer0_outputs(2020) <= not((inputs(72)) or (inputs(88)));
    layer0_outputs(2021) <= inputs(117);
    layer0_outputs(2022) <= not((inputs(205)) or (inputs(99)));
    layer0_outputs(2023) <= not(inputs(116)) or (inputs(235));
    layer0_outputs(2024) <= not(inputs(166));
    layer0_outputs(2025) <= not((inputs(183)) xor (inputs(188)));
    layer0_outputs(2026) <= (inputs(131)) or (inputs(206));
    layer0_outputs(2027) <= (inputs(48)) xor (inputs(85));
    layer0_outputs(2028) <= (inputs(123)) xor (inputs(110));
    layer0_outputs(2029) <= inputs(0);
    layer0_outputs(2030) <= (inputs(144)) or (inputs(173));
    layer0_outputs(2031) <= inputs(44);
    layer0_outputs(2032) <= not((inputs(76)) and (inputs(76)));
    layer0_outputs(2033) <= not(inputs(227)) or (inputs(94));
    layer0_outputs(2034) <= (inputs(250)) or (inputs(238));
    layer0_outputs(2035) <= not(inputs(224));
    layer0_outputs(2036) <= not((inputs(199)) or (inputs(207)));
    layer0_outputs(2037) <= inputs(204);
    layer0_outputs(2038) <= inputs(24);
    layer0_outputs(2039) <= not(inputs(196));
    layer0_outputs(2040) <= not((inputs(87)) or (inputs(173)));
    layer0_outputs(2041) <= inputs(132);
    layer0_outputs(2042) <= inputs(136);
    layer0_outputs(2043) <= '1';
    layer0_outputs(2044) <= not(inputs(106));
    layer0_outputs(2045) <= not((inputs(112)) and (inputs(134)));
    layer0_outputs(2046) <= (inputs(39)) and not (inputs(210));
    layer0_outputs(2047) <= not(inputs(108));
    layer0_outputs(2048) <= (inputs(140)) and not (inputs(28));
    layer0_outputs(2049) <= not((inputs(93)) xor (inputs(77)));
    layer0_outputs(2050) <= (inputs(124)) and not (inputs(29));
    layer0_outputs(2051) <= (inputs(105)) xor (inputs(125));
    layer0_outputs(2052) <= not((inputs(145)) or (inputs(146)));
    layer0_outputs(2053) <= (inputs(216)) and not (inputs(31));
    layer0_outputs(2054) <= not(inputs(88)) or (inputs(204));
    layer0_outputs(2055) <= not(inputs(48));
    layer0_outputs(2056) <= (inputs(139)) xor (inputs(169));
    layer0_outputs(2057) <= not(inputs(134)) or (inputs(33));
    layer0_outputs(2058) <= not((inputs(38)) or (inputs(16)));
    layer0_outputs(2059) <= not(inputs(248)) or (inputs(119));
    layer0_outputs(2060) <= (inputs(87)) xor (inputs(98));
    layer0_outputs(2061) <= not((inputs(14)) or (inputs(150)));
    layer0_outputs(2062) <= not((inputs(7)) xor (inputs(80)));
    layer0_outputs(2063) <= (inputs(89)) and not (inputs(216));
    layer0_outputs(2064) <= not((inputs(60)) or (inputs(254)));
    layer0_outputs(2065) <= inputs(179);
    layer0_outputs(2066) <= (inputs(186)) and not (inputs(15));
    layer0_outputs(2067) <= (inputs(239)) or (inputs(65));
    layer0_outputs(2068) <= not(inputs(104));
    layer0_outputs(2069) <= not(inputs(154)) or (inputs(50));
    layer0_outputs(2070) <= inputs(230);
    layer0_outputs(2071) <= inputs(141);
    layer0_outputs(2072) <= (inputs(164)) xor (inputs(250));
    layer0_outputs(2073) <= not((inputs(94)) or (inputs(68)));
    layer0_outputs(2074) <= inputs(215);
    layer0_outputs(2075) <= not(inputs(40)) or (inputs(235));
    layer0_outputs(2076) <= (inputs(90)) xor (inputs(141));
    layer0_outputs(2077) <= not(inputs(220)) or (inputs(63));
    layer0_outputs(2078) <= (inputs(202)) and not (inputs(30));
    layer0_outputs(2079) <= '1';
    layer0_outputs(2080) <= '0';
    layer0_outputs(2081) <= not(inputs(24)) or (inputs(146));
    layer0_outputs(2082) <= not((inputs(153)) or (inputs(241)));
    layer0_outputs(2083) <= (inputs(141)) or (inputs(60));
    layer0_outputs(2084) <= not(inputs(109)) or (inputs(33));
    layer0_outputs(2085) <= not((inputs(181)) xor (inputs(176)));
    layer0_outputs(2086) <= '0';
    layer0_outputs(2087) <= not(inputs(89));
    layer0_outputs(2088) <= inputs(208);
    layer0_outputs(2089) <= inputs(54);
    layer0_outputs(2090) <= inputs(164);
    layer0_outputs(2091) <= not(inputs(209));
    layer0_outputs(2092) <= (inputs(121)) and (inputs(134));
    layer0_outputs(2093) <= not(inputs(37)) or (inputs(160));
    layer0_outputs(2094) <= inputs(229);
    layer0_outputs(2095) <= (inputs(229)) and (inputs(227));
    layer0_outputs(2096) <= not(inputs(67)) or (inputs(197));
    layer0_outputs(2097) <= (inputs(191)) or (inputs(114));
    layer0_outputs(2098) <= (inputs(220)) or (inputs(193));
    layer0_outputs(2099) <= not(inputs(166));
    layer0_outputs(2100) <= not(inputs(233)) or (inputs(195));
    layer0_outputs(2101) <= not(inputs(181)) or (inputs(5));
    layer0_outputs(2102) <= (inputs(42)) xor (inputs(7));
    layer0_outputs(2103) <= not(inputs(253));
    layer0_outputs(2104) <= (inputs(232)) and not (inputs(137));
    layer0_outputs(2105) <= not(inputs(161));
    layer0_outputs(2106) <= not(inputs(31));
    layer0_outputs(2107) <= inputs(181);
    layer0_outputs(2108) <= (inputs(170)) and not (inputs(241));
    layer0_outputs(2109) <= (inputs(205)) and not (inputs(94));
    layer0_outputs(2110) <= not(inputs(186));
    layer0_outputs(2111) <= not(inputs(41));
    layer0_outputs(2112) <= not((inputs(222)) or (inputs(71)));
    layer0_outputs(2113) <= not(inputs(8));
    layer0_outputs(2114) <= not((inputs(175)) and (inputs(134)));
    layer0_outputs(2115) <= '0';
    layer0_outputs(2116) <= (inputs(163)) and not (inputs(47));
    layer0_outputs(2117) <= inputs(68);
    layer0_outputs(2118) <= not(inputs(81)) or (inputs(186));
    layer0_outputs(2119) <= not(inputs(219));
    layer0_outputs(2120) <= not(inputs(91));
    layer0_outputs(2121) <= not(inputs(4)) or (inputs(146));
    layer0_outputs(2122) <= (inputs(148)) or (inputs(149));
    layer0_outputs(2123) <= not((inputs(206)) xor (inputs(174)));
    layer0_outputs(2124) <= (inputs(134)) and not (inputs(76));
    layer0_outputs(2125) <= (inputs(250)) and not (inputs(150));
    layer0_outputs(2126) <= not((inputs(74)) xor (inputs(14)));
    layer0_outputs(2127) <= not(inputs(93));
    layer0_outputs(2128) <= not(inputs(180)) or (inputs(127));
    layer0_outputs(2129) <= inputs(196);
    layer0_outputs(2130) <= not(inputs(203)) or (inputs(50));
    layer0_outputs(2131) <= (inputs(211)) and not (inputs(37));
    layer0_outputs(2132) <= inputs(19);
    layer0_outputs(2133) <= (inputs(63)) or (inputs(180));
    layer0_outputs(2134) <= not((inputs(252)) or (inputs(94)));
    layer0_outputs(2135) <= inputs(92);
    layer0_outputs(2136) <= not((inputs(118)) and (inputs(200)));
    layer0_outputs(2137) <= (inputs(61)) or (inputs(21));
    layer0_outputs(2138) <= not(inputs(20));
    layer0_outputs(2139) <= not(inputs(104));
    layer0_outputs(2140) <= not(inputs(8)) or (inputs(166));
    layer0_outputs(2141) <= (inputs(175)) or (inputs(64));
    layer0_outputs(2142) <= (inputs(243)) xor (inputs(16));
    layer0_outputs(2143) <= (inputs(146)) xor (inputs(232));
    layer0_outputs(2144) <= not(inputs(147)) or (inputs(77));
    layer0_outputs(2145) <= (inputs(12)) xor (inputs(46));
    layer0_outputs(2146) <= (inputs(156)) or (inputs(102));
    layer0_outputs(2147) <= not((inputs(204)) or (inputs(215)));
    layer0_outputs(2148) <= not((inputs(165)) or (inputs(191)));
    layer0_outputs(2149) <= not((inputs(238)) xor (inputs(49)));
    layer0_outputs(2150) <= not((inputs(57)) xor (inputs(233)));
    layer0_outputs(2151) <= not(inputs(195));
    layer0_outputs(2152) <= inputs(130);
    layer0_outputs(2153) <= (inputs(73)) xor (inputs(56));
    layer0_outputs(2154) <= not(inputs(147));
    layer0_outputs(2155) <= not(inputs(28)) or (inputs(159));
    layer0_outputs(2156) <= (inputs(119)) or (inputs(136));
    layer0_outputs(2157) <= (inputs(200)) and not (inputs(89));
    layer0_outputs(2158) <= (inputs(134)) and not (inputs(180));
    layer0_outputs(2159) <= (inputs(32)) or (inputs(21));
    layer0_outputs(2160) <= '1';
    layer0_outputs(2161) <= not(inputs(9));
    layer0_outputs(2162) <= inputs(45);
    layer0_outputs(2163) <= (inputs(200)) and not (inputs(21));
    layer0_outputs(2164) <= (inputs(105)) or (inputs(135));
    layer0_outputs(2165) <= inputs(136);
    layer0_outputs(2166) <= not((inputs(184)) xor (inputs(2)));
    layer0_outputs(2167) <= not((inputs(158)) or (inputs(142)));
    layer0_outputs(2168) <= (inputs(75)) xor (inputs(181));
    layer0_outputs(2169) <= not((inputs(214)) and (inputs(28)));
    layer0_outputs(2170) <= inputs(183);
    layer0_outputs(2171) <= (inputs(141)) or (inputs(219));
    layer0_outputs(2172) <= (inputs(129)) or (inputs(154));
    layer0_outputs(2173) <= inputs(173);
    layer0_outputs(2174) <= inputs(2);
    layer0_outputs(2175) <= not((inputs(170)) xor (inputs(119)));
    layer0_outputs(2176) <= (inputs(66)) or (inputs(13));
    layer0_outputs(2177) <= not((inputs(3)) or (inputs(224)));
    layer0_outputs(2178) <= not(inputs(59)) or (inputs(146));
    layer0_outputs(2179) <= not((inputs(71)) xor (inputs(97)));
    layer0_outputs(2180) <= not(inputs(92)) or (inputs(174));
    layer0_outputs(2181) <= not(inputs(202));
    layer0_outputs(2182) <= not(inputs(187)) or (inputs(17));
    layer0_outputs(2183) <= inputs(235);
    layer0_outputs(2184) <= (inputs(140)) or (inputs(208));
    layer0_outputs(2185) <= inputs(34);
    layer0_outputs(2186) <= not(inputs(161));
    layer0_outputs(2187) <= not((inputs(104)) and (inputs(106)));
    layer0_outputs(2188) <= not(inputs(176));
    layer0_outputs(2189) <= not(inputs(1));
    layer0_outputs(2190) <= not((inputs(187)) or (inputs(49)));
    layer0_outputs(2191) <= not(inputs(187)) or (inputs(37));
    layer0_outputs(2192) <= inputs(70);
    layer0_outputs(2193) <= inputs(10);
    layer0_outputs(2194) <= (inputs(211)) and not (inputs(89));
    layer0_outputs(2195) <= not((inputs(86)) xor (inputs(200)));
    layer0_outputs(2196) <= (inputs(238)) xor (inputs(210));
    layer0_outputs(2197) <= not(inputs(207));
    layer0_outputs(2198) <= not(inputs(204));
    layer0_outputs(2199) <= (inputs(57)) and not (inputs(83));
    layer0_outputs(2200) <= not(inputs(93));
    layer0_outputs(2201) <= '0';
    layer0_outputs(2202) <= (inputs(234)) and not (inputs(46));
    layer0_outputs(2203) <= (inputs(24)) and (inputs(228));
    layer0_outputs(2204) <= inputs(202);
    layer0_outputs(2205) <= (inputs(227)) and not (inputs(56));
    layer0_outputs(2206) <= not(inputs(245)) or (inputs(107));
    layer0_outputs(2207) <= (inputs(171)) and not (inputs(231));
    layer0_outputs(2208) <= (inputs(225)) or (inputs(148));
    layer0_outputs(2209) <= not(inputs(37)) or (inputs(96));
    layer0_outputs(2210) <= not(inputs(124));
    layer0_outputs(2211) <= (inputs(159)) or (inputs(92));
    layer0_outputs(2212) <= not(inputs(92)) or (inputs(34));
    layer0_outputs(2213) <= (inputs(40)) or (inputs(209));
    layer0_outputs(2214) <= not(inputs(72));
    layer0_outputs(2215) <= (inputs(11)) xor (inputs(29));
    layer0_outputs(2216) <= not(inputs(14)) or (inputs(254));
    layer0_outputs(2217) <= not((inputs(226)) xor (inputs(202)));
    layer0_outputs(2218) <= inputs(3);
    layer0_outputs(2219) <= '1';
    layer0_outputs(2220) <= not(inputs(210));
    layer0_outputs(2221) <= not((inputs(171)) xor (inputs(172)));
    layer0_outputs(2222) <= not((inputs(171)) or (inputs(117)));
    layer0_outputs(2223) <= inputs(161);
    layer0_outputs(2224) <= inputs(197);
    layer0_outputs(2225) <= (inputs(239)) xor (inputs(79));
    layer0_outputs(2226) <= not(inputs(219));
    layer0_outputs(2227) <= not(inputs(96)) or (inputs(190));
    layer0_outputs(2228) <= not(inputs(23));
    layer0_outputs(2229) <= not(inputs(102));
    layer0_outputs(2230) <= (inputs(186)) and not (inputs(63));
    layer0_outputs(2231) <= not((inputs(241)) xor (inputs(149)));
    layer0_outputs(2232) <= (inputs(49)) or (inputs(152));
    layer0_outputs(2233) <= not((inputs(57)) or (inputs(6)));
    layer0_outputs(2234) <= inputs(178);
    layer0_outputs(2235) <= (inputs(248)) or (inputs(16));
    layer0_outputs(2236) <= inputs(194);
    layer0_outputs(2237) <= not(inputs(23)) or (inputs(97));
    layer0_outputs(2238) <= inputs(58);
    layer0_outputs(2239) <= (inputs(196)) and (inputs(233));
    layer0_outputs(2240) <= not((inputs(208)) and (inputs(84)));
    layer0_outputs(2241) <= not((inputs(124)) or (inputs(9)));
    layer0_outputs(2242) <= inputs(141);
    layer0_outputs(2243) <= inputs(196);
    layer0_outputs(2244) <= (inputs(91)) or (inputs(4));
    layer0_outputs(2245) <= not((inputs(199)) or (inputs(30)));
    layer0_outputs(2246) <= not(inputs(93)) or (inputs(185));
    layer0_outputs(2247) <= not((inputs(93)) or (inputs(192)));
    layer0_outputs(2248) <= (inputs(236)) xor (inputs(158));
    layer0_outputs(2249) <= not(inputs(60));
    layer0_outputs(2250) <= not((inputs(18)) or (inputs(55)));
    layer0_outputs(2251) <= inputs(46);
    layer0_outputs(2252) <= (inputs(113)) or (inputs(34));
    layer0_outputs(2253) <= inputs(197);
    layer0_outputs(2254) <= not(inputs(151)) or (inputs(53));
    layer0_outputs(2255) <= not(inputs(236));
    layer0_outputs(2256) <= '0';
    layer0_outputs(2257) <= (inputs(141)) or (inputs(164));
    layer0_outputs(2258) <= (inputs(81)) and (inputs(54));
    layer0_outputs(2259) <= not((inputs(132)) or (inputs(15)));
    layer0_outputs(2260) <= (inputs(153)) and not (inputs(45));
    layer0_outputs(2261) <= (inputs(137)) xor (inputs(233));
    layer0_outputs(2262) <= (inputs(173)) and not (inputs(255));
    layer0_outputs(2263) <= (inputs(151)) and not (inputs(118));
    layer0_outputs(2264) <= not((inputs(123)) or (inputs(10)));
    layer0_outputs(2265) <= not((inputs(148)) xor (inputs(251)));
    layer0_outputs(2266) <= inputs(178);
    layer0_outputs(2267) <= (inputs(237)) and not (inputs(62));
    layer0_outputs(2268) <= not((inputs(11)) or (inputs(30)));
    layer0_outputs(2269) <= inputs(82);
    layer0_outputs(2270) <= not(inputs(24));
    layer0_outputs(2271) <= (inputs(172)) and not (inputs(181));
    layer0_outputs(2272) <= inputs(216);
    layer0_outputs(2273) <= (inputs(66)) and not (inputs(250));
    layer0_outputs(2274) <= not(inputs(197));
    layer0_outputs(2275) <= (inputs(115)) or (inputs(156));
    layer0_outputs(2276) <= inputs(223);
    layer0_outputs(2277) <= inputs(93);
    layer0_outputs(2278) <= inputs(83);
    layer0_outputs(2279) <= (inputs(130)) and not (inputs(80));
    layer0_outputs(2280) <= inputs(60);
    layer0_outputs(2281) <= (inputs(11)) or (inputs(96));
    layer0_outputs(2282) <= (inputs(78)) xor (inputs(2));
    layer0_outputs(2283) <= inputs(6);
    layer0_outputs(2284) <= inputs(40);
    layer0_outputs(2285) <= (inputs(119)) and not (inputs(17));
    layer0_outputs(2286) <= (inputs(138)) and not (inputs(212));
    layer0_outputs(2287) <= inputs(172);
    layer0_outputs(2288) <= not((inputs(176)) or (inputs(195)));
    layer0_outputs(2289) <= not(inputs(76)) or (inputs(158));
    layer0_outputs(2290) <= (inputs(75)) or (inputs(2));
    layer0_outputs(2291) <= (inputs(112)) or (inputs(117));
    layer0_outputs(2292) <= (inputs(78)) xor (inputs(157));
    layer0_outputs(2293) <= not(inputs(9));
    layer0_outputs(2294) <= not(inputs(119)) or (inputs(160));
    layer0_outputs(2295) <= '0';
    layer0_outputs(2296) <= (inputs(40)) xor (inputs(174));
    layer0_outputs(2297) <= (inputs(39)) and not (inputs(74));
    layer0_outputs(2298) <= (inputs(106)) and not (inputs(31));
    layer0_outputs(2299) <= inputs(19);
    layer0_outputs(2300) <= not((inputs(236)) xor (inputs(162)));
    layer0_outputs(2301) <= (inputs(157)) or (inputs(116));
    layer0_outputs(2302) <= inputs(115);
    layer0_outputs(2303) <= (inputs(11)) and not (inputs(150));
    layer0_outputs(2304) <= (inputs(30)) xor (inputs(137));
    layer0_outputs(2305) <= not(inputs(135)) or (inputs(213));
    layer0_outputs(2306) <= not((inputs(111)) xor (inputs(247)));
    layer0_outputs(2307) <= (inputs(38)) xor (inputs(59));
    layer0_outputs(2308) <= inputs(137);
    layer0_outputs(2309) <= (inputs(27)) and not (inputs(97));
    layer0_outputs(2310) <= not((inputs(250)) or (inputs(100)));
    layer0_outputs(2311) <= (inputs(21)) or (inputs(110));
    layer0_outputs(2312) <= (inputs(101)) and not (inputs(214));
    layer0_outputs(2313) <= inputs(133);
    layer0_outputs(2314) <= (inputs(6)) xor (inputs(53));
    layer0_outputs(2315) <= not(inputs(23));
    layer0_outputs(2316) <= not(inputs(89)) or (inputs(211));
    layer0_outputs(2317) <= (inputs(158)) or (inputs(215));
    layer0_outputs(2318) <= (inputs(117)) or (inputs(234));
    layer0_outputs(2319) <= not(inputs(191));
    layer0_outputs(2320) <= not(inputs(107)) or (inputs(228));
    layer0_outputs(2321) <= (inputs(165)) and not (inputs(160));
    layer0_outputs(2322) <= not(inputs(193)) or (inputs(128));
    layer0_outputs(2323) <= not(inputs(55)) or (inputs(49));
    layer0_outputs(2324) <= (inputs(196)) or (inputs(240));
    layer0_outputs(2325) <= not(inputs(124)) or (inputs(197));
    layer0_outputs(2326) <= not(inputs(40));
    layer0_outputs(2327) <= inputs(85);
    layer0_outputs(2328) <= inputs(225);
    layer0_outputs(2329) <= inputs(204);
    layer0_outputs(2330) <= inputs(234);
    layer0_outputs(2331) <= not(inputs(70));
    layer0_outputs(2332) <= (inputs(209)) or (inputs(246));
    layer0_outputs(2333) <= (inputs(75)) and not (inputs(203));
    layer0_outputs(2334) <= inputs(8);
    layer0_outputs(2335) <= not(inputs(38));
    layer0_outputs(2336) <= not(inputs(40)) or (inputs(34));
    layer0_outputs(2337) <= (inputs(148)) or (inputs(102));
    layer0_outputs(2338) <= not((inputs(158)) or (inputs(112)));
    layer0_outputs(2339) <= not(inputs(116)) or (inputs(50));
    layer0_outputs(2340) <= inputs(27);
    layer0_outputs(2341) <= (inputs(12)) or (inputs(224));
    layer0_outputs(2342) <= not((inputs(30)) or (inputs(140)));
    layer0_outputs(2343) <= inputs(135);
    layer0_outputs(2344) <= (inputs(33)) and not (inputs(228));
    layer0_outputs(2345) <= not((inputs(192)) or (inputs(196)));
    layer0_outputs(2346) <= not(inputs(130));
    layer0_outputs(2347) <= '1';
    layer0_outputs(2348) <= inputs(116);
    layer0_outputs(2349) <= not((inputs(29)) or (inputs(13)));
    layer0_outputs(2350) <= (inputs(35)) and not (inputs(31));
    layer0_outputs(2351) <= not((inputs(76)) xor (inputs(60)));
    layer0_outputs(2352) <= not(inputs(231));
    layer0_outputs(2353) <= inputs(65);
    layer0_outputs(2354) <= inputs(63);
    layer0_outputs(2355) <= not((inputs(235)) xor (inputs(177)));
    layer0_outputs(2356) <= not(inputs(57));
    layer0_outputs(2357) <= (inputs(195)) xor (inputs(119));
    layer0_outputs(2358) <= inputs(179);
    layer0_outputs(2359) <= (inputs(157)) or (inputs(187));
    layer0_outputs(2360) <= inputs(179);
    layer0_outputs(2361) <= (inputs(164)) xor (inputs(145));
    layer0_outputs(2362) <= (inputs(228)) and not (inputs(175));
    layer0_outputs(2363) <= not(inputs(125)) or (inputs(249));
    layer0_outputs(2364) <= (inputs(45)) and not (inputs(238));
    layer0_outputs(2365) <= inputs(11);
    layer0_outputs(2366) <= (inputs(70)) or (inputs(50));
    layer0_outputs(2367) <= not(inputs(235));
    layer0_outputs(2368) <= not(inputs(44)) or (inputs(10));
    layer0_outputs(2369) <= inputs(190);
    layer0_outputs(2370) <= not(inputs(251)) or (inputs(57));
    layer0_outputs(2371) <= not((inputs(50)) or (inputs(238)));
    layer0_outputs(2372) <= (inputs(150)) and not (inputs(1));
    layer0_outputs(2373) <= (inputs(100)) and not (inputs(227));
    layer0_outputs(2374) <= not((inputs(34)) and (inputs(131)));
    layer0_outputs(2375) <= not((inputs(213)) or (inputs(176)));
    layer0_outputs(2376) <= inputs(90);
    layer0_outputs(2377) <= not((inputs(133)) or (inputs(253)));
    layer0_outputs(2378) <= not(inputs(139));
    layer0_outputs(2379) <= not((inputs(47)) or (inputs(167)));
    layer0_outputs(2380) <= not((inputs(209)) xor (inputs(20)));
    layer0_outputs(2381) <= (inputs(65)) or (inputs(189));
    layer0_outputs(2382) <= not(inputs(72)) or (inputs(115));
    layer0_outputs(2383) <= not(inputs(100));
    layer0_outputs(2384) <= not(inputs(255)) or (inputs(223));
    layer0_outputs(2385) <= not(inputs(13));
    layer0_outputs(2386) <= (inputs(164)) and not (inputs(86));
    layer0_outputs(2387) <= (inputs(230)) and not (inputs(222));
    layer0_outputs(2388) <= not(inputs(125)) or (inputs(35));
    layer0_outputs(2389) <= not((inputs(8)) xor (inputs(110)));
    layer0_outputs(2390) <= inputs(55);
    layer0_outputs(2391) <= (inputs(64)) xor (inputs(106));
    layer0_outputs(2392) <= (inputs(249)) or (inputs(207));
    layer0_outputs(2393) <= (inputs(250)) and not (inputs(197));
    layer0_outputs(2394) <= (inputs(131)) or (inputs(49));
    layer0_outputs(2395) <= not(inputs(218)) or (inputs(59));
    layer0_outputs(2396) <= inputs(54);
    layer0_outputs(2397) <= (inputs(175)) or (inputs(244));
    layer0_outputs(2398) <= inputs(133);
    layer0_outputs(2399) <= not(inputs(49)) or (inputs(159));
    layer0_outputs(2400) <= not(inputs(75));
    layer0_outputs(2401) <= '1';
    layer0_outputs(2402) <= not(inputs(198));
    layer0_outputs(2403) <= (inputs(199)) and not (inputs(44));
    layer0_outputs(2404) <= inputs(189);
    layer0_outputs(2405) <= not(inputs(163));
    layer0_outputs(2406) <= not((inputs(205)) or (inputs(134)));
    layer0_outputs(2407) <= inputs(162);
    layer0_outputs(2408) <= (inputs(128)) and not (inputs(254));
    layer0_outputs(2409) <= not(inputs(59));
    layer0_outputs(2410) <= inputs(92);
    layer0_outputs(2411) <= inputs(139);
    layer0_outputs(2412) <= not(inputs(119));
    layer0_outputs(2413) <= not((inputs(28)) and (inputs(107)));
    layer0_outputs(2414) <= not(inputs(80));
    layer0_outputs(2415) <= not((inputs(244)) xor (inputs(197)));
    layer0_outputs(2416) <= not(inputs(99)) or (inputs(191));
    layer0_outputs(2417) <= not(inputs(245)) or (inputs(20));
    layer0_outputs(2418) <= inputs(216);
    layer0_outputs(2419) <= inputs(156);
    layer0_outputs(2420) <= (inputs(168)) and (inputs(212));
    layer0_outputs(2421) <= (inputs(8)) or (inputs(223));
    layer0_outputs(2422) <= inputs(210);
    layer0_outputs(2423) <= inputs(168);
    layer0_outputs(2424) <= (inputs(180)) or (inputs(13));
    layer0_outputs(2425) <= not((inputs(243)) and (inputs(36)));
    layer0_outputs(2426) <= inputs(102);
    layer0_outputs(2427) <= not(inputs(88)) or (inputs(18));
    layer0_outputs(2428) <= (inputs(48)) or (inputs(120));
    layer0_outputs(2429) <= not((inputs(209)) xor (inputs(246)));
    layer0_outputs(2430) <= not(inputs(181)) or (inputs(92));
    layer0_outputs(2431) <= not((inputs(43)) xor (inputs(70)));
    layer0_outputs(2432) <= inputs(193);
    layer0_outputs(2433) <= not(inputs(130));
    layer0_outputs(2434) <= not(inputs(101)) or (inputs(89));
    layer0_outputs(2435) <= not(inputs(83)) or (inputs(141));
    layer0_outputs(2436) <= not(inputs(84));
    layer0_outputs(2437) <= (inputs(31)) xor (inputs(44));
    layer0_outputs(2438) <= inputs(177);
    layer0_outputs(2439) <= not((inputs(51)) or (inputs(80)));
    layer0_outputs(2440) <= not(inputs(32));
    layer0_outputs(2441) <= (inputs(196)) xor (inputs(134));
    layer0_outputs(2442) <= not(inputs(173)) or (inputs(0));
    layer0_outputs(2443) <= (inputs(30)) and (inputs(34));
    layer0_outputs(2444) <= (inputs(30)) and not (inputs(177));
    layer0_outputs(2445) <= inputs(62);
    layer0_outputs(2446) <= (inputs(67)) and not (inputs(47));
    layer0_outputs(2447) <= not((inputs(133)) or (inputs(17)));
    layer0_outputs(2448) <= (inputs(93)) and not (inputs(240));
    layer0_outputs(2449) <= (inputs(62)) or (inputs(84));
    layer0_outputs(2450) <= (inputs(81)) xor (inputs(235));
    layer0_outputs(2451) <= (inputs(8)) and (inputs(119));
    layer0_outputs(2452) <= not((inputs(28)) or (inputs(31)));
    layer0_outputs(2453) <= inputs(129);
    layer0_outputs(2454) <= not(inputs(120));
    layer0_outputs(2455) <= not(inputs(120)) or (inputs(4));
    layer0_outputs(2456) <= inputs(86);
    layer0_outputs(2457) <= inputs(33);
    layer0_outputs(2458) <= (inputs(161)) and not (inputs(32));
    layer0_outputs(2459) <= not((inputs(146)) or (inputs(68)));
    layer0_outputs(2460) <= not(inputs(137)) or (inputs(48));
    layer0_outputs(2461) <= inputs(83);
    layer0_outputs(2462) <= not(inputs(180)) or (inputs(113));
    layer0_outputs(2463) <= not(inputs(78)) or (inputs(30));
    layer0_outputs(2464) <= inputs(246);
    layer0_outputs(2465) <= not((inputs(213)) and (inputs(139)));
    layer0_outputs(2466) <= not(inputs(152)) or (inputs(212));
    layer0_outputs(2467) <= (inputs(108)) xor (inputs(44));
    layer0_outputs(2468) <= not((inputs(181)) or (inputs(168)));
    layer0_outputs(2469) <= inputs(177);
    layer0_outputs(2470) <= (inputs(172)) xor (inputs(96));
    layer0_outputs(2471) <= not((inputs(65)) or (inputs(214)));
    layer0_outputs(2472) <= inputs(131);
    layer0_outputs(2473) <= not((inputs(183)) or (inputs(98)));
    layer0_outputs(2474) <= (inputs(96)) or (inputs(52));
    layer0_outputs(2475) <= inputs(220);
    layer0_outputs(2476) <= not(inputs(82));
    layer0_outputs(2477) <= not(inputs(206)) or (inputs(250));
    layer0_outputs(2478) <= not((inputs(240)) or (inputs(0)));
    layer0_outputs(2479) <= (inputs(126)) or (inputs(77));
    layer0_outputs(2480) <= (inputs(109)) or (inputs(4));
    layer0_outputs(2481) <= not(inputs(143)) or (inputs(253));
    layer0_outputs(2482) <= not((inputs(163)) xor (inputs(250)));
    layer0_outputs(2483) <= not((inputs(221)) or (inputs(120)));
    layer0_outputs(2484) <= inputs(238);
    layer0_outputs(2485) <= (inputs(209)) or (inputs(132));
    layer0_outputs(2486) <= inputs(234);
    layer0_outputs(2487) <= (inputs(203)) and not (inputs(254));
    layer0_outputs(2488) <= not(inputs(105)) or (inputs(39));
    layer0_outputs(2489) <= inputs(195);
    layer0_outputs(2490) <= (inputs(187)) or (inputs(220));
    layer0_outputs(2491) <= not(inputs(24)) or (inputs(113));
    layer0_outputs(2492) <= not(inputs(45)) or (inputs(191));
    layer0_outputs(2493) <= not((inputs(100)) or (inputs(250)));
    layer0_outputs(2494) <= inputs(211);
    layer0_outputs(2495) <= inputs(129);
    layer0_outputs(2496) <= not(inputs(211)) or (inputs(88));
    layer0_outputs(2497) <= not(inputs(74));
    layer0_outputs(2498) <= not(inputs(21)) or (inputs(228));
    layer0_outputs(2499) <= inputs(105);
    layer0_outputs(2500) <= (inputs(176)) and not (inputs(234));
    layer0_outputs(2501) <= (inputs(98)) and not (inputs(110));
    layer0_outputs(2502) <= (inputs(224)) and not (inputs(202));
    layer0_outputs(2503) <= (inputs(187)) or (inputs(170));
    layer0_outputs(2504) <= not((inputs(195)) or (inputs(9)));
    layer0_outputs(2505) <= (inputs(19)) and not (inputs(249));
    layer0_outputs(2506) <= inputs(215);
    layer0_outputs(2507) <= inputs(76);
    layer0_outputs(2508) <= not((inputs(137)) and (inputs(152)));
    layer0_outputs(2509) <= inputs(164);
    layer0_outputs(2510) <= inputs(27);
    layer0_outputs(2511) <= not(inputs(170));
    layer0_outputs(2512) <= not(inputs(181));
    layer0_outputs(2513) <= '0';
    layer0_outputs(2514) <= (inputs(22)) and not (inputs(129));
    layer0_outputs(2515) <= not(inputs(197)) or (inputs(81));
    layer0_outputs(2516) <= not(inputs(26)) or (inputs(25));
    layer0_outputs(2517) <= (inputs(214)) or (inputs(201));
    layer0_outputs(2518) <= (inputs(235)) or (inputs(221));
    layer0_outputs(2519) <= not((inputs(237)) or (inputs(116)));
    layer0_outputs(2520) <= (inputs(158)) and not (inputs(48));
    layer0_outputs(2521) <= (inputs(116)) or (inputs(205));
    layer0_outputs(2522) <= not(inputs(160));
    layer0_outputs(2523) <= '0';
    layer0_outputs(2524) <= not((inputs(184)) or (inputs(32)));
    layer0_outputs(2525) <= inputs(125);
    layer0_outputs(2526) <= (inputs(189)) or (inputs(129));
    layer0_outputs(2527) <= (inputs(79)) xor (inputs(192));
    layer0_outputs(2528) <= (inputs(73)) or (inputs(46));
    layer0_outputs(2529) <= not(inputs(153)) or (inputs(64));
    layer0_outputs(2530) <= not(inputs(107));
    layer0_outputs(2531) <= not(inputs(136)) or (inputs(179));
    layer0_outputs(2532) <= (inputs(228)) xor (inputs(213));
    layer0_outputs(2533) <= not((inputs(202)) or (inputs(14)));
    layer0_outputs(2534) <= inputs(230);
    layer0_outputs(2535) <= not(inputs(169)) or (inputs(168));
    layer0_outputs(2536) <= not((inputs(111)) xor (inputs(206)));
    layer0_outputs(2537) <= (inputs(120)) and not (inputs(22));
    layer0_outputs(2538) <= not((inputs(78)) or (inputs(230)));
    layer0_outputs(2539) <= not((inputs(128)) and (inputs(254)));
    layer0_outputs(2540) <= not((inputs(170)) or (inputs(112)));
    layer0_outputs(2541) <= (inputs(13)) xor (inputs(89));
    layer0_outputs(2542) <= not(inputs(243));
    layer0_outputs(2543) <= (inputs(91)) or (inputs(68));
    layer0_outputs(2544) <= not(inputs(148));
    layer0_outputs(2545) <= not(inputs(185)) or (inputs(120));
    layer0_outputs(2546) <= (inputs(68)) or (inputs(159));
    layer0_outputs(2547) <= not((inputs(254)) or (inputs(184)));
    layer0_outputs(2548) <= not(inputs(179));
    layer0_outputs(2549) <= not(inputs(209));
    layer0_outputs(2550) <= not(inputs(245));
    layer0_outputs(2551) <= (inputs(33)) or (inputs(174));
    layer0_outputs(2552) <= not(inputs(78));
    layer0_outputs(2553) <= not(inputs(170)) or (inputs(92));
    layer0_outputs(2554) <= (inputs(16)) or (inputs(2));
    layer0_outputs(2555) <= not(inputs(170));
    layer0_outputs(2556) <= (inputs(31)) and not (inputs(222));
    layer0_outputs(2557) <= '0';
    layer0_outputs(2558) <= '1';
    layer0_outputs(2559) <= (inputs(213)) and not (inputs(32));
    layer0_outputs(2560) <= (inputs(7)) xor (inputs(55));
    layer0_outputs(2561) <= inputs(177);
    layer0_outputs(2562) <= not(inputs(67)) or (inputs(188));
    layer0_outputs(2563) <= inputs(231);
    layer0_outputs(2564) <= inputs(127);
    layer0_outputs(2565) <= (inputs(199)) xor (inputs(202));
    layer0_outputs(2566) <= not(inputs(144));
    layer0_outputs(2567) <= (inputs(163)) and (inputs(136));
    layer0_outputs(2568) <= inputs(99);
    layer0_outputs(2569) <= inputs(230);
    layer0_outputs(2570) <= not((inputs(28)) xor (inputs(45)));
    layer0_outputs(2571) <= (inputs(132)) and (inputs(0));
    layer0_outputs(2572) <= not(inputs(124)) or (inputs(224));
    layer0_outputs(2573) <= (inputs(191)) or (inputs(168));
    layer0_outputs(2574) <= not(inputs(220)) or (inputs(67));
    layer0_outputs(2575) <= not(inputs(42));
    layer0_outputs(2576) <= '0';
    layer0_outputs(2577) <= not((inputs(48)) xor (inputs(0)));
    layer0_outputs(2578) <= inputs(101);
    layer0_outputs(2579) <= (inputs(26)) xor (inputs(114));
    layer0_outputs(2580) <= not((inputs(44)) or (inputs(27)));
    layer0_outputs(2581) <= (inputs(87)) and (inputs(23));
    layer0_outputs(2582) <= (inputs(104)) or (inputs(253));
    layer0_outputs(2583) <= (inputs(20)) xor (inputs(87));
    layer0_outputs(2584) <= not((inputs(127)) or (inputs(226)));
    layer0_outputs(2585) <= not(inputs(209));
    layer0_outputs(2586) <= not((inputs(102)) xor (inputs(144)));
    layer0_outputs(2587) <= (inputs(247)) and not (inputs(28));
    layer0_outputs(2588) <= not(inputs(16));
    layer0_outputs(2589) <= not(inputs(46)) or (inputs(221));
    layer0_outputs(2590) <= '0';
    layer0_outputs(2591) <= not((inputs(1)) or (inputs(175)));
    layer0_outputs(2592) <= not((inputs(244)) and (inputs(58)));
    layer0_outputs(2593) <= inputs(43);
    layer0_outputs(2594) <= '0';
    layer0_outputs(2595) <= not(inputs(198));
    layer0_outputs(2596) <= not((inputs(247)) and (inputs(138)));
    layer0_outputs(2597) <= not(inputs(43));
    layer0_outputs(2598) <= not(inputs(147));
    layer0_outputs(2599) <= (inputs(35)) and not (inputs(178));
    layer0_outputs(2600) <= not((inputs(67)) or (inputs(146)));
    layer0_outputs(2601) <= (inputs(248)) or (inputs(53));
    layer0_outputs(2602) <= (inputs(141)) and not (inputs(49));
    layer0_outputs(2603) <= inputs(232);
    layer0_outputs(2604) <= not((inputs(27)) xor (inputs(59)));
    layer0_outputs(2605) <= inputs(69);
    layer0_outputs(2606) <= not(inputs(69)) or (inputs(77));
    layer0_outputs(2607) <= not((inputs(10)) or (inputs(38)));
    layer0_outputs(2608) <= not((inputs(4)) xor (inputs(43)));
    layer0_outputs(2609) <= not(inputs(37));
    layer0_outputs(2610) <= inputs(25);
    layer0_outputs(2611) <= (inputs(21)) xor (inputs(246));
    layer0_outputs(2612) <= not(inputs(118));
    layer0_outputs(2613) <= (inputs(148)) or (inputs(201));
    layer0_outputs(2614) <= (inputs(191)) or (inputs(160));
    layer0_outputs(2615) <= inputs(150);
    layer0_outputs(2616) <= not(inputs(232));
    layer0_outputs(2617) <= not(inputs(33)) or (inputs(66));
    layer0_outputs(2618) <= inputs(150);
    layer0_outputs(2619) <= not(inputs(130));
    layer0_outputs(2620) <= (inputs(68)) xor (inputs(55));
    layer0_outputs(2621) <= not((inputs(183)) xor (inputs(151)));
    layer0_outputs(2622) <= inputs(25);
    layer0_outputs(2623) <= not(inputs(253)) or (inputs(207));
    layer0_outputs(2624) <= inputs(126);
    layer0_outputs(2625) <= (inputs(17)) xor (inputs(187));
    layer0_outputs(2626) <= (inputs(239)) or (inputs(250));
    layer0_outputs(2627) <= inputs(65);
    layer0_outputs(2628) <= not(inputs(175)) or (inputs(31));
    layer0_outputs(2629) <= (inputs(22)) and not (inputs(109));
    layer0_outputs(2630) <= not((inputs(34)) or (inputs(57)));
    layer0_outputs(2631) <= (inputs(227)) or (inputs(214));
    layer0_outputs(2632) <= inputs(61);
    layer0_outputs(2633) <= not(inputs(107));
    layer0_outputs(2634) <= '0';
    layer0_outputs(2635) <= not(inputs(231));
    layer0_outputs(2636) <= not(inputs(105));
    layer0_outputs(2637) <= inputs(121);
    layer0_outputs(2638) <= (inputs(13)) or (inputs(4));
    layer0_outputs(2639) <= not((inputs(42)) and (inputs(23)));
    layer0_outputs(2640) <= inputs(88);
    layer0_outputs(2641) <= not(inputs(214)) or (inputs(242));
    layer0_outputs(2642) <= (inputs(184)) xor (inputs(122));
    layer0_outputs(2643) <= not(inputs(196)) or (inputs(15));
    layer0_outputs(2644) <= (inputs(237)) and not (inputs(18));
    layer0_outputs(2645) <= inputs(114);
    layer0_outputs(2646) <= (inputs(152)) or (inputs(149));
    layer0_outputs(2647) <= not((inputs(118)) xor (inputs(178)));
    layer0_outputs(2648) <= (inputs(187)) xor (inputs(247));
    layer0_outputs(2649) <= (inputs(80)) xor (inputs(95));
    layer0_outputs(2650) <= not(inputs(135));
    layer0_outputs(2651) <= not(inputs(119)) or (inputs(194));
    layer0_outputs(2652) <= not(inputs(13));
    layer0_outputs(2653) <= inputs(212);
    layer0_outputs(2654) <= inputs(82);
    layer0_outputs(2655) <= (inputs(115)) and not (inputs(20));
    layer0_outputs(2656) <= not((inputs(82)) or (inputs(17)));
    layer0_outputs(2657) <= not((inputs(57)) xor (inputs(86)));
    layer0_outputs(2658) <= inputs(244);
    layer0_outputs(2659) <= not(inputs(184)) or (inputs(27));
    layer0_outputs(2660) <= (inputs(11)) and not (inputs(157));
    layer0_outputs(2661) <= (inputs(157)) or (inputs(158));
    layer0_outputs(2662) <= (inputs(136)) and not (inputs(216));
    layer0_outputs(2663) <= not(inputs(8)) or (inputs(250));
    layer0_outputs(2664) <= (inputs(88)) xor (inputs(119));
    layer0_outputs(2665) <= not((inputs(254)) or (inputs(211)));
    layer0_outputs(2666) <= (inputs(152)) and not (inputs(228));
    layer0_outputs(2667) <= not(inputs(157));
    layer0_outputs(2668) <= inputs(110);
    layer0_outputs(2669) <= not(inputs(214));
    layer0_outputs(2670) <= not(inputs(182));
    layer0_outputs(2671) <= not(inputs(153));
    layer0_outputs(2672) <= not(inputs(193));
    layer0_outputs(2673) <= not(inputs(149)) or (inputs(255));
    layer0_outputs(2674) <= not(inputs(248));
    layer0_outputs(2675) <= not((inputs(46)) or (inputs(132)));
    layer0_outputs(2676) <= not((inputs(105)) or (inputs(16)));
    layer0_outputs(2677) <= not((inputs(231)) and (inputs(77)));
    layer0_outputs(2678) <= (inputs(53)) and not (inputs(114));
    layer0_outputs(2679) <= not(inputs(57));
    layer0_outputs(2680) <= (inputs(56)) and not (inputs(23));
    layer0_outputs(2681) <= inputs(22);
    layer0_outputs(2682) <= inputs(226);
    layer0_outputs(2683) <= inputs(16);
    layer0_outputs(2684) <= '0';
    layer0_outputs(2685) <= inputs(132);
    layer0_outputs(2686) <= not((inputs(211)) or (inputs(121)));
    layer0_outputs(2687) <= (inputs(168)) or (inputs(7));
    layer0_outputs(2688) <= inputs(148);
    layer0_outputs(2689) <= not((inputs(57)) or (inputs(26)));
    layer0_outputs(2690) <= not(inputs(66));
    layer0_outputs(2691) <= not(inputs(22)) or (inputs(218));
    layer0_outputs(2692) <= (inputs(35)) and not (inputs(47));
    layer0_outputs(2693) <= (inputs(238)) or (inputs(165));
    layer0_outputs(2694) <= (inputs(47)) and not (inputs(240));
    layer0_outputs(2695) <= not((inputs(219)) or (inputs(202)));
    layer0_outputs(2696) <= not((inputs(190)) xor (inputs(172)));
    layer0_outputs(2697) <= (inputs(45)) and (inputs(61));
    layer0_outputs(2698) <= not(inputs(101));
    layer0_outputs(2699) <= not(inputs(150));
    layer0_outputs(2700) <= '1';
    layer0_outputs(2701) <= not(inputs(24));
    layer0_outputs(2702) <= not(inputs(252));
    layer0_outputs(2703) <= inputs(44);
    layer0_outputs(2704) <= not((inputs(180)) or (inputs(181)));
    layer0_outputs(2705) <= (inputs(238)) xor (inputs(139));
    layer0_outputs(2706) <= not(inputs(87));
    layer0_outputs(2707) <= not((inputs(37)) xor (inputs(157)));
    layer0_outputs(2708) <= inputs(85);
    layer0_outputs(2709) <= not((inputs(182)) and (inputs(215)));
    layer0_outputs(2710) <= not((inputs(153)) or (inputs(135)));
    layer0_outputs(2711) <= not(inputs(206));
    layer0_outputs(2712) <= not((inputs(100)) xor (inputs(5)));
    layer0_outputs(2713) <= not(inputs(238));
    layer0_outputs(2714) <= (inputs(58)) and not (inputs(29));
    layer0_outputs(2715) <= not(inputs(95));
    layer0_outputs(2716) <= not((inputs(233)) or (inputs(149)));
    layer0_outputs(2717) <= not(inputs(173)) or (inputs(0));
    layer0_outputs(2718) <= not((inputs(102)) xor (inputs(25)));
    layer0_outputs(2719) <= (inputs(89)) or (inputs(164));
    layer0_outputs(2720) <= not(inputs(217)) or (inputs(16));
    layer0_outputs(2721) <= not(inputs(211)) or (inputs(28));
    layer0_outputs(2722) <= not(inputs(232)) or (inputs(224));
    layer0_outputs(2723) <= (inputs(7)) and not (inputs(85));
    layer0_outputs(2724) <= (inputs(205)) and (inputs(222));
    layer0_outputs(2725) <= not(inputs(96));
    layer0_outputs(2726) <= inputs(177);
    layer0_outputs(2727) <= (inputs(49)) and not (inputs(21));
    layer0_outputs(2728) <= not((inputs(103)) or (inputs(238)));
    layer0_outputs(2729) <= (inputs(125)) or (inputs(9));
    layer0_outputs(2730) <= (inputs(199)) or (inputs(34));
    layer0_outputs(2731) <= not((inputs(163)) or (inputs(158)));
    layer0_outputs(2732) <= (inputs(39)) and (inputs(38));
    layer0_outputs(2733) <= not((inputs(127)) or (inputs(62)));
    layer0_outputs(2734) <= (inputs(105)) xor (inputs(76));
    layer0_outputs(2735) <= (inputs(173)) and (inputs(191));
    layer0_outputs(2736) <= not(inputs(218));
    layer0_outputs(2737) <= not(inputs(88)) or (inputs(24));
    layer0_outputs(2738) <= not(inputs(112));
    layer0_outputs(2739) <= not(inputs(39));
    layer0_outputs(2740) <= not(inputs(121)) or (inputs(154));
    layer0_outputs(2741) <= not(inputs(157));
    layer0_outputs(2742) <= not(inputs(210));
    layer0_outputs(2743) <= not(inputs(135)) or (inputs(207));
    layer0_outputs(2744) <= not(inputs(84)) or (inputs(249));
    layer0_outputs(2745) <= inputs(156);
    layer0_outputs(2746) <= (inputs(146)) and not (inputs(223));
    layer0_outputs(2747) <= (inputs(239)) xor (inputs(24));
    layer0_outputs(2748) <= not(inputs(203));
    layer0_outputs(2749) <= not(inputs(105)) or (inputs(27));
    layer0_outputs(2750) <= (inputs(228)) and not (inputs(254));
    layer0_outputs(2751) <= (inputs(54)) and not (inputs(5));
    layer0_outputs(2752) <= not(inputs(112)) or (inputs(140));
    layer0_outputs(2753) <= (inputs(205)) xor (inputs(228));
    layer0_outputs(2754) <= not(inputs(167));
    layer0_outputs(2755) <= not(inputs(106));
    layer0_outputs(2756) <= (inputs(216)) xor (inputs(233));
    layer0_outputs(2757) <= (inputs(169)) and not (inputs(3));
    layer0_outputs(2758) <= not(inputs(115));
    layer0_outputs(2759) <= (inputs(22)) or (inputs(223));
    layer0_outputs(2760) <= not(inputs(129));
    layer0_outputs(2761) <= (inputs(128)) xor (inputs(203));
    layer0_outputs(2762) <= not(inputs(57)) or (inputs(253));
    layer0_outputs(2763) <= not(inputs(119));
    layer0_outputs(2764) <= inputs(9);
    layer0_outputs(2765) <= (inputs(152)) xor (inputs(241));
    layer0_outputs(2766) <= inputs(124);
    layer0_outputs(2767) <= not((inputs(209)) or (inputs(55)));
    layer0_outputs(2768) <= (inputs(77)) or (inputs(62));
    layer0_outputs(2769) <= (inputs(216)) xor (inputs(28));
    layer0_outputs(2770) <= inputs(235);
    layer0_outputs(2771) <= not((inputs(164)) or (inputs(252)));
    layer0_outputs(2772) <= not(inputs(75));
    layer0_outputs(2773) <= not(inputs(200)) or (inputs(144));
    layer0_outputs(2774) <= (inputs(247)) or (inputs(81));
    layer0_outputs(2775) <= (inputs(100)) or (inputs(98));
    layer0_outputs(2776) <= (inputs(73)) or (inputs(70));
    layer0_outputs(2777) <= inputs(3);
    layer0_outputs(2778) <= (inputs(218)) or (inputs(216));
    layer0_outputs(2779) <= not(inputs(24));
    layer0_outputs(2780) <= not((inputs(0)) or (inputs(3)));
    layer0_outputs(2781) <= not((inputs(86)) or (inputs(82)));
    layer0_outputs(2782) <= (inputs(211)) or (inputs(224));
    layer0_outputs(2783) <= not((inputs(112)) or (inputs(145)));
    layer0_outputs(2784) <= not(inputs(191));
    layer0_outputs(2785) <= (inputs(81)) or (inputs(70));
    layer0_outputs(2786) <= inputs(37);
    layer0_outputs(2787) <= not(inputs(115));
    layer0_outputs(2788) <= (inputs(46)) and not (inputs(156));
    layer0_outputs(2789) <= not((inputs(117)) xor (inputs(124)));
    layer0_outputs(2790) <= not(inputs(110)) or (inputs(64));
    layer0_outputs(2791) <= not((inputs(58)) or (inputs(143)));
    layer0_outputs(2792) <= inputs(217);
    layer0_outputs(2793) <= (inputs(159)) xor (inputs(147));
    layer0_outputs(2794) <= inputs(92);
    layer0_outputs(2795) <= not(inputs(250)) or (inputs(31));
    layer0_outputs(2796) <= not(inputs(80));
    layer0_outputs(2797) <= (inputs(133)) and not (inputs(225));
    layer0_outputs(2798) <= not(inputs(216)) or (inputs(207));
    layer0_outputs(2799) <= (inputs(81)) xor (inputs(50));
    layer0_outputs(2800) <= not(inputs(52)) or (inputs(180));
    layer0_outputs(2801) <= not(inputs(187));
    layer0_outputs(2802) <= (inputs(86)) xor (inputs(36));
    layer0_outputs(2803) <= not(inputs(108)) or (inputs(255));
    layer0_outputs(2804) <= not(inputs(204)) or (inputs(242));
    layer0_outputs(2805) <= inputs(123);
    layer0_outputs(2806) <= inputs(222);
    layer0_outputs(2807) <= not(inputs(138)) or (inputs(47));
    layer0_outputs(2808) <= not(inputs(248));
    layer0_outputs(2809) <= (inputs(198)) xor (inputs(109));
    layer0_outputs(2810) <= inputs(120);
    layer0_outputs(2811) <= inputs(85);
    layer0_outputs(2812) <= (inputs(68)) or (inputs(20));
    layer0_outputs(2813) <= (inputs(143)) and not (inputs(168));
    layer0_outputs(2814) <= not((inputs(127)) xor (inputs(124)));
    layer0_outputs(2815) <= (inputs(228)) xor (inputs(35));
    layer0_outputs(2816) <= not(inputs(20));
    layer0_outputs(2817) <= not(inputs(224)) or (inputs(121));
    layer0_outputs(2818) <= (inputs(10)) and not (inputs(254));
    layer0_outputs(2819) <= not(inputs(150)) or (inputs(70));
    layer0_outputs(2820) <= not(inputs(99));
    layer0_outputs(2821) <= not(inputs(107));
    layer0_outputs(2822) <= (inputs(228)) or (inputs(98));
    layer0_outputs(2823) <= not((inputs(64)) or (inputs(37)));
    layer0_outputs(2824) <= (inputs(88)) xor (inputs(28));
    layer0_outputs(2825) <= not(inputs(130));
    layer0_outputs(2826) <= not((inputs(193)) xor (inputs(22)));
    layer0_outputs(2827) <= inputs(26);
    layer0_outputs(2828) <= not((inputs(18)) or (inputs(33)));
    layer0_outputs(2829) <= (inputs(238)) and not (inputs(231));
    layer0_outputs(2830) <= (inputs(147)) and not (inputs(18));
    layer0_outputs(2831) <= not(inputs(36)) or (inputs(2));
    layer0_outputs(2832) <= (inputs(104)) and not (inputs(232));
    layer0_outputs(2833) <= not((inputs(146)) or (inputs(153)));
    layer0_outputs(2834) <= inputs(168);
    layer0_outputs(2835) <= (inputs(120)) and (inputs(40));
    layer0_outputs(2836) <= not((inputs(111)) or (inputs(74)));
    layer0_outputs(2837) <= not((inputs(238)) or (inputs(136)));
    layer0_outputs(2838) <= inputs(30);
    layer0_outputs(2839) <= (inputs(216)) or (inputs(19));
    layer0_outputs(2840) <= not(inputs(97)) or (inputs(207));
    layer0_outputs(2841) <= not((inputs(117)) or (inputs(229)));
    layer0_outputs(2842) <= (inputs(67)) xor (inputs(220));
    layer0_outputs(2843) <= (inputs(30)) or (inputs(69));
    layer0_outputs(2844) <= not((inputs(192)) xor (inputs(19)));
    layer0_outputs(2845) <= inputs(191);
    layer0_outputs(2846) <= not((inputs(254)) or (inputs(186)));
    layer0_outputs(2847) <= not(inputs(19));
    layer0_outputs(2848) <= (inputs(125)) or (inputs(138));
    layer0_outputs(2849) <= (inputs(56)) or (inputs(17));
    layer0_outputs(2850) <= (inputs(252)) or (inputs(93));
    layer0_outputs(2851) <= inputs(91);
    layer0_outputs(2852) <= not(inputs(18));
    layer0_outputs(2853) <= '1';
    layer0_outputs(2854) <= not((inputs(194)) and (inputs(214)));
    layer0_outputs(2855) <= not(inputs(25));
    layer0_outputs(2856) <= (inputs(3)) xor (inputs(33));
    layer0_outputs(2857) <= inputs(89);
    layer0_outputs(2858) <= not(inputs(150)) or (inputs(28));
    layer0_outputs(2859) <= not(inputs(91));
    layer0_outputs(2860) <= not((inputs(238)) xor (inputs(24)));
    layer0_outputs(2861) <= inputs(182);
    layer0_outputs(2862) <= (inputs(64)) xor (inputs(206));
    layer0_outputs(2863) <= not((inputs(251)) xor (inputs(204)));
    layer0_outputs(2864) <= not(inputs(129));
    layer0_outputs(2865) <= not((inputs(24)) and (inputs(118)));
    layer0_outputs(2866) <= not((inputs(170)) xor (inputs(218)));
    layer0_outputs(2867) <= inputs(108);
    layer0_outputs(2868) <= (inputs(233)) and not (inputs(49));
    layer0_outputs(2869) <= (inputs(247)) and not (inputs(241));
    layer0_outputs(2870) <= not(inputs(3));
    layer0_outputs(2871) <= (inputs(2)) or (inputs(236));
    layer0_outputs(2872) <= not((inputs(63)) or (inputs(35)));
    layer0_outputs(2873) <= inputs(239);
    layer0_outputs(2874) <= not((inputs(39)) or (inputs(74)));
    layer0_outputs(2875) <= inputs(148);
    layer0_outputs(2876) <= not(inputs(251));
    layer0_outputs(2877) <= not(inputs(23));
    layer0_outputs(2878) <= not((inputs(151)) or (inputs(7)));
    layer0_outputs(2879) <= not((inputs(135)) or (inputs(44)));
    layer0_outputs(2880) <= (inputs(196)) or (inputs(195));
    layer0_outputs(2881) <= not(inputs(246)) or (inputs(228));
    layer0_outputs(2882) <= not((inputs(99)) or (inputs(157)));
    layer0_outputs(2883) <= (inputs(53)) and (inputs(56));
    layer0_outputs(2884) <= not(inputs(89));
    layer0_outputs(2885) <= not(inputs(237));
    layer0_outputs(2886) <= not((inputs(194)) xor (inputs(197)));
    layer0_outputs(2887) <= (inputs(39)) or (inputs(239));
    layer0_outputs(2888) <= (inputs(154)) xor (inputs(167));
    layer0_outputs(2889) <= not((inputs(229)) or (inputs(100)));
    layer0_outputs(2890) <= (inputs(13)) xor (inputs(23));
    layer0_outputs(2891) <= not((inputs(116)) xor (inputs(36)));
    layer0_outputs(2892) <= not((inputs(244)) xor (inputs(221)));
    layer0_outputs(2893) <= inputs(45);
    layer0_outputs(2894) <= (inputs(254)) or (inputs(178));
    layer0_outputs(2895) <= (inputs(166)) and not (inputs(191));
    layer0_outputs(2896) <= '0';
    layer0_outputs(2897) <= not((inputs(53)) xor (inputs(87)));
    layer0_outputs(2898) <= inputs(82);
    layer0_outputs(2899) <= not(inputs(11));
    layer0_outputs(2900) <= not(inputs(90));
    layer0_outputs(2901) <= inputs(210);
    layer0_outputs(2902) <= not(inputs(197)) or (inputs(248));
    layer0_outputs(2903) <= not(inputs(117));
    layer0_outputs(2904) <= not((inputs(200)) xor (inputs(109)));
    layer0_outputs(2905) <= (inputs(20)) xor (inputs(65));
    layer0_outputs(2906) <= not(inputs(111)) or (inputs(110));
    layer0_outputs(2907) <= (inputs(60)) xor (inputs(9));
    layer0_outputs(2908) <= (inputs(46)) and (inputs(239));
    layer0_outputs(2909) <= (inputs(199)) or (inputs(133));
    layer0_outputs(2910) <= not(inputs(107));
    layer0_outputs(2911) <= (inputs(45)) or (inputs(104));
    layer0_outputs(2912) <= not((inputs(157)) xor (inputs(108)));
    layer0_outputs(2913) <= (inputs(76)) or (inputs(122));
    layer0_outputs(2914) <= (inputs(211)) and not (inputs(33));
    layer0_outputs(2915) <= not((inputs(31)) or (inputs(37)));
    layer0_outputs(2916) <= not(inputs(109));
    layer0_outputs(2917) <= inputs(84);
    layer0_outputs(2918) <= not(inputs(167));
    layer0_outputs(2919) <= (inputs(142)) or (inputs(139));
    layer0_outputs(2920) <= (inputs(26)) or (inputs(194));
    layer0_outputs(2921) <= inputs(167);
    layer0_outputs(2922) <= inputs(84);
    layer0_outputs(2923) <= not(inputs(214)) or (inputs(225));
    layer0_outputs(2924) <= '1';
    layer0_outputs(2925) <= not(inputs(116));
    layer0_outputs(2926) <= not((inputs(41)) or (inputs(254)));
    layer0_outputs(2927) <= not(inputs(142));
    layer0_outputs(2928) <= not(inputs(190)) or (inputs(82));
    layer0_outputs(2929) <= (inputs(73)) xor (inputs(7));
    layer0_outputs(2930) <= not(inputs(201)) or (inputs(212));
    layer0_outputs(2931) <= (inputs(251)) or (inputs(198));
    layer0_outputs(2932) <= (inputs(107)) or (inputs(53));
    layer0_outputs(2933) <= '0';
    layer0_outputs(2934) <= not((inputs(3)) or (inputs(124)));
    layer0_outputs(2935) <= (inputs(57)) and not (inputs(251));
    layer0_outputs(2936) <= inputs(136);
    layer0_outputs(2937) <= (inputs(69)) and not (inputs(55));
    layer0_outputs(2938) <= (inputs(16)) or (inputs(234));
    layer0_outputs(2939) <= (inputs(54)) or (inputs(114));
    layer0_outputs(2940) <= not(inputs(4));
    layer0_outputs(2941) <= inputs(112);
    layer0_outputs(2942) <= inputs(95);
    layer0_outputs(2943) <= not(inputs(87));
    layer0_outputs(2944) <= inputs(25);
    layer0_outputs(2945) <= (inputs(6)) and not (inputs(144));
    layer0_outputs(2946) <= (inputs(86)) or (inputs(255));
    layer0_outputs(2947) <= not(inputs(219)) or (inputs(82));
    layer0_outputs(2948) <= inputs(231);
    layer0_outputs(2949) <= not(inputs(142)) or (inputs(184));
    layer0_outputs(2950) <= (inputs(216)) or (inputs(188));
    layer0_outputs(2951) <= not((inputs(130)) or (inputs(60)));
    layer0_outputs(2952) <= not(inputs(217));
    layer0_outputs(2953) <= inputs(138);
    layer0_outputs(2954) <= inputs(67);
    layer0_outputs(2955) <= not(inputs(70));
    layer0_outputs(2956) <= inputs(209);
    layer0_outputs(2957) <= not((inputs(220)) or (inputs(34)));
    layer0_outputs(2958) <= not(inputs(56));
    layer0_outputs(2959) <= not(inputs(182));
    layer0_outputs(2960) <= not((inputs(48)) or (inputs(225)));
    layer0_outputs(2961) <= '0';
    layer0_outputs(2962) <= (inputs(190)) xor (inputs(138));
    layer0_outputs(2963) <= not(inputs(116));
    layer0_outputs(2964) <= not(inputs(103)) or (inputs(97));
    layer0_outputs(2965) <= not((inputs(55)) xor (inputs(74)));
    layer0_outputs(2966) <= not(inputs(180));
    layer0_outputs(2967) <= not(inputs(194)) or (inputs(112));
    layer0_outputs(2968) <= not((inputs(61)) xor (inputs(115)));
    layer0_outputs(2969) <= inputs(22);
    layer0_outputs(2970) <= (inputs(112)) or (inputs(78));
    layer0_outputs(2971) <= (inputs(212)) xor (inputs(148));
    layer0_outputs(2972) <= (inputs(188)) or (inputs(147));
    layer0_outputs(2973) <= not((inputs(140)) xor (inputs(225)));
    layer0_outputs(2974) <= not(inputs(162));
    layer0_outputs(2975) <= (inputs(201)) and (inputs(171));
    layer0_outputs(2976) <= (inputs(166)) and not (inputs(12));
    layer0_outputs(2977) <= (inputs(232)) xor (inputs(79));
    layer0_outputs(2978) <= not(inputs(42)) or (inputs(181));
    layer0_outputs(2979) <= not(inputs(47)) or (inputs(66));
    layer0_outputs(2980) <= (inputs(125)) and not (inputs(224));
    layer0_outputs(2981) <= (inputs(7)) and not (inputs(189));
    layer0_outputs(2982) <= (inputs(161)) or (inputs(150));
    layer0_outputs(2983) <= not((inputs(99)) or (inputs(128)));
    layer0_outputs(2984) <= (inputs(248)) xor (inputs(146));
    layer0_outputs(2985) <= inputs(161);
    layer0_outputs(2986) <= inputs(106);
    layer0_outputs(2987) <= not(inputs(162));
    layer0_outputs(2988) <= inputs(251);
    layer0_outputs(2989) <= not(inputs(156)) or (inputs(33));
    layer0_outputs(2990) <= not((inputs(180)) or (inputs(97)));
    layer0_outputs(2991) <= not(inputs(165));
    layer0_outputs(2992) <= inputs(193);
    layer0_outputs(2993) <= (inputs(235)) xor (inputs(79));
    layer0_outputs(2994) <= (inputs(86)) xor (inputs(49));
    layer0_outputs(2995) <= (inputs(68)) or (inputs(200));
    layer0_outputs(2996) <= not((inputs(229)) xor (inputs(165)));
    layer0_outputs(2997) <= (inputs(5)) xor (inputs(142));
    layer0_outputs(2998) <= not(inputs(71));
    layer0_outputs(2999) <= (inputs(43)) or (inputs(112));
    layer0_outputs(3000) <= (inputs(32)) or (inputs(49));
    layer0_outputs(3001) <= not(inputs(201));
    layer0_outputs(3002) <= not((inputs(124)) and (inputs(174)));
    layer0_outputs(3003) <= (inputs(104)) xor (inputs(130));
    layer0_outputs(3004) <= not((inputs(217)) xor (inputs(202)));
    layer0_outputs(3005) <= (inputs(44)) and (inputs(219));
    layer0_outputs(3006) <= not((inputs(147)) xor (inputs(119)));
    layer0_outputs(3007) <= not(inputs(106)) or (inputs(15));
    layer0_outputs(3008) <= not((inputs(178)) or (inputs(67)));
    layer0_outputs(3009) <= inputs(128);
    layer0_outputs(3010) <= inputs(96);
    layer0_outputs(3011) <= not((inputs(59)) or (inputs(110)));
    layer0_outputs(3012) <= not(inputs(44)) or (inputs(118));
    layer0_outputs(3013) <= not(inputs(247));
    layer0_outputs(3014) <= (inputs(90)) and not (inputs(128));
    layer0_outputs(3015) <= (inputs(212)) and not (inputs(2));
    layer0_outputs(3016) <= not((inputs(89)) or (inputs(86)));
    layer0_outputs(3017) <= (inputs(53)) xor (inputs(8));
    layer0_outputs(3018) <= not((inputs(114)) xor (inputs(69)));
    layer0_outputs(3019) <= not((inputs(133)) or (inputs(148)));
    layer0_outputs(3020) <= not(inputs(75));
    layer0_outputs(3021) <= inputs(67);
    layer0_outputs(3022) <= inputs(60);
    layer0_outputs(3023) <= not(inputs(202)) or (inputs(9));
    layer0_outputs(3024) <= (inputs(5)) and not (inputs(87));
    layer0_outputs(3025) <= inputs(207);
    layer0_outputs(3026) <= inputs(179);
    layer0_outputs(3027) <= inputs(73);
    layer0_outputs(3028) <= (inputs(79)) xor (inputs(79));
    layer0_outputs(3029) <= not((inputs(31)) or (inputs(97)));
    layer0_outputs(3030) <= not((inputs(116)) or (inputs(85)));
    layer0_outputs(3031) <= (inputs(201)) and not (inputs(27));
    layer0_outputs(3032) <= inputs(244);
    layer0_outputs(3033) <= (inputs(106)) and not (inputs(222));
    layer0_outputs(3034) <= (inputs(51)) or (inputs(188));
    layer0_outputs(3035) <= not((inputs(212)) xor (inputs(219)));
    layer0_outputs(3036) <= inputs(82);
    layer0_outputs(3037) <= not((inputs(185)) xor (inputs(12)));
    layer0_outputs(3038) <= '0';
    layer0_outputs(3039) <= not((inputs(159)) or (inputs(109)));
    layer0_outputs(3040) <= inputs(168);
    layer0_outputs(3041) <= not((inputs(238)) or (inputs(77)));
    layer0_outputs(3042) <= '0';
    layer0_outputs(3043) <= inputs(151);
    layer0_outputs(3044) <= not(inputs(220)) or (inputs(40));
    layer0_outputs(3045) <= not((inputs(141)) or (inputs(234)));
    layer0_outputs(3046) <= not(inputs(154)) or (inputs(226));
    layer0_outputs(3047) <= not(inputs(206));
    layer0_outputs(3048) <= (inputs(100)) and (inputs(124));
    layer0_outputs(3049) <= not(inputs(74));
    layer0_outputs(3050) <= not(inputs(30)) or (inputs(177));
    layer0_outputs(3051) <= not(inputs(141)) or (inputs(221));
    layer0_outputs(3052) <= inputs(44);
    layer0_outputs(3053) <= not((inputs(88)) or (inputs(85)));
    layer0_outputs(3054) <= not(inputs(112));
    layer0_outputs(3055) <= not(inputs(97)) or (inputs(239));
    layer0_outputs(3056) <= inputs(197);
    layer0_outputs(3057) <= not(inputs(181));
    layer0_outputs(3058) <= not((inputs(130)) or (inputs(4)));
    layer0_outputs(3059) <= not(inputs(203));
    layer0_outputs(3060) <= (inputs(198)) and not (inputs(47));
    layer0_outputs(3061) <= inputs(179);
    layer0_outputs(3062) <= not((inputs(198)) xor (inputs(133)));
    layer0_outputs(3063) <= not((inputs(61)) xor (inputs(202)));
    layer0_outputs(3064) <= not((inputs(196)) or (inputs(194)));
    layer0_outputs(3065) <= not((inputs(128)) xor (inputs(116)));
    layer0_outputs(3066) <= not((inputs(65)) or (inputs(105)));
    layer0_outputs(3067) <= not(inputs(177));
    layer0_outputs(3068) <= not(inputs(124)) or (inputs(122));
    layer0_outputs(3069) <= not(inputs(142));
    layer0_outputs(3070) <= not(inputs(142));
    layer0_outputs(3071) <= not(inputs(48)) or (inputs(213));
    layer0_outputs(3072) <= not(inputs(37)) or (inputs(243));
    layer0_outputs(3073) <= (inputs(193)) and not (inputs(201));
    layer0_outputs(3074) <= inputs(229);
    layer0_outputs(3075) <= not((inputs(221)) or (inputs(88)));
    layer0_outputs(3076) <= (inputs(9)) or (inputs(174));
    layer0_outputs(3077) <= not(inputs(117));
    layer0_outputs(3078) <= (inputs(86)) xor (inputs(130));
    layer0_outputs(3079) <= not((inputs(55)) xor (inputs(74)));
    layer0_outputs(3080) <= not(inputs(62));
    layer0_outputs(3081) <= not((inputs(102)) or (inputs(161)));
    layer0_outputs(3082) <= not(inputs(55)) or (inputs(146));
    layer0_outputs(3083) <= inputs(241);
    layer0_outputs(3084) <= (inputs(235)) and not (inputs(61));
    layer0_outputs(3085) <= inputs(117);
    layer0_outputs(3086) <= (inputs(107)) or (inputs(176));
    layer0_outputs(3087) <= '1';
    layer0_outputs(3088) <= not(inputs(101));
    layer0_outputs(3089) <= (inputs(153)) or (inputs(208));
    layer0_outputs(3090) <= (inputs(211)) or (inputs(73));
    layer0_outputs(3091) <= not((inputs(156)) xor (inputs(194)));
    layer0_outputs(3092) <= not(inputs(61));
    layer0_outputs(3093) <= not(inputs(162));
    layer0_outputs(3094) <= inputs(239);
    layer0_outputs(3095) <= (inputs(230)) and not (inputs(18));
    layer0_outputs(3096) <= not(inputs(74)) or (inputs(52));
    layer0_outputs(3097) <= (inputs(122)) and not (inputs(176));
    layer0_outputs(3098) <= '0';
    layer0_outputs(3099) <= inputs(72);
    layer0_outputs(3100) <= (inputs(122)) and not (inputs(250));
    layer0_outputs(3101) <= not(inputs(119)) or (inputs(112));
    layer0_outputs(3102) <= inputs(122);
    layer0_outputs(3103) <= not(inputs(80)) or (inputs(68));
    layer0_outputs(3104) <= inputs(106);
    layer0_outputs(3105) <= (inputs(50)) and not (inputs(169));
    layer0_outputs(3106) <= not((inputs(179)) and (inputs(148)));
    layer0_outputs(3107) <= (inputs(106)) xor (inputs(139));
    layer0_outputs(3108) <= not(inputs(188)) or (inputs(14));
    layer0_outputs(3109) <= not((inputs(1)) xor (inputs(49)));
    layer0_outputs(3110) <= (inputs(230)) and not (inputs(109));
    layer0_outputs(3111) <= inputs(101);
    layer0_outputs(3112) <= inputs(45);
    layer0_outputs(3113) <= inputs(41);
    layer0_outputs(3114) <= inputs(110);
    layer0_outputs(3115) <= inputs(92);
    layer0_outputs(3116) <= inputs(247);
    layer0_outputs(3117) <= not((inputs(255)) xor (inputs(25)));
    layer0_outputs(3118) <= inputs(51);
    layer0_outputs(3119) <= inputs(107);
    layer0_outputs(3120) <= not(inputs(197));
    layer0_outputs(3121) <= not(inputs(118)) or (inputs(129));
    layer0_outputs(3122) <= not(inputs(73)) or (inputs(169));
    layer0_outputs(3123) <= not((inputs(131)) or (inputs(202)));
    layer0_outputs(3124) <= (inputs(1)) and not (inputs(30));
    layer0_outputs(3125) <= (inputs(248)) or (inputs(117));
    layer0_outputs(3126) <= (inputs(59)) xor (inputs(71));
    layer0_outputs(3127) <= not(inputs(64)) or (inputs(127));
    layer0_outputs(3128) <= (inputs(101)) and not (inputs(16));
    layer0_outputs(3129) <= inputs(193);
    layer0_outputs(3130) <= not((inputs(33)) xor (inputs(86)));
    layer0_outputs(3131) <= not(inputs(73));
    layer0_outputs(3132) <= not(inputs(233));
    layer0_outputs(3133) <= (inputs(122)) and not (inputs(234));
    layer0_outputs(3134) <= not((inputs(12)) xor (inputs(155)));
    layer0_outputs(3135) <= not((inputs(44)) or (inputs(23)));
    layer0_outputs(3136) <= not((inputs(9)) or (inputs(144)));
    layer0_outputs(3137) <= inputs(86);
    layer0_outputs(3138) <= not(inputs(95));
    layer0_outputs(3139) <= not(inputs(176)) or (inputs(255));
    layer0_outputs(3140) <= '1';
    layer0_outputs(3141) <= not((inputs(1)) or (inputs(59)));
    layer0_outputs(3142) <= not((inputs(217)) xor (inputs(65)));
    layer0_outputs(3143) <= not((inputs(40)) xor (inputs(91)));
    layer0_outputs(3144) <= inputs(180);
    layer0_outputs(3145) <= inputs(76);
    layer0_outputs(3146) <= not((inputs(161)) xor (inputs(143)));
    layer0_outputs(3147) <= not(inputs(35));
    layer0_outputs(3148) <= (inputs(134)) and not (inputs(255));
    layer0_outputs(3149) <= (inputs(252)) or (inputs(48));
    layer0_outputs(3150) <= inputs(86);
    layer0_outputs(3151) <= not(inputs(129)) or (inputs(224));
    layer0_outputs(3152) <= (inputs(46)) xor (inputs(34));
    layer0_outputs(3153) <= not(inputs(97));
    layer0_outputs(3154) <= (inputs(221)) xor (inputs(167));
    layer0_outputs(3155) <= not(inputs(114));
    layer0_outputs(3156) <= not((inputs(219)) or (inputs(194)));
    layer0_outputs(3157) <= inputs(255);
    layer0_outputs(3158) <= not(inputs(249)) or (inputs(73));
    layer0_outputs(3159) <= (inputs(49)) or (inputs(108));
    layer0_outputs(3160) <= (inputs(125)) and not (inputs(177));
    layer0_outputs(3161) <= (inputs(20)) or (inputs(1));
    layer0_outputs(3162) <= (inputs(223)) xor (inputs(148));
    layer0_outputs(3163) <= (inputs(119)) and not (inputs(58));
    layer0_outputs(3164) <= not(inputs(163));
    layer0_outputs(3165) <= (inputs(171)) and not (inputs(210));
    layer0_outputs(3166) <= (inputs(45)) or (inputs(231));
    layer0_outputs(3167) <= (inputs(205)) and not (inputs(78));
    layer0_outputs(3168) <= not((inputs(218)) or (inputs(236)));
    layer0_outputs(3169) <= not(inputs(56)) or (inputs(125));
    layer0_outputs(3170) <= (inputs(163)) xor (inputs(211));
    layer0_outputs(3171) <= not(inputs(46)) or (inputs(237));
    layer0_outputs(3172) <= not((inputs(154)) or (inputs(251)));
    layer0_outputs(3173) <= (inputs(72)) and not (inputs(227));
    layer0_outputs(3174) <= (inputs(73)) and not (inputs(177));
    layer0_outputs(3175) <= '1';
    layer0_outputs(3176) <= not((inputs(111)) xor (inputs(30)));
    layer0_outputs(3177) <= not(inputs(229));
    layer0_outputs(3178) <= not((inputs(188)) and (inputs(188)));
    layer0_outputs(3179) <= (inputs(36)) xor (inputs(52));
    layer0_outputs(3180) <= not(inputs(198)) or (inputs(93));
    layer0_outputs(3181) <= (inputs(52)) or (inputs(111));
    layer0_outputs(3182) <= (inputs(88)) or (inputs(135));
    layer0_outputs(3183) <= not(inputs(224)) or (inputs(250));
    layer0_outputs(3184) <= not(inputs(109)) or (inputs(236));
    layer0_outputs(3185) <= not(inputs(116)) or (inputs(19));
    layer0_outputs(3186) <= not((inputs(69)) xor (inputs(37)));
    layer0_outputs(3187) <= not((inputs(125)) xor (inputs(45)));
    layer0_outputs(3188) <= not(inputs(152));
    layer0_outputs(3189) <= not(inputs(41));
    layer0_outputs(3190) <= inputs(164);
    layer0_outputs(3191) <= inputs(216);
    layer0_outputs(3192) <= not(inputs(95));
    layer0_outputs(3193) <= (inputs(43)) and not (inputs(250));
    layer0_outputs(3194) <= (inputs(186)) and (inputs(23));
    layer0_outputs(3195) <= not(inputs(233)) or (inputs(211));
    layer0_outputs(3196) <= not(inputs(178));
    layer0_outputs(3197) <= inputs(246);
    layer0_outputs(3198) <= (inputs(163)) and not (inputs(1));
    layer0_outputs(3199) <= (inputs(0)) or (inputs(165));
    layer0_outputs(3200) <= (inputs(84)) or (inputs(7));
    layer0_outputs(3201) <= not(inputs(226));
    layer0_outputs(3202) <= (inputs(88)) xor (inputs(218));
    layer0_outputs(3203) <= (inputs(213)) and not (inputs(23));
    layer0_outputs(3204) <= not(inputs(40)) or (inputs(234));
    layer0_outputs(3205) <= (inputs(83)) or (inputs(5));
    layer0_outputs(3206) <= (inputs(255)) and (inputs(3));
    layer0_outputs(3207) <= (inputs(88)) xor (inputs(136));
    layer0_outputs(3208) <= (inputs(13)) or (inputs(208));
    layer0_outputs(3209) <= (inputs(111)) and not (inputs(36));
    layer0_outputs(3210) <= not(inputs(88)) or (inputs(211));
    layer0_outputs(3211) <= (inputs(214)) or (inputs(196));
    layer0_outputs(3212) <= not((inputs(161)) and (inputs(26)));
    layer0_outputs(3213) <= not(inputs(97));
    layer0_outputs(3214) <= not((inputs(9)) or (inputs(191)));
    layer0_outputs(3215) <= (inputs(20)) or (inputs(31));
    layer0_outputs(3216) <= inputs(124);
    layer0_outputs(3217) <= (inputs(105)) and not (inputs(165));
    layer0_outputs(3218) <= inputs(41);
    layer0_outputs(3219) <= (inputs(147)) and not (inputs(210));
    layer0_outputs(3220) <= (inputs(58)) or (inputs(237));
    layer0_outputs(3221) <= inputs(23);
    layer0_outputs(3222) <= inputs(189);
    layer0_outputs(3223) <= (inputs(7)) and (inputs(125));
    layer0_outputs(3224) <= not(inputs(92));
    layer0_outputs(3225) <= inputs(190);
    layer0_outputs(3226) <= not((inputs(110)) or (inputs(147)));
    layer0_outputs(3227) <= (inputs(95)) and not (inputs(110));
    layer0_outputs(3228) <= (inputs(125)) xor (inputs(165));
    layer0_outputs(3229) <= not(inputs(215));
    layer0_outputs(3230) <= inputs(37);
    layer0_outputs(3231) <= not(inputs(46));
    layer0_outputs(3232) <= not(inputs(21));
    layer0_outputs(3233) <= not(inputs(205));
    layer0_outputs(3234) <= not((inputs(248)) or (inputs(52)));
    layer0_outputs(3235) <= not(inputs(82)) or (inputs(144));
    layer0_outputs(3236) <= (inputs(44)) or (inputs(37));
    layer0_outputs(3237) <= inputs(68);
    layer0_outputs(3238) <= (inputs(86)) or (inputs(130));
    layer0_outputs(3239) <= not((inputs(242)) xor (inputs(59)));
    layer0_outputs(3240) <= '0';
    layer0_outputs(3241) <= (inputs(64)) and (inputs(250));
    layer0_outputs(3242) <= not(inputs(141)) or (inputs(114));
    layer0_outputs(3243) <= not(inputs(54));
    layer0_outputs(3244) <= (inputs(39)) or (inputs(125));
    layer0_outputs(3245) <= not(inputs(31));
    layer0_outputs(3246) <= (inputs(231)) and not (inputs(149));
    layer0_outputs(3247) <= not(inputs(227));
    layer0_outputs(3248) <= (inputs(29)) and not (inputs(80));
    layer0_outputs(3249) <= not(inputs(54));
    layer0_outputs(3250) <= not(inputs(152)) or (inputs(87));
    layer0_outputs(3251) <= not((inputs(88)) xor (inputs(225)));
    layer0_outputs(3252) <= not((inputs(58)) or (inputs(66)));
    layer0_outputs(3253) <= not(inputs(163));
    layer0_outputs(3254) <= (inputs(127)) and not (inputs(208));
    layer0_outputs(3255) <= not((inputs(181)) xor (inputs(140)));
    layer0_outputs(3256) <= (inputs(29)) and not (inputs(107));
    layer0_outputs(3257) <= (inputs(15)) or (inputs(238));
    layer0_outputs(3258) <= not((inputs(62)) or (inputs(0)));
    layer0_outputs(3259) <= (inputs(18)) or (inputs(154));
    layer0_outputs(3260) <= not(inputs(113));
    layer0_outputs(3261) <= not((inputs(128)) or (inputs(120)));
    layer0_outputs(3262) <= inputs(182);
    layer0_outputs(3263) <= inputs(76);
    layer0_outputs(3264) <= not((inputs(223)) and (inputs(186)));
    layer0_outputs(3265) <= not(inputs(173)) or (inputs(85));
    layer0_outputs(3266) <= (inputs(15)) or (inputs(200));
    layer0_outputs(3267) <= not((inputs(36)) or (inputs(160)));
    layer0_outputs(3268) <= (inputs(131)) and not (inputs(192));
    layer0_outputs(3269) <= not((inputs(159)) xor (inputs(36)));
    layer0_outputs(3270) <= inputs(41);
    layer0_outputs(3271) <= inputs(111);
    layer0_outputs(3272) <= inputs(29);
    layer0_outputs(3273) <= not(inputs(181));
    layer0_outputs(3274) <= not(inputs(118)) or (inputs(36));
    layer0_outputs(3275) <= not((inputs(215)) or (inputs(49)));
    layer0_outputs(3276) <= '0';
    layer0_outputs(3277) <= not(inputs(159));
    layer0_outputs(3278) <= (inputs(150)) or (inputs(84));
    layer0_outputs(3279) <= not(inputs(142));
    layer0_outputs(3280) <= (inputs(144)) and not (inputs(18));
    layer0_outputs(3281) <= not(inputs(224));
    layer0_outputs(3282) <= not(inputs(12));
    layer0_outputs(3283) <= not((inputs(147)) and (inputs(80)));
    layer0_outputs(3284) <= (inputs(59)) and (inputs(53));
    layer0_outputs(3285) <= inputs(118);
    layer0_outputs(3286) <= not((inputs(35)) xor (inputs(131)));
    layer0_outputs(3287) <= inputs(227);
    layer0_outputs(3288) <= not(inputs(115));
    layer0_outputs(3289) <= (inputs(247)) or (inputs(132));
    layer0_outputs(3290) <= not((inputs(108)) or (inputs(53)));
    layer0_outputs(3291) <= inputs(13);
    layer0_outputs(3292) <= inputs(84);
    layer0_outputs(3293) <= not(inputs(24)) or (inputs(233));
    layer0_outputs(3294) <= not((inputs(171)) xor (inputs(245)));
    layer0_outputs(3295) <= not(inputs(182));
    layer0_outputs(3296) <= not(inputs(10)) or (inputs(182));
    layer0_outputs(3297) <= not((inputs(74)) or (inputs(159)));
    layer0_outputs(3298) <= (inputs(117)) and not (inputs(227));
    layer0_outputs(3299) <= inputs(140);
    layer0_outputs(3300) <= (inputs(66)) or (inputs(207));
    layer0_outputs(3301) <= not((inputs(211)) or (inputs(65)));
    layer0_outputs(3302) <= not(inputs(231));
    layer0_outputs(3303) <= not((inputs(33)) or (inputs(219)));
    layer0_outputs(3304) <= (inputs(204)) xor (inputs(114));
    layer0_outputs(3305) <= inputs(54);
    layer0_outputs(3306) <= not(inputs(182));
    layer0_outputs(3307) <= not(inputs(163)) or (inputs(48));
    layer0_outputs(3308) <= (inputs(70)) or (inputs(237));
    layer0_outputs(3309) <= not(inputs(21));
    layer0_outputs(3310) <= (inputs(146)) xor (inputs(149));
    layer0_outputs(3311) <= not(inputs(107)) or (inputs(15));
    layer0_outputs(3312) <= (inputs(71)) or (inputs(158));
    layer0_outputs(3313) <= not(inputs(37)) or (inputs(113));
    layer0_outputs(3314) <= not(inputs(253)) or (inputs(174));
    layer0_outputs(3315) <= inputs(114);
    layer0_outputs(3316) <= inputs(160);
    layer0_outputs(3317) <= not(inputs(131));
    layer0_outputs(3318) <= inputs(161);
    layer0_outputs(3319) <= (inputs(140)) xor (inputs(103));
    layer0_outputs(3320) <= not(inputs(157));
    layer0_outputs(3321) <= (inputs(79)) or (inputs(80));
    layer0_outputs(3322) <= (inputs(24)) and (inputs(91));
    layer0_outputs(3323) <= not((inputs(110)) or (inputs(185)));
    layer0_outputs(3324) <= not((inputs(71)) or (inputs(84)));
    layer0_outputs(3325) <= not(inputs(154)) or (inputs(207));
    layer0_outputs(3326) <= (inputs(74)) or (inputs(26));
    layer0_outputs(3327) <= not(inputs(8)) or (inputs(201));
    layer0_outputs(3328) <= not(inputs(37)) or (inputs(58));
    layer0_outputs(3329) <= not(inputs(102)) or (inputs(56));
    layer0_outputs(3330) <= not(inputs(255));
    layer0_outputs(3331) <= not(inputs(2)) or (inputs(240));
    layer0_outputs(3332) <= not(inputs(114));
    layer0_outputs(3333) <= inputs(196);
    layer0_outputs(3334) <= inputs(178);
    layer0_outputs(3335) <= (inputs(36)) or (inputs(39));
    layer0_outputs(3336) <= not((inputs(183)) xor (inputs(192)));
    layer0_outputs(3337) <= inputs(91);
    layer0_outputs(3338) <= (inputs(199)) and not (inputs(136));
    layer0_outputs(3339) <= (inputs(93)) and not (inputs(222));
    layer0_outputs(3340) <= not(inputs(9));
    layer0_outputs(3341) <= '1';
    layer0_outputs(3342) <= not(inputs(236)) or (inputs(114));
    layer0_outputs(3343) <= (inputs(46)) and not (inputs(172));
    layer0_outputs(3344) <= inputs(219);
    layer0_outputs(3345) <= inputs(1);
    layer0_outputs(3346) <= not((inputs(33)) or (inputs(100)));
    layer0_outputs(3347) <= inputs(166);
    layer0_outputs(3348) <= (inputs(106)) and not (inputs(177));
    layer0_outputs(3349) <= (inputs(89)) xor (inputs(215));
    layer0_outputs(3350) <= not(inputs(67)) or (inputs(198));
    layer0_outputs(3351) <= (inputs(43)) and not (inputs(222));
    layer0_outputs(3352) <= (inputs(220)) and not (inputs(184));
    layer0_outputs(3353) <= inputs(156);
    layer0_outputs(3354) <= not(inputs(118)) or (inputs(241));
    layer0_outputs(3355) <= inputs(17);
    layer0_outputs(3356) <= not(inputs(98));
    layer0_outputs(3357) <= (inputs(225)) or (inputs(103));
    layer0_outputs(3358) <= not((inputs(56)) or (inputs(77)));
    layer0_outputs(3359) <= (inputs(139)) xor (inputs(96));
    layer0_outputs(3360) <= (inputs(101)) and not (inputs(161));
    layer0_outputs(3361) <= not(inputs(167));
    layer0_outputs(3362) <= not((inputs(4)) and (inputs(241)));
    layer0_outputs(3363) <= not(inputs(10));
    layer0_outputs(3364) <= (inputs(217)) and not (inputs(49));
    layer0_outputs(3365) <= (inputs(61)) and not (inputs(212));
    layer0_outputs(3366) <= inputs(137);
    layer0_outputs(3367) <= not(inputs(16));
    layer0_outputs(3368) <= inputs(137);
    layer0_outputs(3369) <= inputs(190);
    layer0_outputs(3370) <= not(inputs(215)) or (inputs(185));
    layer0_outputs(3371) <= inputs(107);
    layer0_outputs(3372) <= (inputs(242)) and not (inputs(75));
    layer0_outputs(3373) <= not(inputs(249)) or (inputs(126));
    layer0_outputs(3374) <= (inputs(105)) xor (inputs(80));
    layer0_outputs(3375) <= not(inputs(137));
    layer0_outputs(3376) <= (inputs(186)) or (inputs(50));
    layer0_outputs(3377) <= (inputs(193)) or (inputs(217));
    layer0_outputs(3378) <= (inputs(76)) xor (inputs(27));
    layer0_outputs(3379) <= inputs(169);
    layer0_outputs(3380) <= not(inputs(102));
    layer0_outputs(3381) <= inputs(88);
    layer0_outputs(3382) <= (inputs(246)) and not (inputs(30));
    layer0_outputs(3383) <= (inputs(12)) or (inputs(241));
    layer0_outputs(3384) <= not((inputs(95)) or (inputs(136)));
    layer0_outputs(3385) <= not((inputs(168)) xor (inputs(242)));
    layer0_outputs(3386) <= inputs(245);
    layer0_outputs(3387) <= not(inputs(56)) or (inputs(12));
    layer0_outputs(3388) <= inputs(151);
    layer0_outputs(3389) <= inputs(34);
    layer0_outputs(3390) <= '1';
    layer0_outputs(3391) <= (inputs(117)) or (inputs(138));
    layer0_outputs(3392) <= not((inputs(187)) xor (inputs(251)));
    layer0_outputs(3393) <= (inputs(244)) and not (inputs(94));
    layer0_outputs(3394) <= (inputs(19)) or (inputs(123));
    layer0_outputs(3395) <= not(inputs(227));
    layer0_outputs(3396) <= (inputs(85)) and not (inputs(191));
    layer0_outputs(3397) <= (inputs(56)) xor (inputs(13));
    layer0_outputs(3398) <= (inputs(205)) or (inputs(198));
    layer0_outputs(3399) <= not((inputs(198)) and (inputs(198)));
    layer0_outputs(3400) <= inputs(176);
    layer0_outputs(3401) <= not((inputs(163)) or (inputs(127)));
    layer0_outputs(3402) <= inputs(58);
    layer0_outputs(3403) <= (inputs(76)) and not (inputs(238));
    layer0_outputs(3404) <= not(inputs(24));
    layer0_outputs(3405) <= (inputs(169)) and not (inputs(64));
    layer0_outputs(3406) <= not((inputs(53)) xor (inputs(101)));
    layer0_outputs(3407) <= inputs(129);
    layer0_outputs(3408) <= not((inputs(23)) xor (inputs(55)));
    layer0_outputs(3409) <= not(inputs(159));
    layer0_outputs(3410) <= inputs(47);
    layer0_outputs(3411) <= inputs(237);
    layer0_outputs(3412) <= not(inputs(20)) or (inputs(54));
    layer0_outputs(3413) <= (inputs(5)) or (inputs(52));
    layer0_outputs(3414) <= not((inputs(47)) or (inputs(40)));
    layer0_outputs(3415) <= not((inputs(249)) or (inputs(38)));
    layer0_outputs(3416) <= '1';
    layer0_outputs(3417) <= '1';
    layer0_outputs(3418) <= (inputs(190)) and not (inputs(129));
    layer0_outputs(3419) <= not((inputs(230)) xor (inputs(4)));
    layer0_outputs(3420) <= not(inputs(246)) or (inputs(43));
    layer0_outputs(3421) <= inputs(182);
    layer0_outputs(3422) <= not(inputs(234)) or (inputs(36));
    layer0_outputs(3423) <= not((inputs(22)) and (inputs(43)));
    layer0_outputs(3424) <= not((inputs(213)) or (inputs(64)));
    layer0_outputs(3425) <= not(inputs(149));
    layer0_outputs(3426) <= not((inputs(233)) or (inputs(236)));
    layer0_outputs(3427) <= (inputs(4)) or (inputs(185));
    layer0_outputs(3428) <= not(inputs(65));
    layer0_outputs(3429) <= inputs(26);
    layer0_outputs(3430) <= not((inputs(231)) xor (inputs(140)));
    layer0_outputs(3431) <= not(inputs(18)) or (inputs(143));
    layer0_outputs(3432) <= (inputs(50)) and not (inputs(30));
    layer0_outputs(3433) <= (inputs(169)) and (inputs(139));
    layer0_outputs(3434) <= (inputs(155)) and not (inputs(105));
    layer0_outputs(3435) <= not((inputs(235)) xor (inputs(9)));
    layer0_outputs(3436) <= (inputs(197)) and not (inputs(223));
    layer0_outputs(3437) <= (inputs(7)) or (inputs(64));
    layer0_outputs(3438) <= inputs(34);
    layer0_outputs(3439) <= not(inputs(234));
    layer0_outputs(3440) <= not(inputs(42));
    layer0_outputs(3441) <= not(inputs(159)) or (inputs(174));
    layer0_outputs(3442) <= (inputs(72)) and not (inputs(14));
    layer0_outputs(3443) <= not(inputs(176));
    layer0_outputs(3444) <= inputs(179);
    layer0_outputs(3445) <= not((inputs(4)) and (inputs(12)));
    layer0_outputs(3446) <= not(inputs(111)) or (inputs(32));
    layer0_outputs(3447) <= not((inputs(171)) and (inputs(177)));
    layer0_outputs(3448) <= not((inputs(97)) or (inputs(245)));
    layer0_outputs(3449) <= not((inputs(146)) or (inputs(255)));
    layer0_outputs(3450) <= (inputs(10)) xor (inputs(242));
    layer0_outputs(3451) <= not((inputs(207)) and (inputs(15)));
    layer0_outputs(3452) <= not((inputs(219)) xor (inputs(127)));
    layer0_outputs(3453) <= not((inputs(249)) and (inputs(0)));
    layer0_outputs(3454) <= (inputs(198)) and not (inputs(14));
    layer0_outputs(3455) <= not(inputs(8)) or (inputs(243));
    layer0_outputs(3456) <= inputs(23);
    layer0_outputs(3457) <= (inputs(51)) or (inputs(34));
    layer0_outputs(3458) <= not((inputs(195)) or (inputs(248)));
    layer0_outputs(3459) <= not(inputs(68));
    layer0_outputs(3460) <= (inputs(222)) xor (inputs(147));
    layer0_outputs(3461) <= (inputs(62)) or (inputs(97));
    layer0_outputs(3462) <= (inputs(60)) and not (inputs(17));
    layer0_outputs(3463) <= (inputs(80)) xor (inputs(81));
    layer0_outputs(3464) <= inputs(228);
    layer0_outputs(3465) <= (inputs(58)) xor (inputs(75));
    layer0_outputs(3466) <= (inputs(142)) or (inputs(186));
    layer0_outputs(3467) <= not((inputs(132)) or (inputs(27)));
    layer0_outputs(3468) <= not((inputs(176)) and (inputs(145)));
    layer0_outputs(3469) <= not((inputs(148)) or (inputs(145)));
    layer0_outputs(3470) <= not(inputs(8)) or (inputs(194));
    layer0_outputs(3471) <= inputs(48);
    layer0_outputs(3472) <= not((inputs(120)) and (inputs(224)));
    layer0_outputs(3473) <= (inputs(83)) or (inputs(176));
    layer0_outputs(3474) <= not((inputs(29)) or (inputs(16)));
    layer0_outputs(3475) <= not((inputs(60)) or (inputs(57)));
    layer0_outputs(3476) <= not(inputs(248));
    layer0_outputs(3477) <= inputs(97);
    layer0_outputs(3478) <= not(inputs(218));
    layer0_outputs(3479) <= (inputs(142)) or (inputs(2));
    layer0_outputs(3480) <= (inputs(204)) and not (inputs(81));
    layer0_outputs(3481) <= inputs(99);
    layer0_outputs(3482) <= (inputs(3)) xor (inputs(93));
    layer0_outputs(3483) <= inputs(220);
    layer0_outputs(3484) <= (inputs(122)) and not (inputs(2));
    layer0_outputs(3485) <= not(inputs(168));
    layer0_outputs(3486) <= inputs(235);
    layer0_outputs(3487) <= not(inputs(97));
    layer0_outputs(3488) <= not(inputs(233));
    layer0_outputs(3489) <= not((inputs(170)) or (inputs(237)));
    layer0_outputs(3490) <= not((inputs(208)) or (inputs(211)));
    layer0_outputs(3491) <= (inputs(21)) or (inputs(75));
    layer0_outputs(3492) <= not((inputs(153)) and (inputs(117)));
    layer0_outputs(3493) <= (inputs(145)) or (inputs(196));
    layer0_outputs(3494) <= (inputs(202)) and not (inputs(80));
    layer0_outputs(3495) <= (inputs(230)) xor (inputs(22));
    layer0_outputs(3496) <= (inputs(203)) and not (inputs(16));
    layer0_outputs(3497) <= (inputs(187)) and not (inputs(160));
    layer0_outputs(3498) <= not(inputs(101));
    layer0_outputs(3499) <= not((inputs(250)) xor (inputs(27)));
    layer0_outputs(3500) <= not((inputs(49)) xor (inputs(117)));
    layer0_outputs(3501) <= not(inputs(166)) or (inputs(1));
    layer0_outputs(3502) <= not(inputs(228)) or (inputs(117));
    layer0_outputs(3503) <= not(inputs(140));
    layer0_outputs(3504) <= not(inputs(181));
    layer0_outputs(3505) <= (inputs(223)) xor (inputs(208));
    layer0_outputs(3506) <= (inputs(195)) and not (inputs(94));
    layer0_outputs(3507) <= not((inputs(242)) xor (inputs(167)));
    layer0_outputs(3508) <= (inputs(168)) and not (inputs(243));
    layer0_outputs(3509) <= not((inputs(30)) or (inputs(240)));
    layer0_outputs(3510) <= (inputs(242)) or (inputs(19));
    layer0_outputs(3511) <= not((inputs(92)) xor (inputs(66)));
    layer0_outputs(3512) <= not((inputs(219)) or (inputs(15)));
    layer0_outputs(3513) <= not(inputs(180));
    layer0_outputs(3514) <= (inputs(233)) xor (inputs(27));
    layer0_outputs(3515) <= not(inputs(13)) or (inputs(116));
    layer0_outputs(3516) <= (inputs(200)) and not (inputs(218));
    layer0_outputs(3517) <= not(inputs(140)) or (inputs(78));
    layer0_outputs(3518) <= not(inputs(104));
    layer0_outputs(3519) <= not(inputs(170));
    layer0_outputs(3520) <= (inputs(9)) and not (inputs(251));
    layer0_outputs(3521) <= (inputs(240)) or (inputs(2));
    layer0_outputs(3522) <= inputs(142);
    layer0_outputs(3523) <= not((inputs(128)) or (inputs(29)));
    layer0_outputs(3524) <= not(inputs(151));
    layer0_outputs(3525) <= (inputs(178)) or (inputs(151));
    layer0_outputs(3526) <= not(inputs(43));
    layer0_outputs(3527) <= not(inputs(246));
    layer0_outputs(3528) <= (inputs(207)) or (inputs(148));
    layer0_outputs(3529) <= not((inputs(159)) or (inputs(247)));
    layer0_outputs(3530) <= not(inputs(10)) or (inputs(12));
    layer0_outputs(3531) <= (inputs(214)) and (inputs(92));
    layer0_outputs(3532) <= not(inputs(201));
    layer0_outputs(3533) <= not(inputs(115)) or (inputs(56));
    layer0_outputs(3534) <= inputs(228);
    layer0_outputs(3535) <= not(inputs(101));
    layer0_outputs(3536) <= inputs(223);
    layer0_outputs(3537) <= (inputs(236)) or (inputs(36));
    layer0_outputs(3538) <= (inputs(52)) and not (inputs(32));
    layer0_outputs(3539) <= not(inputs(96)) or (inputs(238));
    layer0_outputs(3540) <= (inputs(195)) or (inputs(194));
    layer0_outputs(3541) <= not((inputs(208)) xor (inputs(1)));
    layer0_outputs(3542) <= not((inputs(174)) xor (inputs(186)));
    layer0_outputs(3543) <= (inputs(61)) and not (inputs(5));
    layer0_outputs(3544) <= not(inputs(104)) or (inputs(3));
    layer0_outputs(3545) <= inputs(145);
    layer0_outputs(3546) <= (inputs(225)) or (inputs(49));
    layer0_outputs(3547) <= not(inputs(78));
    layer0_outputs(3548) <= (inputs(118)) or (inputs(11));
    layer0_outputs(3549) <= inputs(50);
    layer0_outputs(3550) <= not(inputs(7));
    layer0_outputs(3551) <= not((inputs(161)) or (inputs(148)));
    layer0_outputs(3552) <= not(inputs(152)) or (inputs(1));
    layer0_outputs(3553) <= not((inputs(68)) xor (inputs(131)));
    layer0_outputs(3554) <= (inputs(201)) and not (inputs(114));
    layer0_outputs(3555) <= not(inputs(122));
    layer0_outputs(3556) <= not(inputs(104));
    layer0_outputs(3557) <= inputs(20);
    layer0_outputs(3558) <= inputs(137);
    layer0_outputs(3559) <= (inputs(192)) or (inputs(249));
    layer0_outputs(3560) <= not(inputs(178));
    layer0_outputs(3561) <= not(inputs(197));
    layer0_outputs(3562) <= not((inputs(5)) or (inputs(175)));
    layer0_outputs(3563) <= not(inputs(11));
    layer0_outputs(3564) <= not(inputs(121)) or (inputs(189));
    layer0_outputs(3565) <= not(inputs(72)) or (inputs(213));
    layer0_outputs(3566) <= (inputs(100)) and not (inputs(14));
    layer0_outputs(3567) <= not(inputs(78)) or (inputs(72));
    layer0_outputs(3568) <= (inputs(155)) and not (inputs(61));
    layer0_outputs(3569) <= '1';
    layer0_outputs(3570) <= not(inputs(89));
    layer0_outputs(3571) <= (inputs(126)) xor (inputs(116));
    layer0_outputs(3572) <= not(inputs(179)) or (inputs(82));
    layer0_outputs(3573) <= (inputs(71)) and not (inputs(221));
    layer0_outputs(3574) <= (inputs(163)) or (inputs(97));
    layer0_outputs(3575) <= inputs(155);
    layer0_outputs(3576) <= not((inputs(212)) or (inputs(246)));
    layer0_outputs(3577) <= inputs(87);
    layer0_outputs(3578) <= not((inputs(131)) xor (inputs(255)));
    layer0_outputs(3579) <= (inputs(54)) or (inputs(49));
    layer0_outputs(3580) <= not((inputs(234)) xor (inputs(66)));
    layer0_outputs(3581) <= (inputs(70)) or (inputs(145));
    layer0_outputs(3582) <= not(inputs(66));
    layer0_outputs(3583) <= (inputs(59)) and not (inputs(150));
    layer0_outputs(3584) <= (inputs(139)) or (inputs(98));
    layer0_outputs(3585) <= (inputs(49)) or (inputs(159));
    layer0_outputs(3586) <= (inputs(22)) and not (inputs(221));
    layer0_outputs(3587) <= (inputs(236)) or (inputs(172));
    layer0_outputs(3588) <= not(inputs(162));
    layer0_outputs(3589) <= not(inputs(165));
    layer0_outputs(3590) <= (inputs(227)) or (inputs(192));
    layer0_outputs(3591) <= not(inputs(69));
    layer0_outputs(3592) <= not(inputs(91));
    layer0_outputs(3593) <= not(inputs(46)) or (inputs(107));
    layer0_outputs(3594) <= (inputs(30)) or (inputs(46));
    layer0_outputs(3595) <= not((inputs(109)) or (inputs(145)));
    layer0_outputs(3596) <= (inputs(68)) and not (inputs(14));
    layer0_outputs(3597) <= inputs(43);
    layer0_outputs(3598) <= not((inputs(126)) or (inputs(70)));
    layer0_outputs(3599) <= not(inputs(241));
    layer0_outputs(3600) <= (inputs(11)) and not (inputs(156));
    layer0_outputs(3601) <= not(inputs(12)) or (inputs(140));
    layer0_outputs(3602) <= inputs(131);
    layer0_outputs(3603) <= (inputs(125)) and not (inputs(123));
    layer0_outputs(3604) <= (inputs(201)) and not (inputs(43));
    layer0_outputs(3605) <= not((inputs(167)) or (inputs(110)));
    layer0_outputs(3606) <= (inputs(62)) and not (inputs(3));
    layer0_outputs(3607) <= not((inputs(188)) or (inputs(156)));
    layer0_outputs(3608) <= not(inputs(19));
    layer0_outputs(3609) <= (inputs(13)) and (inputs(227));
    layer0_outputs(3610) <= (inputs(122)) and (inputs(226));
    layer0_outputs(3611) <= not(inputs(72));
    layer0_outputs(3612) <= (inputs(94)) or (inputs(174));
    layer0_outputs(3613) <= not(inputs(75)) or (inputs(224));
    layer0_outputs(3614) <= '1';
    layer0_outputs(3615) <= (inputs(62)) or (inputs(232));
    layer0_outputs(3616) <= not((inputs(11)) or (inputs(254)));
    layer0_outputs(3617) <= not(inputs(201)) or (inputs(86));
    layer0_outputs(3618) <= (inputs(162)) and not (inputs(65));
    layer0_outputs(3619) <= inputs(74);
    layer0_outputs(3620) <= inputs(125);
    layer0_outputs(3621) <= (inputs(222)) or (inputs(230));
    layer0_outputs(3622) <= not(inputs(6)) or (inputs(142));
    layer0_outputs(3623) <= inputs(22);
    layer0_outputs(3624) <= not(inputs(181));
    layer0_outputs(3625) <= (inputs(34)) and not (inputs(125));
    layer0_outputs(3626) <= not(inputs(212));
    layer0_outputs(3627) <= not(inputs(151));
    layer0_outputs(3628) <= (inputs(164)) xor (inputs(191));
    layer0_outputs(3629) <= (inputs(86)) and not (inputs(141));
    layer0_outputs(3630) <= not(inputs(47));
    layer0_outputs(3631) <= inputs(249);
    layer0_outputs(3632) <= inputs(95);
    layer0_outputs(3633) <= not((inputs(180)) or (inputs(246)));
    layer0_outputs(3634) <= (inputs(176)) or (inputs(79));
    layer0_outputs(3635) <= not((inputs(152)) or (inputs(130)));
    layer0_outputs(3636) <= (inputs(20)) and not (inputs(176));
    layer0_outputs(3637) <= not(inputs(244));
    layer0_outputs(3638) <= inputs(195);
    layer0_outputs(3639) <= inputs(84);
    layer0_outputs(3640) <= not((inputs(147)) xor (inputs(164)));
    layer0_outputs(3641) <= (inputs(249)) and not (inputs(73));
    layer0_outputs(3642) <= inputs(169);
    layer0_outputs(3643) <= (inputs(73)) and (inputs(64));
    layer0_outputs(3644) <= (inputs(145)) and not (inputs(14));
    layer0_outputs(3645) <= (inputs(59)) xor (inputs(29));
    layer0_outputs(3646) <= inputs(189);
    layer0_outputs(3647) <= not(inputs(30));
    layer0_outputs(3648) <= '1';
    layer0_outputs(3649) <= (inputs(249)) or (inputs(210));
    layer0_outputs(3650) <= not((inputs(37)) and (inputs(108)));
    layer0_outputs(3651) <= not(inputs(28));
    layer0_outputs(3652) <= not((inputs(133)) or (inputs(80)));
    layer0_outputs(3653) <= inputs(29);
    layer0_outputs(3654) <= not(inputs(176)) or (inputs(48));
    layer0_outputs(3655) <= not((inputs(47)) xor (inputs(212)));
    layer0_outputs(3656) <= (inputs(131)) and not (inputs(34));
    layer0_outputs(3657) <= not((inputs(105)) or (inputs(62)));
    layer0_outputs(3658) <= not(inputs(8));
    layer0_outputs(3659) <= inputs(243);
    layer0_outputs(3660) <= (inputs(165)) or (inputs(167));
    layer0_outputs(3661) <= (inputs(226)) and not (inputs(239));
    layer0_outputs(3662) <= not(inputs(24));
    layer0_outputs(3663) <= not(inputs(97));
    layer0_outputs(3664) <= not(inputs(95));
    layer0_outputs(3665) <= '1';
    layer0_outputs(3666) <= not((inputs(128)) or (inputs(201)));
    layer0_outputs(3667) <= not((inputs(32)) or (inputs(36)));
    layer0_outputs(3668) <= not(inputs(2));
    layer0_outputs(3669) <= (inputs(80)) or (inputs(133));
    layer0_outputs(3670) <= not((inputs(218)) xor (inputs(166)));
    layer0_outputs(3671) <= not((inputs(184)) or (inputs(78)));
    layer0_outputs(3672) <= not(inputs(183)) or (inputs(208));
    layer0_outputs(3673) <= not((inputs(140)) or (inputs(33)));
    layer0_outputs(3674) <= not(inputs(146)) or (inputs(227));
    layer0_outputs(3675) <= not(inputs(50)) or (inputs(15));
    layer0_outputs(3676) <= (inputs(161)) and not (inputs(33));
    layer0_outputs(3677) <= (inputs(180)) and not (inputs(143));
    layer0_outputs(3678) <= (inputs(135)) and not (inputs(113));
    layer0_outputs(3679) <= (inputs(93)) xor (inputs(177));
    layer0_outputs(3680) <= not(inputs(72)) or (inputs(222));
    layer0_outputs(3681) <= (inputs(219)) and not (inputs(96));
    layer0_outputs(3682) <= (inputs(246)) xor (inputs(1));
    layer0_outputs(3683) <= (inputs(8)) xor (inputs(28));
    layer0_outputs(3684) <= not(inputs(164));
    layer0_outputs(3685) <= not(inputs(195));
    layer0_outputs(3686) <= not(inputs(21));
    layer0_outputs(3687) <= (inputs(9)) or (inputs(39));
    layer0_outputs(3688) <= inputs(85);
    layer0_outputs(3689) <= not(inputs(93));
    layer0_outputs(3690) <= inputs(114);
    layer0_outputs(3691) <= not(inputs(92));
    layer0_outputs(3692) <= inputs(72);
    layer0_outputs(3693) <= inputs(33);
    layer0_outputs(3694) <= not((inputs(119)) xor (inputs(178)));
    layer0_outputs(3695) <= not((inputs(86)) xor (inputs(50)));
    layer0_outputs(3696) <= not(inputs(200));
    layer0_outputs(3697) <= inputs(208);
    layer0_outputs(3698) <= inputs(101);
    layer0_outputs(3699) <= not(inputs(122));
    layer0_outputs(3700) <= not(inputs(88));
    layer0_outputs(3701) <= not(inputs(172));
    layer0_outputs(3702) <= inputs(101);
    layer0_outputs(3703) <= not((inputs(185)) xor (inputs(83)));
    layer0_outputs(3704) <= inputs(210);
    layer0_outputs(3705) <= (inputs(69)) and not (inputs(35));
    layer0_outputs(3706) <= not(inputs(92));
    layer0_outputs(3707) <= (inputs(89)) xor (inputs(173));
    layer0_outputs(3708) <= (inputs(127)) or (inputs(239));
    layer0_outputs(3709) <= not(inputs(121)) or (inputs(218));
    layer0_outputs(3710) <= not((inputs(59)) or (inputs(44)));
    layer0_outputs(3711) <= inputs(100);
    layer0_outputs(3712) <= (inputs(224)) or (inputs(157));
    layer0_outputs(3713) <= not((inputs(221)) or (inputs(154)));
    layer0_outputs(3714) <= not((inputs(240)) or (inputs(254)));
    layer0_outputs(3715) <= not((inputs(33)) or (inputs(215)));
    layer0_outputs(3716) <= not(inputs(98));
    layer0_outputs(3717) <= (inputs(17)) or (inputs(120));
    layer0_outputs(3718) <= inputs(108);
    layer0_outputs(3719) <= (inputs(131)) and not (inputs(40));
    layer0_outputs(3720) <= not((inputs(209)) or (inputs(208)));
    layer0_outputs(3721) <= (inputs(133)) or (inputs(187));
    layer0_outputs(3722) <= inputs(77);
    layer0_outputs(3723) <= inputs(139);
    layer0_outputs(3724) <= (inputs(242)) or (inputs(250));
    layer0_outputs(3725) <= not(inputs(156)) or (inputs(40));
    layer0_outputs(3726) <= not((inputs(123)) or (inputs(222)));
    layer0_outputs(3727) <= not((inputs(95)) xor (inputs(104)));
    layer0_outputs(3728) <= (inputs(246)) and not (inputs(94));
    layer0_outputs(3729) <= not(inputs(179));
    layer0_outputs(3730) <= not(inputs(49)) or (inputs(11));
    layer0_outputs(3731) <= not((inputs(204)) or (inputs(48)));
    layer0_outputs(3732) <= (inputs(186)) or (inputs(188));
    layer0_outputs(3733) <= (inputs(253)) or (inputs(236));
    layer0_outputs(3734) <= (inputs(180)) or (inputs(111));
    layer0_outputs(3735) <= inputs(192);
    layer0_outputs(3736) <= not((inputs(245)) xor (inputs(204)));
    layer0_outputs(3737) <= (inputs(115)) and not (inputs(224));
    layer0_outputs(3738) <= (inputs(69)) and not (inputs(209));
    layer0_outputs(3739) <= not(inputs(117)) or (inputs(254));
    layer0_outputs(3740) <= (inputs(205)) and not (inputs(193));
    layer0_outputs(3741) <= not(inputs(23));
    layer0_outputs(3742) <= (inputs(243)) or (inputs(63));
    layer0_outputs(3743) <= not(inputs(129));
    layer0_outputs(3744) <= not((inputs(207)) xor (inputs(107)));
    layer0_outputs(3745) <= inputs(140);
    layer0_outputs(3746) <= not((inputs(226)) xor (inputs(138)));
    layer0_outputs(3747) <= not(inputs(117));
    layer0_outputs(3748) <= (inputs(39)) and not (inputs(128));
    layer0_outputs(3749) <= (inputs(251)) or (inputs(184));
    layer0_outputs(3750) <= inputs(153);
    layer0_outputs(3751) <= (inputs(26)) and not (inputs(104));
    layer0_outputs(3752) <= not(inputs(155)) or (inputs(44));
    layer0_outputs(3753) <= not(inputs(146)) or (inputs(191));
    layer0_outputs(3754) <= (inputs(106)) and not (inputs(252));
    layer0_outputs(3755) <= not(inputs(214));
    layer0_outputs(3756) <= not(inputs(105));
    layer0_outputs(3757) <= not((inputs(124)) or (inputs(142)));
    layer0_outputs(3758) <= (inputs(126)) and (inputs(140));
    layer0_outputs(3759) <= (inputs(164)) and (inputs(71));
    layer0_outputs(3760) <= (inputs(135)) and not (inputs(127));
    layer0_outputs(3761) <= inputs(107);
    layer0_outputs(3762) <= (inputs(223)) and (inputs(254));
    layer0_outputs(3763) <= not(inputs(153));
    layer0_outputs(3764) <= not((inputs(218)) or (inputs(205)));
    layer0_outputs(3765) <= not(inputs(148));
    layer0_outputs(3766) <= not(inputs(42)) or (inputs(69));
    layer0_outputs(3767) <= (inputs(123)) and not (inputs(127));
    layer0_outputs(3768) <= (inputs(223)) or (inputs(209));
    layer0_outputs(3769) <= not(inputs(209)) or (inputs(18));
    layer0_outputs(3770) <= not(inputs(246));
    layer0_outputs(3771) <= '0';
    layer0_outputs(3772) <= not((inputs(229)) and (inputs(248)));
    layer0_outputs(3773) <= not((inputs(47)) and (inputs(206)));
    layer0_outputs(3774) <= not((inputs(145)) or (inputs(13)));
    layer0_outputs(3775) <= not(inputs(188)) or (inputs(109));
    layer0_outputs(3776) <= inputs(176);
    layer0_outputs(3777) <= not((inputs(160)) or (inputs(100)));
    layer0_outputs(3778) <= not(inputs(215)) or (inputs(110));
    layer0_outputs(3779) <= (inputs(60)) and not (inputs(220));
    layer0_outputs(3780) <= not((inputs(193)) xor (inputs(221)));
    layer0_outputs(3781) <= inputs(71);
    layer0_outputs(3782) <= (inputs(15)) or (inputs(254));
    layer0_outputs(3783) <= inputs(135);
    layer0_outputs(3784) <= (inputs(155)) or (inputs(129));
    layer0_outputs(3785) <= not(inputs(228)) or (inputs(15));
    layer0_outputs(3786) <= not(inputs(75));
    layer0_outputs(3787) <= (inputs(219)) xor (inputs(154));
    layer0_outputs(3788) <= not(inputs(166));
    layer0_outputs(3789) <= not((inputs(114)) xor (inputs(67)));
    layer0_outputs(3790) <= not(inputs(117));
    layer0_outputs(3791) <= (inputs(131)) or (inputs(188));
    layer0_outputs(3792) <= (inputs(206)) xor (inputs(133));
    layer0_outputs(3793) <= (inputs(43)) and not (inputs(147));
    layer0_outputs(3794) <= inputs(193);
    layer0_outputs(3795) <= not((inputs(49)) xor (inputs(93)));
    layer0_outputs(3796) <= inputs(35);
    layer0_outputs(3797) <= not((inputs(179)) xor (inputs(106)));
    layer0_outputs(3798) <= not((inputs(111)) xor (inputs(98)));
    layer0_outputs(3799) <= not((inputs(186)) or (inputs(242)));
    layer0_outputs(3800) <= inputs(53);
    layer0_outputs(3801) <= (inputs(52)) xor (inputs(82));
    layer0_outputs(3802) <= (inputs(120)) or (inputs(153));
    layer0_outputs(3803) <= inputs(227);
    layer0_outputs(3804) <= not(inputs(166));
    layer0_outputs(3805) <= inputs(124);
    layer0_outputs(3806) <= (inputs(72)) or (inputs(143));
    layer0_outputs(3807) <= (inputs(7)) xor (inputs(52));
    layer0_outputs(3808) <= not(inputs(28)) or (inputs(102));
    layer0_outputs(3809) <= inputs(62);
    layer0_outputs(3810) <= inputs(100);
    layer0_outputs(3811) <= not((inputs(179)) or (inputs(71)));
    layer0_outputs(3812) <= not(inputs(39)) or (inputs(228));
    layer0_outputs(3813) <= not(inputs(128));
    layer0_outputs(3814) <= (inputs(105)) and not (inputs(32));
    layer0_outputs(3815) <= not(inputs(166));
    layer0_outputs(3816) <= not((inputs(166)) and (inputs(168)));
    layer0_outputs(3817) <= (inputs(74)) or (inputs(123));
    layer0_outputs(3818) <= inputs(226);
    layer0_outputs(3819) <= not((inputs(77)) or (inputs(7)));
    layer0_outputs(3820) <= not(inputs(212)) or (inputs(66));
    layer0_outputs(3821) <= (inputs(57)) and not (inputs(144));
    layer0_outputs(3822) <= not((inputs(120)) xor (inputs(87)));
    layer0_outputs(3823) <= not((inputs(98)) or (inputs(163)));
    layer0_outputs(3824) <= (inputs(53)) or (inputs(62));
    layer0_outputs(3825) <= inputs(155);
    layer0_outputs(3826) <= '0';
    layer0_outputs(3827) <= inputs(86);
    layer0_outputs(3828) <= not(inputs(167));
    layer0_outputs(3829) <= inputs(106);
    layer0_outputs(3830) <= not(inputs(213));
    layer0_outputs(3831) <= not((inputs(233)) and (inputs(59)));
    layer0_outputs(3832) <= not(inputs(196)) or (inputs(33));
    layer0_outputs(3833) <= inputs(79);
    layer0_outputs(3834) <= (inputs(205)) xor (inputs(186));
    layer0_outputs(3835) <= inputs(252);
    layer0_outputs(3836) <= not((inputs(143)) or (inputs(145)));
    layer0_outputs(3837) <= inputs(69);
    layer0_outputs(3838) <= not((inputs(234)) or (inputs(18)));
    layer0_outputs(3839) <= '0';
    layer0_outputs(3840) <= '1';
    layer0_outputs(3841) <= inputs(30);
    layer0_outputs(3842) <= not((inputs(102)) or (inputs(49)));
    layer0_outputs(3843) <= (inputs(96)) or (inputs(114));
    layer0_outputs(3844) <= not((inputs(239)) or (inputs(131)));
    layer0_outputs(3845) <= not(inputs(22)) or (inputs(230));
    layer0_outputs(3846) <= not(inputs(222));
    layer0_outputs(3847) <= inputs(41);
    layer0_outputs(3848) <= not(inputs(93));
    layer0_outputs(3849) <= not((inputs(196)) xor (inputs(242)));
    layer0_outputs(3850) <= not(inputs(205));
    layer0_outputs(3851) <= (inputs(30)) or (inputs(117));
    layer0_outputs(3852) <= not((inputs(220)) xor (inputs(6)));
    layer0_outputs(3853) <= not(inputs(105));
    layer0_outputs(3854) <= inputs(1);
    layer0_outputs(3855) <= (inputs(178)) or (inputs(186));
    layer0_outputs(3856) <= not((inputs(50)) xor (inputs(177)));
    layer0_outputs(3857) <= (inputs(127)) or (inputs(122));
    layer0_outputs(3858) <= inputs(99);
    layer0_outputs(3859) <= not((inputs(235)) xor (inputs(61)));
    layer0_outputs(3860) <= (inputs(1)) or (inputs(192));
    layer0_outputs(3861) <= '1';
    layer0_outputs(3862) <= (inputs(189)) or (inputs(174));
    layer0_outputs(3863) <= not((inputs(226)) or (inputs(233)));
    layer0_outputs(3864) <= not(inputs(69));
    layer0_outputs(3865) <= (inputs(66)) xor (inputs(68));
    layer0_outputs(3866) <= inputs(139);
    layer0_outputs(3867) <= (inputs(59)) and not (inputs(237));
    layer0_outputs(3868) <= not(inputs(215));
    layer0_outputs(3869) <= not((inputs(95)) or (inputs(173)));
    layer0_outputs(3870) <= not((inputs(94)) or (inputs(31)));
    layer0_outputs(3871) <= (inputs(37)) xor (inputs(12));
    layer0_outputs(3872) <= inputs(245);
    layer0_outputs(3873) <= (inputs(150)) xor (inputs(107));
    layer0_outputs(3874) <= (inputs(74)) or (inputs(252));
    layer0_outputs(3875) <= inputs(236);
    layer0_outputs(3876) <= not(inputs(69)) or (inputs(77));
    layer0_outputs(3877) <= not(inputs(91)) or (inputs(225));
    layer0_outputs(3878) <= not((inputs(205)) or (inputs(211)));
    layer0_outputs(3879) <= (inputs(209)) and not (inputs(123));
    layer0_outputs(3880) <= not(inputs(99)) or (inputs(64));
    layer0_outputs(3881) <= inputs(115);
    layer0_outputs(3882) <= not(inputs(91));
    layer0_outputs(3883) <= (inputs(85)) and not (inputs(177));
    layer0_outputs(3884) <= not(inputs(232));
    layer0_outputs(3885) <= (inputs(142)) or (inputs(101));
    layer0_outputs(3886) <= (inputs(108)) and not (inputs(15));
    layer0_outputs(3887) <= not((inputs(227)) xor (inputs(24)));
    layer0_outputs(3888) <= not((inputs(239)) or (inputs(189)));
    layer0_outputs(3889) <= (inputs(7)) and not (inputs(1));
    layer0_outputs(3890) <= (inputs(130)) or (inputs(219));
    layer0_outputs(3891) <= (inputs(93)) xor (inputs(53));
    layer0_outputs(3892) <= not(inputs(180));
    layer0_outputs(3893) <= not((inputs(46)) xor (inputs(59)));
    layer0_outputs(3894) <= not(inputs(164)) or (inputs(17));
    layer0_outputs(3895) <= not((inputs(233)) or (inputs(77)));
    layer0_outputs(3896) <= (inputs(160)) or (inputs(190));
    layer0_outputs(3897) <= (inputs(115)) and not (inputs(143));
    layer0_outputs(3898) <= (inputs(50)) or (inputs(31));
    layer0_outputs(3899) <= '1';
    layer0_outputs(3900) <= not(inputs(86));
    layer0_outputs(3901) <= not(inputs(14));
    layer0_outputs(3902) <= (inputs(209)) or (inputs(120));
    layer0_outputs(3903) <= (inputs(102)) and not (inputs(179));
    layer0_outputs(3904) <= not(inputs(238));
    layer0_outputs(3905) <= not(inputs(194)) or (inputs(248));
    layer0_outputs(3906) <= (inputs(191)) or (inputs(224));
    layer0_outputs(3907) <= not((inputs(32)) or (inputs(143)));
    layer0_outputs(3908) <= inputs(230);
    layer0_outputs(3909) <= not((inputs(48)) or (inputs(220)));
    layer0_outputs(3910) <= not((inputs(158)) or (inputs(61)));
    layer0_outputs(3911) <= not((inputs(153)) or (inputs(255)));
    layer0_outputs(3912) <= not(inputs(119)) or (inputs(110));
    layer0_outputs(3913) <= (inputs(30)) or (inputs(37));
    layer0_outputs(3914) <= not(inputs(122));
    layer0_outputs(3915) <= (inputs(48)) or (inputs(11));
    layer0_outputs(3916) <= (inputs(115)) and not (inputs(63));
    layer0_outputs(3917) <= inputs(4);
    layer0_outputs(3918) <= not(inputs(43)) or (inputs(71));
    layer0_outputs(3919) <= not(inputs(68));
    layer0_outputs(3920) <= inputs(167);
    layer0_outputs(3921) <= not((inputs(248)) and (inputs(187)));
    layer0_outputs(3922) <= not((inputs(197)) xor (inputs(1)));
    layer0_outputs(3923) <= (inputs(49)) or (inputs(229));
    layer0_outputs(3924) <= not((inputs(247)) or (inputs(214)));
    layer0_outputs(3925) <= not(inputs(233)) or (inputs(28));
    layer0_outputs(3926) <= not(inputs(213));
    layer0_outputs(3927) <= not(inputs(110));
    layer0_outputs(3928) <= not(inputs(25)) or (inputs(197));
    layer0_outputs(3929) <= not(inputs(249));
    layer0_outputs(3930) <= not((inputs(118)) or (inputs(36)));
    layer0_outputs(3931) <= inputs(101);
    layer0_outputs(3932) <= (inputs(94)) or (inputs(253));
    layer0_outputs(3933) <= inputs(110);
    layer0_outputs(3934) <= (inputs(139)) or (inputs(40));
    layer0_outputs(3935) <= not((inputs(114)) or (inputs(158)));
    layer0_outputs(3936) <= not((inputs(68)) or (inputs(224)));
    layer0_outputs(3937) <= (inputs(73)) or (inputs(72));
    layer0_outputs(3938) <= not((inputs(251)) or (inputs(217)));
    layer0_outputs(3939) <= not(inputs(234));
    layer0_outputs(3940) <= not((inputs(189)) or (inputs(26)));
    layer0_outputs(3941) <= not((inputs(239)) xor (inputs(173)));
    layer0_outputs(3942) <= (inputs(175)) xor (inputs(34));
    layer0_outputs(3943) <= inputs(194);
    layer0_outputs(3944) <= not((inputs(213)) or (inputs(241)));
    layer0_outputs(3945) <= (inputs(111)) or (inputs(52));
    layer0_outputs(3946) <= not(inputs(105));
    layer0_outputs(3947) <= not(inputs(45)) or (inputs(252));
    layer0_outputs(3948) <= inputs(21);
    layer0_outputs(3949) <= not(inputs(119));
    layer0_outputs(3950) <= (inputs(62)) or (inputs(83));
    layer0_outputs(3951) <= (inputs(102)) or (inputs(13));
    layer0_outputs(3952) <= inputs(133);
    layer0_outputs(3953) <= (inputs(132)) or (inputs(241));
    layer0_outputs(3954) <= (inputs(213)) and not (inputs(106));
    layer0_outputs(3955) <= (inputs(73)) and not (inputs(232));
    layer0_outputs(3956) <= (inputs(133)) or (inputs(166));
    layer0_outputs(3957) <= not((inputs(220)) or (inputs(163)));
    layer0_outputs(3958) <= not((inputs(159)) or (inputs(214)));
    layer0_outputs(3959) <= not((inputs(124)) xor (inputs(107)));
    layer0_outputs(3960) <= not(inputs(123)) or (inputs(148));
    layer0_outputs(3961) <= not(inputs(99));
    layer0_outputs(3962) <= (inputs(144)) or (inputs(186));
    layer0_outputs(3963) <= inputs(231);
    layer0_outputs(3964) <= (inputs(231)) xor (inputs(199));
    layer0_outputs(3965) <= (inputs(99)) or (inputs(46));
    layer0_outputs(3966) <= not((inputs(122)) xor (inputs(89)));
    layer0_outputs(3967) <= not((inputs(108)) or (inputs(110)));
    layer0_outputs(3968) <= not(inputs(185)) or (inputs(43));
    layer0_outputs(3969) <= not(inputs(98)) or (inputs(32));
    layer0_outputs(3970) <= inputs(171);
    layer0_outputs(3971) <= not((inputs(44)) xor (inputs(126)));
    layer0_outputs(3972) <= not(inputs(254));
    layer0_outputs(3973) <= (inputs(212)) xor (inputs(11));
    layer0_outputs(3974) <= (inputs(131)) xor (inputs(209));
    layer0_outputs(3975) <= not(inputs(152));
    layer0_outputs(3976) <= inputs(152);
    layer0_outputs(3977) <= not((inputs(189)) xor (inputs(109)));
    layer0_outputs(3978) <= not(inputs(77)) or (inputs(61));
    layer0_outputs(3979) <= inputs(130);
    layer0_outputs(3980) <= inputs(101);
    layer0_outputs(3981) <= not(inputs(226));
    layer0_outputs(3982) <= not(inputs(122));
    layer0_outputs(3983) <= inputs(76);
    layer0_outputs(3984) <= not(inputs(70));
    layer0_outputs(3985) <= inputs(105);
    layer0_outputs(3986) <= (inputs(131)) and not (inputs(48));
    layer0_outputs(3987) <= not(inputs(4));
    layer0_outputs(3988) <= (inputs(168)) and not (inputs(79));
    layer0_outputs(3989) <= (inputs(102)) and not (inputs(174));
    layer0_outputs(3990) <= not((inputs(92)) xor (inputs(126)));
    layer0_outputs(3991) <= (inputs(73)) xor (inputs(94));
    layer0_outputs(3992) <= (inputs(36)) xor (inputs(4));
    layer0_outputs(3993) <= (inputs(64)) or (inputs(108));
    layer0_outputs(3994) <= not(inputs(168));
    layer0_outputs(3995) <= (inputs(234)) and not (inputs(146));
    layer0_outputs(3996) <= not((inputs(192)) or (inputs(223)));
    layer0_outputs(3997) <= not((inputs(219)) and (inputs(229)));
    layer0_outputs(3998) <= (inputs(53)) or (inputs(46));
    layer0_outputs(3999) <= not((inputs(16)) or (inputs(184)));
    layer0_outputs(4000) <= inputs(113);
    layer0_outputs(4001) <= not(inputs(221)) or (inputs(158));
    layer0_outputs(4002) <= not(inputs(92));
    layer0_outputs(4003) <= inputs(23);
    layer0_outputs(4004) <= inputs(24);
    layer0_outputs(4005) <= inputs(164);
    layer0_outputs(4006) <= not(inputs(98));
    layer0_outputs(4007) <= (inputs(147)) and not (inputs(63));
    layer0_outputs(4008) <= inputs(148);
    layer0_outputs(4009) <= inputs(191);
    layer0_outputs(4010) <= not((inputs(221)) xor (inputs(72)));
    layer0_outputs(4011) <= not(inputs(155));
    layer0_outputs(4012) <= (inputs(233)) and not (inputs(18));
    layer0_outputs(4013) <= not((inputs(91)) or (inputs(168)));
    layer0_outputs(4014) <= (inputs(148)) xor (inputs(216));
    layer0_outputs(4015) <= not(inputs(249));
    layer0_outputs(4016) <= inputs(48);
    layer0_outputs(4017) <= not(inputs(70)) or (inputs(35));
    layer0_outputs(4018) <= (inputs(197)) or (inputs(250));
    layer0_outputs(4019) <= not(inputs(76));
    layer0_outputs(4020) <= not((inputs(44)) or (inputs(172)));
    layer0_outputs(4021) <= not((inputs(88)) and (inputs(88)));
    layer0_outputs(4022) <= inputs(14);
    layer0_outputs(4023) <= inputs(164);
    layer0_outputs(4024) <= (inputs(186)) and not (inputs(57));
    layer0_outputs(4025) <= (inputs(74)) and not (inputs(101));
    layer0_outputs(4026) <= '0';
    layer0_outputs(4027) <= not(inputs(21)) or (inputs(144));
    layer0_outputs(4028) <= inputs(59);
    layer0_outputs(4029) <= (inputs(89)) xor (inputs(91));
    layer0_outputs(4030) <= inputs(155);
    layer0_outputs(4031) <= not((inputs(220)) or (inputs(56)));
    layer0_outputs(4032) <= not(inputs(70));
    layer0_outputs(4033) <= inputs(106);
    layer0_outputs(4034) <= (inputs(141)) or (inputs(179));
    layer0_outputs(4035) <= not((inputs(51)) or (inputs(127)));
    layer0_outputs(4036) <= inputs(181);
    layer0_outputs(4037) <= not((inputs(68)) xor (inputs(64)));
    layer0_outputs(4038) <= not((inputs(75)) or (inputs(206)));
    layer0_outputs(4039) <= not(inputs(192)) or (inputs(174));
    layer0_outputs(4040) <= not(inputs(230));
    layer0_outputs(4041) <= not(inputs(124));
    layer0_outputs(4042) <= not(inputs(164));
    layer0_outputs(4043) <= not((inputs(175)) or (inputs(26)));
    layer0_outputs(4044) <= (inputs(96)) xor (inputs(149));
    layer0_outputs(4045) <= inputs(103);
    layer0_outputs(4046) <= (inputs(37)) or (inputs(14));
    layer0_outputs(4047) <= not(inputs(132));
    layer0_outputs(4048) <= not((inputs(159)) or (inputs(161)));
    layer0_outputs(4049) <= not(inputs(177)) or (inputs(254));
    layer0_outputs(4050) <= inputs(73);
    layer0_outputs(4051) <= not((inputs(126)) or (inputs(7)));
    layer0_outputs(4052) <= (inputs(207)) or (inputs(142));
    layer0_outputs(4053) <= not(inputs(189));
    layer0_outputs(4054) <= (inputs(236)) and not (inputs(73));
    layer0_outputs(4055) <= '1';
    layer0_outputs(4056) <= (inputs(195)) or (inputs(2));
    layer0_outputs(4057) <= not(inputs(11)) or (inputs(44));
    layer0_outputs(4058) <= inputs(100);
    layer0_outputs(4059) <= not((inputs(200)) or (inputs(203)));
    layer0_outputs(4060) <= not(inputs(99));
    layer0_outputs(4061) <= not(inputs(102)) or (inputs(192));
    layer0_outputs(4062) <= (inputs(231)) xor (inputs(184));
    layer0_outputs(4063) <= not((inputs(204)) or (inputs(171)));
    layer0_outputs(4064) <= inputs(212);
    layer0_outputs(4065) <= not(inputs(197));
    layer0_outputs(4066) <= not(inputs(218));
    layer0_outputs(4067) <= not((inputs(107)) and (inputs(252)));
    layer0_outputs(4068) <= not((inputs(235)) and (inputs(52)));
    layer0_outputs(4069) <= not(inputs(124));
    layer0_outputs(4070) <= not(inputs(72));
    layer0_outputs(4071) <= not(inputs(236));
    layer0_outputs(4072) <= not((inputs(65)) xor (inputs(227)));
    layer0_outputs(4073) <= (inputs(206)) or (inputs(68));
    layer0_outputs(4074) <= not((inputs(40)) xor (inputs(88)));
    layer0_outputs(4075) <= not((inputs(9)) xor (inputs(56)));
    layer0_outputs(4076) <= (inputs(132)) and not (inputs(227));
    layer0_outputs(4077) <= (inputs(117)) and not (inputs(143));
    layer0_outputs(4078) <= '1';
    layer0_outputs(4079) <= not(inputs(94));
    layer0_outputs(4080) <= not(inputs(45)) or (inputs(239));
    layer0_outputs(4081) <= not(inputs(122));
    layer0_outputs(4082) <= not((inputs(77)) or (inputs(94)));
    layer0_outputs(4083) <= (inputs(246)) xor (inputs(94));
    layer0_outputs(4084) <= inputs(69);
    layer0_outputs(4085) <= not(inputs(102));
    layer0_outputs(4086) <= (inputs(252)) or (inputs(66));
    layer0_outputs(4087) <= (inputs(71)) and not (inputs(171));
    layer0_outputs(4088) <= not((inputs(228)) and (inputs(245)));
    layer0_outputs(4089) <= not(inputs(105)) or (inputs(178));
    layer0_outputs(4090) <= not(inputs(187));
    layer0_outputs(4091) <= not(inputs(107));
    layer0_outputs(4092) <= inputs(172);
    layer0_outputs(4093) <= not((inputs(20)) or (inputs(31)));
    layer0_outputs(4094) <= (inputs(189)) xor (inputs(209));
    layer0_outputs(4095) <= not(inputs(226)) or (inputs(101));
    layer0_outputs(4096) <= (inputs(78)) or (inputs(77));
    layer0_outputs(4097) <= inputs(151);
    layer0_outputs(4098) <= not(inputs(121));
    layer0_outputs(4099) <= not((inputs(18)) xor (inputs(188)));
    layer0_outputs(4100) <= (inputs(46)) or (inputs(192));
    layer0_outputs(4101) <= (inputs(136)) xor (inputs(149));
    layer0_outputs(4102) <= not(inputs(148));
    layer0_outputs(4103) <= not((inputs(184)) xor (inputs(213)));
    layer0_outputs(4104) <= inputs(177);
    layer0_outputs(4105) <= not((inputs(161)) xor (inputs(255)));
    layer0_outputs(4106) <= not((inputs(1)) xor (inputs(136)));
    layer0_outputs(4107) <= (inputs(30)) or (inputs(193));
    layer0_outputs(4108) <= not(inputs(104)) or (inputs(0));
    layer0_outputs(4109) <= inputs(164);
    layer0_outputs(4110) <= not((inputs(242)) or (inputs(19)));
    layer0_outputs(4111) <= not(inputs(94)) or (inputs(44));
    layer0_outputs(4112) <= not((inputs(123)) or (inputs(58)));
    layer0_outputs(4113) <= not(inputs(26));
    layer0_outputs(4114) <= inputs(25);
    layer0_outputs(4115) <= inputs(227);
    layer0_outputs(4116) <= (inputs(205)) or (inputs(201));
    layer0_outputs(4117) <= not(inputs(222));
    layer0_outputs(4118) <= (inputs(195)) and not (inputs(48));
    layer0_outputs(4119) <= (inputs(236)) or (inputs(129));
    layer0_outputs(4120) <= inputs(76);
    layer0_outputs(4121) <= not(inputs(88)) or (inputs(216));
    layer0_outputs(4122) <= not(inputs(166));
    layer0_outputs(4123) <= not((inputs(218)) or (inputs(240)));
    layer0_outputs(4124) <= not((inputs(59)) xor (inputs(105)));
    layer0_outputs(4125) <= not((inputs(217)) or (inputs(175)));
    layer0_outputs(4126) <= (inputs(192)) and not (inputs(254));
    layer0_outputs(4127) <= (inputs(99)) and not (inputs(44));
    layer0_outputs(4128) <= not(inputs(193));
    layer0_outputs(4129) <= (inputs(94)) or (inputs(91));
    layer0_outputs(4130) <= not(inputs(215)) or (inputs(84));
    layer0_outputs(4131) <= not(inputs(212)) or (inputs(28));
    layer0_outputs(4132) <= inputs(91);
    layer0_outputs(4133) <= (inputs(215)) or (inputs(158));
    layer0_outputs(4134) <= (inputs(207)) or (inputs(204));
    layer0_outputs(4135) <= not((inputs(32)) or (inputs(239)));
    layer0_outputs(4136) <= (inputs(244)) and not (inputs(31));
    layer0_outputs(4137) <= not((inputs(65)) or (inputs(213)));
    layer0_outputs(4138) <= not(inputs(205));
    layer0_outputs(4139) <= not(inputs(181));
    layer0_outputs(4140) <= (inputs(48)) and not (inputs(3));
    layer0_outputs(4141) <= not(inputs(38));
    layer0_outputs(4142) <= not(inputs(93));
    layer0_outputs(4143) <= (inputs(224)) or (inputs(254));
    layer0_outputs(4144) <= not(inputs(153));
    layer0_outputs(4145) <= inputs(231);
    layer0_outputs(4146) <= not((inputs(255)) or (inputs(221)));
    layer0_outputs(4147) <= (inputs(248)) and not (inputs(32));
    layer0_outputs(4148) <= (inputs(174)) xor (inputs(217));
    layer0_outputs(4149) <= (inputs(122)) or (inputs(223));
    layer0_outputs(4150) <= (inputs(232)) and not (inputs(110));
    layer0_outputs(4151) <= not(inputs(134));
    layer0_outputs(4152) <= (inputs(120)) and not (inputs(129));
    layer0_outputs(4153) <= (inputs(255)) xor (inputs(208));
    layer0_outputs(4154) <= not((inputs(172)) or (inputs(155)));
    layer0_outputs(4155) <= not(inputs(245));
    layer0_outputs(4156) <= not(inputs(165)) or (inputs(31));
    layer0_outputs(4157) <= '1';
    layer0_outputs(4158) <= not(inputs(26));
    layer0_outputs(4159) <= not((inputs(55)) xor (inputs(225)));
    layer0_outputs(4160) <= not(inputs(247));
    layer0_outputs(4161) <= not((inputs(51)) or (inputs(192)));
    layer0_outputs(4162) <= (inputs(63)) and not (inputs(220));
    layer0_outputs(4163) <= not(inputs(209));
    layer0_outputs(4164) <= not((inputs(249)) or (inputs(94)));
    layer0_outputs(4165) <= not((inputs(110)) xor (inputs(192)));
    layer0_outputs(4166) <= not((inputs(207)) or (inputs(75)));
    layer0_outputs(4167) <= (inputs(186)) and not (inputs(247));
    layer0_outputs(4168) <= not(inputs(98));
    layer0_outputs(4169) <= (inputs(103)) or (inputs(56));
    layer0_outputs(4170) <= not(inputs(99));
    layer0_outputs(4171) <= not(inputs(102)) or (inputs(50));
    layer0_outputs(4172) <= inputs(40);
    layer0_outputs(4173) <= (inputs(91)) xor (inputs(67));
    layer0_outputs(4174) <= '1';
    layer0_outputs(4175) <= not((inputs(245)) xor (inputs(195)));
    layer0_outputs(4176) <= not((inputs(14)) or (inputs(61)));
    layer0_outputs(4177) <= not(inputs(131));
    layer0_outputs(4178) <= (inputs(134)) and not (inputs(172));
    layer0_outputs(4179) <= (inputs(203)) xor (inputs(220));
    layer0_outputs(4180) <= not(inputs(232)) or (inputs(15));
    layer0_outputs(4181) <= (inputs(69)) and not (inputs(32));
    layer0_outputs(4182) <= inputs(225);
    layer0_outputs(4183) <= (inputs(175)) xor (inputs(147));
    layer0_outputs(4184) <= not(inputs(103)) or (inputs(206));
    layer0_outputs(4185) <= (inputs(58)) xor (inputs(119));
    layer0_outputs(4186) <= not(inputs(112));
    layer0_outputs(4187) <= (inputs(217)) or (inputs(203));
    layer0_outputs(4188) <= inputs(98);
    layer0_outputs(4189) <= inputs(116);
    layer0_outputs(4190) <= not((inputs(27)) and (inputs(25)));
    layer0_outputs(4191) <= not((inputs(213)) or (inputs(204)));
    layer0_outputs(4192) <= not((inputs(241)) xor (inputs(50)));
    layer0_outputs(4193) <= inputs(108);
    layer0_outputs(4194) <= not(inputs(70)) or (inputs(5));
    layer0_outputs(4195) <= (inputs(25)) and not (inputs(237));
    layer0_outputs(4196) <= not((inputs(90)) or (inputs(49)));
    layer0_outputs(4197) <= (inputs(171)) xor (inputs(20));
    layer0_outputs(4198) <= not(inputs(67));
    layer0_outputs(4199) <= not(inputs(182));
    layer0_outputs(4200) <= (inputs(149)) and not (inputs(253));
    layer0_outputs(4201) <= (inputs(66)) or (inputs(67));
    layer0_outputs(4202) <= not(inputs(74));
    layer0_outputs(4203) <= inputs(242);
    layer0_outputs(4204) <= not(inputs(213));
    layer0_outputs(4205) <= not((inputs(171)) or (inputs(176)));
    layer0_outputs(4206) <= not((inputs(148)) or (inputs(202)));
    layer0_outputs(4207) <= not((inputs(182)) or (inputs(149)));
    layer0_outputs(4208) <= not((inputs(236)) or (inputs(104)));
    layer0_outputs(4209) <= (inputs(84)) or (inputs(190));
    layer0_outputs(4210) <= not(inputs(26));
    layer0_outputs(4211) <= inputs(120);
    layer0_outputs(4212) <= not((inputs(102)) xor (inputs(154)));
    layer0_outputs(4213) <= inputs(149);
    layer0_outputs(4214) <= not((inputs(145)) or (inputs(51)));
    layer0_outputs(4215) <= (inputs(47)) xor (inputs(0));
    layer0_outputs(4216) <= not(inputs(230));
    layer0_outputs(4217) <= inputs(51);
    layer0_outputs(4218) <= (inputs(134)) xor (inputs(190));
    layer0_outputs(4219) <= (inputs(170)) xor (inputs(184));
    layer0_outputs(4220) <= not((inputs(25)) and (inputs(12)));
    layer0_outputs(4221) <= (inputs(166)) and not (inputs(78));
    layer0_outputs(4222) <= (inputs(53)) and not (inputs(172));
    layer0_outputs(4223) <= (inputs(162)) or (inputs(172));
    layer0_outputs(4224) <= not((inputs(71)) xor (inputs(42)));
    layer0_outputs(4225) <= not(inputs(167));
    layer0_outputs(4226) <= not(inputs(78));
    layer0_outputs(4227) <= not(inputs(210));
    layer0_outputs(4228) <= not((inputs(129)) xor (inputs(133)));
    layer0_outputs(4229) <= (inputs(221)) xor (inputs(236));
    layer0_outputs(4230) <= (inputs(152)) or (inputs(2));
    layer0_outputs(4231) <= not((inputs(189)) or (inputs(164)));
    layer0_outputs(4232) <= (inputs(213)) and not (inputs(17));
    layer0_outputs(4233) <= inputs(104);
    layer0_outputs(4234) <= not(inputs(245)) or (inputs(87));
    layer0_outputs(4235) <= not(inputs(45));
    layer0_outputs(4236) <= not(inputs(206)) or (inputs(128));
    layer0_outputs(4237) <= not(inputs(179));
    layer0_outputs(4238) <= '0';
    layer0_outputs(4239) <= (inputs(205)) and not (inputs(65));
    layer0_outputs(4240) <= not(inputs(52)) or (inputs(152));
    layer0_outputs(4241) <= inputs(153);
    layer0_outputs(4242) <= not((inputs(242)) or (inputs(207)));
    layer0_outputs(4243) <= not((inputs(245)) or (inputs(150)));
    layer0_outputs(4244) <= not(inputs(231)) or (inputs(3));
    layer0_outputs(4245) <= inputs(231);
    layer0_outputs(4246) <= not((inputs(26)) or (inputs(254)));
    layer0_outputs(4247) <= not(inputs(182));
    layer0_outputs(4248) <= not(inputs(85)) or (inputs(191));
    layer0_outputs(4249) <= (inputs(53)) or (inputs(141));
    layer0_outputs(4250) <= (inputs(119)) and not (inputs(35));
    layer0_outputs(4251) <= not((inputs(253)) or (inputs(230)));
    layer0_outputs(4252) <= not(inputs(213)) or (inputs(105));
    layer0_outputs(4253) <= not(inputs(104)) or (inputs(218));
    layer0_outputs(4254) <= inputs(130);
    layer0_outputs(4255) <= inputs(216);
    layer0_outputs(4256) <= (inputs(46)) xor (inputs(225));
    layer0_outputs(4257) <= (inputs(95)) xor (inputs(172));
    layer0_outputs(4258) <= not((inputs(171)) or (inputs(70)));
    layer0_outputs(4259) <= not(inputs(52));
    layer0_outputs(4260) <= (inputs(161)) xor (inputs(25));
    layer0_outputs(4261) <= (inputs(244)) or (inputs(176));
    layer0_outputs(4262) <= not((inputs(167)) or (inputs(103)));
    layer0_outputs(4263) <= (inputs(56)) or (inputs(220));
    layer0_outputs(4264) <= (inputs(58)) xor (inputs(88));
    layer0_outputs(4265) <= (inputs(199)) and not (inputs(81));
    layer0_outputs(4266) <= not(inputs(248));
    layer0_outputs(4267) <= (inputs(93)) xor (inputs(107));
    layer0_outputs(4268) <= (inputs(180)) and not (inputs(61));
    layer0_outputs(4269) <= not(inputs(183)) or (inputs(99));
    layer0_outputs(4270) <= (inputs(148)) xor (inputs(180));
    layer0_outputs(4271) <= not(inputs(21));
    layer0_outputs(4272) <= not(inputs(173)) or (inputs(149));
    layer0_outputs(4273) <= not(inputs(62));
    layer0_outputs(4274) <= (inputs(64)) and not (inputs(232));
    layer0_outputs(4275) <= not(inputs(22)) or (inputs(112));
    layer0_outputs(4276) <= (inputs(14)) and not (inputs(177));
    layer0_outputs(4277) <= inputs(71);
    layer0_outputs(4278) <= not(inputs(139)) or (inputs(123));
    layer0_outputs(4279) <= inputs(156);
    layer0_outputs(4280) <= (inputs(37)) and not (inputs(87));
    layer0_outputs(4281) <= (inputs(109)) or (inputs(9));
    layer0_outputs(4282) <= (inputs(166)) and not (inputs(97));
    layer0_outputs(4283) <= not((inputs(204)) or (inputs(82)));
    layer0_outputs(4284) <= inputs(84);
    layer0_outputs(4285) <= '1';
    layer0_outputs(4286) <= (inputs(193)) or (inputs(33));
    layer0_outputs(4287) <= not(inputs(109)) or (inputs(189));
    layer0_outputs(4288) <= not(inputs(178));
    layer0_outputs(4289) <= not(inputs(247));
    layer0_outputs(4290) <= not((inputs(82)) or (inputs(245)));
    layer0_outputs(4291) <= inputs(166);
    layer0_outputs(4292) <= (inputs(52)) and not (inputs(169));
    layer0_outputs(4293) <= inputs(101);
    layer0_outputs(4294) <= (inputs(210)) and not (inputs(219));
    layer0_outputs(4295) <= inputs(209);
    layer0_outputs(4296) <= (inputs(81)) and (inputs(51));
    layer0_outputs(4297) <= not(inputs(26));
    layer0_outputs(4298) <= (inputs(147)) and not (inputs(124));
    layer0_outputs(4299) <= (inputs(75)) xor (inputs(90));
    layer0_outputs(4300) <= not(inputs(183)) or (inputs(57));
    layer0_outputs(4301) <= (inputs(240)) xor (inputs(148));
    layer0_outputs(4302) <= not(inputs(147));
    layer0_outputs(4303) <= inputs(82);
    layer0_outputs(4304) <= inputs(118);
    layer0_outputs(4305) <= not((inputs(195)) xor (inputs(163)));
    layer0_outputs(4306) <= not(inputs(106)) or (inputs(128));
    layer0_outputs(4307) <= (inputs(45)) xor (inputs(75));
    layer0_outputs(4308) <= inputs(30);
    layer0_outputs(4309) <= inputs(184);
    layer0_outputs(4310) <= inputs(17);
    layer0_outputs(4311) <= '0';
    layer0_outputs(4312) <= not(inputs(198));
    layer0_outputs(4313) <= (inputs(14)) or (inputs(89));
    layer0_outputs(4314) <= not((inputs(189)) or (inputs(251)));
    layer0_outputs(4315) <= not((inputs(230)) xor (inputs(197)));
    layer0_outputs(4316) <= inputs(95);
    layer0_outputs(4317) <= inputs(122);
    layer0_outputs(4318) <= inputs(146);
    layer0_outputs(4319) <= (inputs(194)) and not (inputs(93));
    layer0_outputs(4320) <= not(inputs(175)) or (inputs(62));
    layer0_outputs(4321) <= not(inputs(210));
    layer0_outputs(4322) <= (inputs(167)) or (inputs(208));
    layer0_outputs(4323) <= not(inputs(77));
    layer0_outputs(4324) <= (inputs(60)) and not (inputs(202));
    layer0_outputs(4325) <= not(inputs(120));
    layer0_outputs(4326) <= not(inputs(215));
    layer0_outputs(4327) <= (inputs(63)) and not (inputs(253));
    layer0_outputs(4328) <= not(inputs(180));
    layer0_outputs(4329) <= (inputs(165)) and not (inputs(61));
    layer0_outputs(4330) <= not(inputs(117));
    layer0_outputs(4331) <= not((inputs(34)) or (inputs(102)));
    layer0_outputs(4332) <= (inputs(245)) xor (inputs(76));
    layer0_outputs(4333) <= not(inputs(26));
    layer0_outputs(4334) <= (inputs(61)) xor (inputs(246));
    layer0_outputs(4335) <= (inputs(158)) and not (inputs(12));
    layer0_outputs(4336) <= not(inputs(20)) or (inputs(161));
    layer0_outputs(4337) <= not(inputs(122)) or (inputs(81));
    layer0_outputs(4338) <= (inputs(154)) xor (inputs(68));
    layer0_outputs(4339) <= not((inputs(193)) or (inputs(244)));
    layer0_outputs(4340) <= not(inputs(29)) or (inputs(253));
    layer0_outputs(4341) <= (inputs(254)) or (inputs(137));
    layer0_outputs(4342) <= not(inputs(117));
    layer0_outputs(4343) <= not((inputs(6)) and (inputs(200)));
    layer0_outputs(4344) <= inputs(78);
    layer0_outputs(4345) <= (inputs(240)) and not (inputs(244));
    layer0_outputs(4346) <= (inputs(99)) or (inputs(238));
    layer0_outputs(4347) <= not((inputs(233)) xor (inputs(161)));
    layer0_outputs(4348) <= not(inputs(203)) or (inputs(158));
    layer0_outputs(4349) <= '0';
    layer0_outputs(4350) <= inputs(70);
    layer0_outputs(4351) <= not(inputs(19));
    layer0_outputs(4352) <= inputs(226);
    layer0_outputs(4353) <= not((inputs(11)) or (inputs(254)));
    layer0_outputs(4354) <= not(inputs(225));
    layer0_outputs(4355) <= not(inputs(119));
    layer0_outputs(4356) <= not(inputs(85)) or (inputs(243));
    layer0_outputs(4357) <= (inputs(174)) xor (inputs(206));
    layer0_outputs(4358) <= not((inputs(24)) or (inputs(254)));
    layer0_outputs(4359) <= (inputs(219)) and (inputs(248));
    layer0_outputs(4360) <= not(inputs(233)) or (inputs(16));
    layer0_outputs(4361) <= inputs(90);
    layer0_outputs(4362) <= inputs(130);
    layer0_outputs(4363) <= (inputs(135)) xor (inputs(210));
    layer0_outputs(4364) <= not(inputs(125)) or (inputs(253));
    layer0_outputs(4365) <= not(inputs(166));
    layer0_outputs(4366) <= not(inputs(235)) or (inputs(92));
    layer0_outputs(4367) <= inputs(147);
    layer0_outputs(4368) <= not(inputs(42));
    layer0_outputs(4369) <= not((inputs(191)) or (inputs(11)));
    layer0_outputs(4370) <= inputs(34);
    layer0_outputs(4371) <= (inputs(76)) and not (inputs(65));
    layer0_outputs(4372) <= not(inputs(157));
    layer0_outputs(4373) <= '0';
    layer0_outputs(4374) <= (inputs(131)) and not (inputs(58));
    layer0_outputs(4375) <= not(inputs(84)) or (inputs(228));
    layer0_outputs(4376) <= inputs(151);
    layer0_outputs(4377) <= not(inputs(165));
    layer0_outputs(4378) <= (inputs(227)) or (inputs(87));
    layer0_outputs(4379) <= (inputs(75)) or (inputs(16));
    layer0_outputs(4380) <= inputs(101);
    layer0_outputs(4381) <= inputs(75);
    layer0_outputs(4382) <= not(inputs(149));
    layer0_outputs(4383) <= (inputs(71)) or (inputs(253));
    layer0_outputs(4384) <= (inputs(74)) xor (inputs(72));
    layer0_outputs(4385) <= inputs(145);
    layer0_outputs(4386) <= (inputs(5)) and not (inputs(126));
    layer0_outputs(4387) <= inputs(214);
    layer0_outputs(4388) <= (inputs(91)) and (inputs(241));
    layer0_outputs(4389) <= inputs(165);
    layer0_outputs(4390) <= not((inputs(60)) or (inputs(8)));
    layer0_outputs(4391) <= not((inputs(98)) or (inputs(220)));
    layer0_outputs(4392) <= (inputs(227)) or (inputs(178));
    layer0_outputs(4393) <= (inputs(38)) xor (inputs(155));
    layer0_outputs(4394) <= (inputs(88)) and not (inputs(247));
    layer0_outputs(4395) <= (inputs(63)) or (inputs(66));
    layer0_outputs(4396) <= (inputs(54)) or (inputs(15));
    layer0_outputs(4397) <= not(inputs(209));
    layer0_outputs(4398) <= not((inputs(123)) xor (inputs(15)));
    layer0_outputs(4399) <= not((inputs(26)) or (inputs(41)));
    layer0_outputs(4400) <= (inputs(34)) xor (inputs(0));
    layer0_outputs(4401) <= not((inputs(6)) or (inputs(171)));
    layer0_outputs(4402) <= (inputs(204)) or (inputs(103));
    layer0_outputs(4403) <= (inputs(255)) and not (inputs(93));
    layer0_outputs(4404) <= (inputs(221)) or (inputs(208));
    layer0_outputs(4405) <= not(inputs(199)) or (inputs(31));
    layer0_outputs(4406) <= inputs(235);
    layer0_outputs(4407) <= inputs(92);
    layer0_outputs(4408) <= (inputs(89)) or (inputs(251));
    layer0_outputs(4409) <= (inputs(122)) and not (inputs(226));
    layer0_outputs(4410) <= not(inputs(35)) or (inputs(246));
    layer0_outputs(4411) <= not((inputs(119)) xor (inputs(147)));
    layer0_outputs(4412) <= not((inputs(222)) or (inputs(110)));
    layer0_outputs(4413) <= not(inputs(195));
    layer0_outputs(4414) <= not(inputs(25)) or (inputs(210));
    layer0_outputs(4415) <= '0';
    layer0_outputs(4416) <= inputs(95);
    layer0_outputs(4417) <= (inputs(80)) or (inputs(115));
    layer0_outputs(4418) <= (inputs(129)) or (inputs(179));
    layer0_outputs(4419) <= (inputs(184)) xor (inputs(212));
    layer0_outputs(4420) <= (inputs(219)) and not (inputs(31));
    layer0_outputs(4421) <= (inputs(9)) xor (inputs(174));
    layer0_outputs(4422) <= not((inputs(184)) or (inputs(18)));
    layer0_outputs(4423) <= not((inputs(79)) or (inputs(12)));
    layer0_outputs(4424) <= inputs(102);
    layer0_outputs(4425) <= (inputs(145)) xor (inputs(234));
    layer0_outputs(4426) <= (inputs(145)) xor (inputs(210));
    layer0_outputs(4427) <= not((inputs(190)) or (inputs(143)));
    layer0_outputs(4428) <= (inputs(177)) and not (inputs(47));
    layer0_outputs(4429) <= not((inputs(180)) and (inputs(180)));
    layer0_outputs(4430) <= inputs(144);
    layer0_outputs(4431) <= (inputs(20)) and not (inputs(96));
    layer0_outputs(4432) <= (inputs(159)) or (inputs(45));
    layer0_outputs(4433) <= (inputs(147)) xor (inputs(103));
    layer0_outputs(4434) <= not((inputs(199)) xor (inputs(12)));
    layer0_outputs(4435) <= not((inputs(92)) xor (inputs(43)));
    layer0_outputs(4436) <= inputs(205);
    layer0_outputs(4437) <= not((inputs(127)) or (inputs(149)));
    layer0_outputs(4438) <= (inputs(205)) and not (inputs(76));
    layer0_outputs(4439) <= inputs(179);
    layer0_outputs(4440) <= inputs(230);
    layer0_outputs(4441) <= not((inputs(233)) xor (inputs(143)));
    layer0_outputs(4442) <= not(inputs(85));
    layer0_outputs(4443) <= (inputs(204)) or (inputs(126));
    layer0_outputs(4444) <= not(inputs(75));
    layer0_outputs(4445) <= not(inputs(88)) or (inputs(208));
    layer0_outputs(4446) <= not((inputs(102)) or (inputs(150)));
    layer0_outputs(4447) <= (inputs(91)) and not (inputs(236));
    layer0_outputs(4448) <= not(inputs(21));
    layer0_outputs(4449) <= inputs(126);
    layer0_outputs(4450) <= not(inputs(122)) or (inputs(186));
    layer0_outputs(4451) <= not(inputs(200)) or (inputs(245));
    layer0_outputs(4452) <= (inputs(41)) or (inputs(63));
    layer0_outputs(4453) <= not(inputs(212)) or (inputs(12));
    layer0_outputs(4454) <= inputs(104);
    layer0_outputs(4455) <= not(inputs(161));
    layer0_outputs(4456) <= not(inputs(92)) or (inputs(138));
    layer0_outputs(4457) <= not(inputs(107));
    layer0_outputs(4458) <= not((inputs(47)) xor (inputs(44)));
    layer0_outputs(4459) <= (inputs(131)) and not (inputs(222));
    layer0_outputs(4460) <= (inputs(159)) and (inputs(187));
    layer0_outputs(4461) <= not((inputs(235)) and (inputs(177)));
    layer0_outputs(4462) <= not((inputs(175)) or (inputs(207)));
    layer0_outputs(4463) <= (inputs(246)) or (inputs(215));
    layer0_outputs(4464) <= not(inputs(233));
    layer0_outputs(4465) <= not(inputs(89)) or (inputs(251));
    layer0_outputs(4466) <= not(inputs(150)) or (inputs(234));
    layer0_outputs(4467) <= (inputs(247)) or (inputs(128));
    layer0_outputs(4468) <= not(inputs(235));
    layer0_outputs(4469) <= not((inputs(213)) xor (inputs(253)));
    layer0_outputs(4470) <= (inputs(210)) or (inputs(25));
    layer0_outputs(4471) <= not(inputs(230));
    layer0_outputs(4472) <= (inputs(79)) or (inputs(171));
    layer0_outputs(4473) <= not((inputs(8)) xor (inputs(67)));
    layer0_outputs(4474) <= inputs(38);
    layer0_outputs(4475) <= not(inputs(246));
    layer0_outputs(4476) <= (inputs(121)) and not (inputs(114));
    layer0_outputs(4477) <= not(inputs(22));
    layer0_outputs(4478) <= not(inputs(117));
    layer0_outputs(4479) <= not((inputs(195)) or (inputs(129)));
    layer0_outputs(4480) <= not(inputs(121));
    layer0_outputs(4481) <= not(inputs(110));
    layer0_outputs(4482) <= not(inputs(172));
    layer0_outputs(4483) <= not(inputs(127));
    layer0_outputs(4484) <= not(inputs(55));
    layer0_outputs(4485) <= (inputs(223)) and not (inputs(45));
    layer0_outputs(4486) <= not((inputs(93)) and (inputs(169)));
    layer0_outputs(4487) <= not(inputs(124)) or (inputs(123));
    layer0_outputs(4488) <= not((inputs(143)) or (inputs(185)));
    layer0_outputs(4489) <= (inputs(70)) xor (inputs(21));
    layer0_outputs(4490) <= (inputs(166)) xor (inputs(253));
    layer0_outputs(4491) <= (inputs(201)) and not (inputs(131));
    layer0_outputs(4492) <= not((inputs(247)) xor (inputs(81)));
    layer0_outputs(4493) <= (inputs(232)) and not (inputs(93));
    layer0_outputs(4494) <= not((inputs(106)) xor (inputs(158)));
    layer0_outputs(4495) <= (inputs(57)) or (inputs(95));
    layer0_outputs(4496) <= (inputs(129)) or (inputs(214));
    layer0_outputs(4497) <= not(inputs(41));
    layer0_outputs(4498) <= (inputs(215)) or (inputs(216));
    layer0_outputs(4499) <= inputs(96);
    layer0_outputs(4500) <= (inputs(213)) and not (inputs(158));
    layer0_outputs(4501) <= (inputs(235)) xor (inputs(79));
    layer0_outputs(4502) <= not(inputs(194));
    layer0_outputs(4503) <= not(inputs(50));
    layer0_outputs(4504) <= not((inputs(33)) or (inputs(8)));
    layer0_outputs(4505) <= (inputs(69)) or (inputs(83));
    layer0_outputs(4506) <= not(inputs(233));
    layer0_outputs(4507) <= inputs(42);
    layer0_outputs(4508) <= not((inputs(79)) or (inputs(90)));
    layer0_outputs(4509) <= (inputs(45)) or (inputs(55));
    layer0_outputs(4510) <= (inputs(86)) xor (inputs(93));
    layer0_outputs(4511) <= not((inputs(234)) xor (inputs(121)));
    layer0_outputs(4512) <= '1';
    layer0_outputs(4513) <= (inputs(183)) or (inputs(230));
    layer0_outputs(4514) <= inputs(223);
    layer0_outputs(4515) <= not((inputs(147)) and (inputs(133)));
    layer0_outputs(4516) <= not((inputs(69)) or (inputs(197)));
    layer0_outputs(4517) <= (inputs(127)) and (inputs(225));
    layer0_outputs(4518) <= not((inputs(87)) or (inputs(31)));
    layer0_outputs(4519) <= not(inputs(43));
    layer0_outputs(4520) <= not((inputs(225)) or (inputs(232)));
    layer0_outputs(4521) <= not((inputs(223)) or (inputs(233)));
    layer0_outputs(4522) <= not(inputs(135));
    layer0_outputs(4523) <= inputs(185);
    layer0_outputs(4524) <= (inputs(202)) and not (inputs(128));
    layer0_outputs(4525) <= not(inputs(134));
    layer0_outputs(4526) <= (inputs(86)) or (inputs(209));
    layer0_outputs(4527) <= not(inputs(193));
    layer0_outputs(4528) <= not(inputs(75)) or (inputs(254));
    layer0_outputs(4529) <= not((inputs(18)) or (inputs(10)));
    layer0_outputs(4530) <= not(inputs(117)) or (inputs(187));
    layer0_outputs(4531) <= not((inputs(18)) or (inputs(162)));
    layer0_outputs(4532) <= '0';
    layer0_outputs(4533) <= inputs(228);
    layer0_outputs(4534) <= not(inputs(20)) or (inputs(77));
    layer0_outputs(4535) <= not(inputs(201));
    layer0_outputs(4536) <= not(inputs(235));
    layer0_outputs(4537) <= not((inputs(67)) or (inputs(164)));
    layer0_outputs(4538) <= inputs(8);
    layer0_outputs(4539) <= inputs(187);
    layer0_outputs(4540) <= inputs(88);
    layer0_outputs(4541) <= (inputs(67)) xor (inputs(109));
    layer0_outputs(4542) <= (inputs(143)) or (inputs(162));
    layer0_outputs(4543) <= not((inputs(26)) or (inputs(254)));
    layer0_outputs(4544) <= not(inputs(119));
    layer0_outputs(4545) <= (inputs(96)) or (inputs(202));
    layer0_outputs(4546) <= (inputs(174)) and not (inputs(146));
    layer0_outputs(4547) <= not((inputs(10)) xor (inputs(45)));
    layer0_outputs(4548) <= not(inputs(48));
    layer0_outputs(4549) <= not(inputs(122)) or (inputs(83));
    layer0_outputs(4550) <= not(inputs(46));
    layer0_outputs(4551) <= not(inputs(247));
    layer0_outputs(4552) <= not(inputs(14));
    layer0_outputs(4553) <= not(inputs(132));
    layer0_outputs(4554) <= (inputs(195)) and (inputs(61));
    layer0_outputs(4555) <= inputs(95);
    layer0_outputs(4556) <= (inputs(135)) and not (inputs(114));
    layer0_outputs(4557) <= not(inputs(155)) or (inputs(2));
    layer0_outputs(4558) <= not((inputs(242)) or (inputs(207)));
    layer0_outputs(4559) <= not((inputs(44)) xor (inputs(20)));
    layer0_outputs(4560) <= not(inputs(225)) or (inputs(252));
    layer0_outputs(4561) <= not(inputs(41)) or (inputs(183));
    layer0_outputs(4562) <= (inputs(209)) or (inputs(122));
    layer0_outputs(4563) <= not((inputs(252)) and (inputs(13)));
    layer0_outputs(4564) <= inputs(178);
    layer0_outputs(4565) <= not(inputs(125)) or (inputs(32));
    layer0_outputs(4566) <= not(inputs(68));
    layer0_outputs(4567) <= inputs(26);
    layer0_outputs(4568) <= not((inputs(36)) or (inputs(142)));
    layer0_outputs(4569) <= (inputs(60)) and not (inputs(223));
    layer0_outputs(4570) <= not(inputs(141));
    layer0_outputs(4571) <= not(inputs(104));
    layer0_outputs(4572) <= (inputs(47)) or (inputs(235));
    layer0_outputs(4573) <= not(inputs(234)) or (inputs(95));
    layer0_outputs(4574) <= not(inputs(121));
    layer0_outputs(4575) <= (inputs(49)) or (inputs(226));
    layer0_outputs(4576) <= inputs(204);
    layer0_outputs(4577) <= (inputs(197)) and not (inputs(62));
    layer0_outputs(4578) <= (inputs(176)) xor (inputs(117));
    layer0_outputs(4579) <= (inputs(176)) or (inputs(158));
    layer0_outputs(4580) <= not(inputs(216)) or (inputs(60));
    layer0_outputs(4581) <= not(inputs(95));
    layer0_outputs(4582) <= not((inputs(245)) or (inputs(204)));
    layer0_outputs(4583) <= inputs(23);
    layer0_outputs(4584) <= not((inputs(156)) and (inputs(95)));
    layer0_outputs(4585) <= (inputs(34)) and not (inputs(238));
    layer0_outputs(4586) <= inputs(25);
    layer0_outputs(4587) <= (inputs(130)) xor (inputs(133));
    layer0_outputs(4588) <= not((inputs(144)) or (inputs(88)));
    layer0_outputs(4589) <= (inputs(126)) xor (inputs(206));
    layer0_outputs(4590) <= inputs(173);
    layer0_outputs(4591) <= not((inputs(161)) or (inputs(221)));
    layer0_outputs(4592) <= not(inputs(97));
    layer0_outputs(4593) <= (inputs(56)) and not (inputs(199));
    layer0_outputs(4594) <= (inputs(152)) and not (inputs(16));
    layer0_outputs(4595) <= not(inputs(26));
    layer0_outputs(4596) <= (inputs(108)) xor (inputs(42));
    layer0_outputs(4597) <= not((inputs(111)) or (inputs(182)));
    layer0_outputs(4598) <= not((inputs(109)) xor (inputs(65)));
    layer0_outputs(4599) <= (inputs(119)) and not (inputs(191));
    layer0_outputs(4600) <= not((inputs(128)) xor (inputs(153)));
    layer0_outputs(4601) <= not(inputs(228)) or (inputs(31));
    layer0_outputs(4602) <= not((inputs(150)) and (inputs(118)));
    layer0_outputs(4603) <= not((inputs(105)) xor (inputs(158)));
    layer0_outputs(4604) <= not(inputs(134)) or (inputs(157));
    layer0_outputs(4605) <= (inputs(84)) and not (inputs(73));
    layer0_outputs(4606) <= (inputs(81)) or (inputs(20));
    layer0_outputs(4607) <= (inputs(110)) xor (inputs(37));
    layer0_outputs(4608) <= not(inputs(153));
    layer0_outputs(4609) <= inputs(222);
    layer0_outputs(4610) <= inputs(108);
    layer0_outputs(4611) <= inputs(227);
    layer0_outputs(4612) <= (inputs(165)) and not (inputs(170));
    layer0_outputs(4613) <= not(inputs(58)) or (inputs(203));
    layer0_outputs(4614) <= not((inputs(135)) or (inputs(241)));
    layer0_outputs(4615) <= not(inputs(166));
    layer0_outputs(4616) <= not((inputs(24)) or (inputs(106)));
    layer0_outputs(4617) <= inputs(27);
    layer0_outputs(4618) <= '1';
    layer0_outputs(4619) <= inputs(246);
    layer0_outputs(4620) <= inputs(221);
    layer0_outputs(4621) <= inputs(162);
    layer0_outputs(4622) <= not(inputs(145));
    layer0_outputs(4623) <= not((inputs(52)) xor (inputs(54)));
    layer0_outputs(4624) <= inputs(233);
    layer0_outputs(4625) <= (inputs(231)) xor (inputs(183));
    layer0_outputs(4626) <= (inputs(92)) or (inputs(167));
    layer0_outputs(4627) <= inputs(106);
    layer0_outputs(4628) <= inputs(116);
    layer0_outputs(4629) <= (inputs(154)) or (inputs(162));
    layer0_outputs(4630) <= inputs(162);
    layer0_outputs(4631) <= (inputs(109)) or (inputs(31));
    layer0_outputs(4632) <= not(inputs(9));
    layer0_outputs(4633) <= not((inputs(231)) and (inputs(213)));
    layer0_outputs(4634) <= inputs(134);
    layer0_outputs(4635) <= not(inputs(181));
    layer0_outputs(4636) <= '0';
    layer0_outputs(4637) <= (inputs(15)) or (inputs(45));
    layer0_outputs(4638) <= (inputs(157)) or (inputs(202));
    layer0_outputs(4639) <= not(inputs(105)) or (inputs(13));
    layer0_outputs(4640) <= not(inputs(162)) or (inputs(254));
    layer0_outputs(4641) <= (inputs(23)) and not (inputs(208));
    layer0_outputs(4642) <= not(inputs(221));
    layer0_outputs(4643) <= not((inputs(254)) or (inputs(238)));
    layer0_outputs(4644) <= inputs(214);
    layer0_outputs(4645) <= (inputs(150)) and (inputs(104));
    layer0_outputs(4646) <= inputs(231);
    layer0_outputs(4647) <= not(inputs(229));
    layer0_outputs(4648) <= not((inputs(188)) xor (inputs(65)));
    layer0_outputs(4649) <= inputs(123);
    layer0_outputs(4650) <= (inputs(106)) and not (inputs(200));
    layer0_outputs(4651) <= (inputs(138)) xor (inputs(182));
    layer0_outputs(4652) <= not((inputs(26)) or (inputs(1)));
    layer0_outputs(4653) <= (inputs(173)) and not (inputs(177));
    layer0_outputs(4654) <= (inputs(35)) and not (inputs(12));
    layer0_outputs(4655) <= not((inputs(81)) or (inputs(249)));
    layer0_outputs(4656) <= (inputs(229)) and not (inputs(18));
    layer0_outputs(4657) <= (inputs(95)) xor (inputs(91));
    layer0_outputs(4658) <= not(inputs(102));
    layer0_outputs(4659) <= not(inputs(125));
    layer0_outputs(4660) <= not(inputs(110)) or (inputs(210));
    layer0_outputs(4661) <= not(inputs(220)) or (inputs(234));
    layer0_outputs(4662) <= (inputs(100)) xor (inputs(96));
    layer0_outputs(4663) <= '0';
    layer0_outputs(4664) <= (inputs(249)) or (inputs(93));
    layer0_outputs(4665) <= (inputs(232)) and not (inputs(102));
    layer0_outputs(4666) <= inputs(109);
    layer0_outputs(4667) <= not((inputs(163)) or (inputs(211)));
    layer0_outputs(4668) <= inputs(99);
    layer0_outputs(4669) <= (inputs(61)) xor (inputs(105));
    layer0_outputs(4670) <= (inputs(14)) and (inputs(125));
    layer0_outputs(4671) <= (inputs(47)) xor (inputs(80));
    layer0_outputs(4672) <= not(inputs(32));
    layer0_outputs(4673) <= not(inputs(176)) or (inputs(205));
    layer0_outputs(4674) <= not(inputs(226)) or (inputs(223));
    layer0_outputs(4675) <= (inputs(140)) or (inputs(140));
    layer0_outputs(4676) <= inputs(62);
    layer0_outputs(4677) <= not((inputs(107)) or (inputs(130)));
    layer0_outputs(4678) <= (inputs(161)) or (inputs(189));
    layer0_outputs(4679) <= not((inputs(43)) xor (inputs(42)));
    layer0_outputs(4680) <= inputs(165);
    layer0_outputs(4681) <= (inputs(212)) or (inputs(71));
    layer0_outputs(4682) <= (inputs(7)) or (inputs(96));
    layer0_outputs(4683) <= (inputs(66)) xor (inputs(85));
    layer0_outputs(4684) <= inputs(17);
    layer0_outputs(4685) <= (inputs(52)) xor (inputs(56));
    layer0_outputs(4686) <= inputs(113);
    layer0_outputs(4687) <= not(inputs(45)) or (inputs(242));
    layer0_outputs(4688) <= not(inputs(119)) or (inputs(142));
    layer0_outputs(4689) <= not(inputs(190));
    layer0_outputs(4690) <= (inputs(232)) and not (inputs(239));
    layer0_outputs(4691) <= not(inputs(121)) or (inputs(72));
    layer0_outputs(4692) <= (inputs(251)) or (inputs(192));
    layer0_outputs(4693) <= (inputs(154)) or (inputs(208));
    layer0_outputs(4694) <= (inputs(168)) and not (inputs(42));
    layer0_outputs(4695) <= (inputs(54)) and not (inputs(93));
    layer0_outputs(4696) <= inputs(207);
    layer0_outputs(4697) <= (inputs(102)) and not (inputs(226));
    layer0_outputs(4698) <= not(inputs(230)) or (inputs(162));
    layer0_outputs(4699) <= inputs(23);
    layer0_outputs(4700) <= (inputs(117)) or (inputs(250));
    layer0_outputs(4701) <= not((inputs(219)) and (inputs(197)));
    layer0_outputs(4702) <= not((inputs(220)) or (inputs(198)));
    layer0_outputs(4703) <= inputs(211);
    layer0_outputs(4704) <= (inputs(113)) and (inputs(44));
    layer0_outputs(4705) <= (inputs(49)) or (inputs(200));
    layer0_outputs(4706) <= not((inputs(144)) or (inputs(53)));
    layer0_outputs(4707) <= '0';
    layer0_outputs(4708) <= not((inputs(87)) or (inputs(241)));
    layer0_outputs(4709) <= (inputs(254)) or (inputs(144));
    layer0_outputs(4710) <= inputs(23);
    layer0_outputs(4711) <= (inputs(122)) and (inputs(62));
    layer0_outputs(4712) <= not((inputs(226)) xor (inputs(149)));
    layer0_outputs(4713) <= not(inputs(193));
    layer0_outputs(4714) <= not(inputs(40)) or (inputs(175));
    layer0_outputs(4715) <= not((inputs(199)) and (inputs(214)));
    layer0_outputs(4716) <= inputs(136);
    layer0_outputs(4717) <= inputs(186);
    layer0_outputs(4718) <= (inputs(19)) and not (inputs(33));
    layer0_outputs(4719) <= not(inputs(67)) or (inputs(127));
    layer0_outputs(4720) <= (inputs(74)) and not (inputs(111));
    layer0_outputs(4721) <= not((inputs(125)) xor (inputs(159)));
    layer0_outputs(4722) <= not((inputs(116)) or (inputs(85)));
    layer0_outputs(4723) <= not((inputs(203)) xor (inputs(81)));
    layer0_outputs(4724) <= not((inputs(156)) or (inputs(67)));
    layer0_outputs(4725) <= not(inputs(73)) or (inputs(92));
    layer0_outputs(4726) <= (inputs(173)) xor (inputs(124));
    layer0_outputs(4727) <= inputs(90);
    layer0_outputs(4728) <= not(inputs(214)) or (inputs(82));
    layer0_outputs(4729) <= not(inputs(150));
    layer0_outputs(4730) <= not((inputs(75)) or (inputs(124)));
    layer0_outputs(4731) <= not(inputs(113)) or (inputs(95));
    layer0_outputs(4732) <= not(inputs(204)) or (inputs(3));
    layer0_outputs(4733) <= '0';
    layer0_outputs(4734) <= not((inputs(6)) or (inputs(3)));
    layer0_outputs(4735) <= not((inputs(54)) xor (inputs(102)));
    layer0_outputs(4736) <= '0';
    layer0_outputs(4737) <= not((inputs(80)) or (inputs(234)));
    layer0_outputs(4738) <= not(inputs(77));
    layer0_outputs(4739) <= not(inputs(114));
    layer0_outputs(4740) <= inputs(95);
    layer0_outputs(4741) <= '1';
    layer0_outputs(4742) <= not(inputs(194));
    layer0_outputs(4743) <= not((inputs(120)) or (inputs(134)));
    layer0_outputs(4744) <= not(inputs(239));
    layer0_outputs(4745) <= not(inputs(241));
    layer0_outputs(4746) <= (inputs(138)) or (inputs(128));
    layer0_outputs(4747) <= not(inputs(152)) or (inputs(123));
    layer0_outputs(4748) <= inputs(161);
    layer0_outputs(4749) <= (inputs(186)) or (inputs(196));
    layer0_outputs(4750) <= (inputs(69)) and not (inputs(158));
    layer0_outputs(4751) <= not((inputs(148)) xor (inputs(101)));
    layer0_outputs(4752) <= inputs(90);
    layer0_outputs(4753) <= not(inputs(199)) or (inputs(99));
    layer0_outputs(4754) <= inputs(94);
    layer0_outputs(4755) <= not((inputs(177)) xor (inputs(25)));
    layer0_outputs(4756) <= (inputs(219)) or (inputs(36));
    layer0_outputs(4757) <= not(inputs(25));
    layer0_outputs(4758) <= not((inputs(255)) or (inputs(173)));
    layer0_outputs(4759) <= not((inputs(209)) xor (inputs(218)));
    layer0_outputs(4760) <= inputs(138);
    layer0_outputs(4761) <= inputs(187);
    layer0_outputs(4762) <= not((inputs(143)) xor (inputs(92)));
    layer0_outputs(4763) <= inputs(166);
    layer0_outputs(4764) <= (inputs(7)) or (inputs(10));
    layer0_outputs(4765) <= (inputs(218)) and not (inputs(98));
    layer0_outputs(4766) <= not(inputs(189)) or (inputs(146));
    layer0_outputs(4767) <= (inputs(85)) and not (inputs(32));
    layer0_outputs(4768) <= (inputs(64)) or (inputs(116));
    layer0_outputs(4769) <= not(inputs(240));
    layer0_outputs(4770) <= not(inputs(208)) or (inputs(103));
    layer0_outputs(4771) <= not(inputs(199)) or (inputs(77));
    layer0_outputs(4772) <= not((inputs(104)) xor (inputs(129)));
    layer0_outputs(4773) <= not(inputs(243)) or (inputs(31));
    layer0_outputs(4774) <= inputs(160);
    layer0_outputs(4775) <= not(inputs(29));
    layer0_outputs(4776) <= not((inputs(152)) or (inputs(139)));
    layer0_outputs(4777) <= inputs(203);
    layer0_outputs(4778) <= not((inputs(69)) xor (inputs(236)));
    layer0_outputs(4779) <= not((inputs(181)) or (inputs(0)));
    layer0_outputs(4780) <= inputs(76);
    layer0_outputs(4781) <= inputs(147);
    layer0_outputs(4782) <= (inputs(252)) xor (inputs(80));
    layer0_outputs(4783) <= (inputs(195)) xor (inputs(229));
    layer0_outputs(4784) <= inputs(97);
    layer0_outputs(4785) <= '1';
    layer0_outputs(4786) <= (inputs(240)) xor (inputs(72));
    layer0_outputs(4787) <= not(inputs(119)) or (inputs(111));
    layer0_outputs(4788) <= '1';
    layer0_outputs(4789) <= (inputs(132)) xor (inputs(66));
    layer0_outputs(4790) <= not((inputs(145)) or (inputs(181)));
    layer0_outputs(4791) <= not((inputs(186)) or (inputs(108)));
    layer0_outputs(4792) <= not((inputs(199)) and (inputs(218)));
    layer0_outputs(4793) <= not((inputs(196)) or (inputs(246)));
    layer0_outputs(4794) <= inputs(134);
    layer0_outputs(4795) <= (inputs(205)) xor (inputs(52));
    layer0_outputs(4796) <= not((inputs(158)) or (inputs(236)));
    layer0_outputs(4797) <= not(inputs(198)) or (inputs(93));
    layer0_outputs(4798) <= not(inputs(131));
    layer0_outputs(4799) <= (inputs(19)) or (inputs(210));
    layer0_outputs(4800) <= (inputs(27)) or (inputs(246));
    layer0_outputs(4801) <= not(inputs(199));
    layer0_outputs(4802) <= inputs(9);
    layer0_outputs(4803) <= not((inputs(123)) or (inputs(112)));
    layer0_outputs(4804) <= not(inputs(82));
    layer0_outputs(4805) <= not((inputs(245)) or (inputs(6)));
    layer0_outputs(4806) <= inputs(77);
    layer0_outputs(4807) <= (inputs(133)) xor (inputs(156));
    layer0_outputs(4808) <= not((inputs(48)) xor (inputs(251)));
    layer0_outputs(4809) <= not((inputs(227)) xor (inputs(207)));
    layer0_outputs(4810) <= (inputs(41)) or (inputs(37));
    layer0_outputs(4811) <= not((inputs(239)) or (inputs(238)));
    layer0_outputs(4812) <= '1';
    layer0_outputs(4813) <= not(inputs(69));
    layer0_outputs(4814) <= not((inputs(102)) xor (inputs(179)));
    layer0_outputs(4815) <= not(inputs(131)) or (inputs(89));
    layer0_outputs(4816) <= inputs(75);
    layer0_outputs(4817) <= '1';
    layer0_outputs(4818) <= (inputs(217)) or (inputs(255));
    layer0_outputs(4819) <= not((inputs(132)) xor (inputs(136)));
    layer0_outputs(4820) <= not((inputs(194)) xor (inputs(67)));
    layer0_outputs(4821) <= not((inputs(95)) or (inputs(8)));
    layer0_outputs(4822) <= inputs(126);
    layer0_outputs(4823) <= not(inputs(169)) or (inputs(36));
    layer0_outputs(4824) <= (inputs(134)) xor (inputs(119));
    layer0_outputs(4825) <= not(inputs(99));
    layer0_outputs(4826) <= inputs(152);
    layer0_outputs(4827) <= not((inputs(142)) xor (inputs(163)));
    layer0_outputs(4828) <= not(inputs(90)) or (inputs(11));
    layer0_outputs(4829) <= not(inputs(149));
    layer0_outputs(4830) <= (inputs(229)) and not (inputs(82));
    layer0_outputs(4831) <= inputs(178);
    layer0_outputs(4832) <= not((inputs(177)) or (inputs(204)));
    layer0_outputs(4833) <= (inputs(251)) or (inputs(87));
    layer0_outputs(4834) <= not((inputs(242)) or (inputs(32)));
    layer0_outputs(4835) <= (inputs(193)) xor (inputs(12));
    layer0_outputs(4836) <= not((inputs(191)) or (inputs(245)));
    layer0_outputs(4837) <= not((inputs(32)) xor (inputs(47)));
    layer0_outputs(4838) <= not(inputs(53));
    layer0_outputs(4839) <= not(inputs(90));
    layer0_outputs(4840) <= not(inputs(124));
    layer0_outputs(4841) <= not(inputs(178)) or (inputs(30));
    layer0_outputs(4842) <= inputs(156);
    layer0_outputs(4843) <= not((inputs(225)) or (inputs(57)));
    layer0_outputs(4844) <= not(inputs(24)) or (inputs(166));
    layer0_outputs(4845) <= not((inputs(142)) or (inputs(71)));
    layer0_outputs(4846) <= not(inputs(162));
    layer0_outputs(4847) <= not((inputs(128)) or (inputs(234)));
    layer0_outputs(4848) <= not(inputs(168));
    layer0_outputs(4849) <= inputs(38);
    layer0_outputs(4850) <= inputs(117);
    layer0_outputs(4851) <= '0';
    layer0_outputs(4852) <= not((inputs(62)) or (inputs(191)));
    layer0_outputs(4853) <= (inputs(101)) xor (inputs(154));
    layer0_outputs(4854) <= not((inputs(7)) or (inputs(19)));
    layer0_outputs(4855) <= inputs(34);
    layer0_outputs(4856) <= not(inputs(253));
    layer0_outputs(4857) <= not(inputs(212)) or (inputs(78));
    layer0_outputs(4858) <= (inputs(144)) or (inputs(173));
    layer0_outputs(4859) <= not(inputs(144));
    layer0_outputs(4860) <= (inputs(253)) xor (inputs(133));
    layer0_outputs(4861) <= not((inputs(136)) xor (inputs(168)));
    layer0_outputs(4862) <= not((inputs(79)) xor (inputs(159)));
    layer0_outputs(4863) <= inputs(66);
    layer0_outputs(4864) <= not(inputs(7)) or (inputs(147));
    layer0_outputs(4865) <= not(inputs(106));
    layer0_outputs(4866) <= not(inputs(137));
    layer0_outputs(4867) <= inputs(50);
    layer0_outputs(4868) <= not((inputs(245)) or (inputs(208)));
    layer0_outputs(4869) <= (inputs(255)) or (inputs(205));
    layer0_outputs(4870) <= (inputs(71)) and not (inputs(157));
    layer0_outputs(4871) <= not((inputs(148)) xor (inputs(210)));
    layer0_outputs(4872) <= not((inputs(59)) or (inputs(242)));
    layer0_outputs(4873) <= (inputs(29)) or (inputs(133));
    layer0_outputs(4874) <= (inputs(194)) xor (inputs(235));
    layer0_outputs(4875) <= inputs(165);
    layer0_outputs(4876) <= not(inputs(51));
    layer0_outputs(4877) <= not((inputs(173)) xor (inputs(143)));
    layer0_outputs(4878) <= inputs(229);
    layer0_outputs(4879) <= not(inputs(44));
    layer0_outputs(4880) <= (inputs(88)) or (inputs(142));
    layer0_outputs(4881) <= not((inputs(178)) xor (inputs(237)));
    layer0_outputs(4882) <= (inputs(151)) and not (inputs(17));
    layer0_outputs(4883) <= (inputs(44)) xor (inputs(143));
    layer0_outputs(4884) <= not((inputs(170)) or (inputs(222)));
    layer0_outputs(4885) <= not(inputs(83));
    layer0_outputs(4886) <= not(inputs(100)) or (inputs(4));
    layer0_outputs(4887) <= (inputs(115)) and not (inputs(57));
    layer0_outputs(4888) <= inputs(30);
    layer0_outputs(4889) <= inputs(23);
    layer0_outputs(4890) <= (inputs(194)) and not (inputs(1));
    layer0_outputs(4891) <= inputs(222);
    layer0_outputs(4892) <= not(inputs(74)) or (inputs(53));
    layer0_outputs(4893) <= not(inputs(68));
    layer0_outputs(4894) <= '0';
    layer0_outputs(4895) <= not(inputs(233));
    layer0_outputs(4896) <= (inputs(122)) and not (inputs(32));
    layer0_outputs(4897) <= not((inputs(99)) or (inputs(81)));
    layer0_outputs(4898) <= '1';
    layer0_outputs(4899) <= (inputs(217)) or (inputs(143));
    layer0_outputs(4900) <= (inputs(39)) and not (inputs(252));
    layer0_outputs(4901) <= (inputs(22)) and not (inputs(130));
    layer0_outputs(4902) <= inputs(76);
    layer0_outputs(4903) <= inputs(199);
    layer0_outputs(4904) <= (inputs(154)) and (inputs(183));
    layer0_outputs(4905) <= not((inputs(220)) or (inputs(21)));
    layer0_outputs(4906) <= (inputs(211)) xor (inputs(249));
    layer0_outputs(4907) <= inputs(164);
    layer0_outputs(4908) <= not(inputs(103)) or (inputs(18));
    layer0_outputs(4909) <= not((inputs(38)) or (inputs(39)));
    layer0_outputs(4910) <= inputs(59);
    layer0_outputs(4911) <= inputs(164);
    layer0_outputs(4912) <= inputs(90);
    layer0_outputs(4913) <= (inputs(174)) or (inputs(116));
    layer0_outputs(4914) <= not(inputs(252));
    layer0_outputs(4915) <= (inputs(144)) xor (inputs(136));
    layer0_outputs(4916) <= inputs(114);
    layer0_outputs(4917) <= (inputs(110)) or (inputs(69));
    layer0_outputs(4918) <= not((inputs(175)) or (inputs(88)));
    layer0_outputs(4919) <= inputs(146);
    layer0_outputs(4920) <= inputs(115);
    layer0_outputs(4921) <= (inputs(132)) or (inputs(4));
    layer0_outputs(4922) <= not(inputs(4)) or (inputs(158));
    layer0_outputs(4923) <= not(inputs(183));
    layer0_outputs(4924) <= not(inputs(173)) or (inputs(24));
    layer0_outputs(4925) <= not(inputs(87)) or (inputs(77));
    layer0_outputs(4926) <= not(inputs(204)) or (inputs(29));
    layer0_outputs(4927) <= inputs(185);
    layer0_outputs(4928) <= inputs(232);
    layer0_outputs(4929) <= not((inputs(242)) or (inputs(223)));
    layer0_outputs(4930) <= (inputs(7)) and not (inputs(97));
    layer0_outputs(4931) <= not((inputs(227)) and (inputs(231)));
    layer0_outputs(4932) <= inputs(99);
    layer0_outputs(4933) <= (inputs(23)) xor (inputs(69));
    layer0_outputs(4934) <= not((inputs(106)) or (inputs(45)));
    layer0_outputs(4935) <= not(inputs(105));
    layer0_outputs(4936) <= not((inputs(118)) xor (inputs(145)));
    layer0_outputs(4937) <= not(inputs(161));
    layer0_outputs(4938) <= '0';
    layer0_outputs(4939) <= (inputs(91)) and not (inputs(162));
    layer0_outputs(4940) <= inputs(25);
    layer0_outputs(4941) <= not((inputs(39)) or (inputs(92)));
    layer0_outputs(4942) <= (inputs(198)) and (inputs(206));
    layer0_outputs(4943) <= inputs(155);
    layer0_outputs(4944) <= inputs(58);
    layer0_outputs(4945) <= not(inputs(247));
    layer0_outputs(4946) <= not(inputs(10));
    layer0_outputs(4947) <= not(inputs(147));
    layer0_outputs(4948) <= '1';
    layer0_outputs(4949) <= inputs(11);
    layer0_outputs(4950) <= (inputs(77)) or (inputs(4));
    layer0_outputs(4951) <= (inputs(229)) xor (inputs(40));
    layer0_outputs(4952) <= not(inputs(220)) or (inputs(130));
    layer0_outputs(4953) <= not((inputs(80)) xor (inputs(183)));
    layer0_outputs(4954) <= not((inputs(184)) xor (inputs(191)));
    layer0_outputs(4955) <= (inputs(179)) or (inputs(200));
    layer0_outputs(4956) <= not((inputs(45)) or (inputs(31)));
    layer0_outputs(4957) <= not((inputs(177)) or (inputs(62)));
    layer0_outputs(4958) <= not(inputs(51)) or (inputs(250));
    layer0_outputs(4959) <= inputs(183);
    layer0_outputs(4960) <= (inputs(101)) and not (inputs(143));
    layer0_outputs(4961) <= (inputs(149)) or (inputs(169));
    layer0_outputs(4962) <= not(inputs(253));
    layer0_outputs(4963) <= (inputs(63)) and not (inputs(28));
    layer0_outputs(4964) <= (inputs(255)) or (inputs(44));
    layer0_outputs(4965) <= '0';
    layer0_outputs(4966) <= (inputs(73)) and not (inputs(134));
    layer0_outputs(4967) <= not(inputs(183));
    layer0_outputs(4968) <= not((inputs(32)) or (inputs(205)));
    layer0_outputs(4969) <= not(inputs(95)) or (inputs(253));
    layer0_outputs(4970) <= inputs(24);
    layer0_outputs(4971) <= inputs(138);
    layer0_outputs(4972) <= (inputs(94)) xor (inputs(103));
    layer0_outputs(4973) <= (inputs(210)) and not (inputs(117));
    layer0_outputs(4974) <= inputs(162);
    layer0_outputs(4975) <= not((inputs(132)) xor (inputs(28)));
    layer0_outputs(4976) <= not(inputs(200)) or (inputs(173));
    layer0_outputs(4977) <= not((inputs(239)) or (inputs(120)));
    layer0_outputs(4978) <= (inputs(82)) or (inputs(2));
    layer0_outputs(4979) <= not(inputs(86));
    layer0_outputs(4980) <= not(inputs(232));
    layer0_outputs(4981) <= not((inputs(67)) or (inputs(49)));
    layer0_outputs(4982) <= (inputs(41)) and not (inputs(6));
    layer0_outputs(4983) <= not(inputs(70));
    layer0_outputs(4984) <= inputs(233);
    layer0_outputs(4985) <= inputs(225);
    layer0_outputs(4986) <= (inputs(126)) and not (inputs(251));
    layer0_outputs(4987) <= not((inputs(120)) xor (inputs(86)));
    layer0_outputs(4988) <= not(inputs(127)) or (inputs(31));
    layer0_outputs(4989) <= not(inputs(38));
    layer0_outputs(4990) <= not((inputs(231)) or (inputs(248)));
    layer0_outputs(4991) <= '1';
    layer0_outputs(4992) <= inputs(151);
    layer0_outputs(4993) <= not(inputs(111));
    layer0_outputs(4994) <= not((inputs(198)) xor (inputs(196)));
    layer0_outputs(4995) <= (inputs(65)) or (inputs(34));
    layer0_outputs(4996) <= (inputs(205)) or (inputs(180));
    layer0_outputs(4997) <= not((inputs(180)) xor (inputs(209)));
    layer0_outputs(4998) <= not(inputs(127));
    layer0_outputs(4999) <= not(inputs(33));
    layer0_outputs(5000) <= (inputs(25)) and not (inputs(231));
    layer0_outputs(5001) <= '0';
    layer0_outputs(5002) <= not(inputs(85)) or (inputs(126));
    layer0_outputs(5003) <= not((inputs(34)) or (inputs(16)));
    layer0_outputs(5004) <= inputs(247);
    layer0_outputs(5005) <= (inputs(114)) xor (inputs(122));
    layer0_outputs(5006) <= (inputs(235)) and not (inputs(110));
    layer0_outputs(5007) <= inputs(103);
    layer0_outputs(5008) <= inputs(178);
    layer0_outputs(5009) <= inputs(72);
    layer0_outputs(5010) <= (inputs(208)) xor (inputs(204));
    layer0_outputs(5011) <= (inputs(74)) xor (inputs(92));
    layer0_outputs(5012) <= not(inputs(18)) or (inputs(60));
    layer0_outputs(5013) <= not(inputs(208)) or (inputs(16));
    layer0_outputs(5014) <= not(inputs(61));
    layer0_outputs(5015) <= (inputs(180)) or (inputs(225));
    layer0_outputs(5016) <= (inputs(133)) or (inputs(142));
    layer0_outputs(5017) <= inputs(79);
    layer0_outputs(5018) <= not((inputs(239)) or (inputs(74)));
    layer0_outputs(5019) <= inputs(57);
    layer0_outputs(5020) <= not((inputs(196)) or (inputs(113)));
    layer0_outputs(5021) <= not((inputs(222)) or (inputs(218)));
    layer0_outputs(5022) <= not((inputs(250)) and (inputs(56)));
    layer0_outputs(5023) <= inputs(69);
    layer0_outputs(5024) <= not(inputs(100)) or (inputs(30));
    layer0_outputs(5025) <= not((inputs(190)) or (inputs(34)));
    layer0_outputs(5026) <= not(inputs(103)) or (inputs(246));
    layer0_outputs(5027) <= inputs(146);
    layer0_outputs(5028) <= not(inputs(54));
    layer0_outputs(5029) <= not(inputs(23)) or (inputs(249));
    layer0_outputs(5030) <= (inputs(141)) xor (inputs(173));
    layer0_outputs(5031) <= not(inputs(5));
    layer0_outputs(5032) <= not((inputs(21)) or (inputs(37)));
    layer0_outputs(5033) <= not(inputs(97));
    layer0_outputs(5034) <= not(inputs(8));
    layer0_outputs(5035) <= not(inputs(149));
    layer0_outputs(5036) <= not((inputs(219)) or (inputs(190)));
    layer0_outputs(5037) <= inputs(23);
    layer0_outputs(5038) <= not(inputs(238));
    layer0_outputs(5039) <= not(inputs(108));
    layer0_outputs(5040) <= not(inputs(83)) or (inputs(157));
    layer0_outputs(5041) <= inputs(66);
    layer0_outputs(5042) <= inputs(30);
    layer0_outputs(5043) <= (inputs(113)) or (inputs(133));
    layer0_outputs(5044) <= not(inputs(152)) or (inputs(202));
    layer0_outputs(5045) <= not(inputs(221)) or (inputs(16));
    layer0_outputs(5046) <= not((inputs(34)) and (inputs(35)));
    layer0_outputs(5047) <= not(inputs(36)) or (inputs(232));
    layer0_outputs(5048) <= not(inputs(24));
    layer0_outputs(5049) <= (inputs(164)) xor (inputs(107));
    layer0_outputs(5050) <= (inputs(100)) or (inputs(194));
    layer0_outputs(5051) <= inputs(106);
    layer0_outputs(5052) <= not(inputs(179));
    layer0_outputs(5053) <= not(inputs(157));
    layer0_outputs(5054) <= (inputs(187)) or (inputs(127));
    layer0_outputs(5055) <= (inputs(235)) xor (inputs(30));
    layer0_outputs(5056) <= (inputs(107)) xor (inputs(173));
    layer0_outputs(5057) <= (inputs(137)) and not (inputs(32));
    layer0_outputs(5058) <= (inputs(239)) or (inputs(176));
    layer0_outputs(5059) <= (inputs(86)) and not (inputs(232));
    layer0_outputs(5060) <= not((inputs(183)) or (inputs(97)));
    layer0_outputs(5061) <= (inputs(186)) and not (inputs(102));
    layer0_outputs(5062) <= not(inputs(114)) or (inputs(41));
    layer0_outputs(5063) <= not((inputs(59)) xor (inputs(161)));
    layer0_outputs(5064) <= (inputs(41)) and (inputs(57));
    layer0_outputs(5065) <= not((inputs(137)) xor (inputs(187)));
    layer0_outputs(5066) <= (inputs(166)) and not (inputs(225));
    layer0_outputs(5067) <= not(inputs(116));
    layer0_outputs(5068) <= not(inputs(8));
    layer0_outputs(5069) <= (inputs(246)) or (inputs(0));
    layer0_outputs(5070) <= (inputs(101)) or (inputs(180));
    layer0_outputs(5071) <= inputs(138);
    layer0_outputs(5072) <= inputs(45);
    layer0_outputs(5073) <= inputs(192);
    layer0_outputs(5074) <= (inputs(89)) and not (inputs(87));
    layer0_outputs(5075) <= (inputs(17)) xor (inputs(69));
    layer0_outputs(5076) <= not((inputs(197)) xor (inputs(164)));
    layer0_outputs(5077) <= (inputs(99)) or (inputs(154));
    layer0_outputs(5078) <= not(inputs(131));
    layer0_outputs(5079) <= (inputs(223)) xor (inputs(217));
    layer0_outputs(5080) <= not((inputs(206)) xor (inputs(91)));
    layer0_outputs(5081) <= inputs(132);
    layer0_outputs(5082) <= not(inputs(53)) or (inputs(108));
    layer0_outputs(5083) <= not((inputs(119)) or (inputs(159)));
    layer0_outputs(5084) <= not(inputs(148));
    layer0_outputs(5085) <= (inputs(113)) xor (inputs(216));
    layer0_outputs(5086) <= not(inputs(90));
    layer0_outputs(5087) <= (inputs(105)) and not (inputs(159));
    layer0_outputs(5088) <= not((inputs(123)) or (inputs(42)));
    layer0_outputs(5089) <= not(inputs(138));
    layer0_outputs(5090) <= not((inputs(67)) or (inputs(103)));
    layer0_outputs(5091) <= not(inputs(215)) or (inputs(239));
    layer0_outputs(5092) <= inputs(219);
    layer0_outputs(5093) <= (inputs(228)) and not (inputs(47));
    layer0_outputs(5094) <= '0';
    layer0_outputs(5095) <= not((inputs(64)) or (inputs(135)));
    layer0_outputs(5096) <= not((inputs(237)) or (inputs(105)));
    layer0_outputs(5097) <= not((inputs(52)) or (inputs(26)));
    layer0_outputs(5098) <= not(inputs(132));
    layer0_outputs(5099) <= (inputs(42)) and not (inputs(145));
    layer0_outputs(5100) <= not((inputs(19)) or (inputs(126)));
    layer0_outputs(5101) <= '1';
    layer0_outputs(5102) <= not(inputs(87));
    layer0_outputs(5103) <= not(inputs(116)) or (inputs(125));
    layer0_outputs(5104) <= (inputs(36)) or (inputs(77));
    layer0_outputs(5105) <= inputs(188);
    layer0_outputs(5106) <= not(inputs(23)) or (inputs(112));
    layer0_outputs(5107) <= not((inputs(155)) or (inputs(126)));
    layer0_outputs(5108) <= (inputs(41)) and not (inputs(0));
    layer0_outputs(5109) <= (inputs(133)) xor (inputs(17));
    layer0_outputs(5110) <= not(inputs(22));
    layer0_outputs(5111) <= not((inputs(205)) or (inputs(11)));
    layer0_outputs(5112) <= (inputs(148)) and not (inputs(109));
    layer0_outputs(5113) <= not(inputs(146));
    layer0_outputs(5114) <= inputs(103);
    layer0_outputs(5115) <= (inputs(181)) or (inputs(16));
    layer0_outputs(5116) <= not((inputs(156)) xor (inputs(16)));
    layer0_outputs(5117) <= not(inputs(78));
    layer0_outputs(5118) <= not(inputs(19));
    layer0_outputs(5119) <= inputs(102);
    layer0_outputs(5120) <= not(inputs(84)) or (inputs(55));
    layer0_outputs(5121) <= (inputs(209)) and (inputs(215));
    layer0_outputs(5122) <= not(inputs(75)) or (inputs(8));
    layer0_outputs(5123) <= (inputs(84)) xor (inputs(111));
    layer0_outputs(5124) <= inputs(115);
    layer0_outputs(5125) <= (inputs(121)) and (inputs(143));
    layer0_outputs(5126) <= not((inputs(159)) or (inputs(214)));
    layer0_outputs(5127) <= not((inputs(98)) xor (inputs(74)));
    layer0_outputs(5128) <= not(inputs(139));
    layer0_outputs(5129) <= inputs(19);
    layer0_outputs(5130) <= (inputs(29)) and not (inputs(70));
    layer0_outputs(5131) <= (inputs(90)) and not (inputs(128));
    layer0_outputs(5132) <= not(inputs(58)) or (inputs(177));
    layer0_outputs(5133) <= (inputs(177)) xor (inputs(28));
    layer0_outputs(5134) <= not(inputs(192));
    layer0_outputs(5135) <= '0';
    layer0_outputs(5136) <= (inputs(243)) and not (inputs(0));
    layer0_outputs(5137) <= not((inputs(243)) or (inputs(208)));
    layer0_outputs(5138) <= (inputs(191)) xor (inputs(62));
    layer0_outputs(5139) <= (inputs(9)) xor (inputs(21));
    layer0_outputs(5140) <= inputs(246);
    layer0_outputs(5141) <= not(inputs(182));
    layer0_outputs(5142) <= inputs(217);
    layer0_outputs(5143) <= (inputs(76)) and not (inputs(17));
    layer0_outputs(5144) <= not(inputs(225));
    layer0_outputs(5145) <= inputs(40);
    layer0_outputs(5146) <= not((inputs(98)) xor (inputs(151)));
    layer0_outputs(5147) <= not(inputs(81)) or (inputs(240));
    layer0_outputs(5148) <= not(inputs(178)) or (inputs(155));
    layer0_outputs(5149) <= not(inputs(132));
    layer0_outputs(5150) <= (inputs(194)) and not (inputs(70));
    layer0_outputs(5151) <= (inputs(143)) or (inputs(67));
    layer0_outputs(5152) <= not(inputs(84));
    layer0_outputs(5153) <= not(inputs(99));
    layer0_outputs(5154) <= not(inputs(106)) or (inputs(196));
    layer0_outputs(5155) <= not(inputs(249)) or (inputs(77));
    layer0_outputs(5156) <= inputs(59);
    layer0_outputs(5157) <= '1';
    layer0_outputs(5158) <= not((inputs(163)) or (inputs(210)));
    layer0_outputs(5159) <= (inputs(89)) or (inputs(145));
    layer0_outputs(5160) <= not(inputs(247));
    layer0_outputs(5161) <= not(inputs(58)) or (inputs(252));
    layer0_outputs(5162) <= (inputs(83)) and not (inputs(90));
    layer0_outputs(5163) <= (inputs(124)) xor (inputs(92));
    layer0_outputs(5164) <= inputs(10);
    layer0_outputs(5165) <= inputs(131);
    layer0_outputs(5166) <= '0';
    layer0_outputs(5167) <= not(inputs(51)) or (inputs(145));
    layer0_outputs(5168) <= (inputs(7)) xor (inputs(225));
    layer0_outputs(5169) <= not(inputs(150));
    layer0_outputs(5170) <= (inputs(200)) and not (inputs(11));
    layer0_outputs(5171) <= not((inputs(225)) xor (inputs(179)));
    layer0_outputs(5172) <= inputs(245);
    layer0_outputs(5173) <= inputs(173);
    layer0_outputs(5174) <= not(inputs(217));
    layer0_outputs(5175) <= inputs(206);
    layer0_outputs(5176) <= inputs(228);
    layer0_outputs(5177) <= (inputs(173)) and (inputs(141));
    layer0_outputs(5178) <= not(inputs(245)) or (inputs(17));
    layer0_outputs(5179) <= not((inputs(19)) or (inputs(110)));
    layer0_outputs(5180) <= (inputs(235)) xor (inputs(142));
    layer0_outputs(5181) <= inputs(175);
    layer0_outputs(5182) <= (inputs(155)) or (inputs(149));
    layer0_outputs(5183) <= (inputs(22)) and not (inputs(107));
    layer0_outputs(5184) <= not(inputs(9)) or (inputs(131));
    layer0_outputs(5185) <= not((inputs(126)) xor (inputs(129)));
    layer0_outputs(5186) <= not(inputs(36));
    layer0_outputs(5187) <= not((inputs(172)) and (inputs(192)));
    layer0_outputs(5188) <= (inputs(54)) or (inputs(234));
    layer0_outputs(5189) <= not((inputs(155)) or (inputs(21)));
    layer0_outputs(5190) <= (inputs(232)) and not (inputs(117));
    layer0_outputs(5191) <= not(inputs(231)) or (inputs(240));
    layer0_outputs(5192) <= inputs(53);
    layer0_outputs(5193) <= not(inputs(53));
    layer0_outputs(5194) <= not((inputs(63)) xor (inputs(14)));
    layer0_outputs(5195) <= not(inputs(130)) or (inputs(63));
    layer0_outputs(5196) <= not((inputs(255)) or (inputs(61)));
    layer0_outputs(5197) <= not(inputs(196));
    layer0_outputs(5198) <= not(inputs(217));
    layer0_outputs(5199) <= not((inputs(37)) or (inputs(2)));
    layer0_outputs(5200) <= not((inputs(39)) xor (inputs(76)));
    layer0_outputs(5201) <= not(inputs(75));
    layer0_outputs(5202) <= (inputs(56)) and not (inputs(149));
    layer0_outputs(5203) <= (inputs(214)) and not (inputs(83));
    layer0_outputs(5204) <= (inputs(57)) or (inputs(143));
    layer0_outputs(5205) <= (inputs(215)) or (inputs(147));
    layer0_outputs(5206) <= not(inputs(36)) or (inputs(43));
    layer0_outputs(5207) <= (inputs(151)) and not (inputs(191));
    layer0_outputs(5208) <= '1';
    layer0_outputs(5209) <= not(inputs(164)) or (inputs(32));
    layer0_outputs(5210) <= (inputs(245)) or (inputs(163));
    layer0_outputs(5211) <= not(inputs(236)) or (inputs(179));
    layer0_outputs(5212) <= inputs(242);
    layer0_outputs(5213) <= (inputs(189)) xor (inputs(0));
    layer0_outputs(5214) <= not(inputs(181)) or (inputs(111));
    layer0_outputs(5215) <= not(inputs(231));
    layer0_outputs(5216) <= not(inputs(180));
    layer0_outputs(5217) <= not(inputs(130)) or (inputs(79));
    layer0_outputs(5218) <= not(inputs(232)) or (inputs(127));
    layer0_outputs(5219) <= not(inputs(110));
    layer0_outputs(5220) <= not(inputs(165));
    layer0_outputs(5221) <= not(inputs(55));
    layer0_outputs(5222) <= not((inputs(224)) xor (inputs(29)));
    layer0_outputs(5223) <= (inputs(115)) and (inputs(40));
    layer0_outputs(5224) <= inputs(182);
    layer0_outputs(5225) <= inputs(221);
    layer0_outputs(5226) <= (inputs(164)) and not (inputs(14));
    layer0_outputs(5227) <= inputs(94);
    layer0_outputs(5228) <= inputs(130);
    layer0_outputs(5229) <= inputs(125);
    layer0_outputs(5230) <= (inputs(164)) or (inputs(143));
    layer0_outputs(5231) <= (inputs(157)) or (inputs(116));
    layer0_outputs(5232) <= not(inputs(113));
    layer0_outputs(5233) <= inputs(117);
    layer0_outputs(5234) <= (inputs(249)) or (inputs(229));
    layer0_outputs(5235) <= (inputs(6)) xor (inputs(159));
    layer0_outputs(5236) <= not(inputs(228)) or (inputs(252));
    layer0_outputs(5237) <= not(inputs(135));
    layer0_outputs(5238) <= not(inputs(88));
    layer0_outputs(5239) <= (inputs(236)) xor (inputs(161));
    layer0_outputs(5240) <= (inputs(74)) and (inputs(132));
    layer0_outputs(5241) <= inputs(163);
    layer0_outputs(5242) <= not(inputs(98));
    layer0_outputs(5243) <= not((inputs(17)) or (inputs(221)));
    layer0_outputs(5244) <= (inputs(63)) and not (inputs(4));
    layer0_outputs(5245) <= not(inputs(84)) or (inputs(143));
    layer0_outputs(5246) <= not((inputs(31)) or (inputs(118)));
    layer0_outputs(5247) <= not((inputs(75)) or (inputs(28)));
    layer0_outputs(5248) <= (inputs(21)) and not (inputs(204));
    layer0_outputs(5249) <= (inputs(43)) or (inputs(176));
    layer0_outputs(5250) <= not(inputs(208)) or (inputs(156));
    layer0_outputs(5251) <= inputs(174);
    layer0_outputs(5252) <= '1';
    layer0_outputs(5253) <= (inputs(23)) and (inputs(12));
    layer0_outputs(5254) <= inputs(28);
    layer0_outputs(5255) <= (inputs(62)) and (inputs(124));
    layer0_outputs(5256) <= (inputs(45)) or (inputs(62));
    layer0_outputs(5257) <= not(inputs(26));
    layer0_outputs(5258) <= (inputs(18)) or (inputs(45));
    layer0_outputs(5259) <= not((inputs(124)) or (inputs(59)));
    layer0_outputs(5260) <= not((inputs(232)) xor (inputs(186)));
    layer0_outputs(5261) <= not((inputs(94)) or (inputs(23)));
    layer0_outputs(5262) <= not(inputs(143));
    layer0_outputs(5263) <= inputs(61);
    layer0_outputs(5264) <= not(inputs(34));
    layer0_outputs(5265) <= not((inputs(128)) xor (inputs(116)));
    layer0_outputs(5266) <= (inputs(8)) and not (inputs(98));
    layer0_outputs(5267) <= (inputs(50)) or (inputs(142));
    layer0_outputs(5268) <= inputs(69);
    layer0_outputs(5269) <= not(inputs(120));
    layer0_outputs(5270) <= inputs(90);
    layer0_outputs(5271) <= (inputs(114)) and not (inputs(16));
    layer0_outputs(5272) <= not(inputs(38));
    layer0_outputs(5273) <= not((inputs(147)) or (inputs(130)));
    layer0_outputs(5274) <= inputs(186);
    layer0_outputs(5275) <= inputs(85);
    layer0_outputs(5276) <= inputs(98);
    layer0_outputs(5277) <= inputs(196);
    layer0_outputs(5278) <= (inputs(217)) and not (inputs(167));
    layer0_outputs(5279) <= (inputs(118)) and not (inputs(159));
    layer0_outputs(5280) <= (inputs(85)) and not (inputs(113));
    layer0_outputs(5281) <= (inputs(60)) or (inputs(254));
    layer0_outputs(5282) <= not(inputs(26));
    layer0_outputs(5283) <= not(inputs(208));
    layer0_outputs(5284) <= not(inputs(22));
    layer0_outputs(5285) <= (inputs(17)) and not (inputs(80));
    layer0_outputs(5286) <= inputs(68);
    layer0_outputs(5287) <= not(inputs(151));
    layer0_outputs(5288) <= not(inputs(198)) or (inputs(125));
    layer0_outputs(5289) <= (inputs(159)) xor (inputs(42));
    layer0_outputs(5290) <= not(inputs(226));
    layer0_outputs(5291) <= inputs(5);
    layer0_outputs(5292) <= not(inputs(39)) or (inputs(217));
    layer0_outputs(5293) <= not(inputs(28)) or (inputs(15));
    layer0_outputs(5294) <= not(inputs(137));
    layer0_outputs(5295) <= (inputs(39)) and not (inputs(141));
    layer0_outputs(5296) <= inputs(214);
    layer0_outputs(5297) <= '1';
    layer0_outputs(5298) <= not((inputs(153)) or (inputs(68)));
    layer0_outputs(5299) <= inputs(0);
    layer0_outputs(5300) <= (inputs(163)) and not (inputs(35));
    layer0_outputs(5301) <= inputs(100);
    layer0_outputs(5302) <= (inputs(107)) and not (inputs(112));
    layer0_outputs(5303) <= inputs(91);
    layer0_outputs(5304) <= '1';
    layer0_outputs(5305) <= not(inputs(237));
    layer0_outputs(5306) <= inputs(23);
    layer0_outputs(5307) <= not(inputs(158));
    layer0_outputs(5308) <= not(inputs(9));
    layer0_outputs(5309) <= (inputs(244)) or (inputs(243));
    layer0_outputs(5310) <= not(inputs(186)) or (inputs(239));
    layer0_outputs(5311) <= (inputs(225)) xor (inputs(164));
    layer0_outputs(5312) <= '0';
    layer0_outputs(5313) <= (inputs(226)) xor (inputs(153));
    layer0_outputs(5314) <= (inputs(170)) or (inputs(204));
    layer0_outputs(5315) <= inputs(86);
    layer0_outputs(5316) <= not(inputs(190)) or (inputs(112));
    layer0_outputs(5317) <= '1';
    layer0_outputs(5318) <= (inputs(10)) or (inputs(97));
    layer0_outputs(5319) <= (inputs(105)) or (inputs(16));
    layer0_outputs(5320) <= not(inputs(184));
    layer0_outputs(5321) <= (inputs(69)) xor (inputs(66));
    layer0_outputs(5322) <= inputs(77);
    layer0_outputs(5323) <= (inputs(241)) or (inputs(22));
    layer0_outputs(5324) <= (inputs(157)) and not (inputs(0));
    layer0_outputs(5325) <= inputs(112);
    layer0_outputs(5326) <= not(inputs(10)) or (inputs(32));
    layer0_outputs(5327) <= (inputs(52)) or (inputs(78));
    layer0_outputs(5328) <= not(inputs(134)) or (inputs(138));
    layer0_outputs(5329) <= not((inputs(30)) or (inputs(129)));
    layer0_outputs(5330) <= not((inputs(3)) or (inputs(131)));
    layer0_outputs(5331) <= inputs(87);
    layer0_outputs(5332) <= (inputs(249)) and (inputs(234));
    layer0_outputs(5333) <= (inputs(28)) and not (inputs(159));
    layer0_outputs(5334) <= not((inputs(114)) or (inputs(116)));
    layer0_outputs(5335) <= not(inputs(52));
    layer0_outputs(5336) <= inputs(38);
    layer0_outputs(5337) <= inputs(247);
    layer0_outputs(5338) <= not(inputs(246)) or (inputs(50));
    layer0_outputs(5339) <= '0';
    layer0_outputs(5340) <= (inputs(156)) xor (inputs(176));
    layer0_outputs(5341) <= (inputs(8)) and not (inputs(249));
    layer0_outputs(5342) <= not((inputs(201)) or (inputs(204)));
    layer0_outputs(5343) <= (inputs(108)) and not (inputs(194));
    layer0_outputs(5344) <= not((inputs(150)) or (inputs(191)));
    layer0_outputs(5345) <= not((inputs(127)) or (inputs(54)));
    layer0_outputs(5346) <= inputs(177);
    layer0_outputs(5347) <= '0';
    layer0_outputs(5348) <= not(inputs(82)) or (inputs(56));
    layer0_outputs(5349) <= (inputs(105)) and not (inputs(243));
    layer0_outputs(5350) <= inputs(113);
    layer0_outputs(5351) <= inputs(24);
    layer0_outputs(5352) <= not((inputs(148)) or (inputs(178)));
    layer0_outputs(5353) <= not((inputs(153)) xor (inputs(155)));
    layer0_outputs(5354) <= not((inputs(21)) or (inputs(177)));
    layer0_outputs(5355) <= not((inputs(102)) or (inputs(239)));
    layer0_outputs(5356) <= not(inputs(201)) or (inputs(135));
    layer0_outputs(5357) <= not(inputs(147));
    layer0_outputs(5358) <= not(inputs(60));
    layer0_outputs(5359) <= (inputs(46)) and not (inputs(112));
    layer0_outputs(5360) <= (inputs(41)) or (inputs(30));
    layer0_outputs(5361) <= inputs(171);
    layer0_outputs(5362) <= (inputs(62)) and (inputs(61));
    layer0_outputs(5363) <= inputs(99);
    layer0_outputs(5364) <= (inputs(255)) or (inputs(90));
    layer0_outputs(5365) <= not((inputs(147)) or (inputs(239)));
    layer0_outputs(5366) <= not(inputs(238));
    layer0_outputs(5367) <= (inputs(33)) or (inputs(216));
    layer0_outputs(5368) <= not((inputs(143)) xor (inputs(116)));
    layer0_outputs(5369) <= not((inputs(93)) xor (inputs(56)));
    layer0_outputs(5370) <= (inputs(210)) or (inputs(145));
    layer0_outputs(5371) <= not(inputs(3)) or (inputs(67));
    layer0_outputs(5372) <= not(inputs(106));
    layer0_outputs(5373) <= not(inputs(122));
    layer0_outputs(5374) <= (inputs(59)) or (inputs(28));
    layer0_outputs(5375) <= not((inputs(89)) xor (inputs(45)));
    layer0_outputs(5376) <= (inputs(46)) and (inputs(193));
    layer0_outputs(5377) <= (inputs(123)) or (inputs(89));
    layer0_outputs(5378) <= not(inputs(217));
    layer0_outputs(5379) <= inputs(167);
    layer0_outputs(5380) <= (inputs(141)) and not (inputs(97));
    layer0_outputs(5381) <= not(inputs(225)) or (inputs(147));
    layer0_outputs(5382) <= inputs(103);
    layer0_outputs(5383) <= (inputs(53)) or (inputs(62));
    layer0_outputs(5384) <= not(inputs(108));
    layer0_outputs(5385) <= (inputs(35)) xor (inputs(250));
    layer0_outputs(5386) <= not(inputs(82));
    layer0_outputs(5387) <= not(inputs(152));
    layer0_outputs(5388) <= not((inputs(15)) xor (inputs(46)));
    layer0_outputs(5389) <= not(inputs(59));
    layer0_outputs(5390) <= (inputs(124)) xor (inputs(170));
    layer0_outputs(5391) <= inputs(195);
    layer0_outputs(5392) <= (inputs(33)) or (inputs(3));
    layer0_outputs(5393) <= (inputs(73)) and not (inputs(217));
    layer0_outputs(5394) <= '0';
    layer0_outputs(5395) <= not((inputs(29)) or (inputs(80)));
    layer0_outputs(5396) <= not(inputs(104));
    layer0_outputs(5397) <= (inputs(101)) xor (inputs(144));
    layer0_outputs(5398) <= (inputs(102)) or (inputs(226));
    layer0_outputs(5399) <= not((inputs(132)) or (inputs(126)));
    layer0_outputs(5400) <= not(inputs(163));
    layer0_outputs(5401) <= not((inputs(49)) xor (inputs(86)));
    layer0_outputs(5402) <= not(inputs(192)) or (inputs(207));
    layer0_outputs(5403) <= not(inputs(189));
    layer0_outputs(5404) <= not(inputs(89)) or (inputs(139));
    layer0_outputs(5405) <= inputs(27);
    layer0_outputs(5406) <= (inputs(59)) and not (inputs(254));
    layer0_outputs(5407) <= not((inputs(132)) and (inputs(179)));
    layer0_outputs(5408) <= not((inputs(32)) or (inputs(26)));
    layer0_outputs(5409) <= not((inputs(142)) or (inputs(51)));
    layer0_outputs(5410) <= not(inputs(237));
    layer0_outputs(5411) <= '1';
    layer0_outputs(5412) <= not((inputs(146)) xor (inputs(192)));
    layer0_outputs(5413) <= inputs(205);
    layer0_outputs(5414) <= not(inputs(27)) or (inputs(5));
    layer0_outputs(5415) <= (inputs(233)) or (inputs(66));
    layer0_outputs(5416) <= (inputs(122)) or (inputs(109));
    layer0_outputs(5417) <= not(inputs(118)) or (inputs(192));
    layer0_outputs(5418) <= (inputs(38)) xor (inputs(35));
    layer0_outputs(5419) <= not(inputs(83));
    layer0_outputs(5420) <= not(inputs(72)) or (inputs(1));
    layer0_outputs(5421) <= not(inputs(143));
    layer0_outputs(5422) <= not(inputs(206));
    layer0_outputs(5423) <= not((inputs(143)) or (inputs(112)));
    layer0_outputs(5424) <= inputs(88);
    layer0_outputs(5425) <= not((inputs(8)) and (inputs(75)));
    layer0_outputs(5426) <= not(inputs(182));
    layer0_outputs(5427) <= (inputs(89)) xor (inputs(148));
    layer0_outputs(5428) <= (inputs(190)) or (inputs(133));
    layer0_outputs(5429) <= (inputs(145)) and not (inputs(33));
    layer0_outputs(5430) <= (inputs(214)) or (inputs(233));
    layer0_outputs(5431) <= inputs(122);
    layer0_outputs(5432) <= inputs(148);
    layer0_outputs(5433) <= not(inputs(223)) or (inputs(0));
    layer0_outputs(5434) <= (inputs(23)) and not (inputs(190));
    layer0_outputs(5435) <= not(inputs(173));
    layer0_outputs(5436) <= (inputs(128)) xor (inputs(87));
    layer0_outputs(5437) <= '0';
    layer0_outputs(5438) <= (inputs(160)) and not (inputs(161));
    layer0_outputs(5439) <= not(inputs(247));
    layer0_outputs(5440) <= inputs(183);
    layer0_outputs(5441) <= not((inputs(37)) and (inputs(56)));
    layer0_outputs(5442) <= inputs(231);
    layer0_outputs(5443) <= not((inputs(55)) or (inputs(47)));
    layer0_outputs(5444) <= (inputs(186)) or (inputs(202));
    layer0_outputs(5445) <= not(inputs(92));
    layer0_outputs(5446) <= (inputs(128)) or (inputs(25));
    layer0_outputs(5447) <= not(inputs(162)) or (inputs(87));
    layer0_outputs(5448) <= not(inputs(120)) or (inputs(9));
    layer0_outputs(5449) <= not((inputs(116)) or (inputs(2)));
    layer0_outputs(5450) <= not(inputs(210));
    layer0_outputs(5451) <= not((inputs(196)) xor (inputs(152)));
    layer0_outputs(5452) <= not(inputs(197));
    layer0_outputs(5453) <= not(inputs(181));
    layer0_outputs(5454) <= not(inputs(246));
    layer0_outputs(5455) <= inputs(211);
    layer0_outputs(5456) <= (inputs(248)) and not (inputs(168));
    layer0_outputs(5457) <= inputs(157);
    layer0_outputs(5458) <= '1';
    layer0_outputs(5459) <= (inputs(216)) and not (inputs(134));
    layer0_outputs(5460) <= (inputs(228)) and not (inputs(129));
    layer0_outputs(5461) <= not((inputs(83)) xor (inputs(69)));
    layer0_outputs(5462) <= inputs(209);
    layer0_outputs(5463) <= (inputs(118)) xor (inputs(181));
    layer0_outputs(5464) <= not((inputs(82)) or (inputs(181)));
    layer0_outputs(5465) <= inputs(148);
    layer0_outputs(5466) <= not(inputs(199));
    layer0_outputs(5467) <= not((inputs(60)) or (inputs(108)));
    layer0_outputs(5468) <= not(inputs(231)) or (inputs(163));
    layer0_outputs(5469) <= (inputs(247)) or (inputs(157));
    layer0_outputs(5470) <= not((inputs(101)) xor (inputs(107)));
    layer0_outputs(5471) <= not((inputs(162)) xor (inputs(167)));
    layer0_outputs(5472) <= (inputs(56)) and not (inputs(244));
    layer0_outputs(5473) <= not(inputs(19));
    layer0_outputs(5474) <= not(inputs(1)) or (inputs(162));
    layer0_outputs(5475) <= not(inputs(218));
    layer0_outputs(5476) <= not(inputs(246));
    layer0_outputs(5477) <= not(inputs(235));
    layer0_outputs(5478) <= inputs(236);
    layer0_outputs(5479) <= (inputs(82)) or (inputs(180));
    layer0_outputs(5480) <= inputs(239);
    layer0_outputs(5481) <= not((inputs(10)) or (inputs(27)));
    layer0_outputs(5482) <= (inputs(171)) and not (inputs(13));
    layer0_outputs(5483) <= not(inputs(126)) or (inputs(79));
    layer0_outputs(5484) <= (inputs(13)) and not (inputs(71));
    layer0_outputs(5485) <= (inputs(36)) or (inputs(77));
    layer0_outputs(5486) <= (inputs(4)) xor (inputs(174));
    layer0_outputs(5487) <= (inputs(182)) or (inputs(47));
    layer0_outputs(5488) <= not(inputs(252));
    layer0_outputs(5489) <= inputs(150);
    layer0_outputs(5490) <= inputs(166);
    layer0_outputs(5491) <= (inputs(233)) and not (inputs(39));
    layer0_outputs(5492) <= (inputs(138)) xor (inputs(100));
    layer0_outputs(5493) <= not(inputs(15));
    layer0_outputs(5494) <= not(inputs(152));
    layer0_outputs(5495) <= (inputs(243)) xor (inputs(212));
    layer0_outputs(5496) <= (inputs(246)) and not (inputs(112));
    layer0_outputs(5497) <= not(inputs(98));
    layer0_outputs(5498) <= (inputs(22)) and not (inputs(178));
    layer0_outputs(5499) <= (inputs(85)) or (inputs(164));
    layer0_outputs(5500) <= (inputs(194)) xor (inputs(190));
    layer0_outputs(5501) <= not((inputs(216)) or (inputs(175)));
    layer0_outputs(5502) <= (inputs(165)) xor (inputs(169));
    layer0_outputs(5503) <= (inputs(228)) and not (inputs(75));
    layer0_outputs(5504) <= (inputs(85)) or (inputs(133));
    layer0_outputs(5505) <= (inputs(240)) or (inputs(29));
    layer0_outputs(5506) <= not(inputs(27));
    layer0_outputs(5507) <= (inputs(93)) or (inputs(105));
    layer0_outputs(5508) <= not(inputs(217)) or (inputs(110));
    layer0_outputs(5509) <= (inputs(14)) xor (inputs(194));
    layer0_outputs(5510) <= not(inputs(95)) or (inputs(74));
    layer0_outputs(5511) <= not(inputs(114)) or (inputs(15));
    layer0_outputs(5512) <= (inputs(56)) and not (inputs(116));
    layer0_outputs(5513) <= not((inputs(46)) or (inputs(97)));
    layer0_outputs(5514) <= not(inputs(57));
    layer0_outputs(5515) <= '1';
    layer0_outputs(5516) <= not(inputs(88)) or (inputs(152));
    layer0_outputs(5517) <= not((inputs(5)) xor (inputs(176)));
    layer0_outputs(5518) <= inputs(59);
    layer0_outputs(5519) <= not(inputs(152)) or (inputs(98));
    layer0_outputs(5520) <= '0';
    layer0_outputs(5521) <= not((inputs(255)) or (inputs(39)));
    layer0_outputs(5522) <= not(inputs(168)) or (inputs(149));
    layer0_outputs(5523) <= (inputs(229)) xor (inputs(182));
    layer0_outputs(5524) <= not(inputs(151)) or (inputs(24));
    layer0_outputs(5525) <= (inputs(77)) or (inputs(7));
    layer0_outputs(5526) <= not((inputs(170)) and (inputs(229)));
    layer0_outputs(5527) <= not(inputs(141));
    layer0_outputs(5528) <= not((inputs(238)) or (inputs(206)));
    layer0_outputs(5529) <= not((inputs(255)) or (inputs(252)));
    layer0_outputs(5530) <= not(inputs(74)) or (inputs(71));
    layer0_outputs(5531) <= not(inputs(179));
    layer0_outputs(5532) <= not(inputs(162)) or (inputs(240));
    layer0_outputs(5533) <= (inputs(84)) xor (inputs(227));
    layer0_outputs(5534) <= inputs(115);
    layer0_outputs(5535) <= (inputs(190)) xor (inputs(27));
    layer0_outputs(5536) <= inputs(93);
    layer0_outputs(5537) <= inputs(141);
    layer0_outputs(5538) <= not(inputs(76));
    layer0_outputs(5539) <= inputs(144);
    layer0_outputs(5540) <= (inputs(87)) and not (inputs(238));
    layer0_outputs(5541) <= not((inputs(187)) or (inputs(186)));
    layer0_outputs(5542) <= (inputs(140)) and not (inputs(217));
    layer0_outputs(5543) <= (inputs(253)) or (inputs(180));
    layer0_outputs(5544) <= not((inputs(127)) or (inputs(71)));
    layer0_outputs(5545) <= '1';
    layer0_outputs(5546) <= not(inputs(54));
    layer0_outputs(5547) <= not(inputs(99));
    layer0_outputs(5548) <= not(inputs(193));
    layer0_outputs(5549) <= (inputs(164)) and not (inputs(204));
    layer0_outputs(5550) <= (inputs(63)) or (inputs(3));
    layer0_outputs(5551) <= not((inputs(183)) xor (inputs(175)));
    layer0_outputs(5552) <= (inputs(19)) or (inputs(209));
    layer0_outputs(5553) <= (inputs(51)) and (inputs(220));
    layer0_outputs(5554) <= (inputs(209)) or (inputs(252));
    layer0_outputs(5555) <= (inputs(9)) or (inputs(78));
    layer0_outputs(5556) <= (inputs(250)) or (inputs(161));
    layer0_outputs(5557) <= not((inputs(26)) and (inputs(234)));
    layer0_outputs(5558) <= (inputs(171)) xor (inputs(220));
    layer0_outputs(5559) <= inputs(141);
    layer0_outputs(5560) <= not(inputs(66));
    layer0_outputs(5561) <= (inputs(203)) xor (inputs(62));
    layer0_outputs(5562) <= inputs(178);
    layer0_outputs(5563) <= not(inputs(221));
    layer0_outputs(5564) <= (inputs(149)) or (inputs(17));
    layer0_outputs(5565) <= not(inputs(41));
    layer0_outputs(5566) <= inputs(172);
    layer0_outputs(5567) <= not(inputs(12)) or (inputs(167));
    layer0_outputs(5568) <= not((inputs(171)) and (inputs(249)));
    layer0_outputs(5569) <= inputs(25);
    layer0_outputs(5570) <= (inputs(137)) and not (inputs(96));
    layer0_outputs(5571) <= not(inputs(45));
    layer0_outputs(5572) <= (inputs(12)) xor (inputs(63));
    layer0_outputs(5573) <= not(inputs(56)) or (inputs(16));
    layer0_outputs(5574) <= not(inputs(8)) or (inputs(14));
    layer0_outputs(5575) <= (inputs(93)) or (inputs(85));
    layer0_outputs(5576) <= inputs(46);
    layer0_outputs(5577) <= (inputs(104)) and not (inputs(68));
    layer0_outputs(5578) <= inputs(1);
    layer0_outputs(5579) <= not(inputs(138));
    layer0_outputs(5580) <= (inputs(7)) or (inputs(19));
    layer0_outputs(5581) <= (inputs(12)) or (inputs(167));
    layer0_outputs(5582) <= (inputs(227)) or (inputs(253));
    layer0_outputs(5583) <= inputs(190);
    layer0_outputs(5584) <= not((inputs(158)) or (inputs(147)));
    layer0_outputs(5585) <= not(inputs(118)) or (inputs(177));
    layer0_outputs(5586) <= not((inputs(245)) or (inputs(58)));
    layer0_outputs(5587) <= (inputs(132)) and not (inputs(175));
    layer0_outputs(5588) <= not((inputs(92)) or (inputs(125)));
    layer0_outputs(5589) <= not((inputs(38)) xor (inputs(124)));
    layer0_outputs(5590) <= not((inputs(124)) or (inputs(125)));
    layer0_outputs(5591) <= not((inputs(140)) xor (inputs(174)));
    layer0_outputs(5592) <= not((inputs(190)) or (inputs(34)));
    layer0_outputs(5593) <= inputs(233);
    layer0_outputs(5594) <= (inputs(174)) xor (inputs(70));
    layer0_outputs(5595) <= (inputs(149)) or (inputs(222));
    layer0_outputs(5596) <= inputs(100);
    layer0_outputs(5597) <= '0';
    layer0_outputs(5598) <= not((inputs(157)) and (inputs(247)));
    layer0_outputs(5599) <= (inputs(240)) and not (inputs(63));
    layer0_outputs(5600) <= not((inputs(138)) or (inputs(26)));
    layer0_outputs(5601) <= (inputs(40)) or (inputs(117));
    layer0_outputs(5602) <= (inputs(151)) xor (inputs(171));
    layer0_outputs(5603) <= (inputs(77)) xor (inputs(22));
    layer0_outputs(5604) <= (inputs(11)) xor (inputs(95));
    layer0_outputs(5605) <= inputs(157);
    layer0_outputs(5606) <= not((inputs(63)) xor (inputs(29)));
    layer0_outputs(5607) <= inputs(164);
    layer0_outputs(5608) <= not((inputs(248)) or (inputs(2)));
    layer0_outputs(5609) <= inputs(85);
    layer0_outputs(5610) <= not((inputs(160)) or (inputs(63)));
    layer0_outputs(5611) <= not((inputs(112)) or (inputs(115)));
    layer0_outputs(5612) <= (inputs(77)) or (inputs(34));
    layer0_outputs(5613) <= not((inputs(94)) xor (inputs(92)));
    layer0_outputs(5614) <= inputs(149);
    layer0_outputs(5615) <= (inputs(116)) or (inputs(193));
    layer0_outputs(5616) <= not((inputs(235)) or (inputs(209)));
    layer0_outputs(5617) <= inputs(82);
    layer0_outputs(5618) <= inputs(170);
    layer0_outputs(5619) <= not((inputs(91)) or (inputs(93)));
    layer0_outputs(5620) <= (inputs(196)) or (inputs(13));
    layer0_outputs(5621) <= (inputs(81)) and not (inputs(14));
    layer0_outputs(5622) <= not(inputs(122));
    layer0_outputs(5623) <= not(inputs(39));
    layer0_outputs(5624) <= not((inputs(194)) or (inputs(162)));
    layer0_outputs(5625) <= not((inputs(84)) or (inputs(4)));
    layer0_outputs(5626) <= not(inputs(24)) or (inputs(180));
    layer0_outputs(5627) <= (inputs(153)) xor (inputs(118));
    layer0_outputs(5628) <= not((inputs(107)) and (inputs(121)));
    layer0_outputs(5629) <= not(inputs(22)) or (inputs(160));
    layer0_outputs(5630) <= not((inputs(31)) xor (inputs(134)));
    layer0_outputs(5631) <= not((inputs(88)) or (inputs(195)));
    layer0_outputs(5632) <= '1';
    layer0_outputs(5633) <= (inputs(216)) or (inputs(6));
    layer0_outputs(5634) <= inputs(40);
    layer0_outputs(5635) <= not(inputs(99));
    layer0_outputs(5636) <= '1';
    layer0_outputs(5637) <= not(inputs(248));
    layer0_outputs(5638) <= not(inputs(14)) or (inputs(52));
    layer0_outputs(5639) <= (inputs(151)) and (inputs(166));
    layer0_outputs(5640) <= (inputs(230)) and not (inputs(46));
    layer0_outputs(5641) <= not((inputs(2)) or (inputs(150)));
    layer0_outputs(5642) <= '0';
    layer0_outputs(5643) <= not(inputs(62));
    layer0_outputs(5644) <= not((inputs(220)) or (inputs(95)));
    layer0_outputs(5645) <= (inputs(189)) or (inputs(187));
    layer0_outputs(5646) <= not(inputs(119));
    layer0_outputs(5647) <= (inputs(237)) or (inputs(193));
    layer0_outputs(5648) <= (inputs(212)) xor (inputs(108));
    layer0_outputs(5649) <= not(inputs(142));
    layer0_outputs(5650) <= (inputs(63)) or (inputs(87));
    layer0_outputs(5651) <= (inputs(3)) xor (inputs(46));
    layer0_outputs(5652) <= (inputs(81)) or (inputs(154));
    layer0_outputs(5653) <= (inputs(78)) and not (inputs(239));
    layer0_outputs(5654) <= '0';
    layer0_outputs(5655) <= not((inputs(79)) or (inputs(146)));
    layer0_outputs(5656) <= (inputs(53)) and not (inputs(223));
    layer0_outputs(5657) <= inputs(113);
    layer0_outputs(5658) <= inputs(158);
    layer0_outputs(5659) <= inputs(210);
    layer0_outputs(5660) <= not((inputs(143)) or (inputs(161)));
    layer0_outputs(5661) <= not((inputs(244)) or (inputs(225)));
    layer0_outputs(5662) <= (inputs(114)) or (inputs(104));
    layer0_outputs(5663) <= not(inputs(131));
    layer0_outputs(5664) <= (inputs(101)) and not (inputs(160));
    layer0_outputs(5665) <= '1';
    layer0_outputs(5666) <= not((inputs(67)) xor (inputs(252)));
    layer0_outputs(5667) <= not(inputs(56));
    layer0_outputs(5668) <= (inputs(66)) or (inputs(62));
    layer0_outputs(5669) <= (inputs(242)) and (inputs(169));
    layer0_outputs(5670) <= (inputs(176)) or (inputs(229));
    layer0_outputs(5671) <= (inputs(167)) and not (inputs(239));
    layer0_outputs(5672) <= not(inputs(19));
    layer0_outputs(5673) <= (inputs(39)) and not (inputs(251));
    layer0_outputs(5674) <= not((inputs(145)) or (inputs(79)));
    layer0_outputs(5675) <= (inputs(130)) and not (inputs(49));
    layer0_outputs(5676) <= not(inputs(13));
    layer0_outputs(5677) <= not(inputs(216));
    layer0_outputs(5678) <= not((inputs(1)) or (inputs(198)));
    layer0_outputs(5679) <= inputs(118);
    layer0_outputs(5680) <= not(inputs(11));
    layer0_outputs(5681) <= (inputs(166)) and not (inputs(10));
    layer0_outputs(5682) <= not((inputs(85)) or (inputs(246)));
    layer0_outputs(5683) <= not((inputs(79)) or (inputs(211)));
    layer0_outputs(5684) <= not((inputs(182)) or (inputs(51)));
    layer0_outputs(5685) <= not(inputs(207)) or (inputs(141));
    layer0_outputs(5686) <= (inputs(133)) xor (inputs(186));
    layer0_outputs(5687) <= not(inputs(83));
    layer0_outputs(5688) <= not(inputs(57));
    layer0_outputs(5689) <= not(inputs(152));
    layer0_outputs(5690) <= not(inputs(165));
    layer0_outputs(5691) <= (inputs(56)) and (inputs(61));
    layer0_outputs(5692) <= (inputs(95)) or (inputs(23));
    layer0_outputs(5693) <= not((inputs(247)) and (inputs(216)));
    layer0_outputs(5694) <= inputs(216);
    layer0_outputs(5695) <= not((inputs(219)) xor (inputs(88)));
    layer0_outputs(5696) <= (inputs(140)) and not (inputs(37));
    layer0_outputs(5697) <= not(inputs(140));
    layer0_outputs(5698) <= not(inputs(95));
    layer0_outputs(5699) <= not(inputs(10)) or (inputs(159));
    layer0_outputs(5700) <= (inputs(133)) and not (inputs(136));
    layer0_outputs(5701) <= '1';
    layer0_outputs(5702) <= not(inputs(152));
    layer0_outputs(5703) <= (inputs(73)) or (inputs(73));
    layer0_outputs(5704) <= not(inputs(78)) or (inputs(175));
    layer0_outputs(5705) <= (inputs(154)) or (inputs(50));
    layer0_outputs(5706) <= not(inputs(124)) or (inputs(226));
    layer0_outputs(5707) <= (inputs(160)) or (inputs(190));
    layer0_outputs(5708) <= not((inputs(52)) or (inputs(247)));
    layer0_outputs(5709) <= not(inputs(43));
    layer0_outputs(5710) <= inputs(164);
    layer0_outputs(5711) <= not(inputs(106)) or (inputs(87));
    layer0_outputs(5712) <= inputs(43);
    layer0_outputs(5713) <= (inputs(87)) xor (inputs(47));
    layer0_outputs(5714) <= (inputs(153)) or (inputs(83));
    layer0_outputs(5715) <= (inputs(202)) xor (inputs(253));
    layer0_outputs(5716) <= (inputs(249)) and not (inputs(77));
    layer0_outputs(5717) <= (inputs(10)) and not (inputs(180));
    layer0_outputs(5718) <= inputs(237);
    layer0_outputs(5719) <= (inputs(79)) or (inputs(62));
    layer0_outputs(5720) <= not((inputs(109)) or (inputs(218)));
    layer0_outputs(5721) <= not(inputs(78));
    layer0_outputs(5722) <= not((inputs(48)) or (inputs(253)));
    layer0_outputs(5723) <= inputs(123);
    layer0_outputs(5724) <= not(inputs(153));
    layer0_outputs(5725) <= inputs(72);
    layer0_outputs(5726) <= (inputs(136)) and not (inputs(219));
    layer0_outputs(5727) <= (inputs(130)) and not (inputs(241));
    layer0_outputs(5728) <= '1';
    layer0_outputs(5729) <= (inputs(240)) and (inputs(195));
    layer0_outputs(5730) <= not((inputs(253)) or (inputs(95)));
    layer0_outputs(5731) <= '1';
    layer0_outputs(5732) <= inputs(87);
    layer0_outputs(5733) <= (inputs(133)) or (inputs(84));
    layer0_outputs(5734) <= not(inputs(27));
    layer0_outputs(5735) <= not((inputs(86)) or (inputs(218)));
    layer0_outputs(5736) <= not(inputs(120));
    layer0_outputs(5737) <= not(inputs(89));
    layer0_outputs(5738) <= inputs(232);
    layer0_outputs(5739) <= not(inputs(252));
    layer0_outputs(5740) <= not(inputs(118)) or (inputs(109));
    layer0_outputs(5741) <= not(inputs(149)) or (inputs(63));
    layer0_outputs(5742) <= not((inputs(54)) or (inputs(84)));
    layer0_outputs(5743) <= inputs(232);
    layer0_outputs(5744) <= inputs(166);
    layer0_outputs(5745) <= not((inputs(232)) and (inputs(107)));
    layer0_outputs(5746) <= (inputs(60)) or (inputs(48));
    layer0_outputs(5747) <= inputs(76);
    layer0_outputs(5748) <= (inputs(51)) or (inputs(98));
    layer0_outputs(5749) <= (inputs(41)) or (inputs(78));
    layer0_outputs(5750) <= not(inputs(123)) or (inputs(20));
    layer0_outputs(5751) <= not((inputs(121)) and (inputs(136)));
    layer0_outputs(5752) <= inputs(61);
    layer0_outputs(5753) <= (inputs(190)) or (inputs(70));
    layer0_outputs(5754) <= not((inputs(251)) or (inputs(201)));
    layer0_outputs(5755) <= (inputs(225)) or (inputs(160));
    layer0_outputs(5756) <= (inputs(140)) xor (inputs(207));
    layer0_outputs(5757) <= not(inputs(100));
    layer0_outputs(5758) <= not((inputs(236)) or (inputs(19)));
    layer0_outputs(5759) <= (inputs(150)) or (inputs(137));
    layer0_outputs(5760) <= not(inputs(165));
    layer0_outputs(5761) <= (inputs(237)) and not (inputs(143));
    layer0_outputs(5762) <= not(inputs(206));
    layer0_outputs(5763) <= (inputs(168)) and not (inputs(79));
    layer0_outputs(5764) <= not(inputs(106)) or (inputs(79));
    layer0_outputs(5765) <= not(inputs(215));
    layer0_outputs(5766) <= not((inputs(127)) or (inputs(86)));
    layer0_outputs(5767) <= not((inputs(24)) or (inputs(62)));
    layer0_outputs(5768) <= not(inputs(109)) or (inputs(191));
    layer0_outputs(5769) <= not(inputs(110));
    layer0_outputs(5770) <= (inputs(93)) and not (inputs(223));
    layer0_outputs(5771) <= inputs(21);
    layer0_outputs(5772) <= not((inputs(203)) or (inputs(234)));
    layer0_outputs(5773) <= not(inputs(126)) or (inputs(239));
    layer0_outputs(5774) <= (inputs(195)) and not (inputs(9));
    layer0_outputs(5775) <= not((inputs(77)) xor (inputs(151)));
    layer0_outputs(5776) <= (inputs(188)) xor (inputs(61));
    layer0_outputs(5777) <= not((inputs(221)) xor (inputs(10)));
    layer0_outputs(5778) <= not(inputs(68));
    layer0_outputs(5779) <= (inputs(150)) and not (inputs(160));
    layer0_outputs(5780) <= inputs(52);
    layer0_outputs(5781) <= inputs(167);
    layer0_outputs(5782) <= not(inputs(91));
    layer0_outputs(5783) <= (inputs(188)) and not (inputs(61));
    layer0_outputs(5784) <= (inputs(182)) or (inputs(255));
    layer0_outputs(5785) <= not(inputs(57));
    layer0_outputs(5786) <= inputs(130);
    layer0_outputs(5787) <= not(inputs(168)) or (inputs(37));
    layer0_outputs(5788) <= not(inputs(209));
    layer0_outputs(5789) <= inputs(58);
    layer0_outputs(5790) <= (inputs(231)) and not (inputs(17));
    layer0_outputs(5791) <= inputs(25);
    layer0_outputs(5792) <= not((inputs(65)) or (inputs(149)));
    layer0_outputs(5793) <= (inputs(224)) or (inputs(121));
    layer0_outputs(5794) <= not(inputs(119));
    layer0_outputs(5795) <= (inputs(10)) xor (inputs(75));
    layer0_outputs(5796) <= not(inputs(121));
    layer0_outputs(5797) <= not((inputs(211)) or (inputs(198)));
    layer0_outputs(5798) <= (inputs(28)) xor (inputs(56));
    layer0_outputs(5799) <= inputs(55);
    layer0_outputs(5800) <= not((inputs(30)) or (inputs(195)));
    layer0_outputs(5801) <= inputs(164);
    layer0_outputs(5802) <= (inputs(50)) or (inputs(84));
    layer0_outputs(5803) <= (inputs(221)) xor (inputs(242));
    layer0_outputs(5804) <= not(inputs(115));
    layer0_outputs(5805) <= (inputs(53)) xor (inputs(49));
    layer0_outputs(5806) <= '0';
    layer0_outputs(5807) <= not((inputs(248)) or (inputs(213)));
    layer0_outputs(5808) <= inputs(167);
    layer0_outputs(5809) <= not((inputs(61)) xor (inputs(127)));
    layer0_outputs(5810) <= not(inputs(211));
    layer0_outputs(5811) <= not(inputs(198));
    layer0_outputs(5812) <= not(inputs(212));
    layer0_outputs(5813) <= not((inputs(172)) xor (inputs(23)));
    layer0_outputs(5814) <= not(inputs(238));
    layer0_outputs(5815) <= not(inputs(132)) or (inputs(208));
    layer0_outputs(5816) <= not(inputs(1));
    layer0_outputs(5817) <= inputs(164);
    layer0_outputs(5818) <= inputs(130);
    layer0_outputs(5819) <= not((inputs(187)) or (inputs(207)));
    layer0_outputs(5820) <= not((inputs(109)) xor (inputs(27)));
    layer0_outputs(5821) <= not(inputs(251));
    layer0_outputs(5822) <= inputs(129);
    layer0_outputs(5823) <= inputs(104);
    layer0_outputs(5824) <= not((inputs(167)) or (inputs(57)));
    layer0_outputs(5825) <= (inputs(15)) or (inputs(155));
    layer0_outputs(5826) <= not(inputs(214));
    layer0_outputs(5827) <= inputs(98);
    layer0_outputs(5828) <= inputs(7);
    layer0_outputs(5829) <= not(inputs(243));
    layer0_outputs(5830) <= (inputs(229)) xor (inputs(236));
    layer0_outputs(5831) <= inputs(11);
    layer0_outputs(5832) <= not(inputs(118));
    layer0_outputs(5833) <= not(inputs(228));
    layer0_outputs(5834) <= (inputs(183)) or (inputs(102));
    layer0_outputs(5835) <= inputs(135);
    layer0_outputs(5836) <= not(inputs(100));
    layer0_outputs(5837) <= not((inputs(40)) or (inputs(142)));
    layer0_outputs(5838) <= inputs(88);
    layer0_outputs(5839) <= not((inputs(108)) xor (inputs(44)));
    layer0_outputs(5840) <= (inputs(72)) and not (inputs(128));
    layer0_outputs(5841) <= not(inputs(109));
    layer0_outputs(5842) <= (inputs(217)) xor (inputs(171));
    layer0_outputs(5843) <= inputs(200);
    layer0_outputs(5844) <= (inputs(66)) xor (inputs(227));
    layer0_outputs(5845) <= not((inputs(19)) or (inputs(237)));
    layer0_outputs(5846) <= not(inputs(62)) or (inputs(175));
    layer0_outputs(5847) <= not((inputs(163)) or (inputs(167)));
    layer0_outputs(5848) <= not((inputs(190)) or (inputs(172)));
    layer0_outputs(5849) <= not(inputs(43));
    layer0_outputs(5850) <= not((inputs(142)) or (inputs(39)));
    layer0_outputs(5851) <= inputs(89);
    layer0_outputs(5852) <= (inputs(179)) and not (inputs(143));
    layer0_outputs(5853) <= not(inputs(230)) or (inputs(156));
    layer0_outputs(5854) <= not(inputs(244)) or (inputs(223));
    layer0_outputs(5855) <= not(inputs(198));
    layer0_outputs(5856) <= not((inputs(88)) xor (inputs(103)));
    layer0_outputs(5857) <= inputs(113);
    layer0_outputs(5858) <= not((inputs(120)) or (inputs(79)));
    layer0_outputs(5859) <= not(inputs(212));
    layer0_outputs(5860) <= not((inputs(124)) or (inputs(5)));
    layer0_outputs(5861) <= inputs(135);
    layer0_outputs(5862) <= not(inputs(189));
    layer0_outputs(5863) <= (inputs(133)) or (inputs(139));
    layer0_outputs(5864) <= inputs(152);
    layer0_outputs(5865) <= (inputs(14)) or (inputs(154));
    layer0_outputs(5866) <= not(inputs(183));
    layer0_outputs(5867) <= (inputs(49)) or (inputs(62));
    layer0_outputs(5868) <= not((inputs(30)) xor (inputs(213)));
    layer0_outputs(5869) <= not(inputs(202)) or (inputs(70));
    layer0_outputs(5870) <= (inputs(188)) and not (inputs(244));
    layer0_outputs(5871) <= not(inputs(14));
    layer0_outputs(5872) <= (inputs(47)) and not (inputs(107));
    layer0_outputs(5873) <= not((inputs(5)) or (inputs(217)));
    layer0_outputs(5874) <= not(inputs(220)) or (inputs(68));
    layer0_outputs(5875) <= not((inputs(210)) or (inputs(41)));
    layer0_outputs(5876) <= (inputs(193)) or (inputs(241));
    layer0_outputs(5877) <= (inputs(179)) or (inputs(177));
    layer0_outputs(5878) <= not((inputs(223)) or (inputs(122)));
    layer0_outputs(5879) <= inputs(157);
    layer0_outputs(5880) <= inputs(107);
    layer0_outputs(5881) <= inputs(245);
    layer0_outputs(5882) <= not(inputs(91)) or (inputs(65));
    layer0_outputs(5883) <= (inputs(84)) and not (inputs(233));
    layer0_outputs(5884) <= not((inputs(40)) and (inputs(153)));
    layer0_outputs(5885) <= inputs(161);
    layer0_outputs(5886) <= (inputs(173)) and not (inputs(253));
    layer0_outputs(5887) <= inputs(168);
    layer0_outputs(5888) <= not(inputs(164));
    layer0_outputs(5889) <= not(inputs(118));
    layer0_outputs(5890) <= not(inputs(6)) or (inputs(240));
    layer0_outputs(5891) <= not(inputs(166));
    layer0_outputs(5892) <= (inputs(132)) and not (inputs(90));
    layer0_outputs(5893) <= not(inputs(137));
    layer0_outputs(5894) <= (inputs(249)) xor (inputs(160));
    layer0_outputs(5895) <= (inputs(43)) xor (inputs(92));
    layer0_outputs(5896) <= (inputs(73)) or (inputs(100));
    layer0_outputs(5897) <= not((inputs(121)) or (inputs(120)));
    layer0_outputs(5898) <= (inputs(44)) xor (inputs(131));
    layer0_outputs(5899) <= not(inputs(255));
    layer0_outputs(5900) <= inputs(73);
    layer0_outputs(5901) <= '0';
    layer0_outputs(5902) <= inputs(206);
    layer0_outputs(5903) <= not(inputs(136)) or (inputs(35));
    layer0_outputs(5904) <= not(inputs(214)) or (inputs(46));
    layer0_outputs(5905) <= not(inputs(117)) or (inputs(213));
    layer0_outputs(5906) <= (inputs(154)) xor (inputs(129));
    layer0_outputs(5907) <= (inputs(144)) or (inputs(230));
    layer0_outputs(5908) <= (inputs(171)) and not (inputs(15));
    layer0_outputs(5909) <= '0';
    layer0_outputs(5910) <= inputs(24);
    layer0_outputs(5911) <= not((inputs(172)) xor (inputs(106)));
    layer0_outputs(5912) <= not(inputs(189));
    layer0_outputs(5913) <= (inputs(127)) and not (inputs(221));
    layer0_outputs(5914) <= (inputs(233)) xor (inputs(100));
    layer0_outputs(5915) <= (inputs(40)) and not (inputs(194));
    layer0_outputs(5916) <= not(inputs(15));
    layer0_outputs(5917) <= inputs(219);
    layer0_outputs(5918) <= inputs(34);
    layer0_outputs(5919) <= (inputs(7)) and not (inputs(236));
    layer0_outputs(5920) <= not(inputs(236)) or (inputs(73));
    layer0_outputs(5921) <= not((inputs(11)) or (inputs(122)));
    layer0_outputs(5922) <= not(inputs(152)) or (inputs(159));
    layer0_outputs(5923) <= (inputs(197)) and not (inputs(238));
    layer0_outputs(5924) <= not((inputs(253)) or (inputs(74)));
    layer0_outputs(5925) <= (inputs(121)) or (inputs(122));
    layer0_outputs(5926) <= not(inputs(155)) or (inputs(181));
    layer0_outputs(5927) <= inputs(165);
    layer0_outputs(5928) <= not((inputs(157)) or (inputs(246)));
    layer0_outputs(5929) <= (inputs(246)) xor (inputs(234));
    layer0_outputs(5930) <= not(inputs(148)) or (inputs(64));
    layer0_outputs(5931) <= not((inputs(201)) xor (inputs(138)));
    layer0_outputs(5932) <= inputs(235);
    layer0_outputs(5933) <= not(inputs(124));
    layer0_outputs(5934) <= not(inputs(39)) or (inputs(14));
    layer0_outputs(5935) <= not(inputs(85)) or (inputs(67));
    layer0_outputs(5936) <= not((inputs(188)) xor (inputs(113)));
    layer0_outputs(5937) <= not(inputs(177));
    layer0_outputs(5938) <= inputs(159);
    layer0_outputs(5939) <= inputs(243);
    layer0_outputs(5940) <= not(inputs(169)) or (inputs(44));
    layer0_outputs(5941) <= (inputs(191)) or (inputs(222));
    layer0_outputs(5942) <= (inputs(116)) xor (inputs(148));
    layer0_outputs(5943) <= (inputs(222)) or (inputs(5));
    layer0_outputs(5944) <= (inputs(230)) and not (inputs(135));
    layer0_outputs(5945) <= not(inputs(244)) or (inputs(236));
    layer0_outputs(5946) <= (inputs(240)) and (inputs(16));
    layer0_outputs(5947) <= inputs(74);
    layer0_outputs(5948) <= not((inputs(39)) or (inputs(142)));
    layer0_outputs(5949) <= (inputs(114)) or (inputs(207));
    layer0_outputs(5950) <= not(inputs(87)) or (inputs(48));
    layer0_outputs(5951) <= not(inputs(153));
    layer0_outputs(5952) <= inputs(116);
    layer0_outputs(5953) <= not(inputs(87));
    layer0_outputs(5954) <= not((inputs(31)) xor (inputs(6)));
    layer0_outputs(5955) <= not(inputs(179)) or (inputs(238));
    layer0_outputs(5956) <= not((inputs(61)) or (inputs(73)));
    layer0_outputs(5957) <= (inputs(247)) or (inputs(179));
    layer0_outputs(5958) <= inputs(39);
    layer0_outputs(5959) <= not((inputs(147)) xor (inputs(109)));
    layer0_outputs(5960) <= not((inputs(253)) xor (inputs(195)));
    layer0_outputs(5961) <= not(inputs(128));
    layer0_outputs(5962) <= not(inputs(76)) or (inputs(119));
    layer0_outputs(5963) <= not(inputs(83)) or (inputs(186));
    layer0_outputs(5964) <= (inputs(193)) and not (inputs(111));
    layer0_outputs(5965) <= (inputs(41)) and not (inputs(253));
    layer0_outputs(5966) <= not(inputs(26));
    layer0_outputs(5967) <= inputs(176);
    layer0_outputs(5968) <= not(inputs(19)) or (inputs(155));
    layer0_outputs(5969) <= inputs(146);
    layer0_outputs(5970) <= not((inputs(48)) and (inputs(104)));
    layer0_outputs(5971) <= (inputs(55)) or (inputs(191));
    layer0_outputs(5972) <= not(inputs(253)) or (inputs(52));
    layer0_outputs(5973) <= (inputs(25)) or (inputs(124));
    layer0_outputs(5974) <= (inputs(214)) and not (inputs(17));
    layer0_outputs(5975) <= (inputs(24)) or (inputs(204));
    layer0_outputs(5976) <= (inputs(33)) or (inputs(4));
    layer0_outputs(5977) <= '1';
    layer0_outputs(5978) <= (inputs(115)) or (inputs(154));
    layer0_outputs(5979) <= (inputs(42)) and not (inputs(136));
    layer0_outputs(5980) <= (inputs(151)) and not (inputs(171));
    layer0_outputs(5981) <= inputs(43);
    layer0_outputs(5982) <= (inputs(170)) and not (inputs(247));
    layer0_outputs(5983) <= not((inputs(204)) xor (inputs(132)));
    layer0_outputs(5984) <= (inputs(22)) xor (inputs(126));
    layer0_outputs(5985) <= inputs(228);
    layer0_outputs(5986) <= (inputs(151)) and not (inputs(62));
    layer0_outputs(5987) <= not(inputs(23));
    layer0_outputs(5988) <= inputs(210);
    layer0_outputs(5989) <= not((inputs(250)) or (inputs(120)));
    layer0_outputs(5990) <= not(inputs(104));
    layer0_outputs(5991) <= not(inputs(199)) or (inputs(188));
    layer0_outputs(5992) <= inputs(44);
    layer0_outputs(5993) <= (inputs(204)) and not (inputs(14));
    layer0_outputs(5994) <= not(inputs(158));
    layer0_outputs(5995) <= not(inputs(121)) or (inputs(78));
    layer0_outputs(5996) <= not(inputs(120)) or (inputs(119));
    layer0_outputs(5997) <= (inputs(132)) and not (inputs(190));
    layer0_outputs(5998) <= not(inputs(165)) or (inputs(100));
    layer0_outputs(5999) <= not(inputs(182)) or (inputs(1));
    layer0_outputs(6000) <= (inputs(152)) and (inputs(138));
    layer0_outputs(6001) <= inputs(37);
    layer0_outputs(6002) <= inputs(159);
    layer0_outputs(6003) <= not((inputs(70)) or (inputs(113)));
    layer0_outputs(6004) <= not((inputs(126)) or (inputs(22)));
    layer0_outputs(6005) <= not(inputs(45));
    layer0_outputs(6006) <= inputs(93);
    layer0_outputs(6007) <= (inputs(174)) and (inputs(55));
    layer0_outputs(6008) <= (inputs(108)) or (inputs(140));
    layer0_outputs(6009) <= not((inputs(184)) and (inputs(248)));
    layer0_outputs(6010) <= not(inputs(93));
    layer0_outputs(6011) <= inputs(68);
    layer0_outputs(6012) <= (inputs(236)) xor (inputs(151));
    layer0_outputs(6013) <= (inputs(83)) and not (inputs(16));
    layer0_outputs(6014) <= not(inputs(204));
    layer0_outputs(6015) <= not(inputs(142));
    layer0_outputs(6016) <= not(inputs(204)) or (inputs(212));
    layer0_outputs(6017) <= not(inputs(162)) or (inputs(165));
    layer0_outputs(6018) <= inputs(4);
    layer0_outputs(6019) <= inputs(21);
    layer0_outputs(6020) <= not((inputs(130)) or (inputs(172)));
    layer0_outputs(6021) <= inputs(195);
    layer0_outputs(6022) <= (inputs(103)) and not (inputs(145));
    layer0_outputs(6023) <= not((inputs(175)) xor (inputs(17)));
    layer0_outputs(6024) <= inputs(110);
    layer0_outputs(6025) <= not((inputs(35)) or (inputs(111)));
    layer0_outputs(6026) <= not((inputs(145)) or (inputs(169)));
    layer0_outputs(6027) <= '0';
    layer0_outputs(6028) <= not(inputs(102)) or (inputs(92));
    layer0_outputs(6029) <= (inputs(223)) or (inputs(18));
    layer0_outputs(6030) <= (inputs(33)) or (inputs(5));
    layer0_outputs(6031) <= not(inputs(197)) or (inputs(53));
    layer0_outputs(6032) <= (inputs(176)) or (inputs(59));
    layer0_outputs(6033) <= (inputs(251)) and not (inputs(144));
    layer0_outputs(6034) <= inputs(24);
    layer0_outputs(6035) <= not(inputs(109));
    layer0_outputs(6036) <= (inputs(185)) xor (inputs(122));
    layer0_outputs(6037) <= not((inputs(161)) xor (inputs(119)));
    layer0_outputs(6038) <= (inputs(114)) xor (inputs(19));
    layer0_outputs(6039) <= not(inputs(108)) or (inputs(235));
    layer0_outputs(6040) <= '0';
    layer0_outputs(6041) <= inputs(209);
    layer0_outputs(6042) <= inputs(132);
    layer0_outputs(6043) <= inputs(37);
    layer0_outputs(6044) <= (inputs(97)) or (inputs(255));
    layer0_outputs(6045) <= not(inputs(57)) or (inputs(160));
    layer0_outputs(6046) <= inputs(25);
    layer0_outputs(6047) <= (inputs(0)) or (inputs(3));
    layer0_outputs(6048) <= (inputs(61)) and not (inputs(14));
    layer0_outputs(6049) <= (inputs(58)) xor (inputs(75));
    layer0_outputs(6050) <= (inputs(215)) or (inputs(114));
    layer0_outputs(6051) <= '0';
    layer0_outputs(6052) <= not(inputs(140));
    layer0_outputs(6053) <= inputs(103);
    layer0_outputs(6054) <= not((inputs(203)) or (inputs(187)));
    layer0_outputs(6055) <= not(inputs(10)) or (inputs(176));
    layer0_outputs(6056) <= (inputs(242)) xor (inputs(119));
    layer0_outputs(6057) <= not(inputs(59));
    layer0_outputs(6058) <= (inputs(71)) or (inputs(50));
    layer0_outputs(6059) <= not(inputs(149)) or (inputs(21));
    layer0_outputs(6060) <= (inputs(135)) and not (inputs(36));
    layer0_outputs(6061) <= inputs(78);
    layer0_outputs(6062) <= (inputs(169)) and not (inputs(176));
    layer0_outputs(6063) <= not(inputs(125)) or (inputs(50));
    layer0_outputs(6064) <= not(inputs(58));
    layer0_outputs(6065) <= not(inputs(107));
    layer0_outputs(6066) <= (inputs(215)) xor (inputs(127));
    layer0_outputs(6067) <= (inputs(27)) and not (inputs(87));
    layer0_outputs(6068) <= not(inputs(99));
    layer0_outputs(6069) <= not(inputs(96));
    layer0_outputs(6070) <= not((inputs(244)) or (inputs(227)));
    layer0_outputs(6071) <= not((inputs(46)) xor (inputs(68)));
    layer0_outputs(6072) <= not((inputs(203)) or (inputs(112)));
    layer0_outputs(6073) <= not(inputs(211));
    layer0_outputs(6074) <= (inputs(175)) xor (inputs(171));
    layer0_outputs(6075) <= inputs(94);
    layer0_outputs(6076) <= (inputs(176)) or (inputs(214));
    layer0_outputs(6077) <= (inputs(54)) or (inputs(145));
    layer0_outputs(6078) <= not(inputs(32));
    layer0_outputs(6079) <= not(inputs(146));
    layer0_outputs(6080) <= not((inputs(115)) or (inputs(190)));
    layer0_outputs(6081) <= not(inputs(37)) or (inputs(211));
    layer0_outputs(6082) <= inputs(30);
    layer0_outputs(6083) <= (inputs(158)) and (inputs(47));
    layer0_outputs(6084) <= inputs(82);
    layer0_outputs(6085) <= not((inputs(184)) or (inputs(15)));
    layer0_outputs(6086) <= not(inputs(165));
    layer0_outputs(6087) <= not(inputs(34));
    layer0_outputs(6088) <= (inputs(229)) xor (inputs(183));
    layer0_outputs(6089) <= (inputs(246)) and not (inputs(47));
    layer0_outputs(6090) <= (inputs(6)) or (inputs(10));
    layer0_outputs(6091) <= not(inputs(117)) or (inputs(192));
    layer0_outputs(6092) <= not((inputs(247)) xor (inputs(78)));
    layer0_outputs(6093) <= not((inputs(15)) or (inputs(124)));
    layer0_outputs(6094) <= (inputs(219)) or (inputs(174));
    layer0_outputs(6095) <= not(inputs(167)) or (inputs(111));
    layer0_outputs(6096) <= not((inputs(175)) or (inputs(126)));
    layer0_outputs(6097) <= not((inputs(232)) and (inputs(166)));
    layer0_outputs(6098) <= (inputs(211)) xor (inputs(138));
    layer0_outputs(6099) <= not(inputs(161));
    layer0_outputs(6100) <= inputs(142);
    layer0_outputs(6101) <= (inputs(38)) and not (inputs(94));
    layer0_outputs(6102) <= (inputs(229)) and not (inputs(41));
    layer0_outputs(6103) <= (inputs(133)) or (inputs(146));
    layer0_outputs(6104) <= (inputs(197)) xor (inputs(232));
    layer0_outputs(6105) <= not(inputs(52));
    layer0_outputs(6106) <= (inputs(103)) and not (inputs(85));
    layer0_outputs(6107) <= not(inputs(50));
    layer0_outputs(6108) <= not(inputs(178));
    layer0_outputs(6109) <= not(inputs(36)) or (inputs(72));
    layer0_outputs(6110) <= not(inputs(74));
    layer0_outputs(6111) <= not(inputs(117)) or (inputs(127));
    layer0_outputs(6112) <= inputs(125);
    layer0_outputs(6113) <= not(inputs(152));
    layer0_outputs(6114) <= (inputs(139)) xor (inputs(74));
    layer0_outputs(6115) <= inputs(8);
    layer0_outputs(6116) <= inputs(166);
    layer0_outputs(6117) <= not((inputs(68)) and (inputs(133)));
    layer0_outputs(6118) <= (inputs(158)) or (inputs(100));
    layer0_outputs(6119) <= not(inputs(203)) or (inputs(222));
    layer0_outputs(6120) <= inputs(36);
    layer0_outputs(6121) <= not(inputs(247));
    layer0_outputs(6122) <= not((inputs(33)) xor (inputs(64)));
    layer0_outputs(6123) <= (inputs(230)) and not (inputs(130));
    layer0_outputs(6124) <= (inputs(196)) xor (inputs(154));
    layer0_outputs(6125) <= not((inputs(47)) or (inputs(215)));
    layer0_outputs(6126) <= not((inputs(73)) or (inputs(244)));
    layer0_outputs(6127) <= not(inputs(183)) or (inputs(120));
    layer0_outputs(6128) <= not((inputs(183)) or (inputs(128)));
    layer0_outputs(6129) <= not(inputs(139));
    layer0_outputs(6130) <= inputs(106);
    layer0_outputs(6131) <= inputs(170);
    layer0_outputs(6132) <= not(inputs(151));
    layer0_outputs(6133) <= not(inputs(72));
    layer0_outputs(6134) <= not(inputs(19)) or (inputs(112));
    layer0_outputs(6135) <= inputs(198);
    layer0_outputs(6136) <= not((inputs(99)) or (inputs(225)));
    layer0_outputs(6137) <= not((inputs(62)) or (inputs(123)));
    layer0_outputs(6138) <= not((inputs(33)) or (inputs(192)));
    layer0_outputs(6139) <= not((inputs(71)) xor (inputs(121)));
    layer0_outputs(6140) <= not(inputs(116));
    layer0_outputs(6141) <= (inputs(244)) or (inputs(187));
    layer0_outputs(6142) <= not(inputs(75)) or (inputs(47));
    layer0_outputs(6143) <= not((inputs(88)) xor (inputs(22)));
    layer0_outputs(6144) <= inputs(105);
    layer0_outputs(6145) <= not(inputs(152)) or (inputs(177));
    layer0_outputs(6146) <= (inputs(90)) or (inputs(241));
    layer0_outputs(6147) <= not(inputs(37));
    layer0_outputs(6148) <= not((inputs(127)) or (inputs(40)));
    layer0_outputs(6149) <= not(inputs(214));
    layer0_outputs(6150) <= (inputs(56)) or (inputs(71));
    layer0_outputs(6151) <= (inputs(10)) and (inputs(182));
    layer0_outputs(6152) <= inputs(178);
    layer0_outputs(6153) <= not(inputs(98)) or (inputs(123));
    layer0_outputs(6154) <= (inputs(180)) and not (inputs(116));
    layer0_outputs(6155) <= not(inputs(183));
    layer0_outputs(6156) <= (inputs(229)) and not (inputs(92));
    layer0_outputs(6157) <= (inputs(69)) or (inputs(211));
    layer0_outputs(6158) <= not((inputs(236)) xor (inputs(20)));
    layer0_outputs(6159) <= not(inputs(18));
    layer0_outputs(6160) <= (inputs(247)) and (inputs(139));
    layer0_outputs(6161) <= (inputs(175)) or (inputs(226));
    layer0_outputs(6162) <= (inputs(172)) and not (inputs(64));
    layer0_outputs(6163) <= not(inputs(184)) or (inputs(238));
    layer0_outputs(6164) <= not(inputs(207)) or (inputs(236));
    layer0_outputs(6165) <= not(inputs(218)) or (inputs(53));
    layer0_outputs(6166) <= inputs(241);
    layer0_outputs(6167) <= not(inputs(232));
    layer0_outputs(6168) <= not(inputs(107));
    layer0_outputs(6169) <= not((inputs(13)) xor (inputs(31)));
    layer0_outputs(6170) <= (inputs(161)) or (inputs(12));
    layer0_outputs(6171) <= inputs(165);
    layer0_outputs(6172) <= inputs(135);
    layer0_outputs(6173) <= inputs(182);
    layer0_outputs(6174) <= not(inputs(58));
    layer0_outputs(6175) <= inputs(127);
    layer0_outputs(6176) <= not(inputs(216));
    layer0_outputs(6177) <= (inputs(56)) and not (inputs(56));
    layer0_outputs(6178) <= inputs(189);
    layer0_outputs(6179) <= inputs(230);
    layer0_outputs(6180) <= inputs(167);
    layer0_outputs(6181) <= not(inputs(226));
    layer0_outputs(6182) <= not(inputs(177));
    layer0_outputs(6183) <= (inputs(97)) and not (inputs(32));
    layer0_outputs(6184) <= (inputs(145)) or (inputs(225));
    layer0_outputs(6185) <= not(inputs(149)) or (inputs(74));
    layer0_outputs(6186) <= (inputs(63)) xor (inputs(47));
    layer0_outputs(6187) <= not((inputs(169)) or (inputs(97)));
    layer0_outputs(6188) <= not(inputs(164)) or (inputs(127));
    layer0_outputs(6189) <= (inputs(142)) or (inputs(125));
    layer0_outputs(6190) <= not(inputs(16));
    layer0_outputs(6191) <= inputs(70);
    layer0_outputs(6192) <= (inputs(96)) and not (inputs(96));
    layer0_outputs(6193) <= not(inputs(196)) or (inputs(46));
    layer0_outputs(6194) <= (inputs(126)) or (inputs(21));
    layer0_outputs(6195) <= not(inputs(90));
    layer0_outputs(6196) <= (inputs(55)) and not (inputs(29));
    layer0_outputs(6197) <= (inputs(115)) or (inputs(101));
    layer0_outputs(6198) <= not((inputs(186)) or (inputs(124)));
    layer0_outputs(6199) <= inputs(83);
    layer0_outputs(6200) <= inputs(40);
    layer0_outputs(6201) <= not(inputs(138));
    layer0_outputs(6202) <= (inputs(212)) and not (inputs(76));
    layer0_outputs(6203) <= not(inputs(215));
    layer0_outputs(6204) <= not((inputs(172)) xor (inputs(121)));
    layer0_outputs(6205) <= (inputs(154)) or (inputs(254));
    layer0_outputs(6206) <= not((inputs(3)) or (inputs(74)));
    layer0_outputs(6207) <= (inputs(222)) or (inputs(5));
    layer0_outputs(6208) <= inputs(75);
    layer0_outputs(6209) <= not((inputs(73)) xor (inputs(118)));
    layer0_outputs(6210) <= not(inputs(123)) or (inputs(81));
    layer0_outputs(6211) <= not(inputs(7)) or (inputs(112));
    layer0_outputs(6212) <= (inputs(135)) and (inputs(38));
    layer0_outputs(6213) <= (inputs(116)) or (inputs(162));
    layer0_outputs(6214) <= not((inputs(176)) or (inputs(165)));
    layer0_outputs(6215) <= inputs(70);
    layer0_outputs(6216) <= inputs(87);
    layer0_outputs(6217) <= (inputs(198)) or (inputs(144));
    layer0_outputs(6218) <= (inputs(72)) and not (inputs(253));
    layer0_outputs(6219) <= (inputs(207)) or (inputs(234));
    layer0_outputs(6220) <= not((inputs(182)) or (inputs(237)));
    layer0_outputs(6221) <= not((inputs(115)) or (inputs(132)));
    layer0_outputs(6222) <= (inputs(43)) or (inputs(34));
    layer0_outputs(6223) <= not(inputs(154));
    layer0_outputs(6224) <= not(inputs(85));
    layer0_outputs(6225) <= (inputs(7)) and not (inputs(212));
    layer0_outputs(6226) <= not((inputs(24)) or (inputs(69)));
    layer0_outputs(6227) <= not(inputs(58)) or (inputs(224));
    layer0_outputs(6228) <= not((inputs(206)) and (inputs(182)));
    layer0_outputs(6229) <= not(inputs(134)) or (inputs(95));
    layer0_outputs(6230) <= not((inputs(138)) xor (inputs(18)));
    layer0_outputs(6231) <= not((inputs(20)) or (inputs(185)));
    layer0_outputs(6232) <= inputs(3);
    layer0_outputs(6233) <= not((inputs(141)) or (inputs(197)));
    layer0_outputs(6234) <= not((inputs(232)) or (inputs(251)));
    layer0_outputs(6235) <= (inputs(32)) xor (inputs(75));
    layer0_outputs(6236) <= not((inputs(7)) xor (inputs(194)));
    layer0_outputs(6237) <= (inputs(252)) xor (inputs(171));
    layer0_outputs(6238) <= not(inputs(104));
    layer0_outputs(6239) <= (inputs(72)) xor (inputs(114));
    layer0_outputs(6240) <= (inputs(120)) and not (inputs(253));
    layer0_outputs(6241) <= (inputs(68)) and not (inputs(143));
    layer0_outputs(6242) <= inputs(129);
    layer0_outputs(6243) <= not(inputs(73)) or (inputs(2));
    layer0_outputs(6244) <= not((inputs(240)) xor (inputs(202)));
    layer0_outputs(6245) <= not(inputs(83));
    layer0_outputs(6246) <= inputs(67);
    layer0_outputs(6247) <= not(inputs(151));
    layer0_outputs(6248) <= (inputs(135)) or (inputs(249));
    layer0_outputs(6249) <= (inputs(13)) and not (inputs(210));
    layer0_outputs(6250) <= inputs(158);
    layer0_outputs(6251) <= (inputs(28)) and not (inputs(205));
    layer0_outputs(6252) <= (inputs(238)) or (inputs(147));
    layer0_outputs(6253) <= (inputs(211)) and not (inputs(7));
    layer0_outputs(6254) <= not(inputs(195));
    layer0_outputs(6255) <= '1';
    layer0_outputs(6256) <= not((inputs(129)) or (inputs(12)));
    layer0_outputs(6257) <= not((inputs(24)) xor (inputs(52)));
    layer0_outputs(6258) <= (inputs(198)) and not (inputs(126));
    layer0_outputs(6259) <= (inputs(76)) xor (inputs(108));
    layer0_outputs(6260) <= inputs(166);
    layer0_outputs(6261) <= not((inputs(173)) xor (inputs(198)));
    layer0_outputs(6262) <= inputs(86);
    layer0_outputs(6263) <= inputs(248);
    layer0_outputs(6264) <= not((inputs(185)) xor (inputs(248)));
    layer0_outputs(6265) <= (inputs(22)) xor (inputs(178));
    layer0_outputs(6266) <= not(inputs(218)) or (inputs(91));
    layer0_outputs(6267) <= not(inputs(57));
    layer0_outputs(6268) <= not(inputs(214)) or (inputs(36));
    layer0_outputs(6269) <= not((inputs(174)) or (inputs(22)));
    layer0_outputs(6270) <= not((inputs(169)) or (inputs(241)));
    layer0_outputs(6271) <= inputs(167);
    layer0_outputs(6272) <= not((inputs(77)) or (inputs(138)));
    layer0_outputs(6273) <= not((inputs(87)) xor (inputs(115)));
    layer0_outputs(6274) <= not((inputs(81)) or (inputs(29)));
    layer0_outputs(6275) <= inputs(189);
    layer0_outputs(6276) <= not((inputs(22)) xor (inputs(160)));
    layer0_outputs(6277) <= (inputs(50)) or (inputs(249));
    layer0_outputs(6278) <= (inputs(142)) and not (inputs(254));
    layer0_outputs(6279) <= inputs(51);
    layer0_outputs(6280) <= not((inputs(239)) or (inputs(236)));
    layer0_outputs(6281) <= (inputs(28)) or (inputs(125));
    layer0_outputs(6282) <= not(inputs(177));
    layer0_outputs(6283) <= not(inputs(170)) or (inputs(53));
    layer0_outputs(6284) <= (inputs(203)) and (inputs(243));
    layer0_outputs(6285) <= inputs(40);
    layer0_outputs(6286) <= not((inputs(23)) or (inputs(40)));
    layer0_outputs(6287) <= (inputs(10)) or (inputs(248));
    layer0_outputs(6288) <= (inputs(87)) and not (inputs(224));
    layer0_outputs(6289) <= (inputs(171)) or (inputs(128));
    layer0_outputs(6290) <= (inputs(82)) xor (inputs(45));
    layer0_outputs(6291) <= (inputs(163)) xor (inputs(165));
    layer0_outputs(6292) <= not((inputs(250)) or (inputs(133)));
    layer0_outputs(6293) <= not((inputs(209)) or (inputs(83)));
    layer0_outputs(6294) <= inputs(72);
    layer0_outputs(6295) <= not((inputs(5)) xor (inputs(64)));
    layer0_outputs(6296) <= not(inputs(182));
    layer0_outputs(6297) <= (inputs(63)) and not (inputs(112));
    layer0_outputs(6298) <= not(inputs(39));
    layer0_outputs(6299) <= not((inputs(90)) or (inputs(65)));
    layer0_outputs(6300) <= (inputs(104)) xor (inputs(238));
    layer0_outputs(6301) <= not(inputs(169)) or (inputs(84));
    layer0_outputs(6302) <= not((inputs(212)) xor (inputs(207)));
    layer0_outputs(6303) <= (inputs(209)) or (inputs(226));
    layer0_outputs(6304) <= (inputs(179)) xor (inputs(78));
    layer0_outputs(6305) <= not(inputs(104));
    layer0_outputs(6306) <= not((inputs(230)) xor (inputs(75)));
    layer0_outputs(6307) <= (inputs(34)) xor (inputs(81));
    layer0_outputs(6308) <= inputs(176);
    layer0_outputs(6309) <= not(inputs(219));
    layer0_outputs(6310) <= (inputs(205)) and not (inputs(47));
    layer0_outputs(6311) <= not(inputs(246));
    layer0_outputs(6312) <= (inputs(247)) or (inputs(177));
    layer0_outputs(6313) <= inputs(211);
    layer0_outputs(6314) <= (inputs(197)) and not (inputs(237));
    layer0_outputs(6315) <= not(inputs(197)) or (inputs(172));
    layer0_outputs(6316) <= not(inputs(155));
    layer0_outputs(6317) <= (inputs(247)) and not (inputs(51));
    layer0_outputs(6318) <= not(inputs(67)) or (inputs(29));
    layer0_outputs(6319) <= inputs(230);
    layer0_outputs(6320) <= inputs(187);
    layer0_outputs(6321) <= (inputs(64)) xor (inputs(86));
    layer0_outputs(6322) <= (inputs(51)) xor (inputs(147));
    layer0_outputs(6323) <= inputs(128);
    layer0_outputs(6324) <= inputs(92);
    layer0_outputs(6325) <= inputs(219);
    layer0_outputs(6326) <= (inputs(140)) and not (inputs(18));
    layer0_outputs(6327) <= not(inputs(115)) or (inputs(41));
    layer0_outputs(6328) <= not((inputs(60)) xor (inputs(181)));
    layer0_outputs(6329) <= (inputs(6)) and not (inputs(100));
    layer0_outputs(6330) <= not(inputs(163));
    layer0_outputs(6331) <= inputs(166);
    layer0_outputs(6332) <= not((inputs(33)) or (inputs(61)));
    layer0_outputs(6333) <= not((inputs(195)) xor (inputs(233)));
    layer0_outputs(6334) <= not(inputs(72));
    layer0_outputs(6335) <= not(inputs(119)) or (inputs(157));
    layer0_outputs(6336) <= (inputs(89)) and not (inputs(248));
    layer0_outputs(6337) <= inputs(204);
    layer0_outputs(6338) <= not(inputs(6));
    layer0_outputs(6339) <= not((inputs(173)) xor (inputs(129)));
    layer0_outputs(6340) <= (inputs(86)) and not (inputs(126));
    layer0_outputs(6341) <= not((inputs(169)) xor (inputs(199)));
    layer0_outputs(6342) <= not((inputs(72)) xor (inputs(21)));
    layer0_outputs(6343) <= not(inputs(242));
    layer0_outputs(6344) <= not((inputs(69)) xor (inputs(38)));
    layer0_outputs(6345) <= (inputs(29)) xor (inputs(45));
    layer0_outputs(6346) <= not((inputs(237)) or (inputs(252)));
    layer0_outputs(6347) <= not(inputs(82)) or (inputs(255));
    layer0_outputs(6348) <= not((inputs(105)) or (inputs(13)));
    layer0_outputs(6349) <= not(inputs(101)) or (inputs(191));
    layer0_outputs(6350) <= inputs(235);
    layer0_outputs(6351) <= (inputs(166)) or (inputs(109));
    layer0_outputs(6352) <= (inputs(57)) or (inputs(48));
    layer0_outputs(6353) <= not(inputs(251)) or (inputs(1));
    layer0_outputs(6354) <= not((inputs(169)) or (inputs(153)));
    layer0_outputs(6355) <= (inputs(177)) xor (inputs(191));
    layer0_outputs(6356) <= not(inputs(130));
    layer0_outputs(6357) <= (inputs(201)) or (inputs(189));
    layer0_outputs(6358) <= not(inputs(118)) or (inputs(32));
    layer0_outputs(6359) <= (inputs(203)) or (inputs(15));
    layer0_outputs(6360) <= not((inputs(140)) and (inputs(200)));
    layer0_outputs(6361) <= (inputs(86)) xor (inputs(190));
    layer0_outputs(6362) <= (inputs(60)) and not (inputs(86));
    layer0_outputs(6363) <= inputs(167);
    layer0_outputs(6364) <= not((inputs(21)) or (inputs(47)));
    layer0_outputs(6365) <= not(inputs(85));
    layer0_outputs(6366) <= not(inputs(207)) or (inputs(32));
    layer0_outputs(6367) <= not(inputs(8));
    layer0_outputs(6368) <= not((inputs(196)) or (inputs(93)));
    layer0_outputs(6369) <= not(inputs(115));
    layer0_outputs(6370) <= (inputs(19)) xor (inputs(91));
    layer0_outputs(6371) <= not(inputs(216)) or (inputs(82));
    layer0_outputs(6372) <= not((inputs(66)) xor (inputs(54)));
    layer0_outputs(6373) <= not((inputs(187)) and (inputs(129)));
    layer0_outputs(6374) <= inputs(177);
    layer0_outputs(6375) <= not(inputs(81)) or (inputs(127));
    layer0_outputs(6376) <= (inputs(25)) and not (inputs(112));
    layer0_outputs(6377) <= not(inputs(76));
    layer0_outputs(6378) <= inputs(187);
    layer0_outputs(6379) <= (inputs(184)) or (inputs(189));
    layer0_outputs(6380) <= not((inputs(23)) and (inputs(135)));
    layer0_outputs(6381) <= (inputs(68)) or (inputs(193));
    layer0_outputs(6382) <= not((inputs(93)) xor (inputs(17)));
    layer0_outputs(6383) <= not(inputs(69));
    layer0_outputs(6384) <= not(inputs(228)) or (inputs(88));
    layer0_outputs(6385) <= inputs(135);
    layer0_outputs(6386) <= not((inputs(140)) or (inputs(138)));
    layer0_outputs(6387) <= not(inputs(209));
    layer0_outputs(6388) <= not(inputs(232));
    layer0_outputs(6389) <= (inputs(181)) and not (inputs(32));
    layer0_outputs(6390) <= not(inputs(67)) or (inputs(103));
    layer0_outputs(6391) <= not((inputs(131)) xor (inputs(189)));
    layer0_outputs(6392) <= (inputs(10)) and (inputs(60));
    layer0_outputs(6393) <= inputs(21);
    layer0_outputs(6394) <= (inputs(252)) or (inputs(121));
    layer0_outputs(6395) <= not((inputs(209)) or (inputs(230)));
    layer0_outputs(6396) <= not((inputs(223)) or (inputs(92)));
    layer0_outputs(6397) <= not(inputs(148));
    layer0_outputs(6398) <= inputs(125);
    layer0_outputs(6399) <= not((inputs(11)) and (inputs(99)));
    layer0_outputs(6400) <= (inputs(91)) or (inputs(223));
    layer0_outputs(6401) <= (inputs(69)) and not (inputs(128));
    layer0_outputs(6402) <= not(inputs(87)) or (inputs(229));
    layer0_outputs(6403) <= inputs(229);
    layer0_outputs(6404) <= not(inputs(134));
    layer0_outputs(6405) <= inputs(105);
    layer0_outputs(6406) <= not(inputs(102));
    layer0_outputs(6407) <= not((inputs(151)) or (inputs(128)));
    layer0_outputs(6408) <= inputs(76);
    layer0_outputs(6409) <= (inputs(74)) and not (inputs(224));
    layer0_outputs(6410) <= not((inputs(64)) or (inputs(221)));
    layer0_outputs(6411) <= inputs(39);
    layer0_outputs(6412) <= (inputs(131)) or (inputs(129));
    layer0_outputs(6413) <= not(inputs(92));
    layer0_outputs(6414) <= not((inputs(108)) xor (inputs(181)));
    layer0_outputs(6415) <= (inputs(50)) xor (inputs(52));
    layer0_outputs(6416) <= not((inputs(140)) xor (inputs(171)));
    layer0_outputs(6417) <= inputs(72);
    layer0_outputs(6418) <= not(inputs(28));
    layer0_outputs(6419) <= (inputs(184)) and not (inputs(142));
    layer0_outputs(6420) <= inputs(216);
    layer0_outputs(6421) <= not(inputs(194));
    layer0_outputs(6422) <= not(inputs(148));
    layer0_outputs(6423) <= not((inputs(182)) xor (inputs(174)));
    layer0_outputs(6424) <= not((inputs(250)) or (inputs(175)));
    layer0_outputs(6425) <= not((inputs(134)) or (inputs(95)));
    layer0_outputs(6426) <= inputs(163);
    layer0_outputs(6427) <= (inputs(88)) or (inputs(132));
    layer0_outputs(6428) <= not((inputs(43)) or (inputs(170)));
    layer0_outputs(6429) <= not(inputs(247)) or (inputs(35));
    layer0_outputs(6430) <= (inputs(19)) or (inputs(38));
    layer0_outputs(6431) <= inputs(134);
    layer0_outputs(6432) <= inputs(36);
    layer0_outputs(6433) <= (inputs(167)) and not (inputs(127));
    layer0_outputs(6434) <= (inputs(252)) or (inputs(103));
    layer0_outputs(6435) <= (inputs(144)) or (inputs(70));
    layer0_outputs(6436) <= inputs(166);
    layer0_outputs(6437) <= (inputs(41)) or (inputs(61));
    layer0_outputs(6438) <= not((inputs(176)) xor (inputs(114)));
    layer0_outputs(6439) <= (inputs(25)) or (inputs(3));
    layer0_outputs(6440) <= '0';
    layer0_outputs(6441) <= not(inputs(7)) or (inputs(230));
    layer0_outputs(6442) <= (inputs(52)) and not (inputs(54));
    layer0_outputs(6443) <= not((inputs(120)) or (inputs(124)));
    layer0_outputs(6444) <= not((inputs(192)) xor (inputs(250)));
    layer0_outputs(6445) <= inputs(126);
    layer0_outputs(6446) <= inputs(130);
    layer0_outputs(6447) <= not((inputs(26)) or (inputs(80)));
    layer0_outputs(6448) <= not(inputs(97));
    layer0_outputs(6449) <= '1';
    layer0_outputs(6450) <= '0';
    layer0_outputs(6451) <= not(inputs(254));
    layer0_outputs(6452) <= inputs(105);
    layer0_outputs(6453) <= (inputs(163)) and not (inputs(152));
    layer0_outputs(6454) <= not(inputs(145)) or (inputs(253));
    layer0_outputs(6455) <= not(inputs(242));
    layer0_outputs(6456) <= (inputs(90)) or (inputs(239));
    layer0_outputs(6457) <= (inputs(255)) or (inputs(82));
    layer0_outputs(6458) <= '1';
    layer0_outputs(6459) <= '1';
    layer0_outputs(6460) <= not(inputs(29)) or (inputs(41));
    layer0_outputs(6461) <= (inputs(65)) xor (inputs(20));
    layer0_outputs(6462) <= not(inputs(57));
    layer0_outputs(6463) <= (inputs(219)) and not (inputs(72));
    layer0_outputs(6464) <= not((inputs(198)) xor (inputs(110)));
    layer0_outputs(6465) <= not(inputs(147)) or (inputs(17));
    layer0_outputs(6466) <= (inputs(40)) and not (inputs(208));
    layer0_outputs(6467) <= inputs(48);
    layer0_outputs(6468) <= inputs(43);
    layer0_outputs(6469) <= '1';
    layer0_outputs(6470) <= (inputs(217)) and not (inputs(0));
    layer0_outputs(6471) <= not((inputs(227)) xor (inputs(27)));
    layer0_outputs(6472) <= '0';
    layer0_outputs(6473) <= (inputs(145)) or (inputs(180));
    layer0_outputs(6474) <= inputs(110);
    layer0_outputs(6475) <= not((inputs(199)) xor (inputs(43)));
    layer0_outputs(6476) <= not((inputs(44)) or (inputs(242)));
    layer0_outputs(6477) <= inputs(97);
    layer0_outputs(6478) <= not(inputs(99));
    layer0_outputs(6479) <= not((inputs(198)) or (inputs(238)));
    layer0_outputs(6480) <= (inputs(149)) or (inputs(64));
    layer0_outputs(6481) <= (inputs(86)) or (inputs(202));
    layer0_outputs(6482) <= not((inputs(18)) or (inputs(191)));
    layer0_outputs(6483) <= (inputs(238)) xor (inputs(10));
    layer0_outputs(6484) <= (inputs(141)) or (inputs(59));
    layer0_outputs(6485) <= (inputs(225)) or (inputs(186));
    layer0_outputs(6486) <= (inputs(50)) or (inputs(43));
    layer0_outputs(6487) <= not(inputs(213));
    layer0_outputs(6488) <= '0';
    layer0_outputs(6489) <= inputs(180);
    layer0_outputs(6490) <= not(inputs(133));
    layer0_outputs(6491) <= (inputs(105)) xor (inputs(143));
    layer0_outputs(6492) <= (inputs(37)) and not (inputs(221));
    layer0_outputs(6493) <= inputs(133);
    layer0_outputs(6494) <= (inputs(196)) xor (inputs(227));
    layer0_outputs(6495) <= not((inputs(240)) xor (inputs(87)));
    layer0_outputs(6496) <= (inputs(135)) xor (inputs(237));
    layer0_outputs(6497) <= not((inputs(132)) xor (inputs(37)));
    layer0_outputs(6498) <= not(inputs(213));
    layer0_outputs(6499) <= (inputs(7)) or (inputs(94));
    layer0_outputs(6500) <= (inputs(12)) or (inputs(153));
    layer0_outputs(6501) <= not(inputs(234));
    layer0_outputs(6502) <= not(inputs(230)) or (inputs(122));
    layer0_outputs(6503) <= (inputs(73)) and not (inputs(236));
    layer0_outputs(6504) <= not((inputs(5)) xor (inputs(95)));
    layer0_outputs(6505) <= not(inputs(217)) or (inputs(21));
    layer0_outputs(6506) <= (inputs(194)) and (inputs(204));
    layer0_outputs(6507) <= not((inputs(91)) xor (inputs(94)));
    layer0_outputs(6508) <= not((inputs(46)) or (inputs(57)));
    layer0_outputs(6509) <= (inputs(92)) or (inputs(245));
    layer0_outputs(6510) <= (inputs(162)) and not (inputs(48));
    layer0_outputs(6511) <= not((inputs(188)) xor (inputs(13)));
    layer0_outputs(6512) <= (inputs(43)) and not (inputs(192));
    layer0_outputs(6513) <= not(inputs(227));
    layer0_outputs(6514) <= inputs(176);
    layer0_outputs(6515) <= not(inputs(168));
    layer0_outputs(6516) <= not(inputs(184)) or (inputs(223));
    layer0_outputs(6517) <= (inputs(161)) or (inputs(20));
    layer0_outputs(6518) <= (inputs(171)) and not (inputs(201));
    layer0_outputs(6519) <= not((inputs(113)) or (inputs(216)));
    layer0_outputs(6520) <= inputs(21);
    layer0_outputs(6521) <= not(inputs(141)) or (inputs(108));
    layer0_outputs(6522) <= inputs(47);
    layer0_outputs(6523) <= (inputs(186)) or (inputs(171));
    layer0_outputs(6524) <= inputs(24);
    layer0_outputs(6525) <= not(inputs(74));
    layer0_outputs(6526) <= not(inputs(76));
    layer0_outputs(6527) <= (inputs(137)) and not (inputs(127));
    layer0_outputs(6528) <= (inputs(128)) or (inputs(68));
    layer0_outputs(6529) <= not((inputs(87)) or (inputs(201)));
    layer0_outputs(6530) <= (inputs(66)) and not (inputs(73));
    layer0_outputs(6531) <= inputs(25);
    layer0_outputs(6532) <= not(inputs(30));
    layer0_outputs(6533) <= not((inputs(44)) or (inputs(77)));
    layer0_outputs(6534) <= not(inputs(120));
    layer0_outputs(6535) <= not((inputs(85)) xor (inputs(113)));
    layer0_outputs(6536) <= not((inputs(48)) xor (inputs(4)));
    layer0_outputs(6537) <= not(inputs(86));
    layer0_outputs(6538) <= inputs(101);
    layer0_outputs(6539) <= inputs(120);
    layer0_outputs(6540) <= not(inputs(104));
    layer0_outputs(6541) <= inputs(171);
    layer0_outputs(6542) <= (inputs(156)) or (inputs(98));
    layer0_outputs(6543) <= not((inputs(193)) and (inputs(206)));
    layer0_outputs(6544) <= (inputs(75)) or (inputs(224));
    layer0_outputs(6545) <= not((inputs(213)) and (inputs(20)));
    layer0_outputs(6546) <= (inputs(64)) or (inputs(144));
    layer0_outputs(6547) <= (inputs(41)) or (inputs(194));
    layer0_outputs(6548) <= not(inputs(137)) or (inputs(160));
    layer0_outputs(6549) <= not(inputs(231));
    layer0_outputs(6550) <= not((inputs(19)) or (inputs(244)));
    layer0_outputs(6551) <= not(inputs(128));
    layer0_outputs(6552) <= (inputs(65)) or (inputs(135));
    layer0_outputs(6553) <= not((inputs(77)) or (inputs(111)));
    layer0_outputs(6554) <= not(inputs(231));
    layer0_outputs(6555) <= (inputs(84)) and not (inputs(162));
    layer0_outputs(6556) <= (inputs(6)) and not (inputs(2));
    layer0_outputs(6557) <= not(inputs(84)) or (inputs(224));
    layer0_outputs(6558) <= (inputs(208)) and (inputs(130));
    layer0_outputs(6559) <= inputs(4);
    layer0_outputs(6560) <= (inputs(105)) and not (inputs(149));
    layer0_outputs(6561) <= not(inputs(232)) or (inputs(78));
    layer0_outputs(6562) <= (inputs(137)) xor (inputs(156));
    layer0_outputs(6563) <= not((inputs(35)) or (inputs(14)));
    layer0_outputs(6564) <= not((inputs(161)) or (inputs(101)));
    layer0_outputs(6565) <= inputs(53);
    layer0_outputs(6566) <= (inputs(21)) and not (inputs(83));
    layer0_outputs(6567) <= (inputs(108)) and not (inputs(237));
    layer0_outputs(6568) <= not((inputs(201)) or (inputs(176)));
    layer0_outputs(6569) <= inputs(146);
    layer0_outputs(6570) <= not(inputs(21)) or (inputs(185));
    layer0_outputs(6571) <= not(inputs(92));
    layer0_outputs(6572) <= not((inputs(53)) or (inputs(97)));
    layer0_outputs(6573) <= (inputs(48)) or (inputs(246));
    layer0_outputs(6574) <= inputs(206);
    layer0_outputs(6575) <= inputs(140);
    layer0_outputs(6576) <= inputs(166);
    layer0_outputs(6577) <= not(inputs(227));
    layer0_outputs(6578) <= (inputs(165)) xor (inputs(226));
    layer0_outputs(6579) <= (inputs(221)) or (inputs(190));
    layer0_outputs(6580) <= not(inputs(146));
    layer0_outputs(6581) <= (inputs(35)) or (inputs(89));
    layer0_outputs(6582) <= (inputs(154)) or (inputs(172));
    layer0_outputs(6583) <= (inputs(207)) or (inputs(202));
    layer0_outputs(6584) <= '1';
    layer0_outputs(6585) <= not((inputs(67)) or (inputs(38)));
    layer0_outputs(6586) <= not(inputs(1));
    layer0_outputs(6587) <= not((inputs(222)) or (inputs(2)));
    layer0_outputs(6588) <= not(inputs(117));
    layer0_outputs(6589) <= not(inputs(245));
    layer0_outputs(6590) <= (inputs(189)) or (inputs(201));
    layer0_outputs(6591) <= not(inputs(69)) or (inputs(225));
    layer0_outputs(6592) <= not((inputs(166)) xor (inputs(130)));
    layer0_outputs(6593) <= (inputs(237)) and not (inputs(48));
    layer0_outputs(6594) <= (inputs(60)) and not (inputs(195));
    layer0_outputs(6595) <= not(inputs(50));
    layer0_outputs(6596) <= (inputs(49)) or (inputs(180));
    layer0_outputs(6597) <= inputs(117);
    layer0_outputs(6598) <= not(inputs(84));
    layer0_outputs(6599) <= (inputs(179)) and not (inputs(222));
    layer0_outputs(6600) <= (inputs(22)) or (inputs(126));
    layer0_outputs(6601) <= inputs(86);
    layer0_outputs(6602) <= inputs(216);
    layer0_outputs(6603) <= (inputs(188)) and (inputs(103));
    layer0_outputs(6604) <= not(inputs(82));
    layer0_outputs(6605) <= (inputs(37)) and not (inputs(109));
    layer0_outputs(6606) <= inputs(209);
    layer0_outputs(6607) <= '1';
    layer0_outputs(6608) <= (inputs(104)) xor (inputs(57));
    layer0_outputs(6609) <= not((inputs(253)) or (inputs(99)));
    layer0_outputs(6610) <= inputs(116);
    layer0_outputs(6611) <= not((inputs(11)) or (inputs(110)));
    layer0_outputs(6612) <= not(inputs(200)) or (inputs(159));
    layer0_outputs(6613) <= not(inputs(138)) or (inputs(209));
    layer0_outputs(6614) <= (inputs(102)) or (inputs(178));
    layer0_outputs(6615) <= (inputs(205)) or (inputs(218));
    layer0_outputs(6616) <= not(inputs(232));
    layer0_outputs(6617) <= (inputs(98)) or (inputs(153));
    layer0_outputs(6618) <= inputs(253);
    layer0_outputs(6619) <= (inputs(135)) and not (inputs(17));
    layer0_outputs(6620) <= '0';
    layer0_outputs(6621) <= '0';
    layer0_outputs(6622) <= (inputs(212)) and not (inputs(79));
    layer0_outputs(6623) <= not(inputs(104));
    layer0_outputs(6624) <= not(inputs(79)) or (inputs(65));
    layer0_outputs(6625) <= not(inputs(14));
    layer0_outputs(6626) <= not(inputs(23)) or (inputs(145));
    layer0_outputs(6627) <= not((inputs(115)) or (inputs(135)));
    layer0_outputs(6628) <= inputs(13);
    layer0_outputs(6629) <= inputs(36);
    layer0_outputs(6630) <= '1';
    layer0_outputs(6631) <= (inputs(27)) or (inputs(171));
    layer0_outputs(6632) <= not((inputs(5)) or (inputs(225)));
    layer0_outputs(6633) <= not(inputs(126));
    layer0_outputs(6634) <= not((inputs(135)) xor (inputs(238)));
    layer0_outputs(6635) <= not(inputs(73)) or (inputs(146));
    layer0_outputs(6636) <= (inputs(124)) or (inputs(139));
    layer0_outputs(6637) <= not(inputs(88)) or (inputs(251));
    layer0_outputs(6638) <= not(inputs(247));
    layer0_outputs(6639) <= not((inputs(88)) or (inputs(121)));
    layer0_outputs(6640) <= (inputs(195)) xor (inputs(124));
    layer0_outputs(6641) <= inputs(61);
    layer0_outputs(6642) <= not(inputs(72));
    layer0_outputs(6643) <= inputs(184);
    layer0_outputs(6644) <= (inputs(3)) xor (inputs(31));
    layer0_outputs(6645) <= not(inputs(221)) or (inputs(50));
    layer0_outputs(6646) <= inputs(6);
    layer0_outputs(6647) <= inputs(33);
    layer0_outputs(6648) <= (inputs(99)) and not (inputs(95));
    layer0_outputs(6649) <= (inputs(86)) xor (inputs(52));
    layer0_outputs(6650) <= inputs(117);
    layer0_outputs(6651) <= not(inputs(102)) or (inputs(108));
    layer0_outputs(6652) <= inputs(165);
    layer0_outputs(6653) <= not((inputs(221)) or (inputs(170)));
    layer0_outputs(6654) <= inputs(19);
    layer0_outputs(6655) <= not((inputs(74)) or (inputs(63)));
    layer0_outputs(6656) <= inputs(17);
    layer0_outputs(6657) <= inputs(227);
    layer0_outputs(6658) <= inputs(59);
    layer0_outputs(6659) <= (inputs(158)) and (inputs(200));
    layer0_outputs(6660) <= (inputs(103)) xor (inputs(138));
    layer0_outputs(6661) <= (inputs(246)) and not (inputs(31));
    layer0_outputs(6662) <= (inputs(38)) xor (inputs(71));
    layer0_outputs(6663) <= (inputs(64)) and not (inputs(56));
    layer0_outputs(6664) <= not((inputs(202)) or (inputs(51)));
    layer0_outputs(6665) <= not(inputs(226));
    layer0_outputs(6666) <= (inputs(229)) and not (inputs(89));
    layer0_outputs(6667) <= (inputs(26)) and not (inputs(142));
    layer0_outputs(6668) <= '1';
    layer0_outputs(6669) <= (inputs(73)) or (inputs(28));
    layer0_outputs(6670) <= not(inputs(37));
    layer0_outputs(6671) <= (inputs(8)) or (inputs(173));
    layer0_outputs(6672) <= not((inputs(211)) or (inputs(53)));
    layer0_outputs(6673) <= inputs(179);
    layer0_outputs(6674) <= (inputs(63)) or (inputs(216));
    layer0_outputs(6675) <= inputs(181);
    layer0_outputs(6676) <= not((inputs(173)) or (inputs(64)));
    layer0_outputs(6677) <= inputs(195);
    layer0_outputs(6678) <= not((inputs(22)) or (inputs(122)));
    layer0_outputs(6679) <= (inputs(195)) and not (inputs(55));
    layer0_outputs(6680) <= inputs(83);
    layer0_outputs(6681) <= not(inputs(68)) or (inputs(111));
    layer0_outputs(6682) <= not(inputs(50)) or (inputs(218));
    layer0_outputs(6683) <= (inputs(186)) and not (inputs(136));
    layer0_outputs(6684) <= not(inputs(76));
    layer0_outputs(6685) <= (inputs(106)) and not (inputs(254));
    layer0_outputs(6686) <= (inputs(23)) and not (inputs(233));
    layer0_outputs(6687) <= not((inputs(6)) or (inputs(47)));
    layer0_outputs(6688) <= not(inputs(99));
    layer0_outputs(6689) <= (inputs(166)) xor (inputs(114));
    layer0_outputs(6690) <= inputs(82);
    layer0_outputs(6691) <= (inputs(157)) or (inputs(148));
    layer0_outputs(6692) <= not(inputs(204));
    layer0_outputs(6693) <= (inputs(50)) and (inputs(69));
    layer0_outputs(6694) <= not(inputs(215)) or (inputs(62));
    layer0_outputs(6695) <= not(inputs(197)) or (inputs(0));
    layer0_outputs(6696) <= inputs(212);
    layer0_outputs(6697) <= not((inputs(229)) or (inputs(97)));
    layer0_outputs(6698) <= (inputs(49)) xor (inputs(24));
    layer0_outputs(6699) <= (inputs(31)) or (inputs(106));
    layer0_outputs(6700) <= not((inputs(187)) or (inputs(221)));
    layer0_outputs(6701) <= (inputs(126)) and (inputs(87));
    layer0_outputs(6702) <= inputs(194);
    layer0_outputs(6703) <= (inputs(72)) and (inputs(155));
    layer0_outputs(6704) <= not((inputs(11)) and (inputs(214)));
    layer0_outputs(6705) <= not(inputs(165)) or (inputs(113));
    layer0_outputs(6706) <= not((inputs(71)) xor (inputs(244)));
    layer0_outputs(6707) <= not((inputs(86)) xor (inputs(38)));
    layer0_outputs(6708) <= not((inputs(139)) xor (inputs(218)));
    layer0_outputs(6709) <= not(inputs(230));
    layer0_outputs(6710) <= (inputs(122)) and not (inputs(194));
    layer0_outputs(6711) <= not(inputs(98));
    layer0_outputs(6712) <= not((inputs(196)) xor (inputs(173)));
    layer0_outputs(6713) <= (inputs(47)) and not (inputs(200));
    layer0_outputs(6714) <= inputs(169);
    layer0_outputs(6715) <= (inputs(158)) xor (inputs(221));
    layer0_outputs(6716) <= not((inputs(198)) xor (inputs(244)));
    layer0_outputs(6717) <= not(inputs(163));
    layer0_outputs(6718) <= not(inputs(22));
    layer0_outputs(6719) <= inputs(212);
    layer0_outputs(6720) <= not(inputs(32));
    layer0_outputs(6721) <= not(inputs(125)) or (inputs(42));
    layer0_outputs(6722) <= inputs(220);
    layer0_outputs(6723) <= not(inputs(165));
    layer0_outputs(6724) <= inputs(245);
    layer0_outputs(6725) <= not(inputs(7));
    layer0_outputs(6726) <= not((inputs(14)) or (inputs(31)));
    layer0_outputs(6727) <= (inputs(14)) and not (inputs(38));
    layer0_outputs(6728) <= not((inputs(33)) xor (inputs(157)));
    layer0_outputs(6729) <= not(inputs(93));
    layer0_outputs(6730) <= (inputs(116)) and not (inputs(30));
    layer0_outputs(6731) <= not((inputs(177)) xor (inputs(201)));
    layer0_outputs(6732) <= (inputs(81)) or (inputs(54));
    layer0_outputs(6733) <= (inputs(9)) and not (inputs(118));
    layer0_outputs(6734) <= not(inputs(91));
    layer0_outputs(6735) <= not(inputs(7)) or (inputs(250));
    layer0_outputs(6736) <= inputs(77);
    layer0_outputs(6737) <= not(inputs(30)) or (inputs(240));
    layer0_outputs(6738) <= inputs(162);
    layer0_outputs(6739) <= inputs(253);
    layer0_outputs(6740) <= not((inputs(86)) xor (inputs(112)));
    layer0_outputs(6741) <= not(inputs(124)) or (inputs(56));
    layer0_outputs(6742) <= not(inputs(58)) or (inputs(217));
    layer0_outputs(6743) <= (inputs(20)) and (inputs(54));
    layer0_outputs(6744) <= not((inputs(9)) or (inputs(171)));
    layer0_outputs(6745) <= inputs(196);
    layer0_outputs(6746) <= inputs(227);
    layer0_outputs(6747) <= (inputs(211)) and not (inputs(113));
    layer0_outputs(6748) <= (inputs(50)) and not (inputs(73));
    layer0_outputs(6749) <= (inputs(188)) and not (inputs(128));
    layer0_outputs(6750) <= (inputs(84)) and not (inputs(206));
    layer0_outputs(6751) <= not(inputs(107)) or (inputs(210));
    layer0_outputs(6752) <= '0';
    layer0_outputs(6753) <= not(inputs(25));
    layer0_outputs(6754) <= not(inputs(82)) or (inputs(220));
    layer0_outputs(6755) <= not((inputs(237)) or (inputs(51)));
    layer0_outputs(6756) <= (inputs(209)) or (inputs(197));
    layer0_outputs(6757) <= inputs(135);
    layer0_outputs(6758) <= (inputs(174)) or (inputs(178));
    layer0_outputs(6759) <= inputs(252);
    layer0_outputs(6760) <= (inputs(193)) xor (inputs(247));
    layer0_outputs(6761) <= not(inputs(73));
    layer0_outputs(6762) <= not(inputs(212)) or (inputs(254));
    layer0_outputs(6763) <= (inputs(133)) or (inputs(242));
    layer0_outputs(6764) <= (inputs(178)) or (inputs(254));
    layer0_outputs(6765) <= (inputs(250)) or (inputs(187));
    layer0_outputs(6766) <= inputs(216);
    layer0_outputs(6767) <= (inputs(200)) and not (inputs(7));
    layer0_outputs(6768) <= not((inputs(89)) xor (inputs(252)));
    layer0_outputs(6769) <= (inputs(2)) and not (inputs(175));
    layer0_outputs(6770) <= not(inputs(231));
    layer0_outputs(6771) <= (inputs(151)) and not (inputs(205));
    layer0_outputs(6772) <= inputs(185);
    layer0_outputs(6773) <= inputs(51);
    layer0_outputs(6774) <= not(inputs(118));
    layer0_outputs(6775) <= (inputs(246)) xor (inputs(125));
    layer0_outputs(6776) <= not(inputs(53));
    layer0_outputs(6777) <= not(inputs(144)) or (inputs(247));
    layer0_outputs(6778) <= not(inputs(9)) or (inputs(194));
    layer0_outputs(6779) <= not((inputs(47)) or (inputs(161)));
    layer0_outputs(6780) <= not((inputs(164)) or (inputs(182)));
    layer0_outputs(6781) <= inputs(100);
    layer0_outputs(6782) <= not((inputs(0)) or (inputs(186)));
    layer0_outputs(6783) <= not(inputs(207)) or (inputs(126));
    layer0_outputs(6784) <= not((inputs(38)) or (inputs(144)));
    layer0_outputs(6785) <= (inputs(174)) xor (inputs(240));
    layer0_outputs(6786) <= inputs(147);
    layer0_outputs(6787) <= not(inputs(71));
    layer0_outputs(6788) <= not(inputs(215));
    layer0_outputs(6789) <= not((inputs(177)) or (inputs(231)));
    layer0_outputs(6790) <= inputs(171);
    layer0_outputs(6791) <= (inputs(93)) or (inputs(56));
    layer0_outputs(6792) <= (inputs(157)) or (inputs(61));
    layer0_outputs(6793) <= not(inputs(85));
    layer0_outputs(6794) <= (inputs(151)) xor (inputs(162));
    layer0_outputs(6795) <= not(inputs(99));
    layer0_outputs(6796) <= inputs(3);
    layer0_outputs(6797) <= '0';
    layer0_outputs(6798) <= not(inputs(17));
    layer0_outputs(6799) <= (inputs(158)) or (inputs(247));
    layer0_outputs(6800) <= not(inputs(99));
    layer0_outputs(6801) <= (inputs(250)) and not (inputs(31));
    layer0_outputs(6802) <= (inputs(60)) or (inputs(146));
    layer0_outputs(6803) <= inputs(84);
    layer0_outputs(6804) <= not((inputs(151)) or (inputs(196)));
    layer0_outputs(6805) <= not(inputs(247));
    layer0_outputs(6806) <= not((inputs(159)) or (inputs(187)));
    layer0_outputs(6807) <= not(inputs(105)) or (inputs(144));
    layer0_outputs(6808) <= inputs(143);
    layer0_outputs(6809) <= not((inputs(221)) and (inputs(12)));
    layer0_outputs(6810) <= not(inputs(76)) or (inputs(241));
    layer0_outputs(6811) <= (inputs(176)) or (inputs(202));
    layer0_outputs(6812) <= not((inputs(1)) or (inputs(164)));
    layer0_outputs(6813) <= not(inputs(93)) or (inputs(232));
    layer0_outputs(6814) <= not(inputs(209)) or (inputs(48));
    layer0_outputs(6815) <= not((inputs(47)) or (inputs(122)));
    layer0_outputs(6816) <= (inputs(52)) and not (inputs(23));
    layer0_outputs(6817) <= (inputs(176)) or (inputs(215));
    layer0_outputs(6818) <= (inputs(252)) and not (inputs(175));
    layer0_outputs(6819) <= inputs(83);
    layer0_outputs(6820) <= inputs(25);
    layer0_outputs(6821) <= not(inputs(114));
    layer0_outputs(6822) <= (inputs(242)) and not (inputs(115));
    layer0_outputs(6823) <= (inputs(134)) xor (inputs(81));
    layer0_outputs(6824) <= (inputs(238)) or (inputs(142));
    layer0_outputs(6825) <= inputs(123);
    layer0_outputs(6826) <= inputs(208);
    layer0_outputs(6827) <= (inputs(107)) and not (inputs(57));
    layer0_outputs(6828) <= not((inputs(113)) or (inputs(113)));
    layer0_outputs(6829) <= not(inputs(246));
    layer0_outputs(6830) <= inputs(206);
    layer0_outputs(6831) <= not(inputs(23)) or (inputs(84));
    layer0_outputs(6832) <= not(inputs(175));
    layer0_outputs(6833) <= inputs(167);
    layer0_outputs(6834) <= not((inputs(69)) xor (inputs(2)));
    layer0_outputs(6835) <= not((inputs(121)) and (inputs(68)));
    layer0_outputs(6836) <= (inputs(27)) and (inputs(93));
    layer0_outputs(6837) <= (inputs(94)) or (inputs(183));
    layer0_outputs(6838) <= not((inputs(119)) or (inputs(54)));
    layer0_outputs(6839) <= not(inputs(178));
    layer0_outputs(6840) <= not(inputs(136));
    layer0_outputs(6841) <= (inputs(104)) and not (inputs(164));
    layer0_outputs(6842) <= (inputs(120)) and not (inputs(161));
    layer0_outputs(6843) <= not((inputs(49)) or (inputs(156)));
    layer0_outputs(6844) <= inputs(102);
    layer0_outputs(6845) <= not((inputs(237)) or (inputs(235)));
    layer0_outputs(6846) <= not(inputs(121));
    layer0_outputs(6847) <= not(inputs(112));
    layer0_outputs(6848) <= inputs(99);
    layer0_outputs(6849) <= not(inputs(12));
    layer0_outputs(6850) <= not(inputs(167));
    layer0_outputs(6851) <= (inputs(123)) and not (inputs(115));
    layer0_outputs(6852) <= not(inputs(229));
    layer0_outputs(6853) <= (inputs(232)) and not (inputs(163));
    layer0_outputs(6854) <= (inputs(70)) xor (inputs(99));
    layer0_outputs(6855) <= not(inputs(54));
    layer0_outputs(6856) <= not(inputs(201)) or (inputs(65));
    layer0_outputs(6857) <= (inputs(34)) xor (inputs(5));
    layer0_outputs(6858) <= not(inputs(42));
    layer0_outputs(6859) <= not((inputs(167)) or (inputs(146)));
    layer0_outputs(6860) <= (inputs(46)) or (inputs(21));
    layer0_outputs(6861) <= (inputs(245)) or (inputs(103));
    layer0_outputs(6862) <= not(inputs(217));
    layer0_outputs(6863) <= not(inputs(159));
    layer0_outputs(6864) <= not((inputs(235)) or (inputs(191)));
    layer0_outputs(6865) <= inputs(212);
    layer0_outputs(6866) <= '0';
    layer0_outputs(6867) <= not((inputs(143)) or (inputs(218)));
    layer0_outputs(6868) <= not(inputs(254));
    layer0_outputs(6869) <= inputs(115);
    layer0_outputs(6870) <= not(inputs(215));
    layer0_outputs(6871) <= not(inputs(190)) or (inputs(106));
    layer0_outputs(6872) <= (inputs(23)) xor (inputs(55));
    layer0_outputs(6873) <= not(inputs(75));
    layer0_outputs(6874) <= (inputs(135)) and not (inputs(129));
    layer0_outputs(6875) <= (inputs(213)) or (inputs(20));
    layer0_outputs(6876) <= (inputs(215)) and (inputs(217));
    layer0_outputs(6877) <= not((inputs(235)) and (inputs(210)));
    layer0_outputs(6878) <= not((inputs(214)) and (inputs(236)));
    layer0_outputs(6879) <= inputs(180);
    layer0_outputs(6880) <= not(inputs(96)) or (inputs(191));
    layer0_outputs(6881) <= not(inputs(45));
    layer0_outputs(6882) <= not(inputs(36)) or (inputs(143));
    layer0_outputs(6883) <= not((inputs(193)) and (inputs(107)));
    layer0_outputs(6884) <= (inputs(68)) xor (inputs(70));
    layer0_outputs(6885) <= not((inputs(40)) xor (inputs(28)));
    layer0_outputs(6886) <= not(inputs(85)) or (inputs(158));
    layer0_outputs(6887) <= (inputs(213)) and not (inputs(56));
    layer0_outputs(6888) <= not((inputs(60)) or (inputs(123)));
    layer0_outputs(6889) <= (inputs(24)) and not (inputs(163));
    layer0_outputs(6890) <= (inputs(178)) or (inputs(188));
    layer0_outputs(6891) <= (inputs(234)) xor (inputs(183));
    layer0_outputs(6892) <= not(inputs(22)) or (inputs(162));
    layer0_outputs(6893) <= not(inputs(197)) or (inputs(160));
    layer0_outputs(6894) <= (inputs(11)) xor (inputs(183));
    layer0_outputs(6895) <= not((inputs(199)) or (inputs(243)));
    layer0_outputs(6896) <= inputs(151);
    layer0_outputs(6897) <= not(inputs(53));
    layer0_outputs(6898) <= inputs(239);
    layer0_outputs(6899) <= (inputs(93)) and not (inputs(188));
    layer0_outputs(6900) <= (inputs(77)) and not (inputs(255));
    layer0_outputs(6901) <= not((inputs(104)) xor (inputs(95)));
    layer0_outputs(6902) <= not((inputs(106)) or (inputs(163)));
    layer0_outputs(6903) <= not(inputs(164));
    layer0_outputs(6904) <= inputs(215);
    layer0_outputs(6905) <= not(inputs(50)) or (inputs(30));
    layer0_outputs(6906) <= not(inputs(113));
    layer0_outputs(6907) <= not(inputs(165));
    layer0_outputs(6908) <= not((inputs(130)) or (inputs(45)));
    layer0_outputs(6909) <= not(inputs(51));
    layer0_outputs(6910) <= not(inputs(94)) or (inputs(137));
    layer0_outputs(6911) <= not((inputs(1)) or (inputs(180)));
    layer0_outputs(6912) <= inputs(104);
    layer0_outputs(6913) <= not(inputs(246));
    layer0_outputs(6914) <= (inputs(3)) xor (inputs(198));
    layer0_outputs(6915) <= not(inputs(53));
    layer0_outputs(6916) <= not((inputs(9)) or (inputs(25)));
    layer0_outputs(6917) <= (inputs(9)) xor (inputs(7));
    layer0_outputs(6918) <= not((inputs(52)) or (inputs(109)));
    layer0_outputs(6919) <= (inputs(222)) xor (inputs(141));
    layer0_outputs(6920) <= not((inputs(172)) or (inputs(124)));
    layer0_outputs(6921) <= not(inputs(245));
    layer0_outputs(6922) <= not(inputs(140)) or (inputs(110));
    layer0_outputs(6923) <= inputs(229);
    layer0_outputs(6924) <= (inputs(251)) or (inputs(81));
    layer0_outputs(6925) <= inputs(83);
    layer0_outputs(6926) <= not(inputs(66));
    layer0_outputs(6927) <= (inputs(134)) and (inputs(56));
    layer0_outputs(6928) <= (inputs(95)) xor (inputs(233));
    layer0_outputs(6929) <= (inputs(226)) xor (inputs(200));
    layer0_outputs(6930) <= not((inputs(202)) xor (inputs(138)));
    layer0_outputs(6931) <= (inputs(244)) xor (inputs(22));
    layer0_outputs(6932) <= (inputs(157)) and not (inputs(169));
    layer0_outputs(6933) <= not(inputs(101)) or (inputs(33));
    layer0_outputs(6934) <= (inputs(107)) xor (inputs(110));
    layer0_outputs(6935) <= not(inputs(83));
    layer0_outputs(6936) <= not(inputs(167));
    layer0_outputs(6937) <= (inputs(133)) or (inputs(187));
    layer0_outputs(6938) <= not((inputs(208)) or (inputs(171)));
    layer0_outputs(6939) <= not(inputs(111));
    layer0_outputs(6940) <= inputs(9);
    layer0_outputs(6941) <= not(inputs(199)) or (inputs(64));
    layer0_outputs(6942) <= (inputs(69)) and not (inputs(0));
    layer0_outputs(6943) <= (inputs(173)) or (inputs(219));
    layer0_outputs(6944) <= inputs(163);
    layer0_outputs(6945) <= (inputs(36)) or (inputs(205));
    layer0_outputs(6946) <= (inputs(157)) xor (inputs(123));
    layer0_outputs(6947) <= (inputs(123)) or (inputs(233));
    layer0_outputs(6948) <= not(inputs(114));
    layer0_outputs(6949) <= not((inputs(20)) xor (inputs(204)));
    layer0_outputs(6950) <= not(inputs(67)) or (inputs(143));
    layer0_outputs(6951) <= not((inputs(226)) or (inputs(159)));
    layer0_outputs(6952) <= not((inputs(27)) xor (inputs(230)));
    layer0_outputs(6953) <= not(inputs(179));
    layer0_outputs(6954) <= (inputs(213)) xor (inputs(246));
    layer0_outputs(6955) <= inputs(179);
    layer0_outputs(6956) <= not(inputs(214)) or (inputs(85));
    layer0_outputs(6957) <= not((inputs(182)) xor (inputs(131)));
    layer0_outputs(6958) <= not(inputs(231)) or (inputs(40));
    layer0_outputs(6959) <= (inputs(144)) or (inputs(186));
    layer0_outputs(6960) <= '1';
    layer0_outputs(6961) <= inputs(205);
    layer0_outputs(6962) <= not(inputs(146));
    layer0_outputs(6963) <= not(inputs(72)) or (inputs(170));
    layer0_outputs(6964) <= not(inputs(155));
    layer0_outputs(6965) <= not((inputs(226)) or (inputs(148)));
    layer0_outputs(6966) <= inputs(160);
    layer0_outputs(6967) <= not((inputs(96)) or (inputs(75)));
    layer0_outputs(6968) <= not((inputs(69)) xor (inputs(77)));
    layer0_outputs(6969) <= inputs(80);
    layer0_outputs(6970) <= '0';
    layer0_outputs(6971) <= inputs(0);
    layer0_outputs(6972) <= (inputs(213)) and not (inputs(56));
    layer0_outputs(6973) <= (inputs(122)) and (inputs(107));
    layer0_outputs(6974) <= (inputs(201)) or (inputs(160));
    layer0_outputs(6975) <= inputs(46);
    layer0_outputs(6976) <= (inputs(250)) xor (inputs(154));
    layer0_outputs(6977) <= (inputs(238)) or (inputs(203));
    layer0_outputs(6978) <= not(inputs(22)) or (inputs(163));
    layer0_outputs(6979) <= not((inputs(228)) and (inputs(187)));
    layer0_outputs(6980) <= not(inputs(239));
    layer0_outputs(6981) <= inputs(114);
    layer0_outputs(6982) <= not((inputs(126)) or (inputs(194)));
    layer0_outputs(6983) <= inputs(25);
    layer0_outputs(6984) <= not(inputs(135));
    layer0_outputs(6985) <= not(inputs(182)) or (inputs(157));
    layer0_outputs(6986) <= not((inputs(220)) xor (inputs(6)));
    layer0_outputs(6987) <= not(inputs(39));
    layer0_outputs(6988) <= not(inputs(106));
    layer0_outputs(6989) <= not((inputs(6)) or (inputs(21)));
    layer0_outputs(6990) <= (inputs(252)) xor (inputs(181));
    layer0_outputs(6991) <= not((inputs(11)) or (inputs(185)));
    layer0_outputs(6992) <= (inputs(26)) and (inputs(53));
    layer0_outputs(6993) <= not((inputs(80)) xor (inputs(196)));
    layer0_outputs(6994) <= (inputs(239)) and not (inputs(83));
    layer0_outputs(6995) <= not(inputs(193));
    layer0_outputs(6996) <= inputs(162);
    layer0_outputs(6997) <= '1';
    layer0_outputs(6998) <= not(inputs(68)) or (inputs(175));
    layer0_outputs(6999) <= not(inputs(154)) or (inputs(241));
    layer0_outputs(7000) <= (inputs(247)) and not (inputs(81));
    layer0_outputs(7001) <= not(inputs(9));
    layer0_outputs(7002) <= (inputs(146)) or (inputs(169));
    layer0_outputs(7003) <= (inputs(254)) and not (inputs(241));
    layer0_outputs(7004) <= (inputs(153)) and (inputs(139));
    layer0_outputs(7005) <= inputs(68);
    layer0_outputs(7006) <= inputs(81);
    layer0_outputs(7007) <= not((inputs(152)) and (inputs(220)));
    layer0_outputs(7008) <= inputs(229);
    layer0_outputs(7009) <= not(inputs(169)) or (inputs(229));
    layer0_outputs(7010) <= not(inputs(19));
    layer0_outputs(7011) <= inputs(159);
    layer0_outputs(7012) <= (inputs(138)) or (inputs(253));
    layer0_outputs(7013) <= not(inputs(136)) or (inputs(113));
    layer0_outputs(7014) <= not((inputs(192)) or (inputs(186)));
    layer0_outputs(7015) <= (inputs(213)) or (inputs(229));
    layer0_outputs(7016) <= (inputs(93)) xor (inputs(255));
    layer0_outputs(7017) <= (inputs(183)) or (inputs(14));
    layer0_outputs(7018) <= inputs(98);
    layer0_outputs(7019) <= not(inputs(192));
    layer0_outputs(7020) <= inputs(84);
    layer0_outputs(7021) <= not((inputs(254)) or (inputs(194)));
    layer0_outputs(7022) <= not(inputs(3)) or (inputs(128));
    layer0_outputs(7023) <= not((inputs(200)) xor (inputs(246)));
    layer0_outputs(7024) <= (inputs(115)) and not (inputs(34));
    layer0_outputs(7025) <= not(inputs(249)) or (inputs(60));
    layer0_outputs(7026) <= not(inputs(179)) or (inputs(253));
    layer0_outputs(7027) <= (inputs(103)) or (inputs(118));
    layer0_outputs(7028) <= (inputs(129)) or (inputs(140));
    layer0_outputs(7029) <= inputs(148);
    layer0_outputs(7030) <= inputs(186);
    layer0_outputs(7031) <= inputs(108);
    layer0_outputs(7032) <= not((inputs(44)) or (inputs(58)));
    layer0_outputs(7033) <= inputs(53);
    layer0_outputs(7034) <= (inputs(28)) xor (inputs(156));
    layer0_outputs(7035) <= (inputs(120)) or (inputs(173));
    layer0_outputs(7036) <= not(inputs(90));
    layer0_outputs(7037) <= not(inputs(115)) or (inputs(94));
    layer0_outputs(7038) <= (inputs(190)) xor (inputs(85));
    layer0_outputs(7039) <= not((inputs(222)) or (inputs(231)));
    layer0_outputs(7040) <= not(inputs(208)) or (inputs(41));
    layer0_outputs(7041) <= not((inputs(107)) and (inputs(152)));
    layer0_outputs(7042) <= not((inputs(158)) xor (inputs(176)));
    layer0_outputs(7043) <= not((inputs(171)) and (inputs(73)));
    layer0_outputs(7044) <= not(inputs(183)) or (inputs(88));
    layer0_outputs(7045) <= not(inputs(210)) or (inputs(60));
    layer0_outputs(7046) <= not((inputs(108)) xor (inputs(106)));
    layer0_outputs(7047) <= inputs(12);
    layer0_outputs(7048) <= (inputs(154)) or (inputs(17));
    layer0_outputs(7049) <= (inputs(91)) or (inputs(175));
    layer0_outputs(7050) <= not((inputs(13)) and (inputs(150)));
    layer0_outputs(7051) <= not((inputs(42)) or (inputs(86)));
    layer0_outputs(7052) <= inputs(221);
    layer0_outputs(7053) <= inputs(97);
    layer0_outputs(7054) <= not(inputs(147));
    layer0_outputs(7055) <= inputs(70);
    layer0_outputs(7056) <= (inputs(149)) or (inputs(147));
    layer0_outputs(7057) <= not((inputs(188)) or (inputs(47)));
    layer0_outputs(7058) <= (inputs(82)) and not (inputs(160));
    layer0_outputs(7059) <= (inputs(195)) and not (inputs(13));
    layer0_outputs(7060) <= inputs(118);
    layer0_outputs(7061) <= not(inputs(105));
    layer0_outputs(7062) <= not(inputs(146));
    layer0_outputs(7063) <= inputs(194);
    layer0_outputs(7064) <= not((inputs(148)) xor (inputs(98)));
    layer0_outputs(7065) <= not((inputs(194)) or (inputs(193)));
    layer0_outputs(7066) <= not(inputs(150));
    layer0_outputs(7067) <= (inputs(213)) or (inputs(198));
    layer0_outputs(7068) <= (inputs(30)) and not (inputs(146));
    layer0_outputs(7069) <= not(inputs(125));
    layer0_outputs(7070) <= (inputs(90)) or (inputs(89));
    layer0_outputs(7071) <= inputs(207);
    layer0_outputs(7072) <= not((inputs(149)) xor (inputs(237)));
    layer0_outputs(7073) <= not(inputs(73));
    layer0_outputs(7074) <= not(inputs(19));
    layer0_outputs(7075) <= not((inputs(42)) and (inputs(231)));
    layer0_outputs(7076) <= not(inputs(58)) or (inputs(40));
    layer0_outputs(7077) <= (inputs(203)) xor (inputs(34));
    layer0_outputs(7078) <= (inputs(202)) and not (inputs(95));
    layer0_outputs(7079) <= not((inputs(215)) and (inputs(216)));
    layer0_outputs(7080) <= not(inputs(232));
    layer0_outputs(7081) <= not(inputs(252)) or (inputs(16));
    layer0_outputs(7082) <= (inputs(39)) xor (inputs(173));
    layer0_outputs(7083) <= not(inputs(153));
    layer0_outputs(7084) <= not((inputs(250)) xor (inputs(221)));
    layer0_outputs(7085) <= not(inputs(28));
    layer0_outputs(7086) <= inputs(105);
    layer0_outputs(7087) <= not(inputs(55)) or (inputs(252));
    layer0_outputs(7088) <= not(inputs(5));
    layer0_outputs(7089) <= not((inputs(249)) or (inputs(16)));
    layer0_outputs(7090) <= inputs(17);
    layer0_outputs(7091) <= (inputs(105)) or (inputs(224));
    layer0_outputs(7092) <= not((inputs(1)) or (inputs(177)));
    layer0_outputs(7093) <= inputs(213);
    layer0_outputs(7094) <= inputs(148);
    layer0_outputs(7095) <= (inputs(32)) and not (inputs(24));
    layer0_outputs(7096) <= not((inputs(54)) or (inputs(3)));
    layer0_outputs(7097) <= not(inputs(63)) or (inputs(17));
    layer0_outputs(7098) <= (inputs(8)) and not (inputs(255));
    layer0_outputs(7099) <= (inputs(223)) or (inputs(111));
    layer0_outputs(7100) <= (inputs(14)) xor (inputs(73));
    layer0_outputs(7101) <= inputs(230);
    layer0_outputs(7102) <= (inputs(113)) and not (inputs(15));
    layer0_outputs(7103) <= inputs(68);
    layer0_outputs(7104) <= not((inputs(141)) and (inputs(62)));
    layer0_outputs(7105) <= not(inputs(241)) or (inputs(53));
    layer0_outputs(7106) <= inputs(85);
    layer0_outputs(7107) <= not(inputs(118)) or (inputs(61));
    layer0_outputs(7108) <= '0';
    layer0_outputs(7109) <= not((inputs(16)) or (inputs(209)));
    layer0_outputs(7110) <= inputs(197);
    layer0_outputs(7111) <= not(inputs(76));
    layer0_outputs(7112) <= not((inputs(42)) or (inputs(79)));
    layer0_outputs(7113) <= (inputs(191)) or (inputs(107));
    layer0_outputs(7114) <= inputs(201);
    layer0_outputs(7115) <= (inputs(130)) or (inputs(218));
    layer0_outputs(7116) <= not((inputs(20)) xor (inputs(78)));
    layer0_outputs(7117) <= inputs(21);
    layer0_outputs(7118) <= '0';
    layer0_outputs(7119) <= inputs(25);
    layer0_outputs(7120) <= not(inputs(230)) or (inputs(151));
    layer0_outputs(7121) <= not(inputs(8));
    layer0_outputs(7122) <= not(inputs(192)) or (inputs(143));
    layer0_outputs(7123) <= not((inputs(21)) xor (inputs(174)));
    layer0_outputs(7124) <= not(inputs(164)) or (inputs(143));
    layer0_outputs(7125) <= (inputs(166)) or (inputs(18));
    layer0_outputs(7126) <= not(inputs(68));
    layer0_outputs(7127) <= not((inputs(170)) xor (inputs(187)));
    layer0_outputs(7128) <= (inputs(141)) or (inputs(41));
    layer0_outputs(7129) <= (inputs(91)) and not (inputs(14));
    layer0_outputs(7130) <= not((inputs(245)) or (inputs(253)));
    layer0_outputs(7131) <= not((inputs(184)) or (inputs(113)));
    layer0_outputs(7132) <= (inputs(3)) and not (inputs(127));
    layer0_outputs(7133) <= not((inputs(242)) or (inputs(144)));
    layer0_outputs(7134) <= inputs(140);
    layer0_outputs(7135) <= not((inputs(254)) and (inputs(183)));
    layer0_outputs(7136) <= not(inputs(123)) or (inputs(132));
    layer0_outputs(7137) <= inputs(48);
    layer0_outputs(7138) <= not(inputs(2));
    layer0_outputs(7139) <= not((inputs(136)) xor (inputs(233)));
    layer0_outputs(7140) <= not(inputs(101));
    layer0_outputs(7141) <= (inputs(63)) or (inputs(28));
    layer0_outputs(7142) <= not((inputs(203)) or (inputs(145)));
    layer0_outputs(7143) <= not((inputs(157)) or (inputs(115)));
    layer0_outputs(7144) <= not((inputs(186)) and (inputs(183)));
    layer0_outputs(7145) <= not((inputs(168)) or (inputs(159)));
    layer0_outputs(7146) <= not(inputs(153));
    layer0_outputs(7147) <= inputs(100);
    layer0_outputs(7148) <= inputs(160);
    layer0_outputs(7149) <= not(inputs(99));
    layer0_outputs(7150) <= not(inputs(144)) or (inputs(113));
    layer0_outputs(7151) <= (inputs(169)) and not (inputs(228));
    layer0_outputs(7152) <= inputs(39);
    layer0_outputs(7153) <= not(inputs(139)) or (inputs(21));
    layer0_outputs(7154) <= not(inputs(180));
    layer0_outputs(7155) <= (inputs(229)) or (inputs(132));
    layer0_outputs(7156) <= not((inputs(22)) xor (inputs(195)));
    layer0_outputs(7157) <= (inputs(57)) and not (inputs(83));
    layer0_outputs(7158) <= (inputs(253)) or (inputs(31));
    layer0_outputs(7159) <= not(inputs(154));
    layer0_outputs(7160) <= not(inputs(109)) or (inputs(31));
    layer0_outputs(7161) <= (inputs(26)) and not (inputs(165));
    layer0_outputs(7162) <= not((inputs(179)) xor (inputs(91)));
    layer0_outputs(7163) <= (inputs(69)) or (inputs(231));
    layer0_outputs(7164) <= not(inputs(163)) or (inputs(78));
    layer0_outputs(7165) <= (inputs(187)) and not (inputs(137));
    layer0_outputs(7166) <= (inputs(27)) and not (inputs(35));
    layer0_outputs(7167) <= (inputs(146)) or (inputs(169));
    layer0_outputs(7168) <= not(inputs(120)) or (inputs(198));
    layer0_outputs(7169) <= not(inputs(240)) or (inputs(12));
    layer0_outputs(7170) <= not(inputs(151));
    layer0_outputs(7171) <= (inputs(117)) and not (inputs(90));
    layer0_outputs(7172) <= not((inputs(141)) xor (inputs(17)));
    layer0_outputs(7173) <= not((inputs(124)) xor (inputs(137)));
    layer0_outputs(7174) <= (inputs(229)) and not (inputs(63));
    layer0_outputs(7175) <= inputs(198);
    layer0_outputs(7176) <= not((inputs(134)) or (inputs(79)));
    layer0_outputs(7177) <= (inputs(173)) or (inputs(174));
    layer0_outputs(7178) <= not((inputs(187)) or (inputs(188)));
    layer0_outputs(7179) <= not((inputs(248)) or (inputs(102)));
    layer0_outputs(7180) <= not((inputs(243)) xor (inputs(83)));
    layer0_outputs(7181) <= not(inputs(212));
    layer0_outputs(7182) <= not(inputs(101));
    layer0_outputs(7183) <= not((inputs(129)) xor (inputs(19)));
    layer0_outputs(7184) <= (inputs(35)) xor (inputs(96));
    layer0_outputs(7185) <= (inputs(101)) xor (inputs(165));
    layer0_outputs(7186) <= not(inputs(121)) or (inputs(13));
    layer0_outputs(7187) <= not(inputs(27));
    layer0_outputs(7188) <= (inputs(25)) xor (inputs(205));
    layer0_outputs(7189) <= not(inputs(30));
    layer0_outputs(7190) <= (inputs(116)) and not (inputs(159));
    layer0_outputs(7191) <= (inputs(243)) or (inputs(153));
    layer0_outputs(7192) <= not(inputs(69));
    layer0_outputs(7193) <= not(inputs(146));
    layer0_outputs(7194) <= (inputs(73)) and not (inputs(36));
    layer0_outputs(7195) <= inputs(252);
    layer0_outputs(7196) <= inputs(181);
    layer0_outputs(7197) <= not((inputs(171)) or (inputs(3)));
    layer0_outputs(7198) <= not(inputs(39));
    layer0_outputs(7199) <= (inputs(234)) or (inputs(170));
    layer0_outputs(7200) <= not((inputs(122)) xor (inputs(136)));
    layer0_outputs(7201) <= not(inputs(171));
    layer0_outputs(7202) <= not(inputs(166));
    layer0_outputs(7203) <= (inputs(71)) and (inputs(60));
    layer0_outputs(7204) <= inputs(227);
    layer0_outputs(7205) <= not(inputs(104)) or (inputs(192));
    layer0_outputs(7206) <= not(inputs(76));
    layer0_outputs(7207) <= (inputs(150)) and not (inputs(99));
    layer0_outputs(7208) <= inputs(89);
    layer0_outputs(7209) <= (inputs(200)) and not (inputs(78));
    layer0_outputs(7210) <= not(inputs(114));
    layer0_outputs(7211) <= inputs(187);
    layer0_outputs(7212) <= not(inputs(85));
    layer0_outputs(7213) <= not((inputs(84)) or (inputs(174)));
    layer0_outputs(7214) <= inputs(130);
    layer0_outputs(7215) <= (inputs(203)) xor (inputs(251));
    layer0_outputs(7216) <= not(inputs(156));
    layer0_outputs(7217) <= not(inputs(198)) or (inputs(77));
    layer0_outputs(7218) <= not((inputs(251)) or (inputs(85)));
    layer0_outputs(7219) <= not((inputs(119)) and (inputs(138)));
    layer0_outputs(7220) <= not(inputs(179));
    layer0_outputs(7221) <= not((inputs(56)) xor (inputs(27)));
    layer0_outputs(7222) <= inputs(206);
    layer0_outputs(7223) <= not((inputs(119)) or (inputs(29)));
    layer0_outputs(7224) <= not((inputs(81)) xor (inputs(20)));
    layer0_outputs(7225) <= not(inputs(32)) or (inputs(111));
    layer0_outputs(7226) <= (inputs(196)) xor (inputs(133));
    layer0_outputs(7227) <= not(inputs(4));
    layer0_outputs(7228) <= not((inputs(253)) or (inputs(49)));
    layer0_outputs(7229) <= not((inputs(156)) xor (inputs(125)));
    layer0_outputs(7230) <= (inputs(127)) or (inputs(178));
    layer0_outputs(7231) <= (inputs(233)) and not (inputs(58));
    layer0_outputs(7232) <= not(inputs(57)) or (inputs(137));
    layer0_outputs(7233) <= (inputs(15)) xor (inputs(180));
    layer0_outputs(7234) <= not((inputs(102)) or (inputs(220)));
    layer0_outputs(7235) <= not((inputs(101)) xor (inputs(98)));
    layer0_outputs(7236) <= (inputs(181)) and not (inputs(190));
    layer0_outputs(7237) <= (inputs(236)) or (inputs(134));
    layer0_outputs(7238) <= not((inputs(66)) xor (inputs(196)));
    layer0_outputs(7239) <= not((inputs(144)) xor (inputs(115)));
    layer0_outputs(7240) <= (inputs(55)) and (inputs(48));
    layer0_outputs(7241) <= inputs(65);
    layer0_outputs(7242) <= not((inputs(56)) or (inputs(46)));
    layer0_outputs(7243) <= (inputs(151)) and not (inputs(162));
    layer0_outputs(7244) <= not(inputs(109));
    layer0_outputs(7245) <= (inputs(71)) xor (inputs(118));
    layer0_outputs(7246) <= not(inputs(112));
    layer0_outputs(7247) <= not(inputs(159)) or (inputs(129));
    layer0_outputs(7248) <= not(inputs(21)) or (inputs(86));
    layer0_outputs(7249) <= (inputs(175)) or (inputs(113));
    layer0_outputs(7250) <= not(inputs(74));
    layer0_outputs(7251) <= (inputs(11)) and not (inputs(114));
    layer0_outputs(7252) <= inputs(233);
    layer0_outputs(7253) <= not((inputs(7)) xor (inputs(192)));
    layer0_outputs(7254) <= (inputs(170)) and not (inputs(18));
    layer0_outputs(7255) <= inputs(121);
    layer0_outputs(7256) <= not(inputs(97));
    layer0_outputs(7257) <= not((inputs(151)) xor (inputs(186)));
    layer0_outputs(7258) <= inputs(117);
    layer0_outputs(7259) <= (inputs(92)) and not (inputs(52));
    layer0_outputs(7260) <= not(inputs(126)) or (inputs(113));
    layer0_outputs(7261) <= not(inputs(139)) or (inputs(192));
    layer0_outputs(7262) <= (inputs(123)) xor (inputs(149));
    layer0_outputs(7263) <= not(inputs(35)) or (inputs(111));
    layer0_outputs(7264) <= not(inputs(244));
    layer0_outputs(7265) <= not((inputs(193)) xor (inputs(125)));
    layer0_outputs(7266) <= not(inputs(241));
    layer0_outputs(7267) <= not(inputs(127));
    layer0_outputs(7268) <= not(inputs(38)) or (inputs(188));
    layer0_outputs(7269) <= not((inputs(88)) xor (inputs(50)));
    layer0_outputs(7270) <= not(inputs(57));
    layer0_outputs(7271) <= not(inputs(153)) or (inputs(136));
    layer0_outputs(7272) <= (inputs(77)) or (inputs(70));
    layer0_outputs(7273) <= (inputs(94)) and not (inputs(127));
    layer0_outputs(7274) <= (inputs(246)) and not (inputs(242));
    layer0_outputs(7275) <= (inputs(2)) or (inputs(4));
    layer0_outputs(7276) <= (inputs(227)) and not (inputs(79));
    layer0_outputs(7277) <= not(inputs(103)) or (inputs(144));
    layer0_outputs(7278) <= not(inputs(64)) or (inputs(87));
    layer0_outputs(7279) <= not((inputs(76)) or (inputs(255)));
    layer0_outputs(7280) <= not(inputs(206));
    layer0_outputs(7281) <= inputs(144);
    layer0_outputs(7282) <= inputs(168);
    layer0_outputs(7283) <= (inputs(29)) or (inputs(31));
    layer0_outputs(7284) <= (inputs(36)) or (inputs(37));
    layer0_outputs(7285) <= not((inputs(86)) or (inputs(233)));
    layer0_outputs(7286) <= not((inputs(187)) xor (inputs(201)));
    layer0_outputs(7287) <= not((inputs(167)) or (inputs(200)));
    layer0_outputs(7288) <= not((inputs(157)) xor (inputs(240)));
    layer0_outputs(7289) <= not(inputs(78)) or (inputs(227));
    layer0_outputs(7290) <= not(inputs(192));
    layer0_outputs(7291) <= (inputs(53)) or (inputs(255));
    layer0_outputs(7292) <= not(inputs(214));
    layer0_outputs(7293) <= (inputs(228)) or (inputs(81));
    layer0_outputs(7294) <= not(inputs(35));
    layer0_outputs(7295) <= not(inputs(216)) or (inputs(30));
    layer0_outputs(7296) <= inputs(145);
    layer0_outputs(7297) <= not(inputs(138));
    layer0_outputs(7298) <= '1';
    layer0_outputs(7299) <= inputs(174);
    layer0_outputs(7300) <= '0';
    layer0_outputs(7301) <= (inputs(151)) or (inputs(94));
    layer0_outputs(7302) <= not(inputs(88));
    layer0_outputs(7303) <= not((inputs(208)) and (inputs(45)));
    layer0_outputs(7304) <= not(inputs(78));
    layer0_outputs(7305) <= (inputs(100)) xor (inputs(155));
    layer0_outputs(7306) <= not(inputs(149));
    layer0_outputs(7307) <= inputs(104);
    layer0_outputs(7308) <= not((inputs(56)) or (inputs(140)));
    layer0_outputs(7309) <= (inputs(181)) xor (inputs(210));
    layer0_outputs(7310) <= not(inputs(114));
    layer0_outputs(7311) <= not(inputs(197)) or (inputs(105));
    layer0_outputs(7312) <= not(inputs(23));
    layer0_outputs(7313) <= not((inputs(226)) or (inputs(188)));
    layer0_outputs(7314) <= inputs(66);
    layer0_outputs(7315) <= (inputs(5)) or (inputs(135));
    layer0_outputs(7316) <= not(inputs(2)) or (inputs(160));
    layer0_outputs(7317) <= not((inputs(195)) xor (inputs(187)));
    layer0_outputs(7318) <= (inputs(14)) and not (inputs(32));
    layer0_outputs(7319) <= inputs(206);
    layer0_outputs(7320) <= not(inputs(109)) or (inputs(33));
    layer0_outputs(7321) <= inputs(15);
    layer0_outputs(7322) <= (inputs(178)) xor (inputs(80));
    layer0_outputs(7323) <= not((inputs(150)) or (inputs(122)));
    layer0_outputs(7324) <= not((inputs(77)) xor (inputs(18)));
    layer0_outputs(7325) <= (inputs(42)) or (inputs(55));
    layer0_outputs(7326) <= not(inputs(194));
    layer0_outputs(7327) <= not((inputs(106)) or (inputs(97)));
    layer0_outputs(7328) <= not((inputs(147)) or (inputs(151)));
    layer0_outputs(7329) <= not(inputs(165));
    layer0_outputs(7330) <= inputs(75);
    layer0_outputs(7331) <= inputs(170);
    layer0_outputs(7332) <= (inputs(32)) and (inputs(79));
    layer0_outputs(7333) <= (inputs(213)) or (inputs(31));
    layer0_outputs(7334) <= not((inputs(236)) xor (inputs(232)));
    layer0_outputs(7335) <= not((inputs(155)) and (inputs(90)));
    layer0_outputs(7336) <= not(inputs(255));
    layer0_outputs(7337) <= not((inputs(121)) or (inputs(90)));
    layer0_outputs(7338) <= not((inputs(182)) or (inputs(79)));
    layer0_outputs(7339) <= (inputs(139)) and not (inputs(17));
    layer0_outputs(7340) <= not((inputs(127)) or (inputs(82)));
    layer0_outputs(7341) <= not(inputs(199));
    layer0_outputs(7342) <= not(inputs(194));
    layer0_outputs(7343) <= not(inputs(197));
    layer0_outputs(7344) <= not((inputs(151)) and (inputs(41)));
    layer0_outputs(7345) <= (inputs(227)) or (inputs(177));
    layer0_outputs(7346) <= not(inputs(112)) or (inputs(190));
    layer0_outputs(7347) <= not((inputs(35)) or (inputs(9)));
    layer0_outputs(7348) <= not(inputs(100));
    layer0_outputs(7349) <= (inputs(156)) and not (inputs(238));
    layer0_outputs(7350) <= not(inputs(239)) or (inputs(113));
    layer0_outputs(7351) <= (inputs(212)) and not (inputs(178));
    layer0_outputs(7352) <= not((inputs(60)) and (inputs(25)));
    layer0_outputs(7353) <= '1';
    layer0_outputs(7354) <= not((inputs(213)) or (inputs(249)));
    layer0_outputs(7355) <= not((inputs(184)) or (inputs(3)));
    layer0_outputs(7356) <= not(inputs(211)) or (inputs(0));
    layer0_outputs(7357) <= (inputs(231)) xor (inputs(165));
    layer0_outputs(7358) <= inputs(131);
    layer0_outputs(7359) <= not((inputs(135)) or (inputs(181)));
    layer0_outputs(7360) <= (inputs(32)) or (inputs(188));
    layer0_outputs(7361) <= not((inputs(142)) or (inputs(162)));
    layer0_outputs(7362) <= not(inputs(205)) or (inputs(2));
    layer0_outputs(7363) <= inputs(247);
    layer0_outputs(7364) <= not(inputs(42)) or (inputs(184));
    layer0_outputs(7365) <= (inputs(119)) or (inputs(94));
    layer0_outputs(7366) <= not(inputs(138)) or (inputs(235));
    layer0_outputs(7367) <= (inputs(7)) xor (inputs(58));
    layer0_outputs(7368) <= inputs(203);
    layer0_outputs(7369) <= not((inputs(189)) and (inputs(199)));
    layer0_outputs(7370) <= inputs(197);
    layer0_outputs(7371) <= not((inputs(220)) xor (inputs(1)));
    layer0_outputs(7372) <= not(inputs(133));
    layer0_outputs(7373) <= not((inputs(252)) or (inputs(174)));
    layer0_outputs(7374) <= inputs(38);
    layer0_outputs(7375) <= not((inputs(235)) or (inputs(224)));
    layer0_outputs(7376) <= not((inputs(82)) or (inputs(168)));
    layer0_outputs(7377) <= not(inputs(123)) or (inputs(1));
    layer0_outputs(7378) <= not(inputs(172)) or (inputs(64));
    layer0_outputs(7379) <= not(inputs(86));
    layer0_outputs(7380) <= (inputs(85)) and not (inputs(206));
    layer0_outputs(7381) <= (inputs(194)) and not (inputs(159));
    layer0_outputs(7382) <= not((inputs(130)) xor (inputs(53)));
    layer0_outputs(7383) <= not(inputs(114));
    layer0_outputs(7384) <= '0';
    layer0_outputs(7385) <= not(inputs(81)) or (inputs(240));
    layer0_outputs(7386) <= not(inputs(131)) or (inputs(64));
    layer0_outputs(7387) <= (inputs(53)) and not (inputs(243));
    layer0_outputs(7388) <= inputs(120);
    layer0_outputs(7389) <= (inputs(154)) or (inputs(51));
    layer0_outputs(7390) <= not(inputs(129));
    layer0_outputs(7391) <= not((inputs(76)) and (inputs(88)));
    layer0_outputs(7392) <= inputs(214);
    layer0_outputs(7393) <= (inputs(203)) or (inputs(117));
    layer0_outputs(7394) <= not((inputs(168)) xor (inputs(162)));
    layer0_outputs(7395) <= (inputs(33)) or (inputs(50));
    layer0_outputs(7396) <= not((inputs(175)) or (inputs(189)));
    layer0_outputs(7397) <= not((inputs(128)) xor (inputs(197)));
    layer0_outputs(7398) <= (inputs(130)) or (inputs(147));
    layer0_outputs(7399) <= not((inputs(125)) and (inputs(141)));
    layer0_outputs(7400) <= not((inputs(217)) or (inputs(238)));
    layer0_outputs(7401) <= not((inputs(201)) or (inputs(147)));
    layer0_outputs(7402) <= not(inputs(131)) or (inputs(35));
    layer0_outputs(7403) <= not(inputs(110));
    layer0_outputs(7404) <= not(inputs(184)) or (inputs(103));
    layer0_outputs(7405) <= (inputs(133)) and not (inputs(187));
    layer0_outputs(7406) <= not((inputs(35)) or (inputs(2)));
    layer0_outputs(7407) <= (inputs(127)) or (inputs(18));
    layer0_outputs(7408) <= not(inputs(21));
    layer0_outputs(7409) <= not(inputs(137)) or (inputs(127));
    layer0_outputs(7410) <= not(inputs(219));
    layer0_outputs(7411) <= not(inputs(6));
    layer0_outputs(7412) <= not((inputs(172)) xor (inputs(157)));
    layer0_outputs(7413) <= (inputs(72)) and not (inputs(189));
    layer0_outputs(7414) <= not(inputs(239));
    layer0_outputs(7415) <= (inputs(61)) and (inputs(27));
    layer0_outputs(7416) <= inputs(136);
    layer0_outputs(7417) <= (inputs(4)) and not (inputs(173));
    layer0_outputs(7418) <= inputs(123);
    layer0_outputs(7419) <= (inputs(56)) and not (inputs(77));
    layer0_outputs(7420) <= (inputs(248)) or (inputs(60));
    layer0_outputs(7421) <= not(inputs(114)) or (inputs(39));
    layer0_outputs(7422) <= inputs(68);
    layer0_outputs(7423) <= (inputs(234)) or (inputs(50));
    layer0_outputs(7424) <= (inputs(113)) xor (inputs(83));
    layer0_outputs(7425) <= (inputs(73)) and (inputs(183));
    layer0_outputs(7426) <= (inputs(22)) and not (inputs(144));
    layer0_outputs(7427) <= (inputs(228)) and not (inputs(14));
    layer0_outputs(7428) <= inputs(137);
    layer0_outputs(7429) <= inputs(127);
    layer0_outputs(7430) <= (inputs(215)) and not (inputs(1));
    layer0_outputs(7431) <= not(inputs(211)) or (inputs(0));
    layer0_outputs(7432) <= not((inputs(102)) or (inputs(249)));
    layer0_outputs(7433) <= inputs(254);
    layer0_outputs(7434) <= inputs(178);
    layer0_outputs(7435) <= not((inputs(68)) xor (inputs(113)));
    layer0_outputs(7436) <= not((inputs(74)) xor (inputs(129)));
    layer0_outputs(7437) <= not(inputs(18));
    layer0_outputs(7438) <= not((inputs(69)) xor (inputs(128)));
    layer0_outputs(7439) <= (inputs(1)) or (inputs(2));
    layer0_outputs(7440) <= not((inputs(186)) or (inputs(114)));
    layer0_outputs(7441) <= (inputs(175)) or (inputs(250));
    layer0_outputs(7442) <= not((inputs(145)) xor (inputs(138)));
    layer0_outputs(7443) <= (inputs(165)) xor (inputs(167));
    layer0_outputs(7444) <= not(inputs(100)) or (inputs(111));
    layer0_outputs(7445) <= not((inputs(160)) or (inputs(39)));
    layer0_outputs(7446) <= (inputs(90)) and not (inputs(149));
    layer0_outputs(7447) <= (inputs(48)) xor (inputs(94));
    layer0_outputs(7448) <= (inputs(51)) and not (inputs(216));
    layer0_outputs(7449) <= not(inputs(60)) or (inputs(106));
    layer0_outputs(7450) <= not((inputs(231)) or (inputs(57)));
    layer0_outputs(7451) <= not(inputs(150)) or (inputs(213));
    layer0_outputs(7452) <= inputs(207);
    layer0_outputs(7453) <= not(inputs(151));
    layer0_outputs(7454) <= (inputs(77)) or (inputs(77));
    layer0_outputs(7455) <= not((inputs(168)) and (inputs(242)));
    layer0_outputs(7456) <= (inputs(213)) or (inputs(220));
    layer0_outputs(7457) <= '1';
    layer0_outputs(7458) <= not((inputs(226)) xor (inputs(63)));
    layer0_outputs(7459) <= (inputs(79)) xor (inputs(173));
    layer0_outputs(7460) <= (inputs(42)) or (inputs(3));
    layer0_outputs(7461) <= inputs(176);
    layer0_outputs(7462) <= (inputs(236)) xor (inputs(157));
    layer0_outputs(7463) <= not(inputs(178));
    layer0_outputs(7464) <= not((inputs(30)) and (inputs(237)));
    layer0_outputs(7465) <= not(inputs(120));
    layer0_outputs(7466) <= (inputs(194)) or (inputs(132));
    layer0_outputs(7467) <= not(inputs(40));
    layer0_outputs(7468) <= not((inputs(31)) and (inputs(90)));
    layer0_outputs(7469) <= inputs(104);
    layer0_outputs(7470) <= inputs(4);
    layer0_outputs(7471) <= inputs(14);
    layer0_outputs(7472) <= not(inputs(28));
    layer0_outputs(7473) <= not((inputs(108)) or (inputs(220)));
    layer0_outputs(7474) <= not(inputs(199)) or (inputs(172));
    layer0_outputs(7475) <= inputs(246);
    layer0_outputs(7476) <= (inputs(238)) or (inputs(120));
    layer0_outputs(7477) <= (inputs(227)) xor (inputs(226));
    layer0_outputs(7478) <= (inputs(87)) or (inputs(71));
    layer0_outputs(7479) <= not(inputs(96));
    layer0_outputs(7480) <= not((inputs(175)) xor (inputs(84)));
    layer0_outputs(7481) <= inputs(179);
    layer0_outputs(7482) <= not(inputs(103)) or (inputs(128));
    layer0_outputs(7483) <= (inputs(194)) or (inputs(25));
    layer0_outputs(7484) <= (inputs(9)) and not (inputs(2));
    layer0_outputs(7485) <= (inputs(19)) and not (inputs(145));
    layer0_outputs(7486) <= (inputs(109)) and not (inputs(179));
    layer0_outputs(7487) <= not((inputs(25)) or (inputs(162)));
    layer0_outputs(7488) <= not((inputs(23)) xor (inputs(130)));
    layer0_outputs(7489) <= not((inputs(13)) xor (inputs(161)));
    layer0_outputs(7490) <= (inputs(181)) and (inputs(172));
    layer0_outputs(7491) <= (inputs(192)) xor (inputs(180));
    layer0_outputs(7492) <= inputs(128);
    layer0_outputs(7493) <= not(inputs(227)) or (inputs(97));
    layer0_outputs(7494) <= (inputs(199)) or (inputs(65));
    layer0_outputs(7495) <= not(inputs(212)) or (inputs(129));
    layer0_outputs(7496) <= (inputs(5)) xor (inputs(174));
    layer0_outputs(7497) <= inputs(7);
    layer0_outputs(7498) <= not(inputs(58)) or (inputs(95));
    layer0_outputs(7499) <= not(inputs(83)) or (inputs(121));
    layer0_outputs(7500) <= not((inputs(133)) xor (inputs(146)));
    layer0_outputs(7501) <= '0';
    layer0_outputs(7502) <= not(inputs(234));
    layer0_outputs(7503) <= (inputs(144)) or (inputs(147));
    layer0_outputs(7504) <= inputs(15);
    layer0_outputs(7505) <= not(inputs(58)) or (inputs(98));
    layer0_outputs(7506) <= not(inputs(27));
    layer0_outputs(7507) <= not(inputs(66)) or (inputs(235));
    layer0_outputs(7508) <= '0';
    layer0_outputs(7509) <= '1';
    layer0_outputs(7510) <= not((inputs(70)) or (inputs(12)));
    layer0_outputs(7511) <= (inputs(237)) or (inputs(186));
    layer0_outputs(7512) <= not(inputs(148));
    layer0_outputs(7513) <= not(inputs(212));
    layer0_outputs(7514) <= (inputs(134)) and not (inputs(177));
    layer0_outputs(7515) <= not(inputs(247));
    layer0_outputs(7516) <= not(inputs(66));
    layer0_outputs(7517) <= inputs(230);
    layer0_outputs(7518) <= (inputs(15)) or (inputs(57));
    layer0_outputs(7519) <= not(inputs(237)) or (inputs(4));
    layer0_outputs(7520) <= (inputs(251)) and (inputs(199));
    layer0_outputs(7521) <= not(inputs(209));
    layer0_outputs(7522) <= (inputs(35)) and not (inputs(250));
    layer0_outputs(7523) <= (inputs(178)) or (inputs(196));
    layer0_outputs(7524) <= (inputs(112)) or (inputs(168));
    layer0_outputs(7525) <= not(inputs(171)) or (inputs(64));
    layer0_outputs(7526) <= (inputs(5)) or (inputs(218));
    layer0_outputs(7527) <= not(inputs(184)) or (inputs(132));
    layer0_outputs(7528) <= not((inputs(185)) xor (inputs(157)));
    layer0_outputs(7529) <= inputs(191);
    layer0_outputs(7530) <= (inputs(131)) and not (inputs(239));
    layer0_outputs(7531) <= (inputs(100)) and not (inputs(159));
    layer0_outputs(7532) <= not((inputs(34)) or (inputs(207)));
    layer0_outputs(7533) <= inputs(203);
    layer0_outputs(7534) <= (inputs(251)) and not (inputs(243));
    layer0_outputs(7535) <= inputs(100);
    layer0_outputs(7536) <= not(inputs(30)) or (inputs(142));
    layer0_outputs(7537) <= not(inputs(230)) or (inputs(128));
    layer0_outputs(7538) <= (inputs(233)) xor (inputs(154));
    layer0_outputs(7539) <= inputs(225);
    layer0_outputs(7540) <= not(inputs(200)) or (inputs(127));
    layer0_outputs(7541) <= (inputs(21)) or (inputs(241));
    layer0_outputs(7542) <= not(inputs(68)) or (inputs(58));
    layer0_outputs(7543) <= inputs(203);
    layer0_outputs(7544) <= (inputs(22)) and not (inputs(98));
    layer0_outputs(7545) <= not(inputs(117)) or (inputs(19));
    layer0_outputs(7546) <= not((inputs(228)) or (inputs(78)));
    layer0_outputs(7547) <= not(inputs(230)) or (inputs(57));
    layer0_outputs(7548) <= not((inputs(170)) or (inputs(20)));
    layer0_outputs(7549) <= (inputs(129)) xor (inputs(179));
    layer0_outputs(7550) <= (inputs(68)) or (inputs(46));
    layer0_outputs(7551) <= (inputs(76)) and not (inputs(252));
    layer0_outputs(7552) <= (inputs(210)) or (inputs(229));
    layer0_outputs(7553) <= not((inputs(61)) or (inputs(231)));
    layer0_outputs(7554) <= not(inputs(24));
    layer0_outputs(7555) <= not((inputs(131)) or (inputs(94)));
    layer0_outputs(7556) <= not(inputs(219)) or (inputs(146));
    layer0_outputs(7557) <= (inputs(251)) and not (inputs(175));
    layer0_outputs(7558) <= not((inputs(107)) xor (inputs(158)));
    layer0_outputs(7559) <= not((inputs(243)) xor (inputs(196)));
    layer0_outputs(7560) <= (inputs(69)) xor (inputs(71));
    layer0_outputs(7561) <= not(inputs(228)) or (inputs(63));
    layer0_outputs(7562) <= (inputs(109)) and not (inputs(199));
    layer0_outputs(7563) <= not(inputs(20));
    layer0_outputs(7564) <= (inputs(56)) xor (inputs(12));
    layer0_outputs(7565) <= (inputs(255)) xor (inputs(96));
    layer0_outputs(7566) <= (inputs(176)) and not (inputs(210));
    layer0_outputs(7567) <= (inputs(26)) xor (inputs(132));
    layer0_outputs(7568) <= not(inputs(210));
    layer0_outputs(7569) <= (inputs(198)) and not (inputs(89));
    layer0_outputs(7570) <= '1';
    layer0_outputs(7571) <= not((inputs(158)) xor (inputs(222)));
    layer0_outputs(7572) <= (inputs(173)) xor (inputs(120));
    layer0_outputs(7573) <= (inputs(176)) or (inputs(204));
    layer0_outputs(7574) <= not((inputs(92)) xor (inputs(6)));
    layer0_outputs(7575) <= inputs(181);
    layer0_outputs(7576) <= '1';
    layer0_outputs(7577) <= not(inputs(203));
    layer0_outputs(7578) <= inputs(23);
    layer0_outputs(7579) <= (inputs(154)) and not (inputs(57));
    layer0_outputs(7580) <= (inputs(255)) xor (inputs(220));
    layer0_outputs(7581) <= not((inputs(166)) or (inputs(177)));
    layer0_outputs(7582) <= (inputs(102)) xor (inputs(71));
    layer0_outputs(7583) <= not((inputs(60)) and (inputs(18)));
    layer0_outputs(7584) <= not(inputs(24));
    layer0_outputs(7585) <= inputs(56);
    layer0_outputs(7586) <= inputs(136);
    layer0_outputs(7587) <= (inputs(146)) and not (inputs(240));
    layer0_outputs(7588) <= not(inputs(28)) or (inputs(32));
    layer0_outputs(7589) <= (inputs(89)) and not (inputs(8));
    layer0_outputs(7590) <= not(inputs(104)) or (inputs(254));
    layer0_outputs(7591) <= (inputs(141)) and not (inputs(110));
    layer0_outputs(7592) <= inputs(141);
    layer0_outputs(7593) <= not(inputs(85));
    layer0_outputs(7594) <= not((inputs(205)) xor (inputs(176)));
    layer0_outputs(7595) <= not((inputs(249)) xor (inputs(63)));
    layer0_outputs(7596) <= (inputs(149)) xor (inputs(72));
    layer0_outputs(7597) <= (inputs(142)) or (inputs(180));
    layer0_outputs(7598) <= not(inputs(129));
    layer0_outputs(7599) <= (inputs(198)) and not (inputs(186));
    layer0_outputs(7600) <= inputs(109);
    layer0_outputs(7601) <= not((inputs(112)) or (inputs(141)));
    layer0_outputs(7602) <= not((inputs(65)) and (inputs(254)));
    layer0_outputs(7603) <= (inputs(233)) xor (inputs(224));
    layer0_outputs(7604) <= (inputs(195)) or (inputs(193));
    layer0_outputs(7605) <= (inputs(3)) or (inputs(220));
    layer0_outputs(7606) <= not((inputs(181)) xor (inputs(243)));
    layer0_outputs(7607) <= not(inputs(58)) or (inputs(116));
    layer0_outputs(7608) <= (inputs(10)) and not (inputs(31));
    layer0_outputs(7609) <= inputs(202);
    layer0_outputs(7610) <= (inputs(176)) and not (inputs(17));
    layer0_outputs(7611) <= not((inputs(132)) or (inputs(34)));
    layer0_outputs(7612) <= not(inputs(137));
    layer0_outputs(7613) <= not(inputs(41)) or (inputs(253));
    layer0_outputs(7614) <= (inputs(207)) and not (inputs(12));
    layer0_outputs(7615) <= not(inputs(228));
    layer0_outputs(7616) <= (inputs(160)) or (inputs(79));
    layer0_outputs(7617) <= '1';
    layer0_outputs(7618) <= not((inputs(193)) or (inputs(175)));
    layer0_outputs(7619) <= (inputs(251)) or (inputs(93));
    layer0_outputs(7620) <= (inputs(102)) and not (inputs(38));
    layer0_outputs(7621) <= not(inputs(131));
    layer0_outputs(7622) <= '1';
    layer0_outputs(7623) <= (inputs(87)) and not (inputs(129));
    layer0_outputs(7624) <= (inputs(91)) and not (inputs(3));
    layer0_outputs(7625) <= (inputs(249)) and not (inputs(30));
    layer0_outputs(7626) <= (inputs(217)) and not (inputs(113));
    layer0_outputs(7627) <= (inputs(173)) and not (inputs(210));
    layer0_outputs(7628) <= not((inputs(72)) and (inputs(72)));
    layer0_outputs(7629) <= inputs(12);
    layer0_outputs(7630) <= (inputs(133)) or (inputs(168));
    layer0_outputs(7631) <= inputs(151);
    layer0_outputs(7632) <= not(inputs(253));
    layer0_outputs(7633) <= (inputs(74)) or (inputs(1));
    layer0_outputs(7634) <= (inputs(106)) and not (inputs(241));
    layer0_outputs(7635) <= not((inputs(185)) or (inputs(177)));
    layer0_outputs(7636) <= not(inputs(67));
    layer0_outputs(7637) <= (inputs(168)) and not (inputs(32));
    layer0_outputs(7638) <= (inputs(190)) xor (inputs(3));
    layer0_outputs(7639) <= (inputs(146)) or (inputs(180));
    layer0_outputs(7640) <= inputs(102);
    layer0_outputs(7641) <= not((inputs(169)) and (inputs(205)));
    layer0_outputs(7642) <= inputs(108);
    layer0_outputs(7643) <= not(inputs(228));
    layer0_outputs(7644) <= inputs(204);
    layer0_outputs(7645) <= not(inputs(179));
    layer0_outputs(7646) <= not((inputs(127)) or (inputs(17)));
    layer0_outputs(7647) <= not(inputs(249));
    layer0_outputs(7648) <= (inputs(238)) or (inputs(202));
    layer0_outputs(7649) <= inputs(167);
    layer0_outputs(7650) <= inputs(253);
    layer0_outputs(7651) <= not(inputs(130));
    layer0_outputs(7652) <= (inputs(139)) and not (inputs(250));
    layer0_outputs(7653) <= not(inputs(25)) or (inputs(140));
    layer0_outputs(7654) <= (inputs(34)) xor (inputs(142));
    layer0_outputs(7655) <= not(inputs(100));
    layer0_outputs(7656) <= (inputs(8)) or (inputs(213));
    layer0_outputs(7657) <= (inputs(40)) and not (inputs(52));
    layer0_outputs(7658) <= not((inputs(45)) and (inputs(76)));
    layer0_outputs(7659) <= not(inputs(225)) or (inputs(240));
    layer0_outputs(7660) <= not(inputs(20)) or (inputs(97));
    layer0_outputs(7661) <= not(inputs(197)) or (inputs(115));
    layer0_outputs(7662) <= inputs(68);
    layer0_outputs(7663) <= not(inputs(230)) or (inputs(159));
    layer0_outputs(7664) <= not(inputs(135)) or (inputs(195));
    layer0_outputs(7665) <= (inputs(29)) or (inputs(89));
    layer0_outputs(7666) <= (inputs(132)) xor (inputs(183));
    layer0_outputs(7667) <= (inputs(232)) xor (inputs(196));
    layer0_outputs(7668) <= (inputs(84)) or (inputs(14));
    layer0_outputs(7669) <= not((inputs(152)) or (inputs(44)));
    layer0_outputs(7670) <= inputs(58);
    layer0_outputs(7671) <= (inputs(36)) and (inputs(234));
    layer0_outputs(7672) <= (inputs(212)) or (inputs(248));
    layer0_outputs(7673) <= (inputs(32)) xor (inputs(154));
    layer0_outputs(7674) <= (inputs(241)) and not (inputs(201));
    layer0_outputs(7675) <= (inputs(244)) and not (inputs(145));
    layer0_outputs(7676) <= (inputs(135)) and not (inputs(128));
    layer0_outputs(7677) <= (inputs(105)) and not (inputs(21));
    layer0_outputs(7678) <= not((inputs(15)) xor (inputs(48)));
    layer0_outputs(7679) <= not((inputs(111)) or (inputs(20)));
    outputs(0) <= not((layer0_outputs(4399)) and (layer0_outputs(5849)));
    outputs(1) <= layer0_outputs(4522);
    outputs(2) <= (layer0_outputs(343)) and not (layer0_outputs(6502));
    outputs(3) <= (layer0_outputs(1500)) and not (layer0_outputs(3689));
    outputs(4) <= (layer0_outputs(5387)) and not (layer0_outputs(1181));
    outputs(5) <= layer0_outputs(4574);
    outputs(6) <= not((layer0_outputs(3161)) xor (layer0_outputs(222)));
    outputs(7) <= layer0_outputs(5951);
    outputs(8) <= (layer0_outputs(2212)) xor (layer0_outputs(203));
    outputs(9) <= not((layer0_outputs(3119)) xor (layer0_outputs(748)));
    outputs(10) <= layer0_outputs(5965);
    outputs(11) <= layer0_outputs(3979);
    outputs(12) <= layer0_outputs(7604);
    outputs(13) <= layer0_outputs(3361);
    outputs(14) <= layer0_outputs(441);
    outputs(15) <= not(layer0_outputs(983));
    outputs(16) <= not(layer0_outputs(2145)) or (layer0_outputs(2469));
    outputs(17) <= not(layer0_outputs(3785)) or (layer0_outputs(1627));
    outputs(18) <= (layer0_outputs(2039)) xor (layer0_outputs(2496));
    outputs(19) <= not((layer0_outputs(5368)) and (layer0_outputs(248)));
    outputs(20) <= not(layer0_outputs(6096));
    outputs(21) <= (layer0_outputs(7107)) or (layer0_outputs(6917));
    outputs(22) <= not(layer0_outputs(4241));
    outputs(23) <= layer0_outputs(1126);
    outputs(24) <= layer0_outputs(675);
    outputs(25) <= not((layer0_outputs(3935)) or (layer0_outputs(2618)));
    outputs(26) <= not((layer0_outputs(3184)) and (layer0_outputs(6535)));
    outputs(27) <= not((layer0_outputs(4326)) and (layer0_outputs(3446)));
    outputs(28) <= layer0_outputs(783);
    outputs(29) <= layer0_outputs(6346);
    outputs(30) <= not((layer0_outputs(4750)) xor (layer0_outputs(7432)));
    outputs(31) <= not(layer0_outputs(5980));
    outputs(32) <= (layer0_outputs(2783)) xor (layer0_outputs(5750));
    outputs(33) <= (layer0_outputs(1910)) xor (layer0_outputs(5961));
    outputs(34) <= layer0_outputs(1466);
    outputs(35) <= not((layer0_outputs(4659)) and (layer0_outputs(2522)));
    outputs(36) <= not(layer0_outputs(3684)) or (layer0_outputs(3312));
    outputs(37) <= layer0_outputs(6021);
    outputs(38) <= not(layer0_outputs(6580));
    outputs(39) <= not(layer0_outputs(5765));
    outputs(40) <= layer0_outputs(2284);
    outputs(41) <= (layer0_outputs(4619)) and not (layer0_outputs(142));
    outputs(42) <= not(layer0_outputs(3471));
    outputs(43) <= (layer0_outputs(1490)) and (layer0_outputs(3331));
    outputs(44) <= layer0_outputs(3644);
    outputs(45) <= not((layer0_outputs(3813)) and (layer0_outputs(3664)));
    outputs(46) <= not(layer0_outputs(6405));
    outputs(47) <= layer0_outputs(3339);
    outputs(48) <= (layer0_outputs(3283)) and not (layer0_outputs(166));
    outputs(49) <= not((layer0_outputs(1218)) or (layer0_outputs(4650)));
    outputs(50) <= not((layer0_outputs(6926)) and (layer0_outputs(2923)));
    outputs(51) <= (layer0_outputs(2755)) and not (layer0_outputs(3135));
    outputs(52) <= not(layer0_outputs(7064)) or (layer0_outputs(6558));
    outputs(53) <= layer0_outputs(2089);
    outputs(54) <= not(layer0_outputs(3689));
    outputs(55) <= (layer0_outputs(2489)) and not (layer0_outputs(7508));
    outputs(56) <= layer0_outputs(1677);
    outputs(57) <= layer0_outputs(3280);
    outputs(58) <= (layer0_outputs(6691)) and not (layer0_outputs(5390));
    outputs(59) <= (layer0_outputs(5047)) and (layer0_outputs(228));
    outputs(60) <= layer0_outputs(4445);
    outputs(61) <= not(layer0_outputs(7262));
    outputs(62) <= not(layer0_outputs(2595)) or (layer0_outputs(3375));
    outputs(63) <= (layer0_outputs(4726)) and not (layer0_outputs(2889));
    outputs(64) <= not(layer0_outputs(4177));
    outputs(65) <= (layer0_outputs(291)) or (layer0_outputs(7159));
    outputs(66) <= (layer0_outputs(4132)) and not (layer0_outputs(678));
    outputs(67) <= layer0_outputs(635);
    outputs(68) <= (layer0_outputs(7617)) and (layer0_outputs(6453));
    outputs(69) <= not(layer0_outputs(4502)) or (layer0_outputs(2500));
    outputs(70) <= not((layer0_outputs(7279)) and (layer0_outputs(7403)));
    outputs(71) <= layer0_outputs(7157);
    outputs(72) <= layer0_outputs(7447);
    outputs(73) <= layer0_outputs(5640);
    outputs(74) <= not((layer0_outputs(3067)) and (layer0_outputs(1676)));
    outputs(75) <= (layer0_outputs(5756)) and not (layer0_outputs(6047));
    outputs(76) <= not(layer0_outputs(566)) or (layer0_outputs(927));
    outputs(77) <= layer0_outputs(5796);
    outputs(78) <= layer0_outputs(4459);
    outputs(79) <= (layer0_outputs(6059)) xor (layer0_outputs(6821));
    outputs(80) <= (layer0_outputs(6224)) xor (layer0_outputs(2685));
    outputs(81) <= layer0_outputs(4639);
    outputs(82) <= not(layer0_outputs(3926)) or (layer0_outputs(3129));
    outputs(83) <= layer0_outputs(2152);
    outputs(84) <= (layer0_outputs(491)) and not (layer0_outputs(6913));
    outputs(85) <= not(layer0_outputs(7631));
    outputs(86) <= (layer0_outputs(5237)) and (layer0_outputs(7136));
    outputs(87) <= (layer0_outputs(7325)) and (layer0_outputs(5230));
    outputs(88) <= not(layer0_outputs(3136));
    outputs(89) <= not(layer0_outputs(2737)) or (layer0_outputs(7214));
    outputs(90) <= (layer0_outputs(1933)) or (layer0_outputs(1809));
    outputs(91) <= not(layer0_outputs(4454));
    outputs(92) <= (layer0_outputs(4343)) and (layer0_outputs(5606));
    outputs(93) <= not(layer0_outputs(2538));
    outputs(94) <= not((layer0_outputs(7399)) and (layer0_outputs(3529)));
    outputs(95) <= (layer0_outputs(2464)) or (layer0_outputs(5205));
    outputs(96) <= layer0_outputs(3412);
    outputs(97) <= layer0_outputs(2970);
    outputs(98) <= layer0_outputs(3127);
    outputs(99) <= layer0_outputs(6088);
    outputs(100) <= (layer0_outputs(3231)) and (layer0_outputs(237));
    outputs(101) <= not(layer0_outputs(3051));
    outputs(102) <= not(layer0_outputs(6568));
    outputs(103) <= not((layer0_outputs(546)) xor (layer0_outputs(7050)));
    outputs(104) <= (layer0_outputs(1603)) or (layer0_outputs(4974));
    outputs(105) <= not(layer0_outputs(3456));
    outputs(106) <= not(layer0_outputs(7416));
    outputs(107) <= layer0_outputs(2129);
    outputs(108) <= not(layer0_outputs(2909)) or (layer0_outputs(2867));
    outputs(109) <= not(layer0_outputs(6385));
    outputs(110) <= not(layer0_outputs(5930));
    outputs(111) <= layer0_outputs(2211);
    outputs(112) <= not((layer0_outputs(5203)) xor (layer0_outputs(1976)));
    outputs(113) <= layer0_outputs(1534);
    outputs(114) <= (layer0_outputs(1328)) and not (layer0_outputs(1894));
    outputs(115) <= not(layer0_outputs(2186));
    outputs(116) <= not(layer0_outputs(4438));
    outputs(117) <= (layer0_outputs(3946)) and (layer0_outputs(6877));
    outputs(118) <= (layer0_outputs(4346)) or (layer0_outputs(1673));
    outputs(119) <= not(layer0_outputs(3922)) or (layer0_outputs(931));
    outputs(120) <= (layer0_outputs(2353)) xor (layer0_outputs(4628));
    outputs(121) <= not(layer0_outputs(1539)) or (layer0_outputs(4012));
    outputs(122) <= not(layer0_outputs(2326)) or (layer0_outputs(5569));
    outputs(123) <= not((layer0_outputs(2016)) or (layer0_outputs(999)));
    outputs(124) <= not(layer0_outputs(6318));
    outputs(125) <= layer0_outputs(4571);
    outputs(126) <= layer0_outputs(5387);
    outputs(127) <= not(layer0_outputs(331));
    outputs(128) <= (layer0_outputs(7165)) xor (layer0_outputs(4134));
    outputs(129) <= layer0_outputs(389);
    outputs(130) <= (layer0_outputs(3485)) and (layer0_outputs(7008));
    outputs(131) <= layer0_outputs(7228);
    outputs(132) <= not((layer0_outputs(6642)) and (layer0_outputs(422)));
    outputs(133) <= not(layer0_outputs(289));
    outputs(134) <= (layer0_outputs(2149)) and not (layer0_outputs(3107));
    outputs(135) <= not((layer0_outputs(4519)) and (layer0_outputs(6784)));
    outputs(136) <= not(layer0_outputs(4252));
    outputs(137) <= not(layer0_outputs(6393));
    outputs(138) <= not((layer0_outputs(3401)) and (layer0_outputs(6967)));
    outputs(139) <= not(layer0_outputs(1750)) or (layer0_outputs(844));
    outputs(140) <= (layer0_outputs(6238)) xor (layer0_outputs(6331));
    outputs(141) <= (layer0_outputs(6899)) or (layer0_outputs(4362));
    outputs(142) <= (layer0_outputs(3516)) or (layer0_outputs(72));
    outputs(143) <= not(layer0_outputs(980));
    outputs(144) <= (layer0_outputs(1551)) xor (layer0_outputs(2127));
    outputs(145) <= (layer0_outputs(5629)) xor (layer0_outputs(650));
    outputs(146) <= not(layer0_outputs(360));
    outputs(147) <= not(layer0_outputs(619));
    outputs(148) <= not(layer0_outputs(6552));
    outputs(149) <= not(layer0_outputs(5498));
    outputs(150) <= not(layer0_outputs(5808));
    outputs(151) <= not(layer0_outputs(195));
    outputs(152) <= (layer0_outputs(3960)) and (layer0_outputs(525));
    outputs(153) <= not((layer0_outputs(4992)) or (layer0_outputs(6488)));
    outputs(154) <= layer0_outputs(2547);
    outputs(155) <= not(layer0_outputs(6487)) or (layer0_outputs(7427));
    outputs(156) <= (layer0_outputs(7097)) xor (layer0_outputs(3357));
    outputs(157) <= not(layer0_outputs(2677));
    outputs(158) <= not((layer0_outputs(6704)) xor (layer0_outputs(6404)));
    outputs(159) <= layer0_outputs(5989);
    outputs(160) <= not((layer0_outputs(3157)) or (layer0_outputs(84)));
    outputs(161) <= not(layer0_outputs(3141));
    outputs(162) <= layer0_outputs(762);
    outputs(163) <= layer0_outputs(6917);
    outputs(164) <= (layer0_outputs(6386)) xor (layer0_outputs(5564));
    outputs(165) <= not((layer0_outputs(7127)) xor (layer0_outputs(162)));
    outputs(166) <= not(layer0_outputs(7012));
    outputs(167) <= not((layer0_outputs(7499)) and (layer0_outputs(7402)));
    outputs(168) <= (layer0_outputs(4496)) or (layer0_outputs(6733));
    outputs(169) <= (layer0_outputs(1829)) xor (layer0_outputs(7327));
    outputs(170) <= layer0_outputs(4630);
    outputs(171) <= not(layer0_outputs(1518));
    outputs(172) <= not(layer0_outputs(2788));
    outputs(173) <= not(layer0_outputs(5253)) or (layer0_outputs(2680));
    outputs(174) <= not((layer0_outputs(7441)) xor (layer0_outputs(3300)));
    outputs(175) <= not(layer0_outputs(902));
    outputs(176) <= not((layer0_outputs(6555)) or (layer0_outputs(2781)));
    outputs(177) <= not((layer0_outputs(3317)) or (layer0_outputs(6126)));
    outputs(178) <= not((layer0_outputs(5904)) and (layer0_outputs(1413)));
    outputs(179) <= not(layer0_outputs(145));
    outputs(180) <= not(layer0_outputs(2246));
    outputs(181) <= layer0_outputs(2740);
    outputs(182) <= layer0_outputs(1583);
    outputs(183) <= not((layer0_outputs(3043)) and (layer0_outputs(7335)));
    outputs(184) <= (layer0_outputs(3048)) and not (layer0_outputs(2856));
    outputs(185) <= not(layer0_outputs(4455));
    outputs(186) <= layer0_outputs(6028);
    outputs(187) <= not(layer0_outputs(3802));
    outputs(188) <= not((layer0_outputs(5364)) xor (layer0_outputs(499)));
    outputs(189) <= not(layer0_outputs(4105));
    outputs(190) <= not(layer0_outputs(1520)) or (layer0_outputs(3037));
    outputs(191) <= (layer0_outputs(2557)) or (layer0_outputs(4416));
    outputs(192) <= (layer0_outputs(1886)) and not (layer0_outputs(4540));
    outputs(193) <= not(layer0_outputs(4131)) or (layer0_outputs(1873));
    outputs(194) <= not((layer0_outputs(5440)) and (layer0_outputs(6813)));
    outputs(195) <= (layer0_outputs(3523)) xor (layer0_outputs(7343));
    outputs(196) <= layer0_outputs(2103);
    outputs(197) <= not(layer0_outputs(2626));
    outputs(198) <= not((layer0_outputs(4663)) xor (layer0_outputs(412)));
    outputs(199) <= not(layer0_outputs(364)) or (layer0_outputs(6262));
    outputs(200) <= not((layer0_outputs(484)) xor (layer0_outputs(4973)));
    outputs(201) <= not(layer0_outputs(5627));
    outputs(202) <= (layer0_outputs(4382)) xor (layer0_outputs(3777));
    outputs(203) <= not(layer0_outputs(4990));
    outputs(204) <= layer0_outputs(2425);
    outputs(205) <= (layer0_outputs(245)) and not (layer0_outputs(6713));
    outputs(206) <= (layer0_outputs(3398)) or (layer0_outputs(2257));
    outputs(207) <= not((layer0_outputs(6644)) or (layer0_outputs(6551)));
    outputs(208) <= not(layer0_outputs(3529));
    outputs(209) <= layer0_outputs(7323);
    outputs(210) <= (layer0_outputs(5755)) and not (layer0_outputs(3947));
    outputs(211) <= not((layer0_outputs(6275)) xor (layer0_outputs(2474)));
    outputs(212) <= not((layer0_outputs(5356)) xor (layer0_outputs(4151)));
    outputs(213) <= not(layer0_outputs(1151));
    outputs(214) <= not(layer0_outputs(6818));
    outputs(215) <= not(layer0_outputs(4364));
    outputs(216) <= not(layer0_outputs(4483));
    outputs(217) <= not((layer0_outputs(60)) or (layer0_outputs(5793)));
    outputs(218) <= (layer0_outputs(2553)) and not (layer0_outputs(990));
    outputs(219) <= not((layer0_outputs(1441)) or (layer0_outputs(5343)));
    outputs(220) <= layer0_outputs(62);
    outputs(221) <= not((layer0_outputs(619)) or (layer0_outputs(4270)));
    outputs(222) <= (layer0_outputs(7568)) xor (layer0_outputs(3926));
    outputs(223) <= not(layer0_outputs(7120));
    outputs(224) <= layer0_outputs(4577);
    outputs(225) <= layer0_outputs(4262);
    outputs(226) <= not(layer0_outputs(2582));
    outputs(227) <= not((layer0_outputs(2357)) or (layer0_outputs(3302)));
    outputs(228) <= not(layer0_outputs(2936));
    outputs(229) <= layer0_outputs(5990);
    outputs(230) <= not(layer0_outputs(6896));
    outputs(231) <= not((layer0_outputs(5489)) or (layer0_outputs(302)));
    outputs(232) <= layer0_outputs(5246);
    outputs(233) <= layer0_outputs(4371);
    outputs(234) <= layer0_outputs(6991);
    outputs(235) <= (layer0_outputs(6641)) and (layer0_outputs(2655));
    outputs(236) <= (layer0_outputs(6904)) xor (layer0_outputs(4722));
    outputs(237) <= not(layer0_outputs(7426));
    outputs(238) <= not(layer0_outputs(430)) or (layer0_outputs(1568));
    outputs(239) <= not((layer0_outputs(4483)) and (layer0_outputs(4309)));
    outputs(240) <= (layer0_outputs(4524)) xor (layer0_outputs(6505));
    outputs(241) <= not(layer0_outputs(1957));
    outputs(242) <= not(layer0_outputs(2536));
    outputs(243) <= not((layer0_outputs(1173)) or (layer0_outputs(7614)));
    outputs(244) <= not(layer0_outputs(3102));
    outputs(245) <= (layer0_outputs(1096)) and (layer0_outputs(1773));
    outputs(246) <= not(layer0_outputs(7522)) or (layer0_outputs(6732));
    outputs(247) <= (layer0_outputs(5897)) and not (layer0_outputs(4497));
    outputs(248) <= not((layer0_outputs(2185)) xor (layer0_outputs(3835)));
    outputs(249) <= not((layer0_outputs(2762)) xor (layer0_outputs(6992)));
    outputs(250) <= (layer0_outputs(2197)) and not (layer0_outputs(4684));
    outputs(251) <= not(layer0_outputs(2790));
    outputs(252) <= not((layer0_outputs(1805)) xor (layer0_outputs(6225)));
    outputs(253) <= (layer0_outputs(3845)) and (layer0_outputs(3198));
    outputs(254) <= not((layer0_outputs(3859)) xor (layer0_outputs(4641)));
    outputs(255) <= not(layer0_outputs(5573));
    outputs(256) <= (layer0_outputs(2847)) and not (layer0_outputs(3039));
    outputs(257) <= layer0_outputs(6738);
    outputs(258) <= layer0_outputs(4754);
    outputs(259) <= (layer0_outputs(4686)) and not (layer0_outputs(6022));
    outputs(260) <= layer0_outputs(4316);
    outputs(261) <= not(layer0_outputs(6221));
    outputs(262) <= layer0_outputs(3912);
    outputs(263) <= not((layer0_outputs(5439)) xor (layer0_outputs(4523)));
    outputs(264) <= layer0_outputs(3657);
    outputs(265) <= layer0_outputs(651);
    outputs(266) <= (layer0_outputs(6194)) or (layer0_outputs(7380));
    outputs(267) <= not(layer0_outputs(3419)) or (layer0_outputs(5455));
    outputs(268) <= layer0_outputs(4147);
    outputs(269) <= layer0_outputs(3822);
    outputs(270) <= (layer0_outputs(3114)) or (layer0_outputs(3596));
    outputs(271) <= not((layer0_outputs(1998)) xor (layer0_outputs(1507)));
    outputs(272) <= layer0_outputs(7488);
    outputs(273) <= (layer0_outputs(4604)) and not (layer0_outputs(2806));
    outputs(274) <= not((layer0_outputs(1908)) or (layer0_outputs(381)));
    outputs(275) <= layer0_outputs(6649);
    outputs(276) <= not((layer0_outputs(3199)) xor (layer0_outputs(976)));
    outputs(277) <= layer0_outputs(6494);
    outputs(278) <= layer0_outputs(1433);
    outputs(279) <= (layer0_outputs(6432)) xor (layer0_outputs(3941));
    outputs(280) <= not(layer0_outputs(3592));
    outputs(281) <= not((layer0_outputs(5398)) xor (layer0_outputs(5504)));
    outputs(282) <= not(layer0_outputs(5681));
    outputs(283) <= not((layer0_outputs(7648)) xor (layer0_outputs(45)));
    outputs(284) <= not(layer0_outputs(5759));
    outputs(285) <= (layer0_outputs(2454)) and (layer0_outputs(7375));
    outputs(286) <= not(layer0_outputs(1047));
    outputs(287) <= layer0_outputs(6473);
    outputs(288) <= not(layer0_outputs(314));
    outputs(289) <= layer0_outputs(7044);
    outputs(290) <= not(layer0_outputs(2641)) or (layer0_outputs(5985));
    outputs(291) <= not(layer0_outputs(7091));
    outputs(292) <= not(layer0_outputs(6271));
    outputs(293) <= not(layer0_outputs(239));
    outputs(294) <= not(layer0_outputs(381));
    outputs(295) <= not(layer0_outputs(685));
    outputs(296) <= not(layer0_outputs(4479));
    outputs(297) <= (layer0_outputs(5916)) and not (layer0_outputs(1275));
    outputs(298) <= not((layer0_outputs(3952)) xor (layer0_outputs(230)));
    outputs(299) <= not(layer0_outputs(5407));
    outputs(300) <= not((layer0_outputs(3043)) or (layer0_outputs(6796)));
    outputs(301) <= not((layer0_outputs(879)) or (layer0_outputs(7158)));
    outputs(302) <= (layer0_outputs(5223)) and not (layer0_outputs(2336));
    outputs(303) <= layer0_outputs(3166);
    outputs(304) <= not(layer0_outputs(3976));
    outputs(305) <= layer0_outputs(931);
    outputs(306) <= layer0_outputs(1493);
    outputs(307) <= not(layer0_outputs(6282));
    outputs(308) <= not((layer0_outputs(4626)) and (layer0_outputs(5389)));
    outputs(309) <= (layer0_outputs(571)) and (layer0_outputs(3649));
    outputs(310) <= not(layer0_outputs(2881)) or (layer0_outputs(6278));
    outputs(311) <= (layer0_outputs(2225)) and not (layer0_outputs(1591));
    outputs(312) <= not(layer0_outputs(5779));
    outputs(313) <= not(layer0_outputs(7256)) or (layer0_outputs(6370));
    outputs(314) <= layer0_outputs(2796);
    outputs(315) <= (layer0_outputs(3161)) xor (layer0_outputs(7169));
    outputs(316) <= (layer0_outputs(3901)) and not (layer0_outputs(7494));
    outputs(317) <= (layer0_outputs(4267)) or (layer0_outputs(693));
    outputs(318) <= not((layer0_outputs(1542)) xor (layer0_outputs(2663)));
    outputs(319) <= (layer0_outputs(1898)) xor (layer0_outputs(58));
    outputs(320) <= not(layer0_outputs(6394));
    outputs(321) <= not(layer0_outputs(4979)) or (layer0_outputs(2625));
    outputs(322) <= not((layer0_outputs(6454)) and (layer0_outputs(3455)));
    outputs(323) <= layer0_outputs(2655);
    outputs(324) <= (layer0_outputs(6836)) or (layer0_outputs(1384));
    outputs(325) <= (layer0_outputs(5525)) and not (layer0_outputs(3457));
    outputs(326) <= not(layer0_outputs(3537));
    outputs(327) <= layer0_outputs(2872);
    outputs(328) <= not(layer0_outputs(7237));
    outputs(329) <= not(layer0_outputs(5197));
    outputs(330) <= layer0_outputs(1277);
    outputs(331) <= not((layer0_outputs(7341)) xor (layer0_outputs(6766)));
    outputs(332) <= not(layer0_outputs(1114));
    outputs(333) <= not((layer0_outputs(7014)) or (layer0_outputs(1238)));
    outputs(334) <= layer0_outputs(6678);
    outputs(335) <= (layer0_outputs(1487)) and not (layer0_outputs(2679));
    outputs(336) <= (layer0_outputs(5684)) and not (layer0_outputs(4248));
    outputs(337) <= layer0_outputs(7287);
    outputs(338) <= not(layer0_outputs(3666));
    outputs(339) <= (layer0_outputs(3677)) xor (layer0_outputs(5885));
    outputs(340) <= not(layer0_outputs(5773));
    outputs(341) <= layer0_outputs(4264);
    outputs(342) <= layer0_outputs(7146);
    outputs(343) <= not(layer0_outputs(5049));
    outputs(344) <= not((layer0_outputs(4813)) xor (layer0_outputs(5029)));
    outputs(345) <= layer0_outputs(3933);
    outputs(346) <= layer0_outputs(6923);
    outputs(347) <= not((layer0_outputs(5319)) or (layer0_outputs(3956)));
    outputs(348) <= (layer0_outputs(6304)) or (layer0_outputs(478));
    outputs(349) <= not((layer0_outputs(6733)) xor (layer0_outputs(7216)));
    outputs(350) <= not(layer0_outputs(4804));
    outputs(351) <= not(layer0_outputs(3106));
    outputs(352) <= layer0_outputs(2957);
    outputs(353) <= (layer0_outputs(4236)) and (layer0_outputs(4188));
    outputs(354) <= layer0_outputs(3518);
    outputs(355) <= layer0_outputs(3188);
    outputs(356) <= (layer0_outputs(1102)) and not (layer0_outputs(3703));
    outputs(357) <= not(layer0_outputs(6810));
    outputs(358) <= not((layer0_outputs(4568)) and (layer0_outputs(1038)));
    outputs(359) <= not((layer0_outputs(1840)) or (layer0_outputs(5247)));
    outputs(360) <= not(layer0_outputs(2599));
    outputs(361) <= (layer0_outputs(6085)) and not (layer0_outputs(535));
    outputs(362) <= not(layer0_outputs(4871)) or (layer0_outputs(7016));
    outputs(363) <= not(layer0_outputs(5161));
    outputs(364) <= not((layer0_outputs(3808)) xor (layer0_outputs(2744)));
    outputs(365) <= not(layer0_outputs(2158));
    outputs(366) <= not(layer0_outputs(4055)) or (layer0_outputs(3190));
    outputs(367) <= layer0_outputs(7083);
    outputs(368) <= layer0_outputs(5495);
    outputs(369) <= (layer0_outputs(2807)) and not (layer0_outputs(4988));
    outputs(370) <= not((layer0_outputs(4323)) and (layer0_outputs(987)));
    outputs(371) <= not(layer0_outputs(1381)) or (layer0_outputs(4280));
    outputs(372) <= (layer0_outputs(117)) and not (layer0_outputs(1657));
    outputs(373) <= not((layer0_outputs(2954)) xor (layer0_outputs(1586)));
    outputs(374) <= not(layer0_outputs(3409)) or (layer0_outputs(5866));
    outputs(375) <= layer0_outputs(2671);
    outputs(376) <= layer0_outputs(2144);
    outputs(377) <= (layer0_outputs(4326)) xor (layer0_outputs(3772));
    outputs(378) <= not(layer0_outputs(4017));
    outputs(379) <= not(layer0_outputs(5823)) or (layer0_outputs(6808));
    outputs(380) <= layer0_outputs(7664);
    outputs(381) <= not(layer0_outputs(534)) or (layer0_outputs(5857));
    outputs(382) <= layer0_outputs(6932);
    outputs(383) <= not(layer0_outputs(3848)) or (layer0_outputs(2207));
    outputs(384) <= not((layer0_outputs(6624)) and (layer0_outputs(4320)));
    outputs(385) <= not(layer0_outputs(5379));
    outputs(386) <= not((layer0_outputs(1182)) and (layer0_outputs(4100)));
    outputs(387) <= not((layer0_outputs(5945)) and (layer0_outputs(1403)));
    outputs(388) <= not(layer0_outputs(5627));
    outputs(389) <= layer0_outputs(7323);
    outputs(390) <= (layer0_outputs(2053)) and not (layer0_outputs(2733));
    outputs(391) <= (layer0_outputs(804)) or (layer0_outputs(5811));
    outputs(392) <= not(layer0_outputs(1512));
    outputs(393) <= (layer0_outputs(6482)) and not (layer0_outputs(4171));
    outputs(394) <= not(layer0_outputs(942)) or (layer0_outputs(3797));
    outputs(395) <= layer0_outputs(7551);
    outputs(396) <= (layer0_outputs(2961)) or (layer0_outputs(5692));
    outputs(397) <= not(layer0_outputs(3288)) or (layer0_outputs(3731));
    outputs(398) <= not(layer0_outputs(2842));
    outputs(399) <= not(layer0_outputs(4437));
    outputs(400) <= layer0_outputs(6984);
    outputs(401) <= (layer0_outputs(2563)) and (layer0_outputs(1448));
    outputs(402) <= not(layer0_outputs(7270)) or (layer0_outputs(1271));
    outputs(403) <= not((layer0_outputs(155)) or (layer0_outputs(4570)));
    outputs(404) <= not(layer0_outputs(269));
    outputs(405) <= not(layer0_outputs(4845));
    outputs(406) <= not((layer0_outputs(883)) and (layer0_outputs(1112)));
    outputs(407) <= layer0_outputs(5944);
    outputs(408) <= (layer0_outputs(2940)) and (layer0_outputs(5403));
    outputs(409) <= not(layer0_outputs(4082));
    outputs(410) <= not(layer0_outputs(1505));
    outputs(411) <= layer0_outputs(2649);
    outputs(412) <= (layer0_outputs(3982)) and not (layer0_outputs(577));
    outputs(413) <= not(layer0_outputs(5148)) or (layer0_outputs(4344));
    outputs(414) <= not((layer0_outputs(1227)) or (layer0_outputs(6961)));
    outputs(415) <= not(layer0_outputs(1308));
    outputs(416) <= not(layer0_outputs(4487));
    outputs(417) <= not(layer0_outputs(3750));
    outputs(418) <= not((layer0_outputs(4557)) xor (layer0_outputs(4239)));
    outputs(419) <= layer0_outputs(2279);
    outputs(420) <= not(layer0_outputs(4376));
    outputs(421) <= not(layer0_outputs(4853));
    outputs(422) <= (layer0_outputs(6662)) or (layer0_outputs(2287));
    outputs(423) <= layer0_outputs(5027);
    outputs(424) <= (layer0_outputs(5165)) xor (layer0_outputs(7053));
    outputs(425) <= not(layer0_outputs(2417));
    outputs(426) <= layer0_outputs(4808);
    outputs(427) <= (layer0_outputs(2714)) or (layer0_outputs(5703));
    outputs(428) <= layer0_outputs(3251);
    outputs(429) <= not((layer0_outputs(6518)) or (layer0_outputs(1138)));
    outputs(430) <= not((layer0_outputs(2023)) and (layer0_outputs(1175)));
    outputs(431) <= not(layer0_outputs(2429));
    outputs(432) <= not(layer0_outputs(4079));
    outputs(433) <= not(layer0_outputs(1368)) or (layer0_outputs(1601));
    outputs(434) <= not(layer0_outputs(2338));
    outputs(435) <= not(layer0_outputs(7596));
    outputs(436) <= layer0_outputs(2104);
    outputs(437) <= not(layer0_outputs(2164));
    outputs(438) <= layer0_outputs(4338);
    outputs(439) <= not((layer0_outputs(378)) xor (layer0_outputs(7028)));
    outputs(440) <= not(layer0_outputs(5591));
    outputs(441) <= layer0_outputs(2650);
    outputs(442) <= (layer0_outputs(6142)) xor (layer0_outputs(1103));
    outputs(443) <= not(layer0_outputs(6126));
    outputs(444) <= layer0_outputs(1902);
    outputs(445) <= not(layer0_outputs(5948));
    outputs(446) <= (layer0_outputs(273)) and (layer0_outputs(720));
    outputs(447) <= not((layer0_outputs(7328)) xor (layer0_outputs(5906)));
    outputs(448) <= layer0_outputs(6696);
    outputs(449) <= (layer0_outputs(3482)) or (layer0_outputs(1818));
    outputs(450) <= not(layer0_outputs(5784)) or (layer0_outputs(383));
    outputs(451) <= not((layer0_outputs(7528)) or (layer0_outputs(473)));
    outputs(452) <= layer0_outputs(1244);
    outputs(453) <= not((layer0_outputs(6825)) xor (layer0_outputs(464)));
    outputs(454) <= not(layer0_outputs(6714));
    outputs(455) <= not(layer0_outputs(458));
    outputs(456) <= (layer0_outputs(1705)) and not (layer0_outputs(6328));
    outputs(457) <= (layer0_outputs(2589)) xor (layer0_outputs(3882));
    outputs(458) <= layer0_outputs(265);
    outputs(459) <= not((layer0_outputs(6283)) xor (layer0_outputs(6178)));
    outputs(460) <= layer0_outputs(1905);
    outputs(461) <= (layer0_outputs(4703)) and (layer0_outputs(1573));
    outputs(462) <= layer0_outputs(159);
    outputs(463) <= not(layer0_outputs(7515));
    outputs(464) <= layer0_outputs(5658);
    outputs(465) <= not(layer0_outputs(1221));
    outputs(466) <= not((layer0_outputs(3269)) xor (layer0_outputs(3287)));
    outputs(467) <= not(layer0_outputs(2356));
    outputs(468) <= (layer0_outputs(7094)) or (layer0_outputs(4434));
    outputs(469) <= not(layer0_outputs(1590)) or (layer0_outputs(3334));
    outputs(470) <= (layer0_outputs(4223)) and (layer0_outputs(6884));
    outputs(471) <= (layer0_outputs(885)) or (layer0_outputs(3945));
    outputs(472) <= (layer0_outputs(567)) or (layer0_outputs(6692));
    outputs(473) <= not((layer0_outputs(6697)) and (layer0_outputs(1515)));
    outputs(474) <= (layer0_outputs(7107)) and not (layer0_outputs(5399));
    outputs(475) <= (layer0_outputs(5822)) and not (layer0_outputs(6205));
    outputs(476) <= not(layer0_outputs(2165));
    outputs(477) <= not((layer0_outputs(2217)) and (layer0_outputs(590)));
    outputs(478) <= (layer0_outputs(3745)) or (layer0_outputs(186));
    outputs(479) <= (layer0_outputs(3575)) and (layer0_outputs(2776));
    outputs(480) <= layer0_outputs(4439);
    outputs(481) <= not((layer0_outputs(1727)) and (layer0_outputs(768)));
    outputs(482) <= layer0_outputs(2116);
    outputs(483) <= not(layer0_outputs(4401));
    outputs(484) <= (layer0_outputs(3853)) and not (layer0_outputs(1479));
    outputs(485) <= (layer0_outputs(907)) and not (layer0_outputs(3760));
    outputs(486) <= (layer0_outputs(7274)) and (layer0_outputs(764));
    outputs(487) <= (layer0_outputs(4608)) and not (layer0_outputs(6771));
    outputs(488) <= (layer0_outputs(3267)) xor (layer0_outputs(1349));
    outputs(489) <= not(layer0_outputs(5531));
    outputs(490) <= layer0_outputs(1247);
    outputs(491) <= layer0_outputs(2390);
    outputs(492) <= (layer0_outputs(1483)) and (layer0_outputs(1759));
    outputs(493) <= layer0_outputs(1603);
    outputs(494) <= (layer0_outputs(5985)) and not (layer0_outputs(4088));
    outputs(495) <= layer0_outputs(6348);
    outputs(496) <= not((layer0_outputs(5244)) or (layer0_outputs(4024)));
    outputs(497) <= not((layer0_outputs(6008)) xor (layer0_outputs(969)));
    outputs(498) <= layer0_outputs(4656);
    outputs(499) <= (layer0_outputs(4294)) and not (layer0_outputs(4059));
    outputs(500) <= not(layer0_outputs(2696));
    outputs(501) <= layer0_outputs(5893);
    outputs(502) <= not(layer0_outputs(3927));
    outputs(503) <= not((layer0_outputs(978)) xor (layer0_outputs(668)));
    outputs(504) <= layer0_outputs(7597);
    outputs(505) <= (layer0_outputs(7453)) and not (layer0_outputs(4653));
    outputs(506) <= not(layer0_outputs(1513));
    outputs(507) <= not(layer0_outputs(5781));
    outputs(508) <= (layer0_outputs(5190)) xor (layer0_outputs(5687));
    outputs(509) <= not((layer0_outputs(6920)) xor (layer0_outputs(1214)));
    outputs(510) <= not((layer0_outputs(216)) xor (layer0_outputs(2202)));
    outputs(511) <= layer0_outputs(2863);
    outputs(512) <= not((layer0_outputs(5766)) and (layer0_outputs(3880)));
    outputs(513) <= (layer0_outputs(6013)) xor (layer0_outputs(3633));
    outputs(514) <= (layer0_outputs(3016)) xor (layer0_outputs(4860));
    outputs(515) <= layer0_outputs(7066);
    outputs(516) <= not((layer0_outputs(3790)) or (layer0_outputs(6961)));
    outputs(517) <= layer0_outputs(522);
    outputs(518) <= not(layer0_outputs(1585));
    outputs(519) <= not(layer0_outputs(1217));
    outputs(520) <= layer0_outputs(1668);
    outputs(521) <= (layer0_outputs(6132)) and (layer0_outputs(1216));
    outputs(522) <= not(layer0_outputs(7364)) or (layer0_outputs(1233));
    outputs(523) <= layer0_outputs(7055);
    outputs(524) <= (layer0_outputs(3336)) xor (layer0_outputs(4793));
    outputs(525) <= (layer0_outputs(4284)) xor (layer0_outputs(3951));
    outputs(526) <= layer0_outputs(5522);
    outputs(527) <= layer0_outputs(94);
    outputs(528) <= (layer0_outputs(4687)) and not (layer0_outputs(5642));
    outputs(529) <= (layer0_outputs(5585)) or (layer0_outputs(5274));
    outputs(530) <= (layer0_outputs(4450)) and not (layer0_outputs(358));
    outputs(531) <= not(layer0_outputs(5033)) or (layer0_outputs(6578));
    outputs(532) <= not(layer0_outputs(3561)) or (layer0_outputs(5555));
    outputs(533) <= not(layer0_outputs(5262));
    outputs(534) <= (layer0_outputs(949)) and not (layer0_outputs(5431));
    outputs(535) <= not(layer0_outputs(1822));
    outputs(536) <= (layer0_outputs(2226)) xor (layer0_outputs(6277));
    outputs(537) <= (layer0_outputs(1834)) or (layer0_outputs(5658));
    outputs(538) <= not((layer0_outputs(6970)) xor (layer0_outputs(359)));
    outputs(539) <= not((layer0_outputs(4543)) and (layer0_outputs(5882)));
    outputs(540) <= layer0_outputs(1713);
    outputs(541) <= not(layer0_outputs(6885));
    outputs(542) <= layer0_outputs(6934);
    outputs(543) <= not(layer0_outputs(6071));
    outputs(544) <= not((layer0_outputs(394)) xor (layer0_outputs(4146)));
    outputs(545) <= (layer0_outputs(1546)) and not (layer0_outputs(6173));
    outputs(546) <= (layer0_outputs(6230)) and (layer0_outputs(3986));
    outputs(547) <= layer0_outputs(2379);
    outputs(548) <= not((layer0_outputs(393)) and (layer0_outputs(7075)));
    outputs(549) <= not(layer0_outputs(2059));
    outputs(550) <= not((layer0_outputs(1457)) or (layer0_outputs(3782)));
    outputs(551) <= not(layer0_outputs(5160)) or (layer0_outputs(7530));
    outputs(552) <= not((layer0_outputs(3040)) and (layer0_outputs(2160)));
    outputs(553) <= not(layer0_outputs(4937));
    outputs(554) <= not(layer0_outputs(1975));
    outputs(555) <= (layer0_outputs(2847)) and (layer0_outputs(6517));
    outputs(556) <= layer0_outputs(4544);
    outputs(557) <= not(layer0_outputs(3558));
    outputs(558) <= (layer0_outputs(5535)) and not (layer0_outputs(44));
    outputs(559) <= not((layer0_outputs(2916)) and (layer0_outputs(4840)));
    outputs(560) <= not((layer0_outputs(6298)) xor (layer0_outputs(2341)));
    outputs(561) <= not(layer0_outputs(1352));
    outputs(562) <= not(layer0_outputs(114));
    outputs(563) <= (layer0_outputs(1844)) xor (layer0_outputs(5705));
    outputs(564) <= (layer0_outputs(1253)) and (layer0_outputs(1004));
    outputs(565) <= layer0_outputs(6956);
    outputs(566) <= (layer0_outputs(2467)) and not (layer0_outputs(609));
    outputs(567) <= not(layer0_outputs(3138)) or (layer0_outputs(3048));
    outputs(568) <= layer0_outputs(6220);
    outputs(569) <= (layer0_outputs(7344)) and not (layer0_outputs(4565));
    outputs(570) <= not((layer0_outputs(6774)) xor (layer0_outputs(5673)));
    outputs(571) <= (layer0_outputs(2854)) or (layer0_outputs(627));
    outputs(572) <= not((layer0_outputs(6588)) xor (layer0_outputs(6198)));
    outputs(573) <= not((layer0_outputs(5815)) and (layer0_outputs(3588)));
    outputs(574) <= (layer0_outputs(1554)) xor (layer0_outputs(3484));
    outputs(575) <= not((layer0_outputs(4971)) xor (layer0_outputs(2989)));
    outputs(576) <= (layer0_outputs(3194)) xor (layer0_outputs(7642));
    outputs(577) <= not(layer0_outputs(318)) or (layer0_outputs(4418));
    outputs(578) <= layer0_outputs(5914);
    outputs(579) <= (layer0_outputs(2623)) and not (layer0_outputs(3163));
    outputs(580) <= not(layer0_outputs(288));
    outputs(581) <= layer0_outputs(6966);
    outputs(582) <= (layer0_outputs(3975)) and not (layer0_outputs(6971));
    outputs(583) <= not((layer0_outputs(4693)) or (layer0_outputs(4475)));
    outputs(584) <= layer0_outputs(3462);
    outputs(585) <= not(layer0_outputs(7255));
    outputs(586) <= layer0_outputs(3627);
    outputs(587) <= layer0_outputs(867);
    outputs(588) <= (layer0_outputs(7296)) and not (layer0_outputs(5599));
    outputs(589) <= (layer0_outputs(1862)) and not (layer0_outputs(7052));
    outputs(590) <= not((layer0_outputs(5839)) and (layer0_outputs(5589)));
    outputs(591) <= not(layer0_outputs(992));
    outputs(592) <= layer0_outputs(1809);
    outputs(593) <= not((layer0_outputs(2679)) and (layer0_outputs(4142)));
    outputs(594) <= not(layer0_outputs(831));
    outputs(595) <= not(layer0_outputs(6193));
    outputs(596) <= not(layer0_outputs(134));
    outputs(597) <= not((layer0_outputs(1679)) and (layer0_outputs(3749)));
    outputs(598) <= not(layer0_outputs(5087));
    outputs(599) <= layer0_outputs(4183);
    outputs(600) <= (layer0_outputs(6923)) and (layer0_outputs(556));
    outputs(601) <= (layer0_outputs(6437)) and not (layer0_outputs(7132));
    outputs(602) <= not(layer0_outputs(7442));
    outputs(603) <= layer0_outputs(6677);
    outputs(604) <= not((layer0_outputs(774)) xor (layer0_outputs(1582)));
    outputs(605) <= (layer0_outputs(5579)) and not (layer0_outputs(6857));
    outputs(606) <= layer0_outputs(3270);
    outputs(607) <= (layer0_outputs(4037)) xor (layer0_outputs(6359));
    outputs(608) <= not((layer0_outputs(759)) and (layer0_outputs(7623)));
    outputs(609) <= not(layer0_outputs(7112));
    outputs(610) <= not(layer0_outputs(2381));
    outputs(611) <= not(layer0_outputs(7185)) or (layer0_outputs(1115));
    outputs(612) <= not(layer0_outputs(7645)) or (layer0_outputs(7196));
    outputs(613) <= not((layer0_outputs(3307)) xor (layer0_outputs(6530)));
    outputs(614) <= (layer0_outputs(4236)) and not (layer0_outputs(7528));
    outputs(615) <= not(layer0_outputs(2388));
    outputs(616) <= not(layer0_outputs(6697));
    outputs(617) <= (layer0_outputs(5346)) and not (layer0_outputs(5865));
    outputs(618) <= not(layer0_outputs(2598));
    outputs(619) <= layer0_outputs(7406);
    outputs(620) <= not(layer0_outputs(906));
    outputs(621) <= not(layer0_outputs(3786));
    outputs(622) <= (layer0_outputs(1235)) xor (layer0_outputs(1686));
    outputs(623) <= not((layer0_outputs(63)) and (layer0_outputs(5310)));
    outputs(624) <= layer0_outputs(4299);
    outputs(625) <= not((layer0_outputs(986)) or (layer0_outputs(7046)));
    outputs(626) <= not(layer0_outputs(3898));
    outputs(627) <= layer0_outputs(3975);
    outputs(628) <= layer0_outputs(1432);
    outputs(629) <= not(layer0_outputs(1542)) or (layer0_outputs(5344));
    outputs(630) <= layer0_outputs(1243);
    outputs(631) <= layer0_outputs(3310);
    outputs(632) <= not(layer0_outputs(1446));
    outputs(633) <= not(layer0_outputs(4969));
    outputs(634) <= not((layer0_outputs(4825)) and (layer0_outputs(7541)));
    outputs(635) <= not((layer0_outputs(2673)) xor (layer0_outputs(5462)));
    outputs(636) <= not(layer0_outputs(4601));
    outputs(637) <= (layer0_outputs(6309)) and (layer0_outputs(5696));
    outputs(638) <= not(layer0_outputs(4228));
    outputs(639) <= (layer0_outputs(7170)) and not (layer0_outputs(3226));
    outputs(640) <= not(layer0_outputs(4323));
    outputs(641) <= layer0_outputs(1075);
    outputs(642) <= not(layer0_outputs(1480));
    outputs(643) <= not((layer0_outputs(5117)) xor (layer0_outputs(4036)));
    outputs(644) <= not(layer0_outputs(1307));
    outputs(645) <= layer0_outputs(6807);
    outputs(646) <= not(layer0_outputs(2677)) or (layer0_outputs(3168));
    outputs(647) <= not((layer0_outputs(6390)) and (layer0_outputs(4969)));
    outputs(648) <= layer0_outputs(4986);
    outputs(649) <= layer0_outputs(4811);
    outputs(650) <= (layer0_outputs(5316)) and not (layer0_outputs(3291));
    outputs(651) <= not(layer0_outputs(470)) or (layer0_outputs(1495));
    outputs(652) <= not(layer0_outputs(3836));
    outputs(653) <= not((layer0_outputs(3538)) and (layer0_outputs(1876)));
    outputs(654) <= not(layer0_outputs(1819));
    outputs(655) <= (layer0_outputs(7672)) and not (layer0_outputs(850));
    outputs(656) <= layer0_outputs(4890);
    outputs(657) <= not(layer0_outputs(3055)) or (layer0_outputs(596));
    outputs(658) <= layer0_outputs(5722);
    outputs(659) <= layer0_outputs(7223);
    outputs(660) <= not(layer0_outputs(1863));
    outputs(661) <= not(layer0_outputs(373)) or (layer0_outputs(772));
    outputs(662) <= not((layer0_outputs(6631)) xor (layer0_outputs(5081)));
    outputs(663) <= not(layer0_outputs(3257));
    outputs(664) <= layer0_outputs(5689);
    outputs(665) <= not(layer0_outputs(3990));
    outputs(666) <= layer0_outputs(6209);
    outputs(667) <= layer0_outputs(1483);
    outputs(668) <= not(layer0_outputs(953));
    outputs(669) <= (layer0_outputs(6280)) and (layer0_outputs(1237));
    outputs(670) <= not((layer0_outputs(6297)) xor (layer0_outputs(4167)));
    outputs(671) <= (layer0_outputs(1671)) xor (layer0_outputs(5331));
    outputs(672) <= (layer0_outputs(891)) and not (layer0_outputs(1942));
    outputs(673) <= layer0_outputs(3580);
    outputs(674) <= layer0_outputs(242);
    outputs(675) <= (layer0_outputs(2234)) and not (layer0_outputs(3783));
    outputs(676) <= not(layer0_outputs(4288));
    outputs(677) <= not(layer0_outputs(3252));
    outputs(678) <= not(layer0_outputs(1749)) or (layer0_outputs(3009));
    outputs(679) <= not(layer0_outputs(6910));
    outputs(680) <= layer0_outputs(897);
    outputs(681) <= layer0_outputs(5822);
    outputs(682) <= layer0_outputs(251);
    outputs(683) <= (layer0_outputs(2722)) xor (layer0_outputs(2601));
    outputs(684) <= not(layer0_outputs(4456));
    outputs(685) <= (layer0_outputs(5019)) or (layer0_outputs(5973));
    outputs(686) <= not(layer0_outputs(6114));
    outputs(687) <= (layer0_outputs(6682)) and (layer0_outputs(2211));
    outputs(688) <= layer0_outputs(2238);
    outputs(689) <= not(layer0_outputs(5591));
    outputs(690) <= layer0_outputs(3756);
    outputs(691) <= not((layer0_outputs(2345)) and (layer0_outputs(1653)));
    outputs(692) <= layer0_outputs(787);
    outputs(693) <= layer0_outputs(5470);
    outputs(694) <= not(layer0_outputs(3902)) or (layer0_outputs(5376));
    outputs(695) <= (layer0_outputs(1231)) and (layer0_outputs(3644));
    outputs(696) <= not(layer0_outputs(6525)) or (layer0_outputs(2710));
    outputs(697) <= layer0_outputs(791);
    outputs(698) <= not((layer0_outputs(419)) and (layer0_outputs(3869)));
    outputs(699) <= not((layer0_outputs(2343)) or (layer0_outputs(6914)));
    outputs(700) <= not((layer0_outputs(2951)) or (layer0_outputs(6186)));
    outputs(701) <= not(layer0_outputs(6708));
    outputs(702) <= not(layer0_outputs(4211));
    outputs(703) <= (layer0_outputs(4095)) xor (layer0_outputs(1835));
    outputs(704) <= (layer0_outputs(3937)) or (layer0_outputs(5240));
    outputs(705) <= not(layer0_outputs(7210)) or (layer0_outputs(6089));
    outputs(706) <= layer0_outputs(695);
    outputs(707) <= not(layer0_outputs(2409));
    outputs(708) <= not(layer0_outputs(1846));
    outputs(709) <= layer0_outputs(6410);
    outputs(710) <= not((layer0_outputs(6524)) xor (layer0_outputs(238)));
    outputs(711) <= (layer0_outputs(2082)) and not (layer0_outputs(5191));
    outputs(712) <= (layer0_outputs(4690)) xor (layer0_outputs(5136));
    outputs(713) <= (layer0_outputs(853)) and not (layer0_outputs(636));
    outputs(714) <= (layer0_outputs(2596)) and (layer0_outputs(4440));
    outputs(715) <= not(layer0_outputs(4124)) or (layer0_outputs(4460));
    outputs(716) <= not(layer0_outputs(1811));
    outputs(717) <= not((layer0_outputs(5258)) and (layer0_outputs(878)));
    outputs(718) <= not(layer0_outputs(3895)) or (layer0_outputs(2827));
    outputs(719) <= not(layer0_outputs(794));
    outputs(720) <= layer0_outputs(161);
    outputs(721) <= not(layer0_outputs(6695)) or (layer0_outputs(3046));
    outputs(722) <= not((layer0_outputs(3783)) or (layer0_outputs(7071)));
    outputs(723) <= (layer0_outputs(7393)) and not (layer0_outputs(2176));
    outputs(724) <= layer0_outputs(4507);
    outputs(725) <= (layer0_outputs(6306)) and (layer0_outputs(1006));
    outputs(726) <= not(layer0_outputs(2505));
    outputs(727) <= not(layer0_outputs(5273));
    outputs(728) <= layer0_outputs(6100);
    outputs(729) <= not((layer0_outputs(2331)) xor (layer0_outputs(692)));
    outputs(730) <= (layer0_outputs(590)) xor (layer0_outputs(2008));
    outputs(731) <= not(layer0_outputs(7180));
    outputs(732) <= (layer0_outputs(5315)) xor (layer0_outputs(1883));
    outputs(733) <= not((layer0_outputs(2791)) xor (layer0_outputs(727)));
    outputs(734) <= not(layer0_outputs(3163));
    outputs(735) <= (layer0_outputs(5432)) or (layer0_outputs(5946));
    outputs(736) <= layer0_outputs(5878);
    outputs(737) <= not(layer0_outputs(7390)) or (layer0_outputs(5337));
    outputs(738) <= (layer0_outputs(3314)) and not (layer0_outputs(7388));
    outputs(739) <= (layer0_outputs(3522)) or (layer0_outputs(5240));
    outputs(740) <= layer0_outputs(3627);
    outputs(741) <= not(layer0_outputs(1538)) or (layer0_outputs(1334));
    outputs(742) <= (layer0_outputs(4661)) and (layer0_outputs(5373));
    outputs(743) <= (layer0_outputs(2242)) and not (layer0_outputs(6707));
    outputs(744) <= not(layer0_outputs(4716));
    outputs(745) <= layer0_outputs(4917);
    outputs(746) <= layer0_outputs(5524);
    outputs(747) <= (layer0_outputs(586)) xor (layer0_outputs(1531));
    outputs(748) <= not(layer0_outputs(4205));
    outputs(749) <= (layer0_outputs(1341)) and not (layer0_outputs(7111));
    outputs(750) <= (layer0_outputs(501)) and not (layer0_outputs(6099));
    outputs(751) <= not(layer0_outputs(5854));
    outputs(752) <= not(layer0_outputs(4990)) or (layer0_outputs(7461));
    outputs(753) <= layer0_outputs(3436);
    outputs(754) <= layer0_outputs(357);
    outputs(755) <= (layer0_outputs(6312)) and not (layer0_outputs(402));
    outputs(756) <= (layer0_outputs(5168)) or (layer0_outputs(3115));
    outputs(757) <= not((layer0_outputs(6521)) and (layer0_outputs(477)));
    outputs(758) <= not((layer0_outputs(3350)) xor (layer0_outputs(1010)));
    outputs(759) <= layer0_outputs(1021);
    outputs(760) <= not(layer0_outputs(3093)) or (layer0_outputs(5075));
    outputs(761) <= not(layer0_outputs(1074));
    outputs(762) <= not((layer0_outputs(2446)) xor (layer0_outputs(6422)));
    outputs(763) <= not(layer0_outputs(883));
    outputs(764) <= (layer0_outputs(4576)) xor (layer0_outputs(6983));
    outputs(765) <= (layer0_outputs(7429)) and not (layer0_outputs(5918));
    outputs(766) <= (layer0_outputs(5653)) and not (layer0_outputs(4572));
    outputs(767) <= (layer0_outputs(3235)) and (layer0_outputs(2068));
    outputs(768) <= not((layer0_outputs(7615)) xor (layer0_outputs(6525)));
    outputs(769) <= (layer0_outputs(2133)) xor (layer0_outputs(6476));
    outputs(770) <= layer0_outputs(6929);
    outputs(771) <= not((layer0_outputs(512)) or (layer0_outputs(2694)));
    outputs(772) <= not((layer0_outputs(4518)) or (layer0_outputs(2953)));
    outputs(773) <= not((layer0_outputs(7629)) xor (layer0_outputs(4180)));
    outputs(774) <= not((layer0_outputs(3003)) xor (layer0_outputs(1264)));
    outputs(775) <= not(layer0_outputs(3461)) or (layer0_outputs(3839));
    outputs(776) <= not((layer0_outputs(4984)) xor (layer0_outputs(328)));
    outputs(777) <= (layer0_outputs(6509)) xor (layer0_outputs(6471));
    outputs(778) <= (layer0_outputs(689)) and not (layer0_outputs(3012));
    outputs(779) <= (layer0_outputs(4738)) and not (layer0_outputs(6636));
    outputs(780) <= (layer0_outputs(4067)) and not (layer0_outputs(4257));
    outputs(781) <= (layer0_outputs(2007)) and (layer0_outputs(6888));
    outputs(782) <= not((layer0_outputs(2238)) xor (layer0_outputs(2880)));
    outputs(783) <= (layer0_outputs(1920)) and not (layer0_outputs(3479));
    outputs(784) <= (layer0_outputs(390)) and not (layer0_outputs(2218));
    outputs(785) <= not(layer0_outputs(5552));
    outputs(786) <= not(layer0_outputs(6872));
    outputs(787) <= not((layer0_outputs(4819)) or (layer0_outputs(5669)));
    outputs(788) <= (layer0_outputs(1403)) and (layer0_outputs(5131));
    outputs(789) <= not(layer0_outputs(2146));
    outputs(790) <= (layer0_outputs(5528)) and (layer0_outputs(5703));
    outputs(791) <= (layer0_outputs(5028)) and not (layer0_outputs(3571));
    outputs(792) <= (layer0_outputs(4147)) and (layer0_outputs(1845));
    outputs(793) <= (layer0_outputs(7679)) and not (layer0_outputs(2622));
    outputs(794) <= (layer0_outputs(2580)) and not (layer0_outputs(7295));
    outputs(795) <= not((layer0_outputs(3124)) or (layer0_outputs(3201)));
    outputs(796) <= layer0_outputs(6806);
    outputs(797) <= layer0_outputs(4345);
    outputs(798) <= (layer0_outputs(4957)) and not (layer0_outputs(3215));
    outputs(799) <= not(layer0_outputs(3815));
    outputs(800) <= (layer0_outputs(6485)) xor (layer0_outputs(4905));
    outputs(801) <= (layer0_outputs(2046)) and (layer0_outputs(463));
    outputs(802) <= (layer0_outputs(5922)) xor (layer0_outputs(1070));
    outputs(803) <= (layer0_outputs(2538)) and not (layer0_outputs(1689));
    outputs(804) <= layer0_outputs(330);
    outputs(805) <= (layer0_outputs(1045)) and (layer0_outputs(696));
    outputs(806) <= not((layer0_outputs(7474)) or (layer0_outputs(4638)));
    outputs(807) <= not(layer0_outputs(7184));
    outputs(808) <= (layer0_outputs(2537)) and (layer0_outputs(5424));
    outputs(809) <= not((layer0_outputs(5608)) or (layer0_outputs(4071)));
    outputs(810) <= (layer0_outputs(2994)) xor (layer0_outputs(5273));
    outputs(811) <= (layer0_outputs(1993)) and not (layer0_outputs(3037));
    outputs(812) <= (layer0_outputs(4852)) and not (layer0_outputs(3612));
    outputs(813) <= not((layer0_outputs(6075)) or (layer0_outputs(3304)));
    outputs(814) <= not(layer0_outputs(6451));
    outputs(815) <= (layer0_outputs(4356)) and not (layer0_outputs(2281));
    outputs(816) <= (layer0_outputs(4494)) and not (layer0_outputs(2470));
    outputs(817) <= (layer0_outputs(2231)) and not (layer0_outputs(5475));
    outputs(818) <= not((layer0_outputs(4826)) xor (layer0_outputs(6130)));
    outputs(819) <= (layer0_outputs(7237)) and not (layer0_outputs(4432));
    outputs(820) <= (layer0_outputs(2783)) and (layer0_outputs(5644));
    outputs(821) <= (layer0_outputs(4152)) and not (layer0_outputs(3637));
    outputs(822) <= (layer0_outputs(5355)) xor (layer0_outputs(6881));
    outputs(823) <= layer0_outputs(7092);
    outputs(824) <= not(layer0_outputs(538)) or (layer0_outputs(4870));
    outputs(825) <= not((layer0_outputs(871)) or (layer0_outputs(6851)));
    outputs(826) <= not(layer0_outputs(690));
    outputs(827) <= (layer0_outputs(3517)) and not (layer0_outputs(2092));
    outputs(828) <= not((layer0_outputs(1680)) or (layer0_outputs(1284)));
    outputs(829) <= (layer0_outputs(2621)) and not (layer0_outputs(6442));
    outputs(830) <= (layer0_outputs(3430)) and not (layer0_outputs(5601));
    outputs(831) <= (layer0_outputs(108)) and (layer0_outputs(3448));
    outputs(832) <= not((layer0_outputs(6503)) xor (layer0_outputs(784)));
    outputs(833) <= not((layer0_outputs(4516)) xor (layer0_outputs(4857)));
    outputs(834) <= not((layer0_outputs(5888)) xor (layer0_outputs(1329)));
    outputs(835) <= (layer0_outputs(7488)) and (layer0_outputs(2388));
    outputs(836) <= not(layer0_outputs(4281)) or (layer0_outputs(5063));
    outputs(837) <= (layer0_outputs(344)) and not (layer0_outputs(4693));
    outputs(838) <= '0';
    outputs(839) <= (layer0_outputs(5158)) and not (layer0_outputs(3696));
    outputs(840) <= (layer0_outputs(7652)) xor (layer0_outputs(3258));
    outputs(841) <= (layer0_outputs(7116)) and not (layer0_outputs(2041));
    outputs(842) <= (layer0_outputs(3580)) and not (layer0_outputs(4299));
    outputs(843) <= (layer0_outputs(824)) and (layer0_outputs(4287));
    outputs(844) <= (layer0_outputs(5298)) and (layer0_outputs(5134));
    outputs(845) <= not((layer0_outputs(5887)) or (layer0_outputs(4787)));
    outputs(846) <= not(layer0_outputs(6139));
    outputs(847) <= (layer0_outputs(7206)) and not (layer0_outputs(6575));
    outputs(848) <= not(layer0_outputs(4563)) or (layer0_outputs(6248));
    outputs(849) <= (layer0_outputs(5837)) and not (layer0_outputs(4697));
    outputs(850) <= not((layer0_outputs(3)) or (layer0_outputs(5533)));
    outputs(851) <= (layer0_outputs(3795)) and not (layer0_outputs(3259));
    outputs(852) <= not(layer0_outputs(2301));
    outputs(853) <= (layer0_outputs(3955)) and not (layer0_outputs(5751));
    outputs(854) <= not((layer0_outputs(4141)) xor (layer0_outputs(7194)));
    outputs(855) <= (layer0_outputs(3626)) and not (layer0_outputs(4867));
    outputs(856) <= not((layer0_outputs(1919)) xor (layer0_outputs(5296)));
    outputs(857) <= not(layer0_outputs(2652));
    outputs(858) <= not((layer0_outputs(1184)) or (layer0_outputs(3934)));
    outputs(859) <= (layer0_outputs(4082)) and (layer0_outputs(2804));
    outputs(860) <= (layer0_outputs(4014)) and not (layer0_outputs(2919));
    outputs(861) <= (layer0_outputs(1155)) xor (layer0_outputs(6239));
    outputs(862) <= (layer0_outputs(1375)) and not (layer0_outputs(192));
    outputs(863) <= not((layer0_outputs(2099)) or (layer0_outputs(2008)));
    outputs(864) <= not(layer0_outputs(1431));
    outputs(865) <= not((layer0_outputs(1340)) or (layer0_outputs(6495)));
    outputs(866) <= (layer0_outputs(4389)) and not (layer0_outputs(7267));
    outputs(867) <= not((layer0_outputs(4489)) xor (layer0_outputs(2557)));
    outputs(868) <= (layer0_outputs(1325)) xor (layer0_outputs(2206));
    outputs(869) <= (layer0_outputs(953)) and not (layer0_outputs(1177));
    outputs(870) <= layer0_outputs(2872);
    outputs(871) <= (layer0_outputs(1246)) and (layer0_outputs(5424));
    outputs(872) <= not((layer0_outputs(2905)) or (layer0_outputs(922)));
    outputs(873) <= not((layer0_outputs(5275)) xor (layer0_outputs(4638)));
    outputs(874) <= not((layer0_outputs(5991)) xor (layer0_outputs(6898)));
    outputs(875) <= not(layer0_outputs(975));
    outputs(876) <= not(layer0_outputs(1257));
    outputs(877) <= layer0_outputs(6033);
    outputs(878) <= (layer0_outputs(7348)) and not (layer0_outputs(6145));
    outputs(879) <= not((layer0_outputs(2673)) or (layer0_outputs(6736)));
    outputs(880) <= (layer0_outputs(7555)) and not (layer0_outputs(5015));
    outputs(881) <= not(layer0_outputs(3670));
    outputs(882) <= not(layer0_outputs(2601));
    outputs(883) <= (layer0_outputs(6025)) and (layer0_outputs(6080));
    outputs(884) <= not(layer0_outputs(2206)) or (layer0_outputs(34));
    outputs(885) <= (layer0_outputs(3551)) and not (layer0_outputs(7503));
    outputs(886) <= (layer0_outputs(5600)) and not (layer0_outputs(5886));
    outputs(887) <= layer0_outputs(3126);
    outputs(888) <= not((layer0_outputs(5670)) or (layer0_outputs(4261)));
    outputs(889) <= (layer0_outputs(4988)) and not (layer0_outputs(646));
    outputs(890) <= not(layer0_outputs(1909));
    outputs(891) <= not(layer0_outputs(6494));
    outputs(892) <= layer0_outputs(6054);
    outputs(893) <= (layer0_outputs(6147)) and not (layer0_outputs(6305));
    outputs(894) <= (layer0_outputs(3510)) xor (layer0_outputs(6705));
    outputs(895) <= '0';
    outputs(896) <= layer0_outputs(6626);
    outputs(897) <= not(layer0_outputs(6974)) or (layer0_outputs(777));
    outputs(898) <= not((layer0_outputs(1333)) xor (layer0_outputs(814)));
    outputs(899) <= layer0_outputs(3126);
    outputs(900) <= (layer0_outputs(3935)) and (layer0_outputs(7154));
    outputs(901) <= (layer0_outputs(562)) and not (layer0_outputs(4416));
    outputs(902) <= (layer0_outputs(7220)) and not (layer0_outputs(2842));
    outputs(903) <= (layer0_outputs(3406)) and not (layer0_outputs(2065));
    outputs(904) <= (layer0_outputs(4936)) and not (layer0_outputs(2980));
    outputs(905) <= not((layer0_outputs(3740)) or (layer0_outputs(5105)));
    outputs(906) <= not((layer0_outputs(5922)) or (layer0_outputs(5612)));
    outputs(907) <= (layer0_outputs(6338)) and (layer0_outputs(6448));
    outputs(908) <= not((layer0_outputs(2483)) or (layer0_outputs(2193)));
    outputs(909) <= (layer0_outputs(820)) and not (layer0_outputs(6439));
    outputs(910) <= (layer0_outputs(4402)) and not (layer0_outputs(6008));
    outputs(911) <= not(layer0_outputs(185));
    outputs(912) <= (layer0_outputs(1263)) xor (layer0_outputs(3639));
    outputs(913) <= not(layer0_outputs(6220));
    outputs(914) <= (layer0_outputs(266)) xor (layer0_outputs(5465));
    outputs(915) <= (layer0_outputs(3337)) xor (layer0_outputs(1904));
    outputs(916) <= (layer0_outputs(6842)) and not (layer0_outputs(2337));
    outputs(917) <= not((layer0_outputs(1592)) or (layer0_outputs(5652)));
    outputs(918) <= not(layer0_outputs(1559));
    outputs(919) <= (layer0_outputs(964)) and not (layer0_outputs(2184));
    outputs(920) <= (layer0_outputs(3710)) and not (layer0_outputs(977));
    outputs(921) <= not(layer0_outputs(5975));
    outputs(922) <= not((layer0_outputs(3807)) or (layer0_outputs(3162)));
    outputs(923) <= not((layer0_outputs(2532)) or (layer0_outputs(480)));
    outputs(924) <= not((layer0_outputs(5044)) or (layer0_outputs(7217)));
    outputs(925) <= not((layer0_outputs(5522)) or (layer0_outputs(5333)));
    outputs(926) <= (layer0_outputs(6953)) and not (layer0_outputs(3244));
    outputs(927) <= (layer0_outputs(73)) and not (layer0_outputs(4107));
    outputs(928) <= (layer0_outputs(4364)) and not (layer0_outputs(5016));
    outputs(929) <= (layer0_outputs(1560)) and not (layer0_outputs(687));
    outputs(930) <= (layer0_outputs(2004)) and not (layer0_outputs(2762));
    outputs(931) <= not((layer0_outputs(7517)) or (layer0_outputs(5886)));
    outputs(932) <= not((layer0_outputs(2520)) or (layer0_outputs(811)));
    outputs(933) <= (layer0_outputs(7219)) and not (layer0_outputs(4987));
    outputs(934) <= layer0_outputs(358);
    outputs(935) <= not((layer0_outputs(138)) or (layer0_outputs(1611)));
    outputs(936) <= not((layer0_outputs(277)) xor (layer0_outputs(365)));
    outputs(937) <= layer0_outputs(2769);
    outputs(938) <= not(layer0_outputs(6629));
    outputs(939) <= (layer0_outputs(4770)) and not (layer0_outputs(7038));
    outputs(940) <= layer0_outputs(6927);
    outputs(941) <= layer0_outputs(6276);
    outputs(942) <= not((layer0_outputs(6031)) xor (layer0_outputs(1368)));
    outputs(943) <= not((layer0_outputs(3805)) or (layer0_outputs(7173)));
    outputs(944) <= (layer0_outputs(1810)) and not (layer0_outputs(5151));
    outputs(945) <= not(layer0_outputs(6381));
    outputs(946) <= not(layer0_outputs(3205));
    outputs(947) <= not(layer0_outputs(4312)) or (layer0_outputs(399));
    outputs(948) <= not((layer0_outputs(6799)) or (layer0_outputs(1248)));
    outputs(949) <= '0';
    outputs(950) <= not((layer0_outputs(1954)) or (layer0_outputs(6634)));
    outputs(951) <= (layer0_outputs(5419)) and not (layer0_outputs(1948));
    outputs(952) <= not((layer0_outputs(1272)) or (layer0_outputs(3723)));
    outputs(953) <= not((layer0_outputs(4927)) xor (layer0_outputs(7181)));
    outputs(954) <= layer0_outputs(3348);
    outputs(955) <= (layer0_outputs(4455)) and (layer0_outputs(4751));
    outputs(956) <= (layer0_outputs(6776)) and (layer0_outputs(4205));
    outputs(957) <= not(layer0_outputs(2681));
    outputs(958) <= layer0_outputs(218);
    outputs(959) <= not((layer0_outputs(7200)) or (layer0_outputs(665)));
    outputs(960) <= layer0_outputs(2380);
    outputs(961) <= '0';
    outputs(962) <= not((layer0_outputs(4765)) xor (layer0_outputs(1052)));
    outputs(963) <= (layer0_outputs(3459)) and not (layer0_outputs(6170));
    outputs(964) <= (layer0_outputs(5721)) and (layer0_outputs(2138));
    outputs(965) <= layer0_outputs(5639);
    outputs(966) <= not((layer0_outputs(2461)) or (layer0_outputs(457)));
    outputs(967) <= not((layer0_outputs(3024)) or (layer0_outputs(4395)));
    outputs(968) <= not(layer0_outputs(660)) or (layer0_outputs(3771));
    outputs(969) <= not((layer0_outputs(2973)) xor (layer0_outputs(6005)));
    outputs(970) <= not((layer0_outputs(1438)) xor (layer0_outputs(6946)));
    outputs(971) <= (layer0_outputs(2575)) and (layer0_outputs(4997));
    outputs(972) <= (layer0_outputs(3060)) and not (layer0_outputs(3601));
    outputs(973) <= not((layer0_outputs(1344)) xor (layer0_outputs(3305)));
    outputs(974) <= (layer0_outputs(141)) and not (layer0_outputs(7389));
    outputs(975) <= (layer0_outputs(7413)) and not (layer0_outputs(624));
    outputs(976) <= (layer0_outputs(4998)) and not (layer0_outputs(988));
    outputs(977) <= (layer0_outputs(5189)) and not (layer0_outputs(4621));
    outputs(978) <= not((layer0_outputs(6210)) xor (layer0_outputs(6613)));
    outputs(979) <= (layer0_outputs(5077)) xor (layer0_outputs(6060));
    outputs(980) <= not((layer0_outputs(1397)) xor (layer0_outputs(7207)));
    outputs(981) <= not((layer0_outputs(5099)) xor (layer0_outputs(170)));
    outputs(982) <= (layer0_outputs(3071)) and not (layer0_outputs(5123));
    outputs(983) <= (layer0_outputs(7667)) and not (layer0_outputs(2078));
    outputs(984) <= layer0_outputs(2110);
    outputs(985) <= (layer0_outputs(1502)) and not (layer0_outputs(5267));
    outputs(986) <= layer0_outputs(6397);
    outputs(987) <= not(layer0_outputs(4781));
    outputs(988) <= (layer0_outputs(1721)) and (layer0_outputs(688));
    outputs(989) <= not((layer0_outputs(4357)) or (layer0_outputs(5077)));
    outputs(990) <= '0';
    outputs(991) <= (layer0_outputs(374)) and not (layer0_outputs(7045));
    outputs(992) <= not(layer0_outputs(1268));
    outputs(993) <= not((layer0_outputs(6768)) xor (layer0_outputs(2366)));
    outputs(994) <= not((layer0_outputs(7015)) or (layer0_outputs(4978)));
    outputs(995) <= not(layer0_outputs(2382));
    outputs(996) <= (layer0_outputs(3039)) and not (layer0_outputs(2657));
    outputs(997) <= (layer0_outputs(1463)) and not (layer0_outputs(6411));
    outputs(998) <= not((layer0_outputs(2126)) xor (layer0_outputs(5951)));
    outputs(999) <= not((layer0_outputs(4073)) xor (layer0_outputs(1304)));
    outputs(1000) <= (layer0_outputs(3279)) and (layer0_outputs(7213));
    outputs(1001) <= not((layer0_outputs(5338)) xor (layer0_outputs(1608)));
    outputs(1002) <= (layer0_outputs(5738)) and not (layer0_outputs(3022));
    outputs(1003) <= layer0_outputs(7589);
    outputs(1004) <= (layer0_outputs(2882)) and not (layer0_outputs(3998));
    outputs(1005) <= (layer0_outputs(616)) and not (layer0_outputs(3615));
    outputs(1006) <= not(layer0_outputs(1037));
    outputs(1007) <= (layer0_outputs(4732)) and (layer0_outputs(447));
    outputs(1008) <= (layer0_outputs(7367)) and not (layer0_outputs(3292));
    outputs(1009) <= not((layer0_outputs(6203)) xor (layer0_outputs(4269)));
    outputs(1010) <= not((layer0_outputs(7098)) or (layer0_outputs(2236)));
    outputs(1011) <= (layer0_outputs(1106)) xor (layer0_outputs(4684));
    outputs(1012) <= (layer0_outputs(6299)) and (layer0_outputs(1701));
    outputs(1013) <= layer0_outputs(5577);
    outputs(1014) <= (layer0_outputs(5076)) and not (layer0_outputs(2373));
    outputs(1015) <= (layer0_outputs(829)) xor (layer0_outputs(6544));
    outputs(1016) <= (layer0_outputs(1326)) and not (layer0_outputs(3316));
    outputs(1017) <= '0';
    outputs(1018) <= (layer0_outputs(7109)) and not (layer0_outputs(4521));
    outputs(1019) <= not((layer0_outputs(6662)) or (layer0_outputs(2625)));
    outputs(1020) <= (layer0_outputs(6192)) and not (layer0_outputs(3131));
    outputs(1021) <= (layer0_outputs(7133)) and not (layer0_outputs(4801));
    outputs(1022) <= (layer0_outputs(4206)) and (layer0_outputs(1058));
    outputs(1023) <= (layer0_outputs(6215)) and (layer0_outputs(5564));
    outputs(1024) <= (layer0_outputs(2826)) and not (layer0_outputs(2551));
    outputs(1025) <= not((layer0_outputs(6781)) or (layer0_outputs(2812)));
    outputs(1026) <= (layer0_outputs(854)) and not (layer0_outputs(3473));
    outputs(1027) <= (layer0_outputs(5344)) and not (layer0_outputs(4126));
    outputs(1028) <= (layer0_outputs(6223)) and (layer0_outputs(6017));
    outputs(1029) <= not(layer0_outputs(3284));
    outputs(1030) <= not((layer0_outputs(3330)) xor (layer0_outputs(2307)));
    outputs(1031) <= (layer0_outputs(340)) and not (layer0_outputs(826));
    outputs(1032) <= layer0_outputs(5334);
    outputs(1033) <= (layer0_outputs(7277)) xor (layer0_outputs(5911));
    outputs(1034) <= (layer0_outputs(3393)) and not (layer0_outputs(6370));
    outputs(1035) <= (layer0_outputs(1913)) xor (layer0_outputs(5832));
    outputs(1036) <= (layer0_outputs(7097)) and (layer0_outputs(3232));
    outputs(1037) <= layer0_outputs(140);
    outputs(1038) <= (layer0_outputs(3819)) and (layer0_outputs(6938));
    outputs(1039) <= not((layer0_outputs(7588)) xor (layer0_outputs(4559)));
    outputs(1040) <= (layer0_outputs(7676)) and (layer0_outputs(2780));
    outputs(1041) <= (layer0_outputs(2591)) and not (layer0_outputs(3791));
    outputs(1042) <= not(layer0_outputs(7393));
    outputs(1043) <= not((layer0_outputs(4413)) xor (layer0_outputs(3981)));
    outputs(1044) <= (layer0_outputs(149)) and not (layer0_outputs(486));
    outputs(1045) <= not((layer0_outputs(7188)) or (layer0_outputs(2252)));
    outputs(1046) <= not((layer0_outputs(3885)) xor (layer0_outputs(2879)));
    outputs(1047) <= not((layer0_outputs(4528)) xor (layer0_outputs(5336)));
    outputs(1048) <= not((layer0_outputs(3462)) or (layer0_outputs(3426)));
    outputs(1049) <= not((layer0_outputs(7498)) or (layer0_outputs(7050)));
    outputs(1050) <= (layer0_outputs(2268)) and not (layer0_outputs(85));
    outputs(1051) <= layer0_outputs(889);
    outputs(1052) <= not((layer0_outputs(737)) xor (layer0_outputs(675)));
    outputs(1053) <= (layer0_outputs(25)) and not (layer0_outputs(6355));
    outputs(1054) <= (layer0_outputs(4886)) and not (layer0_outputs(4409));
    outputs(1055) <= not((layer0_outputs(2799)) or (layer0_outputs(2275)));
    outputs(1056) <= not((layer0_outputs(434)) xor (layer0_outputs(7264)));
    outputs(1057) <= (layer0_outputs(91)) and not (layer0_outputs(4209));
    outputs(1058) <= (layer0_outputs(5710)) and (layer0_outputs(3800));
    outputs(1059) <= (layer0_outputs(496)) xor (layer0_outputs(5950));
    outputs(1060) <= (layer0_outputs(6891)) and not (layer0_outputs(1437));
    outputs(1061) <= (layer0_outputs(416)) and (layer0_outputs(1060));
    outputs(1062) <= not((layer0_outputs(972)) or (layer0_outputs(4950)));
    outputs(1063) <= (layer0_outputs(2141)) and not (layer0_outputs(1369));
    outputs(1064) <= not(layer0_outputs(5495));
    outputs(1065) <= (layer0_outputs(1630)) xor (layer0_outputs(2245));
    outputs(1066) <= not((layer0_outputs(4307)) or (layer0_outputs(7031)));
    outputs(1067) <= (layer0_outputs(4305)) and not (layer0_outputs(5561));
    outputs(1068) <= (layer0_outputs(2574)) and not (layer0_outputs(2981));
    outputs(1069) <= not(layer0_outputs(6629));
    outputs(1070) <= not((layer0_outputs(4337)) or (layer0_outputs(5902)));
    outputs(1071) <= (layer0_outputs(24)) and not (layer0_outputs(6803));
    outputs(1072) <= (layer0_outputs(722)) and not (layer0_outputs(5707));
    outputs(1073) <= not((layer0_outputs(4962)) xor (layer0_outputs(1612)));
    outputs(1074) <= not((layer0_outputs(2219)) or (layer0_outputs(7336)));
    outputs(1075) <= (layer0_outputs(2076)) xor (layer0_outputs(4072));
    outputs(1076) <= not((layer0_outputs(3469)) xor (layer0_outputs(1788)));
    outputs(1077) <= not(layer0_outputs(3387)) or (layer0_outputs(1306));
    outputs(1078) <= (layer0_outputs(1321)) and not (layer0_outputs(1841));
    outputs(1079) <= (layer0_outputs(6982)) and not (layer0_outputs(7349));
    outputs(1080) <= not(layer0_outputs(6009));
    outputs(1081) <= (layer0_outputs(3678)) and (layer0_outputs(5262));
    outputs(1082) <= (layer0_outputs(2907)) and (layer0_outputs(81));
    outputs(1083) <= not((layer0_outputs(6314)) xor (layer0_outputs(1202)));
    outputs(1084) <= (layer0_outputs(3139)) and not (layer0_outputs(7177));
    outputs(1085) <= (layer0_outputs(4035)) and (layer0_outputs(1908));
    outputs(1086) <= (layer0_outputs(710)) xor (layer0_outputs(333));
    outputs(1087) <= (layer0_outputs(6909)) and (layer0_outputs(6707));
    outputs(1088) <= (layer0_outputs(4735)) and (layer0_outputs(131));
    outputs(1089) <= layer0_outputs(5708);
    outputs(1090) <= layer0_outputs(3814);
    outputs(1091) <= (layer0_outputs(1533)) and not (layer0_outputs(7496));
    outputs(1092) <= not(layer0_outputs(337));
    outputs(1093) <= layer0_outputs(3408);
    outputs(1094) <= (layer0_outputs(479)) and not (layer0_outputs(1669));
    outputs(1095) <= (layer0_outputs(6097)) and (layer0_outputs(5352));
    outputs(1096) <= not((layer0_outputs(7296)) or (layer0_outputs(3932)));
    outputs(1097) <= (layer0_outputs(4373)) and (layer0_outputs(5704));
    outputs(1098) <= (layer0_outputs(1405)) xor (layer0_outputs(3667));
    outputs(1099) <= (layer0_outputs(6502)) and not (layer0_outputs(295));
    outputs(1100) <= (layer0_outputs(4408)) and (layer0_outputs(6138));
    outputs(1101) <= (layer0_outputs(4852)) and not (layer0_outputs(7627));
    outputs(1102) <= layer0_outputs(1780);
    outputs(1103) <= layer0_outputs(5767);
    outputs(1104) <= (layer0_outputs(6187)) and not (layer0_outputs(5075));
    outputs(1105) <= (layer0_outputs(1966)) and (layer0_outputs(5625));
    outputs(1106) <= (layer0_outputs(898)) and not (layer0_outputs(4474));
    outputs(1107) <= (layer0_outputs(6447)) and not (layer0_outputs(7165));
    outputs(1108) <= (layer0_outputs(7239)) xor (layer0_outputs(2610));
    outputs(1109) <= layer0_outputs(4568);
    outputs(1110) <= not((layer0_outputs(509)) xor (layer0_outputs(5079)));
    outputs(1111) <= not(layer0_outputs(1693));
    outputs(1112) <= not(layer0_outputs(1813));
    outputs(1113) <= (layer0_outputs(1498)) and not (layer0_outputs(7538));
    outputs(1114) <= not((layer0_outputs(7277)) and (layer0_outputs(5428)));
    outputs(1115) <= (layer0_outputs(4101)) and (layer0_outputs(367));
    outputs(1116) <= not((layer0_outputs(3595)) xor (layer0_outputs(664)));
    outputs(1117) <= (layer0_outputs(1840)) and (layer0_outputs(6447));
    outputs(1118) <= (layer0_outputs(5243)) and (layer0_outputs(2003));
    outputs(1119) <= not((layer0_outputs(6907)) xor (layer0_outputs(6590)));
    outputs(1120) <= not((layer0_outputs(6683)) xor (layer0_outputs(2705)));
    outputs(1121) <= (layer0_outputs(4419)) and not (layer0_outputs(6322));
    outputs(1122) <= (layer0_outputs(3989)) xor (layer0_outputs(6004));
    outputs(1123) <= not((layer0_outputs(4249)) or (layer0_outputs(700)));
    outputs(1124) <= (layer0_outputs(2895)) and not (layer0_outputs(1990));
    outputs(1125) <= layer0_outputs(7);
    outputs(1126) <= not((layer0_outputs(7617)) xor (layer0_outputs(6834)));
    outputs(1127) <= (layer0_outputs(6107)) and (layer0_outputs(3384));
    outputs(1128) <= layer0_outputs(7243);
    outputs(1129) <= (layer0_outputs(6216)) and (layer0_outputs(4053));
    outputs(1130) <= (layer0_outputs(4878)) and not (layer0_outputs(5229));
    outputs(1131) <= (layer0_outputs(6316)) and not (layer0_outputs(998));
    outputs(1132) <= not(layer0_outputs(4944));
    outputs(1133) <= not(layer0_outputs(3205));
    outputs(1134) <= not(layer0_outputs(2150));
    outputs(1135) <= (layer0_outputs(3008)) and not (layer0_outputs(5428));
    outputs(1136) <= (layer0_outputs(6214)) xor (layer0_outputs(1663));
    outputs(1137) <= (layer0_outputs(6293)) and not (layer0_outputs(7535));
    outputs(1138) <= layer0_outputs(7311);
    outputs(1139) <= layer0_outputs(1683);
    outputs(1140) <= not((layer0_outputs(5369)) or (layer0_outputs(533)));
    outputs(1141) <= (layer0_outputs(7164)) and not (layer0_outputs(2539));
    outputs(1142) <= (layer0_outputs(4089)) and not (layer0_outputs(1916));
    outputs(1143) <= (layer0_outputs(6861)) and not (layer0_outputs(4439));
    outputs(1144) <= not(layer0_outputs(135)) or (layer0_outputs(6196));
    outputs(1145) <= layer0_outputs(4951);
    outputs(1146) <= (layer0_outputs(4090)) and not (layer0_outputs(6118));
    outputs(1147) <= (layer0_outputs(2447)) and not (layer0_outputs(1116));
    outputs(1148) <= (layer0_outputs(4043)) and not (layer0_outputs(2097));
    outputs(1149) <= not((layer0_outputs(4281)) or (layer0_outputs(80)));
    outputs(1150) <= not((layer0_outputs(2668)) or (layer0_outputs(4834)));
    outputs(1151) <= not((layer0_outputs(3405)) or (layer0_outputs(3304)));
    outputs(1152) <= not((layer0_outputs(3316)) xor (layer0_outputs(7163)));
    outputs(1153) <= (layer0_outputs(6478)) and (layer0_outputs(6611));
    outputs(1154) <= (layer0_outputs(869)) and not (layer0_outputs(5469));
    outputs(1155) <= (layer0_outputs(2190)) and not (layer0_outputs(7368));
    outputs(1156) <= (layer0_outputs(1455)) and not (layer0_outputs(3585));
    outputs(1157) <= not((layer0_outputs(2560)) or (layer0_outputs(2937)));
    outputs(1158) <= (layer0_outputs(2444)) and not (layer0_outputs(3114));
    outputs(1159) <= (layer0_outputs(7347)) xor (layer0_outputs(4119));
    outputs(1160) <= (layer0_outputs(1289)) and not (layer0_outputs(1428));
    outputs(1161) <= not(layer0_outputs(4224));
    outputs(1162) <= (layer0_outputs(2414)) and not (layer0_outputs(5501));
    outputs(1163) <= (layer0_outputs(3068)) and not (layer0_outputs(502));
    outputs(1164) <= not((layer0_outputs(5380)) or (layer0_outputs(1710)));
    outputs(1165) <= not((layer0_outputs(7047)) or (layer0_outputs(4392)));
    outputs(1166) <= (layer0_outputs(4259)) and not (layer0_outputs(139));
    outputs(1167) <= not((layer0_outputs(2168)) or (layer0_outputs(6937)));
    outputs(1168) <= (layer0_outputs(4999)) and not (layer0_outputs(7565));
    outputs(1169) <= (layer0_outputs(6428)) xor (layer0_outputs(7251));
    outputs(1170) <= not((layer0_outputs(7440)) xor (layer0_outputs(3168)));
    outputs(1171) <= (layer0_outputs(2830)) xor (layer0_outputs(6687));
    outputs(1172) <= not((layer0_outputs(3353)) or (layer0_outputs(5569)));
    outputs(1173) <= not((layer0_outputs(2942)) or (layer0_outputs(3896)));
    outputs(1174) <= (layer0_outputs(1524)) and not (layer0_outputs(5620));
    outputs(1175) <= not((layer0_outputs(2890)) xor (layer0_outputs(1193)));
    outputs(1176) <= not((layer0_outputs(5044)) xor (layer0_outputs(3372)));
    outputs(1177) <= not((layer0_outputs(7182)) xor (layer0_outputs(5766)));
    outputs(1178) <= layer0_outputs(3573);
    outputs(1179) <= '0';
    outputs(1180) <= (layer0_outputs(7178)) and (layer0_outputs(4492));
    outputs(1181) <= not(layer0_outputs(5392));
    outputs(1182) <= (layer0_outputs(37)) and not (layer0_outputs(7128));
    outputs(1183) <= (layer0_outputs(552)) and not (layer0_outputs(2692));
    outputs(1184) <= (layer0_outputs(5837)) and not (layer0_outputs(6031));
    outputs(1185) <= layer0_outputs(7623);
    outputs(1186) <= (layer0_outputs(1997)) xor (layer0_outputs(5493));
    outputs(1187) <= (layer0_outputs(5009)) and not (layer0_outputs(3885));
    outputs(1188) <= (layer0_outputs(1452)) xor (layer0_outputs(3074));
    outputs(1189) <= not((layer0_outputs(2031)) xor (layer0_outputs(6114)));
    outputs(1190) <= layer0_outputs(7666);
    outputs(1191) <= (layer0_outputs(899)) and not (layer0_outputs(4270));
    outputs(1192) <= not((layer0_outputs(4411)) xor (layer0_outputs(3887)));
    outputs(1193) <= (layer0_outputs(7385)) and not (layer0_outputs(2480));
    outputs(1194) <= not(layer0_outputs(1771));
    outputs(1195) <= not((layer0_outputs(4726)) or (layer0_outputs(2709)));
    outputs(1196) <= (layer0_outputs(1666)) xor (layer0_outputs(3214));
    outputs(1197) <= (layer0_outputs(128)) xor (layer0_outputs(7033));
    outputs(1198) <= (layer0_outputs(1267)) xor (layer0_outputs(702));
    outputs(1199) <= (layer0_outputs(2888)) and (layer0_outputs(4881));
    outputs(1200) <= not((layer0_outputs(1165)) xor (layer0_outputs(558)));
    outputs(1201) <= (layer0_outputs(13)) and not (layer0_outputs(5908));
    outputs(1202) <= (layer0_outputs(177)) and not (layer0_outputs(5863));
    outputs(1203) <= (layer0_outputs(1722)) and not (layer0_outputs(3632));
    outputs(1204) <= not((layer0_outputs(6045)) or (layer0_outputs(1923)));
    outputs(1205) <= (layer0_outputs(7305)) xor (layer0_outputs(4884));
    outputs(1206) <= (layer0_outputs(3184)) and not (layer0_outputs(5978));
    outputs(1207) <= (layer0_outputs(6981)) and not (layer0_outputs(1104));
    outputs(1208) <= (layer0_outputs(4827)) and (layer0_outputs(1811));
    outputs(1209) <= not((layer0_outputs(2919)) or (layer0_outputs(5914)));
    outputs(1210) <= (layer0_outputs(5345)) and (layer0_outputs(197));
    outputs(1211) <= not((layer0_outputs(2448)) or (layer0_outputs(211)));
    outputs(1212) <= not(layer0_outputs(7245));
    outputs(1213) <= not((layer0_outputs(3929)) or (layer0_outputs(428)));
    outputs(1214) <= not((layer0_outputs(3716)) xor (layer0_outputs(391)));
    outputs(1215) <= (layer0_outputs(1860)) and not (layer0_outputs(6358));
    outputs(1216) <= layer0_outputs(2389);
    outputs(1217) <= layer0_outputs(131);
    outputs(1218) <= not((layer0_outputs(1147)) or (layer0_outputs(7656)));
    outputs(1219) <= (layer0_outputs(5502)) and not (layer0_outputs(5073));
    outputs(1220) <= (layer0_outputs(1696)) and not (layer0_outputs(252));
    outputs(1221) <= not((layer0_outputs(6500)) xor (layer0_outputs(597)));
    outputs(1222) <= (layer0_outputs(234)) xor (layer0_outputs(4320));
    outputs(1223) <= (layer0_outputs(5062)) and (layer0_outputs(836));
    outputs(1224) <= (layer0_outputs(5198)) xor (layer0_outputs(5636));
    outputs(1225) <= layer0_outputs(7589);
    outputs(1226) <= not(layer0_outputs(4747));
    outputs(1227) <= (layer0_outputs(6478)) and not (layer0_outputs(1186));
    outputs(1228) <= not(layer0_outputs(4811));
    outputs(1229) <= not(layer0_outputs(5252));
    outputs(1230) <= (layer0_outputs(6106)) and not (layer0_outputs(2708));
    outputs(1231) <= (layer0_outputs(2825)) and not (layer0_outputs(1126));
    outputs(1232) <= (layer0_outputs(4968)) and not (layer0_outputs(2661));
    outputs(1233) <= (layer0_outputs(2882)) and not (layer0_outputs(4789));
    outputs(1234) <= (layer0_outputs(5020)) xor (layer0_outputs(4488));
    outputs(1235) <= (layer0_outputs(2090)) xor (layer0_outputs(4185));
    outputs(1236) <= not((layer0_outputs(5590)) xor (layer0_outputs(3699)));
    outputs(1237) <= (layer0_outputs(3314)) xor (layer0_outputs(1484));
    outputs(1238) <= (layer0_outputs(6737)) and (layer0_outputs(206));
    outputs(1239) <= (layer0_outputs(1469)) and not (layer0_outputs(1367));
    outputs(1240) <= not((layer0_outputs(2056)) xor (layer0_outputs(1765)));
    outputs(1241) <= layer0_outputs(1511);
    outputs(1242) <= (layer0_outputs(7532)) and not (layer0_outputs(4986));
    outputs(1243) <= (layer0_outputs(6248)) and not (layer0_outputs(6802));
    outputs(1244) <= (layer0_outputs(214)) and (layer0_outputs(4706));
    outputs(1245) <= not((layer0_outputs(414)) or (layer0_outputs(3868)));
    outputs(1246) <= not((layer0_outputs(5691)) or (layer0_outputs(1442)));
    outputs(1247) <= (layer0_outputs(1832)) and not (layer0_outputs(3549));
    outputs(1248) <= (layer0_outputs(3226)) and not (layer0_outputs(7607));
    outputs(1249) <= (layer0_outputs(5872)) and not (layer0_outputs(6821));
    outputs(1250) <= not((layer0_outputs(3550)) xor (layer0_outputs(5573)));
    outputs(1251) <= not((layer0_outputs(5521)) xor (layer0_outputs(7140)));
    outputs(1252) <= layer0_outputs(2868);
    outputs(1253) <= not((layer0_outputs(6531)) or (layer0_outputs(1348)));
    outputs(1254) <= not((layer0_outputs(2438)) or (layer0_outputs(1654)));
    outputs(1255) <= (layer0_outputs(426)) xor (layer0_outputs(6011));
    outputs(1256) <= not((layer0_outputs(4418)) xor (layer0_outputs(5817)));
    outputs(1257) <= (layer0_outputs(306)) and (layer0_outputs(1173));
    outputs(1258) <= not((layer0_outputs(1020)) or (layer0_outputs(7662)));
    outputs(1259) <= (layer0_outputs(6712)) and (layer0_outputs(880));
    outputs(1260) <= not(layer0_outputs(667));
    outputs(1261) <= not((layer0_outputs(4058)) or (layer0_outputs(6706)));
    outputs(1262) <= not((layer0_outputs(5150)) xor (layer0_outputs(645)));
    outputs(1263) <= not((layer0_outputs(7150)) or (layer0_outputs(3069)));
    outputs(1264) <= not(layer0_outputs(2311));
    outputs(1265) <= (layer0_outputs(7534)) and not (layer0_outputs(2313));
    outputs(1266) <= (layer0_outputs(4553)) and not (layer0_outputs(4771));
    outputs(1267) <= not((layer0_outputs(6855)) xor (layer0_outputs(5284)));
    outputs(1268) <= (layer0_outputs(5548)) and not (layer0_outputs(709));
    outputs(1269) <= not((layer0_outputs(3911)) xor (layer0_outputs(1513)));
    outputs(1270) <= (layer0_outputs(6912)) and not (layer0_outputs(3612));
    outputs(1271) <= (layer0_outputs(19)) and not (layer0_outputs(6095));
    outputs(1272) <= '0';
    outputs(1273) <= (layer0_outputs(7234)) and (layer0_outputs(261));
    outputs(1274) <= layer0_outputs(7555);
    outputs(1275) <= not((layer0_outputs(262)) or (layer0_outputs(4092)));
    outputs(1276) <= (layer0_outputs(4097)) and (layer0_outputs(816));
    outputs(1277) <= not((layer0_outputs(6365)) xor (layer0_outputs(2222)));
    outputs(1278) <= (layer0_outputs(6801)) and (layer0_outputs(759));
    outputs(1279) <= layer0_outputs(6835);
    outputs(1280) <= layer0_outputs(3835);
    outputs(1281) <= not((layer0_outputs(144)) xor (layer0_outputs(3944)));
    outputs(1282) <= (layer0_outputs(25)) xor (layer0_outputs(5506));
    outputs(1283) <= (layer0_outputs(286)) and not (layer0_outputs(5418));
    outputs(1284) <= (layer0_outputs(2540)) and not (layer0_outputs(4710));
    outputs(1285) <= not((layer0_outputs(247)) or (layer0_outputs(2412)));
    outputs(1286) <= (layer0_outputs(3930)) and not (layer0_outputs(2193));
    outputs(1287) <= (layer0_outputs(7676)) xor (layer0_outputs(5415));
    outputs(1288) <= not(layer0_outputs(2311));
    outputs(1289) <= (layer0_outputs(399)) and (layer0_outputs(5763));
    outputs(1290) <= not((layer0_outputs(2712)) xor (layer0_outputs(1943)));
    outputs(1291) <= not((layer0_outputs(2252)) or (layer0_outputs(3170)));
    outputs(1292) <= (layer0_outputs(854)) and (layer0_outputs(2102));
    outputs(1293) <= not(layer0_outputs(5446));
    outputs(1294) <= (layer0_outputs(2447)) and (layer0_outputs(2933));
    outputs(1295) <= (layer0_outputs(5089)) and (layer0_outputs(3147));
    outputs(1296) <= (layer0_outputs(6122)) and not (layer0_outputs(6003));
    outputs(1297) <= (layer0_outputs(875)) and not (layer0_outputs(7466));
    outputs(1298) <= not((layer0_outputs(6018)) or (layer0_outputs(6170)));
    outputs(1299) <= (layer0_outputs(33)) and (layer0_outputs(3136));
    outputs(1300) <= not((layer0_outputs(3140)) or (layer0_outputs(6627)));
    outputs(1301) <= (layer0_outputs(4331)) and not (layer0_outputs(845));
    outputs(1302) <= (layer0_outputs(275)) and not (layer0_outputs(5397));
    outputs(1303) <= not((layer0_outputs(1767)) and (layer0_outputs(4614)));
    outputs(1304) <= (layer0_outputs(2944)) xor (layer0_outputs(5232));
    outputs(1305) <= (layer0_outputs(1099)) and not (layer0_outputs(5883));
    outputs(1306) <= not((layer0_outputs(1724)) or (layer0_outputs(1787)));
    outputs(1307) <= layer0_outputs(4722);
    outputs(1308) <= (layer0_outputs(2889)) and (layer0_outputs(4057));
    outputs(1309) <= (layer0_outputs(5048)) and not (layer0_outputs(7454));
    outputs(1310) <= not(layer0_outputs(5231));
    outputs(1311) <= not(layer0_outputs(607));
    outputs(1312) <= (layer0_outputs(591)) xor (layer0_outputs(5355));
    outputs(1313) <= not((layer0_outputs(4930)) xor (layer0_outputs(1869)));
    outputs(1314) <= (layer0_outputs(2199)) and (layer0_outputs(5925));
    outputs(1315) <= (layer0_outputs(4721)) and not (layer0_outputs(7009));
    outputs(1316) <= not(layer0_outputs(6666));
    outputs(1317) <= not((layer0_outputs(1588)) xor (layer0_outputs(6455)));
    outputs(1318) <= (layer0_outputs(5005)) and not (layer0_outputs(689));
    outputs(1319) <= (layer0_outputs(859)) and not (layer0_outputs(1506));
    outputs(1320) <= (layer0_outputs(7179)) xor (layer0_outputs(630));
    outputs(1321) <= (layer0_outputs(3467)) and (layer0_outputs(3502));
    outputs(1322) <= (layer0_outputs(3234)) and not (layer0_outputs(2304));
    outputs(1323) <= (layer0_outputs(3059)) and not (layer0_outputs(3556));
    outputs(1324) <= not((layer0_outputs(1256)) xor (layer0_outputs(2)));
    outputs(1325) <= (layer0_outputs(7216)) and not (layer0_outputs(3376));
    outputs(1326) <= '0';
    outputs(1327) <= (layer0_outputs(4390)) and not (layer0_outputs(5981));
    outputs(1328) <= (layer0_outputs(238)) and not (layer0_outputs(3477));
    outputs(1329) <= layer0_outputs(6082);
    outputs(1330) <= (layer0_outputs(5721)) and not (layer0_outputs(3672));
    outputs(1331) <= (layer0_outputs(3608)) and not (layer0_outputs(1069));
    outputs(1332) <= (layer0_outputs(7378)) and (layer0_outputs(1662));
    outputs(1333) <= (layer0_outputs(6140)) and not (layer0_outputs(647));
    outputs(1334) <= (layer0_outputs(6172)) and (layer0_outputs(2841));
    outputs(1335) <= not((layer0_outputs(3085)) or (layer0_outputs(7483)));
    outputs(1336) <= not((layer0_outputs(2659)) xor (layer0_outputs(7674)));
    outputs(1337) <= layer0_outputs(6497);
    outputs(1338) <= not((layer0_outputs(4748)) or (layer0_outputs(4103)));
    outputs(1339) <= not((layer0_outputs(5821)) xor (layer0_outputs(514)));
    outputs(1340) <= (layer0_outputs(4006)) and (layer0_outputs(5778));
    outputs(1341) <= not((layer0_outputs(1752)) xor (layer0_outputs(4925)));
    outputs(1342) <= (layer0_outputs(5570)) xor (layer0_outputs(740));
    outputs(1343) <= (layer0_outputs(3512)) xor (layer0_outputs(4780));
    outputs(1344) <= (layer0_outputs(3040)) and not (layer0_outputs(3218));
    outputs(1345) <= (layer0_outputs(3914)) xor (layer0_outputs(3204));
    outputs(1346) <= (layer0_outputs(1477)) and not (layer0_outputs(4587));
    outputs(1347) <= not((layer0_outputs(104)) or (layer0_outputs(3096)));
    outputs(1348) <= not((layer0_outputs(5646)) xor (layer0_outputs(2805)));
    outputs(1349) <= not((layer0_outputs(2398)) or (layer0_outputs(671)));
    outputs(1350) <= (layer0_outputs(6854)) and not (layer0_outputs(3812));
    outputs(1351) <= not((layer0_outputs(5949)) xor (layer0_outputs(1951)));
    outputs(1352) <= (layer0_outputs(4277)) or (layer0_outputs(3500));
    outputs(1353) <= not((layer0_outputs(3548)) or (layer0_outputs(5580)));
    outputs(1354) <= not((layer0_outputs(3086)) or (layer0_outputs(3974)));
    outputs(1355) <= not((layer0_outputs(631)) or (layer0_outputs(1804)));
    outputs(1356) <= layer0_outputs(7321);
    outputs(1357) <= (layer0_outputs(7304)) and not (layer0_outputs(2569));
    outputs(1358) <= (layer0_outputs(5928)) xor (layer0_outputs(4265));
    outputs(1359) <= not((layer0_outputs(3169)) or (layer0_outputs(5712)));
    outputs(1360) <= (layer0_outputs(7054)) and (layer0_outputs(5282));
    outputs(1361) <= (layer0_outputs(7197)) and (layer0_outputs(2169));
    outputs(1362) <= (layer0_outputs(4730)) and not (layer0_outputs(2926));
    outputs(1363) <= (layer0_outputs(2855)) and (layer0_outputs(3654));
    outputs(1364) <= (layer0_outputs(637)) xor (layer0_outputs(4253));
    outputs(1365) <= (layer0_outputs(7194)) and (layer0_outputs(6140));
    outputs(1366) <= not((layer0_outputs(7104)) or (layer0_outputs(3110)));
    outputs(1367) <= not((layer0_outputs(6573)) or (layer0_outputs(2448)));
    outputs(1368) <= not(layer0_outputs(3326));
    outputs(1369) <= (layer0_outputs(4150)) and (layer0_outputs(2828));
    outputs(1370) <= not(layer0_outputs(6043));
    outputs(1371) <= not((layer0_outputs(2756)) or (layer0_outputs(1558)));
    outputs(1372) <= not(layer0_outputs(379));
    outputs(1373) <= not(layer0_outputs(3834));
    outputs(1374) <= (layer0_outputs(439)) xor (layer0_outputs(4600));
    outputs(1375) <= not(layer0_outputs(67));
    outputs(1376) <= (layer0_outputs(7124)) xor (layer0_outputs(939));
    outputs(1377) <= not(layer0_outputs(5524));
    outputs(1378) <= (layer0_outputs(5602)) and not (layer0_outputs(3915));
    outputs(1379) <= (layer0_outputs(6137)) and not (layer0_outputs(2027));
    outputs(1380) <= not((layer0_outputs(3159)) or (layer0_outputs(4183)));
    outputs(1381) <= (layer0_outputs(1245)) and not (layer0_outputs(6792));
    outputs(1382) <= (layer0_outputs(1358)) and (layer0_outputs(6911));
    outputs(1383) <= (layer0_outputs(6104)) xor (layer0_outputs(6713));
    outputs(1384) <= (layer0_outputs(910)) and not (layer0_outputs(3034));
    outputs(1385) <= not((layer0_outputs(6541)) or (layer0_outputs(6378)));
    outputs(1386) <= (layer0_outputs(193)) and not (layer0_outputs(5129));
    outputs(1387) <= not(layer0_outputs(5668));
    outputs(1388) <= not((layer0_outputs(196)) or (layer0_outputs(5370)));
    outputs(1389) <= (layer0_outputs(4531)) and not (layer0_outputs(655));
    outputs(1390) <= not(layer0_outputs(2394));
    outputs(1391) <= (layer0_outputs(5342)) xor (layer0_outputs(2057));
    outputs(1392) <= layer0_outputs(769);
    outputs(1393) <= not((layer0_outputs(3685)) xor (layer0_outputs(5840)));
    outputs(1394) <= (layer0_outputs(1156)) and not (layer0_outputs(2204));
    outputs(1395) <= (layer0_outputs(1927)) and (layer0_outputs(1134));
    outputs(1396) <= (layer0_outputs(3041)) and (layer0_outputs(2931));
    outputs(1397) <= (layer0_outputs(5110)) and (layer0_outputs(6354));
    outputs(1398) <= (layer0_outputs(735)) and not (layer0_outputs(4140));
    outputs(1399) <= (layer0_outputs(7564)) and (layer0_outputs(6920));
    outputs(1400) <= (layer0_outputs(89)) xor (layer0_outputs(1382));
    outputs(1401) <= not((layer0_outputs(42)) or (layer0_outputs(1161)));
    outputs(1402) <= (layer0_outputs(53)) and (layer0_outputs(2672));
    outputs(1403) <= layer0_outputs(6263);
    outputs(1404) <= (layer0_outputs(1068)) and not (layer0_outputs(4431));
    outputs(1405) <= not((layer0_outputs(1821)) or (layer0_outputs(4223)));
    outputs(1406) <= (layer0_outputs(1639)) and not (layer0_outputs(4184));
    outputs(1407) <= not((layer0_outputs(7472)) xor (layer0_outputs(390)));
    outputs(1408) <= not((layer0_outputs(7336)) or (layer0_outputs(148)));
    outputs(1409) <= (layer0_outputs(1615)) and not (layer0_outputs(1890));
    outputs(1410) <= (layer0_outputs(2228)) and not (layer0_outputs(280));
    outputs(1411) <= (layer0_outputs(6762)) and not (layer0_outputs(7395));
    outputs(1412) <= (layer0_outputs(1303)) and not (layer0_outputs(3481));
    outputs(1413) <= not(layer0_outputs(6346));
    outputs(1414) <= (layer0_outputs(6812)) xor (layer0_outputs(17));
    outputs(1415) <= not(layer0_outputs(5050));
    outputs(1416) <= (layer0_outputs(1180)) and not (layer0_outputs(7077));
    outputs(1417) <= (layer0_outputs(6111)) and not (layer0_outputs(1261));
    outputs(1418) <= (layer0_outputs(1042)) and not (layer0_outputs(1376));
    outputs(1419) <= (layer0_outputs(6473)) xor (layer0_outputs(4302));
    outputs(1420) <= (layer0_outputs(570)) xor (layer0_outputs(1779));
    outputs(1421) <= (layer0_outputs(6119)) and (layer0_outputs(2675));
    outputs(1422) <= (layer0_outputs(617)) and (layer0_outputs(5538));
    outputs(1423) <= (layer0_outputs(3459)) and not (layer0_outputs(1548));
    outputs(1424) <= (layer0_outputs(4958)) and (layer0_outputs(7679));
    outputs(1425) <= not((layer0_outputs(7371)) xor (layer0_outputs(2600)));
    outputs(1426) <= not((layer0_outputs(2879)) xor (layer0_outputs(776)));
    outputs(1427) <= not((layer0_outputs(2162)) xor (layer0_outputs(4649)));
    outputs(1428) <= layer0_outputs(494);
    outputs(1429) <= not((layer0_outputs(843)) or (layer0_outputs(4030)));
    outputs(1430) <= not(layer0_outputs(3237));
    outputs(1431) <= (layer0_outputs(1005)) and not (layer0_outputs(3389));
    outputs(1432) <= not(layer0_outputs(5552));
    outputs(1433) <= not(layer0_outputs(2384));
    outputs(1434) <= not((layer0_outputs(925)) or (layer0_outputs(1124)));
    outputs(1435) <= (layer0_outputs(5754)) xor (layer0_outputs(6615));
    outputs(1436) <= (layer0_outputs(3018)) and not (layer0_outputs(6042));
    outputs(1437) <= not((layer0_outputs(5956)) or (layer0_outputs(2146)));
    outputs(1438) <= (layer0_outputs(6978)) and not (layer0_outputs(1364));
    outputs(1439) <= (layer0_outputs(5388)) and not (layer0_outputs(427));
    outputs(1440) <= (layer0_outputs(276)) and (layer0_outputs(5933));
    outputs(1441) <= (layer0_outputs(6182)) and not (layer0_outputs(761));
    outputs(1442) <= (layer0_outputs(4712)) and not (layer0_outputs(3634));
    outputs(1443) <= (layer0_outputs(993)) and not (layer0_outputs(2013));
    outputs(1444) <= (layer0_outputs(1959)) and (layer0_outputs(400));
    outputs(1445) <= layer0_outputs(7487);
    outputs(1446) <= (layer0_outputs(6833)) xor (layer0_outputs(2850));
    outputs(1447) <= not((layer0_outputs(4869)) or (layer0_outputs(2546)));
    outputs(1448) <= not((layer0_outputs(2202)) xor (layer0_outputs(3295)));
    outputs(1449) <= not((layer0_outputs(1702)) xor (layer0_outputs(7162)));
    outputs(1450) <= (layer0_outputs(4947)) and not (layer0_outputs(951));
    outputs(1451) <= not(layer0_outputs(3373));
    outputs(1452) <= not((layer0_outputs(5448)) or (layer0_outputs(4052)));
    outputs(1453) <= not((layer0_outputs(3125)) xor (layer0_outputs(7291)));
    outputs(1454) <= (layer0_outputs(2744)) and (layer0_outputs(4391));
    outputs(1455) <= (layer0_outputs(3730)) and (layer0_outputs(4018));
    outputs(1456) <= (layer0_outputs(4859)) and (layer0_outputs(908));
    outputs(1457) <= not(layer0_outputs(1390));
    outputs(1458) <= (layer0_outputs(2247)) and not (layer0_outputs(3700));
    outputs(1459) <= not(layer0_outputs(4892));
    outputs(1460) <= not((layer0_outputs(5315)) xor (layer0_outputs(3200)));
    outputs(1461) <= (layer0_outputs(1013)) and (layer0_outputs(3781));
    outputs(1462) <= not((layer0_outputs(3143)) or (layer0_outputs(1868)));
    outputs(1463) <= (layer0_outputs(6195)) xor (layer0_outputs(7382));
    outputs(1464) <= not((layer0_outputs(6723)) or (layer0_outputs(7331)));
    outputs(1465) <= layer0_outputs(7357);
    outputs(1466) <= (layer0_outputs(5388)) and (layer0_outputs(4783));
    outputs(1467) <= (layer0_outputs(2372)) and (layer0_outputs(2837));
    outputs(1468) <= (layer0_outputs(4227)) and not (layer0_outputs(5695));
    outputs(1469) <= (layer0_outputs(909)) and not (layer0_outputs(5229));
    outputs(1470) <= not((layer0_outputs(3439)) and (layer0_outputs(1095)));
    outputs(1471) <= (layer0_outputs(4981)) and (layer0_outputs(818));
    outputs(1472) <= (layer0_outputs(632)) and not (layer0_outputs(6085));
    outputs(1473) <= (layer0_outputs(253)) and not (layer0_outputs(3016));
    outputs(1474) <= (layer0_outputs(316)) and not (layer0_outputs(5539));
    outputs(1475) <= (layer0_outputs(96)) and not (layer0_outputs(4863));
    outputs(1476) <= not(layer0_outputs(7226));
    outputs(1477) <= (layer0_outputs(3055)) and (layer0_outputs(5354));
    outputs(1478) <= layer0_outputs(1914);
    outputs(1479) <= (layer0_outputs(7046)) and (layer0_outputs(7430));
    outputs(1480) <= not((layer0_outputs(4746)) or (layer0_outputs(5748)));
    outputs(1481) <= not(layer0_outputs(6402));
    outputs(1482) <= not(layer0_outputs(5638));
    outputs(1483) <= (layer0_outputs(1750)) and not (layer0_outputs(4491));
    outputs(1484) <= (layer0_outputs(1180)) and not (layer0_outputs(375));
    outputs(1485) <= (layer0_outputs(6853)) xor (layer0_outputs(672));
    outputs(1486) <= (layer0_outputs(199)) and (layer0_outputs(6710));
    outputs(1487) <= not((layer0_outputs(3144)) xor (layer0_outputs(3236)));
    outputs(1488) <= (layer0_outputs(6012)) and not (layer0_outputs(5145));
    outputs(1489) <= layer0_outputs(5939);
    outputs(1490) <= not((layer0_outputs(6874)) xor (layer0_outputs(7473)));
    outputs(1491) <= layer0_outputs(1871);
    outputs(1492) <= not(layer0_outputs(3970));
    outputs(1493) <= not((layer0_outputs(4052)) or (layer0_outputs(4086)));
    outputs(1494) <= '0';
    outputs(1495) <= layer0_outputs(4532);
    outputs(1496) <= layer0_outputs(23);
    outputs(1497) <= not(layer0_outputs(4917));
    outputs(1498) <= not((layer0_outputs(6623)) or (layer0_outputs(5903)));
    outputs(1499) <= (layer0_outputs(4221)) and not (layer0_outputs(3457));
    outputs(1500) <= not((layer0_outputs(4782)) xor (layer0_outputs(147)));
    outputs(1501) <= not((layer0_outputs(835)) or (layer0_outputs(6565)));
    outputs(1502) <= (layer0_outputs(6782)) and not (layer0_outputs(5645));
    outputs(1503) <= (layer0_outputs(7412)) and not (layer0_outputs(1690));
    outputs(1504) <= not((layer0_outputs(5685)) or (layer0_outputs(4078)));
    outputs(1505) <= not(layer0_outputs(3645));
    outputs(1506) <= (layer0_outputs(368)) and not (layer0_outputs(2303));
    outputs(1507) <= (layer0_outputs(5053)) and (layer0_outputs(7463));
    outputs(1508) <= not(layer0_outputs(185));
    outputs(1509) <= (layer0_outputs(1702)) and not (layer0_outputs(6542));
    outputs(1510) <= not((layer0_outputs(7275)) or (layer0_outputs(7567)));
    outputs(1511) <= not(layer0_outputs(7079));
    outputs(1512) <= not((layer0_outputs(4087)) xor (layer0_outputs(3523)));
    outputs(1513) <= not((layer0_outputs(5456)) or (layer0_outputs(3727)));
    outputs(1514) <= not((layer0_outputs(5876)) or (layer0_outputs(4031)));
    outputs(1515) <= not(layer0_outputs(325));
    outputs(1516) <= (layer0_outputs(52)) and (layer0_outputs(6935));
    outputs(1517) <= (layer0_outputs(4713)) and (layer0_outputs(4252));
    outputs(1518) <= not(layer0_outputs(2203));
    outputs(1519) <= layer0_outputs(7666);
    outputs(1520) <= (layer0_outputs(5502)) and not (layer0_outputs(2815));
    outputs(1521) <= not((layer0_outputs(2721)) xor (layer0_outputs(6968)));
    outputs(1522) <= not((layer0_outputs(3796)) or (layer0_outputs(2254)));
    outputs(1523) <= layer0_outputs(1085);
    outputs(1524) <= (layer0_outputs(579)) and not (layer0_outputs(5136));
    outputs(1525) <= not((layer0_outputs(7609)) or (layer0_outputs(2168)));
    outputs(1526) <= (layer0_outputs(6595)) and (layer0_outputs(2415));
    outputs(1527) <= layer0_outputs(4250);
    outputs(1528) <= not((layer0_outputs(221)) xor (layer0_outputs(3675)));
    outputs(1529) <= (layer0_outputs(2351)) and not (layer0_outputs(5341));
    outputs(1530) <= (layer0_outputs(7347)) and not (layer0_outputs(1882));
    outputs(1531) <= not(layer0_outputs(6631));
    outputs(1532) <= (layer0_outputs(2315)) and (layer0_outputs(3324));
    outputs(1533) <= (layer0_outputs(4462)) and (layer0_outputs(7175));
    outputs(1534) <= (layer0_outputs(5713)) and (layer0_outputs(7455));
    outputs(1535) <= not(layer0_outputs(472));
    outputs(1536) <= not(layer0_outputs(6368));
    outputs(1537) <= not(layer0_outputs(5662));
    outputs(1538) <= not(layer0_outputs(46));
    outputs(1539) <= layer0_outputs(6429);
    outputs(1540) <= (layer0_outputs(5160)) and not (layer0_outputs(154));
    outputs(1541) <= not(layer0_outputs(3851));
    outputs(1542) <= not((layer0_outputs(2425)) and (layer0_outputs(5320)));
    outputs(1543) <= layer0_outputs(7383);
    outputs(1544) <= layer0_outputs(5734);
    outputs(1545) <= not(layer0_outputs(1566));
    outputs(1546) <= not(layer0_outputs(2994));
    outputs(1547) <= (layer0_outputs(155)) or (layer0_outputs(3025));
    outputs(1548) <= not(layer0_outputs(6560));
    outputs(1549) <= not((layer0_outputs(6587)) and (layer0_outputs(2477)));
    outputs(1550) <= (layer0_outputs(2614)) xor (layer0_outputs(533));
    outputs(1551) <= not(layer0_outputs(2986)) or (layer0_outputs(7282));
    outputs(1552) <= (layer0_outputs(5693)) and (layer0_outputs(3065));
    outputs(1553) <= not((layer0_outputs(6569)) xor (layer0_outputs(195)));
    outputs(1554) <= (layer0_outputs(1996)) xor (layer0_outputs(4552));
    outputs(1555) <= (layer0_outputs(2809)) or (layer0_outputs(2194));
    outputs(1556) <= not(layer0_outputs(6477));
    outputs(1557) <= not(layer0_outputs(5177)) or (layer0_outputs(7616));
    outputs(1558) <= layer0_outputs(5975);
    outputs(1559) <= not((layer0_outputs(2534)) xor (layer0_outputs(5139)));
    outputs(1560) <= layer0_outputs(5757);
    outputs(1561) <= (layer0_outputs(2730)) and (layer0_outputs(2246));
    outputs(1562) <= (layer0_outputs(2245)) xor (layer0_outputs(1838));
    outputs(1563) <= not((layer0_outputs(3002)) xor (layer0_outputs(1925)));
    outputs(1564) <= layer0_outputs(7327);
    outputs(1565) <= not(layer0_outputs(5827));
    outputs(1566) <= not((layer0_outputs(471)) xor (layer0_outputs(2772)));
    outputs(1567) <= layer0_outputs(3338);
    outputs(1568) <= not(layer0_outputs(3997));
    outputs(1569) <= not(layer0_outputs(4033)) or (layer0_outputs(4176));
    outputs(1570) <= not((layer0_outputs(4214)) xor (layer0_outputs(5976)));
    outputs(1571) <= (layer0_outputs(1517)) or (layer0_outputs(1116));
    outputs(1572) <= (layer0_outputs(1045)) xor (layer0_outputs(1151));
    outputs(1573) <= layer0_outputs(520);
    outputs(1574) <= layer0_outputs(5039);
    outputs(1575) <= layer0_outputs(4393);
    outputs(1576) <= not(layer0_outputs(3424));
    outputs(1577) <= not(layer0_outputs(5529));
    outputs(1578) <= not((layer0_outputs(3545)) xor (layer0_outputs(7513)));
    outputs(1579) <= (layer0_outputs(2796)) xor (layer0_outputs(3150));
    outputs(1580) <= not((layer0_outputs(2129)) xor (layer0_outputs(4758)));
    outputs(1581) <= (layer0_outputs(210)) xor (layer0_outputs(3686));
    outputs(1582) <= (layer0_outputs(5149)) or (layer0_outputs(423));
    outputs(1583) <= layer0_outputs(6325);
    outputs(1584) <= layer0_outputs(1964);
    outputs(1585) <= layer0_outputs(5876);
    outputs(1586) <= not(layer0_outputs(6127));
    outputs(1587) <= not((layer0_outputs(5713)) and (layer0_outputs(4527)));
    outputs(1588) <= not((layer0_outputs(684)) or (layer0_outputs(3052)));
    outputs(1589) <= not((layer0_outputs(2917)) and (layer0_outputs(5972)));
    outputs(1590) <= layer0_outputs(1947);
    outputs(1591) <= not(layer0_outputs(3104));
    outputs(1592) <= not(layer0_outputs(4233)) or (layer0_outputs(4438));
    outputs(1593) <= not(layer0_outputs(2461));
    outputs(1594) <= not(layer0_outputs(663));
    outputs(1595) <= not(layer0_outputs(7355));
    outputs(1596) <= not(layer0_outputs(5641));
    outputs(1597) <= layer0_outputs(2385);
    outputs(1598) <= (layer0_outputs(6480)) and not (layer0_outputs(208));
    outputs(1599) <= (layer0_outputs(3213)) and not (layer0_outputs(4131));
    outputs(1600) <= (layer0_outputs(6847)) xor (layer0_outputs(3711));
    outputs(1601) <= not((layer0_outputs(1524)) or (layer0_outputs(4385)));
    outputs(1602) <= not(layer0_outputs(5301));
    outputs(1603) <= not(layer0_outputs(6113));
    outputs(1604) <= not(layer0_outputs(561));
    outputs(1605) <= layer0_outputs(3065);
    outputs(1606) <= not(layer0_outputs(3001));
    outputs(1607) <= not((layer0_outputs(1468)) and (layer0_outputs(235)));
    outputs(1608) <= (layer0_outputs(4500)) and not (layer0_outputs(5650));
    outputs(1609) <= not(layer0_outputs(6925));
    outputs(1610) <= not((layer0_outputs(6077)) xor (layer0_outputs(1445)));
    outputs(1611) <= not(layer0_outputs(7410)) or (layer0_outputs(4595));
    outputs(1612) <= (layer0_outputs(225)) and not (layer0_outputs(669));
    outputs(1613) <= (layer0_outputs(6416)) and not (layer0_outputs(2198));
    outputs(1614) <= not(layer0_outputs(7424)) or (layer0_outputs(2561));
    outputs(1615) <= (layer0_outputs(2098)) and not (layer0_outputs(5895));
    outputs(1616) <= layer0_outputs(2170);
    outputs(1617) <= layer0_outputs(6623);
    outputs(1618) <= not((layer0_outputs(307)) and (layer0_outputs(5174)));
    outputs(1619) <= not(layer0_outputs(2220));
    outputs(1620) <= layer0_outputs(7282);
    outputs(1621) <= layer0_outputs(3906);
    outputs(1622) <= not((layer0_outputs(7185)) xor (layer0_outputs(7083)));
    outputs(1623) <= layer0_outputs(4184);
    outputs(1624) <= layer0_outputs(3790);
    outputs(1625) <= not(layer0_outputs(2537));
    outputs(1626) <= not(layer0_outputs(5197)) or (layer0_outputs(1684));
    outputs(1627) <= not((layer0_outputs(698)) xor (layer0_outputs(5439)));
    outputs(1628) <= layer0_outputs(6258);
    outputs(1629) <= layer0_outputs(4465);
    outputs(1630) <= layer0_outputs(1381);
    outputs(1631) <= not((layer0_outputs(3004)) and (layer0_outputs(5758)));
    outputs(1632) <= not(layer0_outputs(4380));
    outputs(1633) <= layer0_outputs(2901);
    outputs(1634) <= layer0_outputs(4289);
    outputs(1635) <= (layer0_outputs(2979)) and not (layer0_outputs(2021));
    outputs(1636) <= (layer0_outputs(2437)) xor (layer0_outputs(5414));
    outputs(1637) <= (layer0_outputs(6067)) or (layer0_outputs(4363));
    outputs(1638) <= layer0_outputs(5015);
    outputs(1639) <= not((layer0_outputs(6859)) and (layer0_outputs(6086)));
    outputs(1640) <= not(layer0_outputs(2817)) or (layer0_outputs(1731));
    outputs(1641) <= layer0_outputs(2687);
    outputs(1642) <= not(layer0_outputs(3950));
    outputs(1643) <= (layer0_outputs(6112)) xor (layer0_outputs(6052));
    outputs(1644) <= not(layer0_outputs(5700));
    outputs(1645) <= layer0_outputs(5348);
    outputs(1646) <= not(layer0_outputs(2866));
    outputs(1647) <= layer0_outputs(5265);
    outputs(1648) <= not(layer0_outputs(2415));
    outputs(1649) <= layer0_outputs(4588);
    outputs(1650) <= not(layer0_outputs(2504));
    outputs(1651) <= not(layer0_outputs(7105)) or (layer0_outputs(3928));
    outputs(1652) <= layer0_outputs(3757);
    outputs(1653) <= (layer0_outputs(4882)) xor (layer0_outputs(5584));
    outputs(1654) <= not(layer0_outputs(1932));
    outputs(1655) <= not((layer0_outputs(2617)) and (layer0_outputs(5912)));
    outputs(1656) <= (layer0_outputs(6456)) xor (layer0_outputs(4717));
    outputs(1657) <= not(layer0_outputs(2967));
    outputs(1658) <= layer0_outputs(2338);
    outputs(1659) <= not((layer0_outputs(6185)) and (layer0_outputs(1071)));
    outputs(1660) <= not((layer0_outputs(4663)) or (layer0_outputs(2937)));
    outputs(1661) <= (layer0_outputs(5781)) and (layer0_outputs(2825));
    outputs(1662) <= layer0_outputs(269);
    outputs(1663) <= layer0_outputs(5808);
    outputs(1664) <= (layer0_outputs(3187)) and not (layer0_outputs(633));
    outputs(1665) <= not(layer0_outputs(7596)) or (layer0_outputs(659));
    outputs(1666) <= not(layer0_outputs(4767));
    outputs(1667) <= not(layer0_outputs(6589)) or (layer0_outputs(2423));
    outputs(1668) <= (layer0_outputs(7544)) and not (layer0_outputs(6290));
    outputs(1669) <= not((layer0_outputs(1853)) and (layer0_outputs(7643)));
    outputs(1670) <= not((layer0_outputs(795)) and (layer0_outputs(4794)));
    outputs(1671) <= not((layer0_outputs(113)) and (layer0_outputs(2134)));
    outputs(1672) <= layer0_outputs(5682);
    outputs(1673) <= not(layer0_outputs(7653)) or (layer0_outputs(206));
    outputs(1674) <= (layer0_outputs(1192)) or (layer0_outputs(6969));
    outputs(1675) <= layer0_outputs(6849);
    outputs(1676) <= (layer0_outputs(4187)) or (layer0_outputs(7496));
    outputs(1677) <= (layer0_outputs(2631)) and not (layer0_outputs(2511));
    outputs(1678) <= layer0_outputs(3621);
    outputs(1679) <= not((layer0_outputs(6523)) xor (layer0_outputs(5989)));
    outputs(1680) <= (layer0_outputs(4291)) or (layer0_outputs(467));
    outputs(1681) <= (layer0_outputs(3531)) xor (layer0_outputs(626));
    outputs(1682) <= not((layer0_outputs(2515)) or (layer0_outputs(1169)));
    outputs(1683) <= (layer0_outputs(3233)) xor (layer0_outputs(3976));
    outputs(1684) <= not((layer0_outputs(3816)) and (layer0_outputs(5119)));
    outputs(1685) <= (layer0_outputs(636)) or (layer0_outputs(2551));
    outputs(1686) <= not(layer0_outputs(6718)) or (layer0_outputs(2674));
    outputs(1687) <= layer0_outputs(5832);
    outputs(1688) <= not(layer0_outputs(3468)) or (layer0_outputs(5490));
    outputs(1689) <= not(layer0_outputs(2771));
    outputs(1690) <= not(layer0_outputs(2611));
    outputs(1691) <= not(layer0_outputs(4932));
    outputs(1692) <= layer0_outputs(1738);
    outputs(1693) <= layer0_outputs(1688);
    outputs(1694) <= layer0_outputs(3739);
    outputs(1695) <= (layer0_outputs(3862)) xor (layer0_outputs(3467));
    outputs(1696) <= not((layer0_outputs(7493)) and (layer0_outputs(4635)));
    outputs(1697) <= layer0_outputs(5804);
    outputs(1698) <= layer0_outputs(6174);
    outputs(1699) <= not((layer0_outputs(5164)) xor (layer0_outputs(2177)));
    outputs(1700) <= (layer0_outputs(7378)) xor (layer0_outputs(1111));
    outputs(1701) <= not(layer0_outputs(2250));
    outputs(1702) <= not(layer0_outputs(1145));
    outputs(1703) <= layer0_outputs(6335);
    outputs(1704) <= (layer0_outputs(3528)) and not (layer0_outputs(6658));
    outputs(1705) <= not((layer0_outputs(143)) xor (layer0_outputs(3216)));
    outputs(1706) <= (layer0_outputs(4592)) and not (layer0_outputs(5275));
    outputs(1707) <= (layer0_outputs(2216)) xor (layer0_outputs(1949));
    outputs(1708) <= not((layer0_outputs(1239)) and (layer0_outputs(4915)));
    outputs(1709) <= not(layer0_outputs(2355));
    outputs(1710) <= not(layer0_outputs(6965));
    outputs(1711) <= (layer0_outputs(2906)) xor (layer0_outputs(1719));
    outputs(1712) <= not((layer0_outputs(2555)) xor (layer0_outputs(1974)));
    outputs(1713) <= not(layer0_outputs(4957)) or (layer0_outputs(1895));
    outputs(1714) <= (layer0_outputs(5191)) xor (layer0_outputs(6098));
    outputs(1715) <= layer0_outputs(6135);
    outputs(1716) <= not(layer0_outputs(2959));
    outputs(1717) <= not((layer0_outputs(5765)) xor (layer0_outputs(3404)));
    outputs(1718) <= layer0_outputs(705);
    outputs(1719) <= (layer0_outputs(2349)) and not (layer0_outputs(1034));
    outputs(1720) <= not(layer0_outputs(4672)) or (layer0_outputs(3427));
    outputs(1721) <= (layer0_outputs(6329)) or (layer0_outputs(840));
    outputs(1722) <= (layer0_outputs(6460)) and not (layer0_outputs(642));
    outputs(1723) <= not(layer0_outputs(5816)) or (layer0_outputs(3601));
    outputs(1724) <= not(layer0_outputs(667));
    outputs(1725) <= (layer0_outputs(2702)) xor (layer0_outputs(3047));
    outputs(1726) <= not(layer0_outputs(620)) or (layer0_outputs(2829));
    outputs(1727) <= (layer0_outputs(6837)) and not (layer0_outputs(3682));
    outputs(1728) <= not(layer0_outputs(3572));
    outputs(1729) <= not((layer0_outputs(6371)) xor (layer0_outputs(5720)));
    outputs(1730) <= not(layer0_outputs(1316));
    outputs(1731) <= layer0_outputs(3398);
    outputs(1732) <= not(layer0_outputs(7635));
    outputs(1733) <= not(layer0_outputs(4204));
    outputs(1734) <= layer0_outputs(4272);
    outputs(1735) <= (layer0_outputs(680)) and (layer0_outputs(1652));
    outputs(1736) <= not(layer0_outputs(4792)) or (layer0_outputs(1306));
    outputs(1737) <= not(layer0_outputs(3867));
    outputs(1738) <= (layer0_outputs(3951)) xor (layer0_outputs(6356));
    outputs(1739) <= not((layer0_outputs(1331)) and (layer0_outputs(1902)));
    outputs(1740) <= not(layer0_outputs(2426));
    outputs(1741) <= not((layer0_outputs(1970)) xor (layer0_outputs(1391)));
    outputs(1742) <= (layer0_outputs(2862)) or (layer0_outputs(6574));
    outputs(1743) <= not((layer0_outputs(6716)) and (layer0_outputs(6995)));
    outputs(1744) <= not((layer0_outputs(4063)) or (layer0_outputs(5450)));
    outputs(1745) <= (layer0_outputs(4192)) xor (layer0_outputs(1735));
    outputs(1746) <= layer0_outputs(4060);
    outputs(1747) <= (layer0_outputs(338)) and not (layer0_outputs(985));
    outputs(1748) <= (layer0_outputs(21)) and not (layer0_outputs(3268));
    outputs(1749) <= (layer0_outputs(1847)) and not (layer0_outputs(936));
    outputs(1750) <= not((layer0_outputs(5537)) xor (layer0_outputs(2153)));
    outputs(1751) <= not(layer0_outputs(1362));
    outputs(1752) <= not(layer0_outputs(1221));
    outputs(1753) <= not((layer0_outputs(3682)) and (layer0_outputs(2620)));
    outputs(1754) <= not(layer0_outputs(4362));
    outputs(1755) <= not(layer0_outputs(1218)) or (layer0_outputs(6093));
    outputs(1756) <= not((layer0_outputs(5374)) and (layer0_outputs(7307)));
    outputs(1757) <= not((layer0_outputs(150)) xor (layer0_outputs(1805)));
    outputs(1758) <= not(layer0_outputs(68));
    outputs(1759) <= not(layer0_outputs(1146));
    outputs(1760) <= not(layer0_outputs(4683));
    outputs(1761) <= (layer0_outputs(4351)) and not (layer0_outputs(4486));
    outputs(1762) <= not(layer0_outputs(7380)) or (layer0_outputs(3334));
    outputs(1763) <= not((layer0_outputs(1496)) xor (layer0_outputs(1451)));
    outputs(1764) <= layer0_outputs(6817);
    outputs(1765) <= layer0_outputs(4389);
    outputs(1766) <= (layer0_outputs(682)) and not (layer0_outputs(6981));
    outputs(1767) <= not(layer0_outputs(585)) or (layer0_outputs(6537));
    outputs(1768) <= layer0_outputs(415);
    outputs(1769) <= layer0_outputs(3787);
    outputs(1770) <= layer0_outputs(942);
    outputs(1771) <= (layer0_outputs(1369)) and not (layer0_outputs(2327));
    outputs(1772) <= not((layer0_outputs(449)) and (layer0_outputs(4797)));
    outputs(1773) <= not(layer0_outputs(3599)) or (layer0_outputs(2386));
    outputs(1774) <= (layer0_outputs(6274)) and (layer0_outputs(202));
    outputs(1775) <= not(layer0_outputs(2526)) or (layer0_outputs(2615));
    outputs(1776) <= (layer0_outputs(6749)) or (layer0_outputs(6955));
    outputs(1777) <= (layer0_outputs(947)) and not (layer0_outputs(736));
    outputs(1778) <= layer0_outputs(1964);
    outputs(1779) <= layer0_outputs(6688);
    outputs(1780) <= not((layer0_outputs(3940)) and (layer0_outputs(55)));
    outputs(1781) <= (layer0_outputs(129)) and (layer0_outputs(7601));
    outputs(1782) <= not(layer0_outputs(892)) or (layer0_outputs(5761));
    outputs(1783) <= (layer0_outputs(6921)) xor (layer0_outputs(888));
    outputs(1784) <= not(layer0_outputs(7021));
    outputs(1785) <= not(layer0_outputs(976));
    outputs(1786) <= not(layer0_outputs(6270));
    outputs(1787) <= not(layer0_outputs(1593)) or (layer0_outputs(6547));
    outputs(1788) <= (layer0_outputs(4985)) or (layer0_outputs(2139));
    outputs(1789) <= not(layer0_outputs(6259));
    outputs(1790) <= layer0_outputs(5460);
    outputs(1791) <= not(layer0_outputs(2255)) or (layer0_outputs(5006));
    outputs(1792) <= layer0_outputs(2183);
    outputs(1793) <= not(layer0_outputs(6344));
    outputs(1794) <= not(layer0_outputs(7519)) or (layer0_outputs(483));
    outputs(1795) <= (layer0_outputs(4197)) or (layer0_outputs(4153));
    outputs(1796) <= (layer0_outputs(4622)) and not (layer0_outputs(6241));
    outputs(1797) <= not(layer0_outputs(2585));
    outputs(1798) <= (layer0_outputs(3758)) or (layer0_outputs(4763));
    outputs(1799) <= (layer0_outputs(226)) or (layer0_outputs(6039));
    outputs(1800) <= (layer0_outputs(5598)) and (layer0_outputs(1367));
    outputs(1801) <= (layer0_outputs(6826)) or (layer0_outputs(1416));
    outputs(1802) <= not((layer0_outputs(3715)) or (layer0_outputs(746)));
    outputs(1803) <= layer0_outputs(1907);
    outputs(1804) <= not(layer0_outputs(4130)) or (layer0_outputs(2116));
    outputs(1805) <= not(layer0_outputs(3315));
    outputs(1806) <= (layer0_outputs(4536)) xor (layer0_outputs(5563));
    outputs(1807) <= not((layer0_outputs(146)) and (layer0_outputs(6878)));
    outputs(1808) <= (layer0_outputs(4228)) and not (layer0_outputs(7038));
    outputs(1809) <= (layer0_outputs(2976)) and (layer0_outputs(5590));
    outputs(1810) <= layer0_outputs(4739);
    outputs(1811) <= not((layer0_outputs(5174)) and (layer0_outputs(7665)));
    outputs(1812) <= not(layer0_outputs(6104)) or (layer0_outputs(3025));
    outputs(1813) <= not((layer0_outputs(7024)) and (layer0_outputs(459)));
    outputs(1814) <= not(layer0_outputs(7034));
    outputs(1815) <= not(layer0_outputs(6832)) or (layer0_outputs(3317));
    outputs(1816) <= not(layer0_outputs(7401));
    outputs(1817) <= layer0_outputs(5242);
    outputs(1818) <= layer0_outputs(2905);
    outputs(1819) <= layer0_outputs(1877);
    outputs(1820) <= layer0_outputs(4575);
    outputs(1821) <= not(layer0_outputs(822)) or (layer0_outputs(739));
    outputs(1822) <= not((layer0_outputs(6933)) xor (layer0_outputs(4897)));
    outputs(1823) <= (layer0_outputs(3088)) and not (layer0_outputs(2449));
    outputs(1824) <= not(layer0_outputs(1195));
    outputs(1825) <= not((layer0_outputs(5427)) and (layer0_outputs(2387)));
    outputs(1826) <= not(layer0_outputs(7641)) or (layer0_outputs(2095));
    outputs(1827) <= layer0_outputs(7402);
    outputs(1828) <= not((layer0_outputs(7643)) xor (layer0_outputs(7503)));
    outputs(1829) <= (layer0_outputs(874)) or (layer0_outputs(5067));
    outputs(1830) <= not(layer0_outputs(1944)) or (layer0_outputs(7630));
    outputs(1831) <= layer0_outputs(6369);
    outputs(1832) <= not((layer0_outputs(7350)) and (layer0_outputs(6700)));
    outputs(1833) <= (layer0_outputs(785)) and (layer0_outputs(3855));
    outputs(1834) <= not(layer0_outputs(3806));
    outputs(1835) <= (layer0_outputs(3506)) and not (layer0_outputs(2278));
    outputs(1836) <= not(layer0_outputs(3315));
    outputs(1837) <= not((layer0_outputs(3803)) xor (layer0_outputs(2188)));
    outputs(1838) <= not(layer0_outputs(2933));
    outputs(1839) <= (layer0_outputs(2187)) and not (layer0_outputs(6513));
    outputs(1840) <= not(layer0_outputs(1503));
    outputs(1841) <= not((layer0_outputs(1044)) and (layer0_outputs(1718)));
    outputs(1842) <= (layer0_outputs(7263)) xor (layer0_outputs(6202));
    outputs(1843) <= layer0_outputs(6747);
    outputs(1844) <= layer0_outputs(7149);
    outputs(1845) <= layer0_outputs(1743);
    outputs(1846) <= not(layer0_outputs(3655));
    outputs(1847) <= not(layer0_outputs(6185)) or (layer0_outputs(6470));
    outputs(1848) <= not((layer0_outputs(5219)) xor (layer0_outputs(2938)));
    outputs(1849) <= not(layer0_outputs(4880));
    outputs(1850) <= (layer0_outputs(2259)) xor (layer0_outputs(7281));
    outputs(1851) <= (layer0_outputs(5543)) and not (layer0_outputs(3256));
    outputs(1852) <= not((layer0_outputs(6146)) xor (layer0_outputs(352)));
    outputs(1853) <= not(layer0_outputs(6783)) or (layer0_outputs(4518));
    outputs(1854) <= (layer0_outputs(30)) and (layer0_outputs(6180));
    outputs(1855) <= not(layer0_outputs(1707));
    outputs(1856) <= layer0_outputs(5976);
    outputs(1857) <= not(layer0_outputs(7081)) or (layer0_outputs(609));
    outputs(1858) <= (layer0_outputs(749)) and not (layer0_outputs(6249));
    outputs(1859) <= not(layer0_outputs(7162));
    outputs(1860) <= not(layer0_outputs(5617));
    outputs(1861) <= layer0_outputs(2361);
    outputs(1862) <= not(layer0_outputs(3594));
    outputs(1863) <= not(layer0_outputs(28)) or (layer0_outputs(5058));
    outputs(1864) <= layer0_outputs(1842);
    outputs(1865) <= not(layer0_outputs(4271));
    outputs(1866) <= not(layer0_outputs(314));
    outputs(1867) <= not((layer0_outputs(5124)) or (layer0_outputs(7028)));
    outputs(1868) <= (layer0_outputs(5635)) and (layer0_outputs(6615));
    outputs(1869) <= not(layer0_outputs(3909));
    outputs(1870) <= layer0_outputs(4006);
    outputs(1871) <= not(layer0_outputs(5657));
    outputs(1872) <= (layer0_outputs(120)) and not (layer0_outputs(370));
    outputs(1873) <= layer0_outputs(842);
    outputs(1874) <= not(layer0_outputs(6084));
    outputs(1875) <= layer0_outputs(2243);
    outputs(1876) <= not((layer0_outputs(4870)) and (layer0_outputs(7362)));
    outputs(1877) <= not(layer0_outputs(5518));
    outputs(1878) <= not(layer0_outputs(214));
    outputs(1879) <= not((layer0_outputs(6673)) xor (layer0_outputs(3773)));
    outputs(1880) <= not((layer0_outputs(2197)) and (layer0_outputs(808)));
    outputs(1881) <= not(layer0_outputs(900));
    outputs(1882) <= not(layer0_outputs(392)) or (layer0_outputs(1061));
    outputs(1883) <= not(layer0_outputs(3180));
    outputs(1884) <= (layer0_outputs(2871)) or (layer0_outputs(7095));
    outputs(1885) <= (layer0_outputs(1188)) or (layer0_outputs(604));
    outputs(1886) <= not(layer0_outputs(2181));
    outputs(1887) <= not(layer0_outputs(7514)) or (layer0_outputs(4564));
    outputs(1888) <= (layer0_outputs(4387)) xor (layer0_outputs(4941));
    outputs(1889) <= (layer0_outputs(2814)) xor (layer0_outputs(840));
    outputs(1890) <= (layer0_outputs(5323)) and not (layer0_outputs(5321));
    outputs(1891) <= not((layer0_outputs(4535)) or (layer0_outputs(6288)));
    outputs(1892) <= (layer0_outputs(4542)) or (layer0_outputs(6643));
    outputs(1893) <= not((layer0_outputs(3779)) or (layer0_outputs(4365)));
    outputs(1894) <= not(layer0_outputs(3513));
    outputs(1895) <= (layer0_outputs(7374)) xor (layer0_outputs(5420));
    outputs(1896) <= not(layer0_outputs(5471));
    outputs(1897) <= layer0_outputs(1012);
    outputs(1898) <= not(layer0_outputs(3502)) or (layer0_outputs(1903));
    outputs(1899) <= (layer0_outputs(4244)) or (layer0_outputs(7654));
    outputs(1900) <= not((layer0_outputs(3620)) xor (layer0_outputs(5025)));
    outputs(1901) <= not(layer0_outputs(3443)) or (layer0_outputs(1872));
    outputs(1902) <= (layer0_outputs(3817)) xor (layer0_outputs(2113));
    outputs(1903) <= (layer0_outputs(6498)) xor (layer0_outputs(3687));
    outputs(1904) <= (layer0_outputs(6919)) and not (layer0_outputs(5163));
    outputs(1905) <= (layer0_outputs(4719)) xor (layer0_outputs(3760));
    outputs(1906) <= layer0_outputs(301);
    outputs(1907) <= not(layer0_outputs(4206));
    outputs(1908) <= (layer0_outputs(4848)) xor (layer0_outputs(7232));
    outputs(1909) <= not((layer0_outputs(763)) or (layer0_outputs(5457)));
    outputs(1910) <= (layer0_outputs(916)) or (layer0_outputs(6091));
    outputs(1911) <= not(layer0_outputs(3008)) or (layer0_outputs(5478));
    outputs(1912) <= (layer0_outputs(4655)) or (layer0_outputs(3677));
    outputs(1913) <= not(layer0_outputs(6845)) or (layer0_outputs(1276));
    outputs(1914) <= not(layer0_outputs(1302));
    outputs(1915) <= layer0_outputs(1394);
    outputs(1916) <= (layer0_outputs(5241)) or (layer0_outputs(1781));
    outputs(1917) <= not(layer0_outputs(5672)) or (layer0_outputs(6764));
    outputs(1918) <= layer0_outputs(5061);
    outputs(1919) <= not(layer0_outputs(1995)) or (layer0_outputs(1366));
    outputs(1920) <= not(layer0_outputs(5644));
    outputs(1921) <= layer0_outputs(7545);
    outputs(1922) <= not((layer0_outputs(1445)) and (layer0_outputs(3059)));
    outputs(1923) <= not((layer0_outputs(4558)) and (layer0_outputs(3057)));
    outputs(1924) <= layer0_outputs(5757);
    outputs(1925) <= layer0_outputs(4329);
    outputs(1926) <= not(layer0_outputs(4448)) or (layer0_outputs(4761));
    outputs(1927) <= not(layer0_outputs(6841)) or (layer0_outputs(6029));
    outputs(1928) <= layer0_outputs(4235);
    outputs(1929) <= layer0_outputs(7655);
    outputs(1930) <= not(layer0_outputs(4144)) or (layer0_outputs(1937));
    outputs(1931) <= (layer0_outputs(2864)) and not (layer0_outputs(4715));
    outputs(1932) <= (layer0_outputs(4034)) or (layer0_outputs(2971));
    outputs(1933) <= layer0_outputs(6154);
    outputs(1934) <= not((layer0_outputs(7292)) and (layer0_outputs(6287)));
    outputs(1935) <= not(layer0_outputs(1128)) or (layer0_outputs(6652));
    outputs(1936) <= not(layer0_outputs(3688));
    outputs(1937) <= (layer0_outputs(1530)) or (layer0_outputs(4743));
    outputs(1938) <= (layer0_outputs(6601)) xor (layer0_outputs(728));
    outputs(1939) <= not(layer0_outputs(5381)) or (layer0_outputs(3089));
    outputs(1940) <= layer0_outputs(1162);
    outputs(1941) <= (layer0_outputs(3532)) xor (layer0_outputs(3335));
    outputs(1942) <= layer0_outputs(2861);
    outputs(1943) <= not((layer0_outputs(1160)) and (layer0_outputs(4768)));
    outputs(1944) <= (layer0_outputs(3971)) and (layer0_outputs(3860));
    outputs(1945) <= not(layer0_outputs(2640));
    outputs(1946) <= (layer0_outputs(784)) or (layer0_outputs(6308));
    outputs(1947) <= not(layer0_outputs(4779));
    outputs(1948) <= (layer0_outputs(4186)) and not (layer0_outputs(7255));
    outputs(1949) <= layer0_outputs(6237);
    outputs(1950) <= (layer0_outputs(5412)) and not (layer0_outputs(656));
    outputs(1951) <= (layer0_outputs(1052)) and not (layer0_outputs(1432));
    outputs(1952) <= layer0_outputs(326);
    outputs(1953) <= (layer0_outputs(7423)) xor (layer0_outputs(1266));
    outputs(1954) <= (layer0_outputs(6935)) and not (layer0_outputs(4880));
    outputs(1955) <= layer0_outputs(5490);
    outputs(1956) <= layer0_outputs(172);
    outputs(1957) <= layer0_outputs(4061);
    outputs(1958) <= (layer0_outputs(2597)) xor (layer0_outputs(554));
    outputs(1959) <= not(layer0_outputs(7280)) or (layer0_outputs(2397));
    outputs(1960) <= not(layer0_outputs(4308)) or (layer0_outputs(2354));
    outputs(1961) <= not(layer0_outputs(6750)) or (layer0_outputs(5120));
    outputs(1962) <= not(layer0_outputs(1746));
    outputs(1963) <= (layer0_outputs(7226)) and not (layer0_outputs(6247));
    outputs(1964) <= (layer0_outputs(3029)) and not (layer0_outputs(7640));
    outputs(1965) <= (layer0_outputs(5326)) and not (layer0_outputs(3146));
    outputs(1966) <= (layer0_outputs(4804)) and not (layer0_outputs(4359));
    outputs(1967) <= layer0_outputs(130);
    outputs(1968) <= not(layer0_outputs(2354));
    outputs(1969) <= (layer0_outputs(4296)) xor (layer0_outputs(1938));
    outputs(1970) <= not(layer0_outputs(2926)) or (layer0_outputs(1968));
    outputs(1971) <= not(layer0_outputs(5106));
    outputs(1972) <= not(layer0_outputs(4535));
    outputs(1973) <= not(layer0_outputs(5510)) or (layer0_outputs(4514));
    outputs(1974) <= layer0_outputs(1411);
    outputs(1975) <= layer0_outputs(3499);
    outputs(1976) <= layer0_outputs(2760);
    outputs(1977) <= (layer0_outputs(3540)) and not (layer0_outputs(3653));
    outputs(1978) <= (layer0_outputs(622)) and not (layer0_outputs(1761));
    outputs(1979) <= (layer0_outputs(1323)) and (layer0_outputs(6037));
    outputs(1980) <= not((layer0_outputs(4380)) and (layer0_outputs(2711)));
    outputs(1981) <= layer0_outputs(7604);
    outputs(1982) <= not(layer0_outputs(2986));
    outputs(1983) <= (layer0_outputs(6871)) xor (layer0_outputs(6725));
    outputs(1984) <= (layer0_outputs(3891)) and not (layer0_outputs(4162));
    outputs(1985) <= not(layer0_outputs(2858)) or (layer0_outputs(3454));
    outputs(1986) <= (layer0_outputs(989)) or (layer0_outputs(1588));
    outputs(1987) <= not((layer0_outputs(3104)) or (layer0_outputs(2941)));
    outputs(1988) <= not((layer0_outputs(1222)) and (layer0_outputs(1099)));
    outputs(1989) <= (layer0_outputs(6772)) and (layer0_outputs(1498));
    outputs(1990) <= not(layer0_outputs(193));
    outputs(1991) <= not(layer0_outputs(1760)) or (layer0_outputs(6977));
    outputs(1992) <= layer0_outputs(4148);
    outputs(1993) <= (layer0_outputs(4859)) xor (layer0_outputs(6522));
    outputs(1994) <= layer0_outputs(2208);
    outputs(1995) <= layer0_outputs(5877);
    outputs(1996) <= layer0_outputs(1726);
    outputs(1997) <= not(layer0_outputs(7554)) or (layer0_outputs(3149));
    outputs(1998) <= not(layer0_outputs(5260));
    outputs(1999) <= not(layer0_outputs(4858));
    outputs(2000) <= layer0_outputs(3716);
    outputs(2001) <= not(layer0_outputs(2885));
    outputs(2002) <= not((layer0_outputs(5404)) xor (layer0_outputs(300)));
    outputs(2003) <= layer0_outputs(3942);
    outputs(2004) <= not((layer0_outputs(5668)) xor (layer0_outputs(6526)));
    outputs(2005) <= (layer0_outputs(4268)) or (layer0_outputs(3735));
    outputs(2006) <= not((layer0_outputs(6552)) xor (layer0_outputs(1485)));
    outputs(2007) <= not(layer0_outputs(4873));
    outputs(2008) <= layer0_outputs(3480);
    outputs(2009) <= layer0_outputs(413);
    outputs(2010) <= not(layer0_outputs(1034));
    outputs(2011) <= not((layer0_outputs(1860)) xor (layer0_outputs(4716)));
    outputs(2012) <= not((layer0_outputs(5261)) xor (layer0_outputs(5971)));
    outputs(2013) <= not(layer0_outputs(5286)) or (layer0_outputs(6093));
    outputs(2014) <= not(layer0_outputs(7471)) or (layer0_outputs(3536));
    outputs(2015) <= not(layer0_outputs(6925));
    outputs(2016) <= not(layer0_outputs(4293));
    outputs(2017) <= (layer0_outputs(4782)) xor (layer0_outputs(4696));
    outputs(2018) <= not((layer0_outputs(5685)) and (layer0_outputs(6353)));
    outputs(2019) <= not((layer0_outputs(3120)) and (layer0_outputs(6902)));
    outputs(2020) <= not(layer0_outputs(2711)) or (layer0_outputs(5582));
    outputs(2021) <= not(layer0_outputs(5363));
    outputs(2022) <= layer0_outputs(4406);
    outputs(2023) <= not((layer0_outputs(7192)) xor (layer0_outputs(6245)));
    outputs(2024) <= not((layer0_outputs(3423)) and (layer0_outputs(6231)));
    outputs(2025) <= layer0_outputs(3195);
    outputs(2026) <= (layer0_outputs(2523)) xor (layer0_outputs(7059));
    outputs(2027) <= layer0_outputs(2239);
    outputs(2028) <= not((layer0_outputs(2234)) xor (layer0_outputs(4360)));
    outputs(2029) <= layer0_outputs(3282);
    outputs(2030) <= not(layer0_outputs(465)) or (layer0_outputs(3000));
    outputs(2031) <= layer0_outputs(1092);
    outputs(2032) <= not((layer0_outputs(6735)) and (layer0_outputs(3784)));
    outputs(2033) <= (layer0_outputs(1595)) xor (layer0_outputs(694));
    outputs(2034) <= layer0_outputs(7052);
    outputs(2035) <= (layer0_outputs(6426)) or (layer0_outputs(6495));
    outputs(2036) <= not(layer0_outputs(7570)) or (layer0_outputs(6041));
    outputs(2037) <= not((layer0_outputs(4958)) xor (layer0_outputs(6184)));
    outputs(2038) <= not((layer0_outputs(3489)) or (layer0_outputs(335)));
    outputs(2039) <= (layer0_outputs(454)) xor (layer0_outputs(970));
    outputs(2040) <= not(layer0_outputs(2654));
    outputs(2041) <= layer0_outputs(2072);
    outputs(2042) <= not(layer0_outputs(6995)) or (layer0_outputs(3471));
    outputs(2043) <= not(layer0_outputs(4348));
    outputs(2044) <= (layer0_outputs(1016)) xor (layer0_outputs(5423));
    outputs(2045) <= layer0_outputs(49);
    outputs(2046) <= (layer0_outputs(693)) or (layer0_outputs(6037));
    outputs(2047) <= not((layer0_outputs(4412)) and (layer0_outputs(5243)));
    outputs(2048) <= not(layer0_outputs(864));
    outputs(2049) <= (layer0_outputs(7205)) and (layer0_outputs(447));
    outputs(2050) <= not(layer0_outputs(3120)) or (layer0_outputs(4589));
    outputs(2051) <= layer0_outputs(5571);
    outputs(2052) <= (layer0_outputs(3281)) xor (layer0_outputs(3622));
    outputs(2053) <= not((layer0_outputs(4190)) xor (layer0_outputs(3045)));
    outputs(2054) <= not((layer0_outputs(4909)) or (layer0_outputs(4227)));
    outputs(2055) <= layer0_outputs(1081);
    outputs(2056) <= not((layer0_outputs(5711)) and (layer0_outputs(73)));
    outputs(2057) <= layer0_outputs(6675);
    outputs(2058) <= not(layer0_outputs(6366)) or (layer0_outputs(4903));
    outputs(2059) <= not((layer0_outputs(1522)) xor (layer0_outputs(4658)));
    outputs(2060) <= (layer0_outputs(3212)) xor (layer0_outputs(4599));
    outputs(2061) <= layer0_outputs(4368);
    outputs(2062) <= (layer0_outputs(6625)) and not (layer0_outputs(4218));
    outputs(2063) <= (layer0_outputs(3565)) xor (layer0_outputs(1563));
    outputs(2064) <= not(layer0_outputs(2300));
    outputs(2065) <= layer0_outputs(3887);
    outputs(2066) <= (layer0_outputs(1189)) and (layer0_outputs(6372));
    outputs(2067) <= not(layer0_outputs(371));
    outputs(2068) <= not(layer0_outputs(3532)) or (layer0_outputs(2264));
    outputs(2069) <= (layer0_outputs(4445)) xor (layer0_outputs(5553));
    outputs(2070) <= not((layer0_outputs(5385)) xor (layer0_outputs(806)));
    outputs(2071) <= (layer0_outputs(3407)) xor (layer0_outputs(6637));
    outputs(2072) <= not(layer0_outputs(1090));
    outputs(2073) <= (layer0_outputs(4675)) xor (layer0_outputs(6729));
    outputs(2074) <= layer0_outputs(1355);
    outputs(2075) <= (layer0_outputs(905)) and (layer0_outputs(1916));
    outputs(2076) <= not(layer0_outputs(7570)) or (layer0_outputs(606));
    outputs(2077) <= not(layer0_outputs(3883));
    outputs(2078) <= (layer0_outputs(1527)) xor (layer0_outputs(2888));
    outputs(2079) <= layer0_outputs(2249);
    outputs(2080) <= not(layer0_outputs(5450));
    outputs(2081) <= layer0_outputs(3274);
    outputs(2082) <= not((layer0_outputs(4578)) or (layer0_outputs(4698)));
    outputs(2083) <= layer0_outputs(346);
    outputs(2084) <= not(layer0_outputs(7521));
    outputs(2085) <= layer0_outputs(7076);
    outputs(2086) <= not((layer0_outputs(6082)) or (layer0_outputs(7405)));
    outputs(2087) <= not(layer0_outputs(411)) or (layer0_outputs(4428));
    outputs(2088) <= not(layer0_outputs(5899)) or (layer0_outputs(3948));
    outputs(2089) <= not((layer0_outputs(2819)) xor (layer0_outputs(6770)));
    outputs(2090) <= (layer0_outputs(939)) and not (layer0_outputs(5831));
    outputs(2091) <= not(layer0_outputs(3584));
    outputs(2092) <= (layer0_outputs(4777)) or (layer0_outputs(4384));
    outputs(2093) <= not(layer0_outputs(421));
    outputs(2094) <= (layer0_outputs(3965)) xor (layer0_outputs(457));
    outputs(2095) <= not(layer0_outputs(3495));
    outputs(2096) <= (layer0_outputs(857)) or (layer0_outputs(3859));
    outputs(2097) <= not(layer0_outputs(3656));
    outputs(2098) <= (layer0_outputs(4616)) and not (layer0_outputs(2731));
    outputs(2099) <= not(layer0_outputs(3731));
    outputs(2100) <= (layer0_outputs(1296)) and (layer0_outputs(1665));
    outputs(2101) <= not(layer0_outputs(6869));
    outputs(2102) <= not((layer0_outputs(4033)) or (layer0_outputs(4467)));
    outputs(2103) <= (layer0_outputs(4666)) xor (layer0_outputs(2692));
    outputs(2104) <= not(layer0_outputs(2694));
    outputs(2105) <= layer0_outputs(3418);
    outputs(2106) <= not((layer0_outputs(2087)) xor (layer0_outputs(1748)));
    outputs(2107) <= layer0_outputs(5467);
    outputs(2108) <= layer0_outputs(3153);
    outputs(2109) <= not((layer0_outputs(1961)) and (layer0_outputs(4096)));
    outputs(2110) <= not(layer0_outputs(4332));
    outputs(2111) <= not(layer0_outputs(4486));
    outputs(2112) <= layer0_outputs(405);
    outputs(2113) <= layer0_outputs(6908);
    outputs(2114) <= not(layer0_outputs(1283));
    outputs(2115) <= not((layer0_outputs(7290)) and (layer0_outputs(5962)));
    outputs(2116) <= not(layer0_outputs(1259));
    outputs(2117) <= (layer0_outputs(7062)) xor (layer0_outputs(5452));
    outputs(2118) <= not((layer0_outputs(4888)) or (layer0_outputs(6522)));
    outputs(2119) <= layer0_outputs(400);
    outputs(2120) <= layer0_outputs(4831);
    outputs(2121) <= not((layer0_outputs(2929)) and (layer0_outputs(5838)));
    outputs(2122) <= layer0_outputs(4830);
    outputs(2123) <= layer0_outputs(981);
    outputs(2124) <= not(layer0_outputs(1552));
    outputs(2125) <= not((layer0_outputs(6240)) and (layer0_outputs(979)));
    outputs(2126) <= not(layer0_outputs(7170));
    outputs(2127) <= not(layer0_outputs(7019));
    outputs(2128) <= layer0_outputs(7427);
    outputs(2129) <= not(layer0_outputs(4971));
    outputs(2130) <= (layer0_outputs(4687)) and not (layer0_outputs(6844));
    outputs(2131) <= (layer0_outputs(4301)) or (layer0_outputs(5180));
    outputs(2132) <= not(layer0_outputs(6073));
    outputs(2133) <= layer0_outputs(6305);
    outputs(2134) <= not((layer0_outputs(1638)) xor (layer0_outputs(1892)));
    outputs(2135) <= layer0_outputs(7511);
    outputs(2136) <= (layer0_outputs(4652)) xor (layer0_outputs(6408));
    outputs(2137) <= not((layer0_outputs(7166)) xor (layer0_outputs(4943)));
    outputs(2138) <= (layer0_outputs(6602)) and not (layer0_outputs(4510));
    outputs(2139) <= (layer0_outputs(5206)) xor (layer0_outputs(2442));
    outputs(2140) <= not(layer0_outputs(3137));
    outputs(2141) <= layer0_outputs(2157);
    outputs(2142) <= layer0_outputs(4743);
    outputs(2143) <= (layer0_outputs(643)) or (layer0_outputs(4136));
    outputs(2144) <= (layer0_outputs(962)) or (layer0_outputs(2324));
    outputs(2145) <= (layer0_outputs(5785)) xor (layer0_outputs(362));
    outputs(2146) <= not(layer0_outputs(2172));
    outputs(2147) <= not(layer0_outputs(1757)) or (layer0_outputs(872));
    outputs(2148) <= not(layer0_outputs(201)) or (layer0_outputs(1129));
    outputs(2149) <= (layer0_outputs(3901)) and (layer0_outputs(1729));
    outputs(2150) <= not((layer0_outputs(6610)) or (layer0_outputs(6257)));
    outputs(2151) <= layer0_outputs(1047);
    outputs(2152) <= (layer0_outputs(1249)) or (layer0_outputs(4974));
    outputs(2153) <= layer0_outputs(836);
    outputs(2154) <= layer0_outputs(4309);
    outputs(2155) <= (layer0_outputs(3598)) and not (layer0_outputs(7400));
    outputs(2156) <= (layer0_outputs(2658)) or (layer0_outputs(2635));
    outputs(2157) <= not(layer0_outputs(1503));
    outputs(2158) <= not((layer0_outputs(788)) xor (layer0_outputs(4799)));
    outputs(2159) <= not(layer0_outputs(5998));
    outputs(2160) <= not(layer0_outputs(4548)) or (layer0_outputs(3535));
    outputs(2161) <= not(layer0_outputs(2536));
    outputs(2162) <= not((layer0_outputs(5426)) and (layer0_outputs(2863)));
    outputs(2163) <= not((layer0_outputs(1228)) xor (layer0_outputs(5825)));
    outputs(2164) <= not((layer0_outputs(5216)) xor (layer0_outputs(6534)));
    outputs(2165) <= layer0_outputs(3332);
    outputs(2166) <= (layer0_outputs(5566)) xor (layer0_outputs(135));
    outputs(2167) <= not(layer0_outputs(5362));
    outputs(2168) <= not(layer0_outputs(2593)) or (layer0_outputs(7636));
    outputs(2169) <= layer0_outputs(7444);
    outputs(2170) <= not((layer0_outputs(6582)) and (layer0_outputs(7065)));
    outputs(2171) <= not(layer0_outputs(4920));
    outputs(2172) <= not((layer0_outputs(4601)) xor (layer0_outputs(757)));
    outputs(2173) <= not((layer0_outputs(2999)) xor (layer0_outputs(890)));
    outputs(2174) <= not((layer0_outputs(5357)) and (layer0_outputs(2081)));
    outputs(2175) <= (layer0_outputs(1790)) xor (layer0_outputs(1112));
    outputs(2176) <= not(layer0_outputs(3519)) or (layer0_outputs(6681));
    outputs(2177) <= (layer0_outputs(3680)) and (layer0_outputs(57));
    outputs(2178) <= (layer0_outputs(3681)) and (layer0_outputs(5153));
    outputs(2179) <= not(layer0_outputs(6296));
    outputs(2180) <= not(layer0_outputs(3584)) or (layer0_outputs(4891));
    outputs(2181) <= layer0_outputs(4266);
    outputs(2182) <= not(layer0_outputs(6368));
    outputs(2183) <= not((layer0_outputs(2511)) and (layer0_outputs(1786)));
    outputs(2184) <= not(layer0_outputs(6529)) or (layer0_outputs(1110));
    outputs(2185) <= not(layer0_outputs(4224)) or (layer0_outputs(5964));
    outputs(2186) <= not((layer0_outputs(5733)) xor (layer0_outputs(4678)));
    outputs(2187) <= not((layer0_outputs(1158)) or (layer0_outputs(1317)));
    outputs(2188) <= not((layer0_outputs(3156)) and (layer0_outputs(780)));
    outputs(2189) <= not(layer0_outputs(168));
    outputs(2190) <= not(layer0_outputs(3062));
    outputs(2191) <= not(layer0_outputs(3465));
    outputs(2192) <= not((layer0_outputs(2365)) xor (layer0_outputs(1868)));
    outputs(2193) <= not(layer0_outputs(1615));
    outputs(2194) <= (layer0_outputs(4291)) or (layer0_outputs(458));
    outputs(2195) <= layer0_outputs(5568);
    outputs(2196) <= layer0_outputs(7598);
    outputs(2197) <= (layer0_outputs(3725)) and not (layer0_outputs(2348));
    outputs(2198) <= layer0_outputs(3695);
    outputs(2199) <= (layer0_outputs(1295)) xor (layer0_outputs(1313));
    outputs(2200) <= not(layer0_outputs(3931));
    outputs(2201) <= layer0_outputs(935);
    outputs(2202) <= not(layer0_outputs(1359));
    outputs(2203) <= (layer0_outputs(2516)) and (layer0_outputs(4699));
    outputs(2204) <= not(layer0_outputs(2467));
    outputs(2205) <= (layer0_outputs(2272)) and not (layer0_outputs(6250));
    outputs(2206) <= (layer0_outputs(2422)) or (layer0_outputs(911));
    outputs(2207) <= (layer0_outputs(5479)) xor (layer0_outputs(2977));
    outputs(2208) <= layer0_outputs(6092);
    outputs(2209) <= (layer0_outputs(4564)) or (layer0_outputs(4282));
    outputs(2210) <= layer0_outputs(3734);
    outputs(2211) <= not(layer0_outputs(4587));
    outputs(2212) <= not(layer0_outputs(7084)) or (layer0_outputs(494));
    outputs(2213) <= not(layer0_outputs(6427));
    outputs(2214) <= (layer0_outputs(4705)) and not (layer0_outputs(6848));
    outputs(2215) <= (layer0_outputs(1978)) or (layer0_outputs(7539));
    outputs(2216) <= not((layer0_outputs(4565)) xor (layer0_outputs(5481)));
    outputs(2217) <= layer0_outputs(1213);
    outputs(2218) <= (layer0_outputs(981)) and not (layer0_outputs(4711));
    outputs(2219) <= not(layer0_outputs(6396)) or (layer0_outputs(3483));
    outputs(2220) <= (layer0_outputs(2864)) xor (layer0_outputs(1556));
    outputs(2221) <= not(layer0_outputs(4161)) or (layer0_outputs(4173));
    outputs(2222) <= layer0_outputs(3088);
    outputs(2223) <= not(layer0_outputs(5038)) or (layer0_outputs(5943));
    outputs(2224) <= not(layer0_outputs(260));
    outputs(2225) <= (layer0_outputs(5863)) xor (layer0_outputs(801));
    outputs(2226) <= not(layer0_outputs(1424));
    outputs(2227) <= not((layer0_outputs(4744)) and (layer0_outputs(4321)));
    outputs(2228) <= not((layer0_outputs(7476)) xor (layer0_outputs(2542)));
    outputs(2229) <= not(layer0_outputs(3617));
    outputs(2230) <= not(layer0_outputs(777));
    outputs(2231) <= not(layer0_outputs(5228));
    outputs(2232) <= not(layer0_outputs(6850));
    outputs(2233) <= not(layer0_outputs(123));
    outputs(2234) <= (layer0_outputs(4491)) and not (layer0_outputs(1342));
    outputs(2235) <= layer0_outputs(7462);
    outputs(2236) <= not((layer0_outputs(760)) xor (layer0_outputs(1444)));
    outputs(2237) <= layer0_outputs(415);
    outputs(2238) <= not((layer0_outputs(5650)) and (layer0_outputs(7225)));
    outputs(2239) <= (layer0_outputs(2329)) xor (layer0_outputs(591));
    outputs(2240) <= not((layer0_outputs(7561)) and (layer0_outputs(1730)));
    outputs(2241) <= not(layer0_outputs(5972)) or (layer0_outputs(2938));
    outputs(2242) <= layer0_outputs(366);
    outputs(2243) <= layer0_outputs(2884);
    outputs(2244) <= layer0_outputs(3818);
    outputs(2245) <= not((layer0_outputs(1417)) xor (layer0_outputs(2381)));
    outputs(2246) <= not(layer0_outputs(3804));
    outputs(2247) <= layer0_outputs(5314);
    outputs(2248) <= layer0_outputs(3961);
    outputs(2249) <= not(layer0_outputs(2302));
    outputs(2250) <= (layer0_outputs(1678)) and (layer0_outputs(1200));
    outputs(2251) <= layer0_outputs(915);
    outputs(2252) <= not((layer0_outputs(4678)) xor (layer0_outputs(7673)));
    outputs(2253) <= (layer0_outputs(4352)) and (layer0_outputs(1033));
    outputs(2254) <= layer0_outputs(3380);
    outputs(2255) <= layer0_outputs(6406);
    outputs(2256) <= (layer0_outputs(4014)) and not (layer0_outputs(2902));
    outputs(2257) <= layer0_outputs(4803);
    outputs(2258) <= not((layer0_outputs(6528)) and (layer0_outputs(661)));
    outputs(2259) <= layer0_outputs(4230);
    outputs(2260) <= not(layer0_outputs(2165)) or (layer0_outputs(85));
    outputs(2261) <= (layer0_outputs(1646)) xor (layer0_outputs(4671));
    outputs(2262) <= not((layer0_outputs(4832)) and (layer0_outputs(4857)));
    outputs(2263) <= not(layer0_outputs(146));
    outputs(2264) <= layer0_outputs(6365);
    outputs(2265) <= (layer0_outputs(3853)) and (layer0_outputs(2339));
    outputs(2266) <= (layer0_outputs(351)) and not (layer0_outputs(1901));
    outputs(2267) <= (layer0_outputs(4398)) and not (layer0_outputs(1561));
    outputs(2268) <= layer0_outputs(2078);
    outputs(2269) <= not(layer0_outputs(4050)) or (layer0_outputs(3222));
    outputs(2270) <= not(layer0_outputs(2773)) or (layer0_outputs(2992));
    outputs(2271) <= not(layer0_outputs(5879));
    outputs(2272) <= not(layer0_outputs(4662));
    outputs(2273) <= layer0_outputs(7276);
    outputs(2274) <= not((layer0_outputs(6343)) and (layer0_outputs(2114)));
    outputs(2275) <= (layer0_outputs(6506)) or (layer0_outputs(3308));
    outputs(2276) <= (layer0_outputs(5188)) xor (layer0_outputs(2125));
    outputs(2277) <= not(layer0_outputs(3684));
    outputs(2278) <= (layer0_outputs(4544)) and not (layer0_outputs(1659));
    outputs(2279) <= layer0_outputs(174);
    outputs(2280) <= (layer0_outputs(1122)) xor (layer0_outputs(448));
    outputs(2281) <= (layer0_outputs(6820)) and (layer0_outputs(1139));
    outputs(2282) <= layer0_outputs(6069);
    outputs(2283) <= not(layer0_outputs(4952)) or (layer0_outputs(4274));
    outputs(2284) <= not(layer0_outputs(5169));
    outputs(2285) <= not(layer0_outputs(4045));
    outputs(2286) <= not(layer0_outputs(2913)) or (layer0_outputs(5459));
    outputs(2287) <= not(layer0_outputs(561));
    outputs(2288) <= not(layer0_outputs(6412));
    outputs(2289) <= not(layer0_outputs(568));
    outputs(2290) <= not(layer0_outputs(5874));
    outputs(2291) <= layer0_outputs(2758);
    outputs(2292) <= not(layer0_outputs(5540));
    outputs(2293) <= not(layer0_outputs(3729)) or (layer0_outputs(80));
    outputs(2294) <= (layer0_outputs(4489)) and not (layer0_outputs(2704));
    outputs(2295) <= not(layer0_outputs(5318)) or (layer0_outputs(3943));
    outputs(2296) <= layer0_outputs(48);
    outputs(2297) <= layer0_outputs(37);
    outputs(2298) <= (layer0_outputs(2651)) and (layer0_outputs(3030));
    outputs(2299) <= (layer0_outputs(6142)) or (layer0_outputs(4194));
    outputs(2300) <= not((layer0_outputs(3977)) xor (layer0_outputs(5894)));
    outputs(2301) <= layer0_outputs(6381);
    outputs(2302) <= not(layer0_outputs(2322)) or (layer0_outputs(3995));
    outputs(2303) <= not((layer0_outputs(3009)) or (layer0_outputs(2402)));
    outputs(2304) <= not((layer0_outputs(5410)) xor (layer0_outputs(2037)));
    outputs(2305) <= not((layer0_outputs(4118)) xor (layer0_outputs(3262)));
    outputs(2306) <= layer0_outputs(6287);
    outputs(2307) <= not((layer0_outputs(1216)) and (layer0_outputs(1995)));
    outputs(2308) <= (layer0_outputs(5820)) and not (layer0_outputs(2001));
    outputs(2309) <= not((layer0_outputs(4066)) and (layer0_outputs(7588)));
    outputs(2310) <= not(layer0_outputs(6944));
    outputs(2311) <= (layer0_outputs(1383)) xor (layer0_outputs(4921));
    outputs(2312) <= layer0_outputs(2473);
    outputs(2313) <= (layer0_outputs(7397)) or (layer0_outputs(3442));
    outputs(2314) <= layer0_outputs(5010);
    outputs(2315) <= not((layer0_outputs(4138)) and (layer0_outputs(2491)));
    outputs(2316) <= (layer0_outputs(7209)) xor (layer0_outputs(6721));
    outputs(2317) <= not(layer0_outputs(6778));
    outputs(2318) <= layer0_outputs(299);
    outputs(2319) <= not(layer0_outputs(1095));
    outputs(2320) <= not(layer0_outputs(2921));
    outputs(2321) <= not((layer0_outputs(6568)) or (layer0_outputs(6679)));
    outputs(2322) <= (layer0_outputs(6872)) and not (layer0_outputs(3666));
    outputs(2323) <= (layer0_outputs(4396)) xor (layer0_outputs(3904));
    outputs(2324) <= not(layer0_outputs(4367));
    outputs(2325) <= (layer0_outputs(1833)) and (layer0_outputs(5249));
    outputs(2326) <= not((layer0_outputs(7431)) or (layer0_outputs(280)));
    outputs(2327) <= (layer0_outputs(1994)) and (layer0_outputs(5888));
    outputs(2328) <= layer0_outputs(6825);
    outputs(2329) <= not(layer0_outputs(6510));
    outputs(2330) <= layer0_outputs(4813);
    outputs(2331) <= not((layer0_outputs(4530)) xor (layer0_outputs(7113)));
    outputs(2332) <= layer0_outputs(7299);
    outputs(2333) <= not((layer0_outputs(891)) xor (layer0_outputs(3917)));
    outputs(2334) <= layer0_outputs(5255);
    outputs(2335) <= not((layer0_outputs(651)) or (layer0_outputs(626)));
    outputs(2336) <= (layer0_outputs(5104)) and (layer0_outputs(4592));
    outputs(2337) <= not(layer0_outputs(1075));
    outputs(2338) <= (layer0_outputs(174)) and not (layer0_outputs(6477));
    outputs(2339) <= (layer0_outputs(7414)) and (layer0_outputs(4900));
    outputs(2340) <= (layer0_outputs(4911)) xor (layer0_outputs(4068));
    outputs(2341) <= not(layer0_outputs(3679));
    outputs(2342) <= (layer0_outputs(4729)) and (layer0_outputs(903));
    outputs(2343) <= not((layer0_outputs(1351)) xor (layer0_outputs(2663)));
    outputs(2344) <= not((layer0_outputs(6388)) or (layer0_outputs(4336)));
    outputs(2345) <= layer0_outputs(7306);
    outputs(2346) <= (layer0_outputs(2714)) and not (layer0_outputs(432));
    outputs(2347) <= (layer0_outputs(674)) and (layer0_outputs(6036));
    outputs(2348) <= layer0_outputs(4981);
    outputs(2349) <= (layer0_outputs(4356)) and not (layer0_outputs(6236));
    outputs(2350) <= (layer0_outputs(5046)) xor (layer0_outputs(6010));
    outputs(2351) <= (layer0_outputs(4665)) and not (layer0_outputs(899));
    outputs(2352) <= layer0_outputs(2911);
    outputs(2353) <= not((layer0_outputs(6398)) xor (layer0_outputs(2691)));
    outputs(2354) <= (layer0_outputs(5635)) and not (layer0_outputs(6576));
    outputs(2355) <= not(layer0_outputs(1185)) or (layer0_outputs(880));
    outputs(2356) <= not(layer0_outputs(3822));
    outputs(2357) <= not(layer0_outputs(1017));
    outputs(2358) <= not((layer0_outputs(1253)) and (layer0_outputs(5083)));
    outputs(2359) <= layer0_outputs(6775);
    outputs(2360) <= not((layer0_outputs(7258)) or (layer0_outputs(3242)));
    outputs(2361) <= layer0_outputs(5891);
    outputs(2362) <= (layer0_outputs(7552)) and (layer0_outputs(4807));
    outputs(2363) <= layer0_outputs(6998);
    outputs(2364) <= not((layer0_outputs(6070)) or (layer0_outputs(7309)));
    outputs(2365) <= not(layer0_outputs(32));
    outputs(2366) <= layer0_outputs(2006);
    outputs(2367) <= not((layer0_outputs(6309)) or (layer0_outputs(2649)));
    outputs(2368) <= (layer0_outputs(7045)) and (layer0_outputs(3672));
    outputs(2369) <= not((layer0_outputs(7649)) or (layer0_outputs(2751)));
    outputs(2370) <= layer0_outputs(5583);
    outputs(2371) <= not((layer0_outputs(6951)) xor (layer0_outputs(6289)));
    outputs(2372) <= layer0_outputs(5430);
    outputs(2373) <= not(layer0_outputs(7437));
    outputs(2374) <= not(layer0_outputs(818)) or (layer0_outputs(4009));
    outputs(2375) <= not((layer0_outputs(497)) and (layer0_outputs(3960)));
    outputs(2376) <= layer0_outputs(2750);
    outputs(2377) <= layer0_outputs(10);
    outputs(2378) <= not(layer0_outputs(1744)) or (layer0_outputs(3834));
    outputs(2379) <= layer0_outputs(706);
    outputs(2380) <= not((layer0_outputs(1952)) and (layer0_outputs(2611)));
    outputs(2381) <= not(layer0_outputs(7531));
    outputs(2382) <= not(layer0_outputs(2939));
    outputs(2383) <= layer0_outputs(5735);
    outputs(2384) <= (layer0_outputs(1106)) and not (layer0_outputs(2748));
    outputs(2385) <= (layer0_outputs(3582)) xor (layer0_outputs(7033));
    outputs(2386) <= layer0_outputs(1579);
    outputs(2387) <= not(layer0_outputs(5875)) or (layer0_outputs(809));
    outputs(2388) <= layer0_outputs(6765);
    outputs(2389) <= layer0_outputs(2213);
    outputs(2390) <= (layer0_outputs(4062)) or (layer0_outputs(3590));
    outputs(2391) <= not((layer0_outputs(4226)) and (layer0_outputs(6562)));
    outputs(2392) <= not(layer0_outputs(4040));
    outputs(2393) <= layer0_outputs(4042);
    outputs(2394) <= not(layer0_outputs(741)) or (layer0_outputs(2573));
    outputs(2395) <= not(layer0_outputs(5628));
    outputs(2396) <= layer0_outputs(926);
    outputs(2397) <= not(layer0_outputs(1497));
    outputs(2398) <= layer0_outputs(310);
    outputs(2399) <= (layer0_outputs(2543)) xor (layer0_outputs(6646));
    outputs(2400) <= (layer0_outputs(143)) and (layer0_outputs(6661));
    outputs(2401) <= layer0_outputs(6049);
    outputs(2402) <= (layer0_outputs(2754)) and not (layer0_outputs(3275));
    outputs(2403) <= layer0_outputs(1364);
    outputs(2404) <= (layer0_outputs(954)) and not (layer0_outputs(4201));
    outputs(2405) <= not(layer0_outputs(5858));
    outputs(2406) <= (layer0_outputs(1711)) and not (layer0_outputs(6649));
    outputs(2407) <= not(layer0_outputs(1427));
    outputs(2408) <= (layer0_outputs(5507)) or (layer0_outputs(1770));
    outputs(2409) <= (layer0_outputs(5190)) xor (layer0_outputs(1193));
    outputs(2410) <= not((layer0_outputs(622)) xor (layer0_outputs(3272)));
    outputs(2411) <= layer0_outputs(6315);
    outputs(2412) <= not(layer0_outputs(2412));
    outputs(2413) <= (layer0_outputs(2301)) and (layer0_outputs(1229));
    outputs(2414) <= (layer0_outputs(3578)) and not (layer0_outputs(1206));
    outputs(2415) <= layer0_outputs(3985);
    outputs(2416) <= not(layer0_outputs(4549));
    outputs(2417) <= not(layer0_outputs(1343));
    outputs(2418) <= (layer0_outputs(3534)) and not (layer0_outputs(7358));
    outputs(2419) <= (layer0_outputs(4488)) or (layer0_outputs(1950));
    outputs(2420) <= (layer0_outputs(4998)) and not (layer0_outputs(6419));
    outputs(2421) <= (layer0_outputs(3653)) or (layer0_outputs(349));
    outputs(2422) <= not(layer0_outputs(1473));
    outputs(2423) <= (layer0_outputs(681)) and not (layer0_outputs(2247));
    outputs(2424) <= not((layer0_outputs(3603)) or (layer0_outputs(5986)));
    outputs(2425) <= layer0_outputs(859);
    outputs(2426) <= not(layer0_outputs(3122));
    outputs(2427) <= not(layer0_outputs(2127)) or (layer0_outputs(1026));
    outputs(2428) <= not(layer0_outputs(6786)) or (layer0_outputs(5624));
    outputs(2429) <= layer0_outputs(1480);
    outputs(2430) <= (layer0_outputs(6736)) and (layer0_outputs(4407));
    outputs(2431) <= (layer0_outputs(6483)) or (layer0_outputs(1836));
    outputs(2432) <= not(layer0_outputs(7032));
    outputs(2433) <= (layer0_outputs(2487)) and not (layer0_outputs(1228));
    outputs(2434) <= not(layer0_outputs(5565)) or (layer0_outputs(7627));
    outputs(2435) <= (layer0_outputs(4512)) xor (layer0_outputs(7639));
    outputs(2436) <= layer0_outputs(3018);
    outputs(2437) <= not((layer0_outputs(330)) xor (layer0_outputs(4046)));
    outputs(2438) <= not((layer0_outputs(7525)) xor (layer0_outputs(4833)));
    outputs(2439) <= not(layer0_outputs(3924));
    outputs(2440) <= not(layer0_outputs(7242));
    outputs(2441) <= (layer0_outputs(5393)) xor (layer0_outputs(2719));
    outputs(2442) <= layer0_outputs(6669);
    outputs(2443) <= not((layer0_outputs(7509)) and (layer0_outputs(5230)));
    outputs(2444) <= layer0_outputs(4169);
    outputs(2445) <= not(layer0_outputs(1919));
    outputs(2446) <= (layer0_outputs(5413)) and not (layer0_outputs(2067));
    outputs(2447) <= not(layer0_outputs(4023));
    outputs(2448) <= (layer0_outputs(5356)) xor (layer0_outputs(5622));
    outputs(2449) <= layer0_outputs(3322);
    outputs(2450) <= (layer0_outputs(6515)) and not (layer0_outputs(7492));
    outputs(2451) <= not((layer0_outputs(4303)) or (layer0_outputs(7167)));
    outputs(2452) <= (layer0_outputs(1723)) xor (layer0_outputs(5413));
    outputs(2453) <= (layer0_outputs(3788)) and not (layer0_outputs(6599));
    outputs(2454) <= not((layer0_outputs(5449)) xor (layer0_outputs(7418)));
    outputs(2455) <= not(layer0_outputs(2380)) or (layer0_outputs(5651));
    outputs(2456) <= (layer0_outputs(5760)) and not (layer0_outputs(1327));
    outputs(2457) <= (layer0_outputs(5035)) and not (layer0_outputs(4350));
    outputs(2458) <= not(layer0_outputs(7335)) or (layer0_outputs(5749));
    outputs(2459) <= not(layer0_outputs(5829)) or (layer0_outputs(252));
    outputs(2460) <= not(layer0_outputs(6867));
    outputs(2461) <= not((layer0_outputs(7590)) or (layer0_outputs(5626)));
    outputs(2462) <= not(layer0_outputs(7409));
    outputs(2463) <= not(layer0_outputs(3187));
    outputs(2464) <= not(layer0_outputs(2647));
    outputs(2465) <= (layer0_outputs(1770)) and (layer0_outputs(997));
    outputs(2466) <= not(layer0_outputs(2424));
    outputs(2467) <= not(layer0_outputs(5737));
    outputs(2468) <= layer0_outputs(2416);
    outputs(2469) <= (layer0_outputs(788)) and (layer0_outputs(623));
    outputs(2470) <= layer0_outputs(803);
    outputs(2471) <= (layer0_outputs(4566)) and (layer0_outputs(1684));
    outputs(2472) <= layer0_outputs(3513);
    outputs(2473) <= not((layer0_outputs(1435)) or (layer0_outputs(7241)));
    outputs(2474) <= not(layer0_outputs(2875));
    outputs(2475) <= layer0_outputs(963);
    outputs(2476) <= layer0_outputs(6479);
    outputs(2477) <= (layer0_outputs(934)) xor (layer0_outputs(2715));
    outputs(2478) <= not((layer0_outputs(5836)) xor (layer0_outputs(6190)));
    outputs(2479) <= (layer0_outputs(1695)) and not (layer0_outputs(7501));
    outputs(2480) <= (layer0_outputs(970)) xor (layer0_outputs(4838));
    outputs(2481) <= (layer0_outputs(584)) and (layer0_outputs(5570));
    outputs(2482) <= (layer0_outputs(1799)) xor (layer0_outputs(4725));
    outputs(2483) <= (layer0_outputs(6775)) and not (layer0_outputs(2605));
    outputs(2484) <= not(layer0_outputs(376));
    outputs(2485) <= (layer0_outputs(5840)) and not (layer0_outputs(4631));
    outputs(2486) <= not(layer0_outputs(3630)) or (layer0_outputs(7000));
    outputs(2487) <= not((layer0_outputs(7040)) xor (layer0_outputs(3094)));
    outputs(2488) <= not(layer0_outputs(420));
    outputs(2489) <= not(layer0_outputs(3781)) or (layer0_outputs(6726));
    outputs(2490) <= (layer0_outputs(3145)) and not (layer0_outputs(589));
    outputs(2491) <= layer0_outputs(4516);
    outputs(2492) <= (layer0_outputs(1688)) xor (layer0_outputs(5674));
    outputs(2493) <= not(layer0_outputs(790));
    outputs(2494) <= not((layer0_outputs(6807)) or (layer0_outputs(1107)));
    outputs(2495) <= layer0_outputs(3427);
    outputs(2496) <= (layer0_outputs(5605)) and (layer0_outputs(2452));
    outputs(2497) <= layer0_outputs(4225);
    outputs(2498) <= not((layer0_outputs(634)) and (layer0_outputs(180)));
    outputs(2499) <= not(layer0_outputs(1637)) or (layer0_outputs(6841));
    outputs(2500) <= layer0_outputs(7636);
    outputs(2501) <= not(layer0_outputs(5268));
    outputs(2502) <= not(layer0_outputs(1934));
    outputs(2503) <= (layer0_outputs(7062)) and (layer0_outputs(6900));
    outputs(2504) <= (layer0_outputs(802)) and (layer0_outputs(1911));
    outputs(2505) <= not(layer0_outputs(2605));
    outputs(2506) <= not((layer0_outputs(2136)) and (layer0_outputs(7225)));
    outputs(2507) <= not(layer0_outputs(2676));
    outputs(2508) <= layer0_outputs(1941);
    outputs(2509) <= not((layer0_outputs(312)) xor (layer0_outputs(7089)));
    outputs(2510) <= layer0_outputs(6464);
    outputs(2511) <= (layer0_outputs(3245)) and (layer0_outputs(2468));
    outputs(2512) <= not(layer0_outputs(1831));
    outputs(2513) <= (layer0_outputs(3361)) xor (layer0_outputs(2624));
    outputs(2514) <= layer0_outputs(5072);
    outputs(2515) <= not(layer0_outputs(6638));
    outputs(2516) <= layer0_outputs(4590);
    outputs(2517) <= layer0_outputs(3306);
    outputs(2518) <= (layer0_outputs(6823)) xor (layer0_outputs(3312));
    outputs(2519) <= (layer0_outputs(4660)) and not (layer0_outputs(4935));
    outputs(2520) <= (layer0_outputs(3482)) and not (layer0_outputs(287));
    outputs(2521) <= (layer0_outputs(6926)) and not (layer0_outputs(324));
    outputs(2522) <= not(layer0_outputs(7658)) or (layer0_outputs(7614));
    outputs(2523) <= not(layer0_outputs(6645)) or (layer0_outputs(4754));
    outputs(2524) <= not((layer0_outputs(52)) xor (layer0_outputs(6372)));
    outputs(2525) <= (layer0_outputs(6449)) xor (layer0_outputs(6831));
    outputs(2526) <= (layer0_outputs(7660)) xor (layer0_outputs(6377));
    outputs(2527) <= (layer0_outputs(4476)) and not (layer0_outputs(1271));
    outputs(2528) <= not((layer0_outputs(1917)) or (layer0_outputs(4482)));
    outputs(2529) <= not((layer0_outputs(325)) xor (layer0_outputs(2580)));
    outputs(2530) <= (layer0_outputs(7259)) or (layer0_outputs(5803));
    outputs(2531) <= not(layer0_outputs(724));
    outputs(2532) <= layer0_outputs(1602);
    outputs(2533) <= (layer0_outputs(2998)) xor (layer0_outputs(3616));
    outputs(2534) <= (layer0_outputs(2173)) or (layer0_outputs(7300));
    outputs(2535) <= not(layer0_outputs(7103));
    outputs(2536) <= (layer0_outputs(7566)) xor (layer0_outputs(2371));
    outputs(2537) <= not((layer0_outputs(542)) xor (layer0_outputs(5215)));
    outputs(2538) <= layer0_outputs(6317);
    outputs(2539) <= (layer0_outputs(4139)) and not (layer0_outputs(4383));
    outputs(2540) <= (layer0_outputs(1385)) xor (layer0_outputs(5799));
    outputs(2541) <= (layer0_outputs(6574)) xor (layer0_outputs(1163));
    outputs(2542) <= layer0_outputs(6275);
    outputs(2543) <= not((layer0_outputs(694)) or (layer0_outputs(4919)));
    outputs(2544) <= not(layer0_outputs(2253));
    outputs(2545) <= not(layer0_outputs(567));
    outputs(2546) <= not(layer0_outputs(5441));
    outputs(2547) <= not(layer0_outputs(3912));
    outputs(2548) <= not((layer0_outputs(4844)) xor (layer0_outputs(6732)));
    outputs(2549) <= not((layer0_outputs(850)) or (layer0_outputs(6205)));
    outputs(2550) <= not(layer0_outputs(3313)) or (layer0_outputs(2235));
    outputs(2551) <= not(layer0_outputs(6689));
    outputs(2552) <= not((layer0_outputs(1078)) xor (layer0_outputs(4214)));
    outputs(2553) <= not((layer0_outputs(240)) and (layer0_outputs(6064)));
    outputs(2554) <= (layer0_outputs(1843)) and (layer0_outputs(1945));
    outputs(2555) <= not(layer0_outputs(7297));
    outputs(2556) <= (layer0_outputs(5386)) and not (layer0_outputs(1875));
    outputs(2557) <= layer0_outputs(4539);
    outputs(2558) <= layer0_outputs(4841);
    outputs(2559) <= (layer0_outputs(5266)) or (layer0_outputs(2344));
    outputs(2560) <= not(layer0_outputs(1575)) or (layer0_outputs(2376));
    outputs(2561) <= not(layer0_outputs(378)) or (layer0_outputs(5719));
    outputs(2562) <= layer0_outputs(7257);
    outputs(2563) <= not(layer0_outputs(2000)) or (layer0_outputs(5074));
    outputs(2564) <= not((layer0_outputs(4015)) and (layer0_outputs(6577)));
    outputs(2565) <= (layer0_outputs(2758)) and not (layer0_outputs(241));
    outputs(2566) <= (layer0_outputs(6671)) and not (layer0_outputs(249));
    outputs(2567) <= layer0_outputs(2459);
    outputs(2568) <= layer0_outputs(3418);
    outputs(2569) <= not(layer0_outputs(2020));
    outputs(2570) <= layer0_outputs(1345);
    outputs(2571) <= not((layer0_outputs(3527)) or (layer0_outputs(133)));
    outputs(2572) <= not(layer0_outputs(6818));
    outputs(2573) <= not(layer0_outputs(7352));
    outputs(2574) <= (layer0_outputs(4515)) and not (layer0_outputs(2968));
    outputs(2575) <= not(layer0_outputs(2122));
    outputs(2576) <= layer0_outputs(4316);
    outputs(2577) <= (layer0_outputs(3663)) and not (layer0_outputs(3256));
    outputs(2578) <= not((layer0_outputs(2668)) or (layer0_outputs(6363)));
    outputs(2579) <= not((layer0_outputs(6783)) and (layer0_outputs(6227)));
    outputs(2580) <= layer0_outputs(3487);
    outputs(2581) <= (layer0_outputs(2434)) and (layer0_outputs(4829));
    outputs(2582) <= (layer0_outputs(2433)) and (layer0_outputs(1971));
    outputs(2583) <= layer0_outputs(6297);
    outputs(2584) <= layer0_outputs(5464);
    outputs(2585) <= not(layer0_outputs(339));
    outputs(2586) <= (layer0_outputs(6543)) and (layer0_outputs(4194));
    outputs(2587) <= (layer0_outputs(507)) and not (layer0_outputs(103));
    outputs(2588) <= not((layer0_outputs(5293)) or (layer0_outputs(7231)));
    outputs(2589) <= (layer0_outputs(7591)) or (layer0_outputs(3634));
    outputs(2590) <= (layer0_outputs(2753)) and not (layer0_outputs(5786));
    outputs(2591) <= layer0_outputs(5798);
    outputs(2592) <= not(layer0_outputs(1649));
    outputs(2593) <= (layer0_outputs(5930)) and (layer0_outputs(5060));
    outputs(2594) <= not((layer0_outputs(2464)) xor (layer0_outputs(7468)));
    outputs(2595) <= (layer0_outputs(3176)) and not (layer0_outputs(7195));
    outputs(2596) <= not(layer0_outputs(1407));
    outputs(2597) <= (layer0_outputs(4886)) xor (layer0_outputs(4855));
    outputs(2598) <= layer0_outputs(4953);
    outputs(2599) <= not(layer0_outputs(6260));
    outputs(2600) <= (layer0_outputs(3968)) and not (layer0_outputs(5827));
    outputs(2601) <= not((layer0_outputs(6334)) xor (layer0_outputs(6795)));
    outputs(2602) <= (layer0_outputs(3967)) and not (layer0_outputs(758));
    outputs(2603) <= layer0_outputs(6002);
    outputs(2604) <= not(layer0_outputs(2501));
    outputs(2605) <= not(layer0_outputs(3142));
    outputs(2606) <= not(layer0_outputs(950));
    outputs(2607) <= (layer0_outputs(4617)) xor (layer0_outputs(605));
    outputs(2608) <= (layer0_outputs(7581)) and not (layer0_outputs(4541));
    outputs(2609) <= layer0_outputs(3964);
    outputs(2610) <= not(layer0_outputs(3026));
    outputs(2611) <= not(layer0_outputs(3036));
    outputs(2612) <= not(layer0_outputs(282));
    outputs(2613) <= layer0_outputs(6712);
    outputs(2614) <= layer0_outputs(2514);
    outputs(2615) <= layer0_outputs(2404);
    outputs(2616) <= layer0_outputs(3610);
    outputs(2617) <= layer0_outputs(5847);
    outputs(2618) <= not((layer0_outputs(3962)) xor (layer0_outputs(7247)));
    outputs(2619) <= (layer0_outputs(588)) and not (layer0_outputs(6735));
    outputs(2620) <= layer0_outputs(5576);
    outputs(2621) <= not((layer0_outputs(1612)) xor (layer0_outputs(3330)));
    outputs(2622) <= not(layer0_outputs(6690));
    outputs(2623) <= not(layer0_outputs(3108));
    outputs(2624) <= layer0_outputs(6466);
    outputs(2625) <= not(layer0_outputs(2237));
    outputs(2626) <= not((layer0_outputs(2881)) and (layer0_outputs(5313)));
    outputs(2627) <= not(layer0_outputs(3858));
    outputs(2628) <= (layer0_outputs(5158)) and not (layer0_outputs(3211));
    outputs(2629) <= layer0_outputs(1310);
    outputs(2630) <= (layer0_outputs(4379)) or (layer0_outputs(6256));
    outputs(2631) <= not(layer0_outputs(4837));
    outputs(2632) <= not(layer0_outputs(6883)) or (layer0_outputs(5291));
    outputs(2633) <= not((layer0_outputs(33)) xor (layer0_outputs(1191)));
    outputs(2634) <= (layer0_outputs(2972)) xor (layer0_outputs(6804));
    outputs(2635) <= not((layer0_outputs(814)) xor (layer0_outputs(3726)));
    outputs(2636) <= (layer0_outputs(1273)) or (layer0_outputs(2383));
    outputs(2637) <= (layer0_outputs(2051)) xor (layer0_outputs(6852));
    outputs(2638) <= (layer0_outputs(2654)) xor (layer0_outputs(2010));
    outputs(2639) <= not(layer0_outputs(4448));
    outputs(2640) <= layer0_outputs(3559);
    outputs(2641) <= layer0_outputs(3892);
    outputs(2642) <= not(layer0_outputs(1734)) or (layer0_outputs(4546));
    outputs(2643) <= layer0_outputs(2945);
    outputs(2644) <= not(layer0_outputs(5068)) or (layer0_outputs(2953));
    outputs(2645) <= layer0_outputs(3222);
    outputs(2646) <= (layer0_outputs(334)) and not (layer0_outputs(4325));
    outputs(2647) <= (layer0_outputs(3071)) and (layer0_outputs(404));
    outputs(2648) <= layer0_outputs(6143);
    outputs(2649) <= not((layer0_outputs(599)) xor (layer0_outputs(4503)));
    outputs(2650) <= not((layer0_outputs(6881)) xor (layer0_outputs(4013)));
    outputs(2651) <= (layer0_outputs(1177)) and not (layer0_outputs(1153));
    outputs(2652) <= layer0_outputs(6800);
    outputs(2653) <= (layer0_outputs(1795)) xor (layer0_outputs(5868));
    outputs(2654) <= not((layer0_outputs(7154)) xor (layer0_outputs(28)));
    outputs(2655) <= not((layer0_outputs(3945)) or (layer0_outputs(1292)));
    outputs(2656) <= (layer0_outputs(1526)) and not (layer0_outputs(1949));
    outputs(2657) <= (layer0_outputs(611)) and (layer0_outputs(3589));
    outputs(2658) <= (layer0_outputs(5386)) and (layer0_outputs(4563));
    outputs(2659) <= layer0_outputs(6799);
    outputs(2660) <= not(layer0_outputs(501));
    outputs(2661) <= layer0_outputs(6688);
    outputs(2662) <= layer0_outputs(5097);
    outputs(2663) <= (layer0_outputs(7386)) and (layer0_outputs(2179));
    outputs(2664) <= layer0_outputs(5255);
    outputs(2665) <= not(layer0_outputs(3021));
    outputs(2666) <= not((layer0_outputs(3413)) xor (layer0_outputs(1433)));
    outputs(2667) <= not(layer0_outputs(5629));
    outputs(2668) <= not(layer0_outputs(3737));
    outputs(2669) <= not((layer0_outputs(1467)) xor (layer0_outputs(7258)));
    outputs(2670) <= layer0_outputs(564);
    outputs(2671) <= not(layer0_outputs(2995));
    outputs(2672) <= not(layer0_outputs(6879));
    outputs(2673) <= not(layer0_outputs(4080));
    outputs(2674) <= (layer0_outputs(2290)) and (layer0_outputs(4250));
    outputs(2675) <= layer0_outputs(3823);
    outputs(2676) <= not(layer0_outputs(3573));
    outputs(2677) <= layer0_outputs(1422);
    outputs(2678) <= layer0_outputs(4815);
    outputs(2679) <= not(layer0_outputs(3878));
    outputs(2680) <= (layer0_outputs(3765)) and not (layer0_outputs(6252));
    outputs(2681) <= not((layer0_outputs(1556)) xor (layer0_outputs(2527)));
    outputs(2682) <= not(layer0_outputs(5563)) or (layer0_outputs(3984));
    outputs(2683) <= not(layer0_outputs(1544));
    outputs(2684) <= not(layer0_outputs(2574));
    outputs(2685) <= (layer0_outputs(821)) and (layer0_outputs(1943));
    outputs(2686) <= not((layer0_outputs(6805)) and (layer0_outputs(3080)));
    outputs(2687) <= not(layer0_outputs(1848));
    outputs(2688) <= not(layer0_outputs(2964));
    outputs(2689) <= not((layer0_outputs(2465)) and (layer0_outputs(3277)));
    outputs(2690) <= (layer0_outputs(3597)) or (layer0_outputs(3917));
    outputs(2691) <= not((layer0_outputs(4757)) or (layer0_outputs(6858)));
    outputs(2692) <= layer0_outputs(1775);
    outputs(2693) <= (layer0_outputs(1534)) xor (layer0_outputs(7069));
    outputs(2694) <= layer0_outputs(2670);
    outputs(2695) <= (layer0_outputs(4853)) or (layer0_outputs(4215));
    outputs(2696) <= not((layer0_outputs(4119)) xor (layer0_outputs(3026)));
    outputs(2697) <= not(layer0_outputs(7266)) or (layer0_outputs(4335));
    outputs(2698) <= not(layer0_outputs(5517)) or (layer0_outputs(7446));
    outputs(2699) <= (layer0_outputs(4933)) and (layer0_outputs(227));
    outputs(2700) <= not(layer0_outputs(4873));
    outputs(2701) <= not(layer0_outputs(1972));
    outputs(2702) <= not((layer0_outputs(5675)) or (layer0_outputs(4868)));
    outputs(2703) <= not((layer0_outputs(6173)) or (layer0_outputs(4084)));
    outputs(2704) <= (layer0_outputs(3543)) and not (layer0_outputs(3759));
    outputs(2705) <= layer0_outputs(7661);
    outputs(2706) <= layer0_outputs(6397);
    outputs(2707) <= not(layer0_outputs(1725));
    outputs(2708) <= not(layer0_outputs(2107));
    outputs(2709) <= not((layer0_outputs(5800)) xor (layer0_outputs(6888)));
    outputs(2710) <= not(layer0_outputs(710));
    outputs(2711) <= not((layer0_outputs(335)) xor (layer0_outputs(1114)));
    outputs(2712) <= not(layer0_outputs(505));
    outputs(2713) <= not((layer0_outputs(449)) xor (layer0_outputs(231)));
    outputs(2714) <= layer0_outputs(799);
    outputs(2715) <= (layer0_outputs(628)) and (layer0_outputs(4815));
    outputs(2716) <= (layer0_outputs(6451)) and (layer0_outputs(5861));
    outputs(2717) <= (layer0_outputs(102)) xor (layer0_outputs(92));
    outputs(2718) <= (layer0_outputs(1648)) and not (layer0_outputs(2734));
    outputs(2719) <= not(layer0_outputs(2809));
    outputs(2720) <= (layer0_outputs(7049)) and not (layer0_outputs(1079));
    outputs(2721) <= layer0_outputs(5172);
    outputs(2722) <= not(layer0_outputs(5745));
    outputs(2723) <= not(layer0_outputs(7556));
    outputs(2724) <= layer0_outputs(5141);
    outputs(2725) <= (layer0_outputs(1234)) xor (layer0_outputs(5459));
    outputs(2726) <= (layer0_outputs(1211)) xor (layer0_outputs(2263));
    outputs(2727) <= not(layer0_outputs(1511)) or (layer0_outputs(851));
    outputs(2728) <= not(layer0_outputs(2589)) or (layer0_outputs(370));
    outputs(2729) <= layer0_outputs(3182);
    outputs(2730) <= (layer0_outputs(7628)) xor (layer0_outputs(2854));
    outputs(2731) <= layer0_outputs(5234);
    outputs(2732) <= not(layer0_outputs(3850));
    outputs(2733) <= (layer0_outputs(6834)) and not (layer0_outputs(663));
    outputs(2734) <= layer0_outputs(1229);
    outputs(2735) <= not(layer0_outputs(2147));
    outputs(2736) <= not(layer0_outputs(1110)) or (layer0_outputs(4331));
    outputs(2737) <= (layer0_outputs(3176)) and not (layer0_outputs(2877));
    outputs(2738) <= (layer0_outputs(4178)) xor (layer0_outputs(4378));
    outputs(2739) <= not(layer0_outputs(3921));
    outputs(2740) <= layer0_outputs(4335);
    outputs(2741) <= (layer0_outputs(1322)) xor (layer0_outputs(5383));
    outputs(2742) <= layer0_outputs(5407);
    outputs(2743) <= layer0_outputs(7611);
    outputs(2744) <= layer0_outputs(6672);
    outputs(2745) <= (layer0_outputs(4747)) xor (layer0_outputs(4301));
    outputs(2746) <= not(layer0_outputs(2033));
    outputs(2747) <= not(layer0_outputs(7236));
    outputs(2748) <= not(layer0_outputs(5499));
    outputs(2749) <= not(layer0_outputs(6));
    outputs(2750) <= not(layer0_outputs(959)) or (layer0_outputs(3610));
    outputs(2751) <= layer0_outputs(6566);
    outputs(2752) <= layer0_outputs(209);
    outputs(2753) <= (layer0_outputs(1385)) or (layer0_outputs(696));
    outputs(2754) <= not(layer0_outputs(7241));
    outputs(2755) <= not((layer0_outputs(1470)) or (layer0_outputs(1826)));
    outputs(2756) <= not((layer0_outputs(5308)) or (layer0_outputs(1535)));
    outputs(2757) <= not(layer0_outputs(5215));
    outputs(2758) <= not(layer0_outputs(4734)) or (layer0_outputs(7430));
    outputs(2759) <= not(layer0_outputs(6577)) or (layer0_outputs(7644));
    outputs(2760) <= not((layer0_outputs(6175)) or (layer0_outputs(3603)));
    outputs(2761) <= not(layer0_outputs(5516));
    outputs(2762) <= layer0_outputs(1334);
    outputs(2763) <= (layer0_outputs(6755)) and (layer0_outputs(4096));
    outputs(2764) <= not(layer0_outputs(5025)) or (layer0_outputs(7485));
    outputs(2765) <= layer0_outputs(3798);
    outputs(2766) <= not((layer0_outputs(7005)) and (layer0_outputs(6334)));
    outputs(2767) <= (layer0_outputs(165)) and not (layer0_outputs(1810));
    outputs(2768) <= not((layer0_outputs(4234)) and (layer0_outputs(7253)));
    outputs(2769) <= (layer0_outputs(945)) and not (layer0_outputs(4605));
    outputs(2770) <= layer0_outputs(230);
    outputs(2771) <= (layer0_outputs(3875)) xor (layer0_outputs(1595));
    outputs(2772) <= not((layer0_outputs(3166)) xor (layer0_outputs(5947)));
    outputs(2773) <= not(layer0_outputs(4582));
    outputs(2774) <= layer0_outputs(1962);
    outputs(2775) <= not(layer0_outputs(2117));
    outputs(2776) <= not((layer0_outputs(526)) and (layer0_outputs(3755)));
    outputs(2777) <= not(layer0_outputs(5053));
    outputs(2778) <= (layer0_outputs(6624)) xor (layer0_outputs(3907));
    outputs(2779) <= (layer0_outputs(1824)) xor (layer0_outputs(3053));
    outputs(2780) <= layer0_outputs(1740);
    outputs(2781) <= layer0_outputs(2096);
    outputs(2782) <= layer0_outputs(611);
    outputs(2783) <= not(layer0_outputs(3183)) or (layer0_outputs(6143));
    outputs(2784) <= layer0_outputs(5140);
    outputs(2785) <= not((layer0_outputs(2846)) xor (layer0_outputs(3649)));
    outputs(2786) <= layer0_outputs(4233);
    outputs(2787) <= not(layer0_outputs(1837)) or (layer0_outputs(2705));
    outputs(2788) <= (layer0_outputs(6709)) xor (layer0_outputs(3420));
    outputs(2789) <= layer0_outputs(1457);
    outputs(2790) <= not(layer0_outputs(2269)) or (layer0_outputs(1577));
    outputs(2791) <= not((layer0_outputs(4135)) xor (layer0_outputs(1018)));
    outputs(2792) <= not(layer0_outputs(3581));
    outputs(2793) <= layer0_outputs(4211);
    outputs(2794) <= not(layer0_outputs(182));
    outputs(2795) <= layer0_outputs(7586);
    outputs(2796) <= not((layer0_outputs(7122)) xor (layer0_outputs(5361)));
    outputs(2797) <= not(layer0_outputs(548));
    outputs(2798) <= layer0_outputs(6187);
    outputs(2799) <= not(layer0_outputs(4773));
    outputs(2800) <= (layer0_outputs(3074)) and not (layer0_outputs(2152));
    outputs(2801) <= (layer0_outputs(2949)) xor (layer0_outputs(866));
    outputs(2802) <= (layer0_outputs(531)) and not (layer0_outputs(6819));
    outputs(2803) <= (layer0_outputs(3306)) and (layer0_outputs(2544));
    outputs(2804) <= layer0_outputs(1378);
    outputs(2805) <= layer0_outputs(5660);
    outputs(2806) <= (layer0_outputs(317)) and not (layer0_outputs(2802));
    outputs(2807) <= (layer0_outputs(914)) xor (layer0_outputs(5680));
    outputs(2808) <= not(layer0_outputs(3737));
    outputs(2809) <= layer0_outputs(3729);
    outputs(2810) <= layer0_outputs(4437);
    outputs(2811) <= (layer0_outputs(7345)) and not (layer0_outputs(4337));
    outputs(2812) <= (layer0_outputs(7084)) and not (layer0_outputs(3358));
    outputs(2813) <= not((layer0_outputs(3625)) or (layer0_outputs(5596)));
    outputs(2814) <= layer0_outputs(3804);
    outputs(2815) <= (layer0_outputs(5009)) and not (layer0_outputs(5489));
    outputs(2816) <= (layer0_outputs(6907)) and not (layer0_outputs(3581));
    outputs(2817) <= (layer0_outputs(6032)) and not (layer0_outputs(1390));
    outputs(2818) <= (layer0_outputs(5674)) xor (layer0_outputs(6567));
    outputs(2819) <= not(layer0_outputs(2696));
    outputs(2820) <= not((layer0_outputs(6651)) and (layer0_outputs(4159)));
    outputs(2821) <= (layer0_outputs(4302)) and not (layer0_outputs(3291));
    outputs(2822) <= not(layer0_outputs(4887));
    outputs(2823) <= layer0_outputs(1893);
    outputs(2824) <= layer0_outputs(1648);
    outputs(2825) <= layer0_outputs(1979);
    outputs(2826) <= (layer0_outputs(7489)) and (layer0_outputs(3876));
    outputs(2827) <= not(layer0_outputs(1140));
    outputs(2828) <= not((layer0_outputs(6469)) xor (layer0_outputs(7428)));
    outputs(2829) <= (layer0_outputs(3754)) and not (layer0_outputs(1002));
    outputs(2830) <= layer0_outputs(5082);
    outputs(2831) <= layer0_outputs(7651);
    outputs(2832) <= not(layer0_outputs(2860));
    outputs(2833) <= not(layer0_outputs(3657));
    outputs(2834) <= (layer0_outputs(304)) xor (layer0_outputs(910));
    outputs(2835) <= not(layer0_outputs(4709));
    outputs(2836) <= not((layer0_outputs(4854)) or (layer0_outputs(2027)));
    outputs(2837) <= not(layer0_outputs(3450));
    outputs(2838) <= layer0_outputs(1999);
    outputs(2839) <= layer0_outputs(2514);
    outputs(2840) <= (layer0_outputs(1763)) and not (layer0_outputs(5620));
    outputs(2841) <= layer0_outputs(5400);
    outputs(2842) <= not(layer0_outputs(2049));
    outputs(2843) <= layer0_outputs(6496);
    outputs(2844) <= (layer0_outputs(2174)) xor (layer0_outputs(7113));
    outputs(2845) <= layer0_outputs(2835);
    outputs(2846) <= layer0_outputs(446);
    outputs(2847) <= (layer0_outputs(4057)) and (layer0_outputs(1894));
    outputs(2848) <= not((layer0_outputs(4863)) or (layer0_outputs(491)));
    outputs(2849) <= not(layer0_outputs(2978));
    outputs(2850) <= not(layer0_outputs(5479));
    outputs(2851) <= layer0_outputs(3717);
    outputs(2852) <= (layer0_outputs(3023)) and not (layer0_outputs(6550));
    outputs(2853) <= not(layer0_outputs(6435));
    outputs(2854) <= not(layer0_outputs(369));
    outputs(2855) <= (layer0_outputs(6557)) and (layer0_outputs(2771));
    outputs(2856) <= (layer0_outputs(4761)) and (layer0_outputs(3213));
    outputs(2857) <= (layer0_outputs(5787)) and not (layer0_outputs(5286));
    outputs(2858) <= layer0_outputs(7392);
    outputs(2859) <= (layer0_outputs(5967)) and not (layer0_outputs(6050));
    outputs(2860) <= layer0_outputs(4168);
    outputs(2861) <= layer0_outputs(313);
    outputs(2862) <= (layer0_outputs(3399)) xor (layer0_outputs(6702));
    outputs(2863) <= (layer0_outputs(4972)) and not (layer0_outputs(6663));
    outputs(2864) <= (layer0_outputs(4446)) or (layer0_outputs(4255));
    outputs(2865) <= not((layer0_outputs(6901)) or (layer0_outputs(6151)));
    outputs(2866) <= not(layer0_outputs(6843));
    outputs(2867) <= not(layer0_outputs(4685));
    outputs(2868) <= not((layer0_outputs(837)) xor (layer0_outputs(2816)));
    outputs(2869) <= layer0_outputs(5792);
    outputs(2870) <= layer0_outputs(2024);
    outputs(2871) <= (layer0_outputs(1742)) xor (layer0_outputs(1249));
    outputs(2872) <= layer0_outputs(683);
    outputs(2873) <= layer0_outputs(5074);
    outputs(2874) <= not((layer0_outputs(1649)) or (layer0_outputs(5980)));
    outputs(2875) <= not((layer0_outputs(476)) and (layer0_outputs(297)));
    outputs(2876) <= not(layer0_outputs(895));
    outputs(2877) <= (layer0_outputs(4622)) and not (layer0_outputs(7036));
    outputs(2878) <= (layer0_outputs(6285)) and not (layer0_outputs(6969));
    outputs(2879) <= (layer0_outputs(554)) and not (layer0_outputs(6446));
    outputs(2880) <= layer0_outputs(671);
    outputs(2881) <= not(layer0_outputs(5422));
    outputs(2882) <= (layer0_outputs(1705)) xor (layer0_outputs(2892));
    outputs(2883) <= not(layer0_outputs(6761));
    outputs(2884) <= layer0_outputs(3017);
    outputs(2885) <= not((layer0_outputs(4695)) xor (layer0_outputs(2278)));
    outputs(2886) <= not(layer0_outputs(3475));
    outputs(2887) <= (layer0_outputs(856)) xor (layer0_outputs(4779));
    outputs(2888) <= not(layer0_outputs(4021));
    outputs(2889) <= not((layer0_outputs(7650)) xor (layer0_outputs(5408)));
    outputs(2890) <= layer0_outputs(1740);
    outputs(2891) <= (layer0_outputs(1579)) and not (layer0_outputs(2358));
    outputs(2892) <= (layer0_outputs(572)) xor (layer0_outputs(7265));
    outputs(2893) <= (layer0_outputs(3510)) or (layer0_outputs(2251));
    outputs(2894) <= (layer0_outputs(592)) and (layer0_outputs(2308));
    outputs(2895) <= layer0_outputs(3712);
    outputs(2896) <= not((layer0_outputs(5878)) and (layer0_outputs(2982)));
    outputs(2897) <= (layer0_outputs(4566)) and not (layer0_outputs(3776));
    outputs(2898) <= not(layer0_outputs(6389));
    outputs(2899) <= not((layer0_outputs(6250)) xor (layer0_outputs(19)));
    outputs(2900) <= layer0_outputs(395);
    outputs(2901) <= layer0_outputs(646);
    outputs(2902) <= not(layer0_outputs(6264));
    outputs(2903) <= (layer0_outputs(3295)) xor (layer0_outputs(1120));
    outputs(2904) <= not(layer0_outputs(2607));
    outputs(2905) <= layer0_outputs(5149);
    outputs(2906) <= (layer0_outputs(4275)) xor (layer0_outputs(4142));
    outputs(2907) <= (layer0_outputs(6703)) xor (layer0_outputs(6488));
    outputs(2908) <= (layer0_outputs(5633)) and not (layer0_outputs(3843));
    outputs(2909) <= (layer0_outputs(427)) or (layer0_outputs(2851));
    outputs(2910) <= layer0_outputs(6751);
    outputs(2911) <= not(layer0_outputs(7103));
    outputs(2912) <= not(layer0_outputs(4791));
    outputs(2913) <= (layer0_outputs(1346)) and not (layer0_outputs(6759));
    outputs(2914) <= not(layer0_outputs(5697)) or (layer0_outputs(1547));
    outputs(2915) <= (layer0_outputs(770)) and not (layer0_outputs(3320));
    outputs(2916) <= (layer0_outputs(2516)) and (layer0_outputs(5319));
    outputs(2917) <= (layer0_outputs(749)) and not (layer0_outputs(5954));
    outputs(2918) <= (layer0_outputs(291)) xor (layer0_outputs(3646));
    outputs(2919) <= (layer0_outputs(2476)) and not (layer0_outputs(3555));
    outputs(2920) <= (layer0_outputs(1328)) or (layer0_outputs(3344));
    outputs(2921) <= not(layer0_outputs(164)) or (layer0_outputs(3207));
    outputs(2922) <= not((layer0_outputs(6922)) and (layer0_outputs(1329)));
    outputs(2923) <= not(layer0_outputs(6727));
    outputs(2924) <= layer0_outputs(4060);
    outputs(2925) <= layer0_outputs(1455);
    outputs(2926) <= not(layer0_outputs(3727));
    outputs(2927) <= not(layer0_outputs(2286));
    outputs(2928) <= not((layer0_outputs(2478)) xor (layer0_outputs(1640)));
    outputs(2929) <= (layer0_outputs(532)) and not (layer0_outputs(1631));
    outputs(2930) <= not(layer0_outputs(5648));
    outputs(2931) <= not((layer0_outputs(4734)) or (layer0_outputs(2553)));
    outputs(2932) <= (layer0_outputs(1683)) and not (layer0_outputs(2590));
    outputs(2933) <= not(layer0_outputs(3131));
    outputs(2934) <= not(layer0_outputs(397)) or (layer0_outputs(7132));
    outputs(2935) <= layer0_outputs(6828);
    outputs(2936) <= layer0_outputs(4199);
    outputs(2937) <= (layer0_outputs(1043)) or (layer0_outputs(7319));
    outputs(2938) <= (layer0_outputs(5195)) and (layer0_outputs(1073));
    outputs(2939) <= layer0_outputs(2070);
    outputs(2940) <= (layer0_outputs(96)) and not (layer0_outputs(161));
    outputs(2941) <= not(layer0_outputs(6058));
    outputs(2942) <= not((layer0_outputs(2090)) or (layer0_outputs(6781)));
    outputs(2943) <= layer0_outputs(7376);
    outputs(2944) <= layer0_outputs(5603);
    outputs(2945) <= layer0_outputs(6671);
    outputs(2946) <= not(layer0_outputs(4505));
    outputs(2947) <= not(layer0_outputs(6210));
    outputs(2948) <= (layer0_outputs(2715)) xor (layer0_outputs(2169));
    outputs(2949) <= not((layer0_outputs(6922)) or (layer0_outputs(886)));
    outputs(2950) <= not(layer0_outputs(7219));
    outputs(2951) <= layer0_outputs(1009);
    outputs(2952) <= not(layer0_outputs(1397));
    outputs(2953) <= layer0_outputs(842);
    outputs(2954) <= (layer0_outputs(3182)) or (layer0_outputs(7307));
    outputs(2955) <= (layer0_outputs(5082)) and not (layer0_outputs(3562));
    outputs(2956) <= (layer0_outputs(2868)) xor (layer0_outputs(22));
    outputs(2957) <= not(layer0_outputs(182));
    outputs(2958) <= (layer0_outputs(3972)) xor (layer0_outputs(4680));
    outputs(2959) <= not(layer0_outputs(6964)) or (layer0_outputs(3394));
    outputs(2960) <= not((layer0_outputs(1289)) or (layer0_outputs(7387)));
    outputs(2961) <= not(layer0_outputs(6295)) or (layer0_outputs(3194));
    outputs(2962) <= (layer0_outputs(3449)) and not (layer0_outputs(2312));
    outputs(2963) <= (layer0_outputs(3167)) xor (layer0_outputs(3809));
    outputs(2964) <= (layer0_outputs(3391)) and (layer0_outputs(5152));
    outputs(2965) <= (layer0_outputs(7621)) and (layer0_outputs(6791));
    outputs(2966) <= (layer0_outputs(7268)) and (layer0_outputs(2410));
    outputs(2967) <= layer0_outputs(6128);
    outputs(2968) <= not(layer0_outputs(1882));
    outputs(2969) <= not(layer0_outputs(6331));
    outputs(2970) <= not((layer0_outputs(93)) xor (layer0_outputs(23)));
    outputs(2971) <= (layer0_outputs(1610)) and (layer0_outputs(929));
    outputs(2972) <= not((layer0_outputs(7354)) xor (layer0_outputs(2011)));
    outputs(2973) <= not(layer0_outputs(1858));
    outputs(2974) <= not((layer0_outputs(5468)) or (layer0_outputs(2224)));
    outputs(2975) <= not((layer0_outputs(737)) or (layer0_outputs(6639)));
    outputs(2976) <= not(layer0_outputs(4766));
    outputs(2977) <= (layer0_outputs(714)) xor (layer0_outputs(3117));
    outputs(2978) <= not((layer0_outputs(3090)) xor (layer0_outputs(3811)));
    outputs(2979) <= not((layer0_outputs(6504)) xor (layer0_outputs(4217)));
    outputs(2980) <= not((layer0_outputs(2466)) xor (layer0_outputs(7621)));
    outputs(2981) <= (layer0_outputs(2794)) and not (layer0_outputs(7553));
    outputs(2982) <= not(layer0_outputs(6489));
    outputs(2983) <= layer0_outputs(7202);
    outputs(2984) <= layer0_outputs(4257);
    outputs(2985) <= not(layer0_outputs(6569));
    outputs(2986) <= not(layer0_outputs(4492));
    outputs(2987) <= not((layer0_outputs(793)) or (layer0_outputs(4217)));
    outputs(2988) <= layer0_outputs(615);
    outputs(2989) <= layer0_outputs(5173);
    outputs(2990) <= not(layer0_outputs(6846));
    outputs(2991) <= layer0_outputs(1313);
    outputs(2992) <= not((layer0_outputs(7313)) or (layer0_outputs(2120)));
    outputs(2993) <= (layer0_outputs(7088)) xor (layer0_outputs(6321));
    outputs(2994) <= not((layer0_outputs(4903)) xor (layer0_outputs(6829)));
    outputs(2995) <= not(layer0_outputs(2895));
    outputs(2996) <= not((layer0_outputs(5316)) and (layer0_outputs(3228)));
    outputs(2997) <= (layer0_outputs(4083)) and not (layer0_outputs(551));
    outputs(2998) <= layer0_outputs(747);
    outputs(2999) <= (layer0_outputs(5725)) and (layer0_outputs(6582));
    outputs(3000) <= not(layer0_outputs(4181));
    outputs(3001) <= (layer0_outputs(7675)) or (layer0_outputs(1681));
    outputs(3002) <= (layer0_outputs(1754)) and (layer0_outputs(6711));
    outputs(3003) <= layer0_outputs(2265);
    outputs(3004) <= not(layer0_outputs(6116));
    outputs(3005) <= (layer0_outputs(382)) and (layer0_outputs(7603));
    outputs(3006) <= not(layer0_outputs(6416));
    outputs(3007) <= (layer0_outputs(3908)) xor (layer0_outputs(4499));
    outputs(3008) <= not((layer0_outputs(593)) or (layer0_outputs(1206)));
    outputs(3009) <= layer0_outputs(5152);
    outputs(3010) <= not(layer0_outputs(3956));
    outputs(3011) <= layer0_outputs(4476);
    outputs(3012) <= (layer0_outputs(7388)) and (layer0_outputs(4994));
    outputs(3013) <= (layer0_outputs(274)) xor (layer0_outputs(5118));
    outputs(3014) <= layer0_outputs(2083);
    outputs(3015) <= (layer0_outputs(2349)) and not (layer0_outputs(6635));
    outputs(3016) <= not(layer0_outputs(7524));
    outputs(3017) <= (layer0_outputs(5382)) and not (layer0_outputs(1881));
    outputs(3018) <= (layer0_outputs(4514)) and (layer0_outputs(1787));
    outputs(3019) <= (layer0_outputs(601)) xor (layer0_outputs(6794));
    outputs(3020) <= not(layer0_outputs(654));
    outputs(3021) <= not((layer0_outputs(2378)) or (layer0_outputs(1492)));
    outputs(3022) <= not(layer0_outputs(3541)) or (layer0_outputs(2350));
    outputs(3023) <= (layer0_outputs(6261)) and (layer0_outputs(1874));
    outputs(3024) <= not(layer0_outputs(1478)) or (layer0_outputs(6685));
    outputs(3025) <= layer0_outputs(3742);
    outputs(3026) <= not(layer0_outputs(1083));
    outputs(3027) <= layer0_outputs(5270);
    outputs(3028) <= (layer0_outputs(371)) and (layer0_outputs(4923));
    outputs(3029) <= layer0_outputs(3225);
    outputs(3030) <= layer0_outputs(5138);
    outputs(3031) <= not(layer0_outputs(620));
    outputs(3032) <= not(layer0_outputs(5224));
    outputs(3033) <= (layer0_outputs(4899)) xor (layer0_outputs(5554));
    outputs(3034) <= layer0_outputs(138);
    outputs(3035) <= (layer0_outputs(18)) and (layer0_outputs(1538));
    outputs(3036) <= (layer0_outputs(3164)) and not (layer0_outputs(6236));
    outputs(3037) <= layer0_outputs(3554);
    outputs(3038) <= not(layer0_outputs(7314));
    outputs(3039) <= (layer0_outputs(7190)) xor (layer0_outputs(7339));
    outputs(3040) <= not(layer0_outputs(7574)) or (layer0_outputs(1776));
    outputs(3041) <= layer0_outputs(6527);
    outputs(3042) <= layer0_outputs(5673);
    outputs(3043) <= layer0_outputs(1735);
    outputs(3044) <= layer0_outputs(2203);
    outputs(3045) <= not(layer0_outputs(7125));
    outputs(3046) <= (layer0_outputs(1149)) xor (layer0_outputs(2287));
    outputs(3047) <= not(layer0_outputs(4632)) or (layer0_outputs(1149));
    outputs(3048) <= (layer0_outputs(5485)) and not (layer0_outputs(284));
    outputs(3049) <= not(layer0_outputs(3881));
    outputs(3050) <= not(layer0_outputs(3278));
    outputs(3051) <= layer0_outputs(920);
    outputs(3052) <= (layer0_outputs(761)) and (layer0_outputs(319));
    outputs(3053) <= not((layer0_outputs(1733)) or (layer0_outputs(5587)));
    outputs(3054) <= not((layer0_outputs(4670)) or (layer0_outputs(3602)));
    outputs(3055) <= layer0_outputs(6074);
    outputs(3056) <= not((layer0_outputs(2708)) xor (layer0_outputs(6044)));
    outputs(3057) <= not(layer0_outputs(249));
    outputs(3058) <= not(layer0_outputs(2491));
    outputs(3059) <= layer0_outputs(7543);
    outputs(3060) <= (layer0_outputs(1550)) and (layer0_outputs(317));
    outputs(3061) <= layer0_outputs(5245);
    outputs(3062) <= not(layer0_outputs(3011));
    outputs(3063) <= not((layer0_outputs(3318)) or (layer0_outputs(2765)));
    outputs(3064) <= not(layer0_outputs(3611)) or (layer0_outputs(2441));
    outputs(3065) <= not((layer0_outputs(3075)) xor (layer0_outputs(2458)));
    outputs(3066) <= not(layer0_outputs(771)) or (layer0_outputs(6696));
    outputs(3067) <= (layer0_outputs(5763)) xor (layer0_outputs(7449));
    outputs(3068) <= layer0_outputs(7202);
    outputs(3069) <= (layer0_outputs(4602)) and (layer0_outputs(7199));
    outputs(3070) <= not((layer0_outputs(1494)) xor (layer0_outputs(3883)));
    outputs(3071) <= not(layer0_outputs(6244));
    outputs(3072) <= not(layer0_outputs(2782));
    outputs(3073) <= (layer0_outputs(1285)) and (layer0_outputs(2844));
    outputs(3074) <= (layer0_outputs(2454)) xor (layer0_outputs(6354));
    outputs(3075) <= not(layer0_outputs(3823));
    outputs(3076) <= (layer0_outputs(3717)) or (layer0_outputs(3219));
    outputs(3077) <= not(layer0_outputs(3605));
    outputs(3078) <= not(layer0_outputs(1685));
    outputs(3079) <= not((layer0_outputs(4686)) xor (layer0_outputs(5433)));
    outputs(3080) <= (layer0_outputs(7553)) or (layer0_outputs(4007));
    outputs(3081) <= layer0_outputs(5567);
    outputs(3082) <= (layer0_outputs(6053)) or (layer0_outputs(7628));
    outputs(3083) <= (layer0_outputs(202)) and (layer0_outputs(5681));
    outputs(3084) <= not((layer0_outputs(4292)) xor (layer0_outputs(5342)));
    outputs(3085) <= not(layer0_outputs(6356)) or (layer0_outputs(3111));
    outputs(3086) <= layer0_outputs(6538);
    outputs(3087) <= (layer0_outputs(3347)) and not (layer0_outputs(5584));
    outputs(3088) <= layer0_outputs(3396);
    outputs(3089) <= layer0_outputs(4175);
    outputs(3090) <= not(layer0_outputs(4061));
    outputs(3091) <= not(layer0_outputs(1877));
    outputs(3092) <= not(layer0_outputs(5372));
    outputs(3093) <= (layer0_outputs(1599)) xor (layer0_outputs(4258));
    outputs(3094) <= not(layer0_outputs(4719)) or (layer0_outputs(7433));
    outputs(3095) <= layer0_outputs(4333);
    outputs(3096) <= layer0_outputs(224);
    outputs(3097) <= layer0_outputs(5688);
    outputs(3098) <= not(layer0_outputs(1847));
    outputs(3099) <= not(layer0_outputs(6200));
    outputs(3100) <= layer0_outputs(328);
    outputs(3101) <= layer0_outputs(805);
    outputs(3102) <= not(layer0_outputs(6600)) or (layer0_outputs(3208));
    outputs(3103) <= (layer0_outputs(3720)) xor (layer0_outputs(4116));
    outputs(3104) <= layer0_outputs(3814);
    outputs(3105) <= layer0_outputs(2767);
    outputs(3106) <= layer0_outputs(3033);
    outputs(3107) <= (layer0_outputs(4160)) and (layer0_outputs(6720));
    outputs(3108) <= (layer0_outputs(5032)) and not (layer0_outputs(7420));
    outputs(3109) <= not((layer0_outputs(475)) xor (layer0_outputs(5933)));
    outputs(3110) <= (layer0_outputs(1623)) and (layer0_outputs(1653));
    outputs(3111) <= (layer0_outputs(1293)) and not (layer0_outputs(4806));
    outputs(3112) <= (layer0_outputs(5465)) and not (layer0_outputs(5621));
    outputs(3113) <= not((layer0_outputs(6280)) xor (layer0_outputs(3913)));
    outputs(3114) <= not(layer0_outputs(4047));
    outputs(3115) <= layer0_outputs(2237);
    outputs(3116) <= not(layer0_outputs(2612));
    outputs(3117) <= layer0_outputs(3662);
    outputs(3118) <= not((layer0_outputs(3264)) and (layer0_outputs(1664)));
    outputs(3119) <= (layer0_outputs(2811)) and not (layer0_outputs(5990));
    outputs(3120) <= (layer0_outputs(6181)) and not (layer0_outputs(3753));
    outputs(3121) <= not((layer0_outputs(4930)) or (layer0_outputs(7447)));
    outputs(3122) <= not(layer0_outputs(263));
    outputs(3123) <= (layer0_outputs(4341)) and (layer0_outputs(4405));
    outputs(3124) <= not((layer0_outputs(4656)) or (layer0_outputs(529)));
    outputs(3125) <= layer0_outputs(6197);
    outputs(3126) <= layer0_outputs(6302);
    outputs(3127) <= (layer0_outputs(1319)) xor (layer0_outputs(596));
    outputs(3128) <= not(layer0_outputs(6059)) or (layer0_outputs(2757));
    outputs(3129) <= layer0_outputs(2302);
    outputs(3130) <= layer0_outputs(5250);
    outputs(3131) <= layer0_outputs(2228);
    outputs(3132) <= layer0_outputs(4317);
    outputs(3133) <= not(layer0_outputs(2094));
    outputs(3134) <= (layer0_outputs(472)) xor (layer0_outputs(6040));
    outputs(3135) <= not(layer0_outputs(2787));
    outputs(3136) <= not(layer0_outputs(2925));
    outputs(3137) <= not(layer0_outputs(2920));
    outputs(3138) <= not(layer0_outputs(6201)) or (layer0_outputs(5507));
    outputs(3139) <= layer0_outputs(5714);
    outputs(3140) <= not(layer0_outputs(6273));
    outputs(3141) <= not(layer0_outputs(1976));
    outputs(3142) <= not(layer0_outputs(7500));
    outputs(3143) <= (layer0_outputs(871)) and not (layer0_outputs(7395));
    outputs(3144) <= layer0_outputs(200);
    outputs(3145) <= not((layer0_outputs(1793)) xor (layer0_outputs(1849)));
    outputs(3146) <= layer0_outputs(2308);
    outputs(3147) <= (layer0_outputs(4972)) xor (layer0_outputs(1808));
    outputs(3148) <= not((layer0_outputs(2631)) and (layer0_outputs(1136)));
    outputs(3149) <= (layer0_outputs(7056)) and not (layer0_outputs(2678));
    outputs(3150) <= layer0_outputs(2326);
    outputs(3151) <= layer0_outputs(3102);
    outputs(3152) <= (layer0_outputs(7613)) and not (layer0_outputs(6795));
    outputs(3153) <= not((layer0_outputs(5553)) or (layer0_outputs(4749)));
    outputs(3154) <= not((layer0_outputs(955)) xor (layer0_outputs(2541)));
    outputs(3155) <= (layer0_outputs(7527)) and not (layer0_outputs(5188));
    outputs(3156) <= not((layer0_outputs(7391)) xor (layer0_outputs(3907)));
    outputs(3157) <= layer0_outputs(6062);
    outputs(3158) <= not(layer0_outputs(6349)) or (layer0_outputs(3719));
    outputs(3159) <= not(layer0_outputs(2038));
    outputs(3160) <= (layer0_outputs(5517)) and (layer0_outputs(6762));
    outputs(3161) <= not(layer0_outputs(4583));
    outputs(3162) <= layer0_outputs(4916);
    outputs(3163) <= not(layer0_outputs(3748));
    outputs(3164) <= not((layer0_outputs(2166)) xor (layer0_outputs(2518)));
    outputs(3165) <= layer0_outputs(2306);
    outputs(3166) <= not(layer0_outputs(1247));
    outputs(3167) <= not(layer0_outputs(6721));
    outputs(3168) <= not(layer0_outputs(4802));
    outputs(3169) <= not((layer0_outputs(5831)) or (layer0_outputs(2532)));
    outputs(3170) <= not(layer0_outputs(3503));
    outputs(3171) <= not(layer0_outputs(199));
    outputs(3172) <= (layer0_outputs(2376)) and not (layer0_outputs(6740));
    outputs(3173) <= (layer0_outputs(7155)) and not (layer0_outputs(1258));
    outputs(3174) <= layer0_outputs(3154);
    outputs(3175) <= (layer0_outputs(5948)) and not (layer0_outputs(1795));
    outputs(3176) <= (layer0_outputs(7597)) and not (layer0_outputs(5116));
    outputs(3177) <= (layer0_outputs(4140)) xor (layer0_outputs(4746));
    outputs(3178) <= layer0_outputs(5290);
    outputs(3179) <= not((layer0_outputs(6625)) and (layer0_outputs(2469)));
    outputs(3180) <= (layer0_outputs(5618)) and (layer0_outputs(7534));
    outputs(3181) <= (layer0_outputs(7100)) or (layer0_outputs(2201));
    outputs(3182) <= (layer0_outputs(2689)) or (layer0_outputs(692));
    outputs(3183) <= (layer0_outputs(5528)) xor (layer0_outputs(5509));
    outputs(3184) <= not((layer0_outputs(1316)) xor (layer0_outputs(6801)));
    outputs(3185) <= not(layer0_outputs(3994)) or (layer0_outputs(4978));
    outputs(3186) <= not((layer0_outputs(74)) or (layer0_outputs(222)));
    outputs(3187) <= (layer0_outputs(6496)) and not (layer0_outputs(3768));
    outputs(3188) <= (layer0_outputs(3165)) xor (layer0_outputs(4222));
    outputs(3189) <= not(layer0_outputs(2764));
    outputs(3190) <= not(layer0_outputs(2387));
    outputs(3191) <= layer0_outputs(928);
    outputs(3192) <= (layer0_outputs(6166)) xor (layer0_outputs(7022));
    outputs(3193) <= layer0_outputs(5727);
    outputs(3194) <= not((layer0_outputs(2880)) or (layer0_outputs(4613)));
    outputs(3195) <= not((layer0_outputs(4058)) xor (layer0_outputs(1250)));
    outputs(3196) <= not((layer0_outputs(5621)) xor (layer0_outputs(1290)));
    outputs(3197) <= layer0_outputs(5997);
    outputs(3198) <= not((layer0_outputs(4553)) or (layer0_outputs(2835)));
    outputs(3199) <= not(layer0_outputs(4094));
    outputs(3200) <= (layer0_outputs(2628)) and (layer0_outputs(4321));
    outputs(3201) <= layer0_outputs(3707);
    outputs(3202) <= layer0_outputs(3629);
    outputs(3203) <= (layer0_outputs(3491)) xor (layer0_outputs(203));
    outputs(3204) <= (layer0_outputs(6810)) and not (layer0_outputs(4182));
    outputs(3205) <= layer0_outputs(642);
    outputs(3206) <= (layer0_outputs(2628)) and not (layer0_outputs(7443));
    outputs(3207) <= layer0_outputs(3238);
    outputs(3208) <= layer0_outputs(2645);
    outputs(3209) <= layer0_outputs(3660);
    outputs(3210) <= (layer0_outputs(5622)) xor (layer0_outputs(6571));
    outputs(3211) <= (layer0_outputs(3992)) xor (layer0_outputs(3539));
    outputs(3212) <= not(layer0_outputs(4791));
    outputs(3213) <= (layer0_outputs(1661)) and not (layer0_outputs(6499));
    outputs(3214) <= not((layer0_outputs(522)) and (layer0_outputs(6726)));
    outputs(3215) <= (layer0_outputs(1360)) and not (layer0_outputs(1419));
    outputs(3216) <= not(layer0_outputs(3661));
    outputs(3217) <= (layer0_outputs(7205)) xor (layer0_outputs(5084));
    outputs(3218) <= not(layer0_outputs(3751));
    outputs(3219) <= not((layer0_outputs(4134)) and (layer0_outputs(4879)));
    outputs(3220) <= (layer0_outputs(683)) xor (layer0_outputs(4288));
    outputs(3221) <= layer0_outputs(1613);
    outputs(3222) <= layer0_outputs(6771);
    outputs(3223) <= layer0_outputs(95);
    outputs(3224) <= not(layer0_outputs(2818));
    outputs(3225) <= not(layer0_outputs(5804)) or (layer0_outputs(7492));
    outputs(3226) <= not(layer0_outputs(7101));
    outputs(3227) <= not((layer0_outputs(5340)) xor (layer0_outputs(4735)));
    outputs(3228) <= not(layer0_outputs(5995)) or (layer0_outputs(2172));
    outputs(3229) <= not(layer0_outputs(6835));
    outputs(3230) <= (layer0_outputs(6340)) and not (layer0_outputs(6151));
    outputs(3231) <= (layer0_outputs(1602)) and not (layer0_outputs(3919));
    outputs(3232) <= not(layer0_outputs(7061));
    outputs(3233) <= not((layer0_outputs(2987)) xor (layer0_outputs(745)));
    outputs(3234) <= not((layer0_outputs(3195)) xor (layer0_outputs(5171)));
    outputs(3235) <= layer0_outputs(471);
    outputs(3236) <= (layer0_outputs(2134)) and (layer0_outputs(2742));
    outputs(3237) <= (layer0_outputs(4760)) xor (layer0_outputs(1494));
    outputs(3238) <= (layer0_outputs(1318)) and not (layer0_outputs(5065));
    outputs(3239) <= (layer0_outputs(1978)) and (layer0_outputs(3108));
    outputs(3240) <= layer0_outputs(5051);
    outputs(3241) <= not((layer0_outputs(6540)) and (layer0_outputs(4800)));
    outputs(3242) <= not(layer0_outputs(3625));
    outputs(3243) <= (layer0_outputs(323)) and (layer0_outputs(2577));
    outputs(3244) <= layer0_outputs(4189);
    outputs(3245) <= (layer0_outputs(3895)) and not (layer0_outputs(5897));
    outputs(3246) <= layer0_outputs(4290);
    outputs(3247) <= not(layer0_outputs(2019));
    outputs(3248) <= (layer0_outputs(1439)) and not (layer0_outputs(2770));
    outputs(3249) <= not(layer0_outputs(5844));
    outputs(3250) <= layer0_outputs(2275);
    outputs(3251) <= (layer0_outputs(5109)) and not (layer0_outputs(1921));
    outputs(3252) <= layer0_outputs(1639);
    outputs(3253) <= not(layer0_outputs(6111));
    outputs(3254) <= not((layer0_outputs(437)) xor (layer0_outputs(7288)));
    outputs(3255) <= (layer0_outputs(2979)) and not (layer0_outputs(7152));
    outputs(3256) <= (layer0_outputs(5810)) and (layer0_outputs(3064));
    outputs(3257) <= (layer0_outputs(5825)) or (layer0_outputs(4188));
    outputs(3258) <= layer0_outputs(6452);
    outputs(3259) <= not(layer0_outputs(3230));
    outputs(3260) <= layer0_outputs(3865);
    outputs(3261) <= not(layer0_outputs(1553));
    outputs(3262) <= not((layer0_outputs(2666)) xor (layer0_outputs(4808)));
    outputs(3263) <= layer0_outputs(2779);
    outputs(3264) <= not(layer0_outputs(5039)) or (layer0_outputs(2662));
    outputs(3265) <= layer0_outputs(2279);
    outputs(3266) <= not((layer0_outputs(5486)) xor (layer0_outputs(6531)));
    outputs(3267) <= not(layer0_outputs(2339));
    outputs(3268) <= layer0_outputs(4333);
    outputs(3269) <= not((layer0_outputs(7425)) or (layer0_outputs(1379)));
    outputs(3270) <= (layer0_outputs(7321)) xor (layer0_outputs(184));
    outputs(3271) <= layer0_outputs(100);
    outputs(3272) <= layer0_outputs(965);
    outputs(3273) <= not(layer0_outputs(4828));
    outputs(3274) <= not((layer0_outputs(7182)) or (layer0_outputs(1459)));
    outputs(3275) <= not(layer0_outputs(6123));
    outputs(3276) <= not((layer0_outputs(4458)) or (layer0_outputs(6352)));
    outputs(3277) <= (layer0_outputs(3761)) and (layer0_outputs(519));
    outputs(3278) <= layer0_outputs(6261);
    outputs(3279) <= not((layer0_outputs(1183)) or (layer0_outputs(1419)));
    outputs(3280) <= layer0_outputs(4313);
    outputs(3281) <= layer0_outputs(7151);
    outputs(3282) <= not((layer0_outputs(1708)) or (layer0_outputs(32)));
    outputs(3283) <= not(layer0_outputs(4617));
    outputs(3284) <= not((layer0_outputs(2948)) or (layer0_outputs(4681)));
    outputs(3285) <= (layer0_outputs(3359)) and not (layer0_outputs(2141));
    outputs(3286) <= not(layer0_outputs(1652)) or (layer0_outputs(7187));
    outputs(3287) <= not((layer0_outputs(1379)) or (layer0_outputs(5782)));
    outputs(3288) <= (layer0_outputs(476)) and not (layer0_outputs(6950));
    outputs(3289) <= not((layer0_outputs(6894)) xor (layer0_outputs(7510)));
    outputs(3290) <= (layer0_outputs(5425)) xor (layer0_outputs(6659));
    outputs(3291) <= (layer0_outputs(4550)) xor (layer0_outputs(2427));
    outputs(3292) <= (layer0_outputs(499)) and not (layer0_outputs(5086));
    outputs(3293) <= not(layer0_outputs(6962));
    outputs(3294) <= layer0_outputs(4088);
    outputs(3295) <= layer0_outputs(2767);
    outputs(3296) <= (layer0_outputs(5144)) and not (layer0_outputs(6758));
    outputs(3297) <= (layer0_outputs(5284)) xor (layer0_outputs(3305));
    outputs(3298) <= not((layer0_outputs(7442)) or (layer0_outputs(5580)));
    outputs(3299) <= (layer0_outputs(4369)) and not (layer0_outputs(4098));
    outputs(3300) <= layer0_outputs(4051);
    outputs(3301) <= (layer0_outputs(26)) and not (layer0_outputs(2095));
    outputs(3302) <= not(layer0_outputs(1532));
    outputs(3303) <= not(layer0_outputs(6095));
    outputs(3304) <= not(layer0_outputs(6754)) or (layer0_outputs(4076));
    outputs(3305) <= layer0_outputs(3780);
    outputs(3306) <= not((layer0_outputs(3096)) xor (layer0_outputs(2333)));
    outputs(3307) <= (layer0_outputs(4606)) xor (layer0_outputs(2064));
    outputs(3308) <= layer0_outputs(2233);
    outputs(3309) <= layer0_outputs(120);
    outputs(3310) <= not((layer0_outputs(382)) xor (layer0_outputs(6919)));
    outputs(3311) <= (layer0_outputs(7449)) and (layer0_outputs(6103));
    outputs(3312) <= layer0_outputs(4311);
    outputs(3313) <= not((layer0_outputs(2903)) or (layer0_outputs(6830)));
    outputs(3314) <= (layer0_outputs(290)) and not (layer0_outputs(5417));
    outputs(3315) <= layer0_outputs(5883);
    outputs(3316) <= not(layer0_outputs(5494));
    outputs(3317) <= not((layer0_outputs(2457)) or (layer0_outputs(1260)));
    outputs(3318) <= (layer0_outputs(613)) or (layer0_outputs(99));
    outputs(3319) <= not(layer0_outputs(4103)) or (layer0_outputs(2050));
    outputs(3320) <= not(layer0_outputs(857));
    outputs(3321) <= (layer0_outputs(6367)) and (layer0_outputs(2669));
    outputs(3322) <= not((layer0_outputs(6918)) xor (layer0_outputs(3031)));
    outputs(3323) <= (layer0_outputs(3620)) and not (layer0_outputs(1953));
    outputs(3324) <= not(layer0_outputs(468));
    outputs(3325) <= not(layer0_outputs(3998)) or (layer0_outputs(151));
    outputs(3326) <= not(layer0_outputs(3674));
    outputs(3327) <= (layer0_outputs(5231)) and not (layer0_outputs(7671));
    outputs(3328) <= not((layer0_outputs(5939)) or (layer0_outputs(2377)));
    outputs(3329) <= layer0_outputs(125);
    outputs(3330) <= layer0_outputs(4673);
    outputs(3331) <= not(layer0_outputs(1356));
    outputs(3332) <= not((layer0_outputs(7612)) or (layer0_outputs(1724)));
    outputs(3333) <= (layer0_outputs(4689)) and (layer0_outputs(5199));
    outputs(3334) <= layer0_outputs(6539);
    outputs(3335) <= (layer0_outputs(6724)) xor (layer0_outputs(4137));
    outputs(3336) <= not((layer0_outputs(2627)) and (layer0_outputs(6630)));
    outputs(3337) <= layer0_outputs(7121);
    outputs(3338) <= not(layer0_outputs(2004));
    outputs(3339) <= (layer0_outputs(1746)) and not (layer0_outputs(539));
    outputs(3340) <= (layer0_outputs(2353)) xor (layer0_outputs(6444));
    outputs(3341) <= (layer0_outputs(4463)) xor (layer0_outputs(40));
    outputs(3342) <= not(layer0_outputs(6200));
    outputs(3343) <= (layer0_outputs(4163)) and not (layer0_outputs(5909));
    outputs(3344) <= layer0_outputs(6462);
    outputs(3345) <= (layer0_outputs(4997)) and not (layer0_outputs(6443));
    outputs(3346) <= not(layer0_outputs(5168));
    outputs(3347) <= not((layer0_outputs(6350)) or (layer0_outputs(1055)));
    outputs(3348) <= (layer0_outputs(7065)) and (layer0_outputs(2042));
    outputs(3349) <= not(layer0_outputs(2983));
    outputs(3350) <= not((layer0_outputs(6415)) xor (layer0_outputs(1011)));
    outputs(3351) <= not(layer0_outputs(1386));
    outputs(3352) <= (layer0_outputs(1065)) xor (layer0_outputs(6674));
    outputs(3353) <= (layer0_outputs(2784)) and not (layer0_outputs(1830));
    outputs(3354) <= not(layer0_outputs(5461));
    outputs(3355) <= (layer0_outputs(1098)) and not (layer0_outputs(4500));
    outputs(3356) <= not(layer0_outputs(2948)) or (layer0_outputs(3132));
    outputs(3357) <= (layer0_outputs(1305)) and not (layer0_outputs(7139));
    outputs(3358) <= not(layer0_outputs(4487)) or (layer0_outputs(4384));
    outputs(3359) <= layer0_outputs(614);
    outputs(3360) <= not((layer0_outputs(2131)) xor (layer0_outputs(4609)));
    outputs(3361) <= layer0_outputs(78);
    outputs(3362) <= not((layer0_outputs(5525)) or (layer0_outputs(5460)));
    outputs(3363) <= not(layer0_outputs(6068));
    outputs(3364) <= not(layer0_outputs(5764));
    outputs(3365) <= (layer0_outputs(6131)) or (layer0_outputs(6323));
    outputs(3366) <= layer0_outputs(4596);
    outputs(3367) <= (layer0_outputs(5759)) and not (layer0_outputs(6609));
    outputs(3368) <= (layer0_outputs(6023)) and not (layer0_outputs(6756));
    outputs(3369) <= not(layer0_outputs(993));
    outputs(3370) <= not(layer0_outputs(2309));
    outputs(3371) <= not(layer0_outputs(7157));
    outputs(3372) <= layer0_outputs(6092);
    outputs(3373) <= not(layer0_outputs(162));
    outputs(3374) <= (layer0_outputs(6563)) xor (layer0_outputs(557));
    outputs(3375) <= layer0_outputs(2398);
    outputs(3376) <= layer0_outputs(4074);
    outputs(3377) <= not((layer0_outputs(2324)) xor (layer0_outputs(7211)));
    outputs(3378) <= layer0_outputs(3371);
    outputs(3379) <= not(layer0_outputs(5663));
    outputs(3380) <= layer0_outputs(4789);
    outputs(3381) <= (layer0_outputs(1100)) xor (layer0_outputs(3888));
    outputs(3382) <= (layer0_outputs(373)) xor (layer0_outputs(2258));
    outputs(3383) <= not(layer0_outputs(5069));
    outputs(3384) <= not((layer0_outputs(5037)) or (layer0_outputs(6785)));
    outputs(3385) <= not((layer0_outputs(6657)) or (layer0_outputs(5088)));
    outputs(3386) <= not((layer0_outputs(4550)) xor (layer0_outputs(3193)));
    outputs(3387) <= not(layer0_outputs(6448)) or (layer0_outputs(4329));
    outputs(3388) <= (layer0_outputs(5506)) and not (layer0_outputs(298));
    outputs(3389) <= not(layer0_outputs(1679)) or (layer0_outputs(4650));
    outputs(3390) <= (layer0_outputs(3692)) xor (layer0_outputs(5068));
    outputs(3391) <= layer0_outputs(4125);
    outputs(3392) <= (layer0_outputs(3097)) and not (layer0_outputs(1373));
    outputs(3393) <= (layer0_outputs(811)) xor (layer0_outputs(1693));
    outputs(3394) <= not(layer0_outputs(2670));
    outputs(3395) <= not(layer0_outputs(3687));
    outputs(3396) <= not((layer0_outputs(5940)) or (layer0_outputs(3800)));
    outputs(3397) <= not(layer0_outputs(7009));
    outputs(3398) <= not((layer0_outputs(1091)) xor (layer0_outputs(1514)));
    outputs(3399) <= not(layer0_outputs(6928)) or (layer0_outputs(7254));
    outputs(3400) <= layer0_outputs(188);
    outputs(3401) <= (layer0_outputs(6570)) and not (layer0_outputs(6319));
    outputs(3402) <= not((layer0_outputs(5958)) or (layer0_outputs(6303)));
    outputs(3403) <= not(layer0_outputs(2368));
    outputs(3404) <= layer0_outputs(5864);
    outputs(3405) <= layer0_outputs(5575);
    outputs(3406) <= layer0_outputs(7080);
    outputs(3407) <= layer0_outputs(2838);
    outputs(3408) <= not(layer0_outputs(2529));
    outputs(3409) <= (layer0_outputs(408)) and (layer0_outputs(3177));
    outputs(3410) <= not((layer0_outputs(2216)) and (layer0_outputs(3559)));
    outputs(3411) <= (layer0_outputs(332)) and not (layer0_outputs(2824));
    outputs(3412) <= not(layer0_outputs(3923));
    outputs(3413) <= not((layer0_outputs(2857)) xor (layer0_outputs(1551)));
    outputs(3414) <= layer0_outputs(4926);
    outputs(3415) <= not((layer0_outputs(1587)) and (layer0_outputs(2912)));
    outputs(3416) <= not(layer0_outputs(118));
    outputs(3417) <= layer0_outputs(2270);
    outputs(3418) <= not(layer0_outputs(4013));
    outputs(3419) <= (layer0_outputs(1910)) and not (layer0_outputs(6743));
    outputs(3420) <= layer0_outputs(2108);
    outputs(3421) <= (layer0_outputs(1788)) and not (layer0_outputs(2569));
    outputs(3422) <= not((layer0_outputs(5298)) or (layer0_outputs(3221)));
    outputs(3423) <= (layer0_outputs(2266)) xor (layer0_outputs(5036));
    outputs(3424) <= not((layer0_outputs(679)) xor (layer0_outputs(424)));
    outputs(3425) <= not(layer0_outputs(1738));
    outputs(3426) <= layer0_outputs(4674);
    outputs(3427) <= layer0_outputs(442);
    outputs(3428) <= layer0_outputs(754);
    outputs(3429) <= not(layer0_outputs(5741));
    outputs(3430) <= not(layer0_outputs(7593));
    outputs(3431) <= not(layer0_outputs(3090));
    outputs(3432) <= not(layer0_outputs(1756));
    outputs(3433) <= not((layer0_outputs(7456)) or (layer0_outputs(657)));
    outputs(3434) <= not((layer0_outputs(126)) or (layer0_outputs(1886)));
    outputs(3435) <= not(layer0_outputs(2764));
    outputs(3436) <= layer0_outputs(4399);
    outputs(3437) <= not((layer0_outputs(2106)) and (layer0_outputs(5320)));
    outputs(3438) <= not((layer0_outputs(6186)) or (layer0_outputs(5988)));
    outputs(3439) <= layer0_outputs(1906);
    outputs(3440) <= not(layer0_outputs(6608));
    outputs(3441) <= (layer0_outputs(4454)) or (layer0_outputs(3825));
    outputs(3442) <= not(layer0_outputs(6936));
    outputs(3443) <= not((layer0_outputs(941)) or (layer0_outputs(5204)));
    outputs(3444) <= not(layer0_outputs(4967)) or (layer0_outputs(7592));
    outputs(3445) <= not(layer0_outputs(6376));
    outputs(3446) <= not((layer0_outputs(704)) and (layer0_outputs(7558)));
    outputs(3447) <= (layer0_outputs(4538)) xor (layer0_outputs(3070));
    outputs(3448) <= not(layer0_outputs(2488)) or (layer0_outputs(3759));
    outputs(3449) <= not((layer0_outputs(2175)) or (layer0_outputs(4995)));
    outputs(3450) <= not((layer0_outputs(7346)) and (layer0_outputs(6999)));
    outputs(3451) <= layer0_outputs(4960);
    outputs(3452) <= not(layer0_outputs(465)) or (layer0_outputs(2578));
    outputs(3453) <= (layer0_outputs(5652)) and (layer0_outputs(4128));
    outputs(3454) <= not((layer0_outputs(2596)) xor (layer0_outputs(5788)));
    outputs(3455) <= layer0_outputs(532);
    outputs(3456) <= layer0_outputs(2848);
    outputs(3457) <= layer0_outputs(5548);
    outputs(3458) <= not(layer0_outputs(4111)) or (layer0_outputs(6286));
    outputs(3459) <= layer0_outputs(348);
    outputs(3460) <= (layer0_outputs(731)) and not (layer0_outputs(6327));
    outputs(3461) <= layer0_outputs(3868);
    outputs(3462) <= layer0_outputs(3989);
    outputs(3463) <= layer0_outputs(5110);
    outputs(3464) <= not(layer0_outputs(3073));
    outputs(3465) <= (layer0_outputs(1330)) xor (layer0_outputs(6754));
    outputs(3466) <= layer0_outputs(1178);
    outputs(3467) <= layer0_outputs(4074);
    outputs(3468) <= (layer0_outputs(4048)) and (layer0_outputs(2504));
    outputs(3469) <= not((layer0_outputs(5332)) or (layer0_outputs(1830)));
    outputs(3470) <= layer0_outputs(4297);
    outputs(3471) <= not(layer0_outputs(2993));
    outputs(3472) <= layer0_outputs(5812);
    outputs(3473) <= not((layer0_outputs(3648)) xor (layer0_outputs(6149)));
    outputs(3474) <= layer0_outputs(5011);
    outputs(3475) <= layer0_outputs(4077);
    outputs(3476) <= not(layer0_outputs(4260));
    outputs(3477) <= (layer0_outputs(5148)) and (layer0_outputs(765));
    outputs(3478) <= not((layer0_outputs(4231)) xor (layer0_outputs(4284)));
    outputs(3479) <= (layer0_outputs(2049)) and not (layer0_outputs(2849));
    outputs(3480) <= (layer0_outputs(5928)) and not (layer0_outputs(5132));
    outputs(3481) <= layer0_outputs(3811);
    outputs(3482) <= layer0_outputs(5772);
    outputs(3483) <= (layer0_outputs(2958)) xor (layer0_outputs(3526));
    outputs(3484) <= (layer0_outputs(7284)) xor (layer0_outputs(5631));
    outputs(3485) <= layer0_outputs(6412);
    outputs(3486) <= not((layer0_outputs(1093)) xor (layer0_outputs(4983)));
    outputs(3487) <= not(layer0_outputs(4172)) or (layer0_outputs(434));
    outputs(3488) <= not((layer0_outputs(3968)) or (layer0_outputs(3432)));
    outputs(3489) <= (layer0_outputs(4462)) and (layer0_outputs(861));
    outputs(3490) <= layer0_outputs(5610);
    outputs(3491) <= not(layer0_outputs(2614));
    outputs(3492) <= not((layer0_outputs(1813)) or (layer0_outputs(3763)));
    outputs(3493) <= (layer0_outputs(4648)) and not (layer0_outputs(6749));
    outputs(3494) <= layer0_outputs(4180);
    outputs(3495) <= not(layer0_outputs(5375));
    outputs(3496) <= not((layer0_outputs(3794)) xor (layer0_outputs(1951)));
    outputs(3497) <= not((layer0_outputs(4002)) or (layer0_outputs(1084)));
    outputs(3498) <= (layer0_outputs(1988)) and not (layer0_outputs(15));
    outputs(3499) <= (layer0_outputs(7521)) and not (layer0_outputs(4644));
    outputs(3500) <= (layer0_outputs(1485)) and not (layer0_outputs(6514));
    outputs(3501) <= not(layer0_outputs(2531));
    outputs(3502) <= layer0_outputs(4841);
    outputs(3503) <= layer0_outputs(2111);
    outputs(3504) <= layer0_outputs(5390);
    outputs(3505) <= layer0_outputs(7445);
    outputs(3506) <= not(layer0_outputs(4012));
    outputs(3507) <= layer0_outputs(3177);
    outputs(3508) <= (layer0_outputs(171)) and not (layer0_outputs(5941));
    outputs(3509) <= not(layer0_outputs(6564));
    outputs(3510) <= not(layer0_outputs(4970));
    outputs(3511) <= not(layer0_outputs(6058));
    outputs(3512) <= layer0_outputs(5031);
    outputs(3513) <= layer0_outputs(121);
    outputs(3514) <= (layer0_outputs(437)) and not (layer0_outputs(4725));
    outputs(3515) <= (layer0_outputs(4113)) and (layer0_outputs(2584));
    outputs(3516) <= (layer0_outputs(7584)) and not (layer0_outputs(4162));
    outputs(3517) <= layer0_outputs(1928);
    outputs(3518) <= layer0_outputs(3690);
    outputs(3519) <= (layer0_outputs(168)) and not (layer0_outputs(6345));
    outputs(3520) <= not(layer0_outputs(3552));
    outputs(3521) <= not(layer0_outputs(4772)) or (layer0_outputs(4807));
    outputs(3522) <= layer0_outputs(5667);
    outputs(3523) <= not(layer0_outputs(344));
    outputs(3524) <= not(layer0_outputs(995));
    outputs(3525) <= not((layer0_outputs(7063)) or (layer0_outputs(7204)));
    outputs(3526) <= layer0_outputs(690);
    outputs(3527) <= not(layer0_outputs(4643));
    outputs(3528) <= not((layer0_outputs(1962)) or (layer0_outputs(4699)));
    outputs(3529) <= layer0_outputs(2946);
    outputs(3530) <= not(layer0_outputs(4849));
    outputs(3531) <= (layer0_outputs(56)) xor (layer0_outputs(2502));
    outputs(3532) <= (layer0_outputs(158)) and (layer0_outputs(4651));
    outputs(3533) <= not(layer0_outputs(1127));
    outputs(3534) <= not(layer0_outputs(1312));
    outputs(3535) <= layer0_outputs(4755);
    outputs(3536) <= not((layer0_outputs(5246)) and (layer0_outputs(7576)));
    outputs(3537) <= (layer0_outputs(223)) and not (layer0_outputs(4677));
    outputs(3538) <= not(layer0_outputs(2586)) or (layer0_outputs(3434));
    outputs(3539) <= not(layer0_outputs(2023)) or (layer0_outputs(5397));
    outputs(3540) <= (layer0_outputs(5354)) and not (layer0_outputs(2418));
    outputs(3541) <= (layer0_outputs(580)) and (layer0_outputs(2967));
    outputs(3542) <= (layer0_outputs(4591)) and not (layer0_outputs(436));
    outputs(3543) <= not(layer0_outputs(2629)) or (layer0_outputs(6996));
    outputs(3544) <= not(layer0_outputs(175));
    outputs(3545) <= (layer0_outputs(2848)) and not (layer0_outputs(1327));
    outputs(3546) <= (layer0_outputs(6870)) and not (layer0_outputs(4403));
    outputs(3547) <= not(layer0_outputs(4047));
    outputs(3548) <= (layer0_outputs(1117)) and not (layer0_outputs(2768));
    outputs(3549) <= not((layer0_outputs(1346)) or (layer0_outputs(2598)));
    outputs(3550) <= layer0_outputs(1013);
    outputs(3551) <= not((layer0_outputs(5938)) and (layer0_outputs(3175)));
    outputs(3552) <= (layer0_outputs(136)) or (layer0_outputs(3628));
    outputs(3553) <= (layer0_outputs(6441)) and not (layer0_outputs(2698));
    outputs(3554) <= not(layer0_outputs(7261)) or (layer0_outputs(1387));
    outputs(3555) <= not(layer0_outputs(4710));
    outputs(3556) <= layer0_outputs(758);
    outputs(3557) <= not(layer0_outputs(2243));
    outputs(3558) <= (layer0_outputs(1051)) xor (layer0_outputs(707));
    outputs(3559) <= not(layer0_outputs(3694));
    outputs(3560) <= not((layer0_outputs(1269)) or (layer0_outputs(7328)));
    outputs(3561) <= (layer0_outputs(2843)) and not (layer0_outputs(2841));
    outputs(3562) <= (layer0_outputs(1700)) xor (layer0_outputs(7465));
    outputs(3563) <= (layer0_outputs(3870)) and not (layer0_outputs(4995));
    outputs(3564) <= not(layer0_outputs(2633));
    outputs(3565) <= (layer0_outputs(4769)) xor (layer0_outputs(4612));
    outputs(3566) <= not((layer0_outputs(2039)) xor (layer0_outputs(2156)));
    outputs(3567) <= not(layer0_outputs(388)) or (layer0_outputs(887));
    outputs(3568) <= layer0_outputs(6295);
    outputs(3569) <= not(layer0_outputs(6265));
    outputs(3570) <= (layer0_outputs(577)) or (layer0_outputs(2861));
    outputs(3571) <= layer0_outputs(5805);
    outputs(3572) <= not(layer0_outputs(3517)) or (layer0_outputs(7058));
    outputs(3573) <= layer0_outputs(1415);
    outputs(3574) <= (layer0_outputs(898)) and (layer0_outputs(951));
    outputs(3575) <= not(layer0_outputs(536));
    outputs(3576) <= (layer0_outputs(5801)) xor (layer0_outputs(114));
    outputs(3577) <= not(layer0_outputs(2612));
    outputs(3578) <= layer0_outputs(7156);
    outputs(3579) <= (layer0_outputs(5051)) and (layer0_outputs(4548));
    outputs(3580) <= not(layer0_outputs(5266));
    outputs(3581) <= not(layer0_outputs(5585));
    outputs(3582) <= not(layer0_outputs(5751));
    outputs(3583) <= layer0_outputs(7317);
    outputs(3584) <= (layer0_outputs(2132)) xor (layer0_outputs(5809));
    outputs(3585) <= not((layer0_outputs(5771)) or (layer0_outputs(5597)));
    outputs(3586) <= layer0_outputs(3940);
    outputs(3587) <= layer0_outputs(3977);
    outputs(3588) <= not(layer0_outputs(2378));
    outputs(3589) <= not(layer0_outputs(5004));
    outputs(3590) <= (layer0_outputs(6523)) xor (layer0_outputs(5655));
    outputs(3591) <= layer0_outputs(4694);
    outputs(3592) <= layer0_outputs(4844);
    outputs(3593) <= not((layer0_outputs(5630)) xor (layer0_outputs(3149)));
    outputs(3594) <= layer0_outputs(1512);
    outputs(3595) <= not(layer0_outputs(4261));
    outputs(3596) <= not((layer0_outputs(4574)) and (layer0_outputs(878)));
    outputs(3597) <= layer0_outputs(3903);
    outputs(3598) <= (layer0_outputs(2462)) and not (layer0_outputs(6411));
    outputs(3599) <= not(layer0_outputs(7664)) or (layer0_outputs(2988));
    outputs(3600) <= (layer0_outputs(2479)) xor (layer0_outputs(1474));
    outputs(3601) <= not(layer0_outputs(5625)) or (layer0_outputs(3267));
    outputs(3602) <= not(layer0_outputs(3553)) or (layer0_outputs(1309));
    outputs(3603) <= not((layer0_outputs(6369)) and (layer0_outputs(3019)));
    outputs(3604) <= not(layer0_outputs(2166)) or (layer0_outputs(7027));
    outputs(3605) <= not((layer0_outputs(6159)) xor (layer0_outputs(1752)));
    outputs(3606) <= layer0_outputs(586);
    outputs(3607) <= (layer0_outputs(5802)) and not (layer0_outputs(144));
    outputs(3608) <= layer0_outputs(4424);
    outputs(3609) <= not(layer0_outputs(2622));
    outputs(3610) <= not(layer0_outputs(5113));
    outputs(3611) <= (layer0_outputs(6987)) and not (layer0_outputs(3246));
    outputs(3612) <= not(layer0_outputs(1373));
    outputs(3613) <= layer0_outputs(5198);
    outputs(3614) <= not(layer0_outputs(5220)) or (layer0_outputs(6084));
    outputs(3615) <= not(layer0_outputs(7210));
    outputs(3616) <= not(layer0_outputs(972));
    outputs(3617) <= layer0_outputs(2495);
    outputs(3618) <= not(layer0_outputs(7310));
    outputs(3619) <= not(layer0_outputs(6596));
    outputs(3620) <= not(layer0_outputs(6068));
    outputs(3621) <= (layer0_outputs(2411)) and (layer0_outputs(4521));
    outputs(3622) <= (layer0_outputs(1142)) xor (layer0_outputs(3328));
    outputs(3623) <= not((layer0_outputs(7246)) xor (layer0_outputs(819)));
    outputs(3624) <= not(layer0_outputs(5348));
    outputs(3625) <= not(layer0_outputs(4283)) or (layer0_outputs(6757));
    outputs(3626) <= not(layer0_outputs(6115));
    outputs(3627) <= (layer0_outputs(340)) and not (layer0_outputs(2451));
    outputs(3628) <= not((layer0_outputs(2198)) xor (layer0_outputs(2036)));
    outputs(3629) <= not(layer0_outputs(6551)) or (layer0_outputs(7418));
    outputs(3630) <= not((layer0_outputs(6534)) or (layer0_outputs(379)));
    outputs(3631) <= layer0_outputs(1267);
    outputs(3632) <= layer0_outputs(3547);
    outputs(3633) <= not(layer0_outputs(1658));
    outputs(3634) <= not((layer0_outputs(905)) xor (layer0_outputs(608)));
    outputs(3635) <= not(layer0_outputs(500));
    outputs(3636) <= not(layer0_outputs(529));
    outputs(3637) <= layer0_outputs(3508);
    outputs(3638) <= not(layer0_outputs(2914));
    outputs(3639) <= (layer0_outputs(3593)) and not (layer0_outputs(1570));
    outputs(3640) <= (layer0_outputs(1224)) and (layer0_outputs(1744));
    outputs(3641) <= layer0_outputs(6446);
    outputs(3642) <= (layer0_outputs(5371)) and (layer0_outputs(7594));
    outputs(3643) <= not(layer0_outputs(3332));
    outputs(3644) <= (layer0_outputs(7126)) xor (layer0_outputs(1977));
    outputs(3645) <= layer0_outputs(3458);
    outputs(3646) <= not((layer0_outputs(658)) or (layer0_outputs(4295)));
    outputs(3647) <= layer0_outputs(4596);
    outputs(3648) <= (layer0_outputs(386)) and not (layer0_outputs(4208));
    outputs(3649) <= (layer0_outputs(3849)) and not (layer0_outputs(5707));
    outputs(3650) <= not((layer0_outputs(7548)) xor (layer0_outputs(2128)));
    outputs(3651) <= layer0_outputs(2701);
    outputs(3652) <= not(layer0_outputs(712));
    outputs(3653) <= (layer0_outputs(1751)) xor (layer0_outputs(5254));
    outputs(3654) <= layer0_outputs(3576);
    outputs(3655) <= (layer0_outputs(124)) and (layer0_outputs(6124));
    outputs(3656) <= not((layer0_outputs(3550)) xor (layer0_outputs(2105)));
    outputs(3657) <= layer0_outputs(5091);
    outputs(3658) <= not((layer0_outputs(7461)) or (layer0_outputs(7539)));
    outputs(3659) <= layer0_outputs(7505);
    outputs(3660) <= not((layer0_outputs(5475)) xor (layer0_outputs(770)));
    outputs(3661) <= (layer0_outputs(926)) xor (layer0_outputs(6528));
    outputs(3662) <= layer0_outputs(4029);
    outputs(3663) <= not(layer0_outputs(4300)) or (layer0_outputs(6942));
    outputs(3664) <= (layer0_outputs(1585)) xor (layer0_outputs(2788));
    outputs(3665) <= (layer0_outputs(2016)) xor (layer0_outputs(178));
    outputs(3666) <= not(layer0_outputs(5738));
    outputs(3667) <= not(layer0_outputs(4263));
    outputs(3668) <= not(layer0_outputs(7656));
    outputs(3669) <= (layer0_outputs(1965)) and not (layer0_outputs(7580));
    outputs(3670) <= (layer0_outputs(3769)) and not (layer0_outputs(6376));
    outputs(3671) <= not(layer0_outputs(4940));
    outputs(3672) <= not(layer0_outputs(3155)) or (layer0_outputs(440));
    outputs(3673) <= (layer0_outputs(935)) and not (layer0_outputs(5391));
    outputs(3674) <= not(layer0_outputs(3179));
    outputs(3675) <= not(layer0_outputs(7459)) or (layer0_outputs(355));
    outputs(3676) <= not(layer0_outputs(104));
    outputs(3677) <= not((layer0_outputs(2706)) xor (layer0_outputs(5111)));
    outputs(3678) <= layer0_outputs(1137);
    outputs(3679) <= not((layer0_outputs(1280)) or (layer0_outputs(6908)));
    outputs(3680) <= not(layer0_outputs(973)) or (layer0_outputs(6000));
    outputs(3681) <= (layer0_outputs(4143)) or (layer0_outputs(4254));
    outputs(3682) <= not(layer0_outputs(2325)) or (layer0_outputs(1291));
    outputs(3683) <= (layer0_outputs(3608)) and not (layer0_outputs(6764));
    outputs(3684) <= not((layer0_outputs(5768)) and (layer0_outputs(1212)));
    outputs(3685) <= (layer0_outputs(3611)) and not (layer0_outputs(1880));
    outputs(3686) <= not((layer0_outputs(4087)) or (layer0_outputs(460)));
    outputs(3687) <= layer0_outputs(1482);
    outputs(3688) <= not(layer0_outputs(624)) or (layer0_outputs(3217));
    outputs(3689) <= (layer0_outputs(4304)) and not (layer0_outputs(634));
    outputs(3690) <= not(layer0_outputs(6034));
    outputs(3691) <= (layer0_outputs(5302)) xor (layer0_outputs(5536));
    outputs(3692) <= not(layer0_outputs(5306));
    outputs(3693) <= not((layer0_outputs(2502)) or (layer0_outputs(1471)));
    outputs(3694) <= not(layer0_outputs(6139));
    outputs(3695) <= not(layer0_outputs(5289));
    outputs(3696) <= not((layer0_outputs(6011)) xor (layer0_outputs(5028)));
    outputs(3697) <= not((layer0_outputs(444)) xor (layer0_outputs(2066)));
    outputs(3698) <= layer0_outputs(7039);
    outputs(3699) <= not(layer0_outputs(7669)) or (layer0_outputs(4888));
    outputs(3700) <= not((layer0_outputs(1767)) and (layer0_outputs(4495)));
    outputs(3701) <= layer0_outputs(5608);
    outputs(3702) <= not(layer0_outputs(276));
    outputs(3703) <= not(layer0_outputs(1633)) or (layer0_outputs(3881));
    outputs(3704) <= not(layer0_outputs(2629));
    outputs(3705) <= layer0_outputs(7579);
    outputs(3706) <= not(layer0_outputs(5351));
    outputs(3707) <= (layer0_outputs(813)) xor (layer0_outputs(1421));
    outputs(3708) <= (layer0_outputs(4597)) xor (layer0_outputs(6605));
    outputs(3709) <= not(layer0_outputs(2792));
    outputs(3710) <= (layer0_outputs(3309)) and not (layer0_outputs(4724));
    outputs(3711) <= layer0_outputs(3626);
    outputs(3712) <= not((layer0_outputs(3276)) xor (layer0_outputs(4003)));
    outputs(3713) <= (layer0_outputs(1833)) and not (layer0_outputs(5296));
    outputs(3714) <= not(layer0_outputs(1641)) or (layer0_outputs(224));
    outputs(3715) <= (layer0_outputs(1279)) or (layer0_outputs(1994));
    outputs(3716) <= (layer0_outputs(452)) xor (layer0_outputs(4624));
    outputs(3717) <= (layer0_outputs(8)) and (layer0_outputs(956));
    outputs(3718) <= (layer0_outputs(7001)) or (layer0_outputs(3381));
    outputs(3719) <= not(layer0_outputs(3185));
    outputs(3720) <= (layer0_outputs(5609)) and (layer0_outputs(4409));
    outputs(3721) <= not((layer0_outputs(3788)) and (layer0_outputs(337)));
    outputs(3722) <= (layer0_outputs(6607)) and (layer0_outputs(6816));
    outputs(3723) <= not((layer0_outputs(7464)) and (layer0_outputs(36)));
    outputs(3724) <= (layer0_outputs(5769)) xor (layer0_outputs(1251));
    outputs(3725) <= (layer0_outputs(3738)) and not (layer0_outputs(5096));
    outputs(3726) <= layer0_outputs(1140);
    outputs(3727) <= (layer0_outputs(4080)) xor (layer0_outputs(5747));
    outputs(3728) <= (layer0_outputs(4123)) or (layer0_outputs(4005));
    outputs(3729) <= not(layer0_outputs(1789));
    outputs(3730) <= not((layer0_outputs(3321)) or (layer0_outputs(4537)));
    outputs(3731) <= (layer0_outputs(6827)) or (layer0_outputs(4318));
    outputs(3732) <= (layer0_outputs(7385)) xor (layer0_outputs(6950));
    outputs(3733) <= layer0_outputs(2765);
    outputs(3734) <= (layer0_outputs(6993)) and not (layer0_outputs(2997));
    outputs(3735) <= not(layer0_outputs(2738)) or (layer0_outputs(2471));
    outputs(3736) <= (layer0_outputs(7007)) and (layer0_outputs(7634));
    outputs(3737) <= layer0_outputs(6870);
    outputs(3738) <= layer0_outputs(2775);
    outputs(3739) <= (layer0_outputs(5955)) and not (layer0_outputs(6486));
    outputs(3740) <= not((layer0_outputs(7141)) or (layer0_outputs(3871)));
    outputs(3741) <= (layer0_outputs(7474)) xor (layer0_outputs(505));
    outputs(3742) <= (layer0_outputs(1001)) and (layer0_outputs(3903));
    outputs(3743) <= not((layer0_outputs(7533)) xor (layer0_outputs(2636)));
    outputs(3744) <= (layer0_outputs(5117)) and (layer0_outputs(6419));
    outputs(3745) <= not(layer0_outputs(706));
    outputs(3746) <= not(layer0_outputs(5523));
    outputs(3747) <= layer0_outputs(5059);
    outputs(3748) <= not((layer0_outputs(4083)) or (layer0_outputs(6954)));
    outputs(3749) <= not(layer0_outputs(480)) or (layer0_outputs(5008));
    outputs(3750) <= not(layer0_outputs(5289));
    outputs(3751) <= layer0_outputs(1990);
    outputs(3752) <= not(layer0_outputs(6715));
    outputs(3753) <= (layer0_outputs(542)) xor (layer0_outputs(5637));
    outputs(3754) <= not(layer0_outputs(839));
    outputs(3755) <= (layer0_outputs(4171)) xor (layer0_outputs(2548));
    outputs(3756) <= layer0_outputs(5043);
    outputs(3757) <= layer0_outputs(7018);
    outputs(3758) <= (layer0_outputs(6784)) and (layer0_outputs(7422));
    outputs(3759) <= layer0_outputs(7238);
    outputs(3760) <= not(layer0_outputs(5558)) or (layer0_outputs(5549));
    outputs(3761) <= not((layer0_outputs(6284)) xor (layer0_outputs(5227)));
    outputs(3762) <= not((layer0_outputs(167)) or (layer0_outputs(2235)));
    outputs(3763) <= not((layer0_outputs(4764)) xor (layer0_outputs(1251)));
    outputs(3764) <= not(layer0_outputs(6392));
    outputs(3765) <= (layer0_outputs(4551)) and (layer0_outputs(5264));
    outputs(3766) <= not((layer0_outputs(7552)) or (layer0_outputs(4104)));
    outputs(3767) <= not(layer0_outputs(4102)) or (layer0_outputs(519));
    outputs(3768) <= not(layer0_outputs(2782));
    outputs(3769) <= not(layer0_outputs(5877)) or (layer0_outputs(865));
    outputs(3770) <= (layer0_outputs(5683)) and (layer0_outputs(7133));
    outputs(3771) <= layer0_outputs(5308);
    outputs(3772) <= layer0_outputs(5363);
    outputs(3773) <= (layer0_outputs(523)) and (layer0_outputs(3002));
    outputs(3774) <= (layer0_outputs(873)) and (layer0_outputs(4672));
    outputs(3775) <= (layer0_outputs(5546)) and not (layer0_outputs(5037));
    outputs(3776) <= (layer0_outputs(5826)) and not (layer0_outputs(3713));
    outputs(3777) <= not((layer0_outputs(5762)) xor (layer0_outputs(1332)));
    outputs(3778) <= not(layer0_outputs(51));
    outputs(3779) <= layer0_outputs(6148);
    outputs(3780) <= layer0_outputs(5934);
    outputs(3781) <= (layer0_outputs(774)) and not (layer0_outputs(5010));
    outputs(3782) <= not(layer0_outputs(1634));
    outputs(3783) <= (layer0_outputs(110)) or (layer0_outputs(3705));
    outputs(3784) <= layer0_outputs(4922);
    outputs(3785) <= (layer0_outputs(7198)) and (layer0_outputs(1567));
    outputs(3786) <= (layer0_outputs(2058)) and not (layer0_outputs(1235));
    outputs(3787) <= layer0_outputs(7546);
    outputs(3788) <= (layer0_outputs(3379)) and not (layer0_outputs(5249));
    outputs(3789) <= (layer0_outputs(751)) xor (layer0_outputs(6670));
    outputs(3790) <= layer0_outputs(3360);
    outputs(3791) <= not(layer0_outputs(559));
    outputs(3792) <= layer0_outputs(5696);
    outputs(3793) <= not(layer0_outputs(3555));
    outputs(3794) <= not((layer0_outputs(7507)) xor (layer0_outputs(865)));
    outputs(3795) <= (layer0_outputs(1940)) xor (layer0_outputs(261));
    outputs(3796) <= not((layer0_outputs(2772)) and (layer0_outputs(2659)));
    outputs(3797) <= not(layer0_outputs(4493));
    outputs(3798) <= (layer0_outputs(1644)) and not (layer0_outputs(6520));
    outputs(3799) <= not(layer0_outputs(2418));
    outputs(3800) <= (layer0_outputs(7414)) and not (layer0_outputs(927));
    outputs(3801) <= not((layer0_outputs(943)) or (layer0_outputs(3333)));
    outputs(3802) <= not(layer0_outputs(4435));
    outputs(3803) <= not(layer0_outputs(6889));
    outputs(3804) <= not((layer0_outputs(5663)) and (layer0_outputs(4803)));
    outputs(3805) <= (layer0_outputs(2124)) or (layer0_outputs(4315));
    outputs(3806) <= layer0_outputs(1279);
    outputs(3807) <= layer0_outputs(5499);
    outputs(3808) <= (layer0_outputs(1647)) and not (layer0_outputs(4525));
    outputs(3809) <= layer0_outputs(5257);
    outputs(3810) <= (layer0_outputs(4242)) and not (layer0_outputs(4899));
    outputs(3811) <= layer0_outputs(4595);
    outputs(3812) <= layer0_outputs(5544);
    outputs(3813) <= not(layer0_outputs(4458));
    outputs(3814) <= not(layer0_outputs(1201));
    outputs(3815) <= not(layer0_outputs(236));
    outputs(3816) <= not(layer0_outputs(1820));
    outputs(3817) <= not(layer0_outputs(4800)) or (layer0_outputs(1956));
    outputs(3818) <= layer0_outputs(6322);
    outputs(3819) <= not(layer0_outputs(5967));
    outputs(3820) <= not(layer0_outputs(84));
    outputs(3821) <= (layer0_outputs(4581)) and not (layer0_outputs(2283));
    outputs(3822) <= layer0_outputs(4505);
    outputs(3823) <= (layer0_outputs(4062)) xor (layer0_outputs(1700));
    outputs(3824) <= (layer0_outputs(7280)) and (layer0_outputs(3817));
    outputs(3825) <= not(layer0_outputs(5217));
    outputs(3826) <= not(layer0_outputs(831)) or (layer0_outputs(7343));
    outputs(3827) <= layer0_outputs(2779);
    outputs(3828) <= not((layer0_outputs(5295)) or (layer0_outputs(1461)));
    outputs(3829) <= not(layer0_outputs(5905));
    outputs(3830) <= not(layer0_outputs(5894));
    outputs(3831) <= (layer0_outputs(4311)) xor (layer0_outputs(1674));
    outputs(3832) <= not(layer0_outputs(6566));
    outputs(3833) <= layer0_outputs(4805);
    outputs(3834) <= not(layer0_outputs(5920)) or (layer0_outputs(7428));
    outputs(3835) <= not(layer0_outputs(7366));
    outputs(3836) <= not(layer0_outputs(2346));
    outputs(3837) <= (layer0_outputs(4102)) xor (layer0_outputs(4893));
    outputs(3838) <= not((layer0_outputs(2554)) xor (layer0_outputs(4949)));
    outputs(3839) <= not((layer0_outputs(1699)) xor (layer0_outputs(4369)));
    outputs(3840) <= layer0_outputs(1009);
    outputs(3841) <= not(layer0_outputs(612));
    outputs(3842) <= not(layer0_outputs(1850));
    outputs(3843) <= layer0_outputs(7076);
    outputs(3844) <= (layer0_outputs(4977)) xor (layer0_outputs(2637));
    outputs(3845) <= not(layer0_outputs(2652)) or (layer0_outputs(553));
    outputs(3846) <= not(layer0_outputs(4542));
    outputs(3847) <= not(layer0_outputs(2525));
    outputs(3848) <= not(layer0_outputs(6153)) or (layer0_outputs(2527));
    outputs(3849) <= not((layer0_outputs(990)) xor (layer0_outputs(3325)));
    outputs(3850) <= (layer0_outputs(649)) and (layer0_outputs(258));
    outputs(3851) <= not(layer0_outputs(5468));
    outputs(3852) <= layer0_outputs(1762);
    outputs(3853) <= not(layer0_outputs(4645));
    outputs(3854) <= (layer0_outputs(1082)) xor (layer0_outputs(6545));
    outputs(3855) <= not(layer0_outputs(3356));
    outputs(3856) <= (layer0_outputs(1993)) and (layer0_outputs(7252));
    outputs(3857) <= not(layer0_outputs(7379));
    outputs(3858) <= not(layer0_outputs(4633));
    outputs(3859) <= (layer0_outputs(3733)) xor (layer0_outputs(5096));
    outputs(3860) <= layer0_outputs(173);
    outputs(3861) <= (layer0_outputs(932)) and (layer0_outputs(3709));
    outputs(3862) <= (layer0_outputs(1593)) and (layer0_outputs(5911));
    outputs(3863) <= not((layer0_outputs(4156)) xor (layer0_outputs(643)));
    outputs(3864) <= not(layer0_outputs(5611));
    outputs(3865) <= not((layer0_outputs(600)) xor (layer0_outputs(4101)));
    outputs(3866) <= layer0_outputs(1854);
    outputs(3867) <= not((layer0_outputs(5282)) xor (layer0_outputs(3606)));
    outputs(3868) <= (layer0_outputs(5999)) xor (layer0_outputs(703));
    outputs(3869) <= (layer0_outputs(7172)) and not (layer0_outputs(3619));
    outputs(3870) <= not(layer0_outputs(1620)) or (layer0_outputs(4571));
    outputs(3871) <= layer0_outputs(1975);
    outputs(3872) <= (layer0_outputs(4549)) and (layer0_outputs(53));
    outputs(3873) <= layer0_outputs(2431);
    outputs(3874) <= (layer0_outputs(6968)) xor (layer0_outputs(1076));
    outputs(3875) <= (layer0_outputs(2483)) and not (layer0_outputs(2248));
    outputs(3876) <= not(layer0_outputs(4820));
    outputs(3877) <= (layer0_outputs(6611)) and (layer0_outputs(4916));
    outputs(3878) <= not((layer0_outputs(5043)) xor (layer0_outputs(443)));
    outputs(3879) <= (layer0_outputs(6233)) and (layer0_outputs(6195));
    outputs(3880) <= layer0_outputs(2560);
    outputs(3881) <= (layer0_outputs(6023)) and not (layer0_outputs(2360));
    outputs(3882) <= not((layer0_outputs(3683)) or (layer0_outputs(5960)));
    outputs(3883) <= not((layer0_outputs(5513)) and (layer0_outputs(6072)));
    outputs(3884) <= (layer0_outputs(4962)) and not (layer0_outputs(5518));
    outputs(3885) <= layer0_outputs(6415);
    outputs(3886) <= not((layer0_outputs(804)) xor (layer0_outputs(7490)));
    outputs(3887) <= not(layer0_outputs(4780));
    outputs(3888) <= (layer0_outputs(6033)) xor (layer0_outputs(817));
    outputs(3889) <= (layer0_outputs(1629)) xor (layer0_outputs(2244));
    outputs(3890) <= not(layer0_outputs(964));
    outputs(3891) <= not((layer0_outputs(640)) xor (layer0_outputs(5997)));
    outputs(3892) <= layer0_outputs(1697);
    outputs(3893) <= not(layer0_outputs(7435));
    outputs(3894) <= not((layer0_outputs(576)) xor (layer0_outputs(3142)));
    outputs(3895) <= (layer0_outputs(2876)) xor (layer0_outputs(5392));
    outputs(3896) <= not((layer0_outputs(5572)) xor (layer0_outputs(6005)));
    outputs(3897) <= not(layer0_outputs(922));
    outputs(3898) <= not((layer0_outputs(5879)) xor (layer0_outputs(1523)));
    outputs(3899) <= not(layer0_outputs(1087));
    outputs(3900) <= layer0_outputs(5086);
    outputs(3901) <= layer0_outputs(2510);
    outputs(3902) <= layer0_outputs(3207);
    outputs(3903) <= (layer0_outputs(1476)) and not (layer0_outputs(6391));
    outputs(3904) <= not((layer0_outputs(4741)) xor (layer0_outputs(6555)));
    outputs(3905) <= not(layer0_outputs(6336));
    outputs(3906) <= not((layer0_outputs(746)) or (layer0_outputs(3701)));
    outputs(3907) <= not((layer0_outputs(5269)) xor (layer0_outputs(6358)));
    outputs(3908) <= not((layer0_outputs(5497)) and (layer0_outputs(1305)));
    outputs(3909) <= not(layer0_outputs(5126));
    outputs(3910) <= not(layer0_outputs(7002));
    outputs(3911) <= not((layer0_outputs(7527)) xor (layer0_outputs(2154)));
    outputs(3912) <= layer0_outputs(3827);
    outputs(3913) <= layer0_outputs(5425);
    outputs(3914) <= layer0_outputs(6403);
    outputs(3915) <= not((layer0_outputs(2232)) or (layer0_outputs(930)));
    outputs(3916) <= not(layer0_outputs(7042));
    outputs(3917) <= layer0_outputs(456);
    outputs(3918) <= not((layer0_outputs(4540)) xor (layer0_outputs(7372)));
    outputs(3919) <= (layer0_outputs(562)) xor (layer0_outputs(7663));
    outputs(3920) <= not(layer0_outputs(2410));
    outputs(3921) <= layer0_outputs(5330);
    outputs(3922) <= not(layer0_outputs(6519));
    outputs(3923) <= (layer0_outputs(2512)) and (layer0_outputs(2313));
    outputs(3924) <= layer0_outputs(641);
    outputs(3925) <= not((layer0_outputs(1665)) xor (layer0_outputs(3061)));
    outputs(3926) <= (layer0_outputs(1326)) and (layer0_outputs(806));
    outputs(3927) <= not((layer0_outputs(1225)) or (layer0_outputs(3301)));
    outputs(3928) <= not((layer0_outputs(4674)) xor (layer0_outputs(2984)));
    outputs(3929) <= layer0_outputs(5332);
    outputs(3930) <= (layer0_outputs(2592)) and (layer0_outputs(946));
    outputs(3931) <= (layer0_outputs(2568)) xor (layer0_outputs(7560));
    outputs(3932) <= not((layer0_outputs(4050)) or (layer0_outputs(4737)));
    outputs(3933) <= layer0_outputs(4750);
    outputs(3934) <= not(layer0_outputs(3663)) or (layer0_outputs(1268));
    outputs(3935) <= (layer0_outputs(1980)) and (layer0_outputs(4051));
    outputs(3936) <= not(layer0_outputs(4626));
    outputs(3937) <= not(layer0_outputs(1207));
    outputs(3938) <= layer0_outputs(702);
    outputs(3939) <= not(layer0_outputs(6545)) or (layer0_outputs(4611));
    outputs(3940) <= layer0_outputs(2802);
    outputs(3941) <= not((layer0_outputs(4202)) xor (layer0_outputs(6373)));
    outputs(3942) <= (layer0_outputs(6061)) xor (layer0_outputs(6193));
    outputs(3943) <= not(layer0_outputs(7633)) or (layer0_outputs(1559));
    outputs(3944) <= (layer0_outputs(5519)) and not (layer0_outputs(248));
    outputs(3945) <= not(layer0_outputs(1942));
    outputs(3946) <= not(layer0_outputs(6306));
    outputs(3947) <= not(layer0_outputs(3871));
    outputs(3948) <= (layer0_outputs(4303)) and (layer0_outputs(6901));
    outputs(3949) <= layer0_outputs(3385);
    outputs(3950) <= not(layer0_outputs(2437));
    outputs(3951) <= not(layer0_outputs(828));
    outputs(3952) <= not(layer0_outputs(5211)) or (layer0_outputs(115));
    outputs(3953) <= (layer0_outputs(896)) xor (layer0_outputs(5966));
    outputs(3954) <= (layer0_outputs(4339)) xor (layer0_outputs(5848));
    outputs(3955) <= not((layer0_outputs(3643)) or (layer0_outputs(4336)));
    outputs(3956) <= not(layer0_outputs(6944));
    outputs(3957) <= (layer0_outputs(6573)) or (layer0_outputs(1501));
    outputs(3958) <= not((layer0_outputs(406)) xor (layer0_outputs(5813)));
    outputs(3959) <= layer0_outputs(6885);
    outputs(3960) <= (layer0_outputs(5329)) xor (layer0_outputs(4591));
    outputs(3961) <= not(layer0_outputs(3722));
    outputs(3962) <= not(layer0_outputs(2314));
    outputs(3963) <= not(layer0_outputs(395));
    outputs(3964) <= layer0_outputs(2530);
    outputs(3965) <= not(layer0_outputs(1144));
    outputs(3966) <= not((layer0_outputs(91)) or (layer0_outputs(3632)));
    outputs(3967) <= (layer0_outputs(3369)) xor (layer0_outputs(5361));
    outputs(3968) <= (layer0_outputs(1591)) xor (layer0_outputs(4502));
    outputs(3969) <= (layer0_outputs(6645)) and not (layer0_outputs(6324));
    outputs(3970) <= (layer0_outputs(7550)) xor (layer0_outputs(5017));
    outputs(3971) <= (layer0_outputs(6065)) and (layer0_outputs(3435));
    outputs(3972) <= not((layer0_outputs(2362)) xor (layer0_outputs(2548)));
    outputs(3973) <= layer0_outputs(6850);
    outputs(3974) <= layer0_outputs(4835);
    outputs(3975) <= layer0_outputs(2922);
    outputs(3976) <= (layer0_outputs(7517)) and (layer0_outputs(6434));
    outputs(3977) <= not(layer0_outputs(653));
    outputs(3978) <= layer0_outputs(7186);
    outputs(3979) <= not((layer0_outputs(4278)) xor (layer0_outputs(6150)));
    outputs(3980) <= (layer0_outputs(5026)) xor (layer0_outputs(3864));
    outputs(3981) <= not(layer0_outputs(1460)) or (layer0_outputs(413));
    outputs(3982) <= layer0_outputs(2965);
    outputs(3983) <= layer0_outputs(1555);
    outputs(3984) <= not(layer0_outputs(5300));
    outputs(3985) <= not(layer0_outputs(587));
    outputs(3986) <= layer0_outputs(6548);
    outputs(3987) <= (layer0_outputs(1712)) xor (layer0_outputs(511));
    outputs(3988) <= not(layer0_outputs(7239));
    outputs(3989) <= (layer0_outputs(885)) xor (layer0_outputs(29));
    outputs(3990) <= layer0_outputs(4762);
    outputs(3991) <= layer0_outputs(2215);
    outputs(3992) <= (layer0_outputs(7342)) xor (layer0_outputs(4805));
    outputs(3993) <= not(layer0_outputs(2525));
    outputs(3994) <= (layer0_outputs(3327)) xor (layer0_outputs(4443));
    outputs(3995) <= not(layer0_outputs(1891));
    outputs(3996) <= not((layer0_outputs(4070)) xor (layer0_outputs(1339)));
    outputs(3997) <= not((layer0_outputs(2724)) xor (layer0_outputs(3591)));
    outputs(3998) <= not(layer0_outputs(1299)) or (layer0_outputs(3010));
    outputs(3999) <= not((layer0_outputs(6983)) xor (layer0_outputs(4923)));
    outputs(4000) <= not(layer0_outputs(5497));
    outputs(4001) <= not((layer0_outputs(4740)) or (layer0_outputs(7615)));
    outputs(4002) <= not(layer0_outputs(2570));
    outputs(4003) <= (layer0_outputs(1915)) or (layer0_outputs(6894));
    outputs(4004) <= not(layer0_outputs(5343));
    outputs(4005) <= (layer0_outputs(4976)) xor (layer0_outputs(2213));
    outputs(4006) <= not((layer0_outputs(3939)) xor (layer0_outputs(3673)));
    outputs(4007) <= (layer0_outputs(3918)) and not (layer0_outputs(965));
    outputs(4008) <= (layer0_outputs(1404)) and not (layer0_outputs(217));
    outputs(4009) <= layer0_outputs(351);
    outputs(4010) <= not((layer0_outputs(1072)) or (layer0_outputs(3119)));
    outputs(4011) <= layer0_outputs(7123);
    outputs(4012) <= not((layer0_outputs(7230)) xor (layer0_outputs(2851)));
    outputs(4013) <= (layer0_outputs(3709)) and (layer0_outputs(6903));
    outputs(4014) <= not(layer0_outputs(5856));
    outputs(4015) <= (layer0_outputs(6046)) xor (layer0_outputs(6218));
    outputs(4016) <= (layer0_outputs(4011)) xor (layer0_outputs(4954));
    outputs(4017) <= layer0_outputs(6859);
    outputs(4018) <= (layer0_outputs(1224)) or (layer0_outputs(3057));
    outputs(4019) <= (layer0_outputs(2741)) xor (layer0_outputs(1638));
    outputs(4020) <= layer0_outputs(3273);
    outputs(4021) <= not(layer0_outputs(6474));
    outputs(4022) <= not(layer0_outputs(875)) or (layer0_outputs(3430));
    outputs(4023) <= not((layer0_outputs(5336)) xor (layer0_outputs(3963)));
    outputs(4024) <= layer0_outputs(5080);
    outputs(4025) <= layer0_outputs(4232);
    outputs(4026) <= not((layer0_outputs(644)) xor (layer0_outputs(4277)));
    outputs(4027) <= not((layer0_outputs(3052)) xor (layer0_outputs(361)));
    outputs(4028) <= layer0_outputs(2363);
    outputs(4029) <= not(layer0_outputs(5833));
    outputs(4030) <= (layer0_outputs(5050)) and not (layer0_outputs(3531));
    outputs(4031) <= layer0_outputs(5795);
    outputs(4032) <= not(layer0_outputs(1179));
    outputs(4033) <= not(layer0_outputs(2321));
    outputs(4034) <= layer0_outputs(5813);
    outputs(4035) <= layer0_outputs(5633);
    outputs(4036) <= (layer0_outputs(5496)) or (layer0_outputs(6129));
    outputs(4037) <= not((layer0_outputs(5872)) xor (layer0_outputs(1400)));
    outputs(4038) <= layer0_outputs(971);
    outputs(4039) <= not((layer0_outputs(1745)) or (layer0_outputs(2729)));
    outputs(4040) <= not((layer0_outputs(5248)) xor (layer0_outputs(81)));
    outputs(4041) <= layer0_outputs(697);
    outputs(4042) <= not((layer0_outputs(1338)) xor (layer0_outputs(6485)));
    outputs(4043) <= not((layer0_outputs(4315)) or (layer0_outputs(3444)));
    outputs(4044) <= layer0_outputs(3010);
    outputs(4045) <= layer0_outputs(274);
    outputs(4046) <= not(layer0_outputs(1392));
    outputs(4047) <= not((layer0_outputs(3476)) xor (layer0_outputs(3508)));
    outputs(4048) <= not((layer0_outputs(7085)) xor (layer0_outputs(4569)));
    outputs(4049) <= not((layer0_outputs(4560)) xor (layer0_outputs(5244)));
    outputs(4050) <= layer0_outputs(7041);
    outputs(4051) <= layer0_outputs(2212);
    outputs(4052) <= not(layer0_outputs(7212)) or (layer0_outputs(4774));
    outputs(4053) <= not(layer0_outputs(7443));
    outputs(4054) <= not(layer0_outputs(503)) or (layer0_outputs(7102));
    outputs(4055) <= not((layer0_outputs(1827)) xor (layer0_outputs(2419)));
    outputs(4056) <= layer0_outputs(3078);
    outputs(4057) <= not(layer0_outputs(255));
    outputs(4058) <= not(layer0_outputs(1587));
    outputs(4059) <= layer0_outputs(1985);
    outputs(4060) <= not((layer0_outputs(236)) xor (layer0_outputs(515)));
    outputs(4061) <= (layer0_outputs(6717)) and not (layer0_outputs(6738));
    outputs(4062) <= not(layer0_outputs(5567)) or (layer0_outputs(4426));
    outputs(4063) <= (layer0_outputs(3681)) and not (layer0_outputs(7003));
    outputs(4064) <= not(layer0_outputs(2604));
    outputs(4065) <= not((layer0_outputs(6152)) xor (layer0_outputs(4490)));
    outputs(4066) <= layer0_outputs(3893);
    outputs(4067) <= layer0_outputs(5690);
    outputs(4068) <= (layer0_outputs(599)) xor (layer0_outputs(4831));
    outputs(4069) <= (layer0_outputs(5121)) or (layer0_outputs(2749));
    outputs(4070) <= layer0_outputs(3595);
    outputs(4071) <= (layer0_outputs(1050)) and (layer0_outputs(1694));
    outputs(4072) <= not((layer0_outputs(7306)) xor (layer0_outputs(5823)));
    outputs(4073) <= layer0_outputs(3519);
    outputs(4074) <= not((layer0_outputs(212)) xor (layer0_outputs(7439)));
    outputs(4075) <= not(layer0_outputs(4705)) or (layer0_outputs(3898));
    outputs(4076) <= layer0_outputs(798);
    outputs(4077) <= layer0_outputs(3524);
    outputs(4078) <= layer0_outputs(1259);
    outputs(4079) <= not((layer0_outputs(77)) xor (layer0_outputs(267)));
    outputs(4080) <= (layer0_outputs(5162)) or (layer0_outputs(1456));
    outputs(4081) <= not((layer0_outputs(7495)) and (layer0_outputs(1613)));
    outputs(4082) <= (layer0_outputs(2320)) and not (layer0_outputs(2048));
    outputs(4083) <= layer0_outputs(6345);
    outputs(4084) <= not(layer0_outputs(994));
    outputs(4085) <= layer0_outputs(7186);
    outputs(4086) <= layer0_outputs(2498);
    outputs(4087) <= (layer0_outputs(3151)) xor (layer0_outputs(2156));
    outputs(4088) <= layer0_outputs(2145);
    outputs(4089) <= not((layer0_outputs(4975)) and (layer0_outputs(1837)));
    outputs(4090) <= (layer0_outputs(7115)) xor (layer0_outputs(5746));
    outputs(4091) <= layer0_outputs(6475);
    outputs(4092) <= (layer0_outputs(6096)) and not (layer0_outputs(1704));
    outputs(4093) <= (layer0_outputs(147)) xor (layer0_outputs(3129));
    outputs(4094) <= layer0_outputs(510);
    outputs(4095) <= layer0_outputs(3046);
    outputs(4096) <= not((layer0_outputs(6131)) xor (layer0_outputs(1991)));
    outputs(4097) <= not((layer0_outputs(3152)) xor (layer0_outputs(0)));
    outputs(4098) <= (layer0_outputs(876)) and not (layer0_outputs(638));
    outputs(4099) <= (layer0_outputs(6222)) xor (layer0_outputs(4573));
    outputs(4100) <= not((layer0_outputs(5472)) xor (layer0_outputs(6217)));
    outputs(4101) <= (layer0_outputs(2362)) xor (layer0_outputs(4557));
    outputs(4102) <= layer0_outputs(5841);
    outputs(4103) <= not(layer0_outputs(7593));
    outputs(4104) <= (layer0_outputs(5934)) and not (layer0_outputs(255));
    outputs(4105) <= (layer0_outputs(7478)) or (layer0_outputs(6748));
    outputs(4106) <= not((layer0_outputs(6027)) xor (layer0_outputs(1499)));
    outputs(4107) <= not(layer0_outputs(3500)) or (layer0_outputs(2638));
    outputs(4108) <= not(layer0_outputs(1986)) or (layer0_outputs(2176));
    outputs(4109) <= layer0_outputs(163);
    outputs(4110) <= not(layer0_outputs(1041));
    outputs(4111) <= layer0_outputs(3020);
    outputs(4112) <= not((layer0_outputs(2391)) and (layer0_outputs(7678)));
    outputs(4113) <= layer0_outputs(7171);
    outputs(4114) <= not(layer0_outputs(1430));
    outputs(4115) <= not((layer0_outputs(1685)) and (layer0_outputs(1647)));
    outputs(4116) <= (layer0_outputs(2666)) xor (layer0_outputs(5141));
    outputs(4117) <= layer0_outputs(4378);
    outputs(4118) <= (layer0_outputs(6086)) xor (layer0_outputs(6445));
    outputs(4119) <= not(layer0_outputs(7131)) or (layer0_outputs(4312));
    outputs(4120) <= not((layer0_outputs(5127)) xor (layer0_outputs(797)));
    outputs(4121) <= layer0_outputs(5430);
    outputs(4122) <= not(layer0_outputs(2719));
    outputs(4123) <= not(layer0_outputs(2160)) or (layer0_outputs(881));
    outputs(4124) <= not(layer0_outputs(1410));
    outputs(4125) <= not(layer0_outputs(1936)) or (layer0_outputs(3592));
    outputs(4126) <= not(layer0_outputs(1215));
    outputs(4127) <= layer0_outputs(983);
    outputs(4128) <= (layer0_outputs(7188)) xor (layer0_outputs(2707));
    outputs(4129) <= not((layer0_outputs(6653)) xor (layer0_outputs(5873)));
    outputs(4130) <= not(layer0_outputs(1573)) or (layer0_outputs(3336));
    outputs(4131) <= not((layer0_outputs(4907)) or (layer0_outputs(1459)));
    outputs(4132) <= not(layer0_outputs(66)) or (layer0_outputs(260));
    outputs(4133) <= layer0_outputs(5572);
    outputs(4134) <= (layer0_outputs(6958)) xor (layer0_outputs(1008));
    outputs(4135) <= (layer0_outputs(5588)) and (layer0_outputs(1222));
    outputs(4136) <= not((layer0_outputs(5263)) xor (layer0_outputs(2814)));
    outputs(4137) <= (layer0_outputs(7646)) and not (layer0_outputs(4478));
    outputs(4138) <= not(layer0_outputs(3179));
    outputs(4139) <= (layer0_outputs(4328)) and (layer0_outputs(1954));
    outputs(4140) <= not((layer0_outputs(5845)) xor (layer0_outputs(4170)));
    outputs(4141) <= (layer0_outputs(113)) xor (layer0_outputs(5842));
    outputs(4142) <= layer0_outputs(1343);
    outputs(4143) <= (layer0_outputs(1851)) and not (layer0_outputs(6808));
    outputs(4144) <= (layer0_outputs(7491)) xor (layer0_outputs(6110));
    outputs(4145) <= layer0_outputs(2785);
    outputs(4146) <= not((layer0_outputs(1065)) xor (layer0_outputs(1572)));
    outputs(4147) <= not((layer0_outputs(6384)) and (layer0_outputs(4341)));
    outputs(4148) <= not((layer0_outputs(3791)) xor (layer0_outputs(6856)));
    outputs(4149) <= not(layer0_outputs(1486)) or (layer0_outputs(6076));
    outputs(4150) <= (layer0_outputs(5613)) and not (layer0_outputs(1493));
    outputs(4151) <= (layer0_outputs(6831)) and not (layer0_outputs(7677));
    outputs(4152) <= not(layer0_outputs(7200));
    outputs(4153) <= layer0_outputs(1581);
    outputs(4154) <= layer0_outputs(3150);
    outputs(4155) <= layer0_outputs(4679);
    outputs(4156) <= (layer0_outputs(4274)) xor (layer0_outputs(4181));
    outputs(4157) <= not(layer0_outputs(6480)) or (layer0_outputs(1497));
    outputs(4158) <= not((layer0_outputs(6873)) xor (layer0_outputs(2566)));
    outputs(4159) <= (layer0_outputs(4220)) xor (layer0_outputs(5395));
    outputs(4160) <= not(layer0_outputs(1741)) or (layer0_outputs(3425));
    outputs(4161) <= (layer0_outputs(2466)) and (layer0_outputs(1791));
    outputs(4162) <= not(layer0_outputs(2648));
    outputs(4163) <= layer0_outputs(6241);
    outputs(4164) <= (layer0_outputs(3292)) or (layer0_outputs(345));
    outputs(4165) <= not(layer0_outputs(6598));
    outputs(4166) <= not(layer0_outputs(5859));
    outputs(4167) <= (layer0_outputs(508)) and (layer0_outputs(6676));
    outputs(4168) <= not(layer0_outputs(6501));
    outputs(4169) <= (layer0_outputs(5655)) xor (layer0_outputs(1428));
    outputs(4170) <= (layer0_outputs(1714)) and not (layer0_outputs(523));
    outputs(4171) <= layer0_outputs(4493);
    outputs(4172) <= not(layer0_outputs(1785)) or (layer0_outputs(1491));
    outputs(4173) <= not(layer0_outputs(7470));
    outputs(4174) <= layer0_outputs(1849);
    outputs(4175) <= not(layer0_outputs(1678)) or (layer0_outputs(7203));
    outputs(4176) <= (layer0_outputs(6939)) and not (layer0_outputs(994));
    outputs(4177) <= (layer0_outputs(936)) or (layer0_outputs(3387));
    outputs(4178) <= layer0_outputs(6010);
    outputs(4179) <= not(layer0_outputs(7301));
    outputs(4180) <= (layer0_outputs(1155)) xor (layer0_outputs(2914));
    outputs(4181) <= layer0_outputs(153);
    outputs(4182) <= not(layer0_outputs(2260));
    outputs(4183) <= not((layer0_outputs(2403)) and (layer0_outputs(1467)));
    outputs(4184) <= not(layer0_outputs(6264));
    outputs(4185) <= not((layer0_outputs(845)) xor (layer0_outputs(5678)));
    outputs(4186) <= (layer0_outputs(4640)) and not (layer0_outputs(4897));
    outputs(4187) <= not((layer0_outputs(4449)) xor (layer0_outputs(2005)));
    outputs(4188) <= not((layer0_outputs(6893)) xor (layer0_outputs(4481)));
    outputs(4189) <= (layer0_outputs(2003)) xor (layer0_outputs(866));
    outputs(4190) <= (layer0_outputs(6845)) and not (layer0_outputs(3190));
    outputs(4191) <= not(layer0_outputs(6900));
    outputs(4192) <= (layer0_outputs(4287)) and (layer0_outputs(6526));
    outputs(4193) <= (layer0_outputs(909)) and (layer0_outputs(1637));
    outputs(4194) <= (layer0_outputs(5509)) and (layer0_outputs(1053));
    outputs(4195) <= (layer0_outputs(3477)) or (layer0_outputs(2291));
    outputs(4196) <= (layer0_outputs(2163)) xor (layer0_outputs(6634));
    outputs(4197) <= not((layer0_outputs(4838)) xor (layer0_outputs(6484)));
    outputs(4198) <= not(layer0_outputs(1565));
    outputs(4199) <= not(layer0_outputs(3856));
    outputs(4200) <= (layer0_outputs(6279)) xor (layer0_outputs(3232));
    outputs(4201) <= (layer0_outputs(6812)) xor (layer0_outputs(6898));
    outputs(4202) <= not(layer0_outputs(3749)) or (layer0_outputs(3506));
    outputs(4203) <= (layer0_outputs(6240)) xor (layer0_outputs(6268));
    outputs(4204) <= layer0_outputs(1086);
    outputs(4205) <= not(layer0_outputs(6814));
    outputs(4206) <= (layer0_outputs(3372)) xor (layer0_outputs(3308));
    outputs(4207) <= layer0_outputs(4603);
    outputs(4208) <= layer0_outputs(5276);
    outputs(4209) <= not((layer0_outputs(7272)) xor (layer0_outputs(6208)));
    outputs(4210) <= (layer0_outputs(5984)) xor (layer0_outputs(4616));
    outputs(4211) <= not(layer0_outputs(7191));
    outputs(4212) <= not(layer0_outputs(1925));
    outputs(4213) <= (layer0_outputs(1636)) and (layer0_outputs(6863));
    outputs(4214) <= (layer0_outputs(743)) xor (layer0_outputs(4579));
    outputs(4215) <= not(layer0_outputs(2890));
    outputs(4216) <= (layer0_outputs(3134)) and not (layer0_outputs(4229));
    outputs(4217) <= (layer0_outputs(3844)) xor (layer0_outputs(5501));
    outputs(4218) <= not((layer0_outputs(1728)) and (layer0_outputs(2706)));
    outputs(4219) <= not((layer0_outputs(1458)) xor (layer0_outputs(2766)));
    outputs(4220) <= (layer0_outputs(3212)) and not (layer0_outputs(6461));
    outputs(4221) <= (layer0_outputs(6035)) and not (layer0_outputs(2248));
    outputs(4222) <= layer0_outputs(1816);
    outputs(4223) <= (layer0_outputs(2044)) and not (layer0_outputs(6786));
    outputs(4224) <= not((layer0_outputs(4367)) or (layer0_outputs(2688)));
    outputs(4225) <= layer0_outputs(6204);
    outputs(4226) <= not((layer0_outputs(5221)) xor (layer0_outputs(6612)));
    outputs(4227) <= (layer0_outputs(2405)) and not (layer0_outputs(3133));
    outputs(4228) <= (layer0_outputs(3436)) xor (layer0_outputs(4918));
    outputs(4229) <= layer0_outputs(1448);
    outputs(4230) <= layer0_outputs(4784);
    outputs(4231) <= not((layer0_outputs(1301)) xor (layer0_outputs(2122)));
    outputs(4232) <= not(layer0_outputs(7619));
    outputs(4233) <= not((layer0_outputs(6941)) xor (layer0_outputs(6760)));
    outputs(4234) <= not((layer0_outputs(6055)) xor (layer0_outputs(177)));
    outputs(4235) <= not((layer0_outputs(2288)) xor (layer0_outputs(7354)));
    outputs(4236) <= not(layer0_outputs(6339)) or (layer0_outputs(2062));
    outputs(4237) <= not(layer0_outputs(6549)) or (layer0_outputs(1517));
    outputs(4238) <= not(layer0_outputs(1699)) or (layer0_outputs(160));
    outputs(4239) <= not(layer0_outputs(2480));
    outputs(4240) <= (layer0_outputs(6761)) xor (layer0_outputs(5719));
    outputs(4241) <= (layer0_outputs(1242)) and (layer0_outputs(1231));
    outputs(4242) <= (layer0_outputs(3095)) and (layer0_outputs(6431));
    outputs(4243) <= not((layer0_outputs(552)) xor (layer0_outputs(6890)));
    outputs(4244) <= (layer0_outputs(5777)) and (layer0_outputs(7366));
    outputs(4245) <= layer0_outputs(6952);
    outputs(4246) <= layer0_outputs(4850);
    outputs(4247) <= layer0_outputs(6357);
    outputs(4248) <= (layer0_outputs(137)) xor (layer0_outputs(2768));
    outputs(4249) <= not((layer0_outputs(3910)) xor (layer0_outputs(4918)));
    outputs(4250) <= (layer0_outputs(1748)) and not (layer0_outputs(7099));
    outputs(4251) <= not((layer0_outputs(3798)) or (layer0_outputs(2624)));
    outputs(4252) <= not(layer0_outputs(5139)) or (layer0_outputs(4022));
    outputs(4253) <= not((layer0_outputs(7070)) xor (layer0_outputs(5181)));
    outputs(4254) <= not(layer0_outputs(4621));
    outputs(4255) <= layer0_outputs(3640);
    outputs(4256) <= not((layer0_outputs(4093)) xor (layer0_outputs(2253)));
    outputs(4257) <= not((layer0_outputs(2268)) and (layer0_outputs(5087)));
    outputs(4258) <= layer0_outputs(4738);
    outputs(4259) <= not(layer0_outputs(6375)) or (layer0_outputs(148));
    outputs(4260) <= (layer0_outputs(819)) or (layer0_outputs(6133));
    outputs(4261) <= not(layer0_outputs(4342)) or (layer0_outputs(3879));
    outputs(4262) <= (layer0_outputs(2576)) xor (layer0_outputs(6538));
    outputs(4263) <= not(layer0_outputs(2025));
    outputs(4264) <= (layer0_outputs(1651)) and not (layer0_outputs(1304));
    outputs(4265) <= (layer0_outputs(3069)) and not (layer0_outputs(6664));
    outputs(4266) <= (layer0_outputs(3021)) and not (layer0_outputs(1866));
    outputs(4267) <= layer0_outputs(4783);
    outputs(4268) <= (layer0_outputs(6768)) and (layer0_outputs(7010));
    outputs(4269) <= layer0_outputs(4457);
    outputs(4270) <= not(layer0_outputs(2383));
    outputs(4271) <= layer0_outputs(4625);
    outputs(4272) <= (layer0_outputs(3981)) xor (layer0_outputs(6564));
    outputs(4273) <= layer0_outputs(2508);
    outputs(4274) <= layer0_outputs(2297);
    outputs(4275) <= not(layer0_outputs(6598));
    outputs(4276) <= layer0_outputs(2024);
    outputs(4277) <= not((layer0_outputs(5679)) xor (layer0_outputs(3855)));
    outputs(4278) <= (layer0_outputs(3544)) and not (layer0_outputs(2800));
    outputs(4279) <= not(layer0_outputs(6049));
    outputs(4280) <= not((layer0_outputs(7592)) xor (layer0_outputs(4649)));
    outputs(4281) <= layer0_outputs(767);
    outputs(4282) <= layer0_outputs(4022);
    outputs(4283) <= not(layer0_outputs(613));
    outputs(4284) <= layer0_outputs(6608);
    outputs(4285) <= not(layer0_outputs(3535));
    outputs(4286) <= layer0_outputs(6729);
    outputs(4287) <= (layer0_outputs(1414)) xor (layer0_outputs(4379));
    outputs(4288) <= not(layer0_outputs(3158));
    outputs(4289) <= (layer0_outputs(7069)) and not (layer0_outputs(208));
    outputs(4290) <= not((layer0_outputs(4126)) xor (layer0_outputs(6109)));
    outputs(4291) <= not(layer0_outputs(4904));
    outputs(4292) <= not((layer0_outputs(1865)) or (layer0_outputs(7458)));
    outputs(4293) <= (layer0_outputs(3728)) xor (layer0_outputs(2241));
    outputs(4294) <= layer0_outputs(5834);
    outputs(4295) <= layer0_outputs(6952);
    outputs(4296) <= not((layer0_outputs(1528)) and (layer0_outputs(6003)));
    outputs(4297) <= not((layer0_outputs(4332)) xor (layer0_outputs(3766)));
    outputs(4298) <= (layer0_outputs(4219)) and not (layer0_outputs(4752));
    outputs(4299) <= layer0_outputs(2052);
    outputs(4300) <= not((layer0_outputs(6421)) xor (layer0_outputs(2214)));
    outputs(4301) <= layer0_outputs(5133);
    outputs(4302) <= not((layer0_outputs(5066)) xor (layer0_outputs(169)));
    outputs(4303) <= layer0_outputs(7394);
    outputs(4304) <= (layer0_outputs(7271)) and not (layer0_outputs(5303));
    outputs(4305) <= layer0_outputs(1977);
    outputs(4306) <= layer0_outputs(1520);
    outputs(4307) <= not(layer0_outputs(5779));
    outputs(4308) <= not(layer0_outputs(4032));
    outputs(4309) <= layer0_outputs(7106);
    outputs(4310) <= (layer0_outputs(7023)) xor (layer0_outputs(3732));
    outputs(4311) <= not(layer0_outputs(6837));
    outputs(4312) <= (layer0_outputs(6160)) or (layer0_outputs(2886));
    outputs(4313) <= layer0_outputs(109);
    outputs(4314) <= layer0_outputs(5942);
    outputs(4315) <= layer0_outputs(1519);
    outputs(4316) <= (layer0_outputs(2636)) xor (layer0_outputs(2359));
    outputs(4317) <= not((layer0_outputs(4778)) xor (layer0_outputs(5218)));
    outputs(4318) <= layer0_outputs(1262);
    outputs(4319) <= layer0_outputs(1749);
    outputs(4320) <= (layer0_outputs(7029)) xor (layer0_outputs(4422));
    outputs(4321) <= layer0_outputs(6330);
    outputs(4322) <= layer0_outputs(6262);
    outputs(4323) <= (layer0_outputs(6468)) xor (layer0_outputs(6787));
    outputs(4324) <= (layer0_outputs(5589)) xor (layer0_outputs(5444));
    outputs(4325) <= layer0_outputs(1330);
    outputs(4326) <= (layer0_outputs(2759)) xor (layer0_outputs(507));
    outputs(4327) <= layer0_outputs(2060);
    outputs(4328) <= not(layer0_outputs(5272));
    outputs(4329) <= not(layer0_outputs(5090));
    outputs(4330) <= (layer0_outputs(1853)) and not (layer0_outputs(7196));
    outputs(4331) <= (layer0_outputs(2671)) and not (layer0_outputs(124));
    outputs(4332) <= (layer0_outputs(541)) and (layer0_outputs(6930));
    outputs(4333) <= layer0_outputs(3605);
    outputs(4334) <= (layer0_outputs(3210)) and not (layer0_outputs(2698));
    outputs(4335) <= not(layer0_outputs(5200));
    outputs(4336) <= not((layer0_outputs(1932)) and (layer0_outputs(6660)));
    outputs(4337) <= not(layer0_outputs(967));
    outputs(4338) <= not((layer0_outputs(5103)) and (layer0_outputs(6444)));
    outputs(4339) <= not((layer0_outputs(422)) and (layer0_outputs(7594)));
    outputs(4340) <= not(layer0_outputs(4010));
    outputs(4341) <= layer0_outputs(1831);
    outputs(4342) <= not((layer0_outputs(2048)) or (layer0_outputs(4680)));
    outputs(4343) <= not((layer0_outputs(4975)) and (layer0_outputs(5683)));
    outputs(4344) <= not((layer0_outputs(1635)) xor (layer0_outputs(6945)));
    outputs(4345) <= not(layer0_outputs(259)) or (layer0_outputs(4054));
    outputs(4346) <= not((layer0_outputs(4778)) and (layer0_outputs(1076)));
    outputs(4347) <= not((layer0_outputs(3872)) xor (layer0_outputs(765)));
    outputs(4348) <= not((layer0_outputs(7397)) xor (layer0_outputs(5958)));
    outputs(4349) <= not(layer0_outputs(5616));
    outputs(4350) <= not(layer0_outputs(695));
    outputs(4351) <= (layer0_outputs(7109)) xor (layer0_outputs(3058));
    outputs(4352) <= not((layer0_outputs(1488)) xor (layer0_outputs(1794)));
    outputs(4353) <= not((layer0_outputs(938)) xor (layer0_outputs(1857)));
    outputs(4354) <= layer0_outputs(5500);
    outputs(4355) <= (layer0_outputs(830)) xor (layer0_outputs(5042));
    outputs(4356) <= (layer0_outputs(7283)) xor (layer0_outputs(3953));
    outputs(4357) <= (layer0_outputs(2291)) and not (layer0_outputs(3533));
    outputs(4358) <= not((layer0_outputs(6785)) or (layer0_outputs(1764)));
    outputs(4359) <= (layer0_outputs(3253)) and not (layer0_outputs(904));
    outputs(4360) <= not((layer0_outputs(2609)) xor (layer0_outputs(3112)));
    outputs(4361) <= not((layer0_outputs(6311)) xor (layer0_outputs(1357)));
    outputs(4362) <= not((layer0_outputs(7383)) and (layer0_outputs(1111)));
    outputs(4363) <= not((layer0_outputs(7595)) and (layer0_outputs(3654)));
    outputs(4364) <= layer0_outputs(4127);
    outputs(4365) <= not(layer0_outputs(5723));
    outputs(4366) <= (layer0_outputs(41)) and not (layer0_outputs(5828));
    outputs(4367) <= (layer0_outputs(6782)) xor (layer0_outputs(6491));
    outputs(4368) <= not(layer0_outputs(3734));
    outputs(4369) <= not(layer0_outputs(4039));
    outputs(4370) <= layer0_outputs(2807);
    outputs(4371) <= not((layer0_outputs(6963)) xor (layer0_outputs(2299)));
    outputs(4372) <= not((layer0_outputs(2367)) xor (layer0_outputs(6511)));
    outputs(4373) <= not((layer0_outputs(2613)) or (layer0_outputs(6714)));
    outputs(4374) <= not((layer0_outputs(4144)) xor (layer0_outputs(3441)));
    outputs(4375) <= not(layer0_outputs(1715));
    outputs(4376) <= not(layer0_outputs(5159));
    outputs(4377) <= not(layer0_outputs(6000));
    outputs(4378) <= (layer0_outputs(7373)) xor (layer0_outputs(5225));
    outputs(4379) <= not((layer0_outputs(5918)) xor (layer0_outputs(6642)));
    outputs(4380) <= not(layer0_outputs(6489)) or (layer0_outputs(7500));
    outputs(4381) <= not(layer0_outputs(1922));
    outputs(4382) <= not((layer0_outputs(4422)) xor (layer0_outputs(2455)));
    outputs(4383) <= layer0_outputs(4433);
    outputs(4384) <= not(layer0_outputs(1544));
    outputs(4385) <= not(layer0_outputs(7536)) or (layer0_outputs(1523));
    outputs(4386) <= not(layer0_outputs(5402));
    outputs(4387) <= layer0_outputs(4334);
    outputs(4388) <= layer0_outputs(7668);
    outputs(4389) <= layer0_outputs(2497);
    outputs(4390) <= layer0_outputs(3377);
    outputs(4391) <= layer0_outputs(6684);
    outputs(4392) <= not((layer0_outputs(4472)) xor (layer0_outputs(6428)));
    outputs(4393) <= not((layer0_outputs(6189)) xor (layer0_outputs(1336)));
    outputs(4394) <= (layer0_outputs(7351)) or (layer0_outputs(604));
    outputs(4395) <= not((layer0_outputs(7159)) xor (layer0_outputs(4834)));
    outputs(4396) <= not((layer0_outputs(915)) xor (layer0_outputs(7293)));
    outputs(4397) <= (layer0_outputs(5531)) and not (layer0_outputs(7508));
    outputs(4398) <= layer0_outputs(5601);
    outputs(4399) <= (layer0_outputs(1066)) xor (layer0_outputs(1666));
    outputs(4400) <= (layer0_outputs(7483)) or (layer0_outputs(4294));
    outputs(4401) <= (layer0_outputs(6753)) xor (layer0_outputs(1873));
    outputs(4402) <= (layer0_outputs(6400)) xor (layer0_outputs(3070));
    outputs(4403) <= layer0_outputs(5768);
    outputs(4404) <= (layer0_outputs(63)) xor (layer0_outputs(1799));
    outputs(4405) <= not((layer0_outputs(1320)) and (layer0_outputs(5314)));
    outputs(4406) <= layer0_outputs(4926);
    outputs(4407) <= not((layer0_outputs(946)) xor (layer0_outputs(3645)));
    outputs(4408) <= not((layer0_outputs(1881)) xor (layer0_outputs(6269)));
    outputs(4409) <= (layer0_outputs(6571)) and (layer0_outputs(4470));
    outputs(4410) <= layer0_outputs(6360);
    outputs(4411) <= layer0_outputs(2907);
    outputs(4412) <= layer0_outputs(7403);
    outputs(4413) <= not(layer0_outputs(48));
    outputs(4414) <= layer0_outputs(4079);
    outputs(4415) <= not((layer0_outputs(1803)) or (layer0_outputs(2832)));
    outputs(4416) <= (layer0_outputs(487)) and not (layer0_outputs(2873));
    outputs(4417) <= not((layer0_outputs(1025)) xor (layer0_outputs(603)));
    outputs(4418) <= (layer0_outputs(7081)) and (layer0_outputs(5845));
    outputs(4419) <= (layer0_outputs(302)) xor (layer0_outputs(4526));
    outputs(4420) <= layer0_outputs(2838);
    outputs(4421) <= not((layer0_outputs(1926)) and (layer0_outputs(6604)));
    outputs(4422) <= layer0_outputs(4866);
    outputs(4423) <= not(layer0_outputs(1143)) or (layer0_outputs(4872));
    outputs(4424) <= not(layer0_outputs(5027));
    outputs(4425) <= (layer0_outputs(4876)) xor (layer0_outputs(1880));
    outputs(4426) <= (layer0_outputs(1332)) or (layer0_outputs(1758));
    outputs(4427) <= layer0_outputs(2265);
    outputs(4428) <= not((layer0_outputs(1080)) and (layer0_outputs(887)));
    outputs(4429) <= not(layer0_outputs(3933));
    outputs(4430) <= not((layer0_outputs(6090)) xor (layer0_outputs(1870)));
    outputs(4431) <= not((layer0_outputs(5194)) and (layer0_outputs(3362)));
    outputs(4432) <= not(layer0_outputs(7462));
    outputs(4433) <= not(layer0_outputs(6672)) or (layer0_outputs(6648));
    outputs(4434) <= (layer0_outputs(2305)) and (layer0_outputs(6063));
    outputs(4435) <= layer0_outputs(3959);
    outputs(4436) <= not(layer0_outputs(2012));
    outputs(4437) <= not(layer0_outputs(4435));
    outputs(4438) <= not(layer0_outputs(7600));
    outputs(4439) <= not(layer0_outputs(3328));
    outputs(4440) <= (layer0_outputs(4713)) xor (layer0_outputs(1109));
    outputs(4441) <= (layer0_outputs(7250)) and not (layer0_outputs(1415));
    outputs(4442) <= not(layer0_outputs(1924));
    outputs(4443) <= not((layer0_outputs(5824)) xor (layer0_outputs(1350)));
    outputs(4444) <= not(layer0_outputs(2606));
    outputs(4445) <= (layer0_outputs(2117)) and (layer0_outputs(4019));
    outputs(4446) <= not((layer0_outputs(7360)) xor (layer0_outputs(6685)));
    outputs(4447) <= not(layer0_outputs(6453));
    outputs(4448) <= layer0_outputs(2837);
    outputs(4449) <= not(layer0_outputs(5313)) or (layer0_outputs(5755));
    outputs(4450) <= not(layer0_outputs(7356));
    outputs(4451) <= layer0_outputs(6004);
    outputs(4452) <= layer0_outputs(324);
    outputs(4453) <= not((layer0_outputs(4673)) and (layer0_outputs(7506)));
    outputs(4454) <= layer0_outputs(6893);
    outputs(4455) <= not((layer0_outputs(662)) xor (layer0_outputs(2036)));
    outputs(4456) <= not(layer0_outputs(6362));
    outputs(4457) <= (layer0_outputs(1031)) xor (layer0_outputs(3543));
    outputs(4458) <= not(layer0_outputs(907));
    outputs(4459) <= not(layer0_outputs(5909));
    outputs(4460) <= layer0_outputs(112);
    outputs(4461) <= not((layer0_outputs(3856)) or (layer0_outputs(673)));
    outputs(4462) <= not(layer0_outputs(5206));
    outputs(4463) <= layer0_outputs(4639);
    outputs(4464) <= (layer0_outputs(1825)) xor (layer0_outputs(6265));
    outputs(4465) <= layer0_outputs(2559);
    outputs(4466) <= (layer0_outputs(5445)) and not (layer0_outputs(3369));
    outputs(4467) <= not(layer0_outputs(1148));
    outputs(4468) <= layer0_outputs(524);
    outputs(4469) <= (layer0_outputs(3828)) and not (layer0_outputs(1914));
    outputs(4470) <= (layer0_outputs(2154)) and (layer0_outputs(2148));
    outputs(4471) <= not((layer0_outputs(1776)) xor (layer0_outputs(3710)));
    outputs(4472) <= (layer0_outputs(5729)) xor (layer0_outputs(1691));
    outputs(4473) <= (layer0_outputs(1628)) and (layer0_outputs(1389));
    outputs(4474) <= layer0_outputs(4243);
    outputs(4475) <= not(layer0_outputs(4589));
    outputs(4476) <= (layer0_outputs(5780)) xor (layer0_outputs(2100));
    outputs(4477) <= not((layer0_outputs(1607)) xor (layer0_outputs(995)));
    outputs(4478) <= (layer0_outputs(4396)) xor (layer0_outputs(4913));
    outputs(4479) <= not(layer0_outputs(1141)) or (layer0_outputs(6838));
    outputs(4480) <= (layer0_outputs(5059)) xor (layer0_outputs(1869));
    outputs(4481) <= (layer0_outputs(7369)) and (layer0_outputs(240));
    outputs(4482) <= not((layer0_outputs(625)) xor (layer0_outputs(2899)));
    outputs(4483) <= not((layer0_outputs(4003)) xor (layer0_outputs(6320)));
    outputs(4484) <= (layer0_outputs(4430)) xor (layer0_outputs(3036));
    outputs(4485) <= (layer0_outputs(1298)) and not (layer0_outputs(198));
    outputs(4486) <= (layer0_outputs(4402)) xor (layer0_outputs(3699));
    outputs(4487) <= layer0_outputs(6817);
    outputs(4488) <= not(layer0_outputs(4032));
    outputs(4489) <= layer0_outputs(1667);
    outputs(4490) <= layer0_outputs(3378);
    outputs(4491) <= layer0_outputs(7574);
    outputs(4492) <= not(layer0_outputs(5002));
    outputs(4493) <= layer0_outputs(3505);
    outputs(4494) <= not(layer0_outputs(785));
    outputs(4495) <= not(layer0_outputs(462));
    outputs(4496) <= layer0_outputs(2836);
    outputs(4497) <= layer0_outputs(5041);
    outputs(4498) <= (layer0_outputs(986)) xor (layer0_outputs(3673));
    outputs(4499) <= layer0_outputs(1747);
    outputs(4500) <= layer0_outputs(3352);
    outputs(4501) <= (layer0_outputs(132)) xor (layer0_outputs(4400));
    outputs(4502) <= (layer0_outputs(4628)) and not (layer0_outputs(549));
    outputs(4503) <= not((layer0_outputs(5792)) xor (layer0_outputs(225)));
    outputs(4504) <= not(layer0_outputs(681));
    outputs(4505) <= not((layer0_outputs(3395)) xor (layer0_outputs(1808)));
    outputs(4506) <= not((layer0_outputs(2499)) and (layer0_outputs(1430)));
    outputs(4507) <= (layer0_outputs(6964)) and not (layer0_outputs(573));
    outputs(4508) <= not(layer0_outputs(2227)) or (layer0_outputs(2775));
    outputs(4509) <= not((layer0_outputs(1619)) and (layer0_outputs(3299)));
    outputs(4510) <= not((layer0_outputs(7322)) xor (layer0_outputs(4354)));
    outputs(4511) <= not(layer0_outputs(5153));
    outputs(4512) <= (layer0_outputs(3343)) and (layer0_outputs(1476));
    outputs(4513) <= not(layer0_outputs(2727));
    outputs(4514) <= not((layer0_outputs(750)) xor (layer0_outputs(2034)));
    outputs(4515) <= layer0_outputs(4671);
    outputs(4516) <= (layer0_outputs(7068)) or (layer0_outputs(3762));
    outputs(4517) <= not(layer0_outputs(2826));
    outputs(4518) <= (layer0_outputs(1262)) and (layer0_outputs(1404));
    outputs(4519) <= (layer0_outputs(921)) and not (layer0_outputs(5476));
    outputs(4520) <= (layer0_outputs(7329)) and not (layer0_outputs(955));
    outputs(4521) <= not((layer0_outputs(2139)) xor (layer0_outputs(4840)));
    outputs(4522) <= (layer0_outputs(4327)) or (layer0_outputs(2751));
    outputs(4523) <= (layer0_outputs(2223)) xor (layer0_outputs(425));
    outputs(4524) <= not(layer0_outputs(807));
    outputs(4525) <= layer0_outputs(1839);
    outputs(4526) <= not(layer0_outputs(4551));
    outputs(4527) <= not((layer0_outputs(2396)) xor (layer0_outputs(3864)));
    outputs(4528) <= not((layer0_outputs(6905)) xor (layer0_outputs(1578)));
    outputs(4529) <= (layer0_outputs(4824)) or (layer0_outputs(1320));
    outputs(4530) <= (layer0_outputs(1608)) xor (layer0_outputs(2878));
    outputs(4531) <= layer0_outputs(713);
    outputs(4532) <= (layer0_outputs(1396)) xor (layer0_outputs(5099));
    outputs(4533) <= not(layer0_outputs(4814));
    outputs(4534) <= not((layer0_outputs(6339)) and (layer0_outputs(1102)));
    outputs(4535) <= not((layer0_outputs(1586)) and (layer0_outputs(2100)));
    outputs(4536) <= not((layer0_outputs(3392)) xor (layer0_outputs(5892)));
    outputs(4537) <= not(layer0_outputs(6048)) or (layer0_outputs(3846));
    outputs(4538) <= (layer0_outputs(2583)) or (layer0_outputs(3746));
    outputs(4539) <= (layer0_outputs(5869)) and not (layer0_outputs(2832));
    outputs(4540) <= not(layer0_outputs(2280)) or (layer0_outputs(5455));
    outputs(4541) <= layer0_outputs(5084);
    outputs(4542) <= not(layer0_outputs(1803));
    outputs(4543) <= not(layer0_outputs(3514));
    outputs(4544) <= not((layer0_outputs(5986)) xor (layer0_outputs(4593)));
    outputs(4545) <= not(layer0_outputs(5963));
    outputs(4546) <= (layer0_outputs(4473)) or (layer0_outputs(5176));
    outputs(4547) <= layer0_outputs(5201);
    outputs(4548) <= layer0_outputs(2032);
    outputs(4549) <= (layer0_outputs(6063)) and not (layer0_outputs(4825));
    outputs(4550) <= not((layer0_outputs(6452)) xor (layer0_outputs(4436)));
    outputs(4551) <= not(layer0_outputs(3139)) or (layer0_outputs(342));
    outputs(4552) <= not(layer0_outputs(7572));
    outputs(4553) <= not(layer0_outputs(6906)) or (layer0_outputs(2521));
    outputs(4554) <= layer0_outputs(3959);
    outputs(4555) <= not(layer0_outputs(5778));
    outputs(4556) <= not((layer0_outputs(6902)) xor (layer0_outputs(5649)));
    outputs(4557) <= layer0_outputs(3272);
    outputs(4558) <= (layer0_outputs(3181)) xor (layer0_outputs(6681));
    outputs(4559) <= (layer0_outputs(2974)) and not (layer0_outputs(3318));
    outputs(4560) <= not(layer0_outputs(6572));
    outputs(4561) <= not(layer0_outputs(7572));
    outputs(4562) <= not((layer0_outputs(5547)) or (layer0_outputs(7650)));
    outputs(4563) <= not(layer0_outputs(4915)) or (layer0_outputs(6253));
    outputs(4564) <= not(layer0_outputs(1931)) or (layer0_outputs(4256));
    outputs(4565) <= layer0_outputs(3609);
    outputs(4566) <= not((layer0_outputs(4028)) xor (layer0_outputs(1646)));
    outputs(4567) <= (layer0_outputs(365)) or (layer0_outputs(4821));
    outputs(4568) <= (layer0_outputs(7359)) xor (layer0_outputs(1239));
    outputs(4569) <= not(layer0_outputs(6874)) or (layer0_outputs(3815));
    outputs(4570) <= layer0_outputs(6101);
    outputs(4571) <= (layer0_outputs(4597)) and not (layer0_outputs(3718));
    outputs(4572) <= (layer0_outputs(2409)) and not (layer0_outputs(6351));
    outputs(4573) <= not((layer0_outputs(7067)) xor (layer0_outputs(3013)));
    outputs(4574) <= not(layer0_outputs(5434)) or (layer0_outputs(2054));
    outputs(4575) <= (layer0_outputs(2501)) or (layer0_outputs(130));
    outputs(4576) <= not(layer0_outputs(7207));
    outputs(4577) <= not(layer0_outputs(3924)) or (layer0_outputs(6269));
    outputs(4578) <= not(layer0_outputs(5222)) or (layer0_outputs(1094));
    outputs(4579) <= layer0_outputs(4646);
    outputs(4580) <= not(layer0_outputs(7265));
    outputs(4581) <= layer0_outputs(6930);
    outputs(4582) <= (layer0_outputs(7134)) xor (layer0_outputs(1360));
    outputs(4583) <= (layer0_outputs(2568)) xor (layer0_outputs(7148));
    outputs(4584) <= not((layer0_outputs(485)) xor (layer0_outputs(5108)));
    outputs(4585) <= not(layer0_outputs(2931));
    outputs(4586) <= layer0_outputs(1963);
    outputs(4587) <= not((layer0_outputs(1946)) and (layer0_outputs(2924)));
    outputs(4588) <= not(layer0_outputs(5227));
    outputs(4589) <= (layer0_outputs(7308)) xor (layer0_outputs(2810));
    outputs(4590) <= not(layer0_outputs(7545));
    outputs(4591) <= not(layer0_outputs(1211));
    outputs(4592) <= not((layer0_outputs(6311)) xor (layer0_outputs(488)));
    outputs(4593) <= (layer0_outputs(7611)) xor (layer0_outputs(789));
    outputs(4594) <= not((layer0_outputs(2207)) or (layer0_outputs(3495)));
    outputs(4595) <= layer0_outputs(7401);
    outputs(4596) <= not(layer0_outputs(4175));
    outputs(4597) <= (layer0_outputs(5889)) xor (layer0_outputs(7482));
    outputs(4598) <= not(layer0_outputs(5049));
    outputs(4599) <= layer0_outputs(7053);
    outputs(4600) <= not((layer0_outputs(3557)) xor (layer0_outputs(6243)));
    outputs(4601) <= layer0_outputs(119);
    outputs(4602) <= not((layer0_outputs(1096)) xor (layer0_outputs(3746)));
    outputs(4603) <= not(layer0_outputs(4381));
    outputs(4604) <= layer0_outputs(5776);
    outputs(4605) <= not((layer0_outputs(1002)) xor (layer0_outputs(7396)));
    outputs(4606) <= (layer0_outputs(531)) xor (layer0_outputs(4569));
    outputs(4607) <= layer0_outputs(6650);
    outputs(4608) <= (layer0_outputs(7224)) and not (layer0_outputs(1635));
    outputs(4609) <= not((layer0_outputs(5941)) xor (layer0_outputs(2917)));
    outputs(4610) <= (layer0_outputs(3421)) or (layer0_outputs(7554));
    outputs(4611) <= (layer0_outputs(838)) and not (layer0_outputs(6400));
    outputs(4612) <= layer0_outputs(377);
    outputs(4613) <= not((layer0_outputs(1885)) or (layer0_outputs(3410)));
    outputs(4614) <= not(layer0_outputs(2731));
    outputs(4615) <= not(layer0_outputs(1759));
    outputs(4616) <= not(layer0_outputs(1801));
    outputs(4617) <= (layer0_outputs(4210)) or (layer0_outputs(3415));
    outputs(4618) <= (layer0_outputs(3209)) xor (layer0_outputs(5105));
    outputs(4619) <= not(layer0_outputs(6437));
    outputs(4620) <= layer0_outputs(1226);
    outputs(4621) <= not(layer0_outputs(3218));
    outputs(4622) <= not(layer0_outputs(6352));
    outputs(4623) <= (layer0_outputs(4876)) and not (layer0_outputs(3339));
    outputs(4624) <= not(layer0_outputs(2085));
    outputs(4625) <= (layer0_outputs(2478)) and not (layer0_outputs(6581));
    outputs(4626) <= (layer0_outputs(5335)) and (layer0_outputs(7254));
    outputs(4627) <= (layer0_outputs(1854)) and (layer0_outputs(5671));
    outputs(4628) <= (layer0_outputs(973)) and (layer0_outputs(7644));
    outputs(4629) <= layer0_outputs(55);
    outputs(4630) <= not(layer0_outputs(4669));
    outputs(4631) <= (layer0_outputs(3567)) and not (layer0_outputs(7100));
    outputs(4632) <= (layer0_outputs(3511)) and not (layer0_outputs(4155));
    outputs(4633) <= (layer0_outputs(6675)) and not (layer0_outputs(4065));
    outputs(4634) <= not(layer0_outputs(3151));
    outputs(4635) <= not(layer0_outputs(3913));
    outputs(4636) <= not(layer0_outputs(1495));
    outputs(4637) <= not(layer0_outputs(3983));
    outputs(4638) <= (layer0_outputs(2406)) xor (layer0_outputs(584));
    outputs(4639) <= not(layer0_outputs(4405));
    outputs(4640) <= layer0_outputs(7199);
    outputs(4641) <= (layer0_outputs(7299)) xor (layer0_outputs(1812));
    outputs(4642) <= (layer0_outputs(7364)) and not (layer0_outputs(4902));
    outputs(4643) <= not(layer0_outputs(6839));
    outputs(4644) <= not(layer0_outputs(1008));
    outputs(4645) <= (layer0_outputs(5782)) and not (layer0_outputs(6856));
    outputs(4646) <= layer0_outputs(5614);
    outputs(4647) <= layer0_outputs(2834);
    outputs(4648) <= not((layer0_outputs(5202)) or (layer0_outputs(5609)));
    outputs(4649) <= not(layer0_outputs(4610));
    outputs(4650) <= (layer0_outputs(7110)) and not (layer0_outputs(2277));
    outputs(4651) <= not((layer0_outputs(3326)) and (layer0_outputs(4114)));
    outputs(4652) <= (layer0_outputs(1029)) xor (layer0_outputs(31));
    outputs(4653) <= (layer0_outputs(7094)) xor (layer0_outputs(2185));
    outputs(4654) <= not(layer0_outputs(1139)) or (layer0_outputs(4319));
    outputs(4655) <= layer0_outputs(2869);
    outputs(4656) <= not(layer0_outputs(2519)) or (layer0_outputs(1056));
    outputs(4657) <= not(layer0_outputs(1215));
    outputs(4658) <= not((layer0_outputs(4541)) or (layer0_outputs(5011)));
    outputs(4659) <= (layer0_outputs(380)) xor (layer0_outputs(1097));
    outputs(4660) <= not((layer0_outputs(6663)) or (layer0_outputs(1719)));
    outputs(4661) <= layer0_outputs(7002);
    outputs(4662) <= not((layer0_outputs(469)) or (layer0_outputs(7667)));
    outputs(4663) <= not(layer0_outputs(4786)) or (layer0_outputs(7408));
    outputs(4664) <= (layer0_outputs(4661)) and not (layer0_outputs(4939));
    outputs(4665) <= not((layer0_outputs(6017)) and (layer0_outputs(3775)));
    outputs(4666) <= not((layer0_outputs(6164)) xor (layer0_outputs(2503)));
    outputs(4667) <= layer0_outputs(5106);
    outputs(4668) <= not(layer0_outputs(1237)) or (layer0_outputs(6253));
    outputs(4669) <= not(layer0_outputs(3172)) or (layer0_outputs(7477));
    outputs(4670) <= not(layer0_outputs(4247));
    outputs(4671) <= not(layer0_outputs(5453));
    outputs(4672) <= not(layer0_outputs(6015)) or (layer0_outputs(2693));
    outputs(4673) <= layer0_outputs(6443);
    outputs(4674) <= not((layer0_outputs(5447)) and (layer0_outputs(1972)));
    outputs(4675) <= (layer0_outputs(4830)) and (layer0_outputs(2865));
    outputs(4676) <= not(layer0_outputs(4216));
    outputs(4677) <= not(layer0_outputs(6483));
    outputs(4678) <= (layer0_outputs(741)) and not (layer0_outputs(3993));
    outputs(4679) <= (layer0_outputs(3192)) and not (layer0_outputs(4046));
    outputs(4680) <= (layer0_outputs(5777)) and not (layer0_outputs(5732));
    outputs(4681) <= not(layer0_outputs(6912));
    outputs(4682) <= (layer0_outputs(4932)) xor (layer0_outputs(5540));
    outputs(4683) <= not(layer0_outputs(3983));
    outputs(4684) <= not((layer0_outputs(868)) or (layer0_outputs(6207)));
    outputs(4685) <= not(layer0_outputs(1801));
    outputs(4686) <= (layer0_outputs(4000)) xor (layer0_outputs(1067));
    outputs(4687) <= not(layer0_outputs(6895));
    outputs(4688) <= not(layer0_outputs(7668)) or (layer0_outputs(1233));
    outputs(4689) <= layer0_outputs(4019);
    outputs(4690) <= not(layer0_outputs(7476));
    outputs(4691) <= (layer0_outputs(2430)) xor (layer0_outputs(2055));
    outputs(4692) <= not(layer0_outputs(1347));
    outputs(4693) <= not(layer0_outputs(4912));
    outputs(4694) <= (layer0_outputs(6896)) xor (layer0_outputs(7674));
    outputs(4695) <= not(layer0_outputs(1137));
    outputs(4696) <= not((layer0_outputs(3752)) and (layer0_outputs(7025)));
    outputs(4697) <= not(layer0_outputs(3892));
    outputs(4698) <= layer0_outputs(175);
    outputs(4699) <= not(layer0_outputs(6079));
    outputs(4700) <= (layer0_outputs(1616)) xor (layer0_outputs(1141));
    outputs(4701) <= (layer0_outputs(1620)) xor (layer0_outputs(4770));
    outputs(4702) <= (layer0_outputs(6293)) xor (layer0_outputs(2746));
    outputs(4703) <= (layer0_outputs(1843)) xor (layer0_outputs(7102));
    outputs(4704) <= layer0_outputs(6267);
    outputs(4705) <= (layer0_outputs(2155)) and (layer0_outputs(4561));
    outputs(4706) <= (layer0_outputs(12)) and (layer0_outputs(6413));
    outputs(4707) <= not(layer0_outputs(7193));
    outputs(4708) <= not(layer0_outputs(1361));
    outputs(4709) <= layer0_outputs(2718);
    outputs(4710) <= (layer0_outputs(5384)) and (layer0_outputs(7475));
    outputs(4711) <= layer0_outputs(5889);
    outputs(4712) <= (layer0_outputs(2413)) and not (layer0_outputs(2935));
    outputs(4713) <= (layer0_outputs(6849)) xor (layer0_outputs(2015));
    outputs(4714) <= not((layer0_outputs(5717)) or (layer0_outputs(2507)));
    outputs(4715) <= (layer0_outputs(988)) or (layer0_outputs(3060));
    outputs(4716) <= not((layer0_outputs(3422)) and (layer0_outputs(3260)));
    outputs(4717) <= not(layer0_outputs(5288)) or (layer0_outputs(2661));
    outputs(4718) <= not(layer0_outputs(7518));
    outputs(4719) <= not(layer0_outputs(1414));
    outputs(4720) <= not((layer0_outputs(1241)) xor (layer0_outputs(3747)));
    outputs(4721) <= (layer0_outputs(2803)) or (layer0_outputs(4158));
    outputs(4722) <= (layer0_outputs(3843)) or (layer0_outputs(4322));
    outputs(4723) <= layer0_outputs(4133);
    outputs(4724) <= (layer0_outputs(780)) and not (layer0_outputs(6073));
    outputs(4725) <= not(layer0_outputs(3047)) or (layer0_outputs(3604));
    outputs(4726) <= layer0_outputs(2859);
    outputs(4727) <= not(layer0_outputs(2428)) or (layer0_outputs(1472));
    outputs(4728) <= not(layer0_outputs(6958));
    outputs(4729) <= layer0_outputs(4613);
    outputs(4730) <= layer0_outputs(4221);
    outputs(4731) <= (layer0_outputs(1004)) or (layer0_outputs(136));
    outputs(4732) <= (layer0_outputs(847)) and (layer0_outputs(1278));
    outputs(4733) <= (layer0_outputs(1785)) and not (layer0_outputs(2932));
    outputs(4734) <= not((layer0_outputs(3501)) and (layer0_outputs(7651)));
    outputs(4735) <= layer0_outputs(2126);
    outputs(4736) <= layer0_outputs(1409);
    outputs(4737) <= not((layer0_outputs(2903)) xor (layer0_outputs(641)));
    outputs(4738) <= layer0_outputs(6202);
    outputs(4739) <= layer0_outputs(563);
    outputs(4740) <= not(layer0_outputs(3925));
    outputs(4741) <= not((layer0_outputs(6155)) or (layer0_outputs(5236)));
    outputs(4742) <= not(layer0_outputs(7356));
    outputs(4743) <= (layer0_outputs(3231)) and not (layer0_outputs(410));
    outputs(4744) <= (layer0_outputs(3927)) and not (layer0_outputs(4980));
    outputs(4745) <= not((layer0_outputs(435)) and (layer0_outputs(3044)));
    outputs(4746) <= (layer0_outputs(7411)) and not (layer0_outputs(5485));
    outputs(4747) <= not(layer0_outputs(6268)) or (layer0_outputs(2131));
    outputs(4748) <= (layer0_outputs(2011)) or (layer0_outputs(6666));
    outputs(4749) <= not(layer0_outputs(4129));
    outputs(4750) <= (layer0_outputs(6918)) and (layer0_outputs(194));
    outputs(4751) <= (layer0_outputs(4268)) and not (layer0_outputs(5218));
    outputs(4752) <= (layer0_outputs(4996)) and (layer0_outputs(1400));
    outputs(4753) <= layer0_outputs(4629);
    outputs(4754) <= not(layer0_outputs(7367)) or (layer0_outputs(4179));
    outputs(4755) <= not((layer0_outputs(1885)) or (layer0_outputs(140)));
    outputs(4756) <= not((layer0_outputs(7068)) or (layer0_outputs(2759)));
    outputs(4757) <= (layer0_outputs(637)) and not (layer0_outputs(469));
    outputs(4758) <= (layer0_outputs(5785)) and (layer0_outputs(912));
    outputs(4759) <= not(layer0_outputs(7129));
    outputs(4760) <= not(layer0_outputs(2481)) or (layer0_outputs(7587));
    outputs(4761) <= not((layer0_outputs(2144)) xor (layer0_outputs(2571)));
    outputs(4762) <= (layer0_outputs(4843)) and not (layer0_outputs(6965));
    outputs(4763) <= layer0_outputs(2032);
    outputs(4764) <= layer0_outputs(3066);
    outputs(4765) <= not(layer0_outputs(7502));
    outputs(4766) <= not(layer0_outputs(1536));
    outputs(4767) <= not(layer0_outputs(232));
    outputs(4768) <= (layer0_outputs(4882)) and (layer0_outputs(7087));
    outputs(4769) <= (layer0_outputs(5247)) and (layer0_outputs(6980));
    outputs(4770) <= not((layer0_outputs(6097)) and (layer0_outputs(1172)));
    outputs(4771) <= layer0_outputs(181);
    outputs(4772) <= layer0_outputs(1514);
    outputs(4773) <= not(layer0_outputs(2273)) or (layer0_outputs(882));
    outputs(4774) <= not(layer0_outputs(1611));
    outputs(4775) <= layer0_outputs(5565);
    outputs(4776) <= not(layer0_outputs(5931));
    outputs(4777) <= not((layer0_outputs(6383)) xor (layer0_outputs(3577)));
    outputs(4778) <= not((layer0_outputs(3969)) and (layer0_outputs(2225)));
    outputs(4779) <= not(layer0_outputs(5171));
    outputs(4780) <= (layer0_outputs(968)) and (layer0_outputs(5860));
    outputs(4781) <= layer0_outputs(3224);
    outputs(4782) <= (layer0_outputs(5730)) and not (layer0_outputs(6030));
    outputs(4783) <= layer0_outputs(2272);
    outputs(4784) <= not(layer0_outputs(4216));
    outputs(4785) <= layer0_outputs(7312);
    outputs(4786) <= not(layer0_outputs(17));
    outputs(4787) <= not(layer0_outputs(1030));
    outputs(4788) <= layer0_outputs(7625);
    outputs(4789) <= not(layer0_outputs(1001));
    outputs(4790) <= (layer0_outputs(4198)) and not (layer0_outputs(6826));
    outputs(4791) <= not(layer0_outputs(2105)) or (layer0_outputs(6632));
    outputs(4792) <= (layer0_outputs(4196)) and (layer0_outputs(5830));
    outputs(4793) <= not((layer0_outputs(2543)) xor (layer0_outputs(5183)));
    outputs(4794) <= (layer0_outputs(7073)) and not (layer0_outputs(2328));
    outputs(4795) <= not((layer0_outputs(2697)) or (layer0_outputs(4580)));
    outputs(4796) <= not((layer0_outputs(3722)) or (layer0_outputs(6895)));
    outputs(4797) <= not((layer0_outputs(3270)) or (layer0_outputs(2581)));
    outputs(4798) <= (layer0_outputs(2047)) and (layer0_outputs(2140));
    outputs(4799) <= not(layer0_outputs(6108)) or (layer0_outputs(3377));
    outputs(4800) <= layer0_outputs(6062);
    outputs(4801) <= not(layer0_outputs(5568)) or (layer0_outputs(1236));
    outputs(4802) <= not(layer0_outputs(2833)) or (layer0_outputs(2026));
    outputs(4803) <= not(layer0_outputs(7287));
    outputs(4804) <= not(layer0_outputs(4691)) or (layer0_outputs(4594));
    outputs(4805) <= not(layer0_outputs(2528));
    outputs(4806) <= not(layer0_outputs(2137));
    outputs(4807) <= (layer0_outputs(3602)) or (layer0_outputs(1817));
    outputs(4808) <= layer0_outputs(3012);
    outputs(4809) <= not(layer0_outputs(782)) or (layer0_outputs(4690));
    outputs(4810) <= not(layer0_outputs(4637));
    outputs(4811) <= layer0_outputs(4145);
    outputs(4812) <= (layer0_outputs(5300)) and not (layer0_outputs(598));
    outputs(4813) <= layer0_outputs(7392);
    outputs(4814) <= (layer0_outputs(3587)) and not (layer0_outputs(4229));
    outputs(4815) <= not(layer0_outputs(3396)) or (layer0_outputs(187));
    outputs(4816) <= (layer0_outputs(4034)) and not (layer0_outputs(839));
    outputs(4817) <= not((layer0_outputs(4267)) or (layer0_outputs(1274)));
    outputs(4818) <= (layer0_outputs(882)) xor (layer0_outputs(2656));
    outputs(4819) <= not((layer0_outputs(7563)) xor (layer0_outputs(6607)));
    outputs(4820) <= (layer0_outputs(5132)) and not (layer0_outputs(1717));
    outputs(4821) <= not(layer0_outputs(1918));
    outputs(4822) <= not((layer0_outputs(3692)) or (layer0_outputs(304)));
    outputs(4823) <= layer0_outputs(1548);
    outputs(4824) <= layer0_outputs(5006);
    outputs(4825) <= (layer0_outputs(2749)) and not (layer0_outputs(701));
    outputs(4826) <= not(layer0_outputs(5526));
    outputs(4827) <= layer0_outputs(7110);
    outputs(4828) <= (layer0_outputs(4681)) and not (layer0_outputs(3302));
    outputs(4829) <= not(layer0_outputs(4727));
    outputs(4830) <= layer0_outputs(2230);
    outputs(4831) <= layer0_outputs(5008);
    outputs(4832) <= not(layer0_outputs(526));
    outputs(4833) <= layer0_outputs(1220);
    outputs(4834) <= layer0_outputs(250);
    outputs(4835) <= layer0_outputs(6156);
    outputs(4836) <= (layer0_outputs(6482)) and not (layer0_outputs(310));
    outputs(4837) <= layer0_outputs(603);
    outputs(4838) <= layer0_outputs(5442);
    outputs(4839) <= layer0_outputs(960);
    outputs(4840) <= (layer0_outputs(6655)) and (layer0_outputs(6344));
    outputs(4841) <= not(layer0_outputs(2507));
    outputs(4842) <= not(layer0_outputs(6009)) or (layer0_outputs(558));
    outputs(4843) <= not((layer0_outputs(6588)) xor (layer0_outputs(7222)));
    outputs(4844) <= not((layer0_outputs(6249)) or (layer0_outputs(2280)));
    outputs(4845) <= not(layer0_outputs(2013));
    outputs(4846) <= layer0_outputs(6159);
    outputs(4847) <= layer0_outputs(4872);
    outputs(4848) <= layer0_outputs(6622);
    outputs(4849) <= layer0_outputs(219);
    outputs(4850) <= (layer0_outputs(2576)) xor (layer0_outputs(1129));
    outputs(4851) <= not((layer0_outputs(892)) and (layer0_outputs(6711)));
    outputs(4852) <= (layer0_outputs(7370)) and not (layer0_outputs(2148));
    outputs(4853) <= (layer0_outputs(3475)) and not (layer0_outputs(4100));
    outputs(4854) <= not((layer0_outputs(2414)) xor (layer0_outputs(1302)));
    outputs(4855) <= layer0_outputs(5908);
    outputs(4856) <= not(layer0_outputs(5258));
    outputs(4857) <= (layer0_outputs(7174)) and not (layer0_outputs(1717));
    outputs(4858) <= not(layer0_outputs(4669));
    outputs(4859) <= layer0_outputs(5923);
    outputs(4860) <= not(layer0_outputs(3156));
    outputs(4861) <= not(layer0_outputs(3779));
    outputs(4862) <= not(layer0_outputs(5405));
    outputs(4863) <= not(layer0_outputs(4633));
    outputs(4864) <= not((layer0_outputs(3051)) xor (layer0_outputs(5566)));
    outputs(4865) <= layer0_outputs(5974);
    outputs(4866) <= not((layer0_outputs(5129)) or (layer0_outputs(45)));
    outputs(4867) <= layer0_outputs(1192);
    outputs(4868) <= not(layer0_outputs(2595)) or (layer0_outputs(3338));
    outputs(4869) <= layer0_outputs(2120);
    outputs(4870) <= layer0_outputs(6102);
    outputs(4871) <= layer0_outputs(1547);
    outputs(4872) <= (layer0_outputs(3726)) and (layer0_outputs(6756));
    outputs(4873) <= layer0_outputs(5055);
    outputs(4874) <= (layer0_outputs(3237)) xor (layer0_outputs(4069));
    outputs(4875) <= not(layer0_outputs(3770));
    outputs(4876) <= not((layer0_outputs(4607)) xor (layer0_outputs(3889)));
    outputs(4877) <= not((layer0_outputs(5220)) and (layer0_outputs(7044)));
    outputs(4878) <= (layer0_outputs(3431)) and (layer0_outputs(4498));
    outputs(4879) <= not(layer0_outputs(3401));
    outputs(4880) <= (layer0_outputs(5956)) xor (layer0_outputs(2873));
    outputs(4881) <= layer0_outputs(6314);
    outputs(4882) <= (layer0_outputs(809)) and (layer0_outputs(49));
    outputs(4883) <= not(layer0_outputs(4889));
    outputs(4884) <= not(layer0_outputs(3713)) or (layer0_outputs(755));
    outputs(4885) <= not((layer0_outputs(3939)) or (layer0_outputs(6235)));
    outputs(4886) <= layer0_outputs(3628);
    outputs(4887) <= (layer0_outputs(2140)) and not (layer0_outputs(6616));
    outputs(4888) <= (layer0_outputs(3756)) and not (layer0_outputs(6392));
    outputs(4889) <= (layer0_outputs(2403)) or (layer0_outputs(4694));
    outputs(4890) <= not(layer0_outputs(5797)) or (layer0_outputs(5277));
    outputs(4891) <= (layer0_outputs(6689)) or (layer0_outputs(6152));
    outputs(4892) <= not(layer0_outputs(3992));
    outputs(4893) <= layer0_outputs(4358);
    outputs(4894) <= not(layer0_outputs(3022));
    outputs(4895) <= (layer0_outputs(1927)) and not (layer0_outputs(3629));
    outputs(4896) <= (layer0_outputs(4150)) and (layer0_outputs(5224));
    outputs(4897) <= not(layer0_outputs(435));
    outputs(4898) <= not(layer0_outputs(3542));
    outputs(4899) <= not((layer0_outputs(5752)) or (layer0_outputs(4910)));
    outputs(4900) <= layer0_outputs(1018);
    outputs(4901) <= not(layer0_outputs(7285));
    outputs(4902) <= layer0_outputs(5516);
    outputs(4903) <= (layer0_outputs(5473)) and (layer0_outputs(1680));
    outputs(4904) <= not(layer0_outputs(1363));
    outputs(4905) <= not(layer0_outputs(4361));
    outputs(4906) <= (layer0_outputs(6533)) and (layer0_outputs(3511));
    outputs(4907) <= layer0_outputs(5887);
    outputs(4908) <= not(layer0_outputs(2971));
    outputs(4909) <= (layer0_outputs(2531)) and not (layer0_outputs(1406));
    outputs(4910) <= not(layer0_outputs(2723));
    outputs(4911) <= not((layer0_outputs(1300)) xor (layer0_outputs(4785)));
    outputs(4912) <= layer0_outputs(403);
    outputs(4913) <= not((layer0_outputs(4847)) or (layer0_outputs(4132)));
    outputs(4914) <= (layer0_outputs(4961)) and not (layer0_outputs(6429));
    outputs(4915) <= not((layer0_outputs(6519)) and (layer0_outputs(2897)));
    outputs(4916) <= layer0_outputs(2955);
    outputs(4917) <= not(layer0_outputs(1202));
    outputs(4918) <= (layer0_outputs(6670)) and not (layer0_outputs(7448));
    outputs(4919) <= not(layer0_outputs(773));
    outputs(4920) <= layer0_outputs(2728);
    outputs(4921) <= layer0_outputs(4457);
    outputs(4922) <= layer0_outputs(4911);
    outputs(4923) <= not(layer0_outputs(5303));
    outputs(4924) <= not((layer0_outputs(5156)) or (layer0_outputs(3606)));
    outputs(4925) <= layer0_outputs(1286);
    outputs(4926) <= not(layer0_outputs(386)) or (layer0_outputs(4920));
    outputs(4927) <= not(layer0_outputs(7161));
    outputs(4928) <= (layer0_outputs(420)) and not (layer0_outputs(5020));
    outputs(4929) <= not((layer0_outputs(5466)) and (layer0_outputs(6301)));
    outputs(4930) <= (layer0_outputs(6384)) xor (layer0_outputs(2223));
    outputs(4931) <= layer0_outputs(4934);
    outputs(4932) <= (layer0_outputs(5176)) and not (layer0_outputs(5771));
    outputs(4933) <= (layer0_outputs(2699)) xor (layer0_outputs(1960));
    outputs(4934) <= layer0_outputs(6661);
    outputs(4935) <= not(layer0_outputs(6254));
    outputs(4936) <= layer0_outputs(7051);
    outputs(4937) <= (layer0_outputs(2289)) and not (layer0_outputs(7117));
    outputs(4938) <= (layer0_outputs(3447)) xor (layer0_outputs(2709));
    outputs(4939) <= (layer0_outputs(6335)) or (layer0_outputs(6541));
    outputs(4940) <= layer0_outputs(5375);
    outputs(4941) <= not((layer0_outputs(4069)) xor (layer0_outputs(5373)));
    outputs(4942) <= (layer0_outputs(7637)) and (layer0_outputs(223));
    outputs(4943) <= not((layer0_outputs(5637)) or (layer0_outputs(1737)));
    outputs(4944) <= not((layer0_outputs(7371)) or (layer0_outputs(1930)));
    outputs(4945) <= not(layer0_outputs(6805));
    outputs(4946) <= (layer0_outputs(3078)) and not (layer0_outputs(6581));
    outputs(4947) <= (layer0_outputs(2104)) or (layer0_outputs(2567));
    outputs(4948) <= (layer0_outputs(6506)) xor (layer0_outputs(1167));
    outputs(4949) <= layer0_outputs(3249);
    outputs(4950) <= layer0_outputs(838);
    outputs(4951) <= not(layer0_outputs(2051)) or (layer0_outputs(6100));
    outputs(4952) <= not((layer0_outputs(1171)) or (layer0_outputs(5919)));
    outputs(4953) <= (layer0_outputs(213)) xor (layer0_outputs(3637));
    outputs(4954) <= not(layer0_outputs(6616));
    outputs(4955) <= (layer0_outputs(1617)) and not (layer0_outputs(1121));
    outputs(4956) <= layer0_outputs(1288);
    outputs(4957) <= layer0_outputs(2018);
    outputs(4958) <= layer0_outputs(6057);
    outputs(4959) <= (layer0_outputs(7022)) and not (layer0_outputs(4867));
    outputs(4960) <= not((layer0_outputs(6228)) and (layer0_outputs(2812)));
    outputs(4961) <= (layer0_outputs(4285)) xor (layer0_outputs(2754));
    outputs(4962) <= (layer0_outputs(1405)) and not (layer0_outputs(1664));
    outputs(4963) <= not(layer0_outputs(1023));
    outputs(4964) <= not(layer0_outputs(132));
    outputs(4965) <= (layer0_outputs(2021)) and not (layer0_outputs(388));
    outputs(4966) <= layer0_outputs(4027);
    outputs(4967) <= (layer0_outputs(316)) and not (layer0_outputs(2621));
    outputs(4968) <= (layer0_outputs(2107)) or (layer0_outputs(1580));
    outputs(4969) <= layer0_outputs(629);
    outputs(4970) <= not(layer0_outputs(4562)) or (layer0_outputs(4385));
    outputs(4971) <= not((layer0_outputs(3432)) or (layer0_outputs(6465)));
    outputs(4972) <= (layer0_outputs(1396)) and not (layer0_outputs(7376));
    outputs(4973) <= (layer0_outputs(982)) and (layer0_outputs(292));
    outputs(4974) <= (layer0_outputs(1866)) xor (layer0_outputs(3425));
    outputs(4975) <= (layer0_outputs(4996)) or (layer0_outputs(2901));
    outputs(4976) <= not(layer0_outputs(1670));
    outputs(4977) <= layer0_outputs(5358);
    outputs(4978) <= not(layer0_outputs(1569));
    outputs(4979) <= layer0_outputs(557);
    outputs(4980) <= (layer0_outputs(4442)) and not (layer0_outputs(1361));
    outputs(4981) <= not(layer0_outputs(1855));
    outputs(4982) <= (layer0_outputs(6626)) and not (layer0_outputs(46));
    outputs(4983) <= (layer0_outputs(1335)) and (layer0_outputs(1786));
    outputs(4984) <= layer0_outputs(589);
    outputs(4985) <= not(layer0_outputs(6544));
    outputs(4986) <= not(layer0_outputs(5508));
    outputs(4987) <= not(layer0_outputs(6461));
    outputs(4988) <= layer0_outputs(4018);
    outputs(4989) <= not((layer0_outputs(5393)) or (layer0_outputs(4901)));
    outputs(4990) <= not(layer0_outputs(4395));
    outputs(4991) <= layer0_outputs(2587);
    outputs(4992) <= (layer0_outputs(3346)) and not (layer0_outputs(5349));
    outputs(4993) <= (layer0_outputs(5112)) or (layer0_outputs(1026));
    outputs(4994) <= layer0_outputs(3744);
    outputs(4995) <= (layer0_outputs(790)) or (layer0_outputs(354));
    outputs(4996) <= layer0_outputs(639);
    outputs(4997) <= layer0_outputs(3224);
    outputs(4998) <= (layer0_outputs(6830)) or (layer0_outputs(6745));
    outputs(4999) <= (layer0_outputs(6532)) and (layer0_outputs(2250));
    outputs(5000) <= not(layer0_outputs(5338));
    outputs(5001) <= not(layer0_outputs(1878));
    outputs(5002) <= not((layer0_outputs(1947)) or (layer0_outputs(6891)));
    outputs(5003) <= not((layer0_outputs(7037)) xor (layer0_outputs(3298)));
    outputs(5004) <= layer0_outputs(6882);
    outputs(5005) <= (layer0_outputs(5092)) and (layer0_outputs(3789));
    outputs(5006) <= layer0_outputs(6291);
    outputs(5007) <= (layer0_outputs(6379)) and not (layer0_outputs(5833));
    outputs(5008) <= layer0_outputs(5384);
    outputs(5009) <= layer0_outputs(1624);
    outputs(5010) <= layer0_outputs(5309);
    outputs(5011) <= layer0_outputs(1420);
    outputs(5012) <= not(layer0_outputs(3044));
    outputs(5013) <= (layer0_outputs(2793)) and (layer0_outputs(3808));
    outputs(5014) <= (layer0_outputs(4679)) and not (layer0_outputs(5195));
    outputs(5015) <= layer0_outputs(2093);
    outputs(5016) <= (layer0_outputs(4935)) xor (layer0_outputs(2686));
    outputs(5017) <= not(layer0_outputs(3850)) or (layer0_outputs(3191));
    outputs(5018) <= not((layer0_outputs(7515)) or (layer0_outputs(7091)));
    outputs(5019) <= not(layer0_outputs(5454));
    outputs(5020) <= layer0_outputs(5026);
    outputs(5021) <= (layer0_outputs(4091)) and not (layer0_outputs(2911));
    outputs(5022) <= not(layer0_outputs(79));
    outputs(5023) <= not((layer0_outputs(1204)) and (layer0_outputs(6019)));
    outputs(5024) <= (layer0_outputs(6134)) and not (layer0_outputs(3820));
    outputs(5025) <= not(layer0_outputs(4453));
    outputs(5026) <= layer0_outputs(3228);
    outputs(5027) <= layer0_outputs(4959);
    outputs(5028) <= (layer0_outputs(7151)) xor (layer0_outputs(4708));
    outputs(5029) <= layer0_outputs(6286);
    outputs(5030) <= (layer0_outputs(4466)) and not (layer0_outputs(429));
    outputs(5031) <= not((layer0_outputs(5302)) or (layer0_outputs(733)));
    outputs(5032) <= layer0_outputs(1535);
    outputs(5033) <= not(layer0_outputs(3836));
    outputs(5034) <= (layer0_outputs(779)) and not (layer0_outputs(1987));
    outputs(5035) <= not(layer0_outputs(2162));
    outputs(5036) <= (layer0_outputs(3162)) and (layer0_outputs(1677));
    outputs(5037) <= not((layer0_outputs(3614)) xor (layer0_outputs(3393)));
    outputs(5038) <= (layer0_outputs(1543)) xor (layer0_outputs(4762));
    outputs(5039) <= not((layer0_outputs(4353)) xor (layer0_outputs(3189)));
    outputs(5040) <= not((layer0_outputs(3093)) and (layer0_outputs(4139)));
    outputs(5041) <= not(layer0_outputs(54));
    outputs(5042) <= layer0_outputs(6887);
    outputs(5043) <= not(layer0_outputs(6266));
    outputs(5044) <= not(layer0_outputs(4790));
    outputs(5045) <= (layer0_outputs(6463)) or (layer0_outputs(4545));
    outputs(5046) <= layer0_outputs(4240);
    outputs(5047) <= (layer0_outputs(2453)) xor (layer0_outputs(2688));
    outputs(5048) <= not(layer0_outputs(5752));
    outputs(5049) <= (layer0_outputs(1197)) xor (layer0_outputs(4308));
    outputs(5050) <= (layer0_outputs(300)) and (layer0_outputs(3870));
    outputs(5051) <= not((layer0_outputs(766)) xor (layer0_outputs(2556)));
    outputs(5052) <= not((layer0_outputs(2121)) xor (layer0_outputs(1769)));
    outputs(5053) <= (layer0_outputs(3916)) and not (layer0_outputs(4201));
    outputs(5054) <= layer0_outputs(3211);
    outputs(5055) <= layer0_outputs(4561);
    outputs(5056) <= not(layer0_outputs(616)) or (layer0_outputs(5002));
    outputs(5057) <= layer0_outputs(3574);
    outputs(5058) <= not(layer0_outputs(6750));
    outputs(5059) <= (layer0_outputs(1226)) or (layer0_outputs(3116));
    outputs(5060) <= not(layer0_outputs(4861));
    outputs(5061) <= layer0_outputs(4864);
    outputs(5062) <= layer0_outputs(5710);
    outputs(5063) <= layer0_outputs(7051);
    outputs(5064) <= not(layer0_outputs(4567));
    outputs(5065) <= layer0_outputs(5196);
    outputs(5066) <= layer0_outputs(7000);
    outputs(5067) <= layer0_outputs(2270);
    outputs(5068) <= not(layer0_outputs(7361)) or (layer0_outputs(5274));
    outputs(5069) <= (layer0_outputs(7293)) and (layer0_outputs(2472));
    outputs(5070) <= layer0_outputs(6765);
    outputs(5071) <= (layer0_outputs(6420)) and not (layer0_outputs(5999));
    outputs(5072) <= (layer0_outputs(1628)) or (layer0_outputs(7620));
    outputs(5073) <= layer0_outputs(7252);
    outputs(5074) <= not(layer0_outputs(2585)) or (layer0_outputs(841));
    outputs(5075) <= not(layer0_outputs(323)) or (layer0_outputs(7167));
    outputs(5076) <= not(layer0_outputs(383));
    outputs(5077) <= (layer0_outputs(1170)) or (layer0_outputs(2173));
    outputs(5078) <= not((layer0_outputs(3285)) xor (layer0_outputs(5660)));
    outputs(5079) <= (layer0_outputs(3706)) and not (layer0_outputs(3263));
    outputs(5080) <= not((layer0_outputs(216)) and (layer0_outputs(3830)));
    outputs(5081) <= (layer0_outputs(3080)) and not (layer0_outputs(3152));
    outputs(5082) <= (layer0_outputs(4698)) xor (layer0_outputs(7655));
    outputs(5083) <= (layer0_outputs(3173)) xor (layer0_outputs(1771));
    outputs(5084) <= not(layer0_outputs(2748));
    outputs(5085) <= not(layer0_outputs(7582));
    outputs(5086) <= layer0_outputs(2900);
    outputs(5087) <= not((layer0_outputs(5981)) or (layer0_outputs(2683)));
    outputs(5088) <= layer0_outputs(7004);
    outputs(5089) <= layer0_outputs(537);
    outputs(5090) <= (layer0_outputs(3568)) or (layer0_outputs(1436));
    outputs(5091) <= not(layer0_outputs(2101));
    outputs(5092) <= layer0_outputs(607);
    outputs(5093) <= not((layer0_outputs(6079)) and (layer0_outputs(4655)));
    outputs(5094) <= not(layer0_outputs(179));
    outputs(5095) <= not(layer0_outputs(5052));
    outputs(5096) <= (layer0_outputs(870)) and (layer0_outputs(5643));
    outputs(5097) <= layer0_outputs(3031);
    outputs(5098) <= not(layer0_outputs(652));
    outputs(5099) <= not((layer0_outputs(2893)) or (layer0_outputs(1682)));
    outputs(5100) <= not(layer0_outputs(1703));
    outputs(5101) <= (layer0_outputs(1135)) and (layer0_outputs(7603));
    outputs(5102) <= (layer0_outputs(7262)) and not (layer0_outputs(2282));
    outputs(5103) <= not((layer0_outputs(2635)) or (layer0_outputs(2887)));
    outputs(5104) <= layer0_outputs(1563);
    outputs(5105) <= (layer0_outputs(2506)) and not (layer0_outputs(4431));
    outputs(5106) <= layer0_outputs(3110);
    outputs(5107) <= layer0_outputs(4232);
    outputs(5108) <= layer0_outputs(2317);
    outputs(5109) <= layer0_outputs(4166);
    outputs(5110) <= (layer0_outputs(1501)) and not (layer0_outputs(6001));
    outputs(5111) <= layer0_outputs(6332);
    outputs(5112) <= (layer0_outputs(813)) and (layer0_outputs(1696));
    outputs(5113) <= not((layer0_outputs(1610)) or (layer0_outputs(2632)));
    outputs(5114) <= not(layer0_outputs(6993)) or (layer0_outputs(5944));
    outputs(5115) <= not(layer0_outputs(3123)) or (layer0_outputs(3794));
    outputs(5116) <= layer0_outputs(6057);
    outputs(5117) <= (layer0_outputs(6586)) and not (layer0_outputs(232));
    outputs(5118) <= (layer0_outputs(2399)) and not (layer0_outputs(1622));
    outputs(5119) <= layer0_outputs(4777);
    outputs(5120) <= layer0_outputs(450);
    outputs(5121) <= layer0_outputs(7067);
    outputs(5122) <= (layer0_outputs(4444)) and not (layer0_outputs(7217));
    outputs(5123) <= (layer0_outputs(6402)) and (layer0_outputs(3493));
    outputs(5124) <= (layer0_outputs(5396)) and (layer0_outputs(2653));
    outputs(5125) <= not(layer0_outputs(1165));
    outputs(5126) <= layer0_outputs(1541);
    outputs(5127) <= not(layer0_outputs(6034)) or (layer0_outputs(5727));
    outputs(5128) <= not(layer0_outputs(1692)) or (layer0_outputs(234));
    outputs(5129) <= not(layer0_outputs(1626));
    outputs(5130) <= layer0_outputs(284);
    outputs(5131) <= (layer0_outputs(6787)) and (layer0_outputs(1131));
    outputs(5132) <= not(layer0_outputs(4647));
    outputs(5133) <= layer0_outputs(4598);
    outputs(5134) <= not((layer0_outputs(7478)) xor (layer0_outputs(2208)));
    outputs(5135) <= layer0_outputs(7279);
    outputs(5136) <= (layer0_outputs(7077)) and not (layer0_outputs(4310));
    outputs(5137) <= (layer0_outputs(4165)) and not (layer0_outputs(1227));
    outputs(5138) <= (layer0_outputs(3954)) and not (layer0_outputs(6780));
    outputs(5139) <= (layer0_outputs(4484)) and (layer0_outputs(126));
    outputs(5140) <= not((layer0_outputs(894)) xor (layer0_outputs(3547)));
    outputs(5141) <= (layer0_outputs(5184)) and not (layer0_outputs(5476));
    outputs(5142) <= (layer0_outputs(3293)) and not (layer0_outputs(3325));
    outputs(5143) <= (layer0_outputs(7183)) and (layer0_outputs(5744));
    outputs(5144) <= not((layer0_outputs(1039)) or (layer0_outputs(1061)));
    outputs(5145) <= not(layer0_outputs(3847)) or (layer0_outputs(7575));
    outputs(5146) <= layer0_outputs(2420);
    outputs(5147) <= not(layer0_outputs(1311));
    outputs(5148) <= layer0_outputs(7112);
    outputs(5149) <= not(layer0_outputs(4889));
    outputs(5150) <= not(layer0_outputs(5322));
    outputs(5151) <= layer0_outputs(6470);
    outputs(5152) <= not(layer0_outputs(2974)) or (layer0_outputs(6767));
    outputs(5153) <= (layer0_outputs(5814)) and (layer0_outputs(731));
    outputs(5154) <= layer0_outputs(7093);
    outputs(5155) <= (layer0_outputs(5234)) and not (layer0_outputs(7670));
    outputs(5156) <= not(layer0_outputs(4264));
    outputs(5157) <= (layer0_outputs(4714)) or (layer0_outputs(88));
    outputs(5158) <= not(layer0_outputs(5060)) or (layer0_outputs(5716));
    outputs(5159) <= not(layer0_outputs(4871));
    outputs(5160) <= not(layer0_outputs(4945));
    outputs(5161) <= layer0_outputs(2844);
    outputs(5162) <= not((layer0_outputs(4276)) xor (layer0_outputs(5281)));
    outputs(5163) <= (layer0_outputs(2983)) xor (layer0_outputs(4073));
    outputs(5164) <= layer0_outputs(3364);
    outputs(5165) <= not(layer0_outputs(3579));
    outputs(5166) <= (layer0_outputs(3050)) and (layer0_outputs(5574));
    outputs(5167) <= (layer0_outputs(266)) xor (layer0_outputs(5900));
    outputs(5168) <= not(layer0_outputs(372)) or (layer0_outputs(5503));
    outputs(5169) <= layer0_outputs(3936);
    outputs(5170) <= not(layer0_outputs(924));
    outputs(5171) <= not((layer0_outputs(3000)) or (layer0_outputs(2703)));
    outputs(5172) <= not(layer0_outputs(6329));
    outputs(5173) <= not((layer0_outputs(7256)) xor (layer0_outputs(7337)));
    outputs(5174) <= not(layer0_outputs(810));
    outputs(5175) <= (layer0_outputs(2334)) xor (layer0_outputs(639));
    outputs(5176) <= (layer0_outputs(220)) and (layer0_outputs(3691));
    outputs(5177) <= not(layer0_outputs(5360));
    outputs(5178) <= (layer0_outputs(3101)) and (layer0_outputs(5022));
    outputs(5179) <= (layer0_outputs(2330)) and not (layer0_outputs(1884));
    outputs(5180) <= layer0_outputs(543);
    outputs(5181) <= layer0_outputs(5180);
    outputs(5182) <= (layer0_outputs(1337)) and (layer0_outputs(5871));
    outputs(5183) <= not(layer0_outputs(6516)) or (layer0_outputs(2205));
    outputs(5184) <= not(layer0_outputs(550));
    outputs(5185) <= not(layer0_outputs(3178));
    outputs(5186) <= not(layer0_outputs(264));
    outputs(5187) <= layer0_outputs(792);
    outputs(5188) <= not((layer0_outputs(2827)) or (layer0_outputs(1203)));
    outputs(5189) <= layer0_outputs(4374);
    outputs(5190) <= layer0_outputs(2064);
    outputs(5191) <= not((layer0_outputs(4775)) xor (layer0_outputs(5737)));
    outputs(5192) <= not(layer0_outputs(1529));
    outputs(5193) <= not(layer0_outputs(3520));
    outputs(5194) <= not((layer0_outputs(2683)) or (layer0_outputs(3356)));
    outputs(5195) <= not(layer0_outputs(1619));
    outputs(5196) <= not((layer0_outputs(4631)) or (layer0_outputs(289)));
    outputs(5197) <= (layer0_outputs(6693)) xor (layer0_outputs(3792));
    outputs(5198) <= not((layer0_outputs(7542)) and (layer0_outputs(3894)));
    outputs(5199) <= not(layer0_outputs(7144)) or (layer0_outputs(1167));
    outputs(5200) <= not(layer0_outputs(4207));
    outputs(5201) <= not((layer0_outputs(2417)) or (layer0_outputs(190)));
    outputs(5202) <= not(layer0_outputs(2462)) or (layer0_outputs(2317));
    outputs(5203) <= layer0_outputs(1525);
    outputs(5204) <= not(layer0_outputs(1711));
    outputs(5205) <= not(layer0_outputs(7647));
    outputs(5206) <= layer0_outputs(1526);
    outputs(5207) <= (layer0_outputs(3109)) and (layer0_outputs(2435));
    outputs(5208) <= not(layer0_outputs(2059));
    outputs(5209) <= (layer0_outputs(1303)) and (layer0_outputs(3333));
    outputs(5210) <= (layer0_outputs(7174)) and (layer0_outputs(7516));
    outputs(5211) <= layer0_outputs(6673);
    outputs(5212) <= not(layer0_outputs(1720));
    outputs(5213) <= layer0_outputs(6364);
    outputs(5214) <= (layer0_outputs(3011)) and (layer0_outputs(377));
    outputs(5215) <= (layer0_outputs(7136)) xor (layer0_outputs(6307));
    outputs(5216) <= (layer0_outputs(6790)) and not (layer0_outputs(5550));
    outputs(5217) <= (layer0_outputs(2778)) and not (layer0_outputs(4447));
    outputs(5218) <= (layer0_outputs(6718)) and not (layer0_outputs(4191));
    outputs(5219) <= layer0_outputs(5221);
    outputs(5220) <= (layer0_outputs(5714)) xor (layer0_outputs(6842));
    outputs(5221) <= not(layer0_outputs(6694));
    outputs(5222) <= not(layer0_outputs(6));
    outputs(5223) <= (layer0_outputs(6012)) xor (layer0_outputs(2142));
    outputs(5224) <= layer0_outputs(6617);
    outputs(5225) <= layer0_outputs(7324);
    outputs(5226) <= not(layer0_outputs(5178));
    outputs(5227) <= (layer0_outputs(5107)) xor (layer0_outputs(738));
    outputs(5228) <= not(layer0_outputs(1966));
    outputs(5229) <= layer0_outputs(4187);
    outputs(5230) <= not(layer0_outputs(2395));
    outputs(5231) <= not(layer0_outputs(6559));
    outputs(5232) <= (layer0_outputs(3185)) xor (layer0_outputs(6633));
    outputs(5233) <= (layer0_outputs(3897)) or (layer0_outputs(2609));
    outputs(5234) <= layer0_outputs(2915);
    outputs(5235) <= not(layer0_outputs(6043));
    outputs(5236) <= (layer0_outputs(3117)) and (layer0_outputs(4928));
    outputs(5237) <= layer0_outputs(5018);
    outputs(5238) <= not((layer0_outputs(4247)) or (layer0_outputs(1357)));
    outputs(5239) <= not(layer0_outputs(3560));
    outputs(5240) <= (layer0_outputs(2056)) and not (layer0_outputs(6539));
    outputs(5241) <= not((layer0_outputs(4606)) xor (layer0_outputs(3209)));
    outputs(5242) <= layer0_outputs(2718);
    outputs(5243) <= not(layer0_outputs(1101));
    outputs(5244) <= (layer0_outputs(1477)) and not (layer0_outputs(7460));
    outputs(5245) <= not(layer0_outputs(4015));
    outputs(5246) <= (layer0_outputs(4914)) and (layer0_outputs(279));
    outputs(5247) <= not(layer0_outputs(4469));
    outputs(5248) <= not((layer0_outputs(595)) and (layer0_outputs(5214)));
    outputs(5249) <= (layer0_outputs(3235)) and not (layer0_outputs(3437));
    outputs(5250) <= layer0_outputs(1453);
    outputs(5251) <= layer0_outputs(4);
    outputs(5252) <= not(layer0_outputs(3832));
    outputs(5253) <= not((layer0_outputs(3718)) and (layer0_outputs(5511)));
    outputs(5254) <= layer0_outputs(1005);
    outputs(5255) <= not(layer0_outputs(59));
    outputs(5256) <= (layer0_outputs(4989)) and (layer0_outputs(2577));
    outputs(5257) <= not(layer0_outputs(6554));
    outputs(5258) <= not(layer0_outputs(2959));
    outputs(5259) <= (layer0_outputs(4135)) and (layer0_outputs(6910));
    outputs(5260) <= not(layer0_outputs(2672)) or (layer0_outputs(7297));
    outputs(5261) <= not(layer0_outputs(3491));
    outputs(5262) <= not((layer0_outputs(6822)) xor (layer0_outputs(4964)));
    outputs(5263) <= (layer0_outputs(3470)) and not (layer0_outputs(8));
    outputs(5264) <= not((layer0_outputs(3986)) xor (layer0_outputs(6401)));
    outputs(5265) <= layer0_outputs(2874);
    outputs(5266) <= not(layer0_outputs(4702));
    outputs(5267) <= (layer0_outputs(7649)) or (layer0_outputs(3566));
    outputs(5268) <= (layer0_outputs(1380)) and not (layer0_outputs(3064));
    outputs(5269) <= not((layer0_outputs(6467)) xor (layer0_outputs(1406)));
    outputs(5270) <= not((layer0_outputs(7470)) or (layer0_outputs(5854)));
    outputs(5271) <= (layer0_outputs(2790)) and (layer0_outputs(5391));
    outputs(5272) <= not(layer0_outputs(6549));
    outputs(5273) <= (layer0_outputs(4127)) and not (layer0_outputs(1566));
    outputs(5274) <= (layer0_outputs(3183)) and not (layer0_outputs(4471));
    outputs(5275) <= not(layer0_outputs(545));
    outputs(5276) <= not(layer0_outputs(7547));
    outputs(5277) <= layer0_outputs(6974);
    outputs(5278) <= (layer0_outputs(3466)) and (layer0_outputs(621));
    outputs(5279) <= (layer0_outputs(7398)) and not (layer0_outputs(3173));
    outputs(5280) <= layer0_outputs(1436);
    outputs(5281) <= layer0_outputs(4984);
    outputs(5282) <= layer0_outputs(2236);
    outputs(5283) <= (layer0_outputs(2087)) and not (layer0_outputs(5383));
    outputs(5284) <= not((layer0_outputs(3488)) and (layer0_outputs(6777)));
    outputs(5285) <= not(layer0_outputs(4427)) or (layer0_outputs(4200));
    outputs(5286) <= not(layer0_outputs(4723));
    outputs(5287) <= (layer0_outputs(6313)) and not (layer0_outputs(6839));
    outputs(5288) <= not(layer0_outputs(904));
    outputs(5289) <= not(layer0_outputs(2747)) or (layer0_outputs(5818));
    outputs(5290) <= not(layer0_outputs(4300)) or (layer0_outputs(2955));
    outputs(5291) <= (layer0_outputs(7294)) and not (layer0_outputs(6975));
    outputs(5292) <= not(layer0_outputs(385)) or (layer0_outputs(7319));
    outputs(5293) <= layer0_outputs(6413);
    outputs(5294) <= not(layer0_outputs(4386));
    outputs(5295) <= layer0_outputs(271);
    outputs(5296) <= layer0_outputs(3509);
    outputs(5297) <= (layer0_outputs(2130)) xor (layer0_outputs(1040));
    outputs(5298) <= layer0_outputs(5491);
    outputs(5299) <= (layer0_outputs(157)) and not (layer0_outputs(474));
    outputs(5300) <= not((layer0_outputs(4847)) and (layer0_outputs(7455)));
    outputs(5301) <= (layer0_outputs(5715)) and not (layer0_outputs(2063));
    outputs(5302) <= not((layer0_outputs(874)) xor (layer0_outputs(438)));
    outputs(5303) <= not(layer0_outputs(5352));
    outputs(5304) <= (layer0_outputs(64)) and not (layer0_outputs(504));
    outputs(5305) <= not((layer0_outputs(3397)) or (layer0_outputs(101)));
    outputs(5306) <= not(layer0_outputs(5746));
    outputs(5307) <= not(layer0_outputs(5155)) or (layer0_outputs(6916));
    outputs(5308) <= not(layer0_outputs(1939));
    outputs(5309) <= layer0_outputs(3203);
    outputs(5310) <= not((layer0_outputs(6211)) xor (layer0_outputs(5510)));
    outputs(5311) <= not(layer0_outputs(5005));
    outputs(5312) <= layer0_outputs(3382);
    outputs(5313) <= not(layer0_outputs(753));
    outputs(5314) <= (layer0_outputs(5167)) and not (layer0_outputs(2541));
    outputs(5315) <= not(layer0_outputs(7164));
    outputs(5316) <= not(layer0_outputs(1446));
    outputs(5317) <= not((layer0_outputs(2033)) or (layer0_outputs(2288)));
    outputs(5318) <= not(layer0_outputs(6497));
    outputs(5319) <= not(layer0_outputs(1157));
    outputs(5320) <= not(layer0_outputs(4222));
    outputs(5321) <= not((layer0_outputs(1015)) xor (layer0_outputs(7026)));
    outputs(5322) <= layer0_outputs(1134);
    outputs(5323) <= (layer0_outputs(7475)) and (layer0_outputs(1541));
    outputs(5324) <= not(layer0_outputs(6860));
    outputs(5325) <= not(layer0_outputs(5349)) or (layer0_outputs(4919));
    outputs(5326) <= not((layer0_outputs(7224)) xor (layer0_outputs(2821)));
    outputs(5327) <= layer0_outputs(3728);
    outputs(5328) <= (layer0_outputs(1690)) and (layer0_outputs(7276));
    outputs(5329) <= layer0_outputs(860);
    outputs(5330) <= (layer0_outputs(242)) and (layer0_outputs(5196));
    outputs(5331) <= not((layer0_outputs(6163)) and (layer0_outputs(97)));
    outputs(5332) <= layer0_outputs(3882);
    outputs(5333) <= not(layer0_outputs(742));
    outputs(5334) <= (layer0_outputs(4179)) and not (layer0_outputs(1668));
    outputs(5335) <= not(layer0_outputs(2710));
    outputs(5336) <= layer0_outputs(6508);
    outputs(5337) <= (layer0_outputs(2563)) and (layer0_outputs(1417));
    outputs(5338) <= not(layer0_outputs(1171)) or (layer0_outputs(5457));
    outputs(5339) <= not(layer0_outputs(2858)) or (layer0_outputs(6691));
    outputs(5340) <= layer0_outputs(5640);
    outputs(5341) <= layer0_outputs(4110);
    outputs(5342) <= layer0_outputs(6179);
    outputs(5343) <= not((layer0_outputs(6638)) or (layer0_outputs(1737)));
    outputs(5344) <= not(layer0_outputs(29));
    outputs(5345) <= not((layer0_outputs(2344)) or (layer0_outputs(2641)));
    outputs(5346) <= not(layer0_outputs(832));
    outputs(5347) <= (layer0_outputs(5004)) and (layer0_outputs(6846));
    outputs(5348) <= not((layer0_outputs(3263)) or (layer0_outputs(1594)));
    outputs(5349) <= not(layer0_outputs(7311));
    outputs(5350) <= not((layer0_outputs(6467)) xor (layer0_outputs(1391)));
    outputs(5351) <= not((layer0_outputs(6693)) or (layer0_outputs(4966)));
    outputs(5352) <= layer0_outputs(215);
    outputs(5353) <= not(layer0_outputs(128)) or (layer0_outputs(792));
    outputs(5354) <= not((layer0_outputs(1348)) or (layer0_outputs(5847)));
    outputs(5355) <= (layer0_outputs(7630)) and not (layer0_outputs(1345));
    outputs(5356) <= (layer0_outputs(6648)) and not (layer0_outputs(3250));
    outputs(5357) <= (layer0_outputs(1374)) and not (layer0_outputs(5202));
    outputs(5358) <= (layer0_outputs(1427)) and not (layer0_outputs(807));
    outputs(5359) <= not(layer0_outputs(3869)) or (layer0_outputs(2985));
    outputs(5360) <= (layer0_outputs(5012)) and not (layer0_outputs(5209));
    outputs(5361) <= not(layer0_outputs(7665));
    outputs(5362) <= layer0_outputs(7231);
    outputs(5363) <= layer0_outputs(5639);
    outputs(5364) <= layer0_outputs(1083);
    outputs(5365) <= not(layer0_outputs(6561));
    outputs(5366) <= layer0_outputs(5503);
    outputs(5367) <= (layer0_outputs(4956)) and (layer0_outputs(1022));
    outputs(5368) <= layer0_outputs(5923);
    outputs(5369) <= not((layer0_outputs(1888)) or (layer0_outputs(4266)));
    outputs(5370) <= layer0_outputs(2205);
    outputs(5371) <= not(layer0_outputs(387));
    outputs(5372) <= (layer0_outputs(3866)) xor (layer0_outputs(6481));
    outputs(5373) <= not(layer0_outputs(6235)) or (layer0_outputs(3879));
    outputs(5374) <= not(layer0_outputs(1363));
    outputs(5375) <= (layer0_outputs(6087)) and not (layer0_outputs(5131));
    outputs(5376) <= not(layer0_outputs(5478));
    outputs(5377) <= not(layer0_outputs(2693)) or (layer0_outputs(4154));
    outputs(5378) <= not(layer0_outputs(5199));
    outputs(5379) <= layer0_outputs(3778);
    outputs(5380) <= not((layer0_outputs(452)) xor (layer0_outputs(3516)));
    outputs(5381) <= layer0_outputs(5056);
    outputs(5382) <= not(layer0_outputs(3125));
    outputs(5383) <= not(layer0_outputs(4104));
    outputs(5384) <= not((layer0_outputs(7363)) or (layer0_outputs(5186)));
    outputs(5385) <= not(layer0_outputs(2575));
    outputs(5386) <= layer0_outputs(6292);
    outputs(5387) <= layer0_outputs(7670);
    outputs(5388) <= (layer0_outputs(6098)) and not (layer0_outputs(7459));
    outputs(5389) <= layer0_outputs(4407);
    outputs(5390) <= not(layer0_outputs(7511));
    outputs(5391) <= (layer0_outputs(1401)) and not (layer0_outputs(6239));
    outputs(5392) <= layer0_outputs(424);
    outputs(5393) <= not(layer0_outputs(6227));
    outputs(5394) <= not((layer0_outputs(3690)) xor (layer0_outputs(2640)));
    outputs(5395) <= (layer0_outputs(2519)) and (layer0_outputs(2616));
    outputs(5396) <= (layer0_outputs(5263)) or (layer0_outputs(35));
    outputs(5397) <= not((layer0_outputs(3662)) or (layer0_outputs(2877)));
    outputs(5398) <= (layer0_outputs(4468)) or (layer0_outputs(2071));
    outputs(5399) <= layer0_outputs(3345);
    outputs(5400) <= not(layer0_outputs(2756));
    outputs(5401) <= not(layer0_outputs(5271));
    outputs(5402) <= (layer0_outputs(5431)) xor (layer0_outputs(4092));
    outputs(5403) <= not(layer0_outputs(5595));
    outputs(5404) <= not(layer0_outputs(7088));
    outputs(5405) <= (layer0_outputs(1152)) and not (layer0_outputs(3404));
    outputs(5406) <= not((layer0_outputs(6897)) or (layer0_outputs(2494)));
    outputs(5407) <= not((layer0_outputs(322)) xor (layer0_outputs(5722)));
    outputs(5408) <= not(layer0_outputs(4539)) or (layer0_outputs(5736));
    outputs(5409) <= not((layer0_outputs(775)) xor (layer0_outputs(3442)));
    outputs(5410) <= (layer0_outputs(5995)) xor (layer0_outputs(4064));
    outputs(5411) <= not(layer0_outputs(5846)) or (layer0_outputs(487));
    outputs(5412) <= (layer0_outputs(7140)) xor (layer0_outputs(42));
    outputs(5413) <= not(layer0_outputs(4298));
    outputs(5414) <= layer0_outputs(7234);
    outputs(5415) <= (layer0_outputs(6072)) and (layer0_outputs(3097));
    outputs(5416) <= not(layer0_outputs(1244));
    outputs(5417) <= not((layer0_outputs(5562)) or (layer0_outputs(4891)));
    outputs(5418) <= (layer0_outputs(1640)) and not (layer0_outputs(5257));
    outputs(5419) <= not(layer0_outputs(7408));
    outputs(5420) <= (layer0_outputs(6176)) and not (layer0_outputs(6027));
    outputs(5421) <= (layer0_outputs(7417)) and not (layer0_outputs(6603));
    outputs(5422) <= layer0_outputs(2031);
    outputs(5423) <= (layer0_outputs(7275)) or (layer0_outputs(6067));
    outputs(5424) <= (layer0_outputs(5401)) and not (layer0_outputs(6493));
    outputs(5425) <= (layer0_outputs(3113)) and not (layer0_outputs(1948));
    outputs(5426) <= not(layer0_outputs(730));
    outputs(5427) <= (layer0_outputs(2319)) and not (layer0_outputs(5921));
    outputs(5428) <= (layer0_outputs(5935)) and not (layer0_outputs(4318));
    outputs(5429) <= not(layer0_outputs(1530));
    outputs(5430) <= not(layer0_outputs(7346)) or (layer0_outputs(6793));
    outputs(5431) <= not(layer0_outputs(7514)) or (layer0_outputs(536));
    outputs(5432) <= layer0_outputs(5021);
    outputs(5433) <= layer0_outputs(6136);
    outputs(5434) <= not(layer0_outputs(11));
    outputs(5435) <= layer0_outputs(1597);
    outputs(5436) <= layer0_outputs(3748);
    outputs(5437) <= not(layer0_outputs(6178));
    outputs(5438) <= not((layer0_outputs(7096)) or (layer0_outputs(7523)));
    outputs(5439) <= (layer0_outputs(394)) and not (layer0_outputs(1292));
    outputs(5440) <= not((layer0_outputs(5504)) or (layer0_outputs(1022)));
    outputs(5441) <= not((layer0_outputs(705)) xor (layer0_outputs(7013)));
    outputs(5442) <= not((layer0_outputs(2346)) xor (layer0_outputs(782)));
    outputs(5443) <= (layer0_outputs(2808)) and (layer0_outputs(3607));
    outputs(5444) <= (layer0_outputs(1706)) and not (layer0_outputs(3504));
    outputs(5445) <= not(layer0_outputs(2691));
    outputs(5446) <= not((layer0_outputs(4625)) or (layer0_outputs(2984)));
    outputs(5447) <= layer0_outputs(7089);
    outputs(5448) <= layer0_outputs(6946);
    outputs(5449) <= layer0_outputs(654);
    outputs(5450) <= (layer0_outputs(2112)) and not (layer0_outputs(4420));
    outputs(5451) <= not(layer0_outputs(3845));
    outputs(5452) <= layer0_outputs(6251);
    outputs(5453) <= layer0_outputs(6351);
    outputs(5454) <= (layer0_outputs(1101)) and (layer0_outputs(1219));
    outputs(5455) <= (layer0_outputs(188)) and (layer0_outputs(4641));
    outputs(5456) <= not(layer0_outputs(3015));
    outputs(5457) <= (layer0_outputs(6181)) xor (layer0_outputs(5927));
    outputs(5458) <= layer0_outputs(2997);
    outputs(5459) <= not(layer0_outputs(1912));
    outputs(5460) <= layer0_outputs(3373);
    outputs(5461) <= not(layer0_outputs(5085));
    outputs(5462) <= not(layer0_outputs(6206));
    outputs(5463) <= not(layer0_outputs(5100));
    outputs(5464) <= (layer0_outputs(1584)) and not (layer0_outputs(4428));
    outputs(5465) <= not(layer0_outputs(2978));
    outputs(5466) <= not((layer0_outputs(7358)) or (layer0_outputs(1200)));
    outputs(5467) <= (layer0_outputs(595)) and not (layer0_outputs(2369));
    outputs(5468) <= (layer0_outputs(2465)) and not (layer0_outputs(1775));
    outputs(5469) <= not(layer0_outputs(254)) or (layer0_outputs(734));
    outputs(5470) <= (layer0_outputs(7375)) and not (layer0_outputs(75));
    outputs(5471) <= (layer0_outputs(3583)) and not (layer0_outputs(4115));
    outputs(5472) <= (layer0_outputs(2375)) and not (layer0_outputs(2830));
    outputs(5473) <= not((layer0_outputs(4748)) or (layer0_outputs(2007)));
    outputs(5474) <= not(layer0_outputs(7192)) or (layer0_outputs(5973));
    outputs(5475) <= not(layer0_outputs(6217));
    outputs(5476) <= layer0_outputs(4025);
    outputs(5477) <= (layer0_outputs(4360)) and not (layer0_outputs(3916));
    outputs(5478) <= not(layer0_outputs(3364));
    outputs(5479) <= (layer0_outputs(7602)) and not (layer0_outputs(6148));
    outputs(5480) <= not(layer0_outputs(5907));
    outputs(5481) <= not((layer0_outputs(6213)) and (layer0_outputs(4999)));
    outputs(5482) <= (layer0_outputs(3426)) and (layer0_outputs(6330));
    outputs(5483) <= not(layer0_outputs(913));
    outputs(5484) <= not(layer0_outputs(4818)) or (layer0_outputs(7486));
    outputs(5485) <= not(layer0_outputs(2664));
    outputs(5486) <= not(layer0_outputs(4008));
    outputs(5487) <= layer0_outputs(2119);
    outputs(5488) <= (layer0_outputs(5260)) and not (layer0_outputs(5251));
    outputs(5489) <= (layer0_outputs(2218)) or (layer0_outputs(4411));
    outputs(5490) <= (layer0_outputs(6627)) xor (layer0_outputs(1528));
    outputs(5491) <= layer0_outputs(2310);
    outputs(5492) <= layer0_outputs(4796);
    outputs(5493) <= not((layer0_outputs(6094)) or (layer0_outputs(1115)));
    outputs(5494) <= (layer0_outputs(7152)) and not (layer0_outputs(3167));
    outputs(5495) <= not(layer0_outputs(6317));
    outputs(5496) <= (layer0_outputs(3539)) and (layer0_outputs(1344));
    outputs(5497) <= (layer0_outputs(6546)) xor (layer0_outputs(5735));
    outputs(5498) <= layer0_outputs(1698);
    outputs(5499) <= not((layer0_outputs(451)) or (layer0_outputs(4887)));
    outputs(5500) <= layer0_outputs(2716);
    outputs(5501) <= (layer0_outputs(7180)) and not (layer0_outputs(6219));
    outputs(5502) <= not((layer0_outputs(4164)) xor (layer0_outputs(1806)));
    outputs(5503) <= not(layer0_outputs(6434));
    outputs(5504) <= layer0_outputs(5692);
    outputs(5505) <= not(layer0_outputs(6206)) or (layer0_outputs(3693));
    outputs(5506) <= (layer0_outputs(6028)) or (layer0_outputs(6934));
    outputs(5507) <= not((layer0_outputs(5988)) or (layer0_outputs(525)));
    outputs(5508) <= (layer0_outputs(374)) xor (layer0_outputs(3154));
    outputs(5509) <= not(layer0_outputs(4259)) or (layer0_outputs(5248));
    outputs(5510) <= (layer0_outputs(4260)) and (layer0_outputs(183));
    outputs(5511) <= layer0_outputs(4495);
    outputs(5512) <= not(layer0_outputs(3095));
    outputs(5513) <= not(layer0_outputs(3638));
    outputs(5514) <= not((layer0_outputs(5902)) or (layer0_outputs(2492)));
    outputs(5515) <= (layer0_outputs(5307)) and not (layer0_outputs(948));
    outputs(5516) <= not(layer0_outputs(2407));
    outputs(5517) <= not(layer0_outputs(6978));
    outputs(5518) <= layer0_outputs(6362);
    outputs(5519) <= (layer0_outputs(5334)) and not (layer0_outputs(5957));
    outputs(5520) <= layer0_outputs(3652);
    outputs(5521) <= not(layer0_outputs(1184));
    outputs(5522) <= not(layer0_outputs(5850));
    outputs(5523) <= layer0_outputs(7512);
    outputs(5524) <= not(layer0_outputs(7607));
    outputs(5525) <= (layer0_outputs(4884)) and not (layer0_outputs(1751));
    outputs(5526) <= (layer0_outputs(4688)) and not (layer0_outputs(6041));
    outputs(5527) <= (layer0_outputs(3542)) and not (layer0_outputs(2526));
    outputs(5528) <= layer0_outputs(6182);
    outputs(5529) <= (layer0_outputs(2801)) and (layer0_outputs(2290));
    outputs(5530) <= layer0_outputs(2299);
    outputs(5531) <= layer0_outputs(2846);
    outputs(5532) <= not((layer0_outputs(825)) or (layer0_outputs(411)));
    outputs(5533) <= (layer0_outputs(7049)) and not (layer0_outputs(7271));
    outputs(5534) <= layer0_outputs(3576);
    outputs(5535) <= (layer0_outputs(6221)) and (layer0_outputs(3395));
    outputs(5536) <= not(layer0_outputs(7244));
    outputs(5537) <= layer0_outputs(2046);
    outputs(5538) <= (layer0_outputs(4240)) xor (layer0_outputs(6315));
    outputs(5539) <= not(layer0_outputs(7060));
    outputs(5540) <= (layer0_outputs(2221)) and not (layer0_outputs(5688));
    outputs(5541) <= layer0_outputs(3247);
    outputs(5542) <= layer0_outputs(7562);
    outputs(5543) <= not((layer0_outputs(1691)) and (layer0_outputs(392)));
    outputs(5544) <= not(layer0_outputs(6081));
    outputs(5545) <= not((layer0_outputs(109)) xor (layer0_outputs(313)));
    outputs(5546) <= (layer0_outputs(3153)) or (layer0_outputs(4327));
    outputs(5547) <= (layer0_outputs(5730)) and not (layer0_outputs(7010));
    outputs(5548) <= not(layer0_outputs(194));
    outputs(5549) <= (layer0_outputs(5950)) and not (layer0_outputs(2432));
    outputs(5550) <= not((layer0_outputs(3827)) or (layer0_outputs(425)));
    outputs(5551) <= layer0_outputs(4689);
    outputs(5552) <= (layer0_outputs(4790)) and not (layer0_outputs(5122));
    outputs(5553) <= not((layer0_outputs(5114)) xor (layer0_outputs(5350)));
    outputs(5554) <= (layer0_outputs(3809)) and not (layer0_outputs(3697));
    outputs(5555) <= not(layer0_outputs(7639));
    outputs(5556) <= not((layer0_outputs(1642)) or (layer0_outputs(5672)));
    outputs(5557) <= not(layer0_outputs(6338));
    outputs(5558) <= (layer0_outputs(2445)) or (layer0_outputs(362));
    outputs(5559) <= not(layer0_outputs(6050));
    outputs(5560) <= not(layer0_outputs(7613));
    outputs(5561) <= (layer0_outputs(2310)) and not (layer0_outputs(4646));
    outputs(5562) <= (layer0_outputs(2929)) and not (layer0_outputs(2956));
    outputs(5563) <= (layer0_outputs(1123)) and not (layer0_outputs(1965));
    outputs(5564) <= not((layer0_outputs(4652)) or (layer0_outputs(517)));
    outputs(5565) <= not((layer0_outputs(95)) or (layer0_outputs(7549)));
    outputs(5566) <= (layer0_outputs(6829)) and not (layer0_outputs(6763));
    outputs(5567) <= (layer0_outputs(5931)) and not (layer0_outputs(5924));
    outputs(5568) <= layer0_outputs(3322);
    outputs(5569) <= not(layer0_outputs(4450)) or (layer0_outputs(5812));
    outputs(5570) <= (layer0_outputs(3736)) and (layer0_outputs(5024));
    outputs(5571) <= (layer0_outputs(272)) and (layer0_outputs(3006));
    outputs(5572) <= not((layer0_outputs(6739)) or (layer0_outputs(4054)));
    outputs(5573) <= not(layer0_outputs(2852));
    outputs(5574) <= layer0_outputs(1438);
    outputs(5575) <= not((layer0_outputs(2811)) or (layer0_outputs(7074)));
    outputs(5576) <= layer0_outputs(2314);
    outputs(5577) <= layer0_outputs(573);
    outputs(5578) <= not(layer0_outputs(6179));
    outputs(5579) <= (layer0_outputs(1130)) and not (layer0_outputs(3141));
    outputs(5580) <= (layer0_outputs(7512)) and (layer0_outputs(6814));
    outputs(5581) <= (layer0_outputs(419)) and (layer0_outputs(832));
    outputs(5582) <= not(layer0_outputs(7653)) or (layer0_outputs(3561));
    outputs(5583) <= (layer0_outputs(5754)) and (layer0_outputs(7119));
    outputs(5584) <= not(layer0_outputs(4075));
    outputs(5585) <= not(layer0_outputs(5408));
    outputs(5586) <= (layer0_outputs(4519)) xor (layer0_outputs(7043));
    outputs(5587) <= not(layer0_outputs(7466));
    outputs(5588) <= layer0_outputs(3107);
    outputs(5589) <= (layer0_outputs(5288)) and not (layer0_outputs(7221));
    outputs(5590) <= layer0_outputs(5856);
    outputs(5591) <= (layer0_outputs(1687)) and not (layer0_outputs(1499));
    outputs(5592) <= not(layer0_outputs(2058));
    outputs(5593) <= (layer0_outputs(3785)) and not (layer0_outputs(2630));
    outputs(5594) <= not((layer0_outputs(7285)) xor (layer0_outputs(5698)));
    outputs(5595) <= (layer0_outputs(7021)) and (layer0_outputs(1425));
    outputs(5596) <= not(layer0_outputs(5233)) or (layer0_outputs(5723));
    outputs(5597) <= (layer0_outputs(5013)) and (layer0_outputs(3863));
    outputs(5598) <= layer0_outputs(297);
    outputs(5599) <= not((layer0_outputs(3643)) xor (layer0_outputs(6590)));
    outputs(5600) <= not((layer0_outputs(4534)) and (layer0_outputs(170)));
    outputs(5601) <= not((layer0_outputs(5659)) or (layer0_outputs(191)));
    outputs(5602) <= layer0_outputs(1901);
    outputs(5603) <= not(layer0_outputs(6134));
    outputs(5604) <= layer0_outputs(2883);
    outputs(5605) <= not(layer0_outputs(486));
    outputs(5606) <= (layer0_outputs(6589)) and not (layer0_outputs(7175));
    outputs(5607) <= (layer0_outputs(5900)) and not (layer0_outputs(5409));
    outputs(5608) <= (layer0_outputs(2528)) and (layer0_outputs(7135));
    outputs(5609) <= layer0_outputs(7120);
    outputs(5610) <= not(layer0_outputs(3050));
    outputs(5611) <= layer0_outputs(4933);
    outputs(5612) <= not(layer0_outputs(6213));
    outputs(5613) <= not((layer0_outputs(7093)) or (layer0_outputs(6493)));
    outputs(5614) <= not((layer0_outputs(160)) or (layer0_outputs(5065)));
    outputs(5615) <= (layer0_outputs(2182)) and not (layer0_outputs(87));
    outputs(5616) <= layer0_outputs(4647);
    outputs(5617) <= layer0_outputs(4280);
    outputs(5618) <= layer0_outputs(7269);
    outputs(5619) <= layer0_outputs(2345);
    outputs(5620) <= not((layer0_outputs(3857)) xor (layer0_outputs(3379)));
    outputs(5621) <= layer0_outputs(7179);
    outputs(5622) <= not((layer0_outputs(1264)) and (layer0_outputs(7104)));
    outputs(5623) <= not((layer0_outputs(3191)) and (layer0_outputs(263)));
    outputs(5624) <= not((layer0_outputs(2037)) or (layer0_outputs(6364)));
    outputs(5625) <= not(layer0_outputs(2950));
    outputs(5626) <= (layer0_outputs(4283)) and not (layer0_outputs(6481));
    outputs(5627) <= (layer0_outputs(3443)) and (layer0_outputs(5612));
    outputs(5628) <= not((layer0_outputs(6089)) and (layer0_outputs(2177)));
    outputs(5629) <= not((layer0_outputs(389)) xor (layer0_outputs(1815)));
    outputs(5630) <= not((layer0_outputs(5753)) xor (layer0_outputs(4414)));
    outputs(5631) <= (layer0_outputs(6547)) xor (layer0_outputs(4890));
    outputs(5632) <= (layer0_outputs(1940)) and not (layer0_outputs(7520));
    outputs(5633) <= (layer0_outputs(4330)) and not (layer0_outputs(5917));
    outputs(5634) <= not(layer0_outputs(6943));
    outputs(5635) <= (layer0_outputs(716)) xor (layer0_outputs(2271));
    outputs(5636) <= layer0_outputs(3841);
    outputs(5637) <= layer0_outputs(430);
    outputs(5638) <= (layer0_outputs(2987)) and not (layer0_outputs(697));
    outputs(5639) <= not((layer0_outputs(5767)) or (layer0_outputs(5647)));
    outputs(5640) <= layer0_outputs(5602);
    outputs(5641) <= layer0_outputs(4339);
    outputs(5642) <= not((layer0_outputs(6899)) xor (layer0_outputs(6570)));
    outputs(5643) <= (layer0_outputs(172)) and (layer0_outputs(1992));
    outputs(5644) <= (layer0_outputs(2159)) and not (layer0_outputs(7071));
    outputs(5645) <= (layer0_outputs(5559)) or (layer0_outputs(669));
    outputs(5646) <= (layer0_outputs(1671)) and not (layer0_outputs(1872));
    outputs(5647) <= (layer0_outputs(3751)) and not (layer0_outputs(2369));
    outputs(5648) <= not((layer0_outputs(4627)) xor (layer0_outputs(4961)));
    outputs(5649) <= not(layer0_outputs(1629));
    outputs(5650) <= layer0_outputs(1720);
    outputs(5651) <= layer0_outputs(5405);
    outputs(5652) <= layer0_outputs(5156);
    outputs(5653) <= not(layer0_outputs(4351));
    outputs(5654) <= not(layer0_outputs(1195));
    outputs(5655) <= layer0_outputs(2586);
    outputs(5656) <= layer0_outputs(3329);
    outputs(5657) <= not(layer0_outputs(6320));
    outputs(5658) <= not(layer0_outputs(4133));
    outputs(5659) <= not(layer0_outputs(4245)) or (layer0_outputs(4651));
    outputs(5660) <= not(layer0_outputs(7437));
    outputs(5661) <= (layer0_outputs(1312)) and (layer0_outputs(4243));
    outputs(5662) <= layer0_outputs(360);
    outputs(5663) <= (layer0_outputs(2786)) and not (layer0_outputs(4077));
    outputs(5664) <= not((layer0_outputs(2453)) xor (layer0_outputs(5264)));
    outputs(5665) <= not((layer0_outputs(5032)) and (layer0_outputs(5194)));
    outputs(5666) <= layer0_outputs(1822);
    outputs(5667) <= (layer0_outputs(7294)) xor (layer0_outputs(7516));
    outputs(5668) <= not((layer0_outputs(520)) or (layer0_outputs(2329)));
    outputs(5669) <= not((layer0_outputs(6698)) xor (layer0_outputs(4141)));
    outputs(5670) <= (layer0_outputs(833)) and not (layer0_outputs(2441));
    outputs(5671) <= (layer0_outputs(5498)) and not (layer0_outputs(3733));
    outputs(5672) <= layer0_outputs(4446);
    outputs(5673) <= not((layer0_outputs(2276)) xor (layer0_outputs(4477)));
    outputs(5674) <= layer0_outputs(5541);
    outputs(5675) <= not(layer0_outputs(5436));
    outputs(5676) <= (layer0_outputs(1049)) and (layer0_outputs(2445));
    outputs(5677) <= (layer0_outputs(5365)) and not (layer0_outputs(6970));
    outputs(5678) <= layer0_outputs(1732);
    outputs(5679) <= (layer0_outputs(672)) xor (layer0_outputs(6214));
    outputs(5680) <= not(layer0_outputs(547));
    outputs(5681) <= not(layer0_outputs(2175));
    outputs(5682) <= (layer0_outputs(5862)) and not (layer0_outputs(2458));
    outputs(5683) <= not((layer0_outputs(3285)) or (layer0_outputs(336)));
    outputs(5684) <= not((layer0_outputs(213)) xor (layer0_outputs(251)));
    outputs(5685) <= not((layer0_outputs(546)) xor (layer0_outputs(2428)));
    outputs(5686) <= (layer0_outputs(489)) and not (layer0_outputs(3473));
    outputs(5687) <= not(layer0_outputs(62));
    outputs(5688) <= (layer0_outputs(3636)) and not (layer0_outputs(1439));
    outputs(5689) <= (layer0_outputs(5821)) and not (layer0_outputs(1089));
    outputs(5690) <= not((layer0_outputs(1197)) or (layer0_outputs(3712)));
    outputs(5691) <= not(layer0_outputs(4202));
    outputs(5692) <= not((layer0_outputs(7481)) xor (layer0_outputs(4319)));
    outputs(5693) <= layer0_outputs(966);
    outputs(5694) <= not(layer0_outputs(3464));
    outputs(5695) <= not((layer0_outputs(2930)) and (layer0_outputs(6928)));
    outputs(5696) <= (layer0_outputs(7350)) and not (layer0_outputs(1818));
    outputs(5697) <= layer0_outputs(7460);
    outputs(5698) <= layer0_outputs(6512);
    outputs(5699) <= not(layer0_outputs(7672));
    outputs(5700) <= layer0_outputs(3251);
    outputs(5701) <= not(layer0_outputs(497));
    outputs(5702) <= (layer0_outputs(1996)) and not (layer0_outputs(7006));
    outputs(5703) <= layer0_outputs(5144);
    outputs(5704) <= not(layer0_outputs(5219)) or (layer0_outputs(5133));
    outputs(5705) <= not(layer0_outputs(2155));
    outputs(5706) <= layer0_outputs(4658);
    outputs(5707) <= not((layer0_outputs(5217)) xor (layer0_outputs(483)));
    outputs(5708) <= layer0_outputs(4231);
    outputs(5709) <= layer0_outputs(6962);
    outputs(5710) <= not(layer0_outputs(4513)) or (layer0_outputs(6517));
    outputs(5711) <= not((layer0_outputs(6357)) xor (layer0_outputs(2845)));
    outputs(5712) <= (layer0_outputs(3894)) and not (layer0_outputs(2485));
    outputs(5713) <= not(layer0_outputs(2664));
    outputs(5714) <= (layer0_outputs(4877)) and (layer0_outputs(2416));
    outputs(5715) <= not((layer0_outputs(4443)) xor (layer0_outputs(6083)));
    outputs(5716) <= not(layer0_outputs(3908));
    outputs(5717) <= not((layer0_outputs(5165)) or (layer0_outputs(2484)));
    outputs(5718) <= (layer0_outputs(2808)) and not (layer0_outputs(947));
    outputs(5719) <= not(layer0_outputs(1331));
    outputs(5720) <= layer0_outputs(1191);
    outputs(5721) <= not(layer0_outputs(6536));
    outputs(5722) <= not((layer0_outputs(3215)) xor (layer0_outputs(1250)));
    outputs(5723) <= (layer0_outputs(2893)) and not (layer0_outputs(5389));
    outputs(5724) <= not((layer0_outputs(2820)) xor (layer0_outputs(468)));
    outputs(5725) <= (layer0_outputs(50)) and (layer0_outputs(7142));
    outputs(5726) <= (layer0_outputs(7387)) or (layer0_outputs(6654));
    outputs(5727) <= (layer0_outputs(6492)) and (layer0_outputs(4931));
    outputs(5728) <= (layer0_outputs(726)) and not (layer0_outputs(4404));
    outputs(5729) <= not(layer0_outputs(1708));
    outputs(5730) <= (layer0_outputs(2427)) and not (layer0_outputs(4392));
    outputs(5731) <= not(layer0_outputs(2010)) or (layer0_outputs(2364));
    outputs(5732) <= not(layer0_outputs(1323));
    outputs(5733) <= layer0_outputs(4177);
    outputs(5734) <= not((layer0_outputs(7063)) or (layer0_outputs(5852)));
    outputs(5735) <= (layer0_outputs(1505)) and not (layer0_outputs(286));
    outputs(5736) <= (layer0_outputs(6194)) and not (layer0_outputs(2276));
    outputs(5737) <= not(layer0_outputs(5443));
    outputs(5738) <= (layer0_outputs(4614)) and (layer0_outputs(78));
    outputs(5739) <= layer0_outputs(1119);
    outputs(5740) <= not((layer0_outputs(5881)) or (layer0_outputs(6403)));
    outputs(5741) <= (layer0_outputs(6398)) or (layer0_outputs(1521));
    outputs(5742) <= not(layer0_outputs(3534));
    outputs(5743) <= not(layer0_outputs(6064)) or (layer0_outputs(1113));
    outputs(5744) <= layer0_outputs(4509);
    outputs(5745) <= (layer0_outputs(1516)) xor (layer0_outputs(3948));
    outputs(5746) <= (layer0_outputs(6868)) and (layer0_outputs(4059));
    outputs(5747) <= not((layer0_outputs(2509)) or (layer0_outputs(268)));
    outputs(5748) <= layer0_outputs(2766);
    outputs(5749) <= layer0_outputs(3380);
    outputs(5750) <= not((layer0_outputs(3100)) xor (layer0_outputs(3138)));
    outputs(5751) <= not(layer0_outputs(528)) or (layer0_outputs(4536));
    outputs(5752) <= not(layer0_outputs(6677));
    outputs(5753) <= (layer0_outputs(5014)) xor (layer0_outputs(5187));
    outputs(5754) <= layer0_outputs(7184);
    outputs(5755) <= (layer0_outputs(6430)) and not (layer0_outputs(754));
    outputs(5756) <= (layer0_outputs(4480)) and not (layer0_outputs(544));
    outputs(5757) <= (layer0_outputs(428)) xor (layer0_outputs(3221));
    outputs(5758) <= not(layer0_outputs(2323)) or (layer0_outputs(7251));
    outputs(5759) <= not((layer0_outputs(5487)) xor (layer0_outputs(3014)));
    outputs(5760) <= layer0_outputs(6860);
    outputs(5761) <= (layer0_outputs(4117)) and not (layer0_outputs(4611));
    outputs(5762) <= (layer0_outputs(1989)) and not (layer0_outputs(4578));
    outputs(5763) <= not((layer0_outputs(6618)) or (layer0_outputs(540)));
    outputs(5764) <= not(layer0_outputs(6763));
    outputs(5765) <= not(layer0_outputs(3092));
    outputs(5766) <= (layer0_outputs(4667)) and not (layer0_outputs(3691));
    outputs(5767) <= (layer0_outputs(5333)) and (layer0_outputs(3075));
    outputs(5768) <= (layer0_outputs(4048)) and not (layer0_outputs(6742));
    outputs(5769) <= not(layer0_outputs(4683));
    outputs(5770) <= not(layer0_outputs(2320));
    outputs(5771) <= not((layer0_outputs(5801)) or (layer0_outputs(1781)));
    outputs(5772) <= layer0_outputs(1077);
    outputs(5773) <= (layer0_outputs(4242)) and not (layer0_outputs(3702));
    outputs(5774) <= not(layer0_outputs(6884));
    outputs(5775) <= not(layer0_outputs(1796));
    outputs(5776) <= (layer0_outputs(2293)) xor (layer0_outputs(7340));
    outputs(5777) <= (layer0_outputs(940)) and not (layer0_outputs(2485));
    outputs(5778) <= not((layer0_outputs(3565)) xor (layer0_outputs(2619)));
    outputs(5779) <= not(layer0_outputs(7467));
    outputs(5780) <= not(layer0_outputs(6045));
    outputs(5781) <= (layer0_outputs(6410)) and not (layer0_outputs(7669));
    outputs(5782) <= not(layer0_outputs(4497)) or (layer0_outputs(6024));
    outputs(5783) <= not((layer0_outputs(585)) or (layer0_outputs(5949)));
    outputs(5784) <= (layer0_outputs(5699)) xor (layer0_outputs(1958));
    outputs(5785) <= not(layer0_outputs(1067));
    outputs(5786) <= (layer0_outputs(4908)) and (layer0_outputs(5853));
    outputs(5787) <= (layer0_outputs(6529)) and not (layer0_outputs(5952));
    outputs(5788) <= (layer0_outputs(6155)) and not (layer0_outputs(3757));
    outputs(5789) <= (layer0_outputs(5749)) and (layer0_outputs(3755));
    outputs(5790) <= layer0_outputs(259);
    outputs(5791) <= (layer0_outputs(1219)) and not (layer0_outputs(5292));
    outputs(5792) <= (layer0_outputs(3921)) and (layer0_outputs(3274));
    outputs(5793) <= layer0_outputs(7522);
    outputs(5794) <= layer0_outputs(3873);
    outputs(5795) <= (layer0_outputs(2229)) and not (layer0_outputs(5774));
    outputs(5796) <= layer0_outputs(1888);
    outputs(5797) <= not((layer0_outputs(3744)) or (layer0_outputs(404)));
    outputs(5798) <= not((layer0_outputs(2368)) and (layer0_outputs(5998)));
    outputs(5799) <= (layer0_outputs(4723)) and (layer0_outputs(1452));
    outputs(5800) <= (layer0_outputs(7578)) and (layer0_outputs(197));
    outputs(5801) <= not((layer0_outputs(2894)) or (layer0_outputs(5482)));
    outputs(5802) <= (layer0_outputs(4753)) and (layer0_outputs(1142));
    outputs(5803) <= layer0_outputs(6561);
    outputs(5804) <= (layer0_outputs(3978)) and not (layer0_outputs(2761));
    outputs(5805) <= layer0_outputs(5903);
    outputs(5806) <= layer0_outputs(1339);
    outputs(5807) <= (layer0_outputs(4637)) and (layer0_outputs(4130));
    outputs(5808) <= (layer0_outputs(2665)) and (layer0_outputs(3745));
    outputs(5809) <= not((layer0_outputs(6015)) xor (layer0_outputs(6251)));
    outputs(5810) <= not((layer0_outputs(6237)) or (layer0_outputs(5346)));
    outputs(5811) <= (layer0_outputs(1614)) and not (layer0_outputs(5896));
    outputs(5812) <= (layer0_outputs(3303)) and (layer0_outputs(1539));
    outputs(5813) <= (layer0_outputs(5461)) and not (layer0_outputs(6060));
    outputs(5814) <= (layer0_outputs(6069)) and (layer0_outputs(7632));
    outputs(5815) <= not((layer0_outputs(1280)) or (layer0_outputs(2264)));
    outputs(5816) <= (layer0_outputs(914)) and (layer0_outputs(5416));
    outputs(5817) <= layer0_outputs(6121);
    outputs(5818) <= (layer0_outputs(4330)) and not (layer0_outputs(4692));
    outputs(5819) <= layer0_outputs(176);
    outputs(5820) <= (layer0_outputs(3900)) and not (layer0_outputs(2194));
    outputs(5821) <= not(layer0_outputs(2209));
    outputs(5822) <= not((layer0_outputs(2869)) or (layer0_outputs(235)));
    outputs(5823) <= not(layer0_outputs(3082));
    outputs(5824) <= (layer0_outputs(5235)) and not (layer0_outputs(348));
    outputs(5825) <= (layer0_outputs(4520)) and not (layer0_outputs(2431));
    outputs(5826) <= not((layer0_outputs(1753)) xor (layer0_outputs(4913)));
    outputs(5827) <= not(layer0_outputs(6798));
    outputs(5828) <= (layer0_outputs(305)) or (layer0_outputs(4447));
    outputs(5829) <= layer0_outputs(6232);
    outputs(5830) <= not(layer0_outputs(5987));
    outputs(5831) <= not(layer0_outputs(5704)) or (layer0_outputs(1944));
    outputs(5832) <= (layer0_outputs(6709)) and not (layer0_outputs(6094));
    outputs(5833) <= layer0_outputs(2966);
    outputs(5834) <= (layer0_outputs(233)) xor (layer0_outputs(3704));
    outputs(5835) <= not((layer0_outputs(750)) xor (layer0_outputs(1269)));
    outputs(5836) <= (layer0_outputs(7310)) and (layer0_outputs(3121));
    outputs(5837) <= not(layer0_outputs(2335));
    outputs(5838) <= (layer0_outputs(3113)) or (layer0_outputs(974));
    outputs(5839) <= (layer0_outputs(7218)) xor (layer0_outputs(7648));
    outputs(5840) <= layer0_outputs(5000);
    outputs(5841) <= not(layer0_outputs(775));
    outputs(5842) <= not(layer0_outputs(6122)) or (layer0_outputs(4029));
    outputs(5843) <= (layer0_outputs(2665)) and (layer0_outputs(1887));
    outputs(5844) <= (layer0_outputs(3101)) or (layer0_outputs(7127));
    outputs(5845) <= layer0_outputs(106);
    outputs(5846) <= not(layer0_outputs(5463));
    outputs(5847) <= not((layer0_outputs(218)) or (layer0_outputs(3128)));
    outputs(5848) <= (layer0_outputs(2747)) and (layer0_outputs(3014));
    outputs(5849) <= layer0_outputs(5691);
    outputs(5850) <= not(layer0_outputs(2739));
    outputs(5851) <= (layer0_outputs(1425)) and (layer0_outputs(3588));
    outputs(5852) <= layer0_outputs(938);
    outputs(5853) <= (layer0_outputs(6793)) and not (layer0_outputs(4700));
    outputs(5854) <= not(layer0_outputs(7289));
    outputs(5855) <= not((layer0_outputs(5261)) or (layer0_outputs(5442)));
    outputs(5856) <= layer0_outputs(4937);
    outputs(5857) <= layer0_outputs(1489);
    outputs(5858) <= (layer0_outputs(1800)) xor (layer0_outputs(58));
    outputs(5859) <= not(layer0_outputs(6156));
    outputs(5860) <= not((layer0_outputs(5)) xor (layer0_outputs(6800)));
    outputs(5861) <= not(layer0_outputs(5844));
    outputs(5862) <= (layer0_outputs(2713)) and not (layer0_outputs(6987));
    outputs(5863) <= not((layer0_outputs(2644)) or (layer0_outputs(3890)));
    outputs(5864) <= not((layer0_outputs(5311)) or (layer0_outputs(7177)));
    outputs(5865) <= (layer0_outputs(6307)) and (layer0_outputs(150));
    outputs(5866) <= not((layer0_outputs(4603)) xor (layer0_outputs(2259)));
    outputs(5867) <= not(layer0_outputs(3243));
    outputs(5868) <= not(layer0_outputs(3931));
    outputs(5869) <= not(layer0_outputs(6252));
    outputs(5870) <= layer0_outputs(1431);
    outputs(5871) <= not(layer0_outputs(3408));
    outputs(5872) <= not((layer0_outputs(5514)) and (layer0_outputs(3893)));
    outputs(5873) <= not(layer0_outputs(5595));
    outputs(5874) <= not(layer0_outputs(6614));
    outputs(5875) <= not((layer0_outputs(1019)) or (layer0_outputs(627)));
    outputs(5876) <= not(layer0_outputs(7308));
    outputs(5877) <= not(layer0_outputs(6137)) or (layer0_outputs(5653));
    outputs(5878) <= not((layer0_outputs(4510)) and (layer0_outputs(7316)));
    outputs(5879) <= not(layer0_outputs(7155));
    outputs(5880) <= (layer0_outputs(7659)) and (layer0_outputs(633));
    outputs(5881) <= not((layer0_outputs(3589)) or (layer0_outputs(3505)));
    outputs(5882) <= layer0_outputs(4908);
    outputs(5883) <= not((layer0_outputs(6955)) or (layer0_outputs(1085)));
    outputs(5884) <= not(layer0_outputs(580)) or (layer0_outputs(6424));
    outputs(5885) <= not(layer0_outputs(70));
    outputs(5886) <= (layer0_outputs(5019)) or (layer0_outputs(2020));
    outputs(5887) <= not((layer0_outputs(565)) or (layer0_outputs(2074)));
    outputs(5888) <= not((layer0_outputs(6022)) or (layer0_outputs(4295)));
    outputs(5889) <= (layer0_outputs(506)) or (layer0_outputs(2505));
    outputs(5890) <= not((layer0_outputs(7048)) xor (layer0_outputs(4558)));
    outputs(5891) <= not(layer0_outputs(20)) or (layer0_outputs(2523));
    outputs(5892) <= not(layer0_outputs(5680)) or (layer0_outputs(2697));
    outputs(5893) <= (layer0_outputs(6848)) xor (layer0_outputs(4731));
    outputs(5894) <= not(layer0_outputs(3313));
    outputs(5895) <= (layer0_outputs(717)) xor (layer0_outputs(3705));
    outputs(5896) <= (layer0_outputs(1127)) and not (layer0_outputs(2075));
    outputs(5897) <= layer0_outputs(2980);
    outputs(5898) <= layer0_outputs(3081);
    outputs(5899) <= not((layer0_outputs(5443)) and (layer0_outputs(7472)));
    outputs(5900) <= (layer0_outputs(3006)) and (layer0_outputs(3019));
    outputs(5901) <= (layer0_outputs(3739)) and not (layer0_outputs(2098));
    outputs(5902) <= (layer0_outputs(4949)) and (layer0_outputs(958));
    outputs(5903) <= (layer0_outputs(6698)) and (layer0_outputs(6014));
    outputs(5904) <= not((layer0_outputs(416)) xor (layer0_outputs(7206)));
    outputs(5905) <= not((layer0_outputs(6892)) or (layer0_outputs(1012)));
    outputs(5906) <= (layer0_outputs(4468)) and not (layer0_outputs(5857));
    outputs(5907) <= not((layer0_outputs(6798)) and (layer0_outputs(1599)));
    outputs(5908) <= (layer0_outputs(5024)) and not (layer0_outputs(1723));
    outputs(5909) <= not(layer0_outputs(2138));
    outputs(5910) <= layer0_outputs(6864);
    outputs(5911) <= (layer0_outputs(7193)) and not (layer0_outputs(6025));
    outputs(5912) <= (layer0_outputs(3920)) xor (layer0_outputs(3321));
    outputs(5913) <= layer0_outputs(3413);
    outputs(5914) <= (layer0_outputs(1626)) and not (layer0_outputs(2946));
    outputs(5915) <= layer0_outputs(5486);
    outputs(5916) <= not((layer0_outputs(2950)) xor (layer0_outputs(700)));
    outputs(5917) <= (layer0_outputs(164)) and not (layer0_outputs(2266));
    outputs(5918) <= (layer0_outputs(5819)) and not (layer0_outputs(2567));
    outputs(5919) <= not(layer0_outputs(640)) or (layer0_outputs(3867));
    outputs(5920) <= not((layer0_outputs(2995)) xor (layer0_outputs(540)));
    outputs(5921) <= not(layer0_outputs(5715)) or (layer0_outputs(4469));
    outputs(5922) <= not(layer0_outputs(66));
    outputs(5923) <= (layer0_outputs(6656)) or (layer0_outputs(2699));
    outputs(5924) <= not(layer0_outputs(3987)) or (layer0_outputs(7439));
    outputs(5925) <= not((layer0_outputs(3157)) or (layer0_outputs(1236)));
    outputs(5926) <= (layer0_outputs(1172)) and (layer0_outputs(612));
    outputs(5927) <= layer0_outputs(709);
    outputs(5928) <= layer0_outputs(906);
    outputs(5929) <= not(layer0_outputs(1889));
    outputs(5930) <= (layer0_outputs(4925)) and not (layer0_outputs(2196));
    outputs(5931) <= not(layer0_outputs(7268));
    outputs(5932) <= not((layer0_outputs(2335)) or (layer0_outputs(1006)));
    outputs(5933) <= layer0_outputs(7161);
    outputs(5934) <= (layer0_outputs(3821)) or (layer0_outputs(2723));
    outputs(5935) <= layer0_outputs(4793);
    outputs(5936) <= (layer0_outputs(787)) or (layer0_outputs(843));
    outputs(5937) <= (layer0_outputs(2040)) and not (layer0_outputs(5376));
    outputs(5938) <= (layer0_outputs(2022)) and not (layer0_outputs(5121));
    outputs(5939) <= not(layer0_outputs(1777)) or (layer0_outputs(6971));
    outputs(5940) <= not((layer0_outputs(5600)) or (layer0_outputs(4533)));
    outputs(5941) <= (layer0_outputs(1297)) and not (layer0_outputs(7573));
    outputs(5942) <= not(layer0_outputs(3698));
    outputs(5943) <= (layer0_outputs(2077)) and not (layer0_outputs(3676));
    outputs(5944) <= (layer0_outputs(1911)) and (layer0_outputs(4244));
    outputs(5945) <= (layer0_outputs(1470)) and (layer0_outputs(7212));
    outputs(5946) <= not((layer0_outputs(5341)) xor (layer0_outputs(2600)));
    outputs(5947) <= not((layer0_outputs(2733)) xor (layer0_outputs(6558)));
    outputs(5948) <= not(layer0_outputs(7260));
    outputs(5949) <= (layer0_outputs(4939)) or (layer0_outputs(6562));
    outputs(5950) <= not(layer0_outputs(2780));
    outputs(5951) <= layer0_outputs(5915);
    outputs(5952) <= not(layer0_outputs(4714));
    outputs(5953) <= not(layer0_outputs(7032));
    outputs(5954) <= not(layer0_outputs(16));
    outputs(5955) <= (layer0_outputs(3351)) or (layer0_outputs(3942));
    outputs(5956) <= layer0_outputs(2799);
    outputs(5957) <= (layer0_outputs(256)) and (layer0_outputs(4068));
    outputs(5958) <= (layer0_outputs(1154)) and not (layer0_outputs(6811));
    outputs(5959) <= (layer0_outputs(3780)) and (layer0_outputs(1900));
    outputs(5960) <= not(layer0_outputs(7316)) or (layer0_outputs(5505));
    outputs(5961) <= not(layer0_outputs(5259)) or (layer0_outputs(2443));
    outputs(5962) <= not(layer0_outputs(5556));
    outputs(5963) <= (layer0_outputs(6537)) and not (layer0_outputs(6276));
    outputs(5964) <= (layer0_outputs(6189)) and (layer0_outputs(4207));
    outputs(5965) <= (layer0_outputs(3753)) and not (layer0_outputs(3890));
    outputs(5966) <= (layer0_outputs(7131)) xor (layer0_outputs(1465));
    outputs(5967) <= layer0_outputs(4105);
    outputs(5968) <= layer0_outputs(4276);
    outputs(5969) <= not(layer0_outputs(3204));
    outputs(5970) <= not((layer0_outputs(6162)) or (layer0_outputs(4112)));
    outputs(5971) <= (layer0_outputs(6117)) and not (layer0_outputs(5186));
    outputs(5972) <= not((layer0_outputs(3403)) xor (layer0_outputs(5451)));
    outputs(5973) <= not(layer0_outputs(7363));
    outputs(5974) <= (layer0_outputs(1204)) and not (layer0_outputs(5029));
    outputs(5975) <= (layer0_outputs(229)) xor (layer0_outputs(4084));
    outputs(5976) <= not((layer0_outputs(5594)) and (layer0_outputs(3331)));
    outputs(5977) <= not((layer0_outputs(6310)) or (layer0_outputs(6578)));
    outputs(5978) <= not(layer0_outputs(1963));
    outputs(5979) <= not((layer0_outputs(5128)) xor (layer0_outputs(6699)));
    outputs(5980) <= (layer0_outputs(4251)) and not (layer0_outputs(4854));
    outputs(5981) <= (layer0_outputs(2550)) and (layer0_outputs(5095));
    outputs(5982) <= not(layer0_outputs(5233));
    outputs(5983) <= not((layer0_outputs(2682)) or (layer0_outputs(3474)));
    outputs(5984) <= not(layer0_outputs(363));
    outputs(5985) <= (layer0_outputs(7451)) and (layer0_outputs(3253));
    outputs(5986) <= (layer0_outputs(133)) xor (layer0_outputs(660));
    outputs(5987) <= layer0_outputs(6466);
    outputs(5988) <= (layer0_outputs(2720)) and not (layer0_outputs(2452));
    outputs(5989) <= not(layer0_outputs(3290));
    outputs(5990) <= not((layer0_outputs(1447)) xor (layer0_outputs(3910)));
    outputs(5991) <= not(layer0_outputs(704));
    outputs(5992) <= layer0_outputs(691);
    outputs(5993) <= layer0_outputs(2732);
    outputs(5994) <= not((layer0_outputs(3084)) or (layer0_outputs(2014)));
    outputs(5995) <= not(layer0_outputs(2318));
    outputs(5996) <= (layer0_outputs(1850)) and (layer0_outputs(2091));
    outputs(5997) <= not(layer0_outputs(984));
    outputs(5998) <= not(layer0_outputs(6158));
    outputs(5999) <= (layer0_outputs(1046)) and not (layer0_outputs(793));
    outputs(6000) <= not(layer0_outputs(6747));
    outputs(6001) <= (layer0_outputs(5102)) and not (layer0_outputs(5172));
    outputs(6002) <= (layer0_outputs(4004)) and (layer0_outputs(3938));
    outputs(6003) <= (layer0_outputs(1741)) and not (layer0_outputs(1798));
    outputs(6004) <= (layer0_outputs(5045)) and not (layer0_outputs(215));
    outputs(6005) <= (layer0_outputs(4757)) xor (layer0_outputs(7601));
    outputs(6006) <= layer0_outputs(538);
    outputs(6007) <= not(layer0_outputs(5122));
    outputs(6008) <= (layer0_outputs(5078)) and not (layer0_outputs(5917));
    outputs(6009) <= not((layer0_outputs(4410)) or (layer0_outputs(4517)));
    outputs(6010) <= layer0_outputs(3805);
    outputs(6011) <= not(layer0_outputs(2774)) or (layer0_outputs(4695));
    outputs(6012) <= layer0_outputs(3389);
    outputs(6013) <= not((layer0_outputs(2940)) and (layer0_outputs(2934)));
    outputs(6014) <= (layer0_outputs(3962)) xor (layer0_outputs(5378));
    outputs(6015) <= not(layer0_outputs(5345));
    outputs(6016) <= layer0_outputs(7444);
    outputs(6017) <= not(layer0_outputs(5107)) or (layer0_outputs(5484));
    outputs(6018) <= not(layer0_outputs(1807));
    outputs(6019) <= not((layer0_outputs(2894)) or (layer0_outputs(2342)));
    outputs(6020) <= not(layer0_outputs(2816));
    outputs(6021) <= (layer0_outputs(5076)) and not (layer0_outputs(1820));
    outputs(6022) <= (layer0_outputs(3586)) and not (layer0_outputs(1301));
    outputs(6023) <= (layer0_outputs(5083)) and not (layer0_outputs(4942));
    outputs(6024) <= (layer0_outputs(4413)) and not (layer0_outputs(3287));
    outputs(6025) <= layer0_outputs(1604);
    outputs(6026) <= (layer0_outputs(6108)) and (layer0_outputs(6498));
    outputs(6027) <= layer0_outputs(6651);
    outputs(6028) <= (layer0_outputs(6789)) and not (layer0_outputs(7433));
    outputs(6029) <= layer0_outputs(6234);
    outputs(6030) <= (layer0_outputs(1023)) xor (layer0_outputs(4361));
    outputs(6031) <= (layer0_outputs(105)) or (layer0_outputs(5322));
    outputs(6032) <= layer0_outputs(3132);
    outputs(6033) <= layer0_outputs(4708);
    outputs(6034) <= not(layer0_outputs(676)) or (layer0_outputs(4883));
    outputs(6035) <= layer0_outputs(2284);
    outputs(6036) <= (layer0_outputs(1618)) and (layer0_outputs(3934));
    outputs(6037) <= not(layer0_outputs(1354));
    outputs(6038) <= layer0_outputs(6406);
    outputs(6039) <= not((layer0_outputs(1979)) or (layer0_outputs(92)));
    outputs(6040) <= (layer0_outputs(736)) xor (layer0_outputs(5864));
    outputs(6041) <= (layer0_outputs(6020)) and not (layer0_outputs(3587));
    outputs(6042) <= not(layer0_outputs(1508));
    outputs(6043) <= (layer0_outputs(1124)) xor (layer0_outputs(1856));
    outputs(6044) <= not((layer0_outputs(6109)) or (layer0_outputs(3918)));
    outputs(6045) <= not(layer0_outputs(2639));
    outputs(6046) <= not((layer0_outputs(2178)) or (layer0_outputs(4440)));
    outputs(6047) <= layer0_outputs(4814);
    outputs(6048) <= (layer0_outputs(4375)) and not (layer0_outputs(3147));
    outputs(6049) <= (layer0_outputs(6164)) and not (layer0_outputs(1904));
    outputs(6050) <= layer0_outputs(211);
    outputs(6051) <= (layer0_outputs(1199)) xor (layer0_outputs(5726));
    outputs(6052) <= layer0_outputs(5000);
    outputs(6053) <= layer0_outputs(5103);
    outputs(6054) <= (layer0_outputs(6188)) and not (layer0_outputs(707));
    outputs(6055) <= not(layer0_outputs(1568));
    outputs(6056) <= (layer0_outputs(6640)) and (layer0_outputs(6296));
    outputs(6057) <= not((layer0_outputs(6722)) or (layer0_outputs(4922)));
    outputs(6058) <= layer0_outputs(1594);
    outputs(6059) <= (layer0_outputs(3778)) and not (layer0_outputs(1132));
    outputs(6060) <= layer0_outputs(1179);
    outputs(6061) <= layer0_outputs(2736);
    outputs(6062) <= not(layer0_outputs(5615));
    outputs(6063) <= layer0_outputs(2493);
    outputs(6064) <= (layer0_outputs(1166)) and not (layer0_outputs(4508));
    outputs(6065) <= not(layer0_outputs(3496));
    outputs(6066) <= (layer0_outputs(5422)) and (layer0_outputs(5102));
    outputs(6067) <= (layer0_outputs(5145)) and not (layer0_outputs(1490));
    outputs(6068) <= not((layer0_outputs(6442)) or (layer0_outputs(553)));
    outputs(6069) <= (layer0_outputs(2734)) and not (layer0_outputs(5718));
    outputs(6070) <= not((layer0_outputs(5855)) xor (layer0_outputs(4122)));
    outputs(6071) <= (layer0_outputs(2167)) xor (layer0_outputs(1287));
    outputs(6072) <= not(layer0_outputs(7248));
    outputs(6073) <= (layer0_outputs(3775)) and not (layer0_outputs(127));
    outputs(6074) <= not(layer0_outputs(7138));
    outputs(6075) <= (layer0_outputs(2488)) and (layer0_outputs(2990));
    outputs(6076) <= not((layer0_outputs(1084)) or (layer0_outputs(5587)));
    outputs(6077) <= (layer0_outputs(5937)) and not (layer0_outputs(2392));
    outputs(6078) <= (layer0_outputs(4701)) and (layer0_outputs(5360));
    outputs(6079) <= not(layer0_outputs(4619));
    outputs(6080) <= (layer0_outputs(5013)) and (layer0_outputs(322));
    outputs(6081) <= layer0_outputs(7426);
    outputs(6082) <= layer0_outputs(6791);
    outputs(6083) <= (layer0_outputs(657)) and not (layer0_outputs(1183));
    outputs(6084) <= not(layer0_outputs(4824));
    outputs(6085) <= (layer0_outputs(4732)) and not (layer0_outputs(4363));
    outputs(6086) <= layer0_outputs(3077);
    outputs(6087) <= not(layer0_outputs(5070));
    outputs(6088) <= (layer0_outputs(6222)) and (layer0_outputs(7571));
    outputs(6089) <= not(layer0_outputs(835));
    outputs(6090) <= not((layer0_outputs(1089)) or (layer0_outputs(1190)));
    outputs(6091) <= (layer0_outputs(2040)) and not (layer0_outputs(5969));
    outputs(6092) <= (layer0_outputs(5740)) and (layer0_outputs(2482));
    outputs(6093) <= not(layer0_outputs(3414));
    outputs(6094) <= not(layer0_outputs(5706));
    outputs(6095) <= not(layer0_outputs(268));
    outputs(6096) <= (layer0_outputs(3900)) and not (layer0_outputs(6876));
    outputs(6097) <= not(layer0_outputs(5993)) or (layer0_outputs(6112));
    outputs(6098) <= not(layer0_outputs(666));
    outputs(6099) <= not(layer0_outputs(2822));
    outputs(6100) <= not(layer0_outputs(1399)) or (layer0_outputs(3299));
    outputs(6101) <= layer0_outputs(6769);
    outputs(6102) <= not(layer0_outputs(3721));
    outputs(6103) <= (layer0_outputs(1959)) and not (layer0_outputs(3423));
    outputs(6104) <= layer0_outputs(4585);
    outputs(6105) <= not((layer0_outputs(1418)) or (layer0_outputs(71)));
    outputs(6106) <= layer0_outputs(2231);
    outputs(6107) <= (layer0_outputs(7005)) xor (layer0_outputs(1641));
    outputs(6108) <= not(layer0_outputs(3255));
    outputs(6109) <= layer0_outputs(1030);
    outputs(6110) <= (layer0_outputs(1324)) and not (layer0_outputs(3979));
    outputs(6111) <= (layer0_outputs(7362)) and not (layer0_outputs(3735));
    outputs(6112) <= (layer0_outputs(5290)) and not (layer0_outputs(4781));
    outputs(6113) <= (layer0_outputs(3846)) and not (layer0_outputs(1407));
    outputs(6114) <= not(layer0_outputs(4176));
    outputs(6115) <= layer0_outputs(1790);
    outputs(6116) <= not(layer0_outputs(191));
    outputs(6117) <= not(layer0_outputs(5527));
    outputs(6118) <= (layer0_outputs(3276)) xor (layer0_outputs(7130));
    outputs(6119) <= (layer0_outputs(1897)) or (layer0_outputs(1376));
    outputs(6120) <= (layer0_outputs(3904)) and not (layer0_outputs(6035));
    outputs(6121) <= (layer0_outputs(2678)) xor (layer0_outputs(5919));
    outputs(6122) <= not((layer0_outputs(4066)) xor (layer0_outputs(7149)));
    outputs(6123) <= layer0_outputs(6281);
    outputs(6124) <= not((layer0_outputs(650)) or (layer0_outputs(7533)));
    outputs(6125) <= (layer0_outputs(412)) and (layer0_outputs(4527));
    outputs(6126) <= not((layer0_outputs(2277)) xor (layer0_outputs(1564)));
    outputs(6127) <= layer0_outputs(4944);
    outputs(6128) <= (layer0_outputs(3599)) and not (layer0_outputs(3407));
    outputs(6129) <= layer0_outputs(917);
    outputs(6130) <= (layer0_outputs(7080)) and (layer0_outputs(824));
    outputs(6131) <= layer0_outputs(1174);
    outputs(6132) <= (layer0_outputs(1454)) and not (layer0_outputs(1145));
    outputs(6133) <= (layer0_outputs(757)) xor (layer0_outputs(1922));
    outputs(6134) <= (layer0_outputs(275)) and not (layer0_outputs(592));
    outputs(6135) <= (layer0_outputs(6055)) xor (layer0_outputs(44));
    outputs(6136) <= not(layer0_outputs(74));
    outputs(6137) <= not(layer0_outputs(6533));
    outputs(6138) <= layer0_outputs(6439);
    outputs(6139) <= (layer0_outputs(743)) and not (layer0_outputs(441));
    outputs(6140) <= layer0_outputs(5656);
    outputs(6141) <= not(layer0_outputs(2357));
    outputs(6142) <= not((layer0_outputs(4955)) or (layer0_outputs(3897)));
    outputs(6143) <= (layer0_outputs(4759)) and not (layer0_outputs(6758));
    outputs(6144) <= (layer0_outputs(7563)) and not (layer0_outputs(756));
    outputs(6145) <= not((layer0_outputs(1663)) and (layer0_outputs(5893)));
    outputs(6146) <= layer0_outputs(1462);
    outputs(6147) <= not(layer0_outputs(579)) or (layer0_outputs(5770));
    outputs(6148) <= layer0_outputs(2815);
    outputs(6149) <= not(layer0_outputs(3268));
    outputs(6150) <= layer0_outputs(4109);
    outputs(6151) <= (layer0_outputs(5469)) and not (layer0_outputs(2460));
    outputs(6152) <= not(layer0_outputs(2892)) or (layer0_outputs(6773));
    outputs(6153) <= not((layer0_outputs(1021)) xor (layer0_outputs(2741)));
    outputs(6154) <= (layer0_outputs(3438)) or (layer0_outputs(656));
    outputs(6155) <= layer0_outputs(2927);
    outputs(6156) <= not((layer0_outputs(4506)) and (layer0_outputs(1388)));
    outputs(6157) <= layer0_outputs(6990);
    outputs(6158) <= not((layer0_outputs(5429)) xor (layer0_outputs(3202)));
    outputs(6159) <= layer0_outputs(7560);
    outputs(6160) <= not(layer0_outputs(5839)) or (layer0_outputs(2988));
    outputs(6161) <= not((layer0_outputs(5558)) or (layer0_outputs(4429)));
    outputs(6162) <= not(layer0_outputs(7663));
    outputs(6163) <= layer0_outputs(6291);
    outputs(6164) <= not(layer0_outputs(6038)) or (layer0_outputs(2521));
    outputs(6165) <= layer0_outputs(2902);
    outputs(6166) <= (layer0_outputs(1709)) xor (layer0_outputs(3702));
    outputs(6167) <= layer0_outputs(5957);
    outputs(6168) <= layer0_outputs(327);
    outputs(6169) <= not((layer0_outputs(7320)) and (layer0_outputs(2608)));
    outputs(6170) <= not(layer0_outputs(4881));
    outputs(6171) <= not((layer0_outputs(341)) xor (layer0_outputs(4482)));
    outputs(6172) <= layer0_outputs(1395);
    outputs(6173) <= (layer0_outputs(6863)) xor (layer0_outputs(3521));
    outputs(6174) <= (layer0_outputs(1010)) or (layer0_outputs(1007));
    outputs(6175) <= not((layer0_outputs(7493)) xor (layer0_outputs(4745)));
    outputs(6176) <= not((layer0_outputs(6723)) or (layer0_outputs(1739)));
    outputs(6177) <= not((layer0_outputs(3352)) xor (layer0_outputs(2373)));
    outputs(6178) <= not(layer0_outputs(1734));
    outputs(6179) <= not(layer0_outputs(6583)) or (layer0_outputs(5403));
    outputs(6180) <= layer0_outputs(4526);
    outputs(6181) <= (layer0_outputs(3818)) or (layer0_outputs(588));
    outputs(6182) <= layer0_outputs(1654);
    outputs(6183) <= layer0_outputs(4701);
    outputs(6184) <= not(layer0_outputs(2399)) or (layer0_outputs(6361));
    outputs(6185) <= not(layer0_outputs(916));
    outputs(6186) <= layer0_outputs(876);
    outputs(6187) <= not(layer0_outputs(7124));
    outputs(6188) <= not(layer0_outputs(2975));
    outputs(6189) <= not((layer0_outputs(5278)) or (layer0_outputs(2935)));
    outputs(6190) <= not(layer0_outputs(7114));
    outputs(6191) <= (layer0_outputs(122)) xor (layer0_outputs(7558));
    outputs(6192) <= not((layer0_outputs(4121)) xor (layer0_outputs(6986)));
    outputs(6193) <= layer0_outputs(610);
    outputs(6194) <= (layer0_outputs(2434)) and not (layer0_outputs(1989));
    outputs(6195) <= (layer0_outputs(649)) or (layer0_outputs(1148));
    outputs(6196) <= not(layer0_outputs(3419)) or (layer0_outputs(7405));
    outputs(6197) <= layer0_outputs(2135);
    outputs(6198) <= (layer0_outputs(6491)) xor (layer0_outputs(6054));
    outputs(6199) <= not((layer0_outputs(6731)) or (layer0_outputs(4508)));
    outputs(6200) <= not((layer0_outputs(3290)) xor (layer0_outputs(6647)));
    outputs(6201) <= layer0_outputs(6056);
    outputs(6202) <= layer0_outputs(296);
    outputs(6203) <= layer0_outputs(2632);
    outputs(6204) <= not(layer0_outputs(3787));
    outputs(6205) <= (layer0_outputs(3098)) or (layer0_outputs(7123));
    outputs(6206) <= layer0_outputs(802);
    outputs(6207) <= (layer0_outputs(6617)) or (layer0_outputs(408));
    outputs(6208) <= not((layer0_outputs(2489)) xor (layer0_outputs(2717)));
    outputs(6209) <= (layer0_outputs(272)) and not (layer0_outputs(5285));
    outputs(6210) <= not((layer0_outputs(7359)) and (layer0_outputs(3551)));
    outputs(6211) <= not((layer0_outputs(4632)) and (layer0_outputs(2124)));
    outputs(6212) <= not(layer0_outputs(4279));
    outputs(6213) <= (layer0_outputs(5535)) xor (layer0_outputs(4125));
    outputs(6214) <= not((layer0_outputs(7600)) and (layer0_outputs(6120)));
    outputs(6215) <= not((layer0_outputs(5709)) xor (layer0_outputs(3343)));
    outputs(6216) <= (layer0_outputs(359)) and (layer0_outputs(4424));
    outputs(6217) <= not(layer0_outputs(647));
    outputs(6218) <= not(layer0_outputs(6029));
    outputs(6219) <= (layer0_outputs(1590)) and not (layer0_outputs(1676));
    outputs(6220) <= not((layer0_outputs(7302)) and (layer0_outputs(1029)));
    outputs(6221) <= not((layer0_outputs(5675)) or (layer0_outputs(1936)));
    outputs(6222) <= not(layer0_outputs(3109)) or (layer0_outputs(919));
    outputs(6223) <= (layer0_outputs(4668)) or (layer0_outputs(2973));
    outputs(6224) <= not(layer0_outputs(2450));
    outputs(6225) <= (layer0_outputs(4833)) or (layer0_outputs(3752));
    outputs(6226) <= not((layer0_outputs(3066)) or (layer0_outputs(7249)));
    outputs(6227) <= layer0_outputs(2565);
    outputs(6228) <= not(layer0_outputs(369));
    outputs(6229) <= not(layer0_outputs(4983));
    outputs(6230) <= not(layer0_outputs(3854));
    outputs(6231) <= layer0_outputs(3600);
    outputs(6232) <= not(layer0_outputs(7286));
    outputs(6233) <= not(layer0_outputs(1028));
    outputs(6234) <= not(layer0_outputs(3782));
    outputs(6235) <= not((layer0_outputs(7381)) xor (layer0_outputs(315)));
    outputs(6236) <= not(layer0_outputs(6425)) or (layer0_outputs(1351));
    outputs(6237) <= not((layer0_outputs(2803)) xor (layer0_outputs(3497)));
    outputs(6238) <= layer0_outputs(6042);
    outputs(6239) <= not(layer0_outputs(3239));
    outputs(6240) <= not(layer0_outputs(1027));
    outputs(6241) <= not(layer0_outputs(7659)) or (layer0_outputs(5280));
    outputs(6242) <= not(layer0_outputs(2436));
    outputs(6243) <= (layer0_outputs(3973)) xor (layer0_outputs(16));
    outputs(6244) <= (layer0_outputs(7208)) xor (layer0_outputs(3402));
    outputs(6245) <= layer0_outputs(7056);
    outputs(6246) <= (layer0_outputs(7204)) xor (layer0_outputs(6157));
    outputs(6247) <= layer0_outputs(3797);
    outputs(6248) <= (layer0_outputs(6641)) xor (layer0_outputs(862));
    outputs(6249) <= (layer0_outputs(2072)) and not (layer0_outputs(2554));
    outputs(6250) <= (layer0_outputs(6006)) or (layer0_outputs(6487));
    outputs(6251) <= layer0_outputs(4860);
    outputs(6252) <= layer0_outputs(6053);
    outputs(6253) <= layer0_outputs(7582);
    outputs(6254) <= layer0_outputs(2285);
    outputs(6255) <= not(layer0_outputs(4537));
    outputs(6256) <= (layer0_outputs(3382)) and not (layer0_outputs(6592));
    outputs(6257) <= not((layer0_outputs(3978)) and (layer0_outputs(1941)));
    outputs(6258) <= (layer0_outputs(5381)) and not (layer0_outputs(587));
    outputs(6259) <= layer0_outputs(674);
    outputs(6260) <= (layer0_outputs(3801)) and (layer0_outputs(2558));
    outputs(6261) <= not(layer0_outputs(2389));
    outputs(6262) <= (layer0_outputs(1230)) xor (layer0_outputs(5433));
    outputs(6263) <= not((layer0_outputs(6602)) xor (layer0_outputs(376)));
    outputs(6264) <= layer0_outputs(3801);
    outputs(6265) <= not(layer0_outputs(3354));
    outputs(6266) <= (layer0_outputs(1929)) xor (layer0_outputs(6016));
    outputs(6267) <= (layer0_outputs(1062)) or (layer0_outputs(3388));
    outputs(6268) <= (layer0_outputs(3714)) and (layer0_outputs(4586));
    outputs(6269) <= not((layer0_outputs(5626)) xor (layer0_outputs(5984)));
    outputs(6270) <= layer0_outputs(5686);
    outputs(6271) <= (layer0_outputs(3740)) xor (layer0_outputs(6128));
    outputs(6272) <= not((layer0_outputs(3489)) xor (layer0_outputs(4864)));
    outputs(6273) <= not(layer0_outputs(6380));
    outputs(6274) <= (layer0_outputs(6399)) and not (layer0_outputs(7465));
    outputs(6275) <= (layer0_outputs(6399)) and not (layer0_outputs(628));
    outputs(6276) <= not((layer0_outputs(3106)) and (layer0_outputs(5953)));
    outputs(6277) <= not(layer0_outputs(1506)) or (layer0_outputs(1168));
    outputs(6278) <= layer0_outputs(2312);
    outputs(6279) <= not(layer0_outputs(1176));
    outputs(6280) <= not((layer0_outputs(4456)) and (layer0_outputs(1245)));
    outputs(6281) <= (layer0_outputs(4739)) xor (layer0_outputs(5213));
    outputs(6282) <= not((layer0_outputs(5557)) and (layer0_outputs(4786)));
    outputs(6283) <= not((layer0_outputs(1162)) xor (layer0_outputs(5935)));
    outputs(6284) <= not(layer0_outputs(5974)) or (layer0_outputs(812));
    outputs(6285) <= layer0_outputs(7416);
    outputs(6286) <= layer0_outputs(5834);
    outputs(6287) <= not(layer0_outputs(617));
    outputs(6288) <= not(layer0_outputs(934));
    outputs(6289) <= not(layer0_outputs(5756));
    outputs(6290) <= layer0_outputs(583);
    outputs(6291) <= not(layer0_outputs(470)) or (layer0_outputs(725));
    outputs(6292) <= not((layer0_outputs(6285)) and (layer0_outputs(4691)));
    outputs(6293) <= not(layer0_outputs(1974));
    outputs(6294) <= not(layer0_outputs(1152)) or (layer0_outputs(3368));
    outputs(6295) <= not(layer0_outputs(3936)) or (layer0_outputs(3112));
    outputs(6296) <= (layer0_outputs(2737)) and not (layer0_outputs(6903));
    outputs(6297) <= not((layer0_outputs(5698)) xor (layer0_outputs(6940)));
    outputs(6298) <= not(layer0_outputs(3720)) or (layer0_outputs(2321));
    outputs(6299) <= layer0_outputs(5007);
    outputs(6300) <= (layer0_outputs(6180)) and (layer0_outputs(2486));
    outputs(6301) <= not((layer0_outputs(2306)) or (layer0_outputs(1733)));
    outputs(6302) <= (layer0_outputs(68)) or (layer0_outputs(5323));
    outputs(6303) <= not(layer0_outputs(1606));
    outputs(6304) <= (layer0_outputs(7469)) or (layer0_outputs(5835));
    outputs(6305) <= (layer0_outputs(1387)) or (layer0_outputs(4676));
    outputs(6306) <= not(layer0_outputs(5130));
    outputs(6307) <= not(layer0_outputs(2604));
    outputs(6308) <= not((layer0_outputs(6609)) xor (layer0_outputs(861)));
    outputs(6309) <= not(layer0_outputs(3504)) or (layer0_outputs(3577));
    outputs(6310) <= (layer0_outputs(5871)) and not (layer0_outputs(7606));
    outputs(6311) <= (layer0_outputs(2052)) or (layer0_outputs(6192));
    outputs(6312) <= not(layer0_outputs(6278));
    outputs(6313) <= layer0_outputs(5530);
    outputs(6314) <= not((layer0_outputs(2680)) or (layer0_outputs(6081)));
    outputs(6315) <= not(layer0_outputs(6960)) or (layer0_outputs(4425));
    outputs(6316) <= not(layer0_outputs(4822));
    outputs(6317) <= not(layer0_outputs(4522));
    outputs(6318) <= not(layer0_outputs(2482));
    outputs(6319) <= not(layer0_outputs(7168));
    outputs(6320) <= not((layer0_outputs(4122)) xor (layer0_outputs(3042)));
    outputs(6321) <= not(layer0_outputs(6998));
    outputs(6322) <= (layer0_outputs(6433)) xor (layer0_outputs(5726));
    outputs(6323) <= not((layer0_outputs(2089)) and (layer0_outputs(5472)));
    outputs(6324) <= not(layer0_outputs(3214));
    outputs(6325) <= (layer0_outputs(841)) and not (layer0_outputs(2355));
    outputs(6326) <= not((layer0_outputs(5661)) xor (layer0_outputs(5624)));
    outputs(6327) <= (layer0_outputs(2137)) and (layer0_outputs(4552));
    outputs(6328) <= layer0_outputs(2110);
    outputs(6329) <= not(layer0_outputs(521));
    outputs(6330) <= not(layer0_outputs(309));
    outputs(6331) <= not((layer0_outputs(4347)) or (layer0_outputs(7419)));
    outputs(6332) <= layer0_outputs(2982);
    outputs(6333) <= not((layer0_outputs(1825)) and (layer0_outputs(2549)));
    outputs(6334) <= not(layer0_outputs(6776)) or (layer0_outputs(848));
    outputs(6335) <= not(layer0_outputs(2943)) or (layer0_outputs(171));
    outputs(6336) <= not(layer0_outputs(2062));
    outputs(6337) <= not((layer0_outputs(5142)) xor (layer0_outputs(7014)));
    outputs(6338) <= layer0_outputs(7399);
    outputs(6339) <= not(layer0_outputs(4355));
    outputs(6340) <= not((layer0_outputs(7138)) xor (layer0_outputs(6532)));
    outputs(6341) <= layer0_outputs(4764);
    outputs(6342) <= not(layer0_outputs(2028));
    outputs(6343) <= not((layer0_outputs(5147)) and (layer0_outputs(3769)));
    outputs(6344) <= not((layer0_outputs(3498)) or (layer0_outputs(198)));
    outputs(6345) <= not((layer0_outputs(798)) xor (layer0_outputs(7577)));
    outputs(6346) <= layer0_outputs(581);
    outputs(6347) <= (layer0_outputs(3638)) and not (layer0_outputs(5097));
    outputs(6348) <= not((layer0_outputs(2578)) xor (layer0_outputs(4654)));
    outputs(6349) <= not(layer0_outputs(64)) or (layer0_outputs(2891));
    outputs(6350) <= not(layer0_outputs(4504));
    outputs(6351) <= not((layer0_outputs(2005)) and (layer0_outputs(7538)));
    outputs(6352) <= (layer0_outputs(6938)) xor (layer0_outputs(893));
    outputs(6353) <= (layer0_outputs(5634)) xor (layer0_outputs(4004));
    outputs(6354) <= not(layer0_outputs(3582));
    outputs(6355) <= (layer0_outputs(2637)) and not (layer0_outputs(5648));
    outputs(6356) <= not((layer0_outputs(1924)) and (layer0_outputs(2476)));
    outputs(6357) <= layer0_outputs(884);
    outputs(6358) <= layer0_outputs(6492);
    outputs(6359) <= not(layer0_outputs(6107)) or (layer0_outputs(527));
    outputs(6360) <= (layer0_outputs(6007)) xor (layer0_outputs(6228));
    outputs(6361) <= (layer0_outputs(952)) xor (layer0_outputs(1273));
    outputs(6362) <= (layer0_outputs(4982)) xor (layer0_outputs(4660));
    outputs(6363) <= not(layer0_outputs(1349));
    outputs(6364) <= not(layer0_outputs(6959)) or (layer0_outputs(5819));
    outputs(6365) <= not((layer0_outputs(6046)) xor (layer0_outputs(7208)));
    outputs(6366) <= not(layer0_outputs(4442));
    outputs(6367) <= not(layer0_outputs(1489)) or (layer0_outputs(6006));
    outputs(6368) <= not(layer0_outputs(3035)) or (layer0_outputs(293));
    outputs(6369) <= not(layer0_outputs(106)) or (layer0_outputs(1758));
    outputs(6370) <= layer0_outputs(7273);
    outputs(6371) <= layer0_outputs(5852);
    outputs(6372) <= layer0_outputs(568);
    outputs(6373) <= not(layer0_outputs(1098));
    outputs(6374) <= layer0_outputs(6499);
    outputs(6375) <= (layer0_outputs(1575)) or (layer0_outputs(2298));
    outputs(6376) <= (layer0_outputs(5193)) xor (layer0_outputs(7041));
    outputs(6377) <= not((layer0_outputs(1707)) or (layer0_outputs(5203)));
    outputs(6378) <= not((layer0_outputs(4752)) xor (layer0_outputs(1857)));
    outputs(6379) <= (layer0_outputs(6674)) xor (layer0_outputs(361));
    outputs(6380) <= not(layer0_outputs(2616)) or (layer0_outputs(1561));
    outputs(6381) <= not((layer0_outputs(398)) or (layer0_outputs(2200)));
    outputs(6382) <= not((layer0_outputs(7304)) and (layer0_outputs(283)));
    outputs(6383) <= not(layer0_outputs(1997)) or (layer0_outputs(6102));
    outputs(6384) <= not((layer0_outputs(4866)) xor (layer0_outputs(1120)));
    outputs(6385) <= not(layer0_outputs(1519));
    outputs(6386) <= not((layer0_outputs(4914)) xor (layer0_outputs(1721)));
    outputs(6387) <= not(layer0_outputs(3350)) or (layer0_outputs(3367));
    outputs(6388) <= layer0_outputs(1934);
    outputs(6389) <= not((layer0_outputs(4263)) xor (layer0_outputs(4728)));
    outputs(6390) <= (layer0_outputs(5292)) xor (layer0_outputs(547));
    outputs(6391) <= layer0_outputs(3680);
    outputs(6392) <= not(layer0_outputs(6535));
    outputs(6393) <= (layer0_outputs(18)) xor (layer0_outputs(4818));
    outputs(6394) <= layer0_outputs(1937);
    outputs(6395) <= not(layer0_outputs(7411)) or (layer0_outputs(4195));
    outputs(6396) <= layer0_outputs(3660);
    outputs(6397) <= not(layer0_outputs(2071));
    outputs(6398) <= not(layer0_outputs(6044)) or (layer0_outputs(4720));
    outputs(6399) <= not(layer0_outputs(2865));
    outputs(6400) <= layer0_outputs(4906);
    outputs(6401) <= (layer0_outputs(3056)) xor (layer0_outputs(6614));
    outputs(6402) <= (layer0_outputs(4461)) and not (layer0_outputs(4365));
    outputs(6403) <= layer0_outputs(2579);
    outputs(6404) <= (layer0_outputs(1282)) and (layer0_outputs(849));
    outputs(6405) <= not(layer0_outputs(1549)) or (layer0_outputs(1181));
    outputs(6406) <= (layer0_outputs(6288)) or (layer0_outputs(6858));
    outputs(6407) <= (layer0_outputs(5882)) and not (layer0_outputs(3544));
    outputs(6408) <= not(layer0_outputs(273));
    outputs(6409) <= not((layer0_outputs(2180)) xor (layer0_outputs(7117)));
    outputs(6410) <= layer0_outputs(426);
    outputs(6411) <= layer0_outputs(6090);
    outputs(6412) <= (layer0_outputs(5402)) xor (layer0_outputs(2081));
    outputs(6413) <= not(layer0_outputs(4530));
    outputs(6414) <= not(layer0_outputs(6540));
    outputs(6415) <= layer0_outputs(7365);
    outputs(6416) <= not(layer0_outputs(6966));
    outputs(6417) <= not(layer0_outputs(3646));
    outputs(6418) <= layer0_outputs(6438);
    outputs(6419) <= (layer0_outputs(2928)) and not (layer0_outputs(2419));
    outputs(6420) <= not((layer0_outputs(5254)) xor (layer0_outputs(5594)));
    outputs(6421) <= not((layer0_outputs(7610)) xor (layer0_outputs(2524)));
    outputs(6422) <= not(layer0_outputs(4900)) or (layer0_outputs(1582));
    outputs(6423) <= not((layer0_outputs(2876)) or (layer0_outputs(3514)));
    outputs(6424) <= (layer0_outputs(1779)) xor (layer0_outputs(4883));
    outputs(6425) <= layer0_outputs(1079);
    outputs(6426) <= not((layer0_outputs(7469)) xor (layer0_outputs(5118)));
    outputs(6427) <= not(layer0_outputs(1307)) or (layer0_outputs(5787));
    outputs(6428) <= layer0_outputs(1461);
    outputs(6429) <= (layer0_outputs(2669)) and not (layer0_outputs(4559));
    outputs(6430) <= not((layer0_outputs(1420)) xor (layer0_outputs(2918)));
    outputs(6431) <= not((layer0_outputs(2990)) xor (layer0_outputs(2065)));
    outputs(6432) <= (layer0_outputs(971)) or (layer0_outputs(3596));
    outputs(6433) <= not(layer0_outputs(3562)) or (layer0_outputs(5412));
    outputs(6434) <= not(layer0_outputs(21)) or (layer0_outputs(246));
    outputs(6435) <= (layer0_outputs(5306)) and (layer0_outputs(4607));
    outputs(6436) <= not((layer0_outputs(4273)) and (layer0_outputs(401)));
    outputs(6437) <= not(layer0_outputs(719));
    outputs(6438) <= layer0_outputs(747);
    outputs(6439) <= not(layer0_outputs(3831));
    outputs(6440) <= (layer0_outputs(3323)) or (layer0_outputs(1178));
    outputs(6441) <= layer0_outputs(2191);
    outputs(6442) <= (layer0_outputs(3240)) xor (layer0_outputs(1574));
    outputs(6443) <= (layer0_outputs(7571)) and not (layer0_outputs(3083));
    outputs(6444) <= not(layer0_outputs(3955));
    outputs(6445) <= (layer0_outputs(2509)) xor (layer0_outputs(209));
    outputs(6446) <= layer0_outputs(7173);
    outputs(6447) <= not(layer0_outputs(3849));
    outputs(6448) <= not((layer0_outputs(6921)) or (layer0_outputs(2806)));
    outputs(6449) <= not(layer0_outputs(3694));
    outputs(6450) <= layer0_outputs(1240);
    outputs(6451) <= not(layer0_outputs(2508)) or (layer0_outputs(6161));
    outputs(6452) <= (layer0_outputs(7047)) xor (layer0_outputs(4929));
    outputs(6453) <= (layer0_outputs(3116)) or (layer0_outputs(610));
    outputs(6454) <= layer0_outputs(5671);
    outputs(6455) <= (layer0_outputs(943)) xor (layer0_outputs(7244));
    outputs(6456) <= layer0_outputs(7197);
    outputs(6457) <= layer0_outputs(111);
    outputs(6458) <= not(layer0_outputs(1281));
    outputs(6459) <= not((layer0_outputs(4584)) xor (layer0_outputs(4715)));
    outputs(6460) <= not((layer0_outputs(1783)) and (layer0_outputs(1890)));
    outputs(6461) <= not(layer0_outputs(339));
    outputs(6462) <= (layer0_outputs(1545)) and not (layer0_outputs(6639));
    outputs(6463) <= not((layer0_outputs(4007)) xor (layer0_outputs(2422)));
    outputs(6464) <= not(layer0_outputs(4039)) or (layer0_outputs(6667));
    outputs(6465) <= not((layer0_outputs(2725)) and (layer0_outputs(2242)));
    outputs(6466) <= layer0_outputs(6260);
    outputs(6467) <= (layer0_outputs(6576)) and not (layer0_outputs(6716));
    outputs(6468) <= (layer0_outputs(2921)) and (layer0_outputs(5961));
    outputs(6469) <= layer0_outputs(2070);
    outputs(6470) <= not(layer0_outputs(6507)) or (layer0_outputs(3546));
    outputs(6471) <= layer0_outputs(1232);
    outputs(6472) <= layer0_outputs(1883);
    outputs(6473) <= (layer0_outputs(2801)) xor (layer0_outputs(5932));
    outputs(6474) <= (layer0_outputs(4213)) and not (layer0_outputs(4545));
    outputs(6475) <= (layer0_outputs(2592)) and not (layer0_outputs(3762));
    outputs(6476) <= not(layer0_outputs(7606));
    outputs(6477) <= layer0_outputs(3447);
    outputs(6478) <= not((layer0_outputs(3063)) xor (layer0_outputs(5775)));
    outputs(6479) <= not((layer0_outputs(116)) and (layer0_outputs(3953)));
    outputs(6480) <= not((layer0_outputs(6628)) xor (layer0_outputs(2296)));
    outputs(6481) <= not((layer0_outputs(2186)) xor (layer0_outputs(5330)));
    outputs(6482) <= layer0_outputs(4200);
    outputs(6483) <= not((layer0_outputs(879)) or (layer0_outputs(5480)));
    outputs(6484) <= (layer0_outputs(4467)) or (layer0_outputs(1282));
    outputs(6485) <= (layer0_outputs(5850)) xor (layer0_outputs(799));
    outputs(6486) <= not(layer0_outputs(5095));
    outputs(6487) <= layer0_outputs(2753);
    outputs(6488) <= not(layer0_outputs(2261));
    outputs(6489) <= layer0_outputs(6565);
    outputs(6490) <= (layer0_outputs(459)) and not (layer0_outputs(5480));
    outputs(6491) <= (layer0_outputs(1806)) and (layer0_outputs(2667));
    outputs(6492) <= not((layer0_outputs(4377)) xor (layer0_outputs(5432)));
    outputs(6493) <= layer0_outputs(2646);
    outputs(6494) <= layer0_outputs(3365);
    outputs(6495) <= (layer0_outputs(1208)) xor (layer0_outputs(4397));
    outputs(6496) <= (layer0_outputs(4910)) or (layer0_outputs(3429));
    outputs(6497) <= (layer0_outputs(6418)) xor (layer0_outputs(3909));
    outputs(6498) <= layer0_outputs(4005);
    outputs(6499) <= not(layer0_outputs(1164)) or (layer0_outputs(180));
    outputs(6500) <= not((layer0_outputs(7379)) and (layer0_outputs(5630)));
    outputs(6501) <= (layer0_outputs(1565)) and not (layer0_outputs(2408));
    outputs(6502) <= not((layer0_outputs(900)) xor (layer0_outputs(855)));
    outputs(6503) <= not((layer0_outputs(5045)) and (layer0_outputs(4382)));
    outputs(6504) <= not(layer0_outputs(2128)) or (layer0_outputs(1449));
    outputs(6505) <= not(layer0_outputs(1059)) or (layer0_outputs(881));
    outputs(6506) <= layer0_outputs(644);
    outputs(6507) <= (layer0_outputs(89)) xor (layer0_outputs(5124));
    outputs(6508) <= not((layer0_outputs(4615)) xor (layer0_outputs(2857)));
    outputs(6509) <= not(layer0_outputs(5471));
    outputs(6510) <= not((layer0_outputs(4608)) and (layer0_outputs(1033)));
    outputs(6511) <= (layer0_outputs(863)) xor (layer0_outputs(7468));
    outputs(6512) <= not(layer0_outputs(5824));
    outputs(6513) <= not((layer0_outputs(2617)) xor (layer0_outputs(5435)));
    outputs(6514) <= not((layer0_outputs(4251)) xor (layer0_outputs(2400)));
    outputs(6515) <= (layer0_outputs(877)) xor (layer0_outputs(1190));
    outputs(6516) <= (layer0_outputs(2188)) xor (layer0_outputs(6341));
    outputs(6517) <= (layer0_outputs(3320)) and (layer0_outputs(5575));
    outputs(6518) <= not(layer0_outputs(3842));
    outputs(6519) <= layer0_outputs(6802);
    outputs(6520) <= (layer0_outputs(6676)) xor (layer0_outputs(3294));
    outputs(6521) <= (layer0_outputs(1983)) and not (layer0_outputs(5578));
    outputs(6522) <= (layer0_outputs(367)) and not (layer0_outputs(22));
    outputs(6523) <= (layer0_outputs(7153)) and (layer0_outputs(2774));
    outputs(6524) <= (layer0_outputs(4149)) xor (layer0_outputs(6066));
    outputs(6525) <= not((layer0_outputs(3874)) xor (layer0_outputs(6207)));
    outputs(6526) <= not((layer0_outputs(2183)) xor (layer0_outputs(3866)));
    outputs(6527) <= not(layer0_outputs(6857)) or (layer0_outputs(2871));
    outputs(6528) <= not(layer0_outputs(2991));
    outputs(6529) <= not((layer0_outputs(355)) xor (layer0_outputs(6132)));
    outputs(6530) <= (layer0_outputs(3484)) and not (layer0_outputs(3028));
    outputs(6531) <= (layer0_outputs(3058)) or (layer0_outputs(7633));
    outputs(6532) <= not(layer0_outputs(439));
    outputs(6533) <= not(layer0_outputs(2831)) or (layer0_outputs(7440));
    outputs(6534) <= not(layer0_outputs(6417)) or (layer0_outputs(6605));
    outputs(6535) <= layer0_outputs(6088);
    outputs(6536) <= not(layer0_outputs(6889)) or (layer0_outputs(4629));
    outputs(6537) <= not(layer0_outputs(3355));
    outputs(6538) <= not(layer0_outputs(6105)) or (layer0_outputs(4123));
    outputs(6539) <= (layer0_outputs(503)) and (layer0_outputs(1971));
    outputs(6540) <= not(layer0_outputs(3708));
    outputs(6541) <= not(layer0_outputs(5596)) or (layer0_outputs(4286));
    outputs(6542) <= (layer0_outputs(6904)) xor (layer0_outputs(2805));
    outputs(6543) <= not((layer0_outputs(3428)) and (layer0_outputs(5120)));
    outputs(6544) <= not(layer0_outputs(5586));
    outputs(6545) <= (layer0_outputs(4570)) and not (layer0_outputs(895));
    outputs(6546) <= (layer0_outputs(137)) and not (layer0_outputs(455));
    outputs(6547) <= layer0_outputs(2143);
    outputs(6548) <= not(layer0_outputs(2341)) or (layer0_outputs(7059));
    outputs(6549) <= layer0_outputs(4041);
    outputs(6550) <= layer0_outputs(1121);
    outputs(6551) <= not((layer0_outputs(5236)) and (layer0_outputs(7263)));
    outputs(6552) <= (layer0_outputs(4434)) and (layer0_outputs(3668));
    outputs(6553) <= layer0_outputs(5205);
    outputs(6554) <= not(layer0_outputs(4128)) or (layer0_outputs(2002));
    outputs(6555) <= not(layer0_outputs(4297)) or (layer0_outputs(918));
    outputs(6556) <= layer0_outputs(5143);
    outputs(6557) <= layer0_outputs(932);
    outputs(6558) <= (layer0_outputs(7222)) xor (layer0_outputs(3197));
    outputs(6559) <= layer0_outputs(51);
    outputs(6560) <= not(layer0_outputs(3192)) or (layer0_outputs(2451));
    outputs(6561) <= not((layer0_outputs(4063)) xor (layer0_outputs(2460)));
    outputs(6562) <= (layer0_outputs(524)) and not (layer0_outputs(350));
    outputs(6563) <= (layer0_outputs(357)) xor (layer0_outputs(7114));
    outputs(6564) <= not(layer0_outputs(1297));
    outputs(6565) <= not((layer0_outputs(3536)) or (layer0_outputs(5064)));
    outputs(6566) <= layer0_outputs(1352);
    outputs(6567) <= not(layer0_outputs(1651));
    outputs(6568) <= (layer0_outputs(1852)) xor (layer0_outputs(5239));
    outputs(6569) <= not(layer0_outputs(4374));
    outputs(6570) <= not((layer0_outputs(1314)) xor (layer0_outputs(3747)));
    outputs(6571) <= not(layer0_outputs(1760));
    outputs(6572) <= (layer0_outputs(4451)) xor (layer0_outputs(4609));
    outputs(6573) <= (layer0_outputs(856)) xor (layer0_outputs(2922));
    outputs(6574) <= layer0_outputs(2913);
    outputs(6575) <= not((layer0_outputs(7532)) xor (layer0_outputs(559)));
    outputs(6576) <= (layer0_outputs(4484)) and not (layer0_outputs(7559));
    outputs(6577) <= (layer0_outputs(7171)) xor (layer0_outputs(3891));
    outputs(6578) <= (layer0_outputs(6191)) or (layer0_outputs(5926));
    outputs(6579) <= not(layer0_outputs(4124));
    outputs(6580) <= not((layer0_outputs(2755)) and (layer0_outputs(6105)));
    outputs(6581) <= not(layer0_outputs(6731));
    outputs(6582) <= not((layer0_outputs(6018)) or (layer0_outputs(3723)));
    outputs(6583) <= (layer0_outputs(5994)) or (layer0_outputs(1632));
    outputs(6584) <= not((layer0_outputs(5071)) and (layer0_outputs(1557)));
    outputs(6585) <= (layer0_outputs(3799)) or (layer0_outputs(4238));
    outputs(6586) <= not(layer0_outputs(6789)) or (layer0_outputs(1953));
    outputs(6587) <= not((layer0_outputs(7564)) xor (layer0_outputs(1716)));
    outputs(6588) <= not(layer0_outputs(4503));
    outputs(6589) <= layer0_outputs(5607);
    outputs(6590) <= (layer0_outputs(1412)) xor (layer0_outputs(86));
    outputs(6591) <= not((layer0_outputs(2789)) xor (layer0_outputs(7463)));
    outputs(6592) <= (layer0_outputs(1281)) xor (layer0_outputs(2340));
    outputs(6593) <= not((layer0_outputs(3099)) and (layer0_outputs(5579)));
    outputs(6594) <= not(layer0_outputs(4787));
    outputs(6595) <= not(layer0_outputs(7394));
    outputs(6596) <= (layer0_outputs(417)) or (layer0_outputs(6389));
    outputs(6597) <= not(layer0_outputs(3530));
    outputs(6598) <= not(layer0_outputs(1421)) or (layer0_outputs(2420));
    outputs(6599) <= not(layer0_outputs(2839)) or (layer0_outputs(6819));
    outputs(6600) <= not(layer0_outputs(2918));
    outputs(6601) <= not(layer0_outputs(7409)) or (layer0_outputs(4794));
    outputs(6602) <= not(layer0_outputs(1754)) or (layer0_outputs(3079));
    outputs(6603) <= layer0_outputs(1201);
    outputs(6604) <= not((layer0_outputs(6687)) or (layer0_outputs(751)));
    outputs(6605) <= not(layer0_outputs(7391)) or (layer0_outputs(1064));
    outputs(6606) <= not((layer0_outputs(2520)) or (layer0_outputs(4167)));
    outputs(6607) <= (layer0_outputs(1773)) and (layer0_outputs(2866));
    outputs(6608) <= not(layer0_outputs(5661)) or (layer0_outputs(2474));
    outputs(6609) <= not(layer0_outputs(1967)) or (layer0_outputs(4657));
    outputs(6610) <= not((layer0_outputs(179)) xor (layer0_outputs(5868)));
    outputs(6611) <= layer0_outputs(6116);
    outputs(6612) <= (layer0_outputs(6746)) or (layer0_outputs(5270));
    outputs(6613) <= not(layer0_outputs(632));
    outputs(6614) <= not(layer0_outputs(2602)) or (layer0_outputs(3400));
    outputs(6615) <= not(layer0_outputs(123));
    outputs(6616) <= layer0_outputs(4186);
    outputs(6617) <= not(layer0_outputs(5560)) or (layer0_outputs(1105));
    outputs(6618) <= layer0_outputs(7248);
    outputs(6619) <= layer0_outputs(5163);
    outputs(6620) <= not(layer0_outputs(6124));
    outputs(6621) <= not((layer0_outputs(2518)) xor (layer0_outputs(6790)));
    outputs(6622) <= not((layer0_outputs(7334)) or (layer0_outputs(7591)));
    outputs(6623) <= (layer0_outputs(1508)) and not (layer0_outputs(3027));
    outputs(6624) <= not((layer0_outputs(958)) or (layer0_outputs(5783)));
    outputs(6625) <= not(layer0_outputs(3186));
    outputs(6626) <= not((layer0_outputs(5269)) and (layer0_outputs(1194)));
    outputs(6627) <= (layer0_outputs(6757)) and (layer0_outputs(6979));
    outputs(6628) <= not((layer0_outputs(7540)) xor (layer0_outputs(3366)));
    outputs(6629) <= layer0_outputs(4643);
    outputs(6630) <= layer0_outputs(6794);
    outputs(6631) <= not((layer0_outputs(246)) xor (layer0_outputs(6643)));
    outputs(6632) <= not((layer0_outputs(3619)) and (layer0_outputs(250)));
    outputs(6633) <= layer0_outputs(6165);
    outputs(6634) <= layer0_outputs(5830);
    outputs(6635) <= (layer0_outputs(3929)) xor (layer0_outputs(372));
    outputs(6636) <= (layer0_outputs(5790)) or (layer0_outputs(6599));
    outputs(6637) <= not((layer0_outputs(4313)) xor (layer0_outputs(1743)));
    outputs(6638) <= not(layer0_outputs(6167)) or (layer0_outputs(5817));
    outputs(6639) <= not(layer0_outputs(3433));
    outputs(6640) <= (layer0_outputs(7420)) and not (layer0_outputs(4085));
    outputs(6641) <= (layer0_outputs(5929)) and not (layer0_outputs(7599));
    outputs(6642) <= not(layer0_outputs(4290)) or (layer0_outputs(5695));
    outputs(6643) <= not(layer0_outputs(3925)) or (layer0_outputs(1983));
    outputs(6644) <= layer0_outputs(4874);
    outputs(6645) <= not(layer0_outputs(4198));
    outputs(6646) <= not(layer0_outputs(1080)) or (layer0_outputs(1290));
    outputs(6647) <= not((layer0_outputs(3464)) xor (layer0_outputs(4204)));
    outputs(6648) <= (layer0_outputs(3906)) xor (layer0_outputs(7143));
    outputs(6649) <= not((layer0_outputs(4809)) and (layer0_outputs(6905)));
    outputs(6650) <= layer0_outputs(4654);
    outputs(6651) <= not((layer0_outputs(903)) and (layer0_outputs(4258)));
    outputs(6652) <= (layer0_outputs(1984)) xor (layer0_outputs(152));
    outputs(6653) <= layer0_outputs(2581);
    outputs(6654) <= not(layer0_outputs(352));
    outputs(6655) <= not(layer0_outputs(4504));
    outputs(6656) <= (layer0_outputs(3260)) and not (layer0_outputs(7487));
    outputs(6657) <= not((layer0_outputs(453)) xor (layer0_outputs(5910)));
    outputs(6658) <= not(layer0_outputs(2690));
    outputs(6659) <= layer0_outputs(5280);
    outputs(6660) <= (layer0_outputs(6374)) or (layer0_outputs(4490));
    outputs(6661) <= not((layer0_outputs(6404)) and (layer0_outputs(2101)));
    outputs(6662) <= not((layer0_outputs(4387)) xor (layer0_outputs(7546)));
    outputs(6663) <= not(layer0_outputs(5740)) or (layer0_outputs(890));
    outputs(6664) <= not(layer0_outputs(3671));
    outputs(6665) <= (layer0_outputs(2304)) or (layer0_outputs(7181));
    outputs(6666) <= layer0_outputs(5697);
    outputs(6667) <= layer0_outputs(1213);
    outputs(6668) <= layer0_outputs(2996);
    outputs(6669) <= layer0_outputs(1998);
    outputs(6670) <= (layer0_outputs(4298)) or (layer0_outputs(2393));
    outputs(6671) <= not(layer0_outputs(271)) or (layer0_outputs(6075));
    outputs(6672) <= not(layer0_outputs(7590)) or (layer0_outputs(2730));
    outputs(6673) <= not(layer0_outputs(7635)) or (layer0_outputs(5406));
    outputs(6674) <= (layer0_outputs(4344)) xor (layer0_outputs(5143));
    outputs(6675) <= not((layer0_outputs(4892)) xor (layer0_outputs(5272)));
    outputs(6676) <= not(layer0_outputs(1108));
    outputs(6677) <= not((layer0_outputs(7096)) xor (layer0_outputs(100)));
    outputs(6678) <= not(layer0_outputs(5146));
    outputs(6679) <= layer0_outputs(4094);
    outputs(6680) <= (layer0_outputs(3286)) and not (layer0_outputs(6715));
    outputs(6681) <= not((layer0_outputs(4170)) xor (layer0_outputs(7057)));
    outputs(6682) <= (layer0_outputs(5062)) and not (layer0_outputs(1143));
    outputs(6683) <= (layer0_outputs(518)) xor (layer0_outputs(7331));
    outputs(6684) <= not(layer0_outputs(1401));
    outputs(6685) <= layer0_outputs(4664);
    outputs(6686) <= not((layer0_outputs(5155)) xor (layer0_outputs(5161)));
    outputs(6687) <= (layer0_outputs(655)) xor (layer0_outputs(7673));
    outputs(6688) <= (layer0_outputs(38)) xor (layer0_outputs(166));
    outputs(6689) <= not((layer0_outputs(5385)) xor (layer0_outputs(3616)));
    outputs(6690) <= layer0_outputs(4245);
    outputs(6691) <= layer0_outputs(3920);
    outputs(6692) <= not(layer0_outputs(7351));
    outputs(6693) <= (layer0_outputs(720)) and not (layer0_outputs(6336));
    outputs(6694) <= not((layer0_outputs(7381)) xor (layer0_outputs(4001)));
    outputs(6695) <= not(layer0_outputs(3081));
    outputs(6696) <= not(layer0_outputs(450)) or (layer0_outputs(1072));
    outputs(6697) <= not((layer0_outputs(492)) xor (layer0_outputs(2798)));
    outputs(6698) <= not((layer0_outputs(3530)) and (layer0_outputs(3121)));
    outputs(6699) <= not(layer0_outputs(490));
    outputs(6700) <= (layer0_outputs(2196)) and (layer0_outputs(7505));
    outputs(6701) <= (layer0_outputs(3549)) or (layer0_outputs(7415));
    outputs(6702) <= (layer0_outputs(701)) xor (layer0_outputs(4370));
    outputs(6703) <= not(layer0_outputs(2305)) or (layer0_outputs(3438));
    outputs(6704) <= not((layer0_outputs(3671)) and (layer0_outputs(3429)));
    outputs(6705) <= not((layer0_outputs(6490)) or (layer0_outputs(6294)));
    outputs(6706) <= not(layer0_outputs(7584));
    outputs(6707) <= layer0_outputs(7424);
    outputs(6708) <= (layer0_outputs(7549)) and not (layer0_outputs(1672));
    outputs(6709) <= (layer0_outputs(5054)) xor (layer0_outputs(2367));
    outputs(6710) <= layer0_outputs(7272);
    outputs(6711) <= layer0_outputs(2042);
    outputs(6712) <= (layer0_outputs(3498)) xor (layer0_outputs(2529));
    outputs(6713) <= not((layer0_outputs(20)) and (layer0_outputs(781)));
    outputs(6714) <= layer0_outputs(6394);
    outputs(6715) <= (layer0_outputs(2927)) and not (layer0_outputs(7011));
    outputs(6716) <= not((layer0_outputs(9)) and (layer0_outputs(5628)));
    outputs(6717) <= layer0_outputs(5895);
    outputs(6718) <= (layer0_outputs(4219)) and not (layer0_outputs(4466));
    outputs(6719) <= not(layer0_outputs(1443)) or (layer0_outputs(4501));
    outputs(6720) <= not(layer0_outputs(742)) or (layer0_outputs(6527));
    outputs(6721) <= (layer0_outputs(4567)) xor (layer0_outputs(6875));
    outputs(6722) <= not(layer0_outputs(3160));
    outputs(6723) <= not(layer0_outputs(846));
    outputs(6724) <= not((layer0_outputs(2763)) or (layer0_outputs(2444)));
    outputs(6725) <= (layer0_outputs(4924)) and not (layer0_outputs(862));
    outputs(6726) <= layer0_outputs(548);
    outputs(6727) <= not(layer0_outputs(815)) or (layer0_outputs(2555));
    outputs(6728) <= not((layer0_outputs(1625)) xor (layer0_outputs(6604)));
    outputs(6729) <= layer0_outputs(2274);
    outputs(6730) <= (layer0_outputs(3515)) and not (layer0_outputs(2029));
    outputs(6731) <= (layer0_outputs(5395)) xor (layer0_outputs(6988));
    outputs(6732) <= (layer0_outputs(6828)) and not (layer0_outputs(7209));
    outputs(6733) <= not((layer0_outputs(7638)) or (layer0_outputs(7581)));
    outputs(6734) <= not((layer0_outputs(2331)) xor (layer0_outputs(5952)));
    outputs(6735) <= not(layer0_outputs(299));
    outputs(6736) <= (layer0_outputs(5488)) xor (layer0_outputs(6423));
    outputs(6737) <= not(layer0_outputs(3947)) or (layer0_outputs(7247));
    outputs(6738) <= not(layer0_outputs(3789));
    outputs(6739) <= (layer0_outputs(4053)) and (layer0_outputs(1154));
    outputs(6740) <= (layer0_outputs(1372)) and (layer0_outputs(4451));
    outputs(6741) <= not((layer0_outputs(2446)) xor (layer0_outputs(5932)));
    outputs(6742) <= (layer0_outputs(75)) or (layer0_outputs(1891));
    outputs(6743) <= (layer0_outputs(6867)) xor (layer0_outputs(1469));
    outputs(6744) <= not(layer0_outputs(1631));
    outputs(6745) <= (layer0_outputs(5187)) and (layer0_outputs(2736));
    outputs(6746) <= layer0_outputs(4511);
    outputs(6747) <= not((layer0_outputs(6323)) or (layer0_outputs(6705)));
    outputs(6748) <= not(layer0_outputs(2099));
    outputs(6749) <= (layer0_outputs(2084)) xor (layer0_outputs(1601));
    outputs(6750) <= not(layer0_outputs(2294));
    outputs(6751) <= not(layer0_outputs(2351));
    outputs(6752) <= layer0_outputs(1895);
    outputs(6753) <= (layer0_outputs(1274)) and not (layer0_outputs(4388));
    outputs(6754) <= not(layer0_outputs(5130));
    outputs(6755) <= not((layer0_outputs(7355)) xor (layer0_outputs(7495)));
    outputs(6756) <= not((layer0_outputs(7090)) xor (layer0_outputs(3841)));
    outputs(6757) <= (layer0_outputs(4968)) and (layer0_outputs(5127));
    outputs(6758) <= not((layer0_outputs(4846)) xor (layer0_outputs(4478)));
    outputs(6759) <= not(layer0_outputs(2429));
    outputs(6760) <= (layer0_outputs(6931)) or (layer0_outputs(6319));
    outputs(6761) <= not((layer0_outputs(5126)) xor (layer0_outputs(722)));
    outputs(6762) <= not((layer0_outputs(5820)) xor (layer0_outputs(2450)));
    outputs(6763) <= layer0_outputs(4154);
    outputs(6764) <= not((layer0_outputs(5760)) or (layer0_outputs(1502)));
    outputs(6765) <= layer0_outputs(3621);
    outputs(6766) <= not((layer0_outputs(2030)) or (layer0_outputs(3448)));
    outputs(6767) <= not((layer0_outputs(4120)) xor (layer0_outputs(5860)));
    outputs(6768) <= not(layer0_outputs(5794));
    outputs(6769) <= (layer0_outputs(1945)) and not (layer0_outputs(384));
    outputs(6770) <= not(layer0_outputs(2073)) or (layer0_outputs(7550));
    outputs(6771) <= (layer0_outputs(6650)) xor (layer0_outputs(2192));
    outputs(6772) <= (layer0_outputs(6986)) xor (layer0_outputs(5271));
    outputs(6773) <= (layer0_outputs(105)) or (layer0_outputs(1726));
    outputs(6774) <= (layer0_outputs(2810)) and not (layer0_outputs(828));
    outputs(6775) <= (layer0_outputs(2746)) xor (layer0_outputs(2135));
    outputs(6776) <= (layer0_outputs(2325)) and (layer0_outputs(5418));
    outputs(6777) <= (layer0_outputs(6230)) and (layer0_outputs(7677));
    outputs(6778) <= (layer0_outputs(5615)) xor (layer0_outputs(6803));
    outputs(6779) <= not(layer0_outputs(4410)) or (layer0_outputs(3683));
    outputs(6780) <= not(layer0_outputs(7432));
    outputs(6781) <= layer0_outputs(2189);
    outputs(6782) <= not(layer0_outputs(521));
    outputs(6783) <= not((layer0_outputs(6425)) or (layer0_outputs(2157)));
    outputs(6784) <= (layer0_outputs(2069)) xor (layer0_outputs(5054));
    outputs(6785) <= (layer0_outputs(4011)) and (layer0_outputs(7129));
    outputs(6786) <= layer0_outputs(5793);
    outputs(6787) <= not(layer0_outputs(4858));
    outputs(6788) <= layer0_outputs(7098);
    outputs(6789) <= '1';
    outputs(6790) <= layer0_outputs(4178);
    outputs(6791) <= (layer0_outputs(90)) or (layer0_outputs(3118));
    outputs(6792) <= layer0_outputs(2123);
    outputs(6793) <= layer0_outputs(1040);
    outputs(6794) <= (layer0_outputs(1198)) and (layer0_outputs(296));
    outputs(6795) <= not((layer0_outputs(4191)) xor (layer0_outputs(2494)));
    outputs(6796) <= not((layer0_outputs(253)) xor (layer0_outputs(3399)));
    outputs(6797) <= not(layer0_outputs(1794));
    outputs(6798) <= layer0_outputs(6340);
    outputs(6799) <= not((layer0_outputs(6427)) xor (layer0_outputs(7013)));
    outputs(6800) <= (layer0_outputs(2643)) xor (layer0_outputs(4065));
    outputs(6801) <= not((layer0_outputs(6796)) and (layer0_outputs(6591)));
    outputs(6802) <= not((layer0_outputs(256)) and (layer0_outputs(4842)));
    outputs(6803) <= not(layer0_outputs(3784));
    outputs(6804) <= not((layer0_outputs(5119)) xor (layer0_outputs(6039)));
    outputs(6805) <= layer0_outputs(5523);
    outputs(6806) <= layer0_outputs(2421);
    outputs(6807) <= not(layer0_outputs(6822));
    outputs(6808) <= (layer0_outputs(4093)) xor (layer0_outputs(1492));
    outputs(6809) <= (layer0_outputs(791)) xor (layer0_outputs(4328));
    outputs(6810) <= not(layer0_outputs(5396));
    outputs(6811) <= (layer0_outputs(6048)) and not (layer0_outputs(295));
    outputs(6812) <= layer0_outputs(1817);
    outputs(6813) <= (layer0_outputs(5744)) and not (layer0_outputs(189));
    outputs(6814) <= not((layer0_outputs(6118)) xor (layer0_outputs(1870)));
    outputs(6815) <= not((layer0_outputs(1928)) and (layer0_outputs(6471)));
    outputs(6816) <= (layer0_outputs(1475)) xor (layer0_outputs(4342));
    outputs(6817) <= not(layer0_outputs(5169));
    outputs(6818) <= not(layer0_outputs(2550));
    outputs(6819) <= (layer0_outputs(1039)) xor (layer0_outputs(1814));
    outputs(6820) <= layer0_outputs(1917);
    outputs(6821) <= (layer0_outputs(5492)) or (layer0_outputs(6510));
    outputs(6822) <= layer0_outputs(6728);
    outputs(6823) <= not((layer0_outputs(4025)) and (layer0_outputs(285)));
    outputs(6824) <= not(layer0_outputs(5853));
    outputs(6825) <= (layer0_outputs(795)) xor (layer0_outputs(6258));
    outputs(6826) <= not(layer0_outputs(7024));
    outputs(6827) <= (layer0_outputs(3923)) xor (layer0_outputs(1056));
    outputs(6828) <= (layer0_outputs(1753)) xor (layer0_outputs(5089));
    outputs(6829) <= not((layer0_outputs(3656)) xor (layer0_outputs(1081)));
    outputs(6830) <= not(layer0_outputs(7605));
    outputs(6831) <= layer0_outputs(292);
    outputs(6832) <= (layer0_outputs(5679)) and not (layer0_outputs(5125));
    outputs(6833) <= not((layer0_outputs(1644)) or (layer0_outputs(102)));
    outputs(6834) <= not((layer0_outputs(6501)) xor (layer0_outputs(3590)));
    outputs(6835) <= (layer0_outputs(7338)) xor (layer0_outputs(6637));
    outputs(6836) <= not(layer0_outputs(5798));
    outputs(6837) <= (layer0_outputs(1164)) xor (layer0_outputs(1864));
    outputs(6838) <= (layer0_outputs(159)) xor (layer0_outputs(4472));
    outputs(6839) <= layer0_outputs(5706);
    outputs(6840) <= layer0_outputs(2060);
    outputs(6841) <= not(layer0_outputs(433)) or (layer0_outputs(6304));
    outputs(6842) <= layer0_outputs(3265);
    outputs(6843) <= (layer0_outputs(1704)) or (layer0_outputs(7422));
    outputs(6844) <= layer0_outputs(6431);
    outputs(6845) <= not(layer0_outputs(6284));
    outputs(6846) <= not(layer0_outputs(5532));
    outputs(6847) <= layer0_outputs(6690);
    outputs(6848) <= (layer0_outputs(2787)) or (layer0_outputs(6939));
    outputs(6849) <= not((layer0_outputs(2721)) xor (layer0_outputs(1109)));
    outputs(6850) <= not((layer0_outputs(7060)) xor (layer0_outputs(7302)));
    outputs(6851) <= not(layer0_outputs(4515)) or (layer0_outputs(2164));
    outputs(6852) <= not((layer0_outputs(3698)) xor (layer0_outputs(920)));
    outputs(6853) <= not(layer0_outputs(4994));
    outputs(6854) <= not(layer0_outputs(1460)) or (layer0_outputs(3525));
    outputs(6855) <= (layer0_outputs(5611)) xor (layer0_outputs(4215));
    outputs(6856) <= (layer0_outputs(3085)) and not (layer0_outputs(4525));
    outputs(6857) <= not(layer0_outputs(6824));
    outputs(6858) <= (layer0_outputs(4008)) or (layer0_outputs(4556));
    outputs(6859) <= (layer0_outputs(122)) xor (layer0_outputs(5193));
    outputs(6860) <= not(layer0_outputs(3957));
    outputs(6861) <= not(layer0_outputs(2068));
    outputs(6862) <= (layer0_outputs(5875)) xor (layer0_outputs(7661));
    outputs(6863) <= not((layer0_outputs(3736)) and (layer0_outputs(6117)));
    outputs(6864) <= layer0_outputs(112);
    outputs(6865) <= not((layer0_outputs(1545)) xor (layer0_outputs(688)));
    outputs(6866) <= not(layer0_outputs(4759)) or (layer0_outputs(5790));
    outputs(6867) <= not(layer0_outputs(7537));
    outputs(6868) <= not((layer0_outputs(7370)) and (layer0_outputs(4868)));
    outputs(6869) <= not((layer0_outputs(3793)) xor (layer0_outputs(889)));
    outputs(6870) <= layer0_outputs(3615);
    outputs(6871) <= (layer0_outputs(6414)) xor (layer0_outputs(5797));
    outputs(6872) <= layer0_outputs(227);
    outputs(6873) <= (layer0_outputs(3347)) or (layer0_outputs(1731));
    outputs(6874) <= layer0_outputs(6724);
    outputs(6875) <= layer0_outputs(3148);
    outputs(6876) <= not(layer0_outputs(4423)) or (layer0_outputs(6924));
    outputs(6877) <= (layer0_outputs(5427)) xor (layer0_outputs(5421));
    outputs(6878) <= not(layer0_outputs(5702));
    outputs(6879) <= layer0_outputs(679);
    outputs(6880) <= layer0_outputs(511);
    outputs(6881) <= not(layer0_outputs(189));
    outputs(6882) <= (layer0_outputs(2870)) and (layer0_outputs(3367));
    outputs(6883) <= layer0_outputs(3678);
    outputs(6884) <= layer0_outputs(5483);
    outputs(6885) <= (layer0_outputs(7042)) xor (layer0_outputs(277));
    outputs(6886) <= not((layer0_outputs(1007)) xor (layer0_outputs(3686)));
    outputs(6887) <= (layer0_outputs(5)) and not (layer0_outputs(6683));
    outputs(6888) <= not((layer0_outputs(4950)) xor (layer0_outputs(1314)));
    outputs(6889) <= (layer0_outputs(3381)) or (layer0_outputs(5279));
    outputs(6890) <= not(layer0_outputs(4161)) or (layer0_outputs(1288));
    outputs(6891) <= not(layer0_outputs(6224));
    outputs(6892) <= not((layer0_outputs(26)) and (layer0_outputs(3203)));
    outputs(6893) <= not((layer0_outputs(1)) or (layer0_outputs(4460)));
    outputs(6894) <= (layer0_outputs(510)) and (layer0_outputs(1946));
    outputs(6895) <= not((layer0_outputs(4832)) xor (layer0_outputs(4116)));
    outputs(6896) <= layer0_outputs(3964);
    outputs(6897) <= not(layer0_outputs(1552));
    outputs(6898) <= (layer0_outputs(7421)) and (layer0_outputs(2989));
    outputs(6899) <= not((layer0_outputs(2267)) and (layer0_outputs(635)));
    outputs(6900) <= not((layer0_outputs(6982)) xor (layer0_outputs(1232)));
    outputs(6901) <= not(layer0_outputs(7122)) or (layer0_outputs(320));
    outputs(6902) <= not(layer0_outputs(4355)) or (layer0_outputs(481));
    outputs(6903) <= not((layer0_outputs(7286)) or (layer0_outputs(1310)));
    outputs(6904) <= not((layer0_outputs(1168)) xor (layer0_outputs(6125)));
    outputs(6905) <= (layer0_outputs(7153)) and not (layer0_outputs(2174));
    outputs(6906) <= (layer0_outputs(7640)) and not (layer0_outputs(1205));
    outputs(6907) <= not(layer0_outputs(7451)) or (layer0_outputs(1062));
    outputs(6908) <= not(layer0_outputs(769));
    outputs(6909) <= not(layer0_outputs(779));
    outputs(6910) <= (layer0_outputs(5851)) xor (layer0_outputs(3371));
    outputs(6911) <= not(layer0_outputs(3133)) or (layer0_outputs(1812));
    outputs(6912) <= (layer0_outputs(7618)) and not (layer0_outputs(4089));
    outputs(6913) <= (layer0_outputs(5788)) and not (layer0_outputs(6514));
    outputs(6914) <= not((layer0_outputs(7357)) xor (layer0_outputs(950)));
    outputs(6915) <= (layer0_outputs(2522)) and (layer0_outputs(6342));
    outputs(6916) <= layer0_outputs(3838);
    outputs(6917) <= (layer0_outputs(488)) xor (layer0_outputs(7413));
    outputs(6918) <= layer0_outputs(4433);
    outputs(6919) <= layer0_outputs(338);
    outputs(6920) <= (layer0_outputs(7189)) and not (layer0_outputs(2241));
    outputs(6921) <= not(layer0_outputs(2517));
    outputs(6922) <= (layer0_outputs(3353)) xor (layer0_outputs(5071));
    outputs(6923) <= layer0_outputs(4945);
    outputs(6924) <= layer0_outputs(6013);
    outputs(6925) <= not((layer0_outputs(2977)) or (layer0_outputs(4946)));
    outputs(6926) <= (layer0_outputs(4895)) and (layer0_outputs(7536));
    outputs(6927) <= not(layer0_outputs(3533));
    outputs(6928) <= (layer0_outputs(1394)) and not (layer0_outputs(3324));
    outputs(6929) <= layer0_outputs(2566);
    outputs(6930) <= (layer0_outputs(711)) xor (layer0_outputs(5416));
    outputs(6931) <= (layer0_outputs(6158)) and (layer0_outputs(1338));
    outputs(6932) <= (layer0_outputs(1182)) and not (layer0_outputs(4546));
    outputs(6933) <= not(layer0_outputs(5277));
    outputs(6934) <= not(layer0_outputs(4121));
    outputs(6935) <= not(layer0_outputs(2132));
    outputs(6936) <= (layer0_outputs(3669)) and not (layer0_outputs(7529));
    outputs(6937) <= not((layer0_outputs(5030)) or (layer0_outputs(2439)));
    outputs(6938) <= layer0_outputs(2657);
    outputs(6939) <= (layer0_outputs(3472)) and not (layer0_outputs(1824));
    outputs(6940) <= not(layer0_outputs(3570));
    outputs(6941) <= not(layer0_outputs(5491));
    outputs(6942) <= not((layer0_outputs(1782)) or (layer0_outputs(2470)));
    outputs(6943) <= (layer0_outputs(7158)) xor (layer0_outputs(1584));
    outputs(6944) <= layer0_outputs(1887);
    outputs(6945) <= (layer0_outputs(2667)) and not (layer0_outputs(5225));
    outputs(6946) <= layer0_outputs(2704);
    outputs(6947) <= layer0_outputs(7245);
    outputs(6948) <= not((layer0_outputs(3518)) and (layer0_outputs(2885)));
    outputs(6949) <= layer0_outputs(4728);
    outputs(6950) <= not((layer0_outputs(5278)) or (layer0_outputs(4585)));
    outputs(6951) <= not(layer0_outputs(5353));
    outputs(6952) <= layer0_outputs(5606);
    outputs(6953) <= not(layer0_outputs(575));
    outputs(6954) <= not(layer0_outputs(1572));
    outputs(6955) <= (layer0_outputs(7577)) and (layer0_outputs(969));
    outputs(6956) <= not((layer0_outputs(4774)) or (layer0_outputs(5783)));
    outputs(6957) <= not(layer0_outputs(1451));
    outputs(6958) <= layer0_outputs(5772);
    outputs(6959) <= (layer0_outputs(5023)) xor (layer0_outputs(5327));
    outputs(6960) <= (layer0_outputs(4956)) xor (layer0_outputs(2757));
    outputs(6961) <= (layer0_outputs(5616)) and not (layer0_outputs(7436));
    outputs(6962) <= not(layer0_outputs(5593));
    outputs(6963) <= (layer0_outputs(265)) and not (layer0_outputs(1136));
    outputs(6964) <= (layer0_outputs(868)) and (layer0_outputs(2695));
    outputs(6965) <= not((layer0_outputs(6272)) xor (layer0_outputs(6150)));
    outputs(6966) <= not(layer0_outputs(1861));
    outputs(6967) <= layer0_outputs(7484);
    outputs(6968) <= not(layer0_outputs(2789)) or (layer0_outputs(6836));
    outputs(6969) <= not(layer0_outputs(4498));
    outputs(6970) <= not(layer0_outputs(2054));
    outputs(6971) <= layer0_outputs(1955);
    outputs(6972) <= (layer0_outputs(6949)) and not (layer0_outputs(5921));
    outputs(6973) <= not(layer0_outputs(560));
    outputs(6974) <= not((layer0_outputs(2096)) and (layer0_outputs(4248)));
    outputs(6975) <= (layer0_outputs(6393)) and not (layer0_outputs(1254));
    outputs(6976) <= (layer0_outputs(2599)) or (layer0_outputs(466));
    outputs(6977) <= not(layer0_outputs(5987));
    outputs(6978) <= not(layer0_outputs(7085));
    outputs(6979) <= (layer0_outputs(712)) xor (layer0_outputs(680));
    outputs(6980) <= (layer0_outputs(4816)) and not (layer0_outputs(346));
    outputs(6981) <= not(layer0_outputs(3741));
    outputs(6982) <= not(layer0_outputs(2316));
    outputs(6983) <= layer0_outputs(270);
    outputs(6984) <= not(layer0_outputs(4543));
    outputs(6985) <= (layer0_outputs(2794)) xor (layer0_outputs(7452));
    outputs(6986) <= layer0_outputs(4896);
    outputs(6987) <= layer0_outputs(6973);
    outputs(6988) <= not((layer0_outputs(1697)) or (layer0_outputs(6915)));
    outputs(6989) <= (layer0_outputs(6665)) and (layer0_outputs(4114));
    outputs(6990) <= not((layer0_outputs(5104)) xor (layer0_outputs(7464)));
    outputs(6991) <= layer0_outputs(2076);
    outputs(6992) <= not((layer0_outputs(2374)) and (layer0_outputs(3635)));
    outputs(6993) <= (layer0_outputs(2545)) and not (layer0_outputs(5115));
    outputs(6994) <= not((layer0_outputs(2088)) or (layer0_outputs(1729)));
    outputs(6995) <= (layer0_outputs(2650)) xor (layer0_outputs(4509));
    outputs(6996) <= not(layer0_outputs(3492)) or (layer0_outputs(5617));
    outputs(6997) <= layer0_outputs(4307);
    outputs(6998) <= not(layer0_outputs(5140));
    outputs(6999) <= (layer0_outputs(1356)) xor (layer0_outputs(4798));
    outputs(7000) <= (layer0_outputs(4942)) xor (layer0_outputs(1627));
    outputs(7001) <= layer0_outputs(7540);
    outputs(7002) <= (layer0_outputs(4856)) xor (layer0_outputs(4412));
    outputs(7003) <= layer0_outputs(1879);
    outputs(7004) <= not(layer0_outputs(1454)) or (layer0_outputs(1823));
    outputs(7005) <= not(layer0_outputs(6725));
    outputs(7006) <= not((layer0_outputs(3049)) or (layer0_outputs(7115)));
    outputs(7007) <= layer0_outputs(3342);
    outputs(7008) <= not((layer0_outputs(1043)) xor (layer0_outputs(572)));
    outputs(7009) <= (layer0_outputs(5631)) xor (layer0_outputs(1060));
    outputs(7010) <= not((layer0_outputs(2681)) xor (layer0_outputs(4769)));
    outputs(7011) <= (layer0_outputs(1113)) xor (layer0_outputs(708));
    outputs(7012) <= (layer0_outputs(2745)) xor (layer0_outputs(5179));
    outputs(7013) <= not((layer0_outputs(7434)) or (layer0_outputs(1935)));
    outputs(7014) <= (layer0_outputs(797)) xor (layer0_outputs(5256));
    outputs(7015) <= not((layer0_outputs(6199)) xor (layer0_outputs(7438)));
    outputs(7016) <= not(layer0_outputs(1188));
    outputs(7017) <= (layer0_outputs(61)) and not (layer0_outputs(823));
    outputs(7018) <= not(layer0_outputs(4928));
    outputs(7019) <= not((layer0_outputs(1265)) or (layer0_outputs(7125)));
    outputs(7020) <= (layer0_outputs(2063)) xor (layer0_outputs(901));
    outputs(7021) <= layer0_outputs(1410);
    outputs(7022) <= (layer0_outputs(3767)) or (layer0_outputs(886));
    outputs(7023) <= (layer0_outputs(2850)) or (layer0_outputs(3298));
    outputs(7024) <= (layer0_outputs(1609)) and not (layer0_outputs(3700));
    outputs(7025) <= not((layer0_outputs(7421)) xor (layer0_outputs(812)));
    outputs(7026) <= (layer0_outputs(2660)) and (layer0_outputs(4843));
    outputs(7027) <= (layer0_outputs(6424)) and (layer0_outputs(3820));
    outputs(7028) <= (layer0_outputs(7229)) and (layer0_outputs(431));
    outputs(7029) <= not((layer0_outputs(3669)) xor (layer0_outputs(4262)));
    outputs(7030) <= (layer0_outputs(5544)) and not (layer0_outputs(5898));
    outputs(7031) <= layer0_outputs(7624);
    outputs(7032) <= (layer0_outputs(6579)) xor (layer0_outputs(5959));
    outputs(7033) <= (layer0_outputs(4560)) and not (layer0_outputs(244));
    outputs(7034) <= layer0_outputs(6246);
    outputs(7035) <= layer0_outputs(3991);
    outputs(7036) <= not(layer0_outputs(3695));
    outputs(7037) <= (layer0_outputs(6854)) or (layer0_outputs(7006));
    outputs(7038) <= not((layer0_outputs(6843)) xor (layer0_outputs(5890)));
    outputs(7039) <= (layer0_outputs(4877)) and not (layer0_outputs(3949));
    outputs(7040) <= (layer0_outputs(2106)) and (layer0_outputs(7618));
    outputs(7041) <= layer0_outputs(5555);
    outputs(7042) <= not(layer0_outputs(6741));
    outputs(7043) <= (layer0_outputs(3987)) and (layer0_outputs(4441));
    outputs(7044) <= not(layer0_outputs(5623)) or (layer0_outputs(5281));
    outputs(7045) <= (layer0_outputs(4667)) and not (layer0_outputs(5669));
    outputs(7046) <= (layer0_outputs(1263)) and not (layer0_outputs(728));
    outputs(7047) <= (layer0_outputs(4827)) and not (layer0_outputs(3525));
    outputs(7048) <= (layer0_outputs(5791)) and (layer0_outputs(7026));
    outputs(7049) <= not(layer0_outputs(7456));
    outputs(7050) <= (layer0_outputs(5036)) xor (layer0_outputs(2618));
    outputs(7051) <= not(layer0_outputs(2332));
    outputs(7052) <= (layer0_outputs(5366)) xor (layer0_outputs(698));
    outputs(7053) <= layer0_outputs(985);
    outputs(7054) <= layer0_outputs(3118);
    outputs(7055) <= layer0_outputs(6197);
    outputs(7056) <= not((layer0_outputs(4239)) or (layer0_outputs(5843)));
    outputs(7057) <= not(layer0_outputs(3293));
    outputs(7058) <= not((layer0_outputs(6879)) or (layer0_outputs(1091)));
    outputs(7059) <= (layer0_outputs(4704)) or (layer0_outputs(1315));
    outputs(7060) <= (layer0_outputs(3446)) xor (layer0_outputs(5340));
    outputs(7061) <= layer0_outputs(3456);
    outputs(7062) <= layer0_outputs(2499);
    outputs(7063) <= layer0_outputs(6395);
    outputs(7064) <= (layer0_outputs(3847)) and not (layer0_outputs(4182));
    outputs(7065) <= layer0_outputs(6710);
    outputs(7066) <= not((layer0_outputs(677)) or (layer0_outputs(4044)));
    outputs(7067) <= layer0_outputs(7064);
    outputs(7068) <= (layer0_outputs(6409)) xor (layer0_outputs(2282));
    outputs(7069) <= (layer0_outputs(4796)) and not (layer0_outputs(2490));
    outputs(7070) <= (layer0_outputs(1450)) and not (layer0_outputs(3227));
    outputs(7071) <= layer0_outputs(4912);
    outputs(7072) <= layer0_outputs(1802);
    outputs(7073) <= (layer0_outputs(4753)) and not (layer0_outputs(4359));
    outputs(7074) <= (layer0_outputs(3971)) and not (layer0_outputs(4023));
    outputs(7075) <= not(layer0_outputs(3030));
    outputs(7076) <= (layer0_outputs(2222)) xor (layer0_outputs(2898));
    outputs(7077) <= not(layer0_outputs(7269));
    outputs(7078) <= layer0_outputs(59);
    outputs(7079) <= (layer0_outputs(5780)) and not (layer0_outputs(305));
    outputs(7080) <= (layer0_outputs(1094)) xor (layer0_outputs(6422));
    outputs(7081) <= layer0_outputs(2061);
    outputs(7082) <= layer0_outputs(4742);
    outputs(7083) <= not((layer0_outputs(406)) xor (layer0_outputs(207)));
    outputs(7084) <= layer0_outputs(4610);
    outputs(7085) <= not(layer0_outputs(2109));
    outputs(7086) <= not((layer0_outputs(4865)) and (layer0_outputs(1187)));
    outputs(7087) <= layer0_outputs(3830);
    outputs(7088) <= not(layer0_outputs(5743));
    outputs(7089) <= not((layer0_outputs(4168)) and (layer0_outputs(397)));
    outputs(7090) <= (layer0_outputs(4802)) and not (layer0_outputs(3631));
    outputs(7091) <= not(layer0_outputs(6886));
    outputs(7092) <= not(layer0_outputs(1710));
    outputs(7093) <= (layer0_outputs(5301)) and not (layer0_outputs(2573));
    outputs(7094) <= layer0_outputs(4234);
    outputs(7095) <= layer0_outputs(998);
    outputs(7096) <= not(layer0_outputs(3613));
    outputs(7097) <= layer0_outputs(3229);
    outputs(7098) <= not((layer0_outputs(3311)) xor (layer0_outputs(2594)));
    outputs(7099) <= not(layer0_outputs(2702));
    outputs(7100) <= (layer0_outputs(456)) and not (layer0_outputs(4798));
    outputs(7101) <= not(layer0_outputs(6778));
    outputs(7102) <= layer0_outputs(1970);
    outputs(7103) <= (layer0_outputs(6223)) xor (layer0_outputs(2229));
    outputs(7104) <= (layer0_outputs(2852)) and not (layer0_outputs(1984));
    outputs(7105) <= not((layer0_outputs(3341)) and (layer0_outputs(4692)));
    outputs(7106) <= (layer0_outputs(6455)) and not (layer0_outputs(3604));
    outputs(7107) <= layer0_outputs(7484);
    outputs(7108) <= not((layer0_outputs(1725)) xor (layer0_outputs(4885)));
    outputs(7109) <= (layer0_outputs(2939)) and not (layer0_outputs(670));
    outputs(7110) <= (layer0_outputs(1618)) xor (layer0_outputs(598));
    outputs(7111) <= not(layer0_outputs(3963));
    outputs(7112) <= layer0_outputs(7023);
    outputs(7113) <= not((layer0_outputs(6597)) xor (layer0_outputs(4021)));
    outputs(7114) <= (layer0_outputs(6300)) and not (layer0_outputs(2093));
    outputs(7115) <= not((layer0_outputs(7407)) or (layer0_outputs(606)));
    outputs(7116) <= not(layer0_outputs(34)) or (layer0_outputs(1049));
    outputs(7117) <= layer0_outputs(3738);
    outputs(7118) <= not((layer0_outputs(498)) xor (layer0_outputs(6215)));
    outputs(7119) <= not(layer0_outputs(3567)) or (layer0_outputs(6279));
    outputs(7120) <= (layer0_outputs(3370)) and not (layer0_outputs(5088));
    outputs(7121) <= not((layer0_outputs(2685)) xor (layer0_outputs(5018)));
    outputs(7122) <= (layer0_outputs(7608)) and not (layer0_outputs(7675));
    outputs(7123) <= layer0_outputs(3993);
    outputs(7124) <= (layer0_outputs(6730)) and (layer0_outputs(5012));
    outputs(7125) <= layer0_outputs(2952);
    outputs(7126) <= not(layer0_outputs(5907));
    outputs(7127) <= (layer0_outputs(6388)) and not (layer0_outputs(6585));
    outputs(7128) <= not((layer0_outputs(4436)) or (layer0_outputs(3208)));
    outputs(7129) <= layer0_outputs(725);
    outputs(7130) <= not(layer0_outputs(5670));
    outputs(7131) <= layer0_outputs(6686);
    outputs(7132) <= (layer0_outputs(3091)) and (layer0_outputs(6212));
    outputs(7133) <= not(layer0_outputs(3130)) or (layer0_outputs(5656));
    outputs(7134) <= not(layer0_outputs(1014));
    outputs(7135) <= (layer0_outputs(50)) and not (layer0_outputs(574));
    outputs(7136) <= not(layer0_outputs(1472));
    outputs(7137) <= not(layer0_outputs(5538));
    outputs(7138) <= (layer0_outputs(1655)) and (layer0_outputs(2960));
    outputs(7139) <= (layer0_outputs(1070)) and (layer0_outputs(5321));
    outputs(7140) <= not(layer0_outputs(1341));
    outputs(7141) <= layer0_outputs(3633);
    outputs(7142) <= (layer0_outputs(6871)) and (layer0_outputs(1533));
    outputs(7143) <= layer0_outputs(5057);
    outputs(7144) <= not((layer0_outputs(353)) xor (layer0_outputs(4020)));
    outputs(7145) <= not(layer0_outputs(4623));
    outputs(7146) <= (layer0_outputs(2740)) xor (layer0_outputs(7377));
    outputs(7147) <= not((layer0_outputs(2390)) or (layer0_outputs(5739)));
    outputs(7148) <= (layer0_outputs(4520)) and (layer0_outputs(6706));
    outputs(7149) <= not(layer0_outputs(2293));
    outputs(7150) <= layer0_outputs(5377);
    outputs(7151) <= (layer0_outputs(3852)) and (layer0_outputs(192));
    outputs(7152) <= (layer0_outputs(495)) xor (layer0_outputs(2408));
    outputs(7153) <= layer0_outputs(5134);
    outputs(7154) <= layer0_outputs(183);
    outputs(7155) <= not(layer0_outputs(752)) or (layer0_outputs(7106));
    outputs(7156) <= (layer0_outputs(1858)) xor (layer0_outputs(4106));
    outputs(7157) <= layer0_outputs(3229);
    outputs(7158) <= (layer0_outputs(4156)) xor (layer0_outputs(5605));
    outputs(7159) <= not((layer0_outputs(2392)) or (layer0_outputs(3776)));
    outputs(7160) <= layer0_outputs(4031);
    outputs(7161) <= layer0_outputs(5434);
    outputs(7162) <= (layer0_outputs(6780)) and not (layer0_outputs(5581));
    outputs(7163) <= (layer0_outputs(4640)) and not (layer0_outputs(82));
    outputs(7164) <= not(layer0_outputs(6273));
    outputs(7165) <= (layer0_outputs(3281)) and (layer0_outputs(570));
    outputs(7166) <= (layer0_outputs(1832)) xor (layer0_outputs(1462));
    outputs(7167) <= (layer0_outputs(7061)) xor (layer0_outputs(1931));
    outputs(7168) <= not(layer0_outputs(5048));
    outputs(7169) <= not(layer0_outputs(7312));
    outputs(7170) <= (layer0_outputs(7146)) xor (layer0_outputs(4265));
    outputs(7171) <= not(layer0_outputs(7160)) or (layer0_outputs(4394));
    outputs(7172) <= not((layer0_outputs(5739)) xor (layer0_outputs(2544)));
    outputs(7173) <= not((layer0_outputs(5741)) xor (layer0_outputs(1175)));
    outputs(7174) <= not(layer0_outputs(3803));
    outputs(7175) <= layer0_outputs(2402);
    outputs(7176) <= (layer0_outputs(1549)) or (layer0_outputs(2897));
    outputs(7177) <= not((layer0_outputs(6865)) or (layer0_outputs(481)));
    outputs(7178) <= not((layer0_outputs(3005)) or (layer0_outputs(4776)));
    outputs(7179) <= not(layer0_outputs(5815)) or (layer0_outputs(7072));
    outputs(7180) <= (layer0_outputs(6557)) xor (layer0_outputs(2463));
    outputs(7181) <= not((layer0_outputs(3414)) or (layer0_outputs(6948)));
    outputs(7182) <= (layer0_outputs(88)) xor (layer0_outputs(5511));
    outputs(7183) <= not(layer0_outputs(3252));
    outputs(7184) <= layer0_outputs(967);
    outputs(7185) <= not(layer0_outputs(115));
    outputs(7186) <= not((layer0_outputs(3553)) and (layer0_outputs(4091)));
    outputs(7187) <= layer0_outputs(6956);
    outputs(7188) <= not(layer0_outputs(3266));
    outputs(7189) <= not(layer0_outputs(2900));
    outputs(7190) <= (layer0_outputs(5702)) and not (layer0_outputs(7));
    outputs(7191) <= not((layer0_outputs(2726)) or (layer0_outputs(1189)));
    outputs(7192) <= layer0_outputs(5983);
    outputs(7193) <= (layer0_outputs(3458)) and not (layer0_outputs(912));
    outputs(7194) <= layer0_outputs(1157);
    outputs(7195) <= not(layer0_outputs(1862));
    outputs(7196) <= (layer0_outputs(1370)) xor (layer0_outputs(1784));
    outputs(7197) <= layer0_outputs(1950);
    outputs(7198) <= (layer0_outputs(2366)) and not (layer0_outputs(3494));
    outputs(7199) <= layer0_outputs(3115);
    outputs(7200) <= (layer0_outputs(7559)) and not (layer0_outputs(5924));
    outputs(7201) <= (layer0_outputs(3501)) and not (layer0_outputs(5285));
    outputs(7202) <= not(layer0_outputs(1600));
    outputs(7203) <= layer0_outputs(1802);
    outputs(7204) <= (layer0_outputs(3003)) and not (layer0_outputs(6232));
    outputs(7205) <= layer0_outputs(4586);
    outputs(7206) <= not((layer0_outputs(6016)) xor (layer0_outputs(6504)));
    outputs(7207) <= layer0_outputs(2729);
    outputs(7208) <= not(layer0_outputs(6161));
    outputs(7209) <= (layer0_outputs(6554)) and not (layer0_outputs(3410));
    outputs(7210) <= not(layer0_outputs(4196));
    outputs(7211) <= not((layer0_outputs(347)) or (layer0_outputs(2475)));
    outputs(7212) <= layer0_outputs(331);
    outputs(7213) <= (layer0_outputs(1755)) and not (layer0_outputs(6303));
    outputs(7214) <= not((layer0_outputs(493)) or (layer0_outputs(5337)));
    outputs(7215) <= not(layer0_outputs(1212));
    outputs(7216) <= layer0_outputs(3255);
    outputs(7217) <= layer0_outputs(281);
    outputs(7218) <= (layer0_outputs(303)) and not (layer0_outputs(4765));
    outputs(7219) <= not(layer0_outputs(1054)) or (layer0_outputs(7537));
    outputs(7220) <= (layer0_outputs(3889)) or (layer0_outputs(2092));
    outputs(7221) <= (layer0_outputs(3607)) or (layer0_outputs(5682));
    outputs(7222) <= layer0_outputs(3886);
    outputs(7223) <= not(layer0_outputs(2142));
    outputs(7224) <= (layer0_outputs(4346)) and not (layer0_outputs(6168));
    outputs(7225) <= (layer0_outputs(210)) and (layer0_outputs(3624));
    outputs(7226) <= (layer0_outputs(4474)) and (layer0_outputs(2784));
    outputs(7227) <= (layer0_outputs(5896)) and (layer0_outputs(2151));
    outputs(7228) <= (layer0_outputs(6283)) and (layer0_outputs(4237));
    outputs(7229) <= not(layer0_outputs(5092));
    outputs(7230) <= not((layer0_outputs(4717)) and (layer0_outputs(2572)));
    outputs(7231) <= not(layer0_outputs(5736));
    outputs(7232) <= layer0_outputs(6788);
    outputs(7233) <= layer0_outputs(3013);
    outputs(7234) <= not((layer0_outputs(2793)) xor (layer0_outputs(201)));
    outputs(7235) <= (layer0_outputs(333)) and not (layer0_outputs(2951));
    outputs(7236) <= not((layer0_outputs(2102)) or (layer0_outputs(3400)));
    outputs(7237) <= not((layer0_outputs(1973)) or (layer0_outputs(5870)));
    outputs(7238) <= not((layer0_outputs(717)) xor (layer0_outputs(5769)));
    outputs(7239) <= layer0_outputs(7016);
    outputs(7240) <= (layer0_outputs(2440)) and (layer0_outputs(2456));
    outputs(7241) <= (layer0_outputs(2720)) and not (layer0_outputs(6734));
    outputs(7242) <= (layer0_outputs(6321)) and (layer0_outputs(3991));
    outputs(7243) <= (layer0_outputs(4348)) or (layer0_outputs(1362));
    outputs(7244) <= not(layer0_outputs(2047));
    outputs(7245) <= (layer0_outputs(753)) and not (layer0_outputs(6746));
    outputs(7246) <= (layer0_outputs(2440)) and not (layer0_outputs(7481));
    outputs(7247) <= not(layer0_outputs(3675)) or (layer0_outputs(1241));
    outputs(7248) <= (layer0_outputs(2760)) xor (layer0_outputs(5210));
    outputs(7249) <= (layer0_outputs(5452)) xor (layer0_outputs(5212));
    outputs(7250) <= layer0_outputs(6138);
    outputs(7251) <= layer0_outputs(4682);
    outputs(7252) <= (layer0_outputs(36)) and (layer0_outputs(4095));
    outputs(7253) <= (layer0_outputs(594)) and (layer0_outputs(2043));
    outputs(7254) <= layer0_outputs(3045);
    outputs(7255) <= (layer0_outputs(1000)) and not (layer0_outputs(631));
    outputs(7256) <= not(layer0_outputs(6678));
    outputs(7257) <= (layer0_outputs(343)) xor (layer0_outputs(7017));
    outputs(7258) <= (layer0_outputs(3670)) xor (layer0_outputs(2224));
    outputs(7259) <= not((layer0_outputs(6353)) xor (layer0_outputs(7099)));
    outputs(7260) <= not(layer0_outputs(6367));
    outputs(7261) <= not((layer0_outputs(2727)) or (layer0_outputs(4533)));
    outputs(7262) <= not(layer0_outputs(6880)) or (layer0_outputs(735));
    outputs(7263) <= not(layer0_outputs(1257));
    outputs(7264) <= layer0_outputs(5880);
    outputs(7265) <= (layer0_outputs(3319)) and not (layer0_outputs(71));
    outputs(7266) <= layer0_outputs(5677);
    outputs(7267) <= not(layer0_outputs(1589)) or (layer0_outputs(5828));
    outputs(7268) <= layer0_outputs(1930);
    outputs(7269) <= layer0_outputs(6556);
    outputs(7270) <= (layer0_outputs(5494)) or (layer0_outputs(6633));
    outputs(7271) <= not((layer0_outputs(4605)) or (layer0_outputs(3405)));
    outputs(7272) <= (layer0_outputs(2817)) xor (layer0_outputs(4210));
    outputs(7273) <= (layer0_outputs(3250)) and not (layer0_outputs(3982));
    outputs(7274) <= (layer0_outputs(4408)) and (layer0_outputs(5003));
    outputs(7275) <= not(layer0_outputs(1063));
    outputs(7276) <= layer0_outputs(3863);
    outputs(7277) <= (layer0_outputs(1574)) and not (layer0_outputs(4406));
    outputs(7278) <= layer0_outputs(4324);
    outputs(7279) <= not(layer0_outputs(992));
    outputs(7280) <= not(layer0_outputs(5055));
    outputs(7281) <= (layer0_outputs(4836)) xor (layer0_outputs(6076));
    outputs(7282) <= layer0_outputs(1205);
    outputs(7283) <= layer0_outputs(5859);
    outputs(7284) <= layer0_outputs(6026);
    outputs(7285) <= layer0_outputs(6246);
    outputs(7286) <= not((layer0_outputs(1366)) xor (layer0_outputs(7368)));
    outputs(7287) <= not(layer0_outputs(341));
    outputs(7288) <= layer0_outputs(6233);
    outputs(7289) <= not(layer0_outputs(482)) or (layer0_outputs(2375));
    outputs(7290) <= (layer0_outputs(6421)) and (layer0_outputs(3655));
    outputs(7291) <= layer0_outputs(3219);
    outputs(7292) <= not(layer0_outputs(2976));
    outputs(7293) <= not(layer0_outputs(5858)) or (layer0_outputs(5137));
    outputs(7294) <= (layer0_outputs(4464)) and not (layer0_outputs(2726));
    outputs(7295) <= (layer0_outputs(4480)) xor (layer0_outputs(7201));
    outputs(7296) <= layer0_outputs(298);
    outputs(7297) <= (layer0_outputs(3217)) and (layer0_outputs(7317));
    outputs(7298) <= (layer0_outputs(2870)) and not (layer0_outputs(2018));
    outputs(7299) <= (layer0_outputs(1878)) and not (layer0_outputs(2109));
    outputs(7300) <= not(layer0_outputs(3197));
    outputs(7301) <= (layer0_outputs(4696)) or (layer0_outputs(1659));
    outputs(7302) <= not(layer0_outputs(5694));
    outputs(7303) <= (layer0_outputs(1230)) xor (layer0_outputs(3303));
    outputs(7304) <= (layer0_outputs(2606)) xor (layer0_outputs(5305));
    outputs(7305) <= (layer0_outputs(3233)) and not (layer0_outputs(4985));
    outputs(7306) <= not((layer0_outputs(4386)) or (layer0_outputs(244)));
    outputs(7307) <= layer0_outputs(3392);
    outputs(7308) <= layer0_outputs(2327);
    outputs(7309) <= layer0_outputs(571);
    outputs(7310) <= layer0_outputs(1747);
    outputs(7311) <= not(layer0_outputs(530));
    outputs(7312) <= layer0_outputs(504);
    outputs(7313) <= not((layer0_outputs(7274)) or (layer0_outputs(5370)));
    outputs(7314) <= not(layer0_outputs(94));
    outputs(7315) <= (layer0_outputs(5423)) xor (layer0_outputs(852));
    outputs(7316) <= layer0_outputs(6125);
    outputs(7317) <= (layer0_outputs(3560)) and (layer0_outputs(1342));
    outputs(7318) <= layer0_outputs(6203);
    outputs(7319) <= layer0_outputs(1429);
    outputs(7320) <= (layer0_outputs(4213)) xor (layer0_outputs(5116));
    outputs(7321) <= (layer0_outputs(6941)) and not (layer0_outputs(5380));
    outputs(7322) <= (layer0_outputs(6292)) and not (layer0_outputs(5181));
    outputs(7323) <= (layer0_outputs(3279)) and not (layer0_outputs(3397));
    outputs(7324) <= (layer0_outputs(6172)) xor (layer0_outputs(5067));
    outputs(7325) <= (layer0_outputs(5870)) xor (layer0_outputs(1353));
    outputs(7326) <= not(layer0_outputs(7372));
    outputs(7327) <= (layer0_outputs(7326)) and (layer0_outputs(996));
    outputs(7328) <= (layer0_outputs(3273)) and not (layer0_outputs(3896));
    outputs(7329) <= (layer0_outputs(5534)) xor (layer0_outputs(5732));
    outputs(7330) <= not(layer0_outputs(929));
    outputs(7331) <= (layer0_outputs(2695)) and not (layer0_outputs(1682));
    outputs(7332) <= not((layer0_outputs(2066)) or (layer0_outputs(4979)));
    outputs(7333) <= (layer0_outputs(6115)) or (layer0_outputs(125));
    outputs(7334) <= (layer0_outputs(1933)) and (layer0_outputs(684));
    outputs(7335) <= (layer0_outputs(7291)) and not (layer0_outputs(3540));
    outputs(7336) <= (layer0_outputs(3277)) and (layer0_outputs(3180));
    outputs(7337) <= (layer0_outputs(7544)) and (layer0_outputs(5551));
    outputs(7338) <= not(layer0_outputs(1258));
    outputs(7339) <= not(layer0_outputs(4108)) or (layer0_outputs(5542));
    outputs(7340) <= not((layer0_outputs(2233)) xor (layer0_outputs(581)));
    outputs(7341) <= (layer0_outputs(3765)) or (layer0_outputs(4193));
    outputs(7342) <= (layer0_outputs(6169)) and not (layer0_outputs(4322));
    outputs(7343) <= layer0_outputs(451);
    outputs(7344) <= (layer0_outputs(1828)) and not (layer0_outputs(6719));
    outputs(7345) <= not(layer0_outputs(2455));
    outputs(7346) <= (layer0_outputs(7176)) xor (layer0_outputs(1088));
    outputs(7347) <= (layer0_outputs(7587)) xor (layer0_outputs(2191));
    outputs(7348) <= layer0_outputs(5848);
    outputs(7349) <= not(layer0_outputs(5154));
    outputs(7350) <= not(layer0_outputs(4286));
    outputs(7351) <= layer0_outputs(6457);
    outputs(7352) <= not((layer0_outputs(156)) and (layer0_outputs(6595)));
    outputs(7353) <= not((layer0_outputs(1377)) xor (layer0_outputs(6242)));
    outputs(7354) <= not((layer0_outputs(5966)) xor (layer0_outputs(6310)));
    outputs(7355) <= not(layer0_outputs(5239));
    outputs(7356) <= (layer0_outputs(716)) and (layer0_outputs(1714));
    outputs(7357) <= (layer0_outputs(7406)) and not (layer0_outputs(3186));
    outputs(7358) <= not((layer0_outputs(3056)) or (layer0_outputs(1064)));
    outputs(7359) <= not((layer0_outputs(2413)) and (layer0_outputs(83)));
    outputs(7360) <= (layer0_outputs(4137)) and not (layer0_outputs(6313));
    outputs(7361) <= (layer0_outputs(157)) xor (layer0_outputs(3383));
    outputs(7362) <= not((layer0_outputs(6816)) or (layer0_outputs(1642)));
    outputs(7363) <= layer0_outputs(1321);
    outputs(7364) <= (layer0_outputs(4160)) and not (layer0_outputs(4212));
    outputs(7365) <= not((layer0_outputs(4756)) xor (layer0_outputs(5235)));
    outputs(7366) <= layer0_outputs(4573);
    outputs(7367) <= (layer0_outputs(7595)) and not (layer0_outputs(2856));
    outputs(7368) <= not(layer0_outputs(2161));
    outputs(7369) <= layer0_outputs(1991);
    outputs(7370) <= (layer0_outputs(4391)) xor (layer0_outputs(1118));
    outputs(7371) <= (layer0_outputs(4795)) xor (layer0_outputs(6435));
    outputs(7372) <= not((layer0_outputs(7073)) or (layer0_outputs(4109)));
    outputs(7373) <= not((layer0_outputs(3123)) xor (layer0_outputs(3764)));
    outputs(7374) <= (layer0_outputs(6536)) and not (layer0_outputs(2438));
    outputs(7375) <= (layer0_outputs(5446)) and not (layer0_outputs(4118));
    outputs(7376) <= (layer0_outputs(6809)) and not (layer0_outputs(4963));
    outputs(7377) <= not(layer0_outputs(1122)) or (layer0_outputs(925));
    outputs(7378) <= (layer0_outputs(4534)) and not (layer0_outputs(418));
    outputs(7379) <= not((layer0_outputs(7015)) or (layer0_outputs(1884)));
    outputs(7380) <= layer0_outputs(190);
    outputs(7381) <= not(layer0_outputs(5232)) or (layer0_outputs(27));
    outputs(7382) <= not(layer0_outputs(786));
    outputs(7383) <= not((layer0_outputs(6853)) or (layer0_outputs(2358)));
    outputs(7384) <= not(layer0_outputs(5574));
    outputs(7385) <= (layer0_outputs(5021)) xor (layer0_outputs(555));
    outputs(7386) <= layer0_outputs(6524);
    outputs(7387) <= (layer0_outputs(5962)) and (layer0_outputs(3100));
    outputs(7388) <= not((layer0_outputs(7261)) or (layer0_outputs(5954)));
    outputs(7389) <= layer0_outputs(600);
    outputs(7390) <= not(layer0_outputs(396));
    outputs(7391) <= not(layer0_outputs(6887));
    outputs(7392) <= not(layer0_outputs(3967));
    outputs(7393) <= not(layer0_outputs(3344));
    outputs(7394) <= layer0_outputs(7330);
    outputs(7395) <= not((layer0_outputs(6967)) or (layer0_outputs(4108)));
    outputs(7396) <= (layer0_outputs(69)) and (layer0_outputs(90));
    outputs(7397) <= not(layer0_outputs(1028));
    outputs(7398) <= not((layer0_outputs(3742)) or (layer0_outputs(1958)));
    outputs(7399) <= (layer0_outputs(4421)) and not (layer0_outputs(4494));
    outputs(7400) <= (layer0_outputs(6653)) or (layer0_outputs(5325));
    outputs(7401) <= not((layer0_outputs(6113)) and (layer0_outputs(4273)));
    outputs(7402) <= (layer0_outputs(5873)) or (layer0_outputs(4417));
    outputs(7403) <= not((layer0_outputs(7438)) or (layer0_outputs(2239)));
    outputs(7404) <= not(layer0_outputs(5711));
    outputs(7405) <= not(layer0_outputs(1912)) or (layer0_outputs(5362));
    outputs(7406) <= layer0_outputs(2352);
    outputs(7407) <= not((layer0_outputs(3877)) or (layer0_outputs(278)));
    outputs(7408) <= (layer0_outputs(3829)) and not (layer0_outputs(4143));
    outputs(7409) <= layer0_outputs(2430);
    outputs(7410) <= (layer0_outputs(1757)) xor (layer0_outputs(4375));
    outputs(7411) <= (layer0_outputs(479)) or (layer0_outputs(2394));
    outputs(7412) <= not(layer0_outputs(6947)) or (layer0_outputs(2286));
    outputs(7413) <= not((layer0_outputs(6019)) xor (layer0_outputs(6120)));
    outputs(7414) <= '0';
    outputs(7415) <= not(layer0_outputs(1580));
    outputs(7416) <= not(layer0_outputs(5366)) or (layer0_outputs(2041));
    outputs(7417) <= not((layer0_outputs(4255)) or (layer0_outputs(6622)));
    outputs(7418) <= not(layer0_outputs(356)) or (layer0_outputs(5942));
    outputs(7419) <= (layer0_outputs(3261)) xor (layer0_outputs(1577));
    outputs(7420) <= not((layer0_outputs(3455)) or (layer0_outputs(5583)));
    outputs(7421) <= (layer0_outputs(7086)) and not (layer0_outputs(2404));
    outputs(7422) <= (layer0_outputs(5816)) and not (layer0_outputs(1027));
    outputs(7423) <= layer0_outputs(4040);
    outputs(7424) <= not(layer0_outputs(5115));
    outputs(7425) <= not((layer0_outputs(6875)) or (layer0_outputs(2813)));
    outputs(7426) <= not((layer0_outputs(3773)) xor (layer0_outputs(7645)));
    outputs(7427) <= not((layer0_outputs(1147)) xor (layer0_outputs(444)));
    outputs(7428) <= (layer0_outputs(2167)) and not (layer0_outputs(4936));
    outputs(7429) <= layer0_outputs(6951);
    outputs(7430) <= (layer0_outputs(5307)) and not (layer0_outputs(2821));
    outputs(7431) <= layer0_outputs(5377);
    outputs(7432) <= layer0_outputs(5807);
    outputs(7433) <= not(layer0_outputs(6742));
    outputs(7434) <= (layer0_outputs(5592)) and not (layer0_outputs(2910));
    outputs(7435) <= layer0_outputs(7119);
    outputs(7436) <= layer0_outputs(5351);
    outputs(7437) <= not((layer0_outputs(3210)) xor (layer0_outputs(4400)));
    outputs(7438) <= (layer0_outputs(7412)) and not (layer0_outputs(1624));
    outputs(7439) <= not(layer0_outputs(5414));
    outputs(7440) <= layer0_outputs(5052);
    outputs(7441) <= not((layer0_outputs(3598)) xor (layer0_outputs(4768)));
    outputs(7442) <= not(layer0_outputs(2200));
    outputs(7443) <= not(layer0_outputs(786));
    outputs(7444) <= not(layer0_outputs(3928));
    outputs(7445) <= not((layer0_outputs(5411)) and (layer0_outputs(5251)));
    outputs(7446) <= (layer0_outputs(7599)) xor (layer0_outputs(4668));
    outputs(7447) <= not((layer0_outputs(2442)) xor (layer0_outputs(3111)));
    outputs(7448) <= layer0_outputs(3244);
    outputs(7449) <= (layer0_outputs(5283)) and (layer0_outputs(6144));
    outputs(7450) <= not(layer0_outputs(4934));
    outputs(7451) <= (layer0_outputs(3591)) xor (layer0_outputs(6572));
    outputs(7452) <= layer0_outputs(409);
    outputs(7453) <= (layer0_outputs(2546)) xor (layer0_outputs(5324));
    outputs(7454) <= not(layer0_outputs(6606));
    outputs(7455) <= not(layer0_outputs(1063)) or (layer0_outputs(5114));
    outputs(7456) <= (layer0_outputs(7404)) or (layer0_outputs(1402));
    outputs(7457) <= not(layer0_outputs(2113));
    outputs(7458) <= layer0_outputs(1481);
    outputs(7459) <= not(layer0_outputs(860));
    outputs(7460) <= (layer0_outputs(2043)) xor (layer0_outputs(3435));
    outputs(7461) <= (layer0_outputs(7290)) and not (layer0_outputs(4501));
    outputs(7462) <= layer0_outputs(3884);
    outputs(7463) <= (layer0_outputs(5429)) xor (layer0_outputs(3439));
    outputs(7464) <= layer0_outputs(821);
    outputs(7465) <= layer0_outputs(4797);
    outputs(7466) <= (layer0_outputs(1656)) and not (layer0_outputs(6318));
    outputs(7467) <= (layer0_outputs(6587)) and (layer0_outputs(6779));
    outputs(7468) <= not((layer0_outputs(285)) xor (layer0_outputs(7374)));
    outputs(7469) <= (layer0_outputs(7150)) and (layer0_outputs(4453));
    outputs(7470) <= (layer0_outputs(5641)) and not (layer0_outputs(3618));
    outputs(7471) <= not((layer0_outputs(4192)) and (layer0_outputs(2964)));
    outputs(7472) <= layer0_outputs(1000);
    outputs(7473) <= not(layer0_outputs(3819)) or (layer0_outputs(1727));
    outputs(7474) <= layer0_outputs(2300);
    outputs(7475) <= layer0_outputs(3337);
    outputs(7476) <= (layer0_outputs(2819)) or (layer0_outputs(6520));
    outputs(7477) <= not(layer0_outputs(1409));
    outputs(7478) <= not(layer0_outputs(6366)) or (layer0_outputs(5936));
    outputs(7479) <= not(layer0_outputs(5562));
    outputs(7480) <= not(layer0_outputs(3658));
    outputs(7481) <= not((layer0_outputs(5913)) or (layer0_outputs(3812)));
    outputs(7482) <= not((layer0_outputs(6316)) xor (layer0_outputs(4041)));
    outputs(7483) <= (layer0_outputs(27)) xor (layer0_outputs(3340));
    outputs(7484) <= not(layer0_outputs(2884));
    outputs(7485) <= not(layer0_outputs(2171));
    outputs(7486) <= not(layer0_outputs(4246));
    outputs(7487) <= layer0_outputs(1701);
    outputs(7488) <= not(layer0_outputs(7101));
    outputs(7489) <= not(layer0_outputs(4148));
    outputs(7490) <= (layer0_outputs(3507)) and not (layer0_outputs(5530));
    outputs(7491) <= (layer0_outputs(4271)) xor (layer0_outputs(204));
    outputs(7492) <= not(layer0_outputs(3072));
    outputs(7493) <= not((layer0_outputs(1416)) or (layer0_outputs(3061)));
    outputs(7494) <= (layer0_outputs(3488)) and not (layer0_outputs(762));
    outputs(7495) <= (layer0_outputs(888)) and (layer0_outputs(2570));
    outputs(7496) <= not(layer0_outputs(1355));
    outputs(7497) <= not(layer0_outputs(543));
    outputs(7498) <= layer0_outputs(6770);
    outputs(7499) <= (layer0_outputs(3247)) and not (layer0_outputs(4056));
    outputs(7500) <= layer0_outputs(961);
    outputs(7501) <= (layer0_outputs(4479)) and (layer0_outputs(1617));
    outputs(7502) <= (layer0_outputs(6597)) xor (layer0_outputs(3289));
    outputs(7503) <= layer0_outputs(1125);
    outputs(7504) <= layer0_outputs(3958);
    outputs(7505) <= (layer0_outputs(7489)) and (layer0_outputs(3668));
    outputs(7506) <= layer0_outputs(1275);
    outputs(7507) <= layer0_outputs(893);
    outputs(7508) <= not(layer0_outputs(1952));
    outputs(7509) <= not(layer0_outputs(2552)) or (layer0_outputs(2833));
    outputs(7510) <= layer0_outputs(1982);
    outputs(7511) <= not(layer0_outputs(6047));
    outputs(7512) <= layer0_outputs(1125);
    outputs(7513) <= not((layer0_outputs(4703)) or (layer0_outputs(5467)));
    outputs(7514) <= layer0_outputs(3490);
    outputs(7515) <= (layer0_outputs(7313)) and not (layer0_outputs(6263));
    outputs(7516) <= not((layer0_outputs(1024)) xor (layer0_outputs(4850)));
    outputs(7517) <= not((layer0_outputs(1504)) xor (layer0_outputs(4960)));
    outputs(7518) <= (layer0_outputs(5477)) and not (layer0_outputs(5946));
    outputs(7519) <= layer0_outputs(2061);
    outputs(7520) <= not((layer0_outputs(7309)) or (layer0_outputs(1658)));
    outputs(7521) <= not(layer0_outputs(537));
    outputs(7522) <= (layer0_outputs(2456)) xor (layer0_outputs(3792));
    outputs(7523) <= not(layer0_outputs(913));
    outputs(7524) <= (layer0_outputs(7660)) and not (layer0_outputs(1968));
    outputs(7525) <= not((layer0_outputs(5500)) or (layer0_outputs(4772)));
    outputs(7526) <= not(layer0_outputs(3460));
    outputs(7527) <= not(layer0_outputs(467));
    outputs(7528) <= layer0_outputs(837);
    outputs(7529) <= not(layer0_outputs(7345));
    outputs(7530) <= layer0_outputs(1521);
    outputs(7531) <= not((layer0_outputs(3786)) or (layer0_outputs(2251)));
    outputs(7532) <= not(layer0_outputs(7235));
    outputs(7533) <= not(layer0_outputs(1903));
    outputs(7534) <= not((layer0_outputs(3969)) or (layer0_outputs(6656)));
    outputs(7535) <= layer0_outputs(539);
    outputs(7536) <= (layer0_outputs(760)) or (layer0_outputs(6199));
    outputs(7537) <= not(layer0_outputs(2179));
    outputs(7538) <= (layer0_outputs(7624)) and (layer0_outputs(3541));
    outputs(7539) <= not(layer0_outputs(2014));
    outputs(7540) <= (layer0_outputs(6959)) xor (layer0_outputs(3647));
    outputs(7541) <= (layer0_outputs(2904)) and (layer0_outputs(7147));
    outputs(7542) <= (layer0_outputs(5329)) xor (layer0_outputs(6996));
    outputs(7543) <= layer0_outputs(3196);
    outputs(7544) <= (layer0_outputs(1032)) and not (layer0_outputs(4532));
    outputs(7545) <= not(layer0_outputs(4075));
    outputs(7546) <= not((layer0_outputs(1194)) xor (layer0_outputs(7249)));
    outputs(7547) <= not(layer0_outputs(3570));
    outputs(7548) <= not((layer0_outputs(4190)) and (layer0_outputs(6441)));
    outputs(7549) <= layer0_outputs(2263);
    outputs(7550) <= layer0_outputs(1437);
    outputs(7551) <= layer0_outputs(2610);
    outputs(7552) <= (layer0_outputs(1839)) xor (layer0_outputs(3411));
    outputs(7553) <= not((layer0_outputs(2823)) or (layer0_outputs(4987)));
    outputs(7554) <= layer0_outputs(3640);
    outputs(7555) <= not(layer0_outputs(7215));
    outputs(7556) <= not(layer0_outputs(3007));
    outputs(7557) <= layer0_outputs(5123);
    outputs(7558) <= (layer0_outputs(2319)) and not (layer0_outputs(1209));
    outputs(7559) <= (layer0_outputs(7141)) xor (layer0_outputs(6225));
    outputs(7560) <= not((layer0_outputs(5970)) xor (layer0_outputs(3624)));
    outputs(7561) <= not((layer0_outputs(956)) and (layer0_outputs(3363)));
    outputs(7562) <= (layer0_outputs(7220)) and not (layer0_outputs(7529));
    outputs(7563) <= (layer0_outputs(3128)) and not (layer0_outputs(6596));
    outputs(7564) <= (layer0_outputs(2785)) and not (layer0_outputs(6701));
    outputs(7565) <= not((layer0_outputs(6740)) or (layer0_outputs(5885)));
    outputs(7566) <= (layer0_outputs(1686)) and not (layer0_outputs(2330));
    outputs(7567) <= layer0_outputs(5791);
    outputs(7568) <= (layer0_outputs(3941)) and (layer0_outputs(7341));
    outputs(7569) <= layer0_outputs(3481);
    outputs(7570) <= not((layer0_outputs(847)) and (layer0_outputs(4878)));
    outputs(7571) <= not((layer0_outputs(5898)) or (layer0_outputs(2332)));
    outputs(7572) <= (layer0_outputs(789)) xor (layer0_outputs(4572));
    outputs(7573) <= layer0_outputs(6121);
    outputs(7574) <= not(layer0_outputs(4623));
    outputs(7575) <= (layer0_outputs(7027)) and not (layer0_outputs(301));
    outputs(7576) <= not(layer0_outputs(2562));
    outputs(7577) <= layer0_outputs(3824);
    outputs(7578) <= layer0_outputs(7116);
    outputs(7579) <= (layer0_outputs(231)) and not (layer0_outputs(3248));
    outputs(7580) <= layer0_outputs(4000);
    outputs(7581) <= (layer0_outputs(1423)) or (layer0_outputs(6417));
    outputs(7582) <= not(layer0_outputs(493));
    outputs(7583) <= not(layer0_outputs(516));
    outputs(7584) <= not(layer0_outputs(4839));
    outputs(7585) <= (layer0_outputs(2112)) and not (layer0_outputs(3724));
    outputs(7586) <= not((layer0_outputs(3469)) xor (layer0_outputs(7147)));
    outputs(7587) <= not((layer0_outputs(3807)) xor (layer0_outputs(6051)));
    outputs(7588) <= (layer0_outputs(1876)) and not (layer0_outputs(1546));
    outputs(7589) <= layer0_outputs(5318);
    outputs(7590) <= not(layer0_outputs(1412));
    outputs(7591) <= not(layer0_outputs(691));
    outputs(7592) <= (layer0_outputs(957)) and not (layer0_outputs(7616));
    outputs(7593) <= not((layer0_outputs(4523)) or (layer0_outputs(2777)));
    outputs(7594) <= layer0_outputs(2981);
    outputs(7595) <= layer0_outputs(7227);
    outputs(7596) <= not(layer0_outputs(6751));
    outputs(7597) <= not(layer0_outputs(2859)) or (layer0_outputs(6594));
    outputs(7598) <= not(layer0_outputs(7632)) or (layer0_outputs(4129));
    outputs(7599) <= layer0_outputs(3348);
    outputs(7600) <= (layer0_outputs(3230)) or (layer0_outputs(7530));
    outputs(7601) <= (layer0_outputs(5968)) and not (layer0_outputs(6734));
    outputs(7602) <= not(layer0_outputs(6886));
    outputs(7603) <= not(layer0_outputs(2689));
    outputs(7604) <= not(layer0_outputs(4577));
    outputs(7605) <= (layer0_outputs(7144)) and not (layer0_outputs(3664));
    outputs(7606) <= (layer0_outputs(3922)) and not (layer0_outputs(7233));
    outputs(7607) <= not((layer0_outputs(2823)) and (layer0_outputs(4081)));
    outputs(7608) <= not(layer0_outputs(1713));
    outputs(7609) <= not((layer0_outputs(6769)) or (layer0_outputs(6915)));
    outputs(7610) <= not(layer0_outputs(6760));
    outputs(7611) <= not(layer0_outputs(3479));
    outputs(7612) <= layer0_outputs(4538);
    outputs(7613) <= (layer0_outputs(4086)) and (layer0_outputs(896));
    outputs(7614) <= not((layer0_outputs(3486)) or (layer0_outputs(2956)));
    outputs(7615) <= not(layer0_outputs(1087));
    outputs(7616) <= layer0_outputs(4602);
    outputs(7617) <= not((layer0_outputs(5031)) xor (layer0_outputs(6820)));
    outputs(7618) <= layer0_outputs(5426);
    outputs(7619) <= (layer0_outputs(4517)) xor (layer0_outputs(2159));
    outputs(7620) <= not((layer0_outputs(2993)) or (layer0_outputs(4941)));
    outputs(7621) <= layer0_outputs(4120);
    outputs(7622) <= layer0_outputs(4895);
    outputs(7623) <= layer0_outputs(5664);
    outputs(7624) <= layer0_outputs(6188);
    outputs(7625) <= not((layer0_outputs(2712)) xor (layer0_outputs(7382)));
    outputs(7626) <= (layer0_outputs(2932)) and (layer0_outputs(6953));
    outputs(7627) <= layer0_outputs(2969);
    outputs(7628) <= not((layer0_outputs(1187)) or (layer0_outputs(1772)));
    outputs(7629) <= not((layer0_outputs(4662)) xor (layer0_outputs(4001)));
    outputs(7630) <= not((layer0_outputs(6243)) xor (layer0_outputs(6474)));
    outputs(7631) <= not(layer0_outputs(2739));
    outputs(7632) <= (layer0_outputs(2421)) and (layer0_outputs(3420));
    outputs(7633) <= not(layer0_outputs(5846)) or (layer0_outputs(4441));
    outputs(7634) <= (layer0_outputs(594)) and not (layer0_outputs(823));
    outputs(7635) <= not(layer0_outputs(2750)) or (layer0_outputs(3105));
    outputs(7636) <= (layer0_outputs(708)) xor (layer0_outputs(5953));
    outputs(7637) <= not(layer0_outputs(2603));
    outputs(7638) <= not(layer0_outputs(4158));
    outputs(7639) <= not((layer0_outputs(1156)) or (layer0_outputs(1793)));
    outputs(7640) <= not((layer0_outputs(4278)) xor (layer0_outputs(1408)));
    outputs(7641) <= (layer0_outputs(5937)) and not (layer0_outputs(4989));
    outputs(7642) <= not(layer0_outputs(2534));
    outputs(7643) <= not((layer0_outputs(1011)) xor (layer0_outputs(5100)));
    outputs(7644) <= not(layer0_outputs(1388));
    outputs(7645) <= not(layer0_outputs(764)) or (layer0_outputs(500));
    outputs(7646) <= not(layer0_outputs(518));
    outputs(7647) <= (layer0_outputs(6942)) and not (layer0_outputs(3261));
    outputs(7648) <= not((layer0_outputs(2559)) or (layer0_outputs(4624)));
    outputs(7649) <= not((layer0_outputs(6890)) or (layer0_outputs(513)));
    outputs(7650) <= (layer0_outputs(2545)) and not (layer0_outputs(1166));
    outputs(7651) <= (layer0_outputs(7058)) and (layer0_outputs(3593));
    outputs(7652) <= (layer0_outputs(3711)) xor (layer0_outputs(4383));
    outputs(7653) <= not(layer0_outputs(220));
    outputs(7654) <= (layer0_outputs(4792)) and not (layer0_outputs(941));
    outputs(7655) <= (layer0_outputs(321)) and not (layer0_outputs(6679));
    outputs(7656) <= not((layer0_outputs(3563)) and (layer0_outputs(3103)));
    outputs(7657) <= (layer0_outputs(2298)) and (layer0_outputs(1844));
    outputs(7658) <= not(layer0_outputs(7325)) or (layer0_outputs(4249));
    outputs(7659) <= not((layer0_outputs(4115)) or (layer0_outputs(5487)));
    outputs(7660) <= not((layer0_outputs(3641)) or (layer0_outputs(4749)));
    outputs(7661) <= (layer0_outputs(648)) and (layer0_outputs(4848));
    outputs(7662) <= not((layer0_outputs(4659)) xor (layer0_outputs(5838)));
    outputs(7663) <= not((layer0_outputs(7638)) or (layer0_outputs(6359)));
    outputs(7664) <= not(layer0_outputs(1907));
    outputs(7665) <= layer0_outputs(772);
    outputs(7666) <= not((layer0_outputs(7654)) xor (layer0_outputs(2030)));
    outputs(7667) <= (layer0_outputs(3145)) and not (layer0_outputs(4246));
    outputs(7668) <= not(layer0_outputs(5699));
    outputs(7669) <= (layer0_outputs(4849)) and not (layer0_outputs(2361));
    outputs(7670) <= not(layer0_outputs(2561));
    outputs(7671) <= (layer0_outputs(39)) and (layer0_outputs(1828));
    outputs(7672) <= (layer0_outputs(980)) xor (layer0_outputs(923));
    outputs(7673) <= not((layer0_outputs(3594)) or (layer0_outputs(6071)));
    outputs(7674) <= not((layer0_outputs(76)) and (layer0_outputs(5996)));
    outputs(7675) <= not((layer0_outputs(2571)) or (layer0_outputs(445)));
    outputs(7676) <= layer0_outputs(5192);
    outputs(7677) <= not((layer0_outputs(5182)) xor (layer0_outputs(4452)));
    outputs(7678) <= (layer0_outputs(3335)) or (layer0_outputs(6804));
    outputs(7679) <= layer0_outputs(3571);

end Behavioral;
