library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs : in std_logic_vector(255 downto 0);
        outputs : out std_logic_vector(2559 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs : std_logic_vector(2559 downto 0);

begin

    layer0_outputs(0) <= inputs(89);
    layer0_outputs(1) <= not(inputs(240));
    layer0_outputs(2) <= (inputs(61)) or (inputs(98));
    layer0_outputs(3) <= not((inputs(59)) or (inputs(94)));
    layer0_outputs(4) <= '0';
    layer0_outputs(5) <= not(inputs(105));
    layer0_outputs(6) <= (inputs(165)) or (inputs(109));
    layer0_outputs(7) <= (inputs(231)) and not (inputs(147));
    layer0_outputs(8) <= (inputs(141)) or (inputs(137));
    layer0_outputs(9) <= not(inputs(244));
    layer0_outputs(10) <= not((inputs(87)) or (inputs(12)));
    layer0_outputs(11) <= not(inputs(147));
    layer0_outputs(12) <= (inputs(237)) or (inputs(124));
    layer0_outputs(13) <= not(inputs(40));
    layer0_outputs(14) <= not(inputs(44)) or (inputs(231));
    layer0_outputs(15) <= not((inputs(98)) or (inputs(97)));
    layer0_outputs(16) <= not(inputs(83));
    layer0_outputs(17) <= (inputs(131)) and not (inputs(55));
    layer0_outputs(18) <= not(inputs(125));
    layer0_outputs(19) <= not(inputs(209));
    layer0_outputs(20) <= not((inputs(36)) or (inputs(10)));
    layer0_outputs(21) <= not((inputs(211)) or (inputs(130)));
    layer0_outputs(22) <= not(inputs(163));
    layer0_outputs(23) <= not((inputs(55)) and (inputs(96)));
    layer0_outputs(24) <= not(inputs(100));
    layer0_outputs(25) <= not(inputs(26));
    layer0_outputs(26) <= inputs(129);
    layer0_outputs(27) <= inputs(131);
    layer0_outputs(28) <= (inputs(20)) and not (inputs(161));
    layer0_outputs(29) <= not(inputs(50));
    layer0_outputs(30) <= not(inputs(191));
    layer0_outputs(31) <= not((inputs(185)) or (inputs(157)));
    layer0_outputs(32) <= (inputs(150)) or (inputs(159));
    layer0_outputs(33) <= inputs(188);
    layer0_outputs(34) <= (inputs(87)) and not (inputs(14));
    layer0_outputs(35) <= inputs(20);
    layer0_outputs(36) <= (inputs(114)) and not (inputs(47));
    layer0_outputs(37) <= not((inputs(251)) or (inputs(141)));
    layer0_outputs(38) <= not(inputs(218));
    layer0_outputs(39) <= not((inputs(204)) xor (inputs(252)));
    layer0_outputs(40) <= (inputs(49)) or (inputs(126));
    layer0_outputs(41) <= not(inputs(183));
    layer0_outputs(42) <= not(inputs(161)) or (inputs(158));
    layer0_outputs(43) <= inputs(101);
    layer0_outputs(44) <= not(inputs(86));
    layer0_outputs(45) <= inputs(10);
    layer0_outputs(46) <= not(inputs(100)) or (inputs(209));
    layer0_outputs(47) <= (inputs(250)) and not (inputs(144));
    layer0_outputs(48) <= not(inputs(61)) or (inputs(221));
    layer0_outputs(49) <= not((inputs(140)) or (inputs(98)));
    layer0_outputs(50) <= (inputs(239)) or (inputs(145));
    layer0_outputs(51) <= inputs(9);
    layer0_outputs(52) <= (inputs(252)) xor (inputs(153));
    layer0_outputs(53) <= (inputs(160)) or (inputs(210));
    layer0_outputs(54) <= not(inputs(119));
    layer0_outputs(55) <= inputs(135);
    layer0_outputs(56) <= inputs(100);
    layer0_outputs(57) <= (inputs(48)) and not (inputs(28));
    layer0_outputs(58) <= (inputs(68)) or (inputs(127));
    layer0_outputs(59) <= not(inputs(230)) or (inputs(106));
    layer0_outputs(60) <= inputs(137);
    layer0_outputs(61) <= inputs(179);
    layer0_outputs(62) <= not(inputs(21));
    layer0_outputs(63) <= not(inputs(21));
    layer0_outputs(64) <= (inputs(43)) and not (inputs(218));
    layer0_outputs(65) <= (inputs(143)) xor (inputs(130));
    layer0_outputs(66) <= not((inputs(241)) xor (inputs(150)));
    layer0_outputs(67) <= not(inputs(189));
    layer0_outputs(68) <= inputs(163);
    layer0_outputs(69) <= inputs(105);
    layer0_outputs(70) <= (inputs(22)) and not (inputs(114));
    layer0_outputs(71) <= not((inputs(27)) or (inputs(11)));
    layer0_outputs(72) <= not(inputs(152));
    layer0_outputs(73) <= not((inputs(92)) or (inputs(64)));
    layer0_outputs(74) <= inputs(146);
    layer0_outputs(75) <= inputs(217);
    layer0_outputs(76) <= not((inputs(149)) or (inputs(35)));
    layer0_outputs(77) <= not(inputs(204));
    layer0_outputs(78) <= not((inputs(232)) or (inputs(227)));
    layer0_outputs(79) <= (inputs(134)) or (inputs(135));
    layer0_outputs(80) <= not((inputs(137)) and (inputs(150)));
    layer0_outputs(81) <= (inputs(255)) or (inputs(70));
    layer0_outputs(82) <= inputs(181);
    layer0_outputs(83) <= not((inputs(196)) or (inputs(161)));
    layer0_outputs(84) <= (inputs(37)) and not (inputs(188));
    layer0_outputs(85) <= '1';
    layer0_outputs(86) <= not(inputs(249)) or (inputs(242));
    layer0_outputs(87) <= (inputs(61)) or (inputs(185));
    layer0_outputs(88) <= (inputs(191)) or (inputs(187));
    layer0_outputs(89) <= inputs(182);
    layer0_outputs(90) <= (inputs(244)) and not (inputs(81));
    layer0_outputs(91) <= not(inputs(87));
    layer0_outputs(92) <= (inputs(209)) xor (inputs(205));
    layer0_outputs(93) <= not(inputs(8)) or (inputs(2));
    layer0_outputs(94) <= (inputs(44)) or (inputs(73));
    layer0_outputs(95) <= '1';
    layer0_outputs(96) <= not(inputs(86));
    layer0_outputs(97) <= not((inputs(75)) xor (inputs(112)));
    layer0_outputs(98) <= not(inputs(211));
    layer0_outputs(99) <= '1';
    layer0_outputs(100) <= inputs(126);
    layer0_outputs(101) <= inputs(68);
    layer0_outputs(102) <= not(inputs(229));
    layer0_outputs(103) <= inputs(22);
    layer0_outputs(104) <= (inputs(22)) and (inputs(254));
    layer0_outputs(105) <= not(inputs(104));
    layer0_outputs(106) <= (inputs(72)) or (inputs(16));
    layer0_outputs(107) <= not(inputs(108));
    layer0_outputs(108) <= not(inputs(98)) or (inputs(79));
    layer0_outputs(109) <= not(inputs(199));
    layer0_outputs(110) <= (inputs(115)) and not (inputs(94));
    layer0_outputs(111) <= not(inputs(179));
    layer0_outputs(112) <= not(inputs(58)) or (inputs(174));
    layer0_outputs(113) <= not(inputs(27));
    layer0_outputs(114) <= not((inputs(117)) or (inputs(226)));
    layer0_outputs(115) <= (inputs(178)) and not (inputs(168));
    layer0_outputs(116) <= inputs(210);
    layer0_outputs(117) <= inputs(194);
    layer0_outputs(118) <= not(inputs(172));
    layer0_outputs(119) <= not(inputs(118));
    layer0_outputs(120) <= not(inputs(216));
    layer0_outputs(121) <= not(inputs(180));
    layer0_outputs(122) <= inputs(165);
    layer0_outputs(123) <= (inputs(180)) or (inputs(250));
    layer0_outputs(124) <= not((inputs(119)) or (inputs(102)));
    layer0_outputs(125) <= inputs(139);
    layer0_outputs(126) <= not(inputs(25));
    layer0_outputs(127) <= not((inputs(179)) or (inputs(78)));
    layer0_outputs(128) <= not((inputs(16)) or (inputs(91)));
    layer0_outputs(129) <= not(inputs(248)) or (inputs(223));
    layer0_outputs(130) <= (inputs(148)) or (inputs(68));
    layer0_outputs(131) <= not(inputs(94));
    layer0_outputs(132) <= inputs(97);
    layer0_outputs(133) <= not((inputs(192)) or (inputs(24)));
    layer0_outputs(134) <= not(inputs(48));
    layer0_outputs(135) <= not(inputs(180));
    layer0_outputs(136) <= inputs(108);
    layer0_outputs(137) <= not(inputs(220));
    layer0_outputs(138) <= inputs(226);
    layer0_outputs(139) <= not(inputs(105)) or (inputs(179));
    layer0_outputs(140) <= (inputs(99)) xor (inputs(208));
    layer0_outputs(141) <= '1';
    layer0_outputs(142) <= not(inputs(154)) or (inputs(10));
    layer0_outputs(143) <= not(inputs(197));
    layer0_outputs(144) <= (inputs(165)) and not (inputs(67));
    layer0_outputs(145) <= not(inputs(60));
    layer0_outputs(146) <= (inputs(19)) or (inputs(44));
    layer0_outputs(147) <= not(inputs(188)) or (inputs(155));
    layer0_outputs(148) <= not(inputs(237)) or (inputs(49));
    layer0_outputs(149) <= not((inputs(79)) or (inputs(5)));
    layer0_outputs(150) <= not((inputs(105)) or (inputs(239)));
    layer0_outputs(151) <= not(inputs(40));
    layer0_outputs(152) <= (inputs(157)) or (inputs(112));
    layer0_outputs(153) <= (inputs(237)) or (inputs(132));
    layer0_outputs(154) <= inputs(246);
    layer0_outputs(155) <= not(inputs(228)) or (inputs(46));
    layer0_outputs(156) <= not((inputs(210)) or (inputs(215)));
    layer0_outputs(157) <= inputs(231);
    layer0_outputs(158) <= not((inputs(23)) and (inputs(53)));
    layer0_outputs(159) <= not((inputs(171)) or (inputs(194)));
    layer0_outputs(160) <= not((inputs(84)) or (inputs(113)));
    layer0_outputs(161) <= not(inputs(149));
    layer0_outputs(162) <= not(inputs(88)) or (inputs(192));
    layer0_outputs(163) <= inputs(151);
    layer0_outputs(164) <= not(inputs(99));
    layer0_outputs(165) <= not(inputs(123)) or (inputs(3));
    layer0_outputs(166) <= not((inputs(72)) and (inputs(201)));
    layer0_outputs(167) <= not(inputs(29));
    layer0_outputs(168) <= inputs(61);
    layer0_outputs(169) <= not((inputs(178)) or (inputs(254)));
    layer0_outputs(170) <= inputs(151);
    layer0_outputs(171) <= not((inputs(25)) or (inputs(101)));
    layer0_outputs(172) <= (inputs(86)) or (inputs(15));
    layer0_outputs(173) <= (inputs(163)) or (inputs(147));
    layer0_outputs(174) <= inputs(59);
    layer0_outputs(175) <= '0';
    layer0_outputs(176) <= not(inputs(234)) or (inputs(5));
    layer0_outputs(177) <= not((inputs(180)) or (inputs(146)));
    layer0_outputs(178) <= (inputs(56)) or (inputs(243));
    layer0_outputs(179) <= inputs(11);
    layer0_outputs(180) <= not(inputs(178)) or (inputs(79));
    layer0_outputs(181) <= inputs(30);
    layer0_outputs(182) <= inputs(245);
    layer0_outputs(183) <= not(inputs(94));
    layer0_outputs(184) <= not(inputs(116));
    layer0_outputs(185) <= not(inputs(218));
    layer0_outputs(186) <= (inputs(1)) or (inputs(205));
    layer0_outputs(187) <= not(inputs(251));
    layer0_outputs(188) <= inputs(117);
    layer0_outputs(189) <= not((inputs(43)) or (inputs(49)));
    layer0_outputs(190) <= inputs(151);
    layer0_outputs(191) <= not((inputs(237)) xor (inputs(222)));
    layer0_outputs(192) <= inputs(140);
    layer0_outputs(193) <= not((inputs(247)) or (inputs(71)));
    layer0_outputs(194) <= not((inputs(191)) or (inputs(150)));
    layer0_outputs(195) <= inputs(117);
    layer0_outputs(196) <= inputs(214);
    layer0_outputs(197) <= (inputs(71)) or (inputs(156));
    layer0_outputs(198) <= not((inputs(3)) or (inputs(62)));
    layer0_outputs(199) <= not(inputs(23)) or (inputs(235));
    layer0_outputs(200) <= not((inputs(159)) or (inputs(252)));
    layer0_outputs(201) <= not(inputs(215)) or (inputs(145));
    layer0_outputs(202) <= (inputs(201)) or (inputs(174));
    layer0_outputs(203) <= (inputs(250)) and not (inputs(127));
    layer0_outputs(204) <= not((inputs(106)) or (inputs(253)));
    layer0_outputs(205) <= (inputs(6)) and not (inputs(221));
    layer0_outputs(206) <= not((inputs(115)) or (inputs(191)));
    layer0_outputs(207) <= not(inputs(39)) or (inputs(161));
    layer0_outputs(208) <= (inputs(231)) or (inputs(179));
    layer0_outputs(209) <= (inputs(204)) xor (inputs(255));
    layer0_outputs(210) <= not(inputs(185));
    layer0_outputs(211) <= not(inputs(119)) or (inputs(205));
    layer0_outputs(212) <= (inputs(98)) or (inputs(11));
    layer0_outputs(213) <= not((inputs(210)) or (inputs(243)));
    layer0_outputs(214) <= not((inputs(72)) and (inputs(5)));
    layer0_outputs(215) <= not((inputs(237)) or (inputs(202)));
    layer0_outputs(216) <= not((inputs(220)) or (inputs(36)));
    layer0_outputs(217) <= inputs(249);
    layer0_outputs(218) <= not(inputs(188));
    layer0_outputs(219) <= (inputs(9)) or (inputs(33));
    layer0_outputs(220) <= not((inputs(48)) or (inputs(172)));
    layer0_outputs(221) <= inputs(60);
    layer0_outputs(222) <= not((inputs(192)) or (inputs(7)));
    layer0_outputs(223) <= not(inputs(182));
    layer0_outputs(224) <= not(inputs(156));
    layer0_outputs(225) <= (inputs(105)) or (inputs(108));
    layer0_outputs(226) <= not(inputs(162));
    layer0_outputs(227) <= not((inputs(20)) or (inputs(56)));
    layer0_outputs(228) <= not(inputs(74)) or (inputs(207));
    layer0_outputs(229) <= not((inputs(120)) or (inputs(116)));
    layer0_outputs(230) <= not(inputs(140));
    layer0_outputs(231) <= inputs(20);
    layer0_outputs(232) <= not((inputs(239)) xor (inputs(173)));
    layer0_outputs(233) <= (inputs(41)) and not (inputs(117));
    layer0_outputs(234) <= (inputs(7)) or (inputs(76));
    layer0_outputs(235) <= (inputs(68)) and not (inputs(211));
    layer0_outputs(236) <= not(inputs(164)) or (inputs(129));
    layer0_outputs(237) <= inputs(75);
    layer0_outputs(238) <= inputs(10);
    layer0_outputs(239) <= not((inputs(227)) or (inputs(229)));
    layer0_outputs(240) <= '0';
    layer0_outputs(241) <= not((inputs(213)) xor (inputs(183)));
    layer0_outputs(242) <= inputs(122);
    layer0_outputs(243) <= inputs(83);
    layer0_outputs(244) <= inputs(5);
    layer0_outputs(245) <= not(inputs(207));
    layer0_outputs(246) <= not((inputs(255)) or (inputs(76)));
    layer0_outputs(247) <= (inputs(229)) or (inputs(209));
    layer0_outputs(248) <= (inputs(172)) xor (inputs(240));
    layer0_outputs(249) <= (inputs(89)) and not (inputs(49));
    layer0_outputs(250) <= inputs(58);
    layer0_outputs(251) <= not(inputs(121));
    layer0_outputs(252) <= (inputs(252)) or (inputs(168));
    layer0_outputs(253) <= not((inputs(47)) or (inputs(122)));
    layer0_outputs(254) <= (inputs(11)) or (inputs(80));
    layer0_outputs(255) <= not(inputs(173)) or (inputs(147));
    layer0_outputs(256) <= not(inputs(104));
    layer0_outputs(257) <= not(inputs(131));
    layer0_outputs(258) <= (inputs(22)) and not (inputs(146));
    layer0_outputs(259) <= not((inputs(166)) or (inputs(140)));
    layer0_outputs(260) <= inputs(181);
    layer0_outputs(261) <= (inputs(83)) or (inputs(80));
    layer0_outputs(262) <= not(inputs(89));
    layer0_outputs(263) <= not(inputs(103)) or (inputs(155));
    layer0_outputs(264) <= not((inputs(240)) xor (inputs(111)));
    layer0_outputs(265) <= not(inputs(110));
    layer0_outputs(266) <= not((inputs(236)) and (inputs(184)));
    layer0_outputs(267) <= (inputs(226)) or (inputs(176));
    layer0_outputs(268) <= not(inputs(97));
    layer0_outputs(269) <= not((inputs(218)) or (inputs(188)));
    layer0_outputs(270) <= not(inputs(228)) or (inputs(128));
    layer0_outputs(271) <= (inputs(97)) xor (inputs(70));
    layer0_outputs(272) <= (inputs(206)) or (inputs(30));
    layer0_outputs(273) <= inputs(22);
    layer0_outputs(274) <= not(inputs(46));
    layer0_outputs(275) <= not((inputs(65)) or (inputs(224)));
    layer0_outputs(276) <= (inputs(85)) and (inputs(40));
    layer0_outputs(277) <= (inputs(3)) or (inputs(156));
    layer0_outputs(278) <= (inputs(168)) and not (inputs(20));
    layer0_outputs(279) <= (inputs(252)) or (inputs(198));
    layer0_outputs(280) <= inputs(77);
    layer0_outputs(281) <= not((inputs(190)) or (inputs(164)));
    layer0_outputs(282) <= not(inputs(61));
    layer0_outputs(283) <= '0';
    layer0_outputs(284) <= inputs(84);
    layer0_outputs(285) <= not(inputs(33));
    layer0_outputs(286) <= inputs(228);
    layer0_outputs(287) <= not((inputs(80)) or (inputs(112)));
    layer0_outputs(288) <= (inputs(142)) or (inputs(146));
    layer0_outputs(289) <= not((inputs(33)) xor (inputs(78)));
    layer0_outputs(290) <= (inputs(26)) or (inputs(37));
    layer0_outputs(291) <= inputs(40);
    layer0_outputs(292) <= not(inputs(244));
    layer0_outputs(293) <= inputs(77);
    layer0_outputs(294) <= not(inputs(224));
    layer0_outputs(295) <= not(inputs(78)) or (inputs(166));
    layer0_outputs(296) <= (inputs(95)) or (inputs(179));
    layer0_outputs(297) <= not((inputs(43)) or (inputs(209)));
    layer0_outputs(298) <= (inputs(26)) and not (inputs(175));
    layer0_outputs(299) <= (inputs(173)) or (inputs(163));
    layer0_outputs(300) <= (inputs(128)) and (inputs(128));
    layer0_outputs(301) <= inputs(40);
    layer0_outputs(302) <= not(inputs(85)) or (inputs(254));
    layer0_outputs(303) <= not(inputs(50));
    layer0_outputs(304) <= not((inputs(0)) xor (inputs(22)));
    layer0_outputs(305) <= (inputs(193)) or (inputs(178));
    layer0_outputs(306) <= not(inputs(220));
    layer0_outputs(307) <= (inputs(122)) and not (inputs(203));
    layer0_outputs(308) <= not(inputs(150));
    layer0_outputs(309) <= not((inputs(97)) or (inputs(17)));
    layer0_outputs(310) <= not((inputs(223)) or (inputs(72)));
    layer0_outputs(311) <= inputs(151);
    layer0_outputs(312) <= inputs(20);
    layer0_outputs(313) <= not(inputs(169));
    layer0_outputs(314) <= not((inputs(253)) or (inputs(85)));
    layer0_outputs(315) <= not(inputs(169));
    layer0_outputs(316) <= (inputs(238)) or (inputs(79));
    layer0_outputs(317) <= inputs(46);
    layer0_outputs(318) <= inputs(44);
    layer0_outputs(319) <= (inputs(187)) or (inputs(67));
    layer0_outputs(320) <= not(inputs(10));
    layer0_outputs(321) <= inputs(246);
    layer0_outputs(322) <= (inputs(33)) xor (inputs(111));
    layer0_outputs(323) <= not(inputs(250));
    layer0_outputs(324) <= not(inputs(171));
    layer0_outputs(325) <= inputs(206);
    layer0_outputs(326) <= inputs(125);
    layer0_outputs(327) <= not((inputs(73)) and (inputs(35)));
    layer0_outputs(328) <= (inputs(229)) or (inputs(219));
    layer0_outputs(329) <= inputs(83);
    layer0_outputs(330) <= (inputs(154)) and not (inputs(76));
    layer0_outputs(331) <= (inputs(245)) or (inputs(204));
    layer0_outputs(332) <= not(inputs(84));
    layer0_outputs(333) <= inputs(75);
    layer0_outputs(334) <= not(inputs(133));
    layer0_outputs(335) <= (inputs(184)) or (inputs(66));
    layer0_outputs(336) <= inputs(110);
    layer0_outputs(337) <= not(inputs(214));
    layer0_outputs(338) <= (inputs(138)) and not (inputs(188));
    layer0_outputs(339) <= not(inputs(122));
    layer0_outputs(340) <= not(inputs(24)) or (inputs(191));
    layer0_outputs(341) <= (inputs(159)) xor (inputs(118));
    layer0_outputs(342) <= not((inputs(4)) or (inputs(82)));
    layer0_outputs(343) <= (inputs(181)) or (inputs(177));
    layer0_outputs(344) <= (inputs(117)) and not (inputs(180));
    layer0_outputs(345) <= inputs(220);
    layer0_outputs(346) <= inputs(246);
    layer0_outputs(347) <= (inputs(136)) or (inputs(191));
    layer0_outputs(348) <= inputs(85);
    layer0_outputs(349) <= not(inputs(70));
    layer0_outputs(350) <= (inputs(166)) and not (inputs(123));
    layer0_outputs(351) <= (inputs(191)) xor (inputs(237));
    layer0_outputs(352) <= (inputs(33)) or (inputs(179));
    layer0_outputs(353) <= inputs(74);
    layer0_outputs(354) <= (inputs(148)) and not (inputs(32));
    layer0_outputs(355) <= not((inputs(179)) xor (inputs(144)));
    layer0_outputs(356) <= (inputs(237)) and not (inputs(48));
    layer0_outputs(357) <= (inputs(199)) and not (inputs(16));
    layer0_outputs(358) <= (inputs(218)) or (inputs(158));
    layer0_outputs(359) <= not(inputs(233));
    layer0_outputs(360) <= inputs(180);
    layer0_outputs(361) <= not((inputs(35)) and (inputs(30)));
    layer0_outputs(362) <= not(inputs(230));
    layer0_outputs(363) <= not(inputs(106)) or (inputs(222));
    layer0_outputs(364) <= inputs(165);
    layer0_outputs(365) <= (inputs(140)) or (inputs(246));
    layer0_outputs(366) <= inputs(132);
    layer0_outputs(367) <= (inputs(237)) or (inputs(102));
    layer0_outputs(368) <= inputs(192);
    layer0_outputs(369) <= (inputs(53)) or (inputs(155));
    layer0_outputs(370) <= not((inputs(75)) or (inputs(143)));
    layer0_outputs(371) <= not(inputs(167)) or (inputs(133));
    layer0_outputs(372) <= not(inputs(102));
    layer0_outputs(373) <= (inputs(52)) or (inputs(96));
    layer0_outputs(374) <= (inputs(87)) and not (inputs(159));
    layer0_outputs(375) <= (inputs(89)) and not (inputs(158));
    layer0_outputs(376) <= not((inputs(117)) or (inputs(162)));
    layer0_outputs(377) <= inputs(217);
    layer0_outputs(378) <= '0';
    layer0_outputs(379) <= not(inputs(54));
    layer0_outputs(380) <= not(inputs(25));
    layer0_outputs(381) <= (inputs(93)) or (inputs(105));
    layer0_outputs(382) <= not((inputs(96)) or (inputs(143)));
    layer0_outputs(383) <= inputs(218);
    layer0_outputs(384) <= (inputs(169)) or (inputs(2));
    layer0_outputs(385) <= not((inputs(106)) or (inputs(19)));
    layer0_outputs(386) <= not(inputs(81)) or (inputs(235));
    layer0_outputs(387) <= (inputs(187)) or (inputs(162));
    layer0_outputs(388) <= (inputs(52)) and not (inputs(16));
    layer0_outputs(389) <= not(inputs(61)) or (inputs(89));
    layer0_outputs(390) <= not(inputs(216));
    layer0_outputs(391) <= inputs(233);
    layer0_outputs(392) <= not(inputs(147));
    layer0_outputs(393) <= not((inputs(78)) or (inputs(51)));
    layer0_outputs(394) <= (inputs(37)) or (inputs(19));
    layer0_outputs(395) <= inputs(195);
    layer0_outputs(396) <= (inputs(124)) and not (inputs(190));
    layer0_outputs(397) <= (inputs(154)) or (inputs(183));
    layer0_outputs(398) <= not((inputs(27)) or (inputs(104)));
    layer0_outputs(399) <= inputs(82);
    layer0_outputs(400) <= (inputs(177)) and not (inputs(221));
    layer0_outputs(401) <= inputs(119);
    layer0_outputs(402) <= inputs(101);
    layer0_outputs(403) <= not((inputs(230)) or (inputs(46)));
    layer0_outputs(404) <= not((inputs(144)) or (inputs(228)));
    layer0_outputs(405) <= inputs(184);
    layer0_outputs(406) <= (inputs(18)) and (inputs(41));
    layer0_outputs(407) <= not(inputs(101));
    layer0_outputs(408) <= (inputs(56)) or (inputs(18));
    layer0_outputs(409) <= not(inputs(27));
    layer0_outputs(410) <= not(inputs(89)) or (inputs(142));
    layer0_outputs(411) <= (inputs(242)) xor (inputs(121));
    layer0_outputs(412) <= not(inputs(134));
    layer0_outputs(413) <= (inputs(84)) and not (inputs(1));
    layer0_outputs(414) <= (inputs(23)) and not (inputs(188));
    layer0_outputs(415) <= (inputs(231)) or (inputs(247));
    layer0_outputs(416) <= inputs(37);
    layer0_outputs(417) <= inputs(178);
    layer0_outputs(418) <= not((inputs(137)) and (inputs(250)));
    layer0_outputs(419) <= inputs(104);
    layer0_outputs(420) <= not((inputs(143)) or (inputs(99)));
    layer0_outputs(421) <= '1';
    layer0_outputs(422) <= not(inputs(130)) or (inputs(223));
    layer0_outputs(423) <= not((inputs(6)) and (inputs(11)));
    layer0_outputs(424) <= not((inputs(20)) and (inputs(19)));
    layer0_outputs(425) <= not(inputs(157));
    layer0_outputs(426) <= inputs(109);
    layer0_outputs(427) <= inputs(97);
    layer0_outputs(428) <= not(inputs(35)) or (inputs(130));
    layer0_outputs(429) <= not(inputs(233)) or (inputs(25));
    layer0_outputs(430) <= (inputs(225)) or (inputs(117));
    layer0_outputs(431) <= inputs(118);
    layer0_outputs(432) <= not((inputs(150)) or (inputs(31)));
    layer0_outputs(433) <= inputs(199);
    layer0_outputs(434) <= inputs(247);
    layer0_outputs(435) <= (inputs(221)) or (inputs(106));
    layer0_outputs(436) <= (inputs(164)) or (inputs(175));
    layer0_outputs(437) <= (inputs(224)) xor (inputs(167));
    layer0_outputs(438) <= (inputs(99)) or (inputs(180));
    layer0_outputs(439) <= (inputs(110)) and (inputs(172));
    layer0_outputs(440) <= not(inputs(228));
    layer0_outputs(441) <= not(inputs(176));
    layer0_outputs(442) <= (inputs(234)) and (inputs(233));
    layer0_outputs(443) <= (inputs(25)) and not (inputs(60));
    layer0_outputs(444) <= not((inputs(226)) or (inputs(91)));
    layer0_outputs(445) <= inputs(83);
    layer0_outputs(446) <= inputs(44);
    layer0_outputs(447) <= not((inputs(186)) and (inputs(199)));
    layer0_outputs(448) <= inputs(75);
    layer0_outputs(449) <= not(inputs(86));
    layer0_outputs(450) <= not((inputs(18)) or (inputs(105)));
    layer0_outputs(451) <= (inputs(146)) xor (inputs(253));
    layer0_outputs(452) <= not(inputs(53));
    layer0_outputs(453) <= not(inputs(100)) or (inputs(0));
    layer0_outputs(454) <= not(inputs(192)) or (inputs(238));
    layer0_outputs(455) <= inputs(28);
    layer0_outputs(456) <= not(inputs(23));
    layer0_outputs(457) <= not(inputs(37));
    layer0_outputs(458) <= not((inputs(85)) xor (inputs(96)));
    layer0_outputs(459) <= not((inputs(229)) and (inputs(106)));
    layer0_outputs(460) <= not((inputs(129)) or (inputs(93)));
    layer0_outputs(461) <= '1';
    layer0_outputs(462) <= (inputs(212)) or (inputs(211));
    layer0_outputs(463) <= (inputs(197)) or (inputs(206));
    layer0_outputs(464) <= (inputs(101)) and not (inputs(15));
    layer0_outputs(465) <= not(inputs(70));
    layer0_outputs(466) <= not((inputs(18)) or (inputs(186)));
    layer0_outputs(467) <= not(inputs(183)) or (inputs(30));
    layer0_outputs(468) <= not(inputs(240));
    layer0_outputs(469) <= not(inputs(135));
    layer0_outputs(470) <= (inputs(190)) or (inputs(233));
    layer0_outputs(471) <= '1';
    layer0_outputs(472) <= not((inputs(168)) or (inputs(33)));
    layer0_outputs(473) <= not(inputs(150));
    layer0_outputs(474) <= (inputs(55)) and not (inputs(54));
    layer0_outputs(475) <= (inputs(186)) and not (inputs(33));
    layer0_outputs(476) <= inputs(132);
    layer0_outputs(477) <= (inputs(115)) and not (inputs(142));
    layer0_outputs(478) <= (inputs(243)) and not (inputs(160));
    layer0_outputs(479) <= not(inputs(67));
    layer0_outputs(480) <= (inputs(115)) and not (inputs(150));
    layer0_outputs(481) <= inputs(102);
    layer0_outputs(482) <= (inputs(181)) and not (inputs(237));
    layer0_outputs(483) <= (inputs(21)) or (inputs(59));
    layer0_outputs(484) <= not(inputs(61));
    layer0_outputs(485) <= not((inputs(156)) or (inputs(69)));
    layer0_outputs(486) <= (inputs(40)) or (inputs(63));
    layer0_outputs(487) <= inputs(38);
    layer0_outputs(488) <= not((inputs(50)) or (inputs(112)));
    layer0_outputs(489) <= not(inputs(137)) or (inputs(207));
    layer0_outputs(490) <= inputs(73);
    layer0_outputs(491) <= (inputs(110)) xor (inputs(4));
    layer0_outputs(492) <= (inputs(13)) xor (inputs(212));
    layer0_outputs(493) <= not((inputs(245)) or (inputs(225)));
    layer0_outputs(494) <= not(inputs(59)) or (inputs(32));
    layer0_outputs(495) <= not(inputs(99));
    layer0_outputs(496) <= inputs(160);
    layer0_outputs(497) <= inputs(73);
    layer0_outputs(498) <= (inputs(15)) xor (inputs(107));
    layer0_outputs(499) <= (inputs(215)) and (inputs(249));
    layer0_outputs(500) <= (inputs(187)) or (inputs(116));
    layer0_outputs(501) <= not(inputs(105));
    layer0_outputs(502) <= (inputs(200)) and not (inputs(15));
    layer0_outputs(503) <= '0';
    layer0_outputs(504) <= (inputs(187)) and not (inputs(254));
    layer0_outputs(505) <= not((inputs(184)) or (inputs(241)));
    layer0_outputs(506) <= not((inputs(187)) or (inputs(154)));
    layer0_outputs(507) <= (inputs(255)) or (inputs(243));
    layer0_outputs(508) <= not(inputs(245));
    layer0_outputs(509) <= inputs(197);
    layer0_outputs(510) <= not(inputs(37));
    layer0_outputs(511) <= not((inputs(217)) or (inputs(211)));
    layer0_outputs(512) <= not((inputs(50)) or (inputs(38)));
    layer0_outputs(513) <= (inputs(130)) and (inputs(183));
    layer0_outputs(514) <= (inputs(115)) xor (inputs(118));
    layer0_outputs(515) <= '0';
    layer0_outputs(516) <= inputs(152);
    layer0_outputs(517) <= '1';
    layer0_outputs(518) <= (inputs(191)) or (inputs(148));
    layer0_outputs(519) <= (inputs(106)) and not (inputs(142));
    layer0_outputs(520) <= (inputs(136)) or (inputs(0));
    layer0_outputs(521) <= not(inputs(168));
    layer0_outputs(522) <= (inputs(233)) or (inputs(66));
    layer0_outputs(523) <= inputs(83);
    layer0_outputs(524) <= not(inputs(28));
    layer0_outputs(525) <= inputs(137);
    layer0_outputs(526) <= not(inputs(183));
    layer0_outputs(527) <= not(inputs(221));
    layer0_outputs(528) <= inputs(221);
    layer0_outputs(529) <= not((inputs(132)) or (inputs(52)));
    layer0_outputs(530) <= not(inputs(88)) or (inputs(241));
    layer0_outputs(531) <= inputs(74);
    layer0_outputs(532) <= (inputs(42)) and not (inputs(202));
    layer0_outputs(533) <= inputs(176);
    layer0_outputs(534) <= not((inputs(224)) or (inputs(218)));
    layer0_outputs(535) <= inputs(108);
    layer0_outputs(536) <= not((inputs(215)) or (inputs(199)));
    layer0_outputs(537) <= not((inputs(61)) xor (inputs(59)));
    layer0_outputs(538) <= not(inputs(92));
    layer0_outputs(539) <= (inputs(114)) or (inputs(36));
    layer0_outputs(540) <= inputs(115);
    layer0_outputs(541) <= (inputs(132)) and (inputs(235));
    layer0_outputs(542) <= not(inputs(102));
    layer0_outputs(543) <= inputs(81);
    layer0_outputs(544) <= inputs(116);
    layer0_outputs(545) <= inputs(77);
    layer0_outputs(546) <= not((inputs(4)) or (inputs(218)));
    layer0_outputs(547) <= not((inputs(0)) or (inputs(183)));
    layer0_outputs(548) <= not((inputs(118)) or (inputs(157)));
    layer0_outputs(549) <= (inputs(150)) and not (inputs(51));
    layer0_outputs(550) <= (inputs(4)) or (inputs(194));
    layer0_outputs(551) <= (inputs(97)) or (inputs(215));
    layer0_outputs(552) <= (inputs(87)) or (inputs(209));
    layer0_outputs(553) <= not(inputs(28)) or (inputs(72));
    layer0_outputs(554) <= not(inputs(2)) or (inputs(159));
    layer0_outputs(555) <= inputs(220);
    layer0_outputs(556) <= not((inputs(212)) xor (inputs(225)));
    layer0_outputs(557) <= (inputs(89)) or (inputs(152));
    layer0_outputs(558) <= not(inputs(68));
    layer0_outputs(559) <= not(inputs(127));
    layer0_outputs(560) <= inputs(212);
    layer0_outputs(561) <= not(inputs(36)) or (inputs(240));
    layer0_outputs(562) <= (inputs(84)) or (inputs(95));
    layer0_outputs(563) <= inputs(230);
    layer0_outputs(564) <= inputs(118);
    layer0_outputs(565) <= (inputs(253)) or (inputs(189));
    layer0_outputs(566) <= inputs(195);
    layer0_outputs(567) <= (inputs(92)) or (inputs(4));
    layer0_outputs(568) <= (inputs(4)) or (inputs(218));
    layer0_outputs(569) <= not(inputs(183));
    layer0_outputs(570) <= not(inputs(223));
    layer0_outputs(571) <= not((inputs(107)) xor (inputs(59)));
    layer0_outputs(572) <= not((inputs(145)) or (inputs(59)));
    layer0_outputs(573) <= not(inputs(169));
    layer0_outputs(574) <= not((inputs(210)) or (inputs(43)));
    layer0_outputs(575) <= (inputs(132)) or (inputs(101));
    layer0_outputs(576) <= inputs(103);
    layer0_outputs(577) <= (inputs(0)) or (inputs(136));
    layer0_outputs(578) <= inputs(104);
    layer0_outputs(579) <= inputs(69);
    layer0_outputs(580) <= (inputs(96)) or (inputs(78));
    layer0_outputs(581) <= (inputs(26)) and (inputs(1));
    layer0_outputs(582) <= not(inputs(84));
    layer0_outputs(583) <= not(inputs(195));
    layer0_outputs(584) <= not(inputs(185));
    layer0_outputs(585) <= not((inputs(14)) or (inputs(243)));
    layer0_outputs(586) <= '0';
    layer0_outputs(587) <= not(inputs(39));
    layer0_outputs(588) <= (inputs(117)) and not (inputs(221));
    layer0_outputs(589) <= not(inputs(86));
    layer0_outputs(590) <= not((inputs(17)) or (inputs(124)));
    layer0_outputs(591) <= (inputs(7)) or (inputs(126));
    layer0_outputs(592) <= not(inputs(130));
    layer0_outputs(593) <= inputs(119);
    layer0_outputs(594) <= not((inputs(109)) or (inputs(45)));
    layer0_outputs(595) <= not((inputs(58)) xor (inputs(91)));
    layer0_outputs(596) <= (inputs(227)) or (inputs(222));
    layer0_outputs(597) <= (inputs(210)) and not (inputs(103));
    layer0_outputs(598) <= not((inputs(48)) xor (inputs(16)));
    layer0_outputs(599) <= (inputs(7)) and not (inputs(253));
    layer0_outputs(600) <= (inputs(188)) or (inputs(189));
    layer0_outputs(601) <= '1';
    layer0_outputs(602) <= inputs(3);
    layer0_outputs(603) <= (inputs(94)) or (inputs(128));
    layer0_outputs(604) <= inputs(90);
    layer0_outputs(605) <= not(inputs(140));
    layer0_outputs(606) <= (inputs(138)) or (inputs(207));
    layer0_outputs(607) <= not(inputs(131));
    layer0_outputs(608) <= inputs(102);
    layer0_outputs(609) <= inputs(201);
    layer0_outputs(610) <= not((inputs(2)) or (inputs(139)));
    layer0_outputs(611) <= (inputs(39)) or (inputs(50));
    layer0_outputs(612) <= (inputs(3)) and not (inputs(247));
    layer0_outputs(613) <= '1';
    layer0_outputs(614) <= (inputs(182)) and not (inputs(18));
    layer0_outputs(615) <= (inputs(107)) or (inputs(165));
    layer0_outputs(616) <= not((inputs(111)) or (inputs(143)));
    layer0_outputs(617) <= not(inputs(59)) or (inputs(245));
    layer0_outputs(618) <= not(inputs(157));
    layer0_outputs(619) <= not((inputs(228)) xor (inputs(233)));
    layer0_outputs(620) <= inputs(34);
    layer0_outputs(621) <= (inputs(251)) or (inputs(77));
    layer0_outputs(622) <= (inputs(67)) and not (inputs(196));
    layer0_outputs(623) <= not((inputs(194)) or (inputs(195)));
    layer0_outputs(624) <= not((inputs(55)) or (inputs(214)));
    layer0_outputs(625) <= not((inputs(83)) or (inputs(176)));
    layer0_outputs(626) <= not((inputs(125)) or (inputs(6)));
    layer0_outputs(627) <= not((inputs(241)) xor (inputs(211)));
    layer0_outputs(628) <= not(inputs(188)) or (inputs(23));
    layer0_outputs(629) <= not(inputs(141));
    layer0_outputs(630) <= not(inputs(195)) or (inputs(129));
    layer0_outputs(631) <= not(inputs(39)) or (inputs(230));
    layer0_outputs(632) <= not((inputs(60)) or (inputs(43)));
    layer0_outputs(633) <= not((inputs(25)) or (inputs(77)));
    layer0_outputs(634) <= not(inputs(31));
    layer0_outputs(635) <= not((inputs(247)) or (inputs(215)));
    layer0_outputs(636) <= not(inputs(26));
    layer0_outputs(637) <= inputs(189);
    layer0_outputs(638) <= not(inputs(99));
    layer0_outputs(639) <= not(inputs(149));
    layer0_outputs(640) <= not((inputs(208)) xor (inputs(241)));
    layer0_outputs(641) <= not((inputs(133)) or (inputs(99)));
    layer0_outputs(642) <= not((inputs(255)) or (inputs(54)));
    layer0_outputs(643) <= not(inputs(210));
    layer0_outputs(644) <= (inputs(5)) or (inputs(206));
    layer0_outputs(645) <= not((inputs(90)) or (inputs(176)));
    layer0_outputs(646) <= (inputs(84)) or (inputs(236));
    layer0_outputs(647) <= not(inputs(212));
    layer0_outputs(648) <= not(inputs(119));
    layer0_outputs(649) <= not((inputs(67)) xor (inputs(48)));
    layer0_outputs(650) <= inputs(117);
    layer0_outputs(651) <= not(inputs(115));
    layer0_outputs(652) <= not(inputs(190));
    layer0_outputs(653) <= inputs(215);
    layer0_outputs(654) <= not(inputs(134));
    layer0_outputs(655) <= not(inputs(42));
    layer0_outputs(656) <= not(inputs(253)) or (inputs(222));
    layer0_outputs(657) <= not(inputs(120)) or (inputs(36));
    layer0_outputs(658) <= inputs(34);
    layer0_outputs(659) <= not(inputs(49)) or (inputs(113));
    layer0_outputs(660) <= not(inputs(118)) or (inputs(138));
    layer0_outputs(661) <= inputs(36);
    layer0_outputs(662) <= (inputs(251)) or (inputs(197));
    layer0_outputs(663) <= inputs(22);
    layer0_outputs(664) <= inputs(136);
    layer0_outputs(665) <= not(inputs(118));
    layer0_outputs(666) <= (inputs(69)) or (inputs(21));
    layer0_outputs(667) <= (inputs(104)) and not (inputs(158));
    layer0_outputs(668) <= '1';
    layer0_outputs(669) <= not(inputs(37));
    layer0_outputs(670) <= inputs(213);
    layer0_outputs(671) <= (inputs(145)) xor (inputs(84));
    layer0_outputs(672) <= not((inputs(77)) or (inputs(245)));
    layer0_outputs(673) <= (inputs(232)) and not (inputs(1));
    layer0_outputs(674) <= (inputs(12)) and not (inputs(176));
    layer0_outputs(675) <= inputs(181);
    layer0_outputs(676) <= not((inputs(235)) or (inputs(32)));
    layer0_outputs(677) <= (inputs(197)) or (inputs(206));
    layer0_outputs(678) <= not((inputs(26)) and (inputs(27)));
    layer0_outputs(679) <= (inputs(142)) or (inputs(141));
    layer0_outputs(680) <= (inputs(14)) or (inputs(218));
    layer0_outputs(681) <= not(inputs(98)) or (inputs(29));
    layer0_outputs(682) <= inputs(20);
    layer0_outputs(683) <= not((inputs(172)) xor (inputs(222)));
    layer0_outputs(684) <= not((inputs(141)) or (inputs(66)));
    layer0_outputs(685) <= not((inputs(164)) or (inputs(224)));
    layer0_outputs(686) <= not((inputs(126)) or (inputs(254)));
    layer0_outputs(687) <= not(inputs(62));
    layer0_outputs(688) <= (inputs(189)) or (inputs(159));
    layer0_outputs(689) <= (inputs(139)) or (inputs(2));
    layer0_outputs(690) <= (inputs(149)) xor (inputs(178));
    layer0_outputs(691) <= not((inputs(109)) or (inputs(164)));
    layer0_outputs(692) <= not(inputs(159));
    layer0_outputs(693) <= not(inputs(20)) or (inputs(189));
    layer0_outputs(694) <= inputs(237);
    layer0_outputs(695) <= (inputs(249)) or (inputs(81));
    layer0_outputs(696) <= not(inputs(85));
    layer0_outputs(697) <= '1';
    layer0_outputs(698) <= not(inputs(52)) or (inputs(253));
    layer0_outputs(699) <= inputs(135);
    layer0_outputs(700) <= not((inputs(243)) or (inputs(202)));
    layer0_outputs(701) <= not(inputs(103)) or (inputs(163));
    layer0_outputs(702) <= inputs(4);
    layer0_outputs(703) <= inputs(194);
    layer0_outputs(704) <= (inputs(165)) and not (inputs(21));
    layer0_outputs(705) <= inputs(159);
    layer0_outputs(706) <= not(inputs(13));
    layer0_outputs(707) <= (inputs(126)) or (inputs(184));
    layer0_outputs(708) <= not(inputs(104));
    layer0_outputs(709) <= not(inputs(120));
    layer0_outputs(710) <= not(inputs(42)) or (inputs(154));
    layer0_outputs(711) <= (inputs(27)) or (inputs(214));
    layer0_outputs(712) <= not(inputs(168)) or (inputs(62));
    layer0_outputs(713) <= not(inputs(56));
    layer0_outputs(714) <= not((inputs(178)) or (inputs(203)));
    layer0_outputs(715) <= not(inputs(35));
    layer0_outputs(716) <= not(inputs(100));
    layer0_outputs(717) <= '1';
    layer0_outputs(718) <= inputs(83);
    layer0_outputs(719) <= not(inputs(189));
    layer0_outputs(720) <= not(inputs(172));
    layer0_outputs(721) <= (inputs(203)) and (inputs(233));
    layer0_outputs(722) <= inputs(213);
    layer0_outputs(723) <= (inputs(182)) and not (inputs(66));
    layer0_outputs(724) <= (inputs(221)) or (inputs(25));
    layer0_outputs(725) <= not(inputs(195));
    layer0_outputs(726) <= not(inputs(102));
    layer0_outputs(727) <= (inputs(193)) or (inputs(202));
    layer0_outputs(728) <= not(inputs(118));
    layer0_outputs(729) <= not((inputs(164)) or (inputs(180)));
    layer0_outputs(730) <= (inputs(218)) or (inputs(203));
    layer0_outputs(731) <= not((inputs(254)) or (inputs(135)));
    layer0_outputs(732) <= (inputs(162)) or (inputs(113));
    layer0_outputs(733) <= not(inputs(164));
    layer0_outputs(734) <= not((inputs(218)) xor (inputs(111)));
    layer0_outputs(735) <= not((inputs(38)) or (inputs(54)));
    layer0_outputs(736) <= not(inputs(51));
    layer0_outputs(737) <= not(inputs(10)) or (inputs(112));
    layer0_outputs(738) <= not(inputs(233)) or (inputs(92));
    layer0_outputs(739) <= (inputs(199)) and not (inputs(231));
    layer0_outputs(740) <= inputs(57);
    layer0_outputs(741) <= not(inputs(195));
    layer0_outputs(742) <= not((inputs(64)) or (inputs(244)));
    layer0_outputs(743) <= not(inputs(225)) or (inputs(40));
    layer0_outputs(744) <= (inputs(45)) xor (inputs(28));
    layer0_outputs(745) <= (inputs(98)) or (inputs(114));
    layer0_outputs(746) <= (inputs(22)) and not (inputs(27));
    layer0_outputs(747) <= not((inputs(174)) and (inputs(255)));
    layer0_outputs(748) <= not(inputs(38));
    layer0_outputs(749) <= not(inputs(153)) or (inputs(210));
    layer0_outputs(750) <= not((inputs(217)) or (inputs(102)));
    layer0_outputs(751) <= not((inputs(188)) xor (inputs(129)));
    layer0_outputs(752) <= inputs(107);
    layer0_outputs(753) <= not(inputs(133)) or (inputs(149));
    layer0_outputs(754) <= not((inputs(188)) or (inputs(63)));
    layer0_outputs(755) <= not((inputs(110)) or (inputs(38)));
    layer0_outputs(756) <= not(inputs(87));
    layer0_outputs(757) <= not(inputs(100));
    layer0_outputs(758) <= inputs(68);
    layer0_outputs(759) <= (inputs(157)) or (inputs(155));
    layer0_outputs(760) <= (inputs(100)) or (inputs(47));
    layer0_outputs(761) <= not(inputs(73)) or (inputs(109));
    layer0_outputs(762) <= not(inputs(12)) or (inputs(53));
    layer0_outputs(763) <= not(inputs(74)) or (inputs(176));
    layer0_outputs(764) <= (inputs(100)) and not (inputs(30));
    layer0_outputs(765) <= inputs(105);
    layer0_outputs(766) <= not((inputs(248)) or (inputs(208)));
    layer0_outputs(767) <= (inputs(172)) and not (inputs(79));
    layer0_outputs(768) <= not(inputs(94));
    layer0_outputs(769) <= (inputs(95)) and not (inputs(237));
    layer0_outputs(770) <= not(inputs(197));
    layer0_outputs(771) <= '0';
    layer0_outputs(772) <= (inputs(204)) and (inputs(199));
    layer0_outputs(773) <= not(inputs(228)) or (inputs(45));
    layer0_outputs(774) <= (inputs(242)) xor (inputs(43));
    layer0_outputs(775) <= not(inputs(106));
    layer0_outputs(776) <= (inputs(160)) or (inputs(129));
    layer0_outputs(777) <= inputs(44);
    layer0_outputs(778) <= not((inputs(240)) and (inputs(9)));
    layer0_outputs(779) <= not((inputs(49)) or (inputs(44)));
    layer0_outputs(780) <= (inputs(37)) and not (inputs(32));
    layer0_outputs(781) <= not(inputs(154)) or (inputs(32));
    layer0_outputs(782) <= not((inputs(144)) or (inputs(42)));
    layer0_outputs(783) <= (inputs(251)) or (inputs(107));
    layer0_outputs(784) <= not((inputs(1)) xor (inputs(123)));
    layer0_outputs(785) <= not(inputs(97));
    layer0_outputs(786) <= (inputs(204)) or (inputs(224));
    layer0_outputs(787) <= not(inputs(90));
    layer0_outputs(788) <= inputs(115);
    layer0_outputs(789) <= inputs(110);
    layer0_outputs(790) <= (inputs(132)) and not (inputs(193));
    layer0_outputs(791) <= not(inputs(234)) or (inputs(144));
    layer0_outputs(792) <= not(inputs(135));
    layer0_outputs(793) <= not(inputs(152)) or (inputs(155));
    layer0_outputs(794) <= not(inputs(151));
    layer0_outputs(795) <= (inputs(184)) or (inputs(147));
    layer0_outputs(796) <= not(inputs(96));
    layer0_outputs(797) <= (inputs(206)) or (inputs(186));
    layer0_outputs(798) <= inputs(212);
    layer0_outputs(799) <= not(inputs(25));
    layer0_outputs(800) <= not(inputs(121)) or (inputs(241));
    layer0_outputs(801) <= '0';
    layer0_outputs(802) <= inputs(243);
    layer0_outputs(803) <= (inputs(129)) or (inputs(115));
    layer0_outputs(804) <= (inputs(69)) and not (inputs(195));
    layer0_outputs(805) <= not(inputs(187));
    layer0_outputs(806) <= not(inputs(155));
    layer0_outputs(807) <= not(inputs(197));
    layer0_outputs(808) <= (inputs(137)) and not (inputs(236));
    layer0_outputs(809) <= inputs(180);
    layer0_outputs(810) <= not((inputs(219)) or (inputs(138)));
    layer0_outputs(811) <= inputs(230);
    layer0_outputs(812) <= not((inputs(166)) and (inputs(25)));
    layer0_outputs(813) <= not((inputs(234)) or (inputs(237)));
    layer0_outputs(814) <= not((inputs(51)) or (inputs(238)));
    layer0_outputs(815) <= '0';
    layer0_outputs(816) <= (inputs(45)) or (inputs(246));
    layer0_outputs(817) <= not(inputs(43)) or (inputs(160));
    layer0_outputs(818) <= not(inputs(118));
    layer0_outputs(819) <= not(inputs(120));
    layer0_outputs(820) <= (inputs(122)) and not (inputs(7));
    layer0_outputs(821) <= inputs(189);
    layer0_outputs(822) <= not(inputs(112));
    layer0_outputs(823) <= not(inputs(124)) or (inputs(52));
    layer0_outputs(824) <= (inputs(104)) and not (inputs(222));
    layer0_outputs(825) <= (inputs(247)) and not (inputs(255));
    layer0_outputs(826) <= (inputs(161)) xor (inputs(133));
    layer0_outputs(827) <= (inputs(91)) and not (inputs(112));
    layer0_outputs(828) <= not(inputs(101)) or (inputs(196));
    layer0_outputs(829) <= not(inputs(167));
    layer0_outputs(830) <= (inputs(185)) or (inputs(201));
    layer0_outputs(831) <= not(inputs(38));
    layer0_outputs(832) <= inputs(183);
    layer0_outputs(833) <= '0';
    layer0_outputs(834) <= inputs(226);
    layer0_outputs(835) <= (inputs(38)) xor (inputs(229));
    layer0_outputs(836) <= not(inputs(57)) or (inputs(163));
    layer0_outputs(837) <= not(inputs(99));
    layer0_outputs(838) <= inputs(105);
    layer0_outputs(839) <= not(inputs(99)) or (inputs(207));
    layer0_outputs(840) <= inputs(140);
    layer0_outputs(841) <= not(inputs(255));
    layer0_outputs(842) <= (inputs(234)) or (inputs(253));
    layer0_outputs(843) <= not((inputs(174)) xor (inputs(254)));
    layer0_outputs(844) <= (inputs(191)) or (inputs(203));
    layer0_outputs(845) <= '0';
    layer0_outputs(846) <= not(inputs(10)) or (inputs(34));
    layer0_outputs(847) <= (inputs(108)) or (inputs(146));
    layer0_outputs(848) <= (inputs(10)) xor (inputs(174));
    layer0_outputs(849) <= not(inputs(114)) or (inputs(50));
    layer0_outputs(850) <= (inputs(88)) and not (inputs(218));
    layer0_outputs(851) <= (inputs(246)) or (inputs(44));
    layer0_outputs(852) <= inputs(93);
    layer0_outputs(853) <= not((inputs(111)) or (inputs(157)));
    layer0_outputs(854) <= not(inputs(99));
    layer0_outputs(855) <= not((inputs(249)) xor (inputs(70)));
    layer0_outputs(856) <= not(inputs(204));
    layer0_outputs(857) <= not((inputs(171)) or (inputs(129)));
    layer0_outputs(858) <= (inputs(89)) or (inputs(0));
    layer0_outputs(859) <= not((inputs(210)) or (inputs(212)));
    layer0_outputs(860) <= inputs(147);
    layer0_outputs(861) <= not(inputs(147));
    layer0_outputs(862) <= not(inputs(25));
    layer0_outputs(863) <= not((inputs(44)) or (inputs(192)));
    layer0_outputs(864) <= (inputs(208)) or (inputs(105));
    layer0_outputs(865) <= (inputs(85)) and not (inputs(191));
    layer0_outputs(866) <= (inputs(161)) and not (inputs(222));
    layer0_outputs(867) <= not(inputs(161));
    layer0_outputs(868) <= (inputs(186)) and not (inputs(236));
    layer0_outputs(869) <= (inputs(28)) and not (inputs(32));
    layer0_outputs(870) <= not(inputs(109)) or (inputs(239));
    layer0_outputs(871) <= inputs(202);
    layer0_outputs(872) <= (inputs(174)) and not (inputs(93));
    layer0_outputs(873) <= inputs(226);
    layer0_outputs(874) <= not(inputs(132));
    layer0_outputs(875) <= not(inputs(103));
    layer0_outputs(876) <= not((inputs(13)) or (inputs(160)));
    layer0_outputs(877) <= inputs(168);
    layer0_outputs(878) <= (inputs(177)) xor (inputs(209));
    layer0_outputs(879) <= not(inputs(231));
    layer0_outputs(880) <= '1';
    layer0_outputs(881) <= (inputs(13)) xor (inputs(126));
    layer0_outputs(882) <= not(inputs(110));
    layer0_outputs(883) <= inputs(153);
    layer0_outputs(884) <= '1';
    layer0_outputs(885) <= inputs(225);
    layer0_outputs(886) <= not((inputs(213)) or (inputs(229)));
    layer0_outputs(887) <= not(inputs(57));
    layer0_outputs(888) <= (inputs(136)) and not (inputs(5));
    layer0_outputs(889) <= inputs(194);
    layer0_outputs(890) <= inputs(115);
    layer0_outputs(891) <= inputs(18);
    layer0_outputs(892) <= (inputs(233)) and (inputs(254));
    layer0_outputs(893) <= (inputs(31)) or (inputs(254));
    layer0_outputs(894) <= inputs(159);
    layer0_outputs(895) <= (inputs(121)) or (inputs(45));
    layer0_outputs(896) <= not(inputs(232));
    layer0_outputs(897) <= inputs(97);
    layer0_outputs(898) <= inputs(114);
    layer0_outputs(899) <= inputs(93);
    layer0_outputs(900) <= inputs(134);
    layer0_outputs(901) <= inputs(104);
    layer0_outputs(902) <= inputs(219);
    layer0_outputs(903) <= not((inputs(239)) xor (inputs(173)));
    layer0_outputs(904) <= inputs(106);
    layer0_outputs(905) <= not(inputs(21));
    layer0_outputs(906) <= (inputs(57)) and not (inputs(209));
    layer0_outputs(907) <= not(inputs(130));
    layer0_outputs(908) <= not((inputs(189)) and (inputs(245)));
    layer0_outputs(909) <= not((inputs(89)) or (inputs(225)));
    layer0_outputs(910) <= not(inputs(133));
    layer0_outputs(911) <= (inputs(21)) or (inputs(61));
    layer0_outputs(912) <= not((inputs(111)) or (inputs(24)));
    layer0_outputs(913) <= not(inputs(97));
    layer0_outputs(914) <= (inputs(138)) and not (inputs(193));
    layer0_outputs(915) <= inputs(167);
    layer0_outputs(916) <= (inputs(158)) or (inputs(117));
    layer0_outputs(917) <= not(inputs(7));
    layer0_outputs(918) <= inputs(117);
    layer0_outputs(919) <= (inputs(221)) or (inputs(182));
    layer0_outputs(920) <= inputs(102);
    layer0_outputs(921) <= '1';
    layer0_outputs(922) <= not((inputs(20)) or (inputs(163)));
    layer0_outputs(923) <= (inputs(243)) or (inputs(209));
    layer0_outputs(924) <= inputs(103);
    layer0_outputs(925) <= '0';
    layer0_outputs(926) <= not((inputs(74)) or (inputs(73)));
    layer0_outputs(927) <= (inputs(250)) or (inputs(87));
    layer0_outputs(928) <= not((inputs(147)) or (inputs(147)));
    layer0_outputs(929) <= not(inputs(163));
    layer0_outputs(930) <= (inputs(182)) or (inputs(188));
    layer0_outputs(931) <= (inputs(241)) or (inputs(77));
    layer0_outputs(932) <= (inputs(34)) xor (inputs(63));
    layer0_outputs(933) <= not((inputs(198)) xor (inputs(96)));
    layer0_outputs(934) <= not((inputs(75)) or (inputs(82)));
    layer0_outputs(935) <= not((inputs(79)) xor (inputs(142)));
    layer0_outputs(936) <= not((inputs(39)) and (inputs(207)));
    layer0_outputs(937) <= (inputs(159)) xor (inputs(88));
    layer0_outputs(938) <= (inputs(204)) or (inputs(202));
    layer0_outputs(939) <= not(inputs(231));
    layer0_outputs(940) <= not((inputs(243)) and (inputs(201)));
    layer0_outputs(941) <= not(inputs(29));
    layer0_outputs(942) <= not(inputs(235)) or (inputs(44));
    layer0_outputs(943) <= not(inputs(63));
    layer0_outputs(944) <= not((inputs(115)) or (inputs(149)));
    layer0_outputs(945) <= not(inputs(160)) or (inputs(2));
    layer0_outputs(946) <= not((inputs(84)) xor (inputs(15)));
    layer0_outputs(947) <= not(inputs(5));
    layer0_outputs(948) <= not(inputs(169)) or (inputs(242));
    layer0_outputs(949) <= not(inputs(123)) or (inputs(191));
    layer0_outputs(950) <= not(inputs(191));
    layer0_outputs(951) <= inputs(99);
    layer0_outputs(952) <= not(inputs(170));
    layer0_outputs(953) <= (inputs(112)) and not (inputs(236));
    layer0_outputs(954) <= (inputs(213)) and not (inputs(17));
    layer0_outputs(955) <= inputs(69);
    layer0_outputs(956) <= inputs(167);
    layer0_outputs(957) <= not((inputs(217)) or (inputs(206)));
    layer0_outputs(958) <= not((inputs(195)) or (inputs(180)));
    layer0_outputs(959) <= not(inputs(82));
    layer0_outputs(960) <= not((inputs(216)) or (inputs(129)));
    layer0_outputs(961) <= not(inputs(208)) or (inputs(129));
    layer0_outputs(962) <= not(inputs(1));
    layer0_outputs(963) <= (inputs(53)) and not (inputs(15));
    layer0_outputs(964) <= not(inputs(13));
    layer0_outputs(965) <= (inputs(161)) or (inputs(231));
    layer0_outputs(966) <= not(inputs(105)) or (inputs(232));
    layer0_outputs(967) <= (inputs(72)) and not (inputs(124));
    layer0_outputs(968) <= inputs(137);
    layer0_outputs(969) <= not((inputs(233)) and (inputs(47)));
    layer0_outputs(970) <= not(inputs(100));
    layer0_outputs(971) <= '1';
    layer0_outputs(972) <= (inputs(136)) and not (inputs(176));
    layer0_outputs(973) <= (inputs(27)) or (inputs(173));
    layer0_outputs(974) <= (inputs(165)) and not (inputs(21));
    layer0_outputs(975) <= not((inputs(206)) or (inputs(162)));
    layer0_outputs(976) <= not((inputs(49)) xor (inputs(223)));
    layer0_outputs(977) <= (inputs(248)) and not (inputs(66));
    layer0_outputs(978) <= (inputs(11)) xor (inputs(73));
    layer0_outputs(979) <= not(inputs(40)) or (inputs(96));
    layer0_outputs(980) <= not(inputs(23)) or (inputs(181));
    layer0_outputs(981) <= not(inputs(162));
    layer0_outputs(982) <= inputs(211);
    layer0_outputs(983) <= not(inputs(95)) or (inputs(144));
    layer0_outputs(984) <= inputs(52);
    layer0_outputs(985) <= not((inputs(129)) or (inputs(158)));
    layer0_outputs(986) <= not((inputs(211)) or (inputs(229)));
    layer0_outputs(987) <= '1';
    layer0_outputs(988) <= not(inputs(135));
    layer0_outputs(989) <= inputs(245);
    layer0_outputs(990) <= not((inputs(18)) or (inputs(230)));
    layer0_outputs(991) <= not(inputs(246));
    layer0_outputs(992) <= (inputs(31)) xor (inputs(55));
    layer0_outputs(993) <= not((inputs(63)) or (inputs(133)));
    layer0_outputs(994) <= inputs(204);
    layer0_outputs(995) <= not((inputs(192)) or (inputs(227)));
    layer0_outputs(996) <= (inputs(81)) or (inputs(53));
    layer0_outputs(997) <= (inputs(64)) or (inputs(252));
    layer0_outputs(998) <= not((inputs(96)) or (inputs(110)));
    layer0_outputs(999) <= not((inputs(128)) or (inputs(183)));
    layer0_outputs(1000) <= not(inputs(84)) or (inputs(32));
    layer0_outputs(1001) <= (inputs(74)) and not (inputs(131));
    layer0_outputs(1002) <= not(inputs(52)) or (inputs(223));
    layer0_outputs(1003) <= not((inputs(89)) xor (inputs(70)));
    layer0_outputs(1004) <= not((inputs(78)) or (inputs(39)));
    layer0_outputs(1005) <= not((inputs(3)) or (inputs(36)));
    layer0_outputs(1006) <= not((inputs(162)) or (inputs(148)));
    layer0_outputs(1007) <= inputs(121);
    layer0_outputs(1008) <= not(inputs(41));
    layer0_outputs(1009) <= not(inputs(254));
    layer0_outputs(1010) <= not(inputs(183));
    layer0_outputs(1011) <= inputs(20);
    layer0_outputs(1012) <= not(inputs(196));
    layer0_outputs(1013) <= not(inputs(231)) or (inputs(22));
    layer0_outputs(1014) <= not((inputs(169)) xor (inputs(155)));
    layer0_outputs(1015) <= inputs(148);
    layer0_outputs(1016) <= inputs(145);
    layer0_outputs(1017) <= not(inputs(106));
    layer0_outputs(1018) <= (inputs(132)) and not (inputs(227));
    layer0_outputs(1019) <= not(inputs(200)) or (inputs(18));
    layer0_outputs(1020) <= not(inputs(16));
    layer0_outputs(1021) <= not(inputs(149)) or (inputs(53));
    layer0_outputs(1022) <= not(inputs(44)) or (inputs(160));
    layer0_outputs(1023) <= (inputs(214)) and not (inputs(90));
    layer0_outputs(1024) <= (inputs(81)) xor (inputs(4));
    layer0_outputs(1025) <= not(inputs(0));
    layer0_outputs(1026) <= (inputs(116)) or (inputs(226));
    layer0_outputs(1027) <= not(inputs(151)) or (inputs(130));
    layer0_outputs(1028) <= (inputs(220)) and not (inputs(123));
    layer0_outputs(1029) <= not(inputs(198)) or (inputs(62));
    layer0_outputs(1030) <= not(inputs(67));
    layer0_outputs(1031) <= (inputs(112)) or (inputs(145));
    layer0_outputs(1032) <= not(inputs(23));
    layer0_outputs(1033) <= not(inputs(211));
    layer0_outputs(1034) <= not((inputs(213)) and (inputs(191)));
    layer0_outputs(1035) <= not(inputs(46));
    layer0_outputs(1036) <= '1';
    layer0_outputs(1037) <= not((inputs(229)) or (inputs(157)));
    layer0_outputs(1038) <= inputs(124);
    layer0_outputs(1039) <= (inputs(185)) or (inputs(140));
    layer0_outputs(1040) <= inputs(138);
    layer0_outputs(1041) <= (inputs(223)) or (inputs(65));
    layer0_outputs(1042) <= not((inputs(51)) or (inputs(211)));
    layer0_outputs(1043) <= not((inputs(222)) or (inputs(208)));
    layer0_outputs(1044) <= (inputs(156)) and not (inputs(176));
    layer0_outputs(1045) <= (inputs(127)) or (inputs(220));
    layer0_outputs(1046) <= not((inputs(49)) or (inputs(122)));
    layer0_outputs(1047) <= inputs(231);
    layer0_outputs(1048) <= not(inputs(108)) or (inputs(208));
    layer0_outputs(1049) <= not(inputs(35)) or (inputs(236));
    layer0_outputs(1050) <= (inputs(83)) or (inputs(69));
    layer0_outputs(1051) <= inputs(4);
    layer0_outputs(1052) <= not((inputs(81)) or (inputs(97)));
    layer0_outputs(1053) <= not(inputs(157));
    layer0_outputs(1054) <= (inputs(13)) and not (inputs(60));
    layer0_outputs(1055) <= not(inputs(70));
    layer0_outputs(1056) <= (inputs(229)) and not (inputs(29));
    layer0_outputs(1057) <= (inputs(164)) or (inputs(206));
    layer0_outputs(1058) <= inputs(14);
    layer0_outputs(1059) <= (inputs(207)) or (inputs(62));
    layer0_outputs(1060) <= (inputs(85)) and not (inputs(190));
    layer0_outputs(1061) <= not((inputs(75)) xor (inputs(107)));
    layer0_outputs(1062) <= (inputs(142)) or (inputs(114));
    layer0_outputs(1063) <= not(inputs(93));
    layer0_outputs(1064) <= not((inputs(37)) xor (inputs(77)));
    layer0_outputs(1065) <= inputs(103);
    layer0_outputs(1066) <= not((inputs(71)) xor (inputs(101)));
    layer0_outputs(1067) <= (inputs(53)) or (inputs(16));
    layer0_outputs(1068) <= (inputs(230)) and not (inputs(0));
    layer0_outputs(1069) <= '1';
    layer0_outputs(1070) <= (inputs(42)) or (inputs(175));
    layer0_outputs(1071) <= (inputs(82)) and not (inputs(61));
    layer0_outputs(1072) <= not(inputs(251));
    layer0_outputs(1073) <= inputs(121);
    layer0_outputs(1074) <= inputs(91);
    layer0_outputs(1075) <= not(inputs(155)) or (inputs(57));
    layer0_outputs(1076) <= not((inputs(179)) or (inputs(173)));
    layer0_outputs(1077) <= not(inputs(207));
    layer0_outputs(1078) <= (inputs(92)) or (inputs(47));
    layer0_outputs(1079) <= not(inputs(41)) or (inputs(71));
    layer0_outputs(1080) <= (inputs(153)) or (inputs(166));
    layer0_outputs(1081) <= not((inputs(161)) or (inputs(64)));
    layer0_outputs(1082) <= (inputs(44)) and not (inputs(58));
    layer0_outputs(1083) <= (inputs(200)) and (inputs(251));
    layer0_outputs(1084) <= inputs(86);
    layer0_outputs(1085) <= inputs(245);
    layer0_outputs(1086) <= (inputs(136)) and not (inputs(224));
    layer0_outputs(1087) <= (inputs(27)) and not (inputs(208));
    layer0_outputs(1088) <= inputs(246);
    layer0_outputs(1089) <= (inputs(238)) or (inputs(107));
    layer0_outputs(1090) <= not((inputs(182)) or (inputs(30)));
    layer0_outputs(1091) <= inputs(154);
    layer0_outputs(1092) <= not(inputs(179));
    layer0_outputs(1093) <= not(inputs(145)) or (inputs(1));
    layer0_outputs(1094) <= inputs(166);
    layer0_outputs(1095) <= (inputs(228)) or (inputs(100));
    layer0_outputs(1096) <= inputs(45);
    layer0_outputs(1097) <= not((inputs(144)) or (inputs(144)));
    layer0_outputs(1098) <= inputs(60);
    layer0_outputs(1099) <= inputs(214);
    layer0_outputs(1100) <= not((inputs(43)) or (inputs(65)));
    layer0_outputs(1101) <= not(inputs(123)) or (inputs(82));
    layer0_outputs(1102) <= '1';
    layer0_outputs(1103) <= (inputs(235)) and (inputs(249));
    layer0_outputs(1104) <= inputs(8);
    layer0_outputs(1105) <= not((inputs(131)) or (inputs(64)));
    layer0_outputs(1106) <= not(inputs(138)) or (inputs(224));
    layer0_outputs(1107) <= not((inputs(88)) xor (inputs(78)));
    layer0_outputs(1108) <= inputs(166);
    layer0_outputs(1109) <= inputs(9);
    layer0_outputs(1110) <= (inputs(228)) and not (inputs(46));
    layer0_outputs(1111) <= inputs(185);
    layer0_outputs(1112) <= (inputs(242)) or (inputs(205));
    layer0_outputs(1113) <= not(inputs(147)) or (inputs(16));
    layer0_outputs(1114) <= not((inputs(2)) and (inputs(244)));
    layer0_outputs(1115) <= inputs(161);
    layer0_outputs(1116) <= not(inputs(226));
    layer0_outputs(1117) <= (inputs(24)) and not (inputs(130));
    layer0_outputs(1118) <= (inputs(58)) or (inputs(191));
    layer0_outputs(1119) <= inputs(178);
    layer0_outputs(1120) <= (inputs(215)) and not (inputs(254));
    layer0_outputs(1121) <= inputs(255);
    layer0_outputs(1122) <= (inputs(67)) or (inputs(169));
    layer0_outputs(1123) <= (inputs(134)) or (inputs(105));
    layer0_outputs(1124) <= (inputs(56)) and not (inputs(252));
    layer0_outputs(1125) <= not(inputs(26));
    layer0_outputs(1126) <= inputs(98);
    layer0_outputs(1127) <= not(inputs(240)) or (inputs(66));
    layer0_outputs(1128) <= inputs(73);
    layer0_outputs(1129) <= not(inputs(103));
    layer0_outputs(1130) <= (inputs(166)) or (inputs(75));
    layer0_outputs(1131) <= not((inputs(54)) or (inputs(113)));
    layer0_outputs(1132) <= (inputs(110)) or (inputs(216));
    layer0_outputs(1133) <= not(inputs(31));
    layer0_outputs(1134) <= (inputs(108)) or (inputs(111));
    layer0_outputs(1135) <= not(inputs(188));
    layer0_outputs(1136) <= (inputs(204)) or (inputs(0));
    layer0_outputs(1137) <= (inputs(236)) and not (inputs(143));
    layer0_outputs(1138) <= not(inputs(247));
    layer0_outputs(1139) <= not(inputs(102)) or (inputs(16));
    layer0_outputs(1140) <= not(inputs(99)) or (inputs(177));
    layer0_outputs(1141) <= inputs(130);
    layer0_outputs(1142) <= (inputs(63)) and not (inputs(126));
    layer0_outputs(1143) <= not((inputs(158)) and (inputs(66)));
    layer0_outputs(1144) <= (inputs(27)) and (inputs(38));
    layer0_outputs(1145) <= (inputs(194)) xor (inputs(187));
    layer0_outputs(1146) <= inputs(105);
    layer0_outputs(1147) <= (inputs(151)) and not (inputs(132));
    layer0_outputs(1148) <= not((inputs(253)) or (inputs(8)));
    layer0_outputs(1149) <= inputs(161);
    layer0_outputs(1150) <= (inputs(77)) or (inputs(186));
    layer0_outputs(1151) <= (inputs(67)) or (inputs(38));
    layer0_outputs(1152) <= (inputs(162)) and not (inputs(40));
    layer0_outputs(1153) <= not(inputs(132));
    layer0_outputs(1154) <= inputs(181);
    layer0_outputs(1155) <= not((inputs(225)) xor (inputs(195)));
    layer0_outputs(1156) <= not(inputs(90));
    layer0_outputs(1157) <= not((inputs(116)) or (inputs(247)));
    layer0_outputs(1158) <= (inputs(199)) and not (inputs(135));
    layer0_outputs(1159) <= not((inputs(81)) and (inputs(135)));
    layer0_outputs(1160) <= not(inputs(235)) or (inputs(15));
    layer0_outputs(1161) <= not(inputs(228)) or (inputs(88));
    layer0_outputs(1162) <= (inputs(103)) or (inputs(207));
    layer0_outputs(1163) <= not(inputs(119));
    layer0_outputs(1164) <= (inputs(71)) or (inputs(72));
    layer0_outputs(1165) <= not(inputs(215)) or (inputs(17));
    layer0_outputs(1166) <= not((inputs(197)) or (inputs(188)));
    layer0_outputs(1167) <= (inputs(155)) or (inputs(253));
    layer0_outputs(1168) <= not((inputs(62)) or (inputs(76)));
    layer0_outputs(1169) <= not((inputs(208)) xor (inputs(196)));
    layer0_outputs(1170) <= (inputs(73)) or (inputs(80));
    layer0_outputs(1171) <= not((inputs(200)) or (inputs(193)));
    layer0_outputs(1172) <= inputs(174);
    layer0_outputs(1173) <= not(inputs(135));
    layer0_outputs(1174) <= not((inputs(144)) xor (inputs(118)));
    layer0_outputs(1175) <= inputs(116);
    layer0_outputs(1176) <= inputs(75);
    layer0_outputs(1177) <= not(inputs(9)) or (inputs(143));
    layer0_outputs(1178) <= not(inputs(156));
    layer0_outputs(1179) <= not(inputs(26));
    layer0_outputs(1180) <= inputs(24);
    layer0_outputs(1181) <= not((inputs(58)) or (inputs(110)));
    layer0_outputs(1182) <= not(inputs(234));
    layer0_outputs(1183) <= not(inputs(146));
    layer0_outputs(1184) <= not(inputs(14));
    layer0_outputs(1185) <= '0';
    layer0_outputs(1186) <= (inputs(103)) xor (inputs(83));
    layer0_outputs(1187) <= not(inputs(52));
    layer0_outputs(1188) <= not((inputs(42)) or (inputs(95)));
    layer0_outputs(1189) <= inputs(75);
    layer0_outputs(1190) <= inputs(239);
    layer0_outputs(1191) <= (inputs(22)) or (inputs(50));
    layer0_outputs(1192) <= (inputs(146)) or (inputs(143));
    layer0_outputs(1193) <= (inputs(230)) and not (inputs(197));
    layer0_outputs(1194) <= (inputs(242)) or (inputs(212));
    layer0_outputs(1195) <= not(inputs(115));
    layer0_outputs(1196) <= (inputs(196)) xor (inputs(227));
    layer0_outputs(1197) <= not((inputs(175)) or (inputs(204)));
    layer0_outputs(1198) <= (inputs(109)) and (inputs(116));
    layer0_outputs(1199) <= inputs(93);
    layer0_outputs(1200) <= '0';
    layer0_outputs(1201) <= not(inputs(168)) or (inputs(2));
    layer0_outputs(1202) <= not(inputs(231)) or (inputs(182));
    layer0_outputs(1203) <= (inputs(128)) or (inputs(63));
    layer0_outputs(1204) <= not((inputs(252)) or (inputs(100)));
    layer0_outputs(1205) <= (inputs(49)) and not (inputs(240));
    layer0_outputs(1206) <= not(inputs(124));
    layer0_outputs(1207) <= (inputs(102)) or (inputs(174));
    layer0_outputs(1208) <= not(inputs(52));
    layer0_outputs(1209) <= (inputs(192)) and not (inputs(47));
    layer0_outputs(1210) <= not(inputs(84));
    layer0_outputs(1211) <= (inputs(75)) and not (inputs(255));
    layer0_outputs(1212) <= not(inputs(205)) or (inputs(159));
    layer0_outputs(1213) <= (inputs(39)) and not (inputs(31));
    layer0_outputs(1214) <= not((inputs(86)) or (inputs(246)));
    layer0_outputs(1215) <= not(inputs(253)) or (inputs(67));
    layer0_outputs(1216) <= not(inputs(89));
    layer0_outputs(1217) <= not(inputs(124));
    layer0_outputs(1218) <= (inputs(173)) and not (inputs(24));
    layer0_outputs(1219) <= not(inputs(209));
    layer0_outputs(1220) <= not((inputs(41)) xor (inputs(249)));
    layer0_outputs(1221) <= (inputs(92)) or (inputs(37));
    layer0_outputs(1222) <= inputs(59);
    layer0_outputs(1223) <= not((inputs(220)) or (inputs(47)));
    layer0_outputs(1224) <= (inputs(156)) and not (inputs(47));
    layer0_outputs(1225) <= inputs(173);
    layer0_outputs(1226) <= inputs(91);
    layer0_outputs(1227) <= not((inputs(1)) or (inputs(108)));
    layer0_outputs(1228) <= not((inputs(242)) or (inputs(222)));
    layer0_outputs(1229) <= inputs(82);
    layer0_outputs(1230) <= not((inputs(201)) xor (inputs(201)));
    layer0_outputs(1231) <= not((inputs(210)) or (inputs(4)));
    layer0_outputs(1232) <= not((inputs(148)) or (inputs(174)));
    layer0_outputs(1233) <= not(inputs(248));
    layer0_outputs(1234) <= not((inputs(21)) or (inputs(10)));
    layer0_outputs(1235) <= inputs(108);
    layer0_outputs(1236) <= not((inputs(215)) and (inputs(51)));
    layer0_outputs(1237) <= inputs(217);
    layer0_outputs(1238) <= not(inputs(134));
    layer0_outputs(1239) <= not(inputs(94));
    layer0_outputs(1240) <= not((inputs(144)) or (inputs(71)));
    layer0_outputs(1241) <= not((inputs(225)) or (inputs(157)));
    layer0_outputs(1242) <= (inputs(198)) and (inputs(94));
    layer0_outputs(1243) <= (inputs(85)) and not (inputs(64));
    layer0_outputs(1244) <= inputs(164);
    layer0_outputs(1245) <= (inputs(170)) and (inputs(214));
    layer0_outputs(1246) <= not(inputs(151));
    layer0_outputs(1247) <= (inputs(15)) or (inputs(212));
    layer0_outputs(1248) <= not((inputs(148)) or (inputs(62)));
    layer0_outputs(1249) <= (inputs(203)) and not (inputs(25));
    layer0_outputs(1250) <= inputs(181);
    layer0_outputs(1251) <= not(inputs(217)) or (inputs(197));
    layer0_outputs(1252) <= inputs(119);
    layer0_outputs(1253) <= not(inputs(153));
    layer0_outputs(1254) <= (inputs(41)) and not (inputs(161));
    layer0_outputs(1255) <= not((inputs(200)) and (inputs(136)));
    layer0_outputs(1256) <= (inputs(126)) and (inputs(52));
    layer0_outputs(1257) <= not(inputs(6)) or (inputs(144));
    layer0_outputs(1258) <= not(inputs(103));
    layer0_outputs(1259) <= (inputs(186)) or (inputs(127));
    layer0_outputs(1260) <= (inputs(248)) xor (inputs(64));
    layer0_outputs(1261) <= not(inputs(24)) or (inputs(71));
    layer0_outputs(1262) <= (inputs(221)) and not (inputs(81));
    layer0_outputs(1263) <= not((inputs(31)) or (inputs(71)));
    layer0_outputs(1264) <= (inputs(25)) and not (inputs(165));
    layer0_outputs(1265) <= not((inputs(35)) or (inputs(64)));
    layer0_outputs(1266) <= inputs(141);
    layer0_outputs(1267) <= not((inputs(184)) or (inputs(181)));
    layer0_outputs(1268) <= not((inputs(238)) or (inputs(225)));
    layer0_outputs(1269) <= (inputs(158)) and not (inputs(240));
    layer0_outputs(1270) <= '0';
    layer0_outputs(1271) <= (inputs(255)) or (inputs(70));
    layer0_outputs(1272) <= (inputs(194)) or (inputs(207));
    layer0_outputs(1273) <= (inputs(30)) and not (inputs(43));
    layer0_outputs(1274) <= (inputs(171)) and not (inputs(106));
    layer0_outputs(1275) <= inputs(104);
    layer0_outputs(1276) <= not(inputs(60)) or (inputs(180));
    layer0_outputs(1277) <= inputs(186);
    layer0_outputs(1278) <= (inputs(49)) or (inputs(220));
    layer0_outputs(1279) <= inputs(155);
    layer0_outputs(1280) <= (inputs(226)) or (inputs(40));
    layer0_outputs(1281) <= (inputs(156)) and not (inputs(156));
    layer0_outputs(1282) <= not((inputs(193)) or (inputs(251)));
    layer0_outputs(1283) <= not(inputs(203));
    layer0_outputs(1284) <= (inputs(168)) and (inputs(229));
    layer0_outputs(1285) <= not((inputs(156)) xor (inputs(125)));
    layer0_outputs(1286) <= not(inputs(196));
    layer0_outputs(1287) <= (inputs(45)) and not (inputs(216));
    layer0_outputs(1288) <= not((inputs(104)) or (inputs(198)));
    layer0_outputs(1289) <= not((inputs(147)) or (inputs(133)));
    layer0_outputs(1290) <= inputs(99);
    layer0_outputs(1291) <= not((inputs(145)) and (inputs(152)));
    layer0_outputs(1292) <= not((inputs(95)) or (inputs(137)));
    layer0_outputs(1293) <= not(inputs(233));
    layer0_outputs(1294) <= inputs(98);
    layer0_outputs(1295) <= inputs(44);
    layer0_outputs(1296) <= (inputs(76)) or (inputs(150));
    layer0_outputs(1297) <= not((inputs(30)) or (inputs(62)));
    layer0_outputs(1298) <= inputs(164);
    layer0_outputs(1299) <= inputs(136);
    layer0_outputs(1300) <= inputs(175);
    layer0_outputs(1301) <= (inputs(172)) or (inputs(164));
    layer0_outputs(1302) <= not(inputs(221));
    layer0_outputs(1303) <= inputs(3);
    layer0_outputs(1304) <= inputs(148);
    layer0_outputs(1305) <= not((inputs(133)) or (inputs(104)));
    layer0_outputs(1306) <= inputs(82);
    layer0_outputs(1307) <= not(inputs(122));
    layer0_outputs(1308) <= not((inputs(55)) or (inputs(190)));
    layer0_outputs(1309) <= (inputs(16)) or (inputs(34));
    layer0_outputs(1310) <= not(inputs(25)) or (inputs(163));
    layer0_outputs(1311) <= inputs(31);
    layer0_outputs(1312) <= (inputs(59)) or (inputs(98));
    layer0_outputs(1313) <= not(inputs(61));
    layer0_outputs(1314) <= not((inputs(34)) or (inputs(51)));
    layer0_outputs(1315) <= (inputs(176)) and not (inputs(34));
    layer0_outputs(1316) <= (inputs(55)) and not (inputs(109));
    layer0_outputs(1317) <= not(inputs(106)) or (inputs(144));
    layer0_outputs(1318) <= not(inputs(166));
    layer0_outputs(1319) <= inputs(153);
    layer0_outputs(1320) <= (inputs(23)) xor (inputs(192));
    layer0_outputs(1321) <= not(inputs(106));
    layer0_outputs(1322) <= inputs(234);
    layer0_outputs(1323) <= not((inputs(255)) or (inputs(219)));
    layer0_outputs(1324) <= (inputs(132)) or (inputs(148));
    layer0_outputs(1325) <= not(inputs(181)) or (inputs(94));
    layer0_outputs(1326) <= (inputs(186)) or (inputs(68));
    layer0_outputs(1327) <= not(inputs(134));
    layer0_outputs(1328) <= (inputs(69)) or (inputs(122));
    layer0_outputs(1329) <= not((inputs(18)) or (inputs(128)));
    layer0_outputs(1330) <= not(inputs(199)) or (inputs(175));
    layer0_outputs(1331) <= '0';
    layer0_outputs(1332) <= (inputs(50)) or (inputs(228));
    layer0_outputs(1333) <= not((inputs(203)) or (inputs(159)));
    layer0_outputs(1334) <= not((inputs(97)) and (inputs(77)));
    layer0_outputs(1335) <= inputs(92);
    layer0_outputs(1336) <= (inputs(114)) and (inputs(151));
    layer0_outputs(1337) <= (inputs(93)) or (inputs(79));
    layer0_outputs(1338) <= not(inputs(197));
    layer0_outputs(1339) <= not((inputs(172)) and (inputs(121)));
    layer0_outputs(1340) <= (inputs(174)) or (inputs(27));
    layer0_outputs(1341) <= '1';
    layer0_outputs(1342) <= not(inputs(76)) or (inputs(4));
    layer0_outputs(1343) <= not(inputs(26));
    layer0_outputs(1344) <= not(inputs(91)) or (inputs(5));
    layer0_outputs(1345) <= not(inputs(92)) or (inputs(76));
    layer0_outputs(1346) <= not((inputs(123)) or (inputs(65)));
    layer0_outputs(1347) <= inputs(55);
    layer0_outputs(1348) <= not((inputs(163)) or (inputs(56)));
    layer0_outputs(1349) <= (inputs(232)) and not (inputs(30));
    layer0_outputs(1350) <= not((inputs(1)) xor (inputs(36)));
    layer0_outputs(1351) <= (inputs(208)) and not (inputs(127));
    layer0_outputs(1352) <= not((inputs(145)) or (inputs(178)));
    layer0_outputs(1353) <= not(inputs(166));
    layer0_outputs(1354) <= not((inputs(35)) or (inputs(227)));
    layer0_outputs(1355) <= inputs(9);
    layer0_outputs(1356) <= not((inputs(89)) or (inputs(77)));
    layer0_outputs(1357) <= not(inputs(163));
    layer0_outputs(1358) <= '0';
    layer0_outputs(1359) <= inputs(106);
    layer0_outputs(1360) <= inputs(99);
    layer0_outputs(1361) <= inputs(60);
    layer0_outputs(1362) <= not(inputs(235));
    layer0_outputs(1363) <= not(inputs(104));
    layer0_outputs(1364) <= inputs(193);
    layer0_outputs(1365) <= not((inputs(192)) or (inputs(248)));
    layer0_outputs(1366) <= inputs(203);
    layer0_outputs(1367) <= inputs(238);
    layer0_outputs(1368) <= not((inputs(18)) or (inputs(136)));
    layer0_outputs(1369) <= (inputs(86)) and not (inputs(0));
    layer0_outputs(1370) <= not(inputs(8));
    layer0_outputs(1371) <= not((inputs(215)) xor (inputs(57)));
    layer0_outputs(1372) <= inputs(65);
    layer0_outputs(1373) <= not((inputs(166)) or (inputs(114)));
    layer0_outputs(1374) <= inputs(101);
    layer0_outputs(1375) <= not((inputs(117)) and (inputs(125)));
    layer0_outputs(1376) <= inputs(164);
    layer0_outputs(1377) <= (inputs(161)) or (inputs(179));
    layer0_outputs(1378) <= inputs(205);
    layer0_outputs(1379) <= not(inputs(36)) or (inputs(198));
    layer0_outputs(1380) <= not(inputs(79)) or (inputs(142));
    layer0_outputs(1381) <= not((inputs(235)) or (inputs(177)));
    layer0_outputs(1382) <= '1';
    layer0_outputs(1383) <= (inputs(43)) and not (inputs(8));
    layer0_outputs(1384) <= (inputs(75)) or (inputs(159));
    layer0_outputs(1385) <= (inputs(3)) or (inputs(89));
    layer0_outputs(1386) <= (inputs(150)) or (inputs(219));
    layer0_outputs(1387) <= inputs(81);
    layer0_outputs(1388) <= not((inputs(159)) or (inputs(158)));
    layer0_outputs(1389) <= inputs(219);
    layer0_outputs(1390) <= not(inputs(101));
    layer0_outputs(1391) <= (inputs(161)) or (inputs(171));
    layer0_outputs(1392) <= (inputs(162)) and not (inputs(168));
    layer0_outputs(1393) <= not(inputs(104)) or (inputs(2));
    layer0_outputs(1394) <= not((inputs(150)) or (inputs(144)));
    layer0_outputs(1395) <= (inputs(152)) and not (inputs(115));
    layer0_outputs(1396) <= not((inputs(156)) or (inputs(98)));
    layer0_outputs(1397) <= inputs(105);
    layer0_outputs(1398) <= not(inputs(234));
    layer0_outputs(1399) <= (inputs(175)) or (inputs(230));
    layer0_outputs(1400) <= not((inputs(253)) or (inputs(21)));
    layer0_outputs(1401) <= not(inputs(9));
    layer0_outputs(1402) <= not(inputs(46));
    layer0_outputs(1403) <= not((inputs(171)) or (inputs(141)));
    layer0_outputs(1404) <= not(inputs(119));
    layer0_outputs(1405) <= not(inputs(199)) or (inputs(93));
    layer0_outputs(1406) <= not(inputs(179));
    layer0_outputs(1407) <= not((inputs(7)) xor (inputs(55)));
    layer0_outputs(1408) <= (inputs(253)) or (inputs(207));
    layer0_outputs(1409) <= not((inputs(239)) or (inputs(135)));
    layer0_outputs(1410) <= inputs(120);
    layer0_outputs(1411) <= not(inputs(110));
    layer0_outputs(1412) <= not((inputs(167)) or (inputs(4)));
    layer0_outputs(1413) <= (inputs(107)) or (inputs(82));
    layer0_outputs(1414) <= inputs(253);
    layer0_outputs(1415) <= not((inputs(29)) or (inputs(219)));
    layer0_outputs(1416) <= inputs(47);
    layer0_outputs(1417) <= (inputs(243)) and not (inputs(145));
    layer0_outputs(1418) <= not(inputs(96)) or (inputs(81));
    layer0_outputs(1419) <= not((inputs(32)) or (inputs(252)));
    layer0_outputs(1420) <= inputs(75);
    layer0_outputs(1421) <= not((inputs(16)) or (inputs(156)));
    layer0_outputs(1422) <= not(inputs(244)) or (inputs(50));
    layer0_outputs(1423) <= inputs(114);
    layer0_outputs(1424) <= inputs(236);
    layer0_outputs(1425) <= not(inputs(78));
    layer0_outputs(1426) <= not(inputs(54));
    layer0_outputs(1427) <= not((inputs(13)) and (inputs(232)));
    layer0_outputs(1428) <= not(inputs(172));
    layer0_outputs(1429) <= (inputs(34)) or (inputs(23));
    layer0_outputs(1430) <= (inputs(41)) and not (inputs(15));
    layer0_outputs(1431) <= (inputs(26)) and not (inputs(88));
    layer0_outputs(1432) <= (inputs(192)) or (inputs(194));
    layer0_outputs(1433) <= not(inputs(111));
    layer0_outputs(1434) <= not(inputs(42));
    layer0_outputs(1435) <= '1';
    layer0_outputs(1436) <= not((inputs(198)) or (inputs(127)));
    layer0_outputs(1437) <= inputs(177);
    layer0_outputs(1438) <= not((inputs(73)) or (inputs(170)));
    layer0_outputs(1439) <= not(inputs(165));
    layer0_outputs(1440) <= (inputs(111)) or (inputs(7));
    layer0_outputs(1441) <= inputs(78);
    layer0_outputs(1442) <= not(inputs(250)) or (inputs(0));
    layer0_outputs(1443) <= not(inputs(177));
    layer0_outputs(1444) <= not(inputs(248));
    layer0_outputs(1445) <= not(inputs(139));
    layer0_outputs(1446) <= not(inputs(185));
    layer0_outputs(1447) <= inputs(193);
    layer0_outputs(1448) <= not(inputs(4));
    layer0_outputs(1449) <= inputs(164);
    layer0_outputs(1450) <= not((inputs(137)) and (inputs(89)));
    layer0_outputs(1451) <= not((inputs(161)) or (inputs(6)));
    layer0_outputs(1452) <= inputs(120);
    layer0_outputs(1453) <= (inputs(220)) and not (inputs(238));
    layer0_outputs(1454) <= not(inputs(130)) or (inputs(239));
    layer0_outputs(1455) <= not(inputs(139)) or (inputs(196));
    layer0_outputs(1456) <= inputs(152);
    layer0_outputs(1457) <= (inputs(121)) xor (inputs(94));
    layer0_outputs(1458) <= (inputs(87)) or (inputs(116));
    layer0_outputs(1459) <= inputs(90);
    layer0_outputs(1460) <= (inputs(162)) and not (inputs(178));
    layer0_outputs(1461) <= not((inputs(20)) or (inputs(48)));
    layer0_outputs(1462) <= inputs(225);
    layer0_outputs(1463) <= (inputs(24)) and (inputs(74));
    layer0_outputs(1464) <= not((inputs(80)) or (inputs(162)));
    layer0_outputs(1465) <= inputs(24);
    layer0_outputs(1466) <= not(inputs(61));
    layer0_outputs(1467) <= not((inputs(128)) or (inputs(160)));
    layer0_outputs(1468) <= not((inputs(39)) or (inputs(192)));
    layer0_outputs(1469) <= (inputs(17)) and not (inputs(229));
    layer0_outputs(1470) <= inputs(188);
    layer0_outputs(1471) <= not((inputs(158)) or (inputs(111)));
    layer0_outputs(1472) <= not(inputs(84));
    layer0_outputs(1473) <= not((inputs(143)) or (inputs(81)));
    layer0_outputs(1474) <= not((inputs(144)) xor (inputs(136)));
    layer0_outputs(1475) <= inputs(81);
    layer0_outputs(1476) <= (inputs(167)) and not (inputs(68));
    layer0_outputs(1477) <= not((inputs(210)) and (inputs(63)));
    layer0_outputs(1478) <= (inputs(126)) or (inputs(127));
    layer0_outputs(1479) <= not(inputs(181));
    layer0_outputs(1480) <= not(inputs(184));
    layer0_outputs(1481) <= '0';
    layer0_outputs(1482) <= not(inputs(156));
    layer0_outputs(1483) <= not(inputs(230));
    layer0_outputs(1484) <= (inputs(141)) or (inputs(16));
    layer0_outputs(1485) <= (inputs(114)) or (inputs(189));
    layer0_outputs(1486) <= not((inputs(240)) or (inputs(9)));
    layer0_outputs(1487) <= inputs(135);
    layer0_outputs(1488) <= inputs(154);
    layer0_outputs(1489) <= not(inputs(167)) or (inputs(30));
    layer0_outputs(1490) <= (inputs(73)) and not (inputs(5));
    layer0_outputs(1491) <= not(inputs(116));
    layer0_outputs(1492) <= (inputs(158)) or (inputs(2));
    layer0_outputs(1493) <= (inputs(163)) or (inputs(71));
    layer0_outputs(1494) <= (inputs(157)) and not (inputs(252));
    layer0_outputs(1495) <= not(inputs(53));
    layer0_outputs(1496) <= not(inputs(13)) or (inputs(204));
    layer0_outputs(1497) <= not(inputs(246)) or (inputs(149));
    layer0_outputs(1498) <= (inputs(156)) and not (inputs(65));
    layer0_outputs(1499) <= not(inputs(41)) or (inputs(225));
    layer0_outputs(1500) <= not(inputs(88));
    layer0_outputs(1501) <= not((inputs(23)) xor (inputs(155)));
    layer0_outputs(1502) <= '0';
    layer0_outputs(1503) <= not((inputs(8)) or (inputs(238)));
    layer0_outputs(1504) <= '1';
    layer0_outputs(1505) <= (inputs(170)) or (inputs(32));
    layer0_outputs(1506) <= (inputs(140)) or (inputs(125));
    layer0_outputs(1507) <= inputs(121);
    layer0_outputs(1508) <= inputs(132);
    layer0_outputs(1509) <= inputs(178);
    layer0_outputs(1510) <= not(inputs(136));
    layer0_outputs(1511) <= inputs(237);
    layer0_outputs(1512) <= not(inputs(56));
    layer0_outputs(1513) <= inputs(71);
    layer0_outputs(1514) <= not(inputs(68));
    layer0_outputs(1515) <= not((inputs(233)) and (inputs(23)));
    layer0_outputs(1516) <= (inputs(185)) or (inputs(111));
    layer0_outputs(1517) <= (inputs(144)) or (inputs(172));
    layer0_outputs(1518) <= not(inputs(248));
    layer0_outputs(1519) <= not(inputs(180));
    layer0_outputs(1520) <= (inputs(167)) xor (inputs(255));
    layer0_outputs(1521) <= not(inputs(162));
    layer0_outputs(1522) <= not(inputs(97)) or (inputs(95));
    layer0_outputs(1523) <= not(inputs(112));
    layer0_outputs(1524) <= not((inputs(114)) or (inputs(181)));
    layer0_outputs(1525) <= inputs(162);
    layer0_outputs(1526) <= not(inputs(194));
    layer0_outputs(1527) <= (inputs(145)) and (inputs(58));
    layer0_outputs(1528) <= not(inputs(87)) or (inputs(205));
    layer0_outputs(1529) <= (inputs(92)) xor (inputs(142));
    layer0_outputs(1530) <= not(inputs(177)) or (inputs(141));
    layer0_outputs(1531) <= inputs(37);
    layer0_outputs(1532) <= not((inputs(17)) or (inputs(190)));
    layer0_outputs(1533) <= not(inputs(127)) or (inputs(64));
    layer0_outputs(1534) <= inputs(205);
    layer0_outputs(1535) <= '1';
    layer0_outputs(1536) <= inputs(248);
    layer0_outputs(1537) <= not(inputs(120));
    layer0_outputs(1538) <= inputs(166);
    layer0_outputs(1539) <= not(inputs(148));
    layer0_outputs(1540) <= inputs(205);
    layer0_outputs(1541) <= not(inputs(38)) or (inputs(193));
    layer0_outputs(1542) <= not(inputs(123));
    layer0_outputs(1543) <= not(inputs(44));
    layer0_outputs(1544) <= not(inputs(20));
    layer0_outputs(1545) <= inputs(9);
    layer0_outputs(1546) <= '1';
    layer0_outputs(1547) <= (inputs(224)) or (inputs(102));
    layer0_outputs(1548) <= '1';
    layer0_outputs(1549) <= not((inputs(195)) or (inputs(33)));
    layer0_outputs(1550) <= not(inputs(56));
    layer0_outputs(1551) <= (inputs(79)) or (inputs(28));
    layer0_outputs(1552) <= inputs(34);
    layer0_outputs(1553) <= (inputs(212)) and not (inputs(93));
    layer0_outputs(1554) <= not(inputs(209));
    layer0_outputs(1555) <= not(inputs(86));
    layer0_outputs(1556) <= not(inputs(202));
    layer0_outputs(1557) <= (inputs(118)) or (inputs(116));
    layer0_outputs(1558) <= inputs(149);
    layer0_outputs(1559) <= (inputs(232)) and not (inputs(0));
    layer0_outputs(1560) <= (inputs(72)) xor (inputs(146));
    layer0_outputs(1561) <= not(inputs(21)) or (inputs(175));
    layer0_outputs(1562) <= inputs(165);
    layer0_outputs(1563) <= not((inputs(209)) or (inputs(216)));
    layer0_outputs(1564) <= (inputs(212)) and not (inputs(141));
    layer0_outputs(1565) <= not((inputs(133)) or (inputs(173)));
    layer0_outputs(1566) <= not(inputs(175));
    layer0_outputs(1567) <= not(inputs(226));
    layer0_outputs(1568) <= not((inputs(219)) xor (inputs(155)));
    layer0_outputs(1569) <= (inputs(23)) and not (inputs(157));
    layer0_outputs(1570) <= inputs(149);
    layer0_outputs(1571) <= inputs(135);
    layer0_outputs(1572) <= (inputs(33)) or (inputs(5));
    layer0_outputs(1573) <= not(inputs(167));
    layer0_outputs(1574) <= not(inputs(89));
    layer0_outputs(1575) <= inputs(123);
    layer0_outputs(1576) <= '1';
    layer0_outputs(1577) <= not(inputs(234));
    layer0_outputs(1578) <= not(inputs(5));
    layer0_outputs(1579) <= not(inputs(125));
    layer0_outputs(1580) <= not((inputs(242)) or (inputs(113)));
    layer0_outputs(1581) <= (inputs(143)) and (inputs(158));
    layer0_outputs(1582) <= inputs(41);
    layer0_outputs(1583) <= not((inputs(133)) or (inputs(96)));
    layer0_outputs(1584) <= not(inputs(174));
    layer0_outputs(1585) <= not(inputs(162));
    layer0_outputs(1586) <= not((inputs(220)) and (inputs(84)));
    layer0_outputs(1587) <= not(inputs(11));
    layer0_outputs(1588) <= not((inputs(129)) or (inputs(182)));
    layer0_outputs(1589) <= not(inputs(119)) or (inputs(179));
    layer0_outputs(1590) <= not((inputs(235)) xor (inputs(26)));
    layer0_outputs(1591) <= (inputs(52)) or (inputs(24));
    layer0_outputs(1592) <= (inputs(202)) and not (inputs(246));
    layer0_outputs(1593) <= inputs(102);
    layer0_outputs(1594) <= not(inputs(193)) or (inputs(13));
    layer0_outputs(1595) <= (inputs(65)) and not (inputs(120));
    layer0_outputs(1596) <= not(inputs(206));
    layer0_outputs(1597) <= inputs(168);
    layer0_outputs(1598) <= not(inputs(163));
    layer0_outputs(1599) <= (inputs(74)) and not (inputs(155));
    layer0_outputs(1600) <= inputs(70);
    layer0_outputs(1601) <= not((inputs(50)) or (inputs(180)));
    layer0_outputs(1602) <= inputs(29);
    layer0_outputs(1603) <= inputs(167);
    layer0_outputs(1604) <= not(inputs(46));
    layer0_outputs(1605) <= (inputs(152)) and not (inputs(154));
    layer0_outputs(1606) <= inputs(22);
    layer0_outputs(1607) <= (inputs(233)) or (inputs(21));
    layer0_outputs(1608) <= not(inputs(248));
    layer0_outputs(1609) <= inputs(31);
    layer0_outputs(1610) <= not(inputs(251)) or (inputs(128));
    layer0_outputs(1611) <= not((inputs(68)) or (inputs(82)));
    layer0_outputs(1612) <= not(inputs(7)) or (inputs(27));
    layer0_outputs(1613) <= not((inputs(119)) or (inputs(46)));
    layer0_outputs(1614) <= inputs(26);
    layer0_outputs(1615) <= inputs(179);
    layer0_outputs(1616) <= (inputs(78)) or (inputs(210));
    layer0_outputs(1617) <= (inputs(184)) or (inputs(167));
    layer0_outputs(1618) <= not(inputs(152));
    layer0_outputs(1619) <= not((inputs(54)) xor (inputs(5)));
    layer0_outputs(1620) <= (inputs(85)) and not (inputs(183));
    layer0_outputs(1621) <= inputs(67);
    layer0_outputs(1622) <= not(inputs(194)) or (inputs(222));
    layer0_outputs(1623) <= inputs(26);
    layer0_outputs(1624) <= (inputs(92)) and not (inputs(226));
    layer0_outputs(1625) <= inputs(61);
    layer0_outputs(1626) <= (inputs(164)) or (inputs(112));
    layer0_outputs(1627) <= (inputs(212)) or (inputs(211));
    layer0_outputs(1628) <= (inputs(28)) and not (inputs(223));
    layer0_outputs(1629) <= not(inputs(210));
    layer0_outputs(1630) <= not((inputs(234)) or (inputs(225)));
    layer0_outputs(1631) <= not(inputs(181));
    layer0_outputs(1632) <= (inputs(90)) or (inputs(252));
    layer0_outputs(1633) <= (inputs(95)) or (inputs(29));
    layer0_outputs(1634) <= inputs(134);
    layer0_outputs(1635) <= not(inputs(131)) or (inputs(2));
    layer0_outputs(1636) <= not(inputs(53));
    layer0_outputs(1637) <= (inputs(107)) or (inputs(35));
    layer0_outputs(1638) <= inputs(149);
    layer0_outputs(1639) <= inputs(66);
    layer0_outputs(1640) <= not((inputs(94)) or (inputs(57)));
    layer0_outputs(1641) <= (inputs(172)) and not (inputs(167));
    layer0_outputs(1642) <= inputs(146);
    layer0_outputs(1643) <= not(inputs(40));
    layer0_outputs(1644) <= (inputs(211)) and not (inputs(119));
    layer0_outputs(1645) <= not(inputs(236));
    layer0_outputs(1646) <= (inputs(246)) and not (inputs(138));
    layer0_outputs(1647) <= inputs(223);
    layer0_outputs(1648) <= not((inputs(176)) or (inputs(1)));
    layer0_outputs(1649) <= not((inputs(193)) or (inputs(108)));
    layer0_outputs(1650) <= inputs(43);
    layer0_outputs(1651) <= not(inputs(131));
    layer0_outputs(1652) <= not((inputs(178)) or (inputs(154)));
    layer0_outputs(1653) <= (inputs(226)) or (inputs(65));
    layer0_outputs(1654) <= inputs(9);
    layer0_outputs(1655) <= not(inputs(35)) or (inputs(113));
    layer0_outputs(1656) <= not((inputs(221)) xor (inputs(251)));
    layer0_outputs(1657) <= not(inputs(105)) or (inputs(211));
    layer0_outputs(1658) <= (inputs(229)) and (inputs(62));
    layer0_outputs(1659) <= not(inputs(108)) or (inputs(199));
    layer0_outputs(1660) <= (inputs(213)) or (inputs(235));
    layer0_outputs(1661) <= (inputs(236)) and not (inputs(12));
    layer0_outputs(1662) <= not(inputs(75));
    layer0_outputs(1663) <= not(inputs(233));
    layer0_outputs(1664) <= not(inputs(102)) or (inputs(239));
    layer0_outputs(1665) <= not((inputs(85)) or (inputs(162)));
    layer0_outputs(1666) <= (inputs(129)) or (inputs(153));
    layer0_outputs(1667) <= (inputs(124)) or (inputs(83));
    layer0_outputs(1668) <= not(inputs(173)) or (inputs(182));
    layer0_outputs(1669) <= inputs(138);
    layer0_outputs(1670) <= inputs(68);
    layer0_outputs(1671) <= (inputs(19)) xor (inputs(93));
    layer0_outputs(1672) <= not((inputs(76)) or (inputs(121)));
    layer0_outputs(1673) <= inputs(233);
    layer0_outputs(1674) <= (inputs(221)) xor (inputs(17));
    layer0_outputs(1675) <= not(inputs(146));
    layer0_outputs(1676) <= '1';
    layer0_outputs(1677) <= inputs(94);
    layer0_outputs(1678) <= (inputs(95)) or (inputs(253));
    layer0_outputs(1679) <= (inputs(250)) or (inputs(131));
    layer0_outputs(1680) <= inputs(2);
    layer0_outputs(1681) <= not((inputs(167)) or (inputs(123)));
    layer0_outputs(1682) <= not(inputs(82));
    layer0_outputs(1683) <= not((inputs(74)) or (inputs(62)));
    layer0_outputs(1684) <= (inputs(127)) xor (inputs(156));
    layer0_outputs(1685) <= not(inputs(223));
    layer0_outputs(1686) <= inputs(125);
    layer0_outputs(1687) <= inputs(126);
    layer0_outputs(1688) <= '1';
    layer0_outputs(1689) <= inputs(115);
    layer0_outputs(1690) <= not((inputs(128)) or (inputs(65)));
    layer0_outputs(1691) <= inputs(117);
    layer0_outputs(1692) <= not((inputs(174)) or (inputs(17)));
    layer0_outputs(1693) <= not((inputs(4)) or (inputs(33)));
    layer0_outputs(1694) <= (inputs(31)) and not (inputs(95));
    layer0_outputs(1695) <= not((inputs(144)) or (inputs(82)));
    layer0_outputs(1696) <= not((inputs(92)) or (inputs(100)));
    layer0_outputs(1697) <= (inputs(250)) or (inputs(134));
    layer0_outputs(1698) <= inputs(37);
    layer0_outputs(1699) <= inputs(203);
    layer0_outputs(1700) <= (inputs(193)) or (inputs(242));
    layer0_outputs(1701) <= not(inputs(116)) or (inputs(2));
    layer0_outputs(1702) <= not(inputs(161));
    layer0_outputs(1703) <= inputs(18);
    layer0_outputs(1704) <= not(inputs(57));
    layer0_outputs(1705) <= not((inputs(15)) or (inputs(196)));
    layer0_outputs(1706) <= not(inputs(91));
    layer0_outputs(1707) <= not(inputs(123));
    layer0_outputs(1708) <= not(inputs(230));
    layer0_outputs(1709) <= not(inputs(102));
    layer0_outputs(1710) <= inputs(215);
    layer0_outputs(1711) <= (inputs(90)) or (inputs(245));
    layer0_outputs(1712) <= (inputs(8)) and not (inputs(165));
    layer0_outputs(1713) <= not(inputs(95));
    layer0_outputs(1714) <= (inputs(174)) or (inputs(147));
    layer0_outputs(1715) <= (inputs(161)) or (inputs(166));
    layer0_outputs(1716) <= '0';
    layer0_outputs(1717) <= (inputs(214)) or (inputs(232));
    layer0_outputs(1718) <= (inputs(28)) or (inputs(242));
    layer0_outputs(1719) <= (inputs(234)) or (inputs(31));
    layer0_outputs(1720) <= not(inputs(224));
    layer0_outputs(1721) <= not(inputs(108)) or (inputs(193));
    layer0_outputs(1722) <= not(inputs(14));
    layer0_outputs(1723) <= (inputs(64)) or (inputs(21));
    layer0_outputs(1724) <= not(inputs(247));
    layer0_outputs(1725) <= not(inputs(92));
    layer0_outputs(1726) <= (inputs(181)) and not (inputs(17));
    layer0_outputs(1727) <= not(inputs(143));
    layer0_outputs(1728) <= not((inputs(80)) or (inputs(78)));
    layer0_outputs(1729) <= inputs(60);
    layer0_outputs(1730) <= not((inputs(87)) or (inputs(119)));
    layer0_outputs(1731) <= '1';
    layer0_outputs(1732) <= (inputs(95)) or (inputs(170));
    layer0_outputs(1733) <= (inputs(186)) or (inputs(43));
    layer0_outputs(1734) <= (inputs(178)) xor (inputs(160));
    layer0_outputs(1735) <= (inputs(132)) or (inputs(101));
    layer0_outputs(1736) <= inputs(202);
    layer0_outputs(1737) <= (inputs(37)) and not (inputs(207));
    layer0_outputs(1738) <= not((inputs(245)) or (inputs(113)));
    layer0_outputs(1739) <= inputs(173);
    layer0_outputs(1740) <= inputs(195);
    layer0_outputs(1741) <= inputs(58);
    layer0_outputs(1742) <= (inputs(163)) or (inputs(146));
    layer0_outputs(1743) <= not((inputs(52)) or (inputs(112)));
    layer0_outputs(1744) <= inputs(76);
    layer0_outputs(1745) <= not((inputs(169)) or (inputs(201)));
    layer0_outputs(1746) <= (inputs(138)) and not (inputs(39));
    layer0_outputs(1747) <= inputs(38);
    layer0_outputs(1748) <= inputs(67);
    layer0_outputs(1749) <= inputs(131);
    layer0_outputs(1750) <= (inputs(133)) and not (inputs(191));
    layer0_outputs(1751) <= (inputs(37)) or (inputs(67));
    layer0_outputs(1752) <= (inputs(112)) or (inputs(66));
    layer0_outputs(1753) <= not(inputs(120)) or (inputs(34));
    layer0_outputs(1754) <= inputs(85);
    layer0_outputs(1755) <= (inputs(85)) or (inputs(81));
    layer0_outputs(1756) <= not(inputs(131));
    layer0_outputs(1757) <= not(inputs(107)) or (inputs(194));
    layer0_outputs(1758) <= not((inputs(45)) or (inputs(28)));
    layer0_outputs(1759) <= (inputs(38)) and not (inputs(162));
    layer0_outputs(1760) <= (inputs(137)) and not (inputs(161));
    layer0_outputs(1761) <= inputs(230);
    layer0_outputs(1762) <= not(inputs(173)) or (inputs(14));
    layer0_outputs(1763) <= not((inputs(128)) or (inputs(171)));
    layer0_outputs(1764) <= not(inputs(1));
    layer0_outputs(1765) <= not((inputs(183)) or (inputs(238)));
    layer0_outputs(1766) <= not((inputs(2)) or (inputs(42)));
    layer0_outputs(1767) <= not((inputs(24)) or (inputs(219)));
    layer0_outputs(1768) <= not(inputs(254));
    layer0_outputs(1769) <= not(inputs(120)) or (inputs(113));
    layer0_outputs(1770) <= (inputs(120)) and not (inputs(178));
    layer0_outputs(1771) <= not(inputs(29));
    layer0_outputs(1772) <= not(inputs(149)) or (inputs(114));
    layer0_outputs(1773) <= inputs(208);
    layer0_outputs(1774) <= not((inputs(247)) or (inputs(56)));
    layer0_outputs(1775) <= (inputs(83)) or (inputs(113));
    layer0_outputs(1776) <= inputs(28);
    layer0_outputs(1777) <= not(inputs(179)) or (inputs(128));
    layer0_outputs(1778) <= (inputs(34)) or (inputs(208));
    layer0_outputs(1779) <= inputs(79);
    layer0_outputs(1780) <= not((inputs(255)) or (inputs(189)));
    layer0_outputs(1781) <= not(inputs(26));
    layer0_outputs(1782) <= not(inputs(102));
    layer0_outputs(1783) <= not(inputs(29));
    layer0_outputs(1784) <= (inputs(238)) or (inputs(200));
    layer0_outputs(1785) <= (inputs(96)) and (inputs(41));
    layer0_outputs(1786) <= (inputs(203)) xor (inputs(207));
    layer0_outputs(1787) <= not(inputs(247)) or (inputs(75));
    layer0_outputs(1788) <= (inputs(35)) or (inputs(224));
    layer0_outputs(1789) <= not(inputs(166));
    layer0_outputs(1790) <= inputs(155);
    layer0_outputs(1791) <= not(inputs(178)) or (inputs(238));
    layer0_outputs(1792) <= not(inputs(19));
    layer0_outputs(1793) <= not(inputs(182));
    layer0_outputs(1794) <= not((inputs(246)) or (inputs(137)));
    layer0_outputs(1795) <= inputs(227);
    layer0_outputs(1796) <= (inputs(52)) and not (inputs(113));
    layer0_outputs(1797) <= (inputs(117)) or (inputs(213));
    layer0_outputs(1798) <= not((inputs(76)) or (inputs(32)));
    layer0_outputs(1799) <= not(inputs(70));
    layer0_outputs(1800) <= (inputs(13)) and not (inputs(111));
    layer0_outputs(1801) <= not(inputs(99));
    layer0_outputs(1802) <= '1';
    layer0_outputs(1803) <= not(inputs(232));
    layer0_outputs(1804) <= not(inputs(129));
    layer0_outputs(1805) <= not(inputs(83));
    layer0_outputs(1806) <= (inputs(77)) and not (inputs(45));
    layer0_outputs(1807) <= not(inputs(247));
    layer0_outputs(1808) <= '1';
    layer0_outputs(1809) <= not((inputs(64)) or (inputs(92)));
    layer0_outputs(1810) <= inputs(165);
    layer0_outputs(1811) <= not(inputs(249));
    layer0_outputs(1812) <= (inputs(182)) and not (inputs(108));
    layer0_outputs(1813) <= inputs(179);
    layer0_outputs(1814) <= (inputs(223)) xor (inputs(186));
    layer0_outputs(1815) <= not(inputs(211)) or (inputs(11));
    layer0_outputs(1816) <= (inputs(219)) or (inputs(179));
    layer0_outputs(1817) <= not(inputs(131)) or (inputs(70));
    layer0_outputs(1818) <= (inputs(179)) and not (inputs(253));
    layer0_outputs(1819) <= not(inputs(126));
    layer0_outputs(1820) <= not(inputs(20)) or (inputs(239));
    layer0_outputs(1821) <= (inputs(121)) and not (inputs(176));
    layer0_outputs(1822) <= (inputs(84)) or (inputs(76));
    layer0_outputs(1823) <= '1';
    layer0_outputs(1824) <= inputs(73);
    layer0_outputs(1825) <= not(inputs(74));
    layer0_outputs(1826) <= not(inputs(85));
    layer0_outputs(1827) <= (inputs(105)) xor (inputs(182));
    layer0_outputs(1828) <= not(inputs(214)) or (inputs(60));
    layer0_outputs(1829) <= not((inputs(247)) or (inputs(130)));
    layer0_outputs(1830) <= not((inputs(128)) or (inputs(189)));
    layer0_outputs(1831) <= '1';
    layer0_outputs(1832) <= not(inputs(53)) or (inputs(146));
    layer0_outputs(1833) <= not((inputs(1)) xor (inputs(171)));
    layer0_outputs(1834) <= (inputs(10)) and not (inputs(172));
    layer0_outputs(1835) <= not(inputs(155));
    layer0_outputs(1836) <= not(inputs(230)) or (inputs(184));
    layer0_outputs(1837) <= '1';
    layer0_outputs(1838) <= inputs(69);
    layer0_outputs(1839) <= (inputs(103)) or (inputs(247));
    layer0_outputs(1840) <= (inputs(36)) and not (inputs(128));
    layer0_outputs(1841) <= not(inputs(19));
    layer0_outputs(1842) <= not((inputs(25)) and (inputs(39)));
    layer0_outputs(1843) <= not(inputs(194));
    layer0_outputs(1844) <= inputs(117);
    layer0_outputs(1845) <= not((inputs(248)) or (inputs(29)));
    layer0_outputs(1846) <= not(inputs(56));
    layer0_outputs(1847) <= (inputs(53)) or (inputs(46));
    layer0_outputs(1848) <= not(inputs(143)) or (inputs(253));
    layer0_outputs(1849) <= inputs(181);
    layer0_outputs(1850) <= (inputs(92)) xor (inputs(19));
    layer0_outputs(1851) <= not(inputs(7));
    layer0_outputs(1852) <= (inputs(65)) or (inputs(63));
    layer0_outputs(1853) <= not((inputs(141)) or (inputs(124)));
    layer0_outputs(1854) <= (inputs(152)) and not (inputs(5));
    layer0_outputs(1855) <= inputs(90);
    layer0_outputs(1856) <= (inputs(47)) or (inputs(52));
    layer0_outputs(1857) <= '0';
    layer0_outputs(1858) <= inputs(8);
    layer0_outputs(1859) <= not(inputs(208)) or (inputs(145));
    layer0_outputs(1860) <= '1';
    layer0_outputs(1861) <= not((inputs(62)) xor (inputs(24)));
    layer0_outputs(1862) <= not(inputs(134));
    layer0_outputs(1863) <= not(inputs(192));
    layer0_outputs(1864) <= inputs(115);
    layer0_outputs(1865) <= not(inputs(216)) or (inputs(98));
    layer0_outputs(1866) <= not((inputs(121)) or (inputs(97)));
    layer0_outputs(1867) <= (inputs(90)) or (inputs(80));
    layer0_outputs(1868) <= not(inputs(55)) or (inputs(101));
    layer0_outputs(1869) <= '0';
    layer0_outputs(1870) <= not(inputs(7)) or (inputs(56));
    layer0_outputs(1871) <= (inputs(88)) and not (inputs(48));
    layer0_outputs(1872) <= not(inputs(41));
    layer0_outputs(1873) <= not(inputs(84)) or (inputs(125));
    layer0_outputs(1874) <= not(inputs(25)) or (inputs(193));
    layer0_outputs(1875) <= (inputs(141)) and not (inputs(148));
    layer0_outputs(1876) <= '1';
    layer0_outputs(1877) <= (inputs(135)) and not (inputs(111));
    layer0_outputs(1878) <= not(inputs(88));
    layer0_outputs(1879) <= not((inputs(251)) or (inputs(137)));
    layer0_outputs(1880) <= not(inputs(145));
    layer0_outputs(1881) <= (inputs(195)) or (inputs(31));
    layer0_outputs(1882) <= inputs(28);
    layer0_outputs(1883) <= inputs(178);
    layer0_outputs(1884) <= (inputs(234)) and not (inputs(0));
    layer0_outputs(1885) <= (inputs(88)) and not (inputs(122));
    layer0_outputs(1886) <= (inputs(195)) and not (inputs(253));
    layer0_outputs(1887) <= not(inputs(248)) or (inputs(182));
    layer0_outputs(1888) <= not((inputs(195)) or (inputs(116)));
    layer0_outputs(1889) <= '1';
    layer0_outputs(1890) <= not(inputs(137)) or (inputs(42));
    layer0_outputs(1891) <= not((inputs(19)) or (inputs(31)));
    layer0_outputs(1892) <= not((inputs(146)) or (inputs(165)));
    layer0_outputs(1893) <= (inputs(144)) or (inputs(94));
    layer0_outputs(1894) <= inputs(8);
    layer0_outputs(1895) <= not(inputs(217)) or (inputs(156));
    layer0_outputs(1896) <= inputs(209);
    layer0_outputs(1897) <= (inputs(54)) and not (inputs(249));
    layer0_outputs(1898) <= (inputs(184)) or (inputs(175));
    layer0_outputs(1899) <= '0';
    layer0_outputs(1900) <= '1';
    layer0_outputs(1901) <= not(inputs(104)) or (inputs(112));
    layer0_outputs(1902) <= '1';
    layer0_outputs(1903) <= inputs(232);
    layer0_outputs(1904) <= (inputs(170)) or (inputs(176));
    layer0_outputs(1905) <= not(inputs(164)) or (inputs(5));
    layer0_outputs(1906) <= (inputs(145)) or (inputs(163));
    layer0_outputs(1907) <= not((inputs(89)) and (inputs(167)));
    layer0_outputs(1908) <= inputs(12);
    layer0_outputs(1909) <= (inputs(97)) and (inputs(44));
    layer0_outputs(1910) <= not(inputs(182));
    layer0_outputs(1911) <= (inputs(10)) and not (inputs(96));
    layer0_outputs(1912) <= not(inputs(230));
    layer0_outputs(1913) <= inputs(197);
    layer0_outputs(1914) <= (inputs(48)) or (inputs(94));
    layer0_outputs(1915) <= inputs(205);
    layer0_outputs(1916) <= inputs(155);
    layer0_outputs(1917) <= inputs(135);
    layer0_outputs(1918) <= not(inputs(133));
    layer0_outputs(1919) <= (inputs(65)) or (inputs(48));
    layer0_outputs(1920) <= (inputs(37)) or (inputs(118));
    layer0_outputs(1921) <= (inputs(110)) and not (inputs(224));
    layer0_outputs(1922) <= not(inputs(71)) or (inputs(17));
    layer0_outputs(1923) <= (inputs(153)) and not (inputs(239));
    layer0_outputs(1924) <= not((inputs(157)) and (inputs(111)));
    layer0_outputs(1925) <= (inputs(83)) and not (inputs(3));
    layer0_outputs(1926) <= (inputs(15)) or (inputs(107));
    layer0_outputs(1927) <= (inputs(85)) and not (inputs(221));
    layer0_outputs(1928) <= inputs(170);
    layer0_outputs(1929) <= not(inputs(36)) or (inputs(224));
    layer0_outputs(1930) <= not(inputs(142));
    layer0_outputs(1931) <= not((inputs(146)) or (inputs(59)));
    layer0_outputs(1932) <= (inputs(16)) or (inputs(59));
    layer0_outputs(1933) <= not((inputs(86)) and (inputs(19)));
    layer0_outputs(1934) <= not((inputs(69)) xor (inputs(149)));
    layer0_outputs(1935) <= not((inputs(224)) xor (inputs(232)));
    layer0_outputs(1936) <= not(inputs(202)) or (inputs(139));
    layer0_outputs(1937) <= not((inputs(214)) or (inputs(164)));
    layer0_outputs(1938) <= not((inputs(171)) or (inputs(100)));
    layer0_outputs(1939) <= not(inputs(11)) or (inputs(188));
    layer0_outputs(1940) <= (inputs(227)) and not (inputs(197));
    layer0_outputs(1941) <= not(inputs(202));
    layer0_outputs(1942) <= (inputs(42)) and not (inputs(63));
    layer0_outputs(1943) <= '0';
    layer0_outputs(1944) <= (inputs(0)) xor (inputs(78));
    layer0_outputs(1945) <= (inputs(179)) or (inputs(34));
    layer0_outputs(1946) <= not(inputs(38)) or (inputs(214));
    layer0_outputs(1947) <= (inputs(150)) and not (inputs(121));
    layer0_outputs(1948) <= (inputs(227)) and (inputs(197));
    layer0_outputs(1949) <= not((inputs(247)) or (inputs(91)));
    layer0_outputs(1950) <= not((inputs(80)) or (inputs(210)));
    layer0_outputs(1951) <= inputs(129);
    layer0_outputs(1952) <= not(inputs(74));
    layer0_outputs(1953) <= (inputs(186)) or (inputs(70));
    layer0_outputs(1954) <= not((inputs(97)) or (inputs(248)));
    layer0_outputs(1955) <= not((inputs(147)) or (inputs(109)));
    layer0_outputs(1956) <= (inputs(58)) and not (inputs(82));
    layer0_outputs(1957) <= not(inputs(147));
    layer0_outputs(1958) <= (inputs(11)) and not (inputs(223));
    layer0_outputs(1959) <= not((inputs(0)) xor (inputs(78)));
    layer0_outputs(1960) <= not(inputs(131));
    layer0_outputs(1961) <= (inputs(53)) and not (inputs(241));
    layer0_outputs(1962) <= not(inputs(208));
    layer0_outputs(1963) <= inputs(237);
    layer0_outputs(1964) <= '1';
    layer0_outputs(1965) <= not(inputs(76));
    layer0_outputs(1966) <= not(inputs(152));
    layer0_outputs(1967) <= not(inputs(146)) or (inputs(15));
    layer0_outputs(1968) <= not(inputs(226));
    layer0_outputs(1969) <= not((inputs(174)) or (inputs(43)));
    layer0_outputs(1970) <= not(inputs(166));
    layer0_outputs(1971) <= not((inputs(169)) or (inputs(2)));
    layer0_outputs(1972) <= (inputs(123)) and not (inputs(194));
    layer0_outputs(1973) <= not((inputs(129)) or (inputs(133)));
    layer0_outputs(1974) <= inputs(118);
    layer0_outputs(1975) <= not(inputs(213));
    layer0_outputs(1976) <= not(inputs(22)) or (inputs(162));
    layer0_outputs(1977) <= not(inputs(227));
    layer0_outputs(1978) <= not(inputs(234));
    layer0_outputs(1979) <= not(inputs(180));
    layer0_outputs(1980) <= not(inputs(134));
    layer0_outputs(1981) <= not((inputs(3)) and (inputs(79)));
    layer0_outputs(1982) <= not((inputs(55)) or (inputs(148)));
    layer0_outputs(1983) <= (inputs(250)) xor (inputs(255));
    layer0_outputs(1984) <= '1';
    layer0_outputs(1985) <= not(inputs(139));
    layer0_outputs(1986) <= not((inputs(99)) or (inputs(202)));
    layer0_outputs(1987) <= not(inputs(62));
    layer0_outputs(1988) <= not(inputs(3));
    layer0_outputs(1989) <= not(inputs(228));
    layer0_outputs(1990) <= not(inputs(230)) or (inputs(91));
    layer0_outputs(1991) <= (inputs(187)) or (inputs(80));
    layer0_outputs(1992) <= not((inputs(228)) or (inputs(81)));
    layer0_outputs(1993) <= not(inputs(138));
    layer0_outputs(1994) <= not((inputs(134)) xor (inputs(104)));
    layer0_outputs(1995) <= (inputs(50)) or (inputs(16));
    layer0_outputs(1996) <= not(inputs(111));
    layer0_outputs(1997) <= not(inputs(163)) or (inputs(220));
    layer0_outputs(1998) <= (inputs(1)) and not (inputs(90));
    layer0_outputs(1999) <= (inputs(44)) or (inputs(50));
    layer0_outputs(2000) <= (inputs(96)) or (inputs(209));
    layer0_outputs(2001) <= inputs(183);
    layer0_outputs(2002) <= (inputs(35)) and not (inputs(193));
    layer0_outputs(2003) <= not(inputs(194));
    layer0_outputs(2004) <= (inputs(160)) or (inputs(2));
    layer0_outputs(2005) <= not(inputs(181)) or (inputs(101));
    layer0_outputs(2006) <= inputs(69);
    layer0_outputs(2007) <= not(inputs(85));
    layer0_outputs(2008) <= not((inputs(24)) and (inputs(214)));
    layer0_outputs(2009) <= not((inputs(94)) or (inputs(224)));
    layer0_outputs(2010) <= inputs(167);
    layer0_outputs(2011) <= not(inputs(231)) or (inputs(6));
    layer0_outputs(2012) <= inputs(121);
    layer0_outputs(2013) <= (inputs(42)) or (inputs(124));
    layer0_outputs(2014) <= not((inputs(22)) or (inputs(84)));
    layer0_outputs(2015) <= inputs(50);
    layer0_outputs(2016) <= not(inputs(51)) or (inputs(144));
    layer0_outputs(2017) <= (inputs(252)) and not (inputs(39));
    layer0_outputs(2018) <= (inputs(154)) and not (inputs(62));
    layer0_outputs(2019) <= not((inputs(177)) or (inputs(247)));
    layer0_outputs(2020) <= not(inputs(51));
    layer0_outputs(2021) <= (inputs(180)) and not (inputs(107));
    layer0_outputs(2022) <= not(inputs(79)) or (inputs(152));
    layer0_outputs(2023) <= not(inputs(26));
    layer0_outputs(2024) <= (inputs(34)) or (inputs(54));
    layer0_outputs(2025) <= not((inputs(174)) and (inputs(175)));
    layer0_outputs(2026) <= not(inputs(148));
    layer0_outputs(2027) <= not(inputs(146));
    layer0_outputs(2028) <= not(inputs(230)) or (inputs(71));
    layer0_outputs(2029) <= not(inputs(233));
    layer0_outputs(2030) <= (inputs(131)) and not (inputs(8));
    layer0_outputs(2031) <= not(inputs(245));
    layer0_outputs(2032) <= inputs(141);
    layer0_outputs(2033) <= (inputs(211)) or (inputs(8));
    layer0_outputs(2034) <= (inputs(176)) and not (inputs(127));
    layer0_outputs(2035) <= not(inputs(225));
    layer0_outputs(2036) <= not((inputs(7)) or (inputs(159)));
    layer0_outputs(2037) <= inputs(169);
    layer0_outputs(2038) <= not((inputs(77)) or (inputs(192)));
    layer0_outputs(2039) <= not((inputs(60)) or (inputs(252)));
    layer0_outputs(2040) <= (inputs(165)) or (inputs(5));
    layer0_outputs(2041) <= (inputs(113)) or (inputs(29));
    layer0_outputs(2042) <= not((inputs(239)) or (inputs(186)));
    layer0_outputs(2043) <= not((inputs(123)) or (inputs(117)));
    layer0_outputs(2044) <= (inputs(118)) or (inputs(203));
    layer0_outputs(2045) <= not(inputs(147)) or (inputs(150));
    layer0_outputs(2046) <= inputs(183);
    layer0_outputs(2047) <= not(inputs(177));
    layer0_outputs(2048) <= (inputs(143)) or (inputs(131));
    layer0_outputs(2049) <= not((inputs(196)) or (inputs(227)));
    layer0_outputs(2050) <= not(inputs(68));
    layer0_outputs(2051) <= '0';
    layer0_outputs(2052) <= not(inputs(110)) or (inputs(15));
    layer0_outputs(2053) <= not((inputs(58)) or (inputs(107)));
    layer0_outputs(2054) <= '0';
    layer0_outputs(2055) <= not((inputs(120)) or (inputs(121)));
    layer0_outputs(2056) <= not(inputs(173)) or (inputs(126));
    layer0_outputs(2057) <= not((inputs(224)) or (inputs(238)));
    layer0_outputs(2058) <= (inputs(246)) or (inputs(128));
    layer0_outputs(2059) <= (inputs(28)) or (inputs(92));
    layer0_outputs(2060) <= not(inputs(214));
    layer0_outputs(2061) <= (inputs(108)) or (inputs(224));
    layer0_outputs(2062) <= (inputs(7)) and not (inputs(97));
    layer0_outputs(2063) <= not((inputs(164)) xor (inputs(200)));
    layer0_outputs(2064) <= not(inputs(229)) or (inputs(252));
    layer0_outputs(2065) <= inputs(100);
    layer0_outputs(2066) <= (inputs(107)) and not (inputs(131));
    layer0_outputs(2067) <= not((inputs(225)) and (inputs(240)));
    layer0_outputs(2068) <= inputs(91);
    layer0_outputs(2069) <= not(inputs(190));
    layer0_outputs(2070) <= inputs(218);
    layer0_outputs(2071) <= not((inputs(112)) xor (inputs(186)));
    layer0_outputs(2072) <= not(inputs(98));
    layer0_outputs(2073) <= inputs(217);
    layer0_outputs(2074) <= inputs(180);
    layer0_outputs(2075) <= not((inputs(167)) or (inputs(48)));
    layer0_outputs(2076) <= not(inputs(235));
    layer0_outputs(2077) <= inputs(130);
    layer0_outputs(2078) <= inputs(177);
    layer0_outputs(2079) <= not(inputs(52));
    layer0_outputs(2080) <= not(inputs(122));
    layer0_outputs(2081) <= (inputs(201)) and not (inputs(213));
    layer0_outputs(2082) <= not((inputs(147)) or (inputs(236)));
    layer0_outputs(2083) <= (inputs(37)) and not (inputs(209));
    layer0_outputs(2084) <= inputs(196);
    layer0_outputs(2085) <= inputs(69);
    layer0_outputs(2086) <= not((inputs(46)) or (inputs(35)));
    layer0_outputs(2087) <= not((inputs(1)) or (inputs(34)));
    layer0_outputs(2088) <= inputs(52);
    layer0_outputs(2089) <= not((inputs(74)) or (inputs(237)));
    layer0_outputs(2090) <= inputs(210);
    layer0_outputs(2091) <= (inputs(99)) and not (inputs(50));
    layer0_outputs(2092) <= not(inputs(230));
    layer0_outputs(2093) <= not(inputs(133));
    layer0_outputs(2094) <= (inputs(232)) xor (inputs(236));
    layer0_outputs(2095) <= (inputs(23)) and not (inputs(141));
    layer0_outputs(2096) <= not(inputs(234)) or (inputs(104));
    layer0_outputs(2097) <= not(inputs(223)) or (inputs(14));
    layer0_outputs(2098) <= not(inputs(4)) or (inputs(96));
    layer0_outputs(2099) <= not((inputs(101)) xor (inputs(177)));
    layer0_outputs(2100) <= not((inputs(35)) or (inputs(191)));
    layer0_outputs(2101) <= (inputs(56)) and not (inputs(22));
    layer0_outputs(2102) <= (inputs(123)) and not (inputs(47));
    layer0_outputs(2103) <= not((inputs(203)) and (inputs(216)));
    layer0_outputs(2104) <= (inputs(116)) or (inputs(222));
    layer0_outputs(2105) <= not(inputs(154));
    layer0_outputs(2106) <= (inputs(139)) or (inputs(204));
    layer0_outputs(2107) <= not(inputs(17)) or (inputs(214));
    layer0_outputs(2108) <= inputs(39);
    layer0_outputs(2109) <= inputs(65);
    layer0_outputs(2110) <= not(inputs(13));
    layer0_outputs(2111) <= not(inputs(58)) or (inputs(88));
    layer0_outputs(2112) <= inputs(165);
    layer0_outputs(2113) <= inputs(248);
    layer0_outputs(2114) <= inputs(79);
    layer0_outputs(2115) <= (inputs(101)) and not (inputs(125));
    layer0_outputs(2116) <= inputs(130);
    layer0_outputs(2117) <= not((inputs(94)) or (inputs(76)));
    layer0_outputs(2118) <= not(inputs(192));
    layer0_outputs(2119) <= not((inputs(200)) or (inputs(239)));
    layer0_outputs(2120) <= not(inputs(29));
    layer0_outputs(2121) <= not(inputs(171));
    layer0_outputs(2122) <= (inputs(87)) and not (inputs(177));
    layer0_outputs(2123) <= not(inputs(146));
    layer0_outputs(2124) <= (inputs(73)) or (inputs(198));
    layer0_outputs(2125) <= not((inputs(202)) or (inputs(113)));
    layer0_outputs(2126) <= (inputs(233)) or (inputs(161));
    layer0_outputs(2127) <= (inputs(210)) xor (inputs(190));
    layer0_outputs(2128) <= not((inputs(43)) or (inputs(47)));
    layer0_outputs(2129) <= inputs(225);
    layer0_outputs(2130) <= inputs(222);
    layer0_outputs(2131) <= not(inputs(131));
    layer0_outputs(2132) <= (inputs(81)) or (inputs(70));
    layer0_outputs(2133) <= inputs(225);
    layer0_outputs(2134) <= (inputs(217)) and not (inputs(78));
    layer0_outputs(2135) <= not(inputs(40)) or (inputs(45));
    layer0_outputs(2136) <= (inputs(31)) xor (inputs(40));
    layer0_outputs(2137) <= not(inputs(181)) or (inputs(67));
    layer0_outputs(2138) <= inputs(119);
    layer0_outputs(2139) <= (inputs(233)) and not (inputs(4));
    layer0_outputs(2140) <= not(inputs(233));
    layer0_outputs(2141) <= not(inputs(140));
    layer0_outputs(2142) <= not(inputs(33));
    layer0_outputs(2143) <= (inputs(195)) or (inputs(190));
    layer0_outputs(2144) <= not(inputs(213));
    layer0_outputs(2145) <= (inputs(113)) and not (inputs(255));
    layer0_outputs(2146) <= not((inputs(106)) or (inputs(240)));
    layer0_outputs(2147) <= (inputs(212)) or (inputs(255));
    layer0_outputs(2148) <= not(inputs(120));
    layer0_outputs(2149) <= (inputs(196)) or (inputs(46));
    layer0_outputs(2150) <= not(inputs(234)) or (inputs(14));
    layer0_outputs(2151) <= (inputs(12)) and not (inputs(3));
    layer0_outputs(2152) <= (inputs(142)) or (inputs(250));
    layer0_outputs(2153) <= (inputs(115)) or (inputs(142));
    layer0_outputs(2154) <= inputs(100);
    layer0_outputs(2155) <= inputs(88);
    layer0_outputs(2156) <= not(inputs(218));
    layer0_outputs(2157) <= (inputs(159)) or (inputs(142));
    layer0_outputs(2158) <= not(inputs(24)) or (inputs(113));
    layer0_outputs(2159) <= (inputs(42)) and not (inputs(204));
    layer0_outputs(2160) <= (inputs(148)) or (inputs(236));
    layer0_outputs(2161) <= not(inputs(91));
    layer0_outputs(2162) <= (inputs(8)) and not (inputs(197));
    layer0_outputs(2163) <= not((inputs(49)) or (inputs(91)));
    layer0_outputs(2164) <= not(inputs(83));
    layer0_outputs(2165) <= not(inputs(170));
    layer0_outputs(2166) <= not((inputs(80)) or (inputs(162)));
    layer0_outputs(2167) <= not(inputs(25)) or (inputs(84));
    layer0_outputs(2168) <= not(inputs(91));
    layer0_outputs(2169) <= not(inputs(196));
    layer0_outputs(2170) <= '0';
    layer0_outputs(2171) <= not(inputs(68)) or (inputs(125));
    layer0_outputs(2172) <= '1';
    layer0_outputs(2173) <= (inputs(168)) and not (inputs(253));
    layer0_outputs(2174) <= not((inputs(63)) xor (inputs(207)));
    layer0_outputs(2175) <= inputs(116);
    layer0_outputs(2176) <= inputs(195);
    layer0_outputs(2177) <= inputs(219);
    layer0_outputs(2178) <= not(inputs(145)) or (inputs(17));
    layer0_outputs(2179) <= not(inputs(40));
    layer0_outputs(2180) <= not(inputs(69)) or (inputs(241));
    layer0_outputs(2181) <= not((inputs(157)) or (inputs(5)));
    layer0_outputs(2182) <= '1';
    layer0_outputs(2183) <= not((inputs(169)) or (inputs(80)));
    layer0_outputs(2184) <= not(inputs(142));
    layer0_outputs(2185) <= inputs(17);
    layer0_outputs(2186) <= not(inputs(91));
    layer0_outputs(2187) <= inputs(234);
    layer0_outputs(2188) <= not(inputs(199)) or (inputs(52));
    layer0_outputs(2189) <= not((inputs(72)) xor (inputs(42)));
    layer0_outputs(2190) <= not(inputs(227));
    layer0_outputs(2191) <= inputs(245);
    layer0_outputs(2192) <= not(inputs(139));
    layer0_outputs(2193) <= (inputs(244)) and not (inputs(132));
    layer0_outputs(2194) <= (inputs(7)) and not (inputs(49));
    layer0_outputs(2195) <= not(inputs(101)) or (inputs(174));
    layer0_outputs(2196) <= inputs(98);
    layer0_outputs(2197) <= not((inputs(188)) xor (inputs(250)));
    layer0_outputs(2198) <= (inputs(209)) or (inputs(18));
    layer0_outputs(2199) <= not(inputs(89));
    layer0_outputs(2200) <= not((inputs(145)) or (inputs(116)));
    layer0_outputs(2201) <= inputs(203);
    layer0_outputs(2202) <= (inputs(149)) and not (inputs(51));
    layer0_outputs(2203) <= (inputs(12)) xor (inputs(109));
    layer0_outputs(2204) <= inputs(227);
    layer0_outputs(2205) <= not((inputs(254)) or (inputs(3)));
    layer0_outputs(2206) <= not(inputs(164));
    layer0_outputs(2207) <= inputs(82);
    layer0_outputs(2208) <= (inputs(255)) or (inputs(92));
    layer0_outputs(2209) <= '1';
    layer0_outputs(2210) <= not((inputs(112)) xor (inputs(116)));
    layer0_outputs(2211) <= not(inputs(19));
    layer0_outputs(2212) <= (inputs(219)) or (inputs(203));
    layer0_outputs(2213) <= (inputs(17)) or (inputs(238));
    layer0_outputs(2214) <= not(inputs(154));
    layer0_outputs(2215) <= (inputs(196)) and not (inputs(30));
    layer0_outputs(2216) <= not((inputs(187)) or (inputs(17)));
    layer0_outputs(2217) <= inputs(55);
    layer0_outputs(2218) <= not(inputs(33)) or (inputs(150));
    layer0_outputs(2219) <= not(inputs(215)) or (inputs(142));
    layer0_outputs(2220) <= (inputs(189)) and not (inputs(18));
    layer0_outputs(2221) <= (inputs(174)) or (inputs(27));
    layer0_outputs(2222) <= inputs(231);
    layer0_outputs(2223) <= not(inputs(68)) or (inputs(79));
    layer0_outputs(2224) <= inputs(212);
    layer0_outputs(2225) <= (inputs(103)) and not (inputs(15));
    layer0_outputs(2226) <= (inputs(27)) or (inputs(11));
    layer0_outputs(2227) <= '1';
    layer0_outputs(2228) <= not(inputs(20));
    layer0_outputs(2229) <= inputs(68);
    layer0_outputs(2230) <= not((inputs(220)) xor (inputs(187)));
    layer0_outputs(2231) <= not(inputs(219)) or (inputs(237));
    layer0_outputs(2232) <= inputs(153);
    layer0_outputs(2233) <= inputs(122);
    layer0_outputs(2234) <= not((inputs(123)) or (inputs(48)));
    layer0_outputs(2235) <= not(inputs(249));
    layer0_outputs(2236) <= inputs(184);
    layer0_outputs(2237) <= inputs(232);
    layer0_outputs(2238) <= (inputs(243)) or (inputs(22));
    layer0_outputs(2239) <= not((inputs(158)) or (inputs(127)));
    layer0_outputs(2240) <= (inputs(53)) and (inputs(45));
    layer0_outputs(2241) <= not(inputs(213)) or (inputs(241));
    layer0_outputs(2242) <= inputs(64);
    layer0_outputs(2243) <= inputs(155);
    layer0_outputs(2244) <= (inputs(9)) or (inputs(41));
    layer0_outputs(2245) <= (inputs(14)) or (inputs(206));
    layer0_outputs(2246) <= inputs(249);
    layer0_outputs(2247) <= '0';
    layer0_outputs(2248) <= not(inputs(114));
    layer0_outputs(2249) <= not(inputs(120));
    layer0_outputs(2250) <= (inputs(63)) or (inputs(232));
    layer0_outputs(2251) <= (inputs(31)) or (inputs(19));
    layer0_outputs(2252) <= (inputs(66)) and not (inputs(75));
    layer0_outputs(2253) <= (inputs(30)) and not (inputs(185));
    layer0_outputs(2254) <= not((inputs(194)) or (inputs(67)));
    layer0_outputs(2255) <= (inputs(105)) and not (inputs(85));
    layer0_outputs(2256) <= not(inputs(182)) or (inputs(1));
    layer0_outputs(2257) <= '1';
    layer0_outputs(2258) <= inputs(237);
    layer0_outputs(2259) <= inputs(144);
    layer0_outputs(2260) <= inputs(25);
    layer0_outputs(2261) <= not(inputs(137));
    layer0_outputs(2262) <= '0';
    layer0_outputs(2263) <= not(inputs(78));
    layer0_outputs(2264) <= inputs(23);
    layer0_outputs(2265) <= (inputs(3)) or (inputs(197));
    layer0_outputs(2266) <= not(inputs(238));
    layer0_outputs(2267) <= (inputs(172)) and (inputs(172));
    layer0_outputs(2268) <= not(inputs(35)) or (inputs(177));
    layer0_outputs(2269) <= not(inputs(137));
    layer0_outputs(2270) <= inputs(198);
    layer0_outputs(2271) <= inputs(23);
    layer0_outputs(2272) <= not((inputs(4)) or (inputs(205)));
    layer0_outputs(2273) <= (inputs(10)) and not (inputs(175));
    layer0_outputs(2274) <= (inputs(198)) and not (inputs(218));
    layer0_outputs(2275) <= (inputs(203)) or (inputs(79));
    layer0_outputs(2276) <= not((inputs(114)) or (inputs(130)));
    layer0_outputs(2277) <= not(inputs(244));
    layer0_outputs(2278) <= not(inputs(25));
    layer0_outputs(2279) <= inputs(6);
    layer0_outputs(2280) <= (inputs(23)) or (inputs(47));
    layer0_outputs(2281) <= not(inputs(213)) or (inputs(105));
    layer0_outputs(2282) <= '1';
    layer0_outputs(2283) <= (inputs(177)) or (inputs(117));
    layer0_outputs(2284) <= inputs(84);
    layer0_outputs(2285) <= not((inputs(70)) or (inputs(166)));
    layer0_outputs(2286) <= not((inputs(143)) or (inputs(194)));
    layer0_outputs(2287) <= not(inputs(84));
    layer0_outputs(2288) <= inputs(82);
    layer0_outputs(2289) <= not((inputs(124)) xor (inputs(158)));
    layer0_outputs(2290) <= not((inputs(221)) or (inputs(123)));
    layer0_outputs(2291) <= not(inputs(153)) or (inputs(241));
    layer0_outputs(2292) <= (inputs(138)) and not (inputs(46));
    layer0_outputs(2293) <= '1';
    layer0_outputs(2294) <= inputs(204);
    layer0_outputs(2295) <= not((inputs(31)) or (inputs(122)));
    layer0_outputs(2296) <= inputs(197);
    layer0_outputs(2297) <= not(inputs(227));
    layer0_outputs(2298) <= (inputs(212)) or (inputs(107));
    layer0_outputs(2299) <= inputs(7);
    layer0_outputs(2300) <= not(inputs(87));
    layer0_outputs(2301) <= '0';
    layer0_outputs(2302) <= not((inputs(31)) or (inputs(33)));
    layer0_outputs(2303) <= not(inputs(23)) or (inputs(192));
    layer0_outputs(2304) <= (inputs(217)) or (inputs(192));
    layer0_outputs(2305) <= not((inputs(152)) or (inputs(125)));
    layer0_outputs(2306) <= '1';
    layer0_outputs(2307) <= (inputs(206)) or (inputs(57));
    layer0_outputs(2308) <= not(inputs(118));
    layer0_outputs(2309) <= (inputs(24)) and not (inputs(249));
    layer0_outputs(2310) <= not(inputs(247));
    layer0_outputs(2311) <= (inputs(28)) and not (inputs(222));
    layer0_outputs(2312) <= (inputs(116)) or (inputs(186));
    layer0_outputs(2313) <= (inputs(165)) and not (inputs(47));
    layer0_outputs(2314) <= not(inputs(88));
    layer0_outputs(2315) <= not(inputs(90));
    layer0_outputs(2316) <= not(inputs(91));
    layer0_outputs(2317) <= (inputs(211)) or (inputs(190));
    layer0_outputs(2318) <= not(inputs(179));
    layer0_outputs(2319) <= not((inputs(11)) and (inputs(46)));
    layer0_outputs(2320) <= not(inputs(187)) or (inputs(254));
    layer0_outputs(2321) <= (inputs(59)) or (inputs(246));
    layer0_outputs(2322) <= not((inputs(82)) or (inputs(154)));
    layer0_outputs(2323) <= inputs(8);
    layer0_outputs(2324) <= inputs(94);
    layer0_outputs(2325) <= inputs(248);
    layer0_outputs(2326) <= not(inputs(6)) or (inputs(75));
    layer0_outputs(2327) <= not((inputs(169)) and (inputs(198)));
    layer0_outputs(2328) <= not(inputs(19)) or (inputs(76));
    layer0_outputs(2329) <= inputs(121);
    layer0_outputs(2330) <= (inputs(228)) or (inputs(139));
    layer0_outputs(2331) <= (inputs(217)) and not (inputs(49));
    layer0_outputs(2332) <= not(inputs(151));
    layer0_outputs(2333) <= not(inputs(194));
    layer0_outputs(2334) <= inputs(170);
    layer0_outputs(2335) <= (inputs(157)) and (inputs(186));
    layer0_outputs(2336) <= not((inputs(111)) xor (inputs(90)));
    layer0_outputs(2337) <= not(inputs(100));
    layer0_outputs(2338) <= not(inputs(114));
    layer0_outputs(2339) <= (inputs(75)) and not (inputs(163));
    layer0_outputs(2340) <= inputs(106);
    layer0_outputs(2341) <= (inputs(98)) or (inputs(185));
    layer0_outputs(2342) <= not(inputs(200));
    layer0_outputs(2343) <= not((inputs(40)) xor (inputs(42)));
    layer0_outputs(2344) <= inputs(166);
    layer0_outputs(2345) <= not(inputs(55)) or (inputs(2));
    layer0_outputs(2346) <= (inputs(222)) xor (inputs(140));
    layer0_outputs(2347) <= not((inputs(47)) or (inputs(71)));
    layer0_outputs(2348) <= not((inputs(246)) or (inputs(158)));
    layer0_outputs(2349) <= inputs(120);
    layer0_outputs(2350) <= not(inputs(122));
    layer0_outputs(2351) <= not(inputs(132));
    layer0_outputs(2352) <= not((inputs(6)) or (inputs(106)));
    layer0_outputs(2353) <= not((inputs(156)) or (inputs(143)));
    layer0_outputs(2354) <= not(inputs(93));
    layer0_outputs(2355) <= not(inputs(234));
    layer0_outputs(2356) <= not(inputs(117));
    layer0_outputs(2357) <= not((inputs(113)) or (inputs(48)));
    layer0_outputs(2358) <= (inputs(131)) or (inputs(140));
    layer0_outputs(2359) <= not(inputs(20));
    layer0_outputs(2360) <= not(inputs(195));
    layer0_outputs(2361) <= inputs(152);
    layer0_outputs(2362) <= (inputs(228)) or (inputs(176));
    layer0_outputs(2363) <= inputs(56);
    layer0_outputs(2364) <= inputs(132);
    layer0_outputs(2365) <= not(inputs(120));
    layer0_outputs(2366) <= not((inputs(126)) or (inputs(114)));
    layer0_outputs(2367) <= (inputs(139)) xor (inputs(121));
    layer0_outputs(2368) <= not(inputs(205)) or (inputs(14));
    layer0_outputs(2369) <= not(inputs(212));
    layer0_outputs(2370) <= not(inputs(134));
    layer0_outputs(2371) <= not((inputs(3)) xor (inputs(222)));
    layer0_outputs(2372) <= not((inputs(75)) xor (inputs(89)));
    layer0_outputs(2373) <= not(inputs(207));
    layer0_outputs(2374) <= not(inputs(90));
    layer0_outputs(2375) <= not(inputs(27)) or (inputs(189));
    layer0_outputs(2376) <= (inputs(229)) or (inputs(133));
    layer0_outputs(2377) <= (inputs(76)) or (inputs(22));
    layer0_outputs(2378) <= inputs(100);
    layer0_outputs(2379) <= not(inputs(231));
    layer0_outputs(2380) <= (inputs(124)) or (inputs(78));
    layer0_outputs(2381) <= '1';
    layer0_outputs(2382) <= inputs(159);
    layer0_outputs(2383) <= inputs(212);
    layer0_outputs(2384) <= not((inputs(76)) or (inputs(45)));
    layer0_outputs(2385) <= not(inputs(244)) or (inputs(19));
    layer0_outputs(2386) <= (inputs(225)) or (inputs(158));
    layer0_outputs(2387) <= (inputs(198)) or (inputs(193));
    layer0_outputs(2388) <= not((inputs(250)) or (inputs(37)));
    layer0_outputs(2389) <= not(inputs(198));
    layer0_outputs(2390) <= not(inputs(140));
    layer0_outputs(2391) <= (inputs(216)) and not (inputs(129));
    layer0_outputs(2392) <= not((inputs(72)) or (inputs(42)));
    layer0_outputs(2393) <= not(inputs(39)) or (inputs(63));
    layer0_outputs(2394) <= not(inputs(79)) or (inputs(189));
    layer0_outputs(2395) <= not((inputs(42)) or (inputs(159)));
    layer0_outputs(2396) <= (inputs(234)) and not (inputs(130));
    layer0_outputs(2397) <= not(inputs(190));
    layer0_outputs(2398) <= not(inputs(232));
    layer0_outputs(2399) <= not(inputs(118));
    layer0_outputs(2400) <= not((inputs(143)) or (inputs(231)));
    layer0_outputs(2401) <= (inputs(232)) and not (inputs(15));
    layer0_outputs(2402) <= inputs(132);
    layer0_outputs(2403) <= (inputs(133)) and not (inputs(109));
    layer0_outputs(2404) <= (inputs(246)) or (inputs(76));
    layer0_outputs(2405) <= inputs(164);
    layer0_outputs(2406) <= (inputs(72)) and not (inputs(33));
    layer0_outputs(2407) <= (inputs(4)) and not (inputs(208));
    layer0_outputs(2408) <= (inputs(180)) and not (inputs(192));
    layer0_outputs(2409) <= (inputs(14)) and not (inputs(242));
    layer0_outputs(2410) <= (inputs(160)) xor (inputs(39));
    layer0_outputs(2411) <= '1';
    layer0_outputs(2412) <= inputs(41);
    layer0_outputs(2413) <= (inputs(65)) or (inputs(80));
    layer0_outputs(2414) <= (inputs(24)) or (inputs(213));
    layer0_outputs(2415) <= inputs(25);
    layer0_outputs(2416) <= inputs(48);
    layer0_outputs(2417) <= (inputs(204)) and not (inputs(170));
    layer0_outputs(2418) <= not(inputs(4));
    layer0_outputs(2419) <= not(inputs(129));
    layer0_outputs(2420) <= not((inputs(103)) or (inputs(169)));
    layer0_outputs(2421) <= '1';
    layer0_outputs(2422) <= inputs(16);
    layer0_outputs(2423) <= (inputs(223)) or (inputs(116));
    layer0_outputs(2424) <= inputs(151);
    layer0_outputs(2425) <= (inputs(99)) or (inputs(124));
    layer0_outputs(2426) <= (inputs(115)) or (inputs(27));
    layer0_outputs(2427) <= not(inputs(162));
    layer0_outputs(2428) <= not(inputs(170));
    layer0_outputs(2429) <= not(inputs(87)) or (inputs(171));
    layer0_outputs(2430) <= not((inputs(17)) or (inputs(160)));
    layer0_outputs(2431) <= (inputs(157)) and not (inputs(29));
    layer0_outputs(2432) <= inputs(160);
    layer0_outputs(2433) <= (inputs(89)) and not (inputs(50));
    layer0_outputs(2434) <= inputs(227);
    layer0_outputs(2435) <= not(inputs(136)) or (inputs(96));
    layer0_outputs(2436) <= (inputs(98)) or (inputs(109));
    layer0_outputs(2437) <= not(inputs(238));
    layer0_outputs(2438) <= inputs(172);
    layer0_outputs(2439) <= (inputs(50)) or (inputs(151));
    layer0_outputs(2440) <= (inputs(125)) or (inputs(160));
    layer0_outputs(2441) <= not((inputs(207)) or (inputs(222)));
    layer0_outputs(2442) <= not(inputs(26)) or (inputs(139));
    layer0_outputs(2443) <= not(inputs(141)) or (inputs(107));
    layer0_outputs(2444) <= (inputs(51)) or (inputs(13));
    layer0_outputs(2445) <= not(inputs(100));
    layer0_outputs(2446) <= inputs(147);
    layer0_outputs(2447) <= inputs(2);
    layer0_outputs(2448) <= not((inputs(244)) and (inputs(134)));
    layer0_outputs(2449) <= inputs(215);
    layer0_outputs(2450) <= inputs(106);
    layer0_outputs(2451) <= not(inputs(211)) or (inputs(16));
    layer0_outputs(2452) <= not(inputs(220));
    layer0_outputs(2453) <= not(inputs(200));
    layer0_outputs(2454) <= (inputs(244)) or (inputs(173));
    layer0_outputs(2455) <= not(inputs(181));
    layer0_outputs(2456) <= inputs(154);
    layer0_outputs(2457) <= not((inputs(223)) or (inputs(141)));
    layer0_outputs(2458) <= inputs(38);
    layer0_outputs(2459) <= not((inputs(65)) and (inputs(132)));
    layer0_outputs(2460) <= not((inputs(8)) or (inputs(236)));
    layer0_outputs(2461) <= not((inputs(38)) or (inputs(49)));
    layer0_outputs(2462) <= (inputs(247)) and not (inputs(49));
    layer0_outputs(2463) <= (inputs(193)) and not (inputs(127));
    layer0_outputs(2464) <= not(inputs(133)) or (inputs(36));
    layer0_outputs(2465) <= not(inputs(126));
    layer0_outputs(2466) <= (inputs(5)) or (inputs(20));
    layer0_outputs(2467) <= (inputs(38)) and (inputs(122));
    layer0_outputs(2468) <= not(inputs(227));
    layer0_outputs(2469) <= (inputs(112)) or (inputs(159));
    layer0_outputs(2470) <= not(inputs(184));
    layer0_outputs(2471) <= (inputs(122)) and not (inputs(218));
    layer0_outputs(2472) <= (inputs(140)) or (inputs(3));
    layer0_outputs(2473) <= not(inputs(248)) or (inputs(91));
    layer0_outputs(2474) <= (inputs(226)) and not (inputs(138));
    layer0_outputs(2475) <= inputs(216);
    layer0_outputs(2476) <= not(inputs(122));
    layer0_outputs(2477) <= not(inputs(121));
    layer0_outputs(2478) <= not((inputs(60)) or (inputs(226)));
    layer0_outputs(2479) <= not(inputs(93));
    layer0_outputs(2480) <= (inputs(77)) or (inputs(175));
    layer0_outputs(2481) <= not(inputs(90));
    layer0_outputs(2482) <= (inputs(41)) or (inputs(33));
    layer0_outputs(2483) <= inputs(148);
    layer0_outputs(2484) <= not(inputs(68)) or (inputs(60));
    layer0_outputs(2485) <= not((inputs(238)) xor (inputs(24)));
    layer0_outputs(2486) <= (inputs(42)) and not (inputs(152));
    layer0_outputs(2487) <= not((inputs(182)) or (inputs(146)));
    layer0_outputs(2488) <= (inputs(173)) or (inputs(69));
    layer0_outputs(2489) <= not(inputs(226));
    layer0_outputs(2490) <= '1';
    layer0_outputs(2491) <= '1';
    layer0_outputs(2492) <= not(inputs(234));
    layer0_outputs(2493) <= inputs(115);
    layer0_outputs(2494) <= not((inputs(119)) and (inputs(230)));
    layer0_outputs(2495) <= not(inputs(151));
    layer0_outputs(2496) <= not(inputs(136));
    layer0_outputs(2497) <= not((inputs(13)) or (inputs(190)));
    layer0_outputs(2498) <= (inputs(130)) or (inputs(236));
    layer0_outputs(2499) <= not(inputs(66));
    layer0_outputs(2500) <= (inputs(86)) and (inputs(63));
    layer0_outputs(2501) <= not(inputs(74));
    layer0_outputs(2502) <= (inputs(229)) or (inputs(247));
    layer0_outputs(2503) <= inputs(196);
    layer0_outputs(2504) <= not((inputs(151)) or (inputs(185)));
    layer0_outputs(2505) <= inputs(58);
    layer0_outputs(2506) <= (inputs(34)) or (inputs(3));
    layer0_outputs(2507) <= (inputs(255)) or (inputs(225));
    layer0_outputs(2508) <= not(inputs(220)) or (inputs(15));
    layer0_outputs(2509) <= not((inputs(246)) or (inputs(15)));
    layer0_outputs(2510) <= '1';
    layer0_outputs(2511) <= not(inputs(57));
    layer0_outputs(2512) <= (inputs(61)) and not (inputs(130));
    layer0_outputs(2513) <= (inputs(232)) xor (inputs(208));
    layer0_outputs(2514) <= not(inputs(82));
    layer0_outputs(2515) <= (inputs(225)) or (inputs(202));
    layer0_outputs(2516) <= not(inputs(216));
    layer0_outputs(2517) <= not(inputs(26)) or (inputs(206));
    layer0_outputs(2518) <= (inputs(47)) or (inputs(101));
    layer0_outputs(2519) <= (inputs(251)) or (inputs(152));
    layer0_outputs(2520) <= (inputs(182)) xor (inputs(244));
    layer0_outputs(2521) <= not((inputs(77)) and (inputs(11)));
    layer0_outputs(2522) <= inputs(212);
    layer0_outputs(2523) <= not((inputs(128)) or (inputs(110)));
    layer0_outputs(2524) <= (inputs(219)) or (inputs(32));
    layer0_outputs(2525) <= (inputs(249)) or (inputs(87));
    layer0_outputs(2526) <= not(inputs(140));
    layer0_outputs(2527) <= (inputs(183)) and not (inputs(113));
    layer0_outputs(2528) <= not((inputs(200)) or (inputs(98)));
    layer0_outputs(2529) <= (inputs(69)) or (inputs(181));
    layer0_outputs(2530) <= (inputs(180)) and not (inputs(32));
    layer0_outputs(2531) <= not(inputs(196));
    layer0_outputs(2532) <= (inputs(218)) and not (inputs(115));
    layer0_outputs(2533) <= not((inputs(98)) or (inputs(169)));
    layer0_outputs(2534) <= inputs(68);
    layer0_outputs(2535) <= not((inputs(235)) or (inputs(220)));
    layer0_outputs(2536) <= not(inputs(85));
    layer0_outputs(2537) <= (inputs(208)) or (inputs(15));
    layer0_outputs(2538) <= inputs(61);
    layer0_outputs(2539) <= (inputs(90)) or (inputs(207));
    layer0_outputs(2540) <= not((inputs(145)) or (inputs(130)));
    layer0_outputs(2541) <= not(inputs(90));
    layer0_outputs(2542) <= (inputs(71)) xor (inputs(165));
    layer0_outputs(2543) <= not(inputs(9)) or (inputs(83));
    layer0_outputs(2544) <= (inputs(92)) or (inputs(189));
    layer0_outputs(2545) <= (inputs(85)) and not (inputs(158));
    layer0_outputs(2546) <= not(inputs(147));
    layer0_outputs(2547) <= '0';
    layer0_outputs(2548) <= (inputs(171)) and not (inputs(32));
    layer0_outputs(2549) <= not((inputs(249)) or (inputs(70)));
    layer0_outputs(2550) <= not(inputs(47)) or (inputs(73));
    layer0_outputs(2551) <= (inputs(234)) or (inputs(127));
    layer0_outputs(2552) <= inputs(21);
    layer0_outputs(2553) <= (inputs(191)) or (inputs(187));
    layer0_outputs(2554) <= inputs(198);
    layer0_outputs(2555) <= not(inputs(229));
    layer0_outputs(2556) <= inputs(54);
    layer0_outputs(2557) <= not((inputs(166)) or (inputs(149)));
    layer0_outputs(2558) <= not(inputs(248));
    layer0_outputs(2559) <= not((inputs(200)) or (inputs(209)));
    outputs(0) <= not((layer0_outputs(278)) or (layer0_outputs(1468)));
    outputs(1) <= (layer0_outputs(868)) or (layer0_outputs(2515));
    outputs(2) <= not(layer0_outputs(404));
    outputs(3) <= not(layer0_outputs(699));
    outputs(4) <= not(layer0_outputs(1239));
    outputs(5) <= layer0_outputs(1901);
    outputs(6) <= (layer0_outputs(1828)) and (layer0_outputs(1559));
    outputs(7) <= (layer0_outputs(1765)) and not (layer0_outputs(2046));
    outputs(8) <= (layer0_outputs(2271)) xor (layer0_outputs(831));
    outputs(9) <= not((layer0_outputs(2456)) and (layer0_outputs(2394)));
    outputs(10) <= layer0_outputs(2504);
    outputs(11) <= not(layer0_outputs(1252));
    outputs(12) <= not(layer0_outputs(2263)) or (layer0_outputs(1384));
    outputs(13) <= not(layer0_outputs(2117));
    outputs(14) <= not(layer0_outputs(1064)) or (layer0_outputs(653));
    outputs(15) <= (layer0_outputs(761)) and not (layer0_outputs(2019));
    outputs(16) <= (layer0_outputs(527)) and (layer0_outputs(464));
    outputs(17) <= not(layer0_outputs(1092));
    outputs(18) <= (layer0_outputs(1764)) and not (layer0_outputs(1155));
    outputs(19) <= (layer0_outputs(1685)) and not (layer0_outputs(2549));
    outputs(20) <= not(layer0_outputs(520));
    outputs(21) <= not(layer0_outputs(1975));
    outputs(22) <= (layer0_outputs(1213)) and not (layer0_outputs(47));
    outputs(23) <= not(layer0_outputs(945));
    outputs(24) <= layer0_outputs(202);
    outputs(25) <= not(layer0_outputs(864));
    outputs(26) <= (layer0_outputs(2459)) and not (layer0_outputs(956));
    outputs(27) <= not(layer0_outputs(904));
    outputs(28) <= not((layer0_outputs(2509)) and (layer0_outputs(1248)));
    outputs(29) <= (layer0_outputs(1754)) and not (layer0_outputs(1703));
    outputs(30) <= layer0_outputs(412);
    outputs(31) <= not(layer0_outputs(2179));
    outputs(32) <= not(layer0_outputs(1385)) or (layer0_outputs(304));
    outputs(33) <= not((layer0_outputs(1895)) xor (layer0_outputs(475)));
    outputs(34) <= layer0_outputs(1478);
    outputs(35) <= not(layer0_outputs(2465));
    outputs(36) <= layer0_outputs(1016);
    outputs(37) <= not(layer0_outputs(1774));
    outputs(38) <= layer0_outputs(533);
    outputs(39) <= (layer0_outputs(1228)) and not (layer0_outputs(1426));
    outputs(40) <= not(layer0_outputs(265));
    outputs(41) <= not((layer0_outputs(1091)) or (layer0_outputs(404)));
    outputs(42) <= (layer0_outputs(2435)) and (layer0_outputs(142));
    outputs(43) <= not((layer0_outputs(311)) or (layer0_outputs(2049)));
    outputs(44) <= not((layer0_outputs(330)) or (layer0_outputs(1252)));
    outputs(45) <= not((layer0_outputs(1168)) or (layer0_outputs(83)));
    outputs(46) <= not(layer0_outputs(2027));
    outputs(47) <= (layer0_outputs(2084)) and not (layer0_outputs(1774));
    outputs(48) <= not(layer0_outputs(1960)) or (layer0_outputs(2431));
    outputs(49) <= (layer0_outputs(1416)) xor (layer0_outputs(2149));
    outputs(50) <= not(layer0_outputs(1425));
    outputs(51) <= not((layer0_outputs(1967)) and (layer0_outputs(1930)));
    outputs(52) <= (layer0_outputs(2522)) and not (layer0_outputs(49));
    outputs(53) <= not((layer0_outputs(2395)) or (layer0_outputs(1562)));
    outputs(54) <= not(layer0_outputs(782));
    outputs(55) <= not((layer0_outputs(1443)) or (layer0_outputs(615)));
    outputs(56) <= not(layer0_outputs(883));
    outputs(57) <= layer0_outputs(2105);
    outputs(58) <= not(layer0_outputs(606));
    outputs(59) <= not(layer0_outputs(907)) or (layer0_outputs(603));
    outputs(60) <= (layer0_outputs(1694)) xor (layer0_outputs(1610));
    outputs(61) <= not(layer0_outputs(177));
    outputs(62) <= not(layer0_outputs(2233));
    outputs(63) <= not(layer0_outputs(1299));
    outputs(64) <= not((layer0_outputs(882)) or (layer0_outputs(2010)));
    outputs(65) <= not(layer0_outputs(1454));
    outputs(66) <= layer0_outputs(1620);
    outputs(67) <= not(layer0_outputs(163));
    outputs(68) <= layer0_outputs(280);
    outputs(69) <= layer0_outputs(553);
    outputs(70) <= not(layer0_outputs(557));
    outputs(71) <= layer0_outputs(1646);
    outputs(72) <= layer0_outputs(1667);
    outputs(73) <= layer0_outputs(826);
    outputs(74) <= not(layer0_outputs(981));
    outputs(75) <= not((layer0_outputs(1267)) xor (layer0_outputs(423)));
    outputs(76) <= (layer0_outputs(1230)) xor (layer0_outputs(1756));
    outputs(77) <= layer0_outputs(2048);
    outputs(78) <= layer0_outputs(2215);
    outputs(79) <= layer0_outputs(526);
    outputs(80) <= not((layer0_outputs(1704)) and (layer0_outputs(534)));
    outputs(81) <= not(layer0_outputs(1550));
    outputs(82) <= not(layer0_outputs(1568));
    outputs(83) <= (layer0_outputs(361)) and not (layer0_outputs(2489));
    outputs(84) <= not(layer0_outputs(1697));
    outputs(85) <= not(layer0_outputs(1397));
    outputs(86) <= not((layer0_outputs(2255)) or (layer0_outputs(1181)));
    outputs(87) <= layer0_outputs(504);
    outputs(88) <= not(layer0_outputs(460));
    outputs(89) <= not((layer0_outputs(1511)) or (layer0_outputs(867)));
    outputs(90) <= (layer0_outputs(423)) and not (layer0_outputs(1342));
    outputs(91) <= not(layer0_outputs(2210));
    outputs(92) <= not(layer0_outputs(2400));
    outputs(93) <= layer0_outputs(1134);
    outputs(94) <= (layer0_outputs(1014)) and not (layer0_outputs(683));
    outputs(95) <= (layer0_outputs(950)) xor (layer0_outputs(1278));
    outputs(96) <= (layer0_outputs(2513)) and (layer0_outputs(328));
    outputs(97) <= not(layer0_outputs(1471)) or (layer0_outputs(2402));
    outputs(98) <= not((layer0_outputs(782)) or (layer0_outputs(658)));
    outputs(99) <= (layer0_outputs(1072)) and not (layer0_outputs(1397));
    outputs(100) <= layer0_outputs(92);
    outputs(101) <= layer0_outputs(2065);
    outputs(102) <= not(layer0_outputs(2393)) or (layer0_outputs(2432));
    outputs(103) <= (layer0_outputs(869)) or (layer0_outputs(963));
    outputs(104) <= not((layer0_outputs(1279)) xor (layer0_outputs(1978)));
    outputs(105) <= (layer0_outputs(1027)) and not (layer0_outputs(127));
    outputs(106) <= layer0_outputs(2420);
    outputs(107) <= (layer0_outputs(2425)) and not (layer0_outputs(2450));
    outputs(108) <= not(layer0_outputs(1123));
    outputs(109) <= not(layer0_outputs(877));
    outputs(110) <= layer0_outputs(2091);
    outputs(111) <= not(layer0_outputs(2392));
    outputs(112) <= not(layer0_outputs(1571));
    outputs(113) <= (layer0_outputs(294)) and (layer0_outputs(2229));
    outputs(114) <= layer0_outputs(547);
    outputs(115) <= (layer0_outputs(313)) and not (layer0_outputs(2253));
    outputs(116) <= not((layer0_outputs(2506)) or (layer0_outputs(855)));
    outputs(117) <= layer0_outputs(2269);
    outputs(118) <= not(layer0_outputs(710)) or (layer0_outputs(94));
    outputs(119) <= not(layer0_outputs(995)) or (layer0_outputs(844));
    outputs(120) <= not(layer0_outputs(2179));
    outputs(121) <= (layer0_outputs(2269)) and (layer0_outputs(263));
    outputs(122) <= layer0_outputs(2321);
    outputs(123) <= not(layer0_outputs(2022)) or (layer0_outputs(1883));
    outputs(124) <= not(layer0_outputs(564)) or (layer0_outputs(835));
    outputs(125) <= (layer0_outputs(327)) and not (layer0_outputs(409));
    outputs(126) <= (layer0_outputs(2401)) and (layer0_outputs(1050));
    outputs(127) <= not(layer0_outputs(0));
    outputs(128) <= not(layer0_outputs(1146));
    outputs(129) <= not(layer0_outputs(1319));
    outputs(130) <= (layer0_outputs(745)) and not (layer0_outputs(974));
    outputs(131) <= not((layer0_outputs(1065)) or (layer0_outputs(2344)));
    outputs(132) <= layer0_outputs(731);
    outputs(133) <= layer0_outputs(1392);
    outputs(134) <= layer0_outputs(794);
    outputs(135) <= (layer0_outputs(247)) and not (layer0_outputs(1974));
    outputs(136) <= (layer0_outputs(2389)) and not (layer0_outputs(744));
    outputs(137) <= not((layer0_outputs(230)) and (layer0_outputs(616)));
    outputs(138) <= not(layer0_outputs(1342)) or (layer0_outputs(26));
    outputs(139) <= (layer0_outputs(2137)) and not (layer0_outputs(1308));
    outputs(140) <= (layer0_outputs(2550)) and (layer0_outputs(852));
    outputs(141) <= (layer0_outputs(61)) or (layer0_outputs(597));
    outputs(142) <= not(layer0_outputs(1080));
    outputs(143) <= layer0_outputs(1412);
    outputs(144) <= layer0_outputs(1430);
    outputs(145) <= layer0_outputs(2302);
    outputs(146) <= (layer0_outputs(1687)) and not (layer0_outputs(1190));
    outputs(147) <= not(layer0_outputs(1108));
    outputs(148) <= (layer0_outputs(1610)) and (layer0_outputs(1910));
    outputs(149) <= not(layer0_outputs(903));
    outputs(150) <= (layer0_outputs(1016)) or (layer0_outputs(2446));
    outputs(151) <= not(layer0_outputs(1359));
    outputs(152) <= (layer0_outputs(1427)) and not (layer0_outputs(2200));
    outputs(153) <= (layer0_outputs(333)) or (layer0_outputs(400));
    outputs(154) <= (layer0_outputs(361)) xor (layer0_outputs(901));
    outputs(155) <= not(layer0_outputs(559)) or (layer0_outputs(562));
    outputs(156) <= not(layer0_outputs(1396));
    outputs(157) <= layer0_outputs(1510);
    outputs(158) <= not(layer0_outputs(641)) or (layer0_outputs(1374));
    outputs(159) <= (layer0_outputs(598)) and not (layer0_outputs(21));
    outputs(160) <= layer0_outputs(480);
    outputs(161) <= (layer0_outputs(2033)) and (layer0_outputs(2502));
    outputs(162) <= (layer0_outputs(1980)) and not (layer0_outputs(1483));
    outputs(163) <= (layer0_outputs(825)) or (layer0_outputs(1300));
    outputs(164) <= (layer0_outputs(1818)) and not (layer0_outputs(2213));
    outputs(165) <= not(layer0_outputs(1406));
    outputs(166) <= not(layer0_outputs(768));
    outputs(167) <= (layer0_outputs(1211)) or (layer0_outputs(76));
    outputs(168) <= (layer0_outputs(759)) and not (layer0_outputs(1024));
    outputs(169) <= not((layer0_outputs(879)) and (layer0_outputs(908)));
    outputs(170) <= (layer0_outputs(1994)) and (layer0_outputs(1455));
    outputs(171) <= not(layer0_outputs(583)) or (layer0_outputs(789));
    outputs(172) <= layer0_outputs(2420);
    outputs(173) <= not(layer0_outputs(655));
    outputs(174) <= (layer0_outputs(1258)) and (layer0_outputs(1618));
    outputs(175) <= not(layer0_outputs(725));
    outputs(176) <= layer0_outputs(866);
    outputs(177) <= not(layer0_outputs(2443)) or (layer0_outputs(1644));
    outputs(178) <= (layer0_outputs(1739)) or (layer0_outputs(1132));
    outputs(179) <= layer0_outputs(1582);
    outputs(180) <= layer0_outputs(1498);
    outputs(181) <= (layer0_outputs(253)) and (layer0_outputs(2214));
    outputs(182) <= layer0_outputs(1681);
    outputs(183) <= layer0_outputs(580);
    outputs(184) <= not(layer0_outputs(69));
    outputs(185) <= not(layer0_outputs(572));
    outputs(186) <= not((layer0_outputs(857)) or (layer0_outputs(1100)));
    outputs(187) <= not(layer0_outputs(2347)) or (layer0_outputs(1574));
    outputs(188) <= layer0_outputs(1196);
    outputs(189) <= not((layer0_outputs(612)) or (layer0_outputs(1538)));
    outputs(190) <= not((layer0_outputs(1334)) and (layer0_outputs(870)));
    outputs(191) <= (layer0_outputs(1409)) and (layer0_outputs(266));
    outputs(192) <= layer0_outputs(992);
    outputs(193) <= layer0_outputs(2085);
    outputs(194) <= layer0_outputs(250);
    outputs(195) <= layer0_outputs(851);
    outputs(196) <= not(layer0_outputs(1483));
    outputs(197) <= not(layer0_outputs(525));
    outputs(198) <= not((layer0_outputs(1997)) and (layer0_outputs(164)));
    outputs(199) <= (layer0_outputs(448)) and not (layer0_outputs(2360));
    outputs(200) <= not(layer0_outputs(397));
    outputs(201) <= (layer0_outputs(2221)) and (layer0_outputs(1768));
    outputs(202) <= (layer0_outputs(976)) and not (layer0_outputs(1094));
    outputs(203) <= (layer0_outputs(204)) and not (layer0_outputs(1414));
    outputs(204) <= not(layer0_outputs(1240));
    outputs(205) <= layer0_outputs(2522);
    outputs(206) <= (layer0_outputs(1494)) and (layer0_outputs(285));
    outputs(207) <= layer0_outputs(336);
    outputs(208) <= (layer0_outputs(874)) xor (layer0_outputs(796));
    outputs(209) <= not(layer0_outputs(2045));
    outputs(210) <= not(layer0_outputs(1309));
    outputs(211) <= layer0_outputs(703);
    outputs(212) <= not(layer0_outputs(2329));
    outputs(213) <= not(layer0_outputs(111));
    outputs(214) <= layer0_outputs(115);
    outputs(215) <= (layer0_outputs(2352)) and not (layer0_outputs(364));
    outputs(216) <= layer0_outputs(2098);
    outputs(217) <= not((layer0_outputs(2320)) or (layer0_outputs(485)));
    outputs(218) <= layer0_outputs(769);
    outputs(219) <= not(layer0_outputs(226));
    outputs(220) <= (layer0_outputs(2513)) and not (layer0_outputs(1367));
    outputs(221) <= not(layer0_outputs(1567)) or (layer0_outputs(897));
    outputs(222) <= not(layer0_outputs(838));
    outputs(223) <= (layer0_outputs(860)) and not (layer0_outputs(1632));
    outputs(224) <= not(layer0_outputs(1116)) or (layer0_outputs(798));
    outputs(225) <= not((layer0_outputs(83)) or (layer0_outputs(1726)));
    outputs(226) <= layer0_outputs(385);
    outputs(227) <= (layer0_outputs(1382)) and not (layer0_outputs(904));
    outputs(228) <= layer0_outputs(1494);
    outputs(229) <= not(layer0_outputs(370));
    outputs(230) <= not((layer0_outputs(1598)) and (layer0_outputs(2276)));
    outputs(231) <= layer0_outputs(938);
    outputs(232) <= layer0_outputs(2126);
    outputs(233) <= not(layer0_outputs(1422)) or (layer0_outputs(496));
    outputs(234) <= not(layer0_outputs(1799));
    outputs(235) <= not((layer0_outputs(1986)) or (layer0_outputs(1284)));
    outputs(236) <= not(layer0_outputs(741));
    outputs(237) <= not(layer0_outputs(1622));
    outputs(238) <= (layer0_outputs(673)) and (layer0_outputs(187));
    outputs(239) <= layer0_outputs(308);
    outputs(240) <= layer0_outputs(1212);
    outputs(241) <= layer0_outputs(497);
    outputs(242) <= (layer0_outputs(1293)) xor (layer0_outputs(1604));
    outputs(243) <= not(layer0_outputs(664));
    outputs(244) <= not(layer0_outputs(625));
    outputs(245) <= layer0_outputs(521);
    outputs(246) <= not(layer0_outputs(1507));
    outputs(247) <= not(layer0_outputs(1572)) or (layer0_outputs(329));
    outputs(248) <= (layer0_outputs(897)) or (layer0_outputs(1085));
    outputs(249) <= layer0_outputs(1897);
    outputs(250) <= layer0_outputs(1641);
    outputs(251) <= layer0_outputs(1350);
    outputs(252) <= not(layer0_outputs(282)) or (layer0_outputs(1658));
    outputs(253) <= not(layer0_outputs(1058));
    outputs(254) <= not(layer0_outputs(1762)) or (layer0_outputs(2382));
    outputs(255) <= not(layer0_outputs(849)) or (layer0_outputs(1932));
    outputs(256) <= (layer0_outputs(1780)) and not (layer0_outputs(603));
    outputs(257) <= not(layer0_outputs(1858));
    outputs(258) <= not((layer0_outputs(1944)) or (layer0_outputs(1437)));
    outputs(259) <= not((layer0_outputs(1788)) or (layer0_outputs(790)));
    outputs(260) <= (layer0_outputs(1924)) and not (layer0_outputs(774));
    outputs(261) <= (layer0_outputs(1817)) and not (layer0_outputs(1916));
    outputs(262) <= (layer0_outputs(2430)) and (layer0_outputs(1709));
    outputs(263) <= (layer0_outputs(62)) and (layer0_outputs(433));
    outputs(264) <= (layer0_outputs(171)) and not (layer0_outputs(1136));
    outputs(265) <= (layer0_outputs(1236)) and not (layer0_outputs(1165));
    outputs(266) <= (layer0_outputs(2042)) and not (layer0_outputs(1328));
    outputs(267) <= (layer0_outputs(2182)) and not (layer0_outputs(1732));
    outputs(268) <= (layer0_outputs(76)) and (layer0_outputs(1448));
    outputs(269) <= not((layer0_outputs(192)) or (layer0_outputs(540)));
    outputs(270) <= (layer0_outputs(200)) and (layer0_outputs(2478));
    outputs(271) <= '0';
    outputs(272) <= (layer0_outputs(2289)) and not (layer0_outputs(1920));
    outputs(273) <= (layer0_outputs(1186)) and (layer0_outputs(1292));
    outputs(274) <= not((layer0_outputs(2553)) or (layer0_outputs(709)));
    outputs(275) <= (layer0_outputs(735)) and not (layer0_outputs(1923));
    outputs(276) <= (layer0_outputs(1388)) and not (layer0_outputs(53));
    outputs(277) <= (layer0_outputs(37)) and not (layer0_outputs(415));
    outputs(278) <= not((layer0_outputs(829)) or (layer0_outputs(804)));
    outputs(279) <= (layer0_outputs(1352)) and not (layer0_outputs(689));
    outputs(280) <= (layer0_outputs(2183)) and not (layer0_outputs(622));
    outputs(281) <= (layer0_outputs(1314)) and (layer0_outputs(1202));
    outputs(282) <= (layer0_outputs(97)) and not (layer0_outputs(2376));
    outputs(283) <= (layer0_outputs(2086)) and not (layer0_outputs(1773));
    outputs(284) <= (layer0_outputs(2234)) and (layer0_outputs(2484));
    outputs(285) <= (layer0_outputs(1565)) and not (layer0_outputs(2382));
    outputs(286) <= not((layer0_outputs(1408)) or (layer0_outputs(2341)));
    outputs(287) <= (layer0_outputs(1048)) and not (layer0_outputs(1059));
    outputs(288) <= not(layer0_outputs(606));
    outputs(289) <= (layer0_outputs(1490)) and not (layer0_outputs(611));
    outputs(290) <= not((layer0_outputs(1670)) or (layer0_outputs(2059)));
    outputs(291) <= (layer0_outputs(1835)) and (layer0_outputs(252));
    outputs(292) <= (layer0_outputs(2231)) and not (layer0_outputs(875));
    outputs(293) <= (layer0_outputs(856)) and not (layer0_outputs(1528));
    outputs(294) <= not((layer0_outputs(611)) or (layer0_outputs(1266)));
    outputs(295) <= (layer0_outputs(1473)) and (layer0_outputs(2038));
    outputs(296) <= not(layer0_outputs(2280));
    outputs(297) <= layer0_outputs(1993);
    outputs(298) <= (layer0_outputs(1139)) and (layer0_outputs(1419));
    outputs(299) <= not((layer0_outputs(2275)) or (layer0_outputs(2544)));
    outputs(300) <= (layer0_outputs(1652)) and not (layer0_outputs(256));
    outputs(301) <= layer0_outputs(1234);
    outputs(302) <= (layer0_outputs(714)) and not (layer0_outputs(1661));
    outputs(303) <= (layer0_outputs(993)) and not (layer0_outputs(1995));
    outputs(304) <= (layer0_outputs(31)) and (layer0_outputs(287));
    outputs(305) <= (layer0_outputs(1415)) and not (layer0_outputs(602));
    outputs(306) <= (layer0_outputs(180)) and not (layer0_outputs(891));
    outputs(307) <= layer0_outputs(1871);
    outputs(308) <= (layer0_outputs(1938)) and not (layer0_outputs(1207));
    outputs(309) <= not((layer0_outputs(1723)) or (layer0_outputs(272)));
    outputs(310) <= (layer0_outputs(1223)) and not (layer0_outputs(1529));
    outputs(311) <= (layer0_outputs(1106)) and not (layer0_outputs(2498));
    outputs(312) <= (layer0_outputs(96)) and not (layer0_outputs(840));
    outputs(313) <= not(layer0_outputs(816));
    outputs(314) <= not(layer0_outputs(241));
    outputs(315) <= (layer0_outputs(29)) and (layer0_outputs(2296));
    outputs(316) <= layer0_outputs(401);
    outputs(317) <= (layer0_outputs(886)) and not (layer0_outputs(1209));
    outputs(318) <= (layer0_outputs(114)) and (layer0_outputs(1619));
    outputs(319) <= (layer0_outputs(775)) and not (layer0_outputs(2454));
    outputs(320) <= layer0_outputs(1108);
    outputs(321) <= (layer0_outputs(1987)) and (layer0_outputs(906));
    outputs(322) <= (layer0_outputs(2419)) and not (layer0_outputs(819));
    outputs(323) <= (layer0_outputs(1105)) and not (layer0_outputs(994));
    outputs(324) <= not((layer0_outputs(2544)) or (layer0_outputs(130)));
    outputs(325) <= not(layer0_outputs(2377));
    outputs(326) <= layer0_outputs(106);
    outputs(327) <= (layer0_outputs(187)) and (layer0_outputs(937));
    outputs(328) <= (layer0_outputs(2203)) xor (layer0_outputs(270));
    outputs(329) <= (layer0_outputs(1419)) and not (layer0_outputs(2539));
    outputs(330) <= (layer0_outputs(1248)) and not (layer0_outputs(1259));
    outputs(331) <= (layer0_outputs(627)) and not (layer0_outputs(2466));
    outputs(332) <= not((layer0_outputs(1553)) or (layer0_outputs(2185)));
    outputs(333) <= (layer0_outputs(2485)) and not (layer0_outputs(1907));
    outputs(334) <= (layer0_outputs(837)) and not (layer0_outputs(792));
    outputs(335) <= layer0_outputs(1234);
    outputs(336) <= layer0_outputs(403);
    outputs(337) <= (layer0_outputs(1285)) and (layer0_outputs(1451));
    outputs(338) <= (layer0_outputs(2295)) and not (layer0_outputs(173));
    outputs(339) <= (layer0_outputs(2357)) and not (layer0_outputs(2512));
    outputs(340) <= (layer0_outputs(1960)) and (layer0_outputs(922));
    outputs(341) <= (layer0_outputs(905)) and (layer0_outputs(1585));
    outputs(342) <= (layer0_outputs(1665)) and not (layer0_outputs(2285));
    outputs(343) <= (layer0_outputs(2322)) and not (layer0_outputs(1858));
    outputs(344) <= not((layer0_outputs(591)) or (layer0_outputs(2312)));
    outputs(345) <= not((layer0_outputs(1589)) or (layer0_outputs(730)));
    outputs(346) <= (layer0_outputs(2278)) and not (layer0_outputs(745));
    outputs(347) <= not((layer0_outputs(2503)) or (layer0_outputs(296)));
    outputs(348) <= not((layer0_outputs(2500)) or (layer0_outputs(761)));
    outputs(349) <= (layer0_outputs(813)) and not (layer0_outputs(1325));
    outputs(350) <= (layer0_outputs(1997)) and (layer0_outputs(667));
    outputs(351) <= (layer0_outputs(2477)) and not (layer0_outputs(701));
    outputs(352) <= (layer0_outputs(1503)) and not (layer0_outputs(1915));
    outputs(353) <= not((layer0_outputs(492)) or (layer0_outputs(1405)));
    outputs(354) <= (layer0_outputs(2508)) and not (layer0_outputs(2199));
    outputs(355) <= (layer0_outputs(206)) and (layer0_outputs(1037));
    outputs(356) <= layer0_outputs(350);
    outputs(357) <= not((layer0_outputs(1718)) or (layer0_outputs(1459)));
    outputs(358) <= (layer0_outputs(642)) and not (layer0_outputs(1991));
    outputs(359) <= (layer0_outputs(309)) and not (layer0_outputs(328));
    outputs(360) <= (layer0_outputs(1992)) and (layer0_outputs(649));
    outputs(361) <= (layer0_outputs(805)) and (layer0_outputs(1826));
    outputs(362) <= (layer0_outputs(393)) and (layer0_outputs(1146));
    outputs(363) <= not(layer0_outputs(35));
    outputs(364) <= (layer0_outputs(853)) and (layer0_outputs(1804));
    outputs(365) <= (layer0_outputs(1164)) and (layer0_outputs(814));
    outputs(366) <= not(layer0_outputs(932));
    outputs(367) <= (layer0_outputs(2142)) and (layer0_outputs(499));
    outputs(368) <= (layer0_outputs(962)) and (layer0_outputs(2014));
    outputs(369) <= (layer0_outputs(1892)) and not (layer0_outputs(1883));
    outputs(370) <= not((layer0_outputs(1393)) or (layer0_outputs(1506)));
    outputs(371) <= (layer0_outputs(2428)) and not (layer0_outputs(1822));
    outputs(372) <= (layer0_outputs(1232)) and not (layer0_outputs(2341));
    outputs(373) <= (layer0_outputs(692)) and (layer0_outputs(1381));
    outputs(374) <= (layer0_outputs(1239)) and (layer0_outputs(1128));
    outputs(375) <= (layer0_outputs(751)) and not (layer0_outputs(2551));
    outputs(376) <= (layer0_outputs(1767)) and not (layer0_outputs(1517));
    outputs(377) <= (layer0_outputs(743)) and (layer0_outputs(34));
    outputs(378) <= (layer0_outputs(2163)) and (layer0_outputs(922));
    outputs(379) <= (layer0_outputs(645)) and not (layer0_outputs(1163));
    outputs(380) <= (layer0_outputs(1471)) and not (layer0_outputs(2429));
    outputs(381) <= (layer0_outputs(1402)) and not (layer0_outputs(1626));
    outputs(382) <= not((layer0_outputs(1041)) or (layer0_outputs(1733)));
    outputs(383) <= not((layer0_outputs(2)) or (layer0_outputs(1173)));
    outputs(384) <= (layer0_outputs(1870)) and not (layer0_outputs(2518));
    outputs(385) <= not((layer0_outputs(2004)) or (layer0_outputs(1450)));
    outputs(386) <= (layer0_outputs(1476)) and not (layer0_outputs(1606));
    outputs(387) <= (layer0_outputs(2239)) and (layer0_outputs(672));
    outputs(388) <= (layer0_outputs(548)) and not (layer0_outputs(836));
    outputs(389) <= not((layer0_outputs(663)) or (layer0_outputs(2015)));
    outputs(390) <= (layer0_outputs(2531)) and not (layer0_outputs(530));
    outputs(391) <= not((layer0_outputs(1878)) or (layer0_outputs(27)));
    outputs(392) <= (layer0_outputs(877)) and (layer0_outputs(863));
    outputs(393) <= layer0_outputs(2254);
    outputs(394) <= not(layer0_outputs(1966));
    outputs(395) <= (layer0_outputs(855)) and (layer0_outputs(2433));
    outputs(396) <= (layer0_outputs(1042)) and (layer0_outputs(73));
    outputs(397) <= (layer0_outputs(538)) and not (layer0_outputs(1689));
    outputs(398) <= (layer0_outputs(159)) and not (layer0_outputs(1460));
    outputs(399) <= (layer0_outputs(734)) and not (layer0_outputs(286));
    outputs(400) <= not(layer0_outputs(211));
    outputs(401) <= (layer0_outputs(2151)) and (layer0_outputs(1008));
    outputs(402) <= (layer0_outputs(230)) and not (layer0_outputs(53));
    outputs(403) <= (layer0_outputs(134)) and not (layer0_outputs(619));
    outputs(404) <= '0';
    outputs(405) <= (layer0_outputs(1168)) and not (layer0_outputs(764));
    outputs(406) <= (layer0_outputs(2535)) and not (layer0_outputs(539));
    outputs(407) <= (layer0_outputs(958)) and not (layer0_outputs(1229));
    outputs(408) <= not((layer0_outputs(1789)) or (layer0_outputs(1698)));
    outputs(409) <= not((layer0_outputs(1850)) or (layer0_outputs(1067)));
    outputs(410) <= (layer0_outputs(1987)) and not (layer0_outputs(1499));
    outputs(411) <= (layer0_outputs(1151)) xor (layer0_outputs(323));
    outputs(412) <= (layer0_outputs(2026)) and not (layer0_outputs(568));
    outputs(413) <= not((layer0_outputs(235)) or (layer0_outputs(52)));
    outputs(414) <= (layer0_outputs(470)) xor (layer0_outputs(482));
    outputs(415) <= (layer0_outputs(1299)) and not (layer0_outputs(316));
    outputs(416) <= (layer0_outputs(910)) and (layer0_outputs(1780));
    outputs(417) <= (layer0_outputs(1425)) and (layer0_outputs(1971));
    outputs(418) <= layer0_outputs(2554);
    outputs(419) <= (layer0_outputs(149)) and not (layer0_outputs(140));
    outputs(420) <= (layer0_outputs(1805)) and not (layer0_outputs(600));
    outputs(421) <= not((layer0_outputs(162)) or (layer0_outputs(1062)));
    outputs(422) <= (layer0_outputs(813)) and not (layer0_outputs(43));
    outputs(423) <= (layer0_outputs(342)) and (layer0_outputs(1725));
    outputs(424) <= (layer0_outputs(2047)) and not (layer0_outputs(1040));
    outputs(425) <= layer0_outputs(0);
    outputs(426) <= (layer0_outputs(1427)) and (layer0_outputs(2542));
    outputs(427) <= (layer0_outputs(583)) and not (layer0_outputs(1337));
    outputs(428) <= (layer0_outputs(723)) and not (layer0_outputs(2432));
    outputs(429) <= (layer0_outputs(1973)) and not (layer0_outputs(1384));
    outputs(430) <= (layer0_outputs(2366)) and not (layer0_outputs(2044));
    outputs(431) <= (layer0_outputs(585)) xor (layer0_outputs(2345));
    outputs(432) <= not((layer0_outputs(1753)) or (layer0_outputs(2323)));
    outputs(433) <= '0';
    outputs(434) <= not((layer0_outputs(325)) or (layer0_outputs(522)));
    outputs(435) <= (layer0_outputs(912)) and (layer0_outputs(1495));
    outputs(436) <= not((layer0_outputs(1500)) or (layer0_outputs(2534)));
    outputs(437) <= (layer0_outputs(1957)) and (layer0_outputs(1105));
    outputs(438) <= not((layer0_outputs(1779)) or (layer0_outputs(1201)));
    outputs(439) <= (layer0_outputs(1885)) and not (layer0_outputs(436));
    outputs(440) <= not((layer0_outputs(2507)) or (layer0_outputs(271)));
    outputs(441) <= not((layer0_outputs(1300)) or (layer0_outputs(1149)));
    outputs(442) <= (layer0_outputs(862)) and not (layer0_outputs(2153));
    outputs(443) <= not((layer0_outputs(1719)) or (layer0_outputs(411)));
    outputs(444) <= not((layer0_outputs(1129)) xor (layer0_outputs(2054)));
    outputs(445) <= (layer0_outputs(1833)) and not (layer0_outputs(1175));
    outputs(446) <= not(layer0_outputs(918));
    outputs(447) <= (layer0_outputs(943)) and not (layer0_outputs(377));
    outputs(448) <= (layer0_outputs(278)) and not (layer0_outputs(368));
    outputs(449) <= (layer0_outputs(2181)) and not (layer0_outputs(1904));
    outputs(450) <= (layer0_outputs(750)) and not (layer0_outputs(504));
    outputs(451) <= not((layer0_outputs(50)) or (layer0_outputs(1547)));
    outputs(452) <= not((layer0_outputs(890)) or (layer0_outputs(1271)));
    outputs(453) <= not((layer0_outputs(40)) or (layer0_outputs(1492)));
    outputs(454) <= (layer0_outputs(1182)) and not (layer0_outputs(1904));
    outputs(455) <= (layer0_outputs(584)) and not (layer0_outputs(132));
    outputs(456) <= (layer0_outputs(1605)) and (layer0_outputs(1467));
    outputs(457) <= (layer0_outputs(665)) and not (layer0_outputs(599));
    outputs(458) <= (layer0_outputs(1611)) and not (layer0_outputs(1945));
    outputs(459) <= (layer0_outputs(420)) and not (layer0_outputs(2304));
    outputs(460) <= layer0_outputs(474);
    outputs(461) <= (layer0_outputs(2173)) and (layer0_outputs(2100));
    outputs(462) <= (layer0_outputs(1794)) and not (layer0_outputs(2109));
    outputs(463) <= layer0_outputs(2156);
    outputs(464) <= not((layer0_outputs(2265)) xor (layer0_outputs(1711)));
    outputs(465) <= (layer0_outputs(784)) and (layer0_outputs(520));
    outputs(466) <= (layer0_outputs(437)) and not (layer0_outputs(844));
    outputs(467) <= (layer0_outputs(2437)) and not (layer0_outputs(1922));
    outputs(468) <= not((layer0_outputs(2212)) or (layer0_outputs(2330)));
    outputs(469) <= layer0_outputs(1812);
    outputs(470) <= not((layer0_outputs(2524)) or (layer0_outputs(2095)));
    outputs(471) <= not((layer0_outputs(1600)) or (layer0_outputs(1852)));
    outputs(472) <= (layer0_outputs(841)) and not (layer0_outputs(2132));
    outputs(473) <= not((layer0_outputs(2377)) or (layer0_outputs(1972)));
    outputs(474) <= (layer0_outputs(2274)) and not (layer0_outputs(543));
    outputs(475) <= layer0_outputs(845);
    outputs(476) <= (layer0_outputs(382)) and not (layer0_outputs(1240));
    outputs(477) <= not((layer0_outputs(81)) or (layer0_outputs(87)));
    outputs(478) <= (layer0_outputs(1055)) and not (layer0_outputs(1679));
    outputs(479) <= not(layer0_outputs(1320));
    outputs(480) <= not((layer0_outputs(492)) or (layer0_outputs(1505)));
    outputs(481) <= (layer0_outputs(686)) and not (layer0_outputs(1110));
    outputs(482) <= not((layer0_outputs(470)) or (layer0_outputs(1953)));
    outputs(483) <= not((layer0_outputs(436)) or (layer0_outputs(2219)));
    outputs(484) <= (layer0_outputs(985)) and not (layer0_outputs(1575));
    outputs(485) <= (layer0_outputs(1097)) and (layer0_outputs(787));
    outputs(486) <= (layer0_outputs(444)) and (layer0_outputs(73));
    outputs(487) <= layer0_outputs(1187);
    outputs(488) <= (layer0_outputs(177)) and not (layer0_outputs(624));
    outputs(489) <= (layer0_outputs(2079)) and not (layer0_outputs(830));
    outputs(490) <= (layer0_outputs(255)) and (layer0_outputs(253));
    outputs(491) <= (layer0_outputs(617)) and (layer0_outputs(714));
    outputs(492) <= (layer0_outputs(634)) and not (layer0_outputs(2436));
    outputs(493) <= not((layer0_outputs(262)) or (layer0_outputs(152)));
    outputs(494) <= (layer0_outputs(159)) and not (layer0_outputs(1983));
    outputs(495) <= not(layer0_outputs(2470));
    outputs(496) <= not((layer0_outputs(938)) or (layer0_outputs(373)));
    outputs(497) <= (layer0_outputs(1973)) and (layer0_outputs(216));
    outputs(498) <= not((layer0_outputs(2537)) or (layer0_outputs(221)));
    outputs(499) <= (layer0_outputs(684)) and (layer0_outputs(2468));
    outputs(500) <= not((layer0_outputs(153)) or (layer0_outputs(568)));
    outputs(501) <= (layer0_outputs(2394)) and (layer0_outputs(901));
    outputs(502) <= '0';
    outputs(503) <= not((layer0_outputs(1748)) or (layer0_outputs(1572)));
    outputs(504) <= (layer0_outputs(2287)) and not (layer0_outputs(1003));
    outputs(505) <= (layer0_outputs(98)) and not (layer0_outputs(1895));
    outputs(506) <= not((layer0_outputs(690)) or (layer0_outputs(2532)));
    outputs(507) <= (layer0_outputs(2501)) and not (layer0_outputs(1259));
    outputs(508) <= (layer0_outputs(605)) and (layer0_outputs(1578));
    outputs(509) <= (layer0_outputs(1166)) and not (layer0_outputs(2313));
    outputs(510) <= not((layer0_outputs(319)) or (layer0_outputs(1940)));
    outputs(511) <= (layer0_outputs(576)) and (layer0_outputs(867));
    outputs(512) <= not((layer0_outputs(2240)) or (layer0_outputs(2065)));
    outputs(513) <= not((layer0_outputs(3)) xor (layer0_outputs(362)));
    outputs(514) <= not((layer0_outputs(705)) xor (layer0_outputs(1532)));
    outputs(515) <= layer0_outputs(1432);
    outputs(516) <= not(layer0_outputs(471)) or (layer0_outputs(479));
    outputs(517) <= layer0_outputs(1080);
    outputs(518) <= not((layer0_outputs(1793)) and (layer0_outputs(1594)));
    outputs(519) <= layer0_outputs(572);
    outputs(520) <= not(layer0_outputs(445));
    outputs(521) <= (layer0_outputs(491)) or (layer0_outputs(1035));
    outputs(522) <= layer0_outputs(229);
    outputs(523) <= not(layer0_outputs(19));
    outputs(524) <= layer0_outputs(2524);
    outputs(525) <= not((layer0_outputs(1685)) and (layer0_outputs(2328)));
    outputs(526) <= not(layer0_outputs(276));
    outputs(527) <= not(layer0_outputs(2518));
    outputs(528) <= not(layer0_outputs(1885)) or (layer0_outputs(1303));
    outputs(529) <= (layer0_outputs(1053)) and (layer0_outputs(363));
    outputs(530) <= (layer0_outputs(1981)) and not (layer0_outputs(2077));
    outputs(531) <= not((layer0_outputs(191)) and (layer0_outputs(1631)));
    outputs(532) <= not((layer0_outputs(541)) or (layer0_outputs(1439)));
    outputs(533) <= layer0_outputs(1424);
    outputs(534) <= not(layer0_outputs(1092));
    outputs(535) <= not(layer0_outputs(1745));
    outputs(536) <= not((layer0_outputs(2272)) and (layer0_outputs(2211)));
    outputs(537) <= not(layer0_outputs(135));
    outputs(538) <= not((layer0_outputs(2469)) or (layer0_outputs(1261)));
    outputs(539) <= layer0_outputs(2338);
    outputs(540) <= layer0_outputs(70);
    outputs(541) <= layer0_outputs(1866);
    outputs(542) <= layer0_outputs(696);
    outputs(543) <= not(layer0_outputs(1044));
    outputs(544) <= layer0_outputs(1753);
    outputs(545) <= not(layer0_outputs(289)) or (layer0_outputs(2130));
    outputs(546) <= not(layer0_outputs(2097)) or (layer0_outputs(322));
    outputs(547) <= not((layer0_outputs(1265)) xor (layer0_outputs(1082)));
    outputs(548) <= not(layer0_outputs(473));
    outputs(549) <= (layer0_outputs(1533)) and not (layer0_outputs(575));
    outputs(550) <= not(layer0_outputs(2089)) or (layer0_outputs(1897));
    outputs(551) <= not((layer0_outputs(1556)) and (layer0_outputs(2321)));
    outputs(552) <= layer0_outputs(2131);
    outputs(553) <= not((layer0_outputs(2495)) and (layer0_outputs(1517)));
    outputs(554) <= not(layer0_outputs(172));
    outputs(555) <= (layer0_outputs(422)) and (layer0_outputs(595));
    outputs(556) <= layer0_outputs(746);
    outputs(557) <= (layer0_outputs(2276)) and not (layer0_outputs(581));
    outputs(558) <= not(layer0_outputs(42)) or (layer0_outputs(350));
    outputs(559) <= (layer0_outputs(1097)) and (layer0_outputs(670));
    outputs(560) <= not(layer0_outputs(2389)) or (layer0_outputs(2034));
    outputs(561) <= not(layer0_outputs(2318));
    outputs(562) <= (layer0_outputs(2239)) and (layer0_outputs(2223));
    outputs(563) <= not(layer0_outputs(30)) or (layer0_outputs(617));
    outputs(564) <= not((layer0_outputs(1576)) xor (layer0_outputs(1592)));
    outputs(565) <= not(layer0_outputs(1843));
    outputs(566) <= not(layer0_outputs(1410));
    outputs(567) <= not(layer0_outputs(285)) or (layer0_outputs(1653));
    outputs(568) <= not(layer0_outputs(472));
    outputs(569) <= (layer0_outputs(970)) and (layer0_outputs(1889));
    outputs(570) <= not((layer0_outputs(1684)) xor (layer0_outputs(185)));
    outputs(571) <= not((layer0_outputs(2430)) xor (layer0_outputs(2061)));
    outputs(572) <= layer0_outputs(1137);
    outputs(573) <= not((layer0_outputs(1679)) or (layer0_outputs(2273)));
    outputs(574) <= (layer0_outputs(644)) or (layer0_outputs(739));
    outputs(575) <= (layer0_outputs(896)) and (layer0_outputs(1848));
    outputs(576) <= layer0_outputs(2310);
    outputs(577) <= layer0_outputs(542);
    outputs(578) <= not((layer0_outputs(842)) xor (layer0_outputs(2353)));
    outputs(579) <= not((layer0_outputs(843)) xor (layer0_outputs(2396)));
    outputs(580) <= not(layer0_outputs(1215)) or (layer0_outputs(1157));
    outputs(581) <= not(layer0_outputs(1027));
    outputs(582) <= (layer0_outputs(1659)) and (layer0_outputs(902));
    outputs(583) <= not(layer0_outputs(1656));
    outputs(584) <= layer0_outputs(1262);
    outputs(585) <= not(layer0_outputs(2538));
    outputs(586) <= not(layer0_outputs(55)) or (layer0_outputs(619));
    outputs(587) <= not((layer0_outputs(2290)) or (layer0_outputs(1536)));
    outputs(588) <= not(layer0_outputs(505)) or (layer0_outputs(1364));
    outputs(589) <= not(layer0_outputs(1573));
    outputs(590) <= not(layer0_outputs(324)) or (layer0_outputs(2465));
    outputs(591) <= not(layer0_outputs(1243));
    outputs(592) <= not(layer0_outputs(2041));
    outputs(593) <= not((layer0_outputs(2122)) or (layer0_outputs(700)));
    outputs(594) <= layer0_outputs(1213);
    outputs(595) <= not((layer0_outputs(598)) and (layer0_outputs(972)));
    outputs(596) <= layer0_outputs(727);
    outputs(597) <= not(layer0_outputs(1207));
    outputs(598) <= (layer0_outputs(1913)) or (layer0_outputs(354));
    outputs(599) <= layer0_outputs(528);
    outputs(600) <= not(layer0_outputs(770));
    outputs(601) <= not(layer0_outputs(424)) or (layer0_outputs(2509));
    outputs(602) <= (layer0_outputs(530)) and not (layer0_outputs(493));
    outputs(603) <= layer0_outputs(160);
    outputs(604) <= not(layer0_outputs(1989)) or (layer0_outputs(330));
    outputs(605) <= not(layer0_outputs(1530)) or (layer0_outputs(2129));
    outputs(606) <= (layer0_outputs(1784)) and (layer0_outputs(2351));
    outputs(607) <= layer0_outputs(48);
    outputs(608) <= not(layer0_outputs(1186));
    outputs(609) <= layer0_outputs(116);
    outputs(610) <= not(layer0_outputs(685));
    outputs(611) <= not((layer0_outputs(975)) or (layer0_outputs(1642)));
    outputs(612) <= not(layer0_outputs(975));
    outputs(613) <= not(layer0_outputs(1649)) or (layer0_outputs(2034));
    outputs(614) <= not(layer0_outputs(1950));
    outputs(615) <= not(layer0_outputs(1636)) or (layer0_outputs(1030));
    outputs(616) <= layer0_outputs(279);
    outputs(617) <= not((layer0_outputs(132)) or (layer0_outputs(544)));
    outputs(618) <= not(layer0_outputs(2119));
    outputs(619) <= not((layer0_outputs(526)) and (layer0_outputs(1302)));
    outputs(620) <= not(layer0_outputs(2393)) or (layer0_outputs(251));
    outputs(621) <= (layer0_outputs(657)) and (layer0_outputs(458));
    outputs(622) <= not(layer0_outputs(1971));
    outputs(623) <= not(layer0_outputs(236));
    outputs(624) <= layer0_outputs(1701);
    outputs(625) <= (layer0_outputs(1440)) or (layer0_outputs(1862));
    outputs(626) <= not(layer0_outputs(2098)) or (layer0_outputs(836));
    outputs(627) <= not(layer0_outputs(1348));
    outputs(628) <= not((layer0_outputs(1756)) xor (layer0_outputs(1467)));
    outputs(629) <= not((layer0_outputs(1802)) xor (layer0_outputs(1511)));
    outputs(630) <= not(layer0_outputs(26));
    outputs(631) <= not(layer0_outputs(133));
    outputs(632) <= not(layer0_outputs(2441)) or (layer0_outputs(1813));
    outputs(633) <= (layer0_outputs(2337)) and not (layer0_outputs(2169));
    outputs(634) <= (layer0_outputs(589)) and not (layer0_outputs(824));
    outputs(635) <= not(layer0_outputs(1312));
    outputs(636) <= not(layer0_outputs(402));
    outputs(637) <= not((layer0_outputs(881)) or (layer0_outputs(1937)));
    outputs(638) <= not(layer0_outputs(1832)) or (layer0_outputs(746));
    outputs(639) <= layer0_outputs(122);
    outputs(640) <= (layer0_outputs(46)) and (layer0_outputs(2338));
    outputs(641) <= not(layer0_outputs(1033));
    outputs(642) <= layer0_outputs(548);
    outputs(643) <= (layer0_outputs(1195)) and not (layer0_outputs(212));
    outputs(644) <= layer0_outputs(1682);
    outputs(645) <= layer0_outputs(2213);
    outputs(646) <= not((layer0_outputs(926)) and (layer0_outputs(1955)));
    outputs(647) <= not(layer0_outputs(1951));
    outputs(648) <= (layer0_outputs(668)) xor (layer0_outputs(1609));
    outputs(649) <= layer0_outputs(509);
    outputs(650) <= (layer0_outputs(1695)) and (layer0_outputs(279));
    outputs(651) <= not(layer0_outputs(161)) or (layer0_outputs(2527));
    outputs(652) <= not(layer0_outputs(2368)) or (layer0_outputs(2133));
    outputs(653) <= not(layer0_outputs(1161));
    outputs(654) <= layer0_outputs(1390);
    outputs(655) <= not((layer0_outputs(1844)) or (layer0_outputs(1256)));
    outputs(656) <= (layer0_outputs(494)) and not (layer0_outputs(1224));
    outputs(657) <= not(layer0_outputs(631)) or (layer0_outputs(1309));
    outputs(658) <= layer0_outputs(1617);
    outputs(659) <= not(layer0_outputs(1282));
    outputs(660) <= (layer0_outputs(1657)) and not (layer0_outputs(955));
    outputs(661) <= not((layer0_outputs(1554)) and (layer0_outputs(1863)));
    outputs(662) <= (layer0_outputs(138)) and not (layer0_outputs(2145));
    outputs(663) <= not(layer0_outputs(467)) or (layer0_outputs(889));
    outputs(664) <= not(layer0_outputs(2426)) or (layer0_outputs(1740));
    outputs(665) <= (layer0_outputs(2164)) and not (layer0_outputs(1383));
    outputs(666) <= layer0_outputs(730);
    outputs(667) <= (layer0_outputs(1113)) xor (layer0_outputs(1777));
    outputs(668) <= layer0_outputs(417);
    outputs(669) <= layer0_outputs(739);
    outputs(670) <= not(layer0_outputs(1871));
    outputs(671) <= (layer0_outputs(607)) and not (layer0_outputs(808));
    outputs(672) <= (layer0_outputs(2447)) or (layer0_outputs(2365));
    outputs(673) <= not(layer0_outputs(2008)) or (layer0_outputs(2201));
    outputs(674) <= not(layer0_outputs(630));
    outputs(675) <= not(layer0_outputs(2005));
    outputs(676) <= (layer0_outputs(839)) and not (layer0_outputs(1231));
    outputs(677) <= not(layer0_outputs(217));
    outputs(678) <= not(layer0_outputs(1526)) or (layer0_outputs(1417));
    outputs(679) <= layer0_outputs(726);
    outputs(680) <= not((layer0_outputs(2479)) xor (layer0_outputs(632)));
    outputs(681) <= (layer0_outputs(2087)) xor (layer0_outputs(983));
    outputs(682) <= (layer0_outputs(1111)) and not (layer0_outputs(576));
    outputs(683) <= layer0_outputs(1210);
    outputs(684) <= layer0_outputs(1174);
    outputs(685) <= layer0_outputs(2110);
    outputs(686) <= (layer0_outputs(1644)) or (layer0_outputs(1028));
    outputs(687) <= not(layer0_outputs(341));
    outputs(688) <= layer0_outputs(2348);
    outputs(689) <= (layer0_outputs(2347)) or (layer0_outputs(186));
    outputs(690) <= layer0_outputs(716);
    outputs(691) <= layer0_outputs(420);
    outputs(692) <= not((layer0_outputs(77)) xor (layer0_outputs(1172)));
    outputs(693) <= not(layer0_outputs(916));
    outputs(694) <= (layer0_outputs(1305)) and not (layer0_outputs(300));
    outputs(695) <= (layer0_outputs(439)) or (layer0_outputs(993));
    outputs(696) <= not(layer0_outputs(807));
    outputs(697) <= not((layer0_outputs(1469)) xor (layer0_outputs(791)));
    outputs(698) <= not(layer0_outputs(284));
    outputs(699) <= not(layer0_outputs(1596)) or (layer0_outputs(555));
    outputs(700) <= not(layer0_outputs(390)) or (layer0_outputs(797));
    outputs(701) <= (layer0_outputs(2298)) and (layer0_outputs(832));
    outputs(702) <= (layer0_outputs(1743)) xor (layer0_outputs(2155));
    outputs(703) <= not(layer0_outputs(810));
    outputs(704) <= layer0_outputs(405);
    outputs(705) <= layer0_outputs(1136);
    outputs(706) <= not(layer0_outputs(217));
    outputs(707) <= not(layer0_outputs(155)) or (layer0_outputs(872));
    outputs(708) <= not((layer0_outputs(2233)) xor (layer0_outputs(1346)));
    outputs(709) <= not(layer0_outputs(99)) or (layer0_outputs(2064));
    outputs(710) <= (layer0_outputs(2176)) or (layer0_outputs(1163));
    outputs(711) <= (layer0_outputs(1724)) or (layer0_outputs(1949));
    outputs(712) <= layer0_outputs(2536);
    outputs(713) <= not(layer0_outputs(275));
    outputs(714) <= not(layer0_outputs(2118)) or (layer0_outputs(28));
    outputs(715) <= (layer0_outputs(2464)) and not (layer0_outputs(773));
    outputs(716) <= not((layer0_outputs(161)) and (layer0_outputs(676)));
    outputs(717) <= not((layer0_outputs(1287)) or (layer0_outputs(865)));
    outputs(718) <= not((layer0_outputs(281)) and (layer0_outputs(2452)));
    outputs(719) <= not(layer0_outputs(1228)) or (layer0_outputs(1948));
    outputs(720) <= not(layer0_outputs(2303)) or (layer0_outputs(387));
    outputs(721) <= not(layer0_outputs(1215)) or (layer0_outputs(946));
    outputs(722) <= not(layer0_outputs(1970));
    outputs(723) <= not((layer0_outputs(2284)) or (layer0_outputs(188)));
    outputs(724) <= layer0_outputs(260);
    outputs(725) <= not(layer0_outputs(920));
    outputs(726) <= not(layer0_outputs(264)) or (layer0_outputs(178));
    outputs(727) <= layer0_outputs(1277);
    outputs(728) <= layer0_outputs(2143);
    outputs(729) <= not(layer0_outputs(2342)) or (layer0_outputs(384));
    outputs(730) <= (layer0_outputs(2362)) and (layer0_outputs(15));
    outputs(731) <= layer0_outputs(830);
    outputs(732) <= layer0_outputs(2515);
    outputs(733) <= not(layer0_outputs(1318));
    outputs(734) <= layer0_outputs(597);
    outputs(735) <= not(layer0_outputs(812)) or (layer0_outputs(260));
    outputs(736) <= not(layer0_outputs(1962)) or (layer0_outputs(286));
    outputs(737) <= not(layer0_outputs(1563)) or (layer0_outputs(772));
    outputs(738) <= (layer0_outputs(618)) and not (layer0_outputs(1908));
    outputs(739) <= layer0_outputs(422);
    outputs(740) <= not(layer0_outputs(2159)) or (layer0_outputs(1758));
    outputs(741) <= (layer0_outputs(2045)) and not (layer0_outputs(1438));
    outputs(742) <= layer0_outputs(923);
    outputs(743) <= not((layer0_outputs(1081)) and (layer0_outputs(1645)));
    outputs(744) <= layer0_outputs(123);
    outputs(745) <= not(layer0_outputs(2166));
    outputs(746) <= layer0_outputs(233);
    outputs(747) <= (layer0_outputs(1850)) or (layer0_outputs(2078));
    outputs(748) <= (layer0_outputs(211)) xor (layer0_outputs(1469));
    outputs(749) <= not(layer0_outputs(2441));
    outputs(750) <= layer0_outputs(560);
    outputs(751) <= not(layer0_outputs(536));
    outputs(752) <= not((layer0_outputs(1134)) xor (layer0_outputs(512)));
    outputs(753) <= (layer0_outputs(1220)) xor (layer0_outputs(2412));
    outputs(754) <= not((layer0_outputs(1939)) xor (layer0_outputs(1696)));
    outputs(755) <= layer0_outputs(122);
    outputs(756) <= (layer0_outputs(1778)) or (layer0_outputs(2463));
    outputs(757) <= not(layer0_outputs(2426));
    outputs(758) <= layer0_outputs(1377);
    outputs(759) <= not(layer0_outputs(1927));
    outputs(760) <= layer0_outputs(1829);
    outputs(761) <= not(layer0_outputs(695));
    outputs(762) <= (layer0_outputs(57)) or (layer0_outputs(1112));
    outputs(763) <= not(layer0_outputs(2075));
    outputs(764) <= not(layer0_outputs(788));
    outputs(765) <= not((layer0_outputs(1693)) and (layer0_outputs(2437)));
    outputs(766) <= layer0_outputs(1963);
    outputs(767) <= layer0_outputs(677);
    outputs(768) <= not(layer0_outputs(2326)) or (layer0_outputs(593));
    outputs(769) <= (layer0_outputs(1799)) and not (layer0_outputs(758));
    outputs(770) <= (layer0_outputs(264)) and (layer0_outputs(1637));
    outputs(771) <= not(layer0_outputs(1678));
    outputs(772) <= not((layer0_outputs(503)) xor (layer0_outputs(2167)));
    outputs(773) <= not(layer0_outputs(823)) or (layer0_outputs(293));
    outputs(774) <= not(layer0_outputs(1851));
    outputs(775) <= not(layer0_outputs(881));
    outputs(776) <= not((layer0_outputs(590)) or (layer0_outputs(1175)));
    outputs(777) <= not((layer0_outputs(2439)) and (layer0_outputs(1584)));
    outputs(778) <= (layer0_outputs(365)) and (layer0_outputs(2180));
    outputs(779) <= (layer0_outputs(1038)) and (layer0_outputs(498));
    outputs(780) <= not(layer0_outputs(935));
    outputs(781) <= layer0_outputs(41);
    outputs(782) <= (layer0_outputs(2340)) and not (layer0_outputs(1663));
    outputs(783) <= not(layer0_outputs(763));
    outputs(784) <= layer0_outputs(858);
    outputs(785) <= not((layer0_outputs(1810)) or (layer0_outputs(2207)));
    outputs(786) <= (layer0_outputs(59)) and not (layer0_outputs(1874));
    outputs(787) <= layer0_outputs(2287);
    outputs(788) <= (layer0_outputs(1587)) and not (layer0_outputs(954));
    outputs(789) <= (layer0_outputs(465)) and not (layer0_outputs(171));
    outputs(790) <= not((layer0_outputs(1963)) xor (layer0_outputs(1833)));
    outputs(791) <= not(layer0_outputs(118));
    outputs(792) <= not(layer0_outputs(1566));
    outputs(793) <= (layer0_outputs(1410)) and not (layer0_outputs(1423));
    outputs(794) <= not((layer0_outputs(2140)) or (layer0_outputs(543)));
    outputs(795) <= not((layer0_outputs(1031)) or (layer0_outputs(179)));
    outputs(796) <= (layer0_outputs(1911)) or (layer0_outputs(1660));
    outputs(797) <= not((layer0_outputs(984)) or (layer0_outputs(348)));
    outputs(798) <= layer0_outputs(1588);
    outputs(799) <= (layer0_outputs(2357)) and not (layer0_outputs(635));
    outputs(800) <= not(layer0_outputs(1372));
    outputs(801) <= layer0_outputs(607);
    outputs(802) <= not(layer0_outputs(1258));
    outputs(803) <= (layer0_outputs(234)) and not (layer0_outputs(1135));
    outputs(804) <= not((layer0_outputs(2148)) or (layer0_outputs(2249)));
    outputs(805) <= layer0_outputs(2391);
    outputs(806) <= not(layer0_outputs(2031)) or (layer0_outputs(209));
    outputs(807) <= not((layer0_outputs(2252)) or (layer0_outputs(1367)));
    outputs(808) <= not(layer0_outputs(1750)) or (layer0_outputs(2301));
    outputs(809) <= not(layer0_outputs(1570));
    outputs(810) <= layer0_outputs(2417);
    outputs(811) <= (layer0_outputs(928)) and not (layer0_outputs(402));
    outputs(812) <= (layer0_outputs(1729)) or (layer0_outputs(994));
    outputs(813) <= not(layer0_outputs(440));
    outputs(814) <= layer0_outputs(1264);
    outputs(815) <= not((layer0_outputs(38)) or (layer0_outputs(2259)));
    outputs(816) <= not(layer0_outputs(2392));
    outputs(817) <= (layer0_outputs(1628)) and not (layer0_outputs(1800));
    outputs(818) <= not(layer0_outputs(255));
    outputs(819) <= not(layer0_outputs(662));
    outputs(820) <= not(layer0_outputs(2352));
    outputs(821) <= not(layer0_outputs(2457));
    outputs(822) <= (layer0_outputs(1389)) and not (layer0_outputs(1121));
    outputs(823) <= not((layer0_outputs(810)) or (layer0_outputs(2477)));
    outputs(824) <= layer0_outputs(453);
    outputs(825) <= (layer0_outputs(824)) and not (layer0_outputs(1813));
    outputs(826) <= not((layer0_outputs(1733)) xor (layer0_outputs(465)));
    outputs(827) <= layer0_outputs(2020);
    outputs(828) <= not(layer0_outputs(2399));
    outputs(829) <= (layer0_outputs(1351)) or (layer0_outputs(1779));
    outputs(830) <= (layer0_outputs(757)) and not (layer0_outputs(784));
    outputs(831) <= (layer0_outputs(1010)) and (layer0_outputs(268));
    outputs(832) <= not(layer0_outputs(1129));
    outputs(833) <= not((layer0_outputs(1400)) or (layer0_outputs(2158)));
    outputs(834) <= (layer0_outputs(488)) and (layer0_outputs(1330));
    outputs(835) <= (layer0_outputs(2360)) and not (layer0_outputs(766));
    outputs(836) <= layer0_outputs(1068);
    outputs(837) <= (layer0_outputs(1394)) and (layer0_outputs(2540));
    outputs(838) <= (layer0_outputs(2063)) and (layer0_outputs(2528));
    outputs(839) <= layer0_outputs(1956);
    outputs(840) <= (layer0_outputs(181)) or (layer0_outputs(2152));
    outputs(841) <= not(layer0_outputs(1362));
    outputs(842) <= (layer0_outputs(1934)) and not (layer0_outputs(1363));
    outputs(843) <= not((layer0_outputs(1380)) xor (layer0_outputs(51)));
    outputs(844) <= layer0_outputs(2162);
    outputs(845) <= (layer0_outputs(925)) xor (layer0_outputs(2532));
    outputs(846) <= layer0_outputs(1267);
    outputs(847) <= not(layer0_outputs(2112));
    outputs(848) <= layer0_outputs(2291);
    outputs(849) <= (layer0_outputs(736)) and not (layer0_outputs(1060));
    outputs(850) <= not(layer0_outputs(2290));
    outputs(851) <= not(layer0_outputs(91)) or (layer0_outputs(1795));
    outputs(852) <= layer0_outputs(1131);
    outputs(853) <= not((layer0_outputs(1807)) and (layer0_outputs(652)));
    outputs(854) <= not(layer0_outputs(1662)) or (layer0_outputs(623));
    outputs(855) <= not((layer0_outputs(2001)) or (layer0_outputs(89)));
    outputs(856) <= not(layer0_outputs(2006));
    outputs(857) <= not(layer0_outputs(2353)) or (layer0_outputs(2548));
    outputs(858) <= layer0_outputs(248);
    outputs(859) <= (layer0_outputs(2071)) and not (layer0_outputs(433));
    outputs(860) <= layer0_outputs(1253);
    outputs(861) <= (layer0_outputs(2050)) and not (layer0_outputs(2043));
    outputs(862) <= not(layer0_outputs(546));
    outputs(863) <= layer0_outputs(1088);
    outputs(864) <= not((layer0_outputs(1119)) or (layer0_outputs(1231)));
    outputs(865) <= layer0_outputs(2166);
    outputs(866) <= not(layer0_outputs(1360));
    outputs(867) <= (layer0_outputs(2453)) and not (layer0_outputs(1838));
    outputs(868) <= (layer0_outputs(814)) and not (layer0_outputs(1032));
    outputs(869) <= not(layer0_outputs(173));
    outputs(870) <= (layer0_outputs(314)) and not (layer0_outputs(1192));
    outputs(871) <= not(layer0_outputs(2400));
    outputs(872) <= layer0_outputs(2193);
    outputs(873) <= layer0_outputs(724);
    outputs(874) <= not(layer0_outputs(1849));
    outputs(875) <= layer0_outputs(2307);
    outputs(876) <= (layer0_outputs(2106)) and (layer0_outputs(435));
    outputs(877) <= not((layer0_outputs(1558)) or (layer0_outputs(2460)));
    outputs(878) <= not(layer0_outputs(67));
    outputs(879) <= (layer0_outputs(1274)) xor (layer0_outputs(2480));
    outputs(880) <= (layer0_outputs(1524)) and not (layer0_outputs(909));
    outputs(881) <= not(layer0_outputs(456));
    outputs(882) <= (layer0_outputs(169)) and (layer0_outputs(2325));
    outputs(883) <= (layer0_outputs(287)) and not (layer0_outputs(2021));
    outputs(884) <= layer0_outputs(1463);
    outputs(885) <= not((layer0_outputs(775)) and (layer0_outputs(2541)));
    outputs(886) <= (layer0_outputs(1452)) and (layer0_outputs(828));
    outputs(887) <= not(layer0_outputs(5));
    outputs(888) <= layer0_outputs(16);
    outputs(889) <= not(layer0_outputs(2308));
    outputs(890) <= not(layer0_outputs(130));
    outputs(891) <= not(layer0_outputs(1612));
    outputs(892) <= not(layer0_outputs(1497));
    outputs(893) <= layer0_outputs(2466);
    outputs(894) <= not((layer0_outputs(243)) or (layer0_outputs(68)));
    outputs(895) <= not((layer0_outputs(925)) or (layer0_outputs(1126)));
    outputs(896) <= not((layer0_outputs(2364)) or (layer0_outputs(1537)));
    outputs(897) <= not(layer0_outputs(1860)) or (layer0_outputs(578));
    outputs(898) <= not(layer0_outputs(2192));
    outputs(899) <= not(layer0_outputs(1823)) or (layer0_outputs(452));
    outputs(900) <= (layer0_outputs(529)) and not (layer0_outputs(1520));
    outputs(901) <= (layer0_outputs(1839)) and not (layer0_outputs(2378));
    outputs(902) <= (layer0_outputs(332)) and (layer0_outputs(1601));
    outputs(903) <= not(layer0_outputs(1402)) or (layer0_outputs(1739));
    outputs(904) <= (layer0_outputs(1888)) and not (layer0_outputs(239));
    outputs(905) <= not(layer0_outputs(2374)) or (layer0_outputs(2012));
    outputs(906) <= not(layer0_outputs(438));
    outputs(907) <= layer0_outputs(1373);
    outputs(908) <= not(layer0_outputs(1061));
    outputs(909) <= (layer0_outputs(223)) and not (layer0_outputs(2236));
    outputs(910) <= layer0_outputs(2514);
    outputs(911) <= layer0_outputs(755);
    outputs(912) <= not((layer0_outputs(2056)) and (layer0_outputs(969)));
    outputs(913) <= (layer0_outputs(1226)) and not (layer0_outputs(351));
    outputs(914) <= not((layer0_outputs(1421)) and (layer0_outputs(1504)));
    outputs(915) <= not(layer0_outputs(1276));
    outputs(916) <= not(layer0_outputs(707));
    outputs(917) <= (layer0_outputs(1464)) and not (layer0_outputs(652));
    outputs(918) <= (layer0_outputs(1375)) and not (layer0_outputs(2259));
    outputs(919) <= (layer0_outputs(495)) and not (layer0_outputs(2249));
    outputs(920) <= not((layer0_outputs(1340)) xor (layer0_outputs(1230)));
    outputs(921) <= (layer0_outputs(854)) and not (layer0_outputs(732));
    outputs(922) <= not(layer0_outputs(476));
    outputs(923) <= not((layer0_outputs(1404)) and (layer0_outputs(1477)));
    outputs(924) <= (layer0_outputs(854)) and (layer0_outputs(1123));
    outputs(925) <= not(layer0_outputs(1887)) or (layer0_outputs(2438));
    outputs(926) <= not(layer0_outputs(737));
    outputs(927) <= not((layer0_outputs(2218)) and (layer0_outputs(610)));
    outputs(928) <= (layer0_outputs(2470)) and (layer0_outputs(2546));
    outputs(929) <= (layer0_outputs(2282)) xor (layer0_outputs(2435));
    outputs(930) <= (layer0_outputs(599)) and not (layer0_outputs(416));
    outputs(931) <= (layer0_outputs(628)) and not (layer0_outputs(425));
    outputs(932) <= not((layer0_outputs(1841)) and (layer0_outputs(289)));
    outputs(933) <= layer0_outputs(1373);
    outputs(934) <= (layer0_outputs(2516)) xor (layer0_outputs(1518));
    outputs(935) <= (layer0_outputs(552)) and (layer0_outputs(2169));
    outputs(936) <= (layer0_outputs(169)) and not (layer0_outputs(2088));
    outputs(937) <= not((layer0_outputs(2227)) and (layer0_outputs(1597)));
    outputs(938) <= (layer0_outputs(1009)) and not (layer0_outputs(218));
    outputs(939) <= (layer0_outputs(1394)) and not (layer0_outputs(1154));
    outputs(940) <= (layer0_outputs(443)) and (layer0_outputs(1150));
    outputs(941) <= layer0_outputs(349);
    outputs(942) <= not((layer0_outputs(2418)) and (layer0_outputs(222)));
    outputs(943) <= layer0_outputs(1636);
    outputs(944) <= layer0_outputs(2533);
    outputs(945) <= not(layer0_outputs(754));
    outputs(946) <= not(layer0_outputs(1477)) or (layer0_outputs(1760));
    outputs(947) <= (layer0_outputs(569)) and (layer0_outputs(1260));
    outputs(948) <= not((layer0_outputs(1198)) or (layer0_outputs(252)));
    outputs(949) <= (layer0_outputs(573)) and not (layer0_outputs(1317));
    outputs(950) <= not(layer0_outputs(753)) or (layer0_outputs(1940));
    outputs(951) <= not(layer0_outputs(734));
    outputs(952) <= layer0_outputs(1464);
    outputs(953) <= layer0_outputs(1225);
    outputs(954) <= not((layer0_outputs(633)) or (layer0_outputs(1015)));
    outputs(955) <= not(layer0_outputs(1542));
    outputs(956) <= not(layer0_outputs(708));
    outputs(957) <= (layer0_outputs(1266)) or (layer0_outputs(735));
    outputs(958) <= layer0_outputs(236);
    outputs(959) <= (layer0_outputs(1446)) and not (layer0_outputs(1475));
    outputs(960) <= not(layer0_outputs(1304));
    outputs(961) <= layer0_outputs(2502);
    outputs(962) <= (layer0_outputs(1338)) and (layer0_outputs(839));
    outputs(963) <= not(layer0_outputs(2140));
    outputs(964) <= (layer0_outputs(1711)) and not (layer0_outputs(1752));
    outputs(965) <= not((layer0_outputs(2545)) or (layer0_outputs(1460)));
    outputs(966) <= layer0_outputs(2487);
    outputs(967) <= not(layer0_outputs(1017));
    outputs(968) <= not(layer0_outputs(2064));
    outputs(969) <= not((layer0_outputs(2148)) or (layer0_outputs(1806)));
    outputs(970) <= not(layer0_outputs(2048));
    outputs(971) <= not((layer0_outputs(506)) or (layer0_outputs(1755)));
    outputs(972) <= not((layer0_outputs(399)) or (layer0_outputs(450)));
    outputs(973) <= layer0_outputs(7);
    outputs(974) <= not(layer0_outputs(224));
    outputs(975) <= (layer0_outputs(2225)) and (layer0_outputs(2345));
    outputs(976) <= (layer0_outputs(932)) and not (layer0_outputs(2288));
    outputs(977) <= (layer0_outputs(1357)) and (layer0_outputs(1671));
    outputs(978) <= layer0_outputs(797);
    outputs(979) <= not(layer0_outputs(909));
    outputs(980) <= layer0_outputs(1254);
    outputs(981) <= not(layer0_outputs(1339));
    outputs(982) <= (layer0_outputs(1353)) and not (layer0_outputs(1708));
    outputs(983) <= (layer0_outputs(569)) and not (layer0_outputs(2236));
    outputs(984) <= not(layer0_outputs(1304));
    outputs(985) <= not(layer0_outputs(1126));
    outputs(986) <= not((layer0_outputs(728)) or (layer0_outputs(1621)));
    outputs(987) <= (layer0_outputs(965)) and not (layer0_outputs(2030));
    outputs(988) <= (layer0_outputs(2138)) and not (layer0_outputs(1244));
    outputs(989) <= not(layer0_outputs(133));
    outputs(990) <= layer0_outputs(2332);
    outputs(991) <= layer0_outputs(1204);
    outputs(992) <= layer0_outputs(637);
    outputs(993) <= not(layer0_outputs(1283)) or (layer0_outputs(1378));
    outputs(994) <= (layer0_outputs(1819)) and not (layer0_outputs(2485));
    outputs(995) <= not(layer0_outputs(459));
    outputs(996) <= not((layer0_outputs(2494)) or (layer0_outputs(2074)));
    outputs(997) <= not(layer0_outputs(2278));
    outputs(998) <= layer0_outputs(2504);
    outputs(999) <= not(layer0_outputs(2397));
    outputs(1000) <= not(layer0_outputs(292));
    outputs(1001) <= not((layer0_outputs(295)) and (layer0_outputs(1515)));
    outputs(1002) <= not(layer0_outputs(2350));
    outputs(1003) <= not((layer0_outputs(269)) or (layer0_outputs(58)));
    outputs(1004) <= not(layer0_outputs(1629));
    outputs(1005) <= layer0_outputs(959);
    outputs(1006) <= not((layer0_outputs(102)) or (layer0_outputs(445)));
    outputs(1007) <= (layer0_outputs(793)) and (layer0_outputs(1029));
    outputs(1008) <= not(layer0_outputs(89));
    outputs(1009) <= (layer0_outputs(1073)) and not (layer0_outputs(1639));
    outputs(1010) <= layer0_outputs(1480);
    outputs(1011) <= not((layer0_outputs(1279)) xor (layer0_outputs(2107)));
    outputs(1012) <= layer0_outputs(1507);
    outputs(1013) <= not((layer0_outputs(1639)) or (layer0_outputs(579)));
    outputs(1014) <= not(layer0_outputs(2476));
    outputs(1015) <= (layer0_outputs(1044)) or (layer0_outputs(977));
    outputs(1016) <= not(layer0_outputs(2085));
    outputs(1017) <= (layer0_outputs(2067)) and (layer0_outputs(1675));
    outputs(1018) <= layer0_outputs(1040);
    outputs(1019) <= (layer0_outputs(1330)) and (layer0_outputs(1052));
    outputs(1020) <= layer0_outputs(432);
    outputs(1021) <= layer0_outputs(2012);
    outputs(1022) <= not(layer0_outputs(2028));
    outputs(1023) <= (layer0_outputs(2499)) and (layer0_outputs(16));
    outputs(1024) <= not(layer0_outputs(749));
    outputs(1025) <= (layer0_outputs(1365)) and not (layer0_outputs(70));
    outputs(1026) <= not((layer0_outputs(848)) or (layer0_outputs(339)));
    outputs(1027) <= not((layer0_outputs(1757)) and (layer0_outputs(558)));
    outputs(1028) <= not(layer0_outputs(928));
    outputs(1029) <= layer0_outputs(2023);
    outputs(1030) <= not(layer0_outputs(24));
    outputs(1031) <= layer0_outputs(288);
    outputs(1032) <= (layer0_outputs(1596)) and (layer0_outputs(2188));
    outputs(1033) <= (layer0_outputs(852)) xor (layer0_outputs(221));
    outputs(1034) <= not(layer0_outputs(2412)) or (layer0_outputs(513));
    outputs(1035) <= layer0_outputs(56);
    outputs(1036) <= layer0_outputs(1333);
    outputs(1037) <= layer0_outputs(1630);
    outputs(1038) <= layer0_outputs(986);
    outputs(1039) <= not(layer0_outputs(811));
    outputs(1040) <= layer0_outputs(1689);
    outputs(1041) <= (layer0_outputs(704)) or (layer0_outputs(1484));
    outputs(1042) <= (layer0_outputs(2373)) and not (layer0_outputs(108));
    outputs(1043) <= not(layer0_outputs(1582));
    outputs(1044) <= layer0_outputs(366);
    outputs(1045) <= (layer0_outputs(307)) and (layer0_outputs(2468));
    outputs(1046) <= (layer0_outputs(2052)) and (layer0_outputs(750));
    outputs(1047) <= layer0_outputs(1359);
    outputs(1048) <= not(layer0_outputs(2501));
    outputs(1049) <= (layer0_outputs(1857)) or (layer0_outputs(1074));
    outputs(1050) <= layer0_outputs(2077);
    outputs(1051) <= (layer0_outputs(1020)) and not (layer0_outputs(988));
    outputs(1052) <= (layer0_outputs(125)) and not (layer0_outputs(1716));
    outputs(1053) <= (layer0_outputs(683)) and (layer0_outputs(2306));
    outputs(1054) <= (layer0_outputs(2111)) xor (layer0_outputs(2120));
    outputs(1055) <= not(layer0_outputs(1660));
    outputs(1056) <= layer0_outputs(366);
    outputs(1057) <= layer0_outputs(2519);
    outputs(1058) <= not(layer0_outputs(164));
    outputs(1059) <= not(layer0_outputs(1905));
    outputs(1060) <= not(layer0_outputs(821));
    outputs(1061) <= not(layer0_outputs(2525));
    outputs(1062) <= (layer0_outputs(1629)) and not (layer0_outputs(641));
    outputs(1063) <= layer0_outputs(1638);
    outputs(1064) <= layer0_outputs(1275);
    outputs(1065) <= not(layer0_outputs(103));
    outputs(1066) <= not((layer0_outputs(929)) or (layer0_outputs(729)));
    outputs(1067) <= not(layer0_outputs(2434));
    outputs(1068) <= not(layer0_outputs(712));
    outputs(1069) <= (layer0_outputs(60)) and not (layer0_outputs(767));
    outputs(1070) <= not(layer0_outputs(1445));
    outputs(1071) <= not(layer0_outputs(1801));
    outputs(1072) <= not(layer0_outputs(1355));
    outputs(1073) <= layer0_outputs(790);
    outputs(1074) <= not(layer0_outputs(184));
    outputs(1075) <= layer0_outputs(587);
    outputs(1076) <= layer0_outputs(2555);
    outputs(1077) <= layer0_outputs(1770);
    outputs(1078) <= (layer0_outputs(1979)) and not (layer0_outputs(1674));
    outputs(1079) <= not((layer0_outputs(1826)) and (layer0_outputs(1159)));
    outputs(1080) <= not(layer0_outputs(1966));
    outputs(1081) <= not(layer0_outputs(259));
    outputs(1082) <= (layer0_outputs(2128)) or (layer0_outputs(1301));
    outputs(1083) <= not(layer0_outputs(653));
    outputs(1084) <= not((layer0_outputs(786)) or (layer0_outputs(1119)));
    outputs(1085) <= not(layer0_outputs(257));
    outputs(1086) <= not((layer0_outputs(1804)) and (layer0_outputs(656)));
    outputs(1087) <= layer0_outputs(1306);
    outputs(1088) <= not((layer0_outputs(1534)) or (layer0_outputs(1581)));
    outputs(1089) <= not((layer0_outputs(722)) or (layer0_outputs(1390)));
    outputs(1090) <= (layer0_outputs(2297)) and (layer0_outputs(1803));
    outputs(1091) <= layer0_outputs(424);
    outputs(1092) <= (layer0_outputs(435)) and not (layer0_outputs(154));
    outputs(1093) <= not((layer0_outputs(1671)) or (layer0_outputs(931)));
    outputs(1094) <= layer0_outputs(127);
    outputs(1095) <= layer0_outputs(1141);
    outputs(1096) <= layer0_outputs(1012);
    outputs(1097) <= not((layer0_outputs(964)) or (layer0_outputs(374)));
    outputs(1098) <= not((layer0_outputs(2250)) or (layer0_outputs(1806)));
    outputs(1099) <= not((layer0_outputs(2387)) or (layer0_outputs(2105)));
    outputs(1100) <= not((layer0_outputs(1728)) xor (layer0_outputs(554)));
    outputs(1101) <= layer0_outputs(1520);
    outputs(1102) <= layer0_outputs(951);
    outputs(1103) <= not(layer0_outputs(1106));
    outputs(1104) <= (layer0_outputs(1050)) and not (layer0_outputs(138));
    outputs(1105) <= not(layer0_outputs(721));
    outputs(1106) <= not(layer0_outputs(1184)) or (layer0_outputs(831));
    outputs(1107) <= not((layer0_outputs(2194)) or (layer0_outputs(1000)));
    outputs(1108) <= (layer0_outputs(1361)) or (layer0_outputs(2056));
    outputs(1109) <= layer0_outputs(2379);
    outputs(1110) <= (layer0_outputs(1872)) and (layer0_outputs(2368));
    outputs(1111) <= not(layer0_outputs(1047));
    outputs(1112) <= not((layer0_outputs(1246)) xor (layer0_outputs(1857)));
    outputs(1113) <= not(layer0_outputs(1985));
    outputs(1114) <= (layer0_outputs(295)) and not (layer0_outputs(1616));
    outputs(1115) <= (layer0_outputs(1550)) and (layer0_outputs(546));
    outputs(1116) <= (layer0_outputs(2423)) and not (layer0_outputs(219));
    outputs(1117) <= layer0_outputs(2060);
    outputs(1118) <= (layer0_outputs(660)) and not (layer0_outputs(2195));
    outputs(1119) <= layer0_outputs(820);
    outputs(1120) <= (layer0_outputs(1456)) and not (layer0_outputs(967));
    outputs(1121) <= (layer0_outputs(1601)) and not (layer0_outputs(1470));
    outputs(1122) <= not(layer0_outputs(550));
    outputs(1123) <= not((layer0_outputs(580)) or (layer0_outputs(2212)));
    outputs(1124) <= not(layer0_outputs(721));
    outputs(1125) <= not(layer0_outputs(334)) or (layer0_outputs(2288));
    outputs(1126) <= not((layer0_outputs(1785)) or (layer0_outputs(1462)));
    outputs(1127) <= (layer0_outputs(2385)) and not (layer0_outputs(1672));
    outputs(1128) <= not(layer0_outputs(2372));
    outputs(1129) <= not((layer0_outputs(2082)) and (layer0_outputs(959)));
    outputs(1130) <= not(layer0_outputs(2434));
    outputs(1131) <= not(layer0_outputs(1993));
    outputs(1132) <= (layer0_outputs(1508)) and not (layer0_outputs(892));
    outputs(1133) <= not(layer0_outputs(1075)) or (layer0_outputs(58));
    outputs(1134) <= (layer0_outputs(659)) and not (layer0_outputs(224));
    outputs(1135) <= not(layer0_outputs(1607));
    outputs(1136) <= (layer0_outputs(2232)) and not (layer0_outputs(2062));
    outputs(1137) <= (layer0_outputs(1236)) and (layer0_outputs(1968));
    outputs(1138) <= layer0_outputs(1935);
    outputs(1139) <= layer0_outputs(397);
    outputs(1140) <= layer0_outputs(647);
    outputs(1141) <= not(layer0_outputs(1454));
    outputs(1142) <= not(layer0_outputs(408));
    outputs(1143) <= not(layer0_outputs(2244));
    outputs(1144) <= layer0_outputs(1348);
    outputs(1145) <= not(layer0_outputs(596));
    outputs(1146) <= not((layer0_outputs(651)) or (layer0_outputs(2500)));
    outputs(1147) <= not(layer0_outputs(949)) or (layer0_outputs(1152));
    outputs(1148) <= not(layer0_outputs(2195));
    outputs(1149) <= layer0_outputs(270);
    outputs(1150) <= (layer0_outputs(945)) and not (layer0_outputs(2130));
    outputs(1151) <= (layer0_outputs(755)) and not (layer0_outputs(2114));
    outputs(1152) <= layer0_outputs(2511);
    outputs(1153) <= not(layer0_outputs(2304));
    outputs(1154) <= not((layer0_outputs(2198)) or (layer0_outputs(1472)));
    outputs(1155) <= not((layer0_outputs(2108)) or (layer0_outputs(273)));
    outputs(1156) <= not((layer0_outputs(1514)) and (layer0_outputs(829)));
    outputs(1157) <= (layer0_outputs(1273)) and not (layer0_outputs(891));
    outputs(1158) <= (layer0_outputs(82)) xor (layer0_outputs(950));
    outputs(1159) <= (layer0_outputs(1530)) and (layer0_outputs(990));
    outputs(1160) <= not((layer0_outputs(2525)) or (layer0_outputs(2073)));
    outputs(1161) <= (layer0_outputs(1043)) and (layer0_outputs(1841));
    outputs(1162) <= (layer0_outputs(468)) and not (layer0_outputs(51));
    outputs(1163) <= not(layer0_outputs(1140));
    outputs(1164) <= not(layer0_outputs(2264));
    outputs(1165) <= not(layer0_outputs(434));
    outputs(1166) <= layer0_outputs(690);
    outputs(1167) <= not(layer0_outputs(2454));
    outputs(1168) <= not(layer0_outputs(2527));
    outputs(1169) <= (layer0_outputs(2145)) or (layer0_outputs(1290));
    outputs(1170) <= (layer0_outputs(1302)) and not (layer0_outputs(800));
    outputs(1171) <= layer0_outputs(1549);
    outputs(1172) <= layer0_outputs(968);
    outputs(1173) <= not(layer0_outputs(2414));
    outputs(1174) <= layer0_outputs(17);
    outputs(1175) <= layer0_outputs(1324);
    outputs(1176) <= not((layer0_outputs(2279)) or (layer0_outputs(108)));
    outputs(1177) <= layer0_outputs(744);
    outputs(1178) <= layer0_outputs(2063);
    outputs(1179) <= (layer0_outputs(113)) and not (layer0_outputs(2401));
    outputs(1180) <= not(layer0_outputs(2250));
    outputs(1181) <= (layer0_outputs(1444)) and not (layer0_outputs(1349));
    outputs(1182) <= layer0_outputs(2036);
    outputs(1183) <= layer0_outputs(626);
    outputs(1184) <= not(layer0_outputs(2187));
    outputs(1185) <= not(layer0_outputs(251));
    outputs(1186) <= layer0_outputs(1926);
    outputs(1187) <= not(layer0_outputs(2415));
    outputs(1188) <= not(layer0_outputs(785));
    outputs(1189) <= not((layer0_outputs(704)) xor (layer0_outputs(1522)));
    outputs(1190) <= not(layer0_outputs(1761));
    outputs(1191) <= (layer0_outputs(1039)) and not (layer0_outputs(1945));
    outputs(1192) <= layer0_outputs(887);
    outputs(1193) <= not((layer0_outputs(1985)) and (layer0_outputs(2510)));
    outputs(1194) <= not(layer0_outputs(2224));
    outputs(1195) <= layer0_outputs(1557);
    outputs(1196) <= not(layer0_outputs(989));
    outputs(1197) <= (layer0_outputs(1512)) and not (layer0_outputs(2386));
    outputs(1198) <= not(layer0_outputs(196));
    outputs(1199) <= (layer0_outputs(2263)) and not (layer0_outputs(1396));
    outputs(1200) <= (layer0_outputs(189)) and (layer0_outputs(1241));
    outputs(1201) <= (layer0_outputs(2403)) or (layer0_outputs(413));
    outputs(1202) <= not(layer0_outputs(919)) or (layer0_outputs(893));
    outputs(1203) <= layer0_outputs(2037);
    outputs(1204) <= (layer0_outputs(2030)) or (layer0_outputs(2081));
    outputs(1205) <= layer0_outputs(2052);
    outputs(1206) <= not(layer0_outputs(2530));
    outputs(1207) <= layer0_outputs(516);
    outputs(1208) <= (layer0_outputs(2150)) and not (layer0_outputs(1896));
    outputs(1209) <= (layer0_outputs(964)) xor (layer0_outputs(94));
    outputs(1210) <= (layer0_outputs(275)) and (layer0_outputs(1138));
    outputs(1211) <= layer0_outputs(1587);
    outputs(1212) <= (layer0_outputs(860)) and not (layer0_outputs(115));
    outputs(1213) <= layer0_outputs(222);
    outputs(1214) <= (layer0_outputs(917)) and not (layer0_outputs(2350));
    outputs(1215) <= (layer0_outputs(373)) xor (layer0_outputs(1544));
    outputs(1216) <= layer0_outputs(1749);
    outputs(1217) <= layer0_outputs(39);
    outputs(1218) <= layer0_outputs(227);
    outputs(1219) <= layer0_outputs(1669);
    outputs(1220) <= layer0_outputs(1755);
    outputs(1221) <= not((layer0_outputs(1347)) or (layer0_outputs(49)));
    outputs(1222) <= not(layer0_outputs(301));
    outputs(1223) <= not((layer0_outputs(2217)) or (layer0_outputs(2383)));
    outputs(1224) <= not((layer0_outputs(1957)) or (layer0_outputs(117)));
    outputs(1225) <= (layer0_outputs(1626)) or (layer0_outputs(826));
    outputs(1226) <= not(layer0_outputs(1272));
    outputs(1227) <= not(layer0_outputs(2093));
    outputs(1228) <= (layer0_outputs(2439)) and not (layer0_outputs(368));
    outputs(1229) <= not((layer0_outputs(1913)) or (layer0_outputs(2053)));
    outputs(1230) <= not(layer0_outputs(711));
    outputs(1231) <= (layer0_outputs(1863)) and not (layer0_outputs(1194));
    outputs(1232) <= not(layer0_outputs(1879));
    outputs(1233) <= (layer0_outputs(1224)) and not (layer0_outputs(872));
    outputs(1234) <= (layer0_outputs(98)) and not (layer0_outputs(1056));
    outputs(1235) <= (layer0_outputs(1018)) and (layer0_outputs(213));
    outputs(1236) <= (layer0_outputs(1770)) and not (layer0_outputs(1260));
    outputs(1237) <= (layer0_outputs(143)) and (layer0_outputs(23));
    outputs(1238) <= layer0_outputs(799);
    outputs(1239) <= layer0_outputs(1167);
    outputs(1240) <= not(layer0_outputs(973));
    outputs(1241) <= not(layer0_outputs(1607));
    outputs(1242) <= layer0_outputs(151);
    outputs(1243) <= not((layer0_outputs(684)) xor (layer0_outputs(866)));
    outputs(1244) <= (layer0_outputs(1286)) and not (layer0_outputs(276));
    outputs(1245) <= layer0_outputs(847);
    outputs(1246) <= (layer0_outputs(1791)) and not (layer0_outputs(1321));
    outputs(1247) <= layer0_outputs(2190);
    outputs(1248) <= (layer0_outputs(2035)) and not (layer0_outputs(2261));
    outputs(1249) <= (layer0_outputs(1909)) or (layer0_outputs(1974));
    outputs(1250) <= layer0_outputs(655);
    outputs(1251) <= layer0_outputs(2446);
    outputs(1252) <= (layer0_outputs(2208)) or (layer0_outputs(1298));
    outputs(1253) <= layer0_outputs(635);
    outputs(1254) <= not(layer0_outputs(2270));
    outputs(1255) <= layer0_outputs(369);
    outputs(1256) <= not(layer0_outputs(2271));
    outputs(1257) <= not(layer0_outputs(2026)) or (layer0_outputs(1620));
    outputs(1258) <= layer0_outputs(1042);
    outputs(1259) <= not((layer0_outputs(489)) or (layer0_outputs(305)));
    outputs(1260) <= not((layer0_outputs(336)) or (layer0_outputs(490)));
    outputs(1261) <= layer0_outputs(362);
    outputs(1262) <= (layer0_outputs(1752)) and (layer0_outputs(1380));
    outputs(1263) <= layer0_outputs(1975);
    outputs(1264) <= (layer0_outputs(1735)) and not (layer0_outputs(1700));
    outputs(1265) <= (layer0_outputs(1990)) and (layer0_outputs(1541));
    outputs(1266) <= layer0_outputs(2003);
    outputs(1267) <= layer0_outputs(1936);
    outputs(1268) <= not((layer0_outputs(1147)) and (layer0_outputs(1473)));
    outputs(1269) <= layer0_outputs(126);
    outputs(1270) <= (layer0_outputs(2326)) and (layer0_outputs(1370));
    outputs(1271) <= (layer0_outputs(24)) xor (layer0_outputs(517));
    outputs(1272) <= not(layer0_outputs(2027));
    outputs(1273) <= (layer0_outputs(120)) and not (layer0_outputs(1316));
    outputs(1274) <= (layer0_outputs(441)) and not (layer0_outputs(2237));
    outputs(1275) <= not(layer0_outputs(2033));
    outputs(1276) <= (layer0_outputs(1323)) and not (layer0_outputs(873));
    outputs(1277) <= not(layer0_outputs(1981));
    outputs(1278) <= (layer0_outputs(2277)) and not (layer0_outputs(2317));
    outputs(1279) <= layer0_outputs(359);
    outputs(1280) <= layer0_outputs(760);
    outputs(1281) <= layer0_outputs(2403);
    outputs(1282) <= layer0_outputs(2410);
    outputs(1283) <= (layer0_outputs(214)) and not (layer0_outputs(915));
    outputs(1284) <= (layer0_outputs(2257)) and not (layer0_outputs(1130));
    outputs(1285) <= not(layer0_outputs(497));
    outputs(1286) <= not(layer0_outputs(1335));
    outputs(1287) <= not(layer0_outputs(1298));
    outputs(1288) <= not((layer0_outputs(1765)) xor (layer0_outputs(282)));
    outputs(1289) <= not(layer0_outputs(1873));
    outputs(1290) <= (layer0_outputs(487)) or (layer0_outputs(1455));
    outputs(1291) <= not(layer0_outputs(334)) or (layer0_outputs(1778));
    outputs(1292) <= not(layer0_outputs(1235));
    outputs(1293) <= not(layer0_outputs(2399));
    outputs(1294) <= not((layer0_outputs(1661)) or (layer0_outputs(1014)));
    outputs(1295) <= not(layer0_outputs(1192));
    outputs(1296) <= (layer0_outputs(281)) and not (layer0_outputs(899));
    outputs(1297) <= (layer0_outputs(1021)) and not (layer0_outputs(835));
    outputs(1298) <= not((layer0_outputs(1218)) or (layer0_outputs(6)));
    outputs(1299) <= not(layer0_outputs(1699));
    outputs(1300) <= not((layer0_outputs(1917)) and (layer0_outputs(1407)));
    outputs(1301) <= layer0_outputs(1793);
    outputs(1302) <= layer0_outputs(2168);
    outputs(1303) <= (layer0_outputs(1717)) xor (layer0_outputs(2046));
    outputs(1304) <= not((layer0_outputs(2447)) xor (layer0_outputs(2258)));
    outputs(1305) <= layer0_outputs(1276);
    outputs(1306) <= not(layer0_outputs(102));
    outputs(1307) <= not((layer0_outputs(209)) xor (layer0_outputs(2467)));
    outputs(1308) <= (layer0_outputs(629)) and not (layer0_outputs(1052));
    outputs(1309) <= (layer0_outputs(2000)) and (layer0_outputs(1713));
    outputs(1310) <= (layer0_outputs(1113)) and (layer0_outputs(1865));
    outputs(1311) <= (layer0_outputs(1890)) and (layer0_outputs(1847));
    outputs(1312) <= layer0_outputs(2127);
    outputs(1313) <= not((layer0_outputs(1815)) xor (layer0_outputs(345)));
    outputs(1314) <= layer0_outputs(1856);
    outputs(1315) <= layer0_outputs(2343);
    outputs(1316) <= not(layer0_outputs(10)) or (layer0_outputs(1767));
    outputs(1317) <= (layer0_outputs(505)) and not (layer0_outputs(174));
    outputs(1318) <= layer0_outputs(413);
    outputs(1319) <= layer0_outputs(1246);
    outputs(1320) <= (layer0_outputs(327)) and (layer0_outputs(1227));
    outputs(1321) <= not(layer0_outputs(1724)) or (layer0_outputs(1017));
    outputs(1322) <= not(layer0_outputs(1604));
    outputs(1323) <= (layer0_outputs(128)) and (layer0_outputs(981));
    outputs(1324) <= (layer0_outputs(1160)) xor (layer0_outputs(2471));
    outputs(1325) <= (layer0_outputs(1882)) and not (layer0_outputs(136));
    outputs(1326) <= not((layer0_outputs(1783)) or (layer0_outputs(2017)));
    outputs(1327) <= layer0_outputs(2161);
    outputs(1328) <= not(layer0_outputs(1045));
    outputs(1329) <= not((layer0_outputs(2484)) or (layer0_outputs(1157)));
    outputs(1330) <= not(layer0_outputs(1263));
    outputs(1331) <= layer0_outputs(107);
    outputs(1332) <= not((layer0_outputs(2444)) xor (layer0_outputs(1622)));
    outputs(1333) <= not((layer0_outputs(942)) or (layer0_outputs(1998)));
    outputs(1334) <= (layer0_outputs(268)) xor (layer0_outputs(1526));
    outputs(1335) <= not(layer0_outputs(980));
    outputs(1336) <= not(layer0_outputs(859));
    outputs(1337) <= layer0_outputs(898);
    outputs(1338) <= layer0_outputs(1952);
    outputs(1339) <= (layer0_outputs(1612)) and (layer0_outputs(2117));
    outputs(1340) <= not(layer0_outputs(91)) or (layer0_outputs(2240));
    outputs(1341) <= (layer0_outputs(371)) and (layer0_outputs(18));
    outputs(1342) <= not(layer0_outputs(1771));
    outputs(1343) <= not(layer0_outputs(2160)) or (layer0_outputs(1595));
    outputs(1344) <= layer0_outputs(1840);
    outputs(1345) <= (layer0_outputs(861)) and not (layer0_outputs(545));
    outputs(1346) <= layer0_outputs(1026);
    outputs(1347) <= (layer0_outputs(429)) and not (layer0_outputs(1855));
    outputs(1348) <= not(layer0_outputs(349));
    outputs(1349) <= not(layer0_outputs(190));
    outputs(1350) <= layer0_outputs(544);
    outputs(1351) <= layer0_outputs(1183);
    outputs(1352) <= not((layer0_outputs(995)) and (layer0_outputs(2369)));
    outputs(1353) <= (layer0_outputs(461)) and (layer0_outputs(1521));
    outputs(1354) <= not((layer0_outputs(2505)) xor (layer0_outputs(216)));
    outputs(1355) <= layer0_outputs(2196);
    outputs(1356) <= (layer0_outputs(2205)) and not (layer0_outputs(914));
    outputs(1357) <= (layer0_outputs(999)) and not (layer0_outputs(1824));
    outputs(1358) <= not((layer0_outputs(638)) and (layer0_outputs(1758)));
    outputs(1359) <= (layer0_outputs(2463)) and not (layer0_outputs(2335));
    outputs(1360) <= not((layer0_outputs(2008)) xor (layer0_outputs(720)));
    outputs(1361) <= (layer0_outputs(2175)) and not (layer0_outputs(360));
    outputs(1362) <= layer0_outputs(2123);
    outputs(1363) <= not((layer0_outputs(1125)) or (layer0_outputs(426)));
    outputs(1364) <= (layer0_outputs(101)) or (layer0_outputs(1203));
    outputs(1365) <= not(layer0_outputs(556)) or (layer0_outputs(2129));
    outputs(1366) <= layer0_outputs(1294);
    outputs(1367) <= layer0_outputs(733);
    outputs(1368) <= not((layer0_outputs(2069)) xor (layer0_outputs(629)));
    outputs(1369) <= (layer0_outputs(666)) and not (layer0_outputs(1729));
    outputs(1370) <= not(layer0_outputs(44));
    outputs(1371) <= (layer0_outputs(267)) and not (layer0_outputs(2551));
    outputs(1372) <= layer0_outputs(1474);
    outputs(1373) <= not((layer0_outputs(1803)) xor (layer0_outputs(1333)));
    outputs(1374) <= not((layer0_outputs(1478)) or (layer0_outputs(353)));
    outputs(1375) <= layer0_outputs(1142);
    outputs(1376) <= not(layer0_outputs(1990));
    outputs(1377) <= (layer0_outputs(1769)) and (layer0_outputs(1019));
    outputs(1378) <= (layer0_outputs(1403)) xor (layer0_outputs(1465));
    outputs(1379) <= not(layer0_outputs(1709));
    outputs(1380) <= not(layer0_outputs(2367));
    outputs(1381) <= (layer0_outputs(72)) and not (layer0_outputs(1861));
    outputs(1382) <= not((layer0_outputs(1698)) xor (layer0_outputs(2126)));
    outputs(1383) <= (layer0_outputs(1931)) and not (layer0_outputs(1361));
    outputs(1384) <= not(layer0_outputs(2492)) or (layer0_outputs(590));
    outputs(1385) <= not(layer0_outputs(529));
    outputs(1386) <= layer0_outputs(2154);
    outputs(1387) <= (layer0_outputs(1326)) and not (layer0_outputs(1592));
    outputs(1388) <= not(layer0_outputs(207));
    outputs(1389) <= (layer0_outputs(1625)) xor (layer0_outputs(1737));
    outputs(1390) <= not(layer0_outputs(1859));
    outputs(1391) <= not(layer0_outputs(858));
    outputs(1392) <= not(layer0_outputs(582));
    outputs(1393) <= not(layer0_outputs(19)) or (layer0_outputs(2358));
    outputs(1394) <= layer0_outputs(2481);
    outputs(1395) <= (layer0_outputs(1196)) or (layer0_outputs(2252));
    outputs(1396) <= (layer0_outputs(266)) and not (layer0_outputs(651));
    outputs(1397) <= not((layer0_outputs(710)) and (layer0_outputs(2019)));
    outputs(1398) <= not(layer0_outputs(1147));
    outputs(1399) <= not(layer0_outputs(511));
    outputs(1400) <= layer0_outputs(80);
    outputs(1401) <= (layer0_outputs(1844)) xor (layer0_outputs(1716));
    outputs(1402) <= not((layer0_outputs(2314)) xor (layer0_outputs(178)));
    outputs(1403) <= not(layer0_outputs(454)) or (layer0_outputs(1838));
    outputs(1404) <= not(layer0_outputs(249));
    outputs(1405) <= (layer0_outputs(1026)) and not (layer0_outputs(225));
    outputs(1406) <= (layer0_outputs(168)) xor (layer0_outputs(1280));
    outputs(1407) <= not(layer0_outputs(516)) or (layer0_outputs(1315));
    outputs(1408) <= not(layer0_outputs(2194));
    outputs(1409) <= not(layer0_outputs(2499));
    outputs(1410) <= layer0_outputs(1060);
    outputs(1411) <= (layer0_outputs(1054)) and not (layer0_outputs(1625));
    outputs(1412) <= layer0_outputs(1547);
    outputs(1413) <= not(layer0_outputs(604));
    outputs(1414) <= (layer0_outputs(646)) and not (layer0_outputs(356));
    outputs(1415) <= not(layer0_outputs(2111)) or (layer0_outputs(1479));
    outputs(1416) <= (layer0_outputs(982)) and (layer0_outputs(2455));
    outputs(1417) <= not((layer0_outputs(1441)) or (layer0_outputs(2072)));
    outputs(1418) <= layer0_outputs(355);
    outputs(1419) <= (layer0_outputs(95)) and not (layer0_outputs(1226));
    outputs(1420) <= (layer0_outputs(1564)) or (layer0_outputs(442));
    outputs(1421) <= not(layer0_outputs(648));
    outputs(1422) <= not(layer0_outputs(2035));
    outputs(1423) <= (layer0_outputs(1307)) and not (layer0_outputs(299));
    outputs(1424) <= (layer0_outputs(1789)) and (layer0_outputs(1374));
    outputs(1425) <= not(layer0_outputs(1677));
    outputs(1426) <= layer0_outputs(608);
    outputs(1427) <= layer0_outputs(1598);
    outputs(1428) <= (layer0_outputs(291)) and (layer0_outputs(1232));
    outputs(1429) <= layer0_outputs(1979);
    outputs(1430) <= not((layer0_outputs(8)) or (layer0_outputs(2408)));
    outputs(1431) <= layer0_outputs(1775);
    outputs(1432) <= (layer0_outputs(1029)) and (layer0_outputs(1486));
    outputs(1433) <= layer0_outputs(2493);
    outputs(1434) <= (layer0_outputs(1370)) and not (layer0_outputs(88));
    outputs(1435) <= layer0_outputs(72);
    outputs(1436) <= layer0_outputs(1071);
    outputs(1437) <= (layer0_outputs(2251)) or (layer0_outputs(1364));
    outputs(1438) <= layer0_outputs(477);
    outputs(1439) <= layer0_outputs(481);
    outputs(1440) <= not((layer0_outputs(640)) and (layer0_outputs(2171)));
    outputs(1441) <= (layer0_outputs(1368)) or (layer0_outputs(2101));
    outputs(1442) <= (layer0_outputs(2266)) and not (layer0_outputs(1064));
    outputs(1443) <= not(layer0_outputs(2480));
    outputs(1444) <= not((layer0_outputs(1133)) and (layer0_outputs(941)));
    outputs(1445) <= layer0_outputs(2229);
    outputs(1446) <= layer0_outputs(344);
    outputs(1447) <= layer0_outputs(1564);
    outputs(1448) <= not((layer0_outputs(441)) or (layer0_outputs(894)));
    outputs(1449) <= (layer0_outputs(320)) xor (layer0_outputs(47));
    outputs(1450) <= layer0_outputs(1631);
    outputs(1451) <= (layer0_outputs(1009)) and not (layer0_outputs(1989));
    outputs(1452) <= (layer0_outputs(527)) xor (layer0_outputs(326));
    outputs(1453) <= (layer0_outputs(907)) and not (layer0_outputs(1603));
    outputs(1454) <= not(layer0_outputs(1184)) or (layer0_outputs(1107));
    outputs(1455) <= not(layer0_outputs(1994));
    outputs(1456) <= not(layer0_outputs(847));
    outputs(1457) <= not((layer0_outputs(1647)) or (layer0_outputs(986)));
    outputs(1458) <= not((layer0_outputs(2255)) or (layer0_outputs(2313)));
    outputs(1459) <= not(layer0_outputs(1686));
    outputs(1460) <= not(layer0_outputs(2160));
    outputs(1461) <= (layer0_outputs(214)) and not (layer0_outputs(1732));
    outputs(1462) <= layer0_outputs(1006);
    outputs(1463) <= (layer0_outputs(1314)) xor (layer0_outputs(654));
    outputs(1464) <= not(layer0_outputs(1251)) or (layer0_outputs(2496));
    outputs(1465) <= layer0_outputs(1156);
    outputs(1466) <= layer0_outputs(1864);
    outputs(1467) <= (layer0_outputs(1371)) and not (layer0_outputs(1414));
    outputs(1468) <= not(layer0_outputs(1000));
    outputs(1469) <= layer0_outputs(691);
    outputs(1470) <= not((layer0_outputs(1488)) and (layer0_outputs(1580)));
    outputs(1471) <= not(layer0_outputs(379));
    outputs(1472) <= not((layer0_outputs(2260)) xor (layer0_outputs(1800)));
    outputs(1473) <= (layer0_outputs(1727)) and (layer0_outputs(450));
    outputs(1474) <= not((layer0_outputs(61)) or (layer0_outputs(1643)));
    outputs(1475) <= layer0_outputs(265);
    outputs(1476) <= layer0_outputs(1588);
    outputs(1477) <= not(layer0_outputs(1783));
    outputs(1478) <= not(layer0_outputs(1950));
    outputs(1479) <= not(layer0_outputs(10)) or (layer0_outputs(1347));
    outputs(1480) <= not(layer0_outputs(1057));
    outputs(1481) <= not(layer0_outputs(615));
    outputs(1482) <= not((layer0_outputs(1956)) or (layer0_outputs(508)));
    outputs(1483) <= (layer0_outputs(656)) and not (layer0_outputs(2094));
    outputs(1484) <= not(layer0_outputs(783));
    outputs(1485) <= layer0_outputs(2165);
    outputs(1486) <= (layer0_outputs(832)) xor (layer0_outputs(563));
    outputs(1487) <= layer0_outputs(2457);
    outputs(1488) <= layer0_outputs(2289);
    outputs(1489) <= (layer0_outputs(1900)) and not (layer0_outputs(1376));
    outputs(1490) <= not((layer0_outputs(2152)) or (layer0_outputs(1395)));
    outputs(1491) <= not(layer0_outputs(2043));
    outputs(1492) <= (layer0_outputs(727)) and not (layer0_outputs(621));
    outputs(1493) <= not(layer0_outputs(1491));
    outputs(1494) <= (layer0_outputs(1063)) and not (layer0_outputs(1354));
    outputs(1495) <= not(layer0_outputs(2081));
    outputs(1496) <= (layer0_outputs(1896)) or (layer0_outputs(2245));
    outputs(1497) <= (layer0_outputs(254)) or (layer0_outputs(1568));
    outputs(1498) <= layer0_outputs(1590);
    outputs(1499) <= not(layer0_outputs(1842));
    outputs(1500) <= (layer0_outputs(2546)) and not (layer0_outputs(1948));
    outputs(1501) <= not(layer0_outputs(2340));
    outputs(1502) <= (layer0_outputs(1340)) and not (layer0_outputs(848));
    outputs(1503) <= (layer0_outputs(1691)) and not (layer0_outputs(675));
    outputs(1504) <= not(layer0_outputs(706)) or (layer0_outputs(194));
    outputs(1505) <= (layer0_outputs(626)) and not (layer0_outputs(1185));
    outputs(1506) <= not(layer0_outputs(2232));
    outputs(1507) <= (layer0_outputs(1969)) and (layer0_outputs(1127));
    outputs(1508) <= layer0_outputs(1706);
    outputs(1509) <= not((layer0_outputs(724)) or (layer0_outputs(1190)));
    outputs(1510) <= (layer0_outputs(2371)) and (layer0_outputs(215));
    outputs(1511) <= (layer0_outputs(633)) xor (layer0_outputs(713));
    outputs(1512) <= (layer0_outputs(2427)) and not (layer0_outputs(1581));
    outputs(1513) <= (layer0_outputs(443)) and (layer0_outputs(1519));
    outputs(1514) <= not((layer0_outputs(2235)) and (layer0_outputs(2062)));
    outputs(1515) <= layer0_outputs(878);
    outputs(1516) <= layer0_outputs(1748);
    outputs(1517) <= not((layer0_outputs(1627)) xor (layer0_outputs(2013)));
    outputs(1518) <= not(layer0_outputs(1199));
    outputs(1519) <= not((layer0_outputs(1482)) xor (layer0_outputs(86)));
    outputs(1520) <= (layer0_outputs(2479)) and (layer0_outputs(2371));
    outputs(1521) <= not((layer0_outputs(333)) or (layer0_outputs(937)));
    outputs(1522) <= (layer0_outputs(80)) and (layer0_outputs(890));
    outputs(1523) <= not(layer0_outputs(1154));
    outputs(1524) <= not(layer0_outputs(2223));
    outputs(1525) <= not(layer0_outputs(1089));
    outputs(1526) <= (layer0_outputs(2055)) xor (layer0_outputs(1366));
    outputs(1527) <= not(layer0_outputs(531)) or (layer0_outputs(117));
    outputs(1528) <= not((layer0_outputs(1746)) or (layer0_outputs(1744)));
    outputs(1529) <= not((layer0_outputs(2264)) and (layer0_outputs(2459)));
    outputs(1530) <= not((layer0_outputs(2182)) xor (layer0_outputs(2280)));
    outputs(1531) <= (layer0_outputs(2374)) and not (layer0_outputs(1038));
    outputs(1532) <= layer0_outputs(2557);
    outputs(1533) <= (layer0_outputs(537)) and (layer0_outputs(2427));
    outputs(1534) <= (layer0_outputs(501)) and not (layer0_outputs(612));
    outputs(1535) <= layer0_outputs(1955);
    outputs(1536) <= (layer0_outputs(2530)) or (layer0_outputs(614));
    outputs(1537) <= not(layer0_outputs(991));
    outputs(1538) <= layer0_outputs(1046);
    outputs(1539) <= not(layer0_outputs(419));
    outputs(1540) <= (layer0_outputs(204)) and not (layer0_outputs(2380));
    outputs(1541) <= (layer0_outputs(20)) and not (layer0_outputs(1311));
    outputs(1542) <= not(layer0_outputs(1165));
    outputs(1543) <= layer0_outputs(1249);
    outputs(1544) <= (layer0_outputs(1868)) and not (layer0_outputs(1169));
    outputs(1545) <= layer0_outputs(2296);
    outputs(1546) <= not((layer0_outputs(84)) or (layer0_outputs(28)));
    outputs(1547) <= (layer0_outputs(537)) and (layer0_outputs(1965));
    outputs(1548) <= not((layer0_outputs(712)) or (layer0_outputs(353)));
    outputs(1549) <= (layer0_outputs(1638)) and not (layer0_outputs(2552));
    outputs(1550) <= layer0_outputs(2461);
    outputs(1551) <= (layer0_outputs(105)) and not (layer0_outputs(2539));
    outputs(1552) <= not(layer0_outputs(1074));
    outputs(1553) <= not((layer0_outputs(997)) or (layer0_outputs(315)));
    outputs(1554) <= (layer0_outputs(882)) and (layer0_outputs(1666));
    outputs(1555) <= (layer0_outputs(182)) and not (layer0_outputs(948));
    outputs(1556) <= (layer0_outputs(1976)) and not (layer0_outputs(1096));
    outputs(1557) <= not(layer0_outputs(2096)) or (layer0_outputs(475));
    outputs(1558) <= (layer0_outputs(246)) and not (layer0_outputs(777));
    outputs(1559) <= not(layer0_outputs(1791));
    outputs(1560) <= (layer0_outputs(1903)) and (layer0_outputs(563));
    outputs(1561) <= (layer0_outputs(2319)) and not (layer0_outputs(1312));
    outputs(1562) <= not(layer0_outputs(1828));
    outputs(1563) <= not(layer0_outputs(958)) or (layer0_outputs(772));
    outputs(1564) <= not((layer0_outputs(498)) or (layer0_outputs(1978)));
    outputs(1565) <= not((layer0_outputs(1012)) and (layer0_outputs(2333)));
    outputs(1566) <= not(layer0_outputs(2099));
    outputs(1567) <= layer0_outputs(2243);
    outputs(1568) <= (layer0_outputs(1593)) and (layer0_outputs(538));
    outputs(1569) <= not(layer0_outputs(577));
    outputs(1570) <= (layer0_outputs(1120)) and (layer0_outputs(1313));
    outputs(1571) <= not(layer0_outputs(618)) or (layer0_outputs(1557));
    outputs(1572) <= not((layer0_outputs(2241)) or (layer0_outputs(1098)));
    outputs(1573) <= layer0_outputs(1400);
    outputs(1574) <= not(layer0_outputs(2108));
    outputs(1575) <= layer0_outputs(1683);
    outputs(1576) <= not(layer0_outputs(1912));
    outputs(1577) <= (layer0_outputs(979)) or (layer0_outputs(1173));
    outputs(1578) <= not(layer0_outputs(176));
    outputs(1579) <= not(layer0_outputs(719)) or (layer0_outputs(2246));
    outputs(1580) <= layer0_outputs(1816);
    outputs(1581) <= not((layer0_outputs(1420)) or (layer0_outputs(2416)));
    outputs(1582) <= (layer0_outputs(197)) and not (layer0_outputs(317));
    outputs(1583) <= not(layer0_outputs(1413));
    outputs(1584) <= (layer0_outputs(1900)) and not (layer0_outputs(1489));
    outputs(1585) <= layer0_outputs(2010);
    outputs(1586) <= not(layer0_outputs(381));
    outputs(1587) <= not(layer0_outputs(874)) or (layer0_outputs(1509));
    outputs(1588) <= layer0_outputs(2021);
    outputs(1589) <= layer0_outputs(1057);
    outputs(1590) <= not((layer0_outputs(1970)) or (layer0_outputs(491)));
    outputs(1591) <= layer0_outputs(3);
    outputs(1592) <= (layer0_outputs(2414)) and not (layer0_outputs(396));
    outputs(1593) <= not(layer0_outputs(146));
    outputs(1594) <= not(layer0_outputs(1606));
    outputs(1595) <= not(layer0_outputs(237));
    outputs(1596) <= layer0_outputs(1536);
    outputs(1597) <= layer0_outputs(1965);
    outputs(1598) <= layer0_outputs(2554);
    outputs(1599) <= not(layer0_outputs(2531));
    outputs(1600) <= (layer0_outputs(2462)) and not (layer0_outputs(1001));
    outputs(1601) <= (layer0_outputs(2134)) and not (layer0_outputs(957));
    outputs(1602) <= (layer0_outputs(415)) and (layer0_outputs(1375));
    outputs(1603) <= not((layer0_outputs(97)) xor (layer0_outputs(1523)));
    outputs(1604) <= (layer0_outputs(199)) or (layer0_outputs(2519));
    outputs(1605) <= not(layer0_outputs(1614));
    outputs(1606) <= (layer0_outputs(559)) xor (layer0_outputs(1139));
    outputs(1607) <= layer0_outputs(1391);
    outputs(1608) <= (layer0_outputs(936)) and not (layer0_outputs(978));
    outputs(1609) <= (layer0_outputs(1188)) and not (layer0_outputs(2409));
    outputs(1610) <= layer0_outputs(1486);
    outputs(1611) <= (layer0_outputs(1115)) xor (layer0_outputs(2483));
    outputs(1612) <= (layer0_outputs(778)) and not (layer0_outputs(2474));
    outputs(1613) <= (layer0_outputs(1020)) and (layer0_outputs(2462));
    outputs(1614) <= layer0_outputs(1657);
    outputs(1615) <= layer0_outputs(594);
    outputs(1616) <= not((layer0_outputs(233)) or (layer0_outputs(535)));
    outputs(1617) <= not(layer0_outputs(146));
    outputs(1618) <= layer0_outputs(1825);
    outputs(1619) <= not((layer0_outputs(2146)) xor (layer0_outputs(998)));
    outputs(1620) <= layer0_outputs(2315);
    outputs(1621) <= not((layer0_outputs(1640)) xor (layer0_outputs(162)));
    outputs(1622) <= (layer0_outputs(88)) and not (layer0_outputs(312));
    outputs(1623) <= (layer0_outputs(52)) and not (layer0_outputs(1943));
    outputs(1624) <= (layer0_outputs(2078)) xor (layer0_outputs(2460));
    outputs(1625) <= not(layer0_outputs(1357)) or (layer0_outputs(1269));
    outputs(1626) <= not(layer0_outputs(1738));
    outputs(1627) <= not(layer0_outputs(180));
    outputs(1628) <= layer0_outputs(1809);
    outputs(1629) <= (layer0_outputs(1008)) xor (layer0_outputs(1369));
    outputs(1630) <= layer0_outputs(2058);
    outputs(1631) <= (layer0_outputs(1722)) and not (layer0_outputs(773));
    outputs(1632) <= not(layer0_outputs(1521));
    outputs(1633) <= (layer0_outputs(2189)) and not (layer0_outputs(2144));
    outputs(1634) <= not(layer0_outputs(111));
    outputs(1635) <= layer0_outputs(1757);
    outputs(1636) <= (layer0_outputs(1898)) and not (layer0_outputs(2024));
    outputs(1637) <= (layer0_outputs(722)) and not (layer0_outputs(1189));
    outputs(1638) <= (layer0_outputs(1790)) and not (layer0_outputs(1633));
    outputs(1639) <= not(layer0_outputs(738));
    outputs(1640) <= not(layer0_outputs(1166));
    outputs(1641) <= not((layer0_outputs(2324)) or (layer0_outputs(2210)));
    outputs(1642) <= (layer0_outputs(2174)) and not (layer0_outputs(318));
    outputs(1643) <= (layer0_outputs(2094)) and (layer0_outputs(2128));
    outputs(1644) <= not(layer0_outputs(663)) or (layer0_outputs(1249));
    outputs(1645) <= not((layer0_outputs(2474)) or (layer0_outputs(1198)));
    outputs(1646) <= layer0_outputs(2186);
    outputs(1647) <= layer0_outputs(2089);
    outputs(1648) <= layer0_outputs(1740);
    outputs(1649) <= not(layer0_outputs(1135));
    outputs(1650) <= not((layer0_outputs(2323)) or (layer0_outputs(406)));
    outputs(1651) <= (layer0_outputs(342)) and not (layer0_outputs(394));
    outputs(1652) <= not(layer0_outputs(1076));
    outputs(1653) <= not(layer0_outputs(181));
    outputs(1654) <= (layer0_outputs(2266)) and not (layer0_outputs(2011));
    outputs(1655) <= (layer0_outputs(1613)) and (layer0_outputs(1461));
    outputs(1656) <= (layer0_outputs(150)) and not (layer0_outputs(658));
    outputs(1657) <= (layer0_outputs(425)) xor (layer0_outputs(1936));
    outputs(1658) <= layer0_outputs(1781);
    outputs(1659) <= layer0_outputs(2220);
    outputs(1660) <= not(layer0_outputs(1577)) or (layer0_outputs(1004));
    outputs(1661) <= not((layer0_outputs(1776)) or (layer0_outputs(1153)));
    outputs(1662) <= not(layer0_outputs(483));
    outputs(1663) <= not(layer0_outputs(1233));
    outputs(1664) <= not(layer0_outputs(1654)) or (layer0_outputs(2040));
    outputs(1665) <= not(layer0_outputs(1387)) or (layer0_outputs(203));
    outputs(1666) <= not(layer0_outputs(1013)) or (layer0_outputs(1270));
    outputs(1667) <= layer0_outputs(1673);
    outputs(1668) <= not((layer0_outputs(392)) or (layer0_outputs(1296)));
    outputs(1669) <= (layer0_outputs(2218)) and not (layer0_outputs(1759));
    outputs(1670) <= layer0_outputs(1560);
    outputs(1671) <= layer0_outputs(1659);
    outputs(1672) <= layer0_outputs(1769);
    outputs(1673) <= not(layer0_outputs(219));
    outputs(1674) <= layer0_outputs(2316);
    outputs(1675) <= layer0_outputs(357);
    outputs(1676) <= not(layer0_outputs(1811));
    outputs(1677) <= (layer0_outputs(1924)) and (layer0_outputs(926));
    outputs(1678) <= layer0_outputs(391);
    outputs(1679) <= not(layer0_outputs(1089));
    outputs(1680) <= not(layer0_outputs(718)) or (layer0_outputs(90));
    outputs(1681) <= not(layer0_outputs(237));
    outputs(1682) <= layer0_outputs(977);
    outputs(1683) <= (layer0_outputs(469)) and not (layer0_outputs(1104));
    outputs(1684) <= not((layer0_outputs(1087)) xor (layer0_outputs(1054)));
    outputs(1685) <= not(layer0_outputs(11));
    outputs(1686) <= not(layer0_outputs(1577));
    outputs(1687) <= not(layer0_outputs(168));
    outputs(1688) <= layer0_outputs(1110);
    outputs(1689) <= not(layer0_outputs(1286)) or (layer0_outputs(513));
    outputs(1690) <= (layer0_outputs(1301)) and not (layer0_outputs(1096));
    outputs(1691) <= not(layer0_outputs(1007));
    outputs(1692) <= (layer0_outputs(354)) and not (layer0_outputs(2170));
    outputs(1693) <= (layer0_outputs(1786)) and not (layer0_outputs(1201));
    outputs(1694) <= not(layer0_outputs(1178));
    outputs(1695) <= layer0_outputs(145);
    outputs(1696) <= not((layer0_outputs(2443)) xor (layer0_outputs(1274)));
    outputs(1697) <= not(layer0_outputs(2071)) or (layer0_outputs(1525));
    outputs(1698) <= not((layer0_outputs(1713)) xor (layer0_outputs(1025)));
    outputs(1699) <= (layer0_outputs(779)) and (layer0_outputs(1));
    outputs(1700) <= not((layer0_outputs(780)) or (layer0_outputs(960)));
    outputs(1701) <= not(layer0_outputs(2320)) or (layer0_outputs(2143));
    outputs(1702) <= (layer0_outputs(131)) and not (layer0_outputs(2558));
    outputs(1703) <= not((layer0_outputs(1420)) or (layer0_outputs(939)));
    outputs(1704) <= not((layer0_outputs(1128)) xor (layer0_outputs(1602)));
    outputs(1705) <= not((layer0_outputs(223)) and (layer0_outputs(392)));
    outputs(1706) <= not((layer0_outputs(1418)) xor (layer0_outputs(2408)));
    outputs(1707) <= (layer0_outputs(902)) and not (layer0_outputs(1894));
    outputs(1708) <= layer0_outputs(1458);
    outputs(1709) <= not((layer0_outputs(991)) or (layer0_outputs(1059)));
    outputs(1710) <= layer0_outputs(1349);
    outputs(1711) <= layer0_outputs(2087);
    outputs(1712) <= (layer0_outputs(1959)) and not (layer0_outputs(2281));
    outputs(1713) <= not(layer0_outputs(1289));
    outputs(1714) <= layer0_outputs(1798);
    outputs(1715) <= not(layer0_outputs(1440));
    outputs(1716) <= (layer0_outputs(1866)) and (layer0_outputs(514));
    outputs(1717) <= (layer0_outputs(2057)) and not (layer0_outputs(1919));
    outputs(1718) <= layer0_outputs(2146);
    outputs(1719) <= layer0_outputs(395);
    outputs(1720) <= (layer0_outputs(1543)) and (layer0_outputs(1901));
    outputs(1721) <= not(layer0_outputs(1751));
    outputs(1722) <= not(layer0_outputs(1712));
    outputs(1723) <= not(layer0_outputs(1518)) or (layer0_outputs(1714));
    outputs(1724) <= layer0_outputs(1056);
    outputs(1725) <= layer0_outputs(462);
    outputs(1726) <= not(layer0_outputs(944));
    outputs(1727) <= (layer0_outputs(2354)) and (layer0_outputs(182));
    outputs(1728) <= (layer0_outputs(1818)) and not (layer0_outputs(174));
    outputs(1729) <= layer0_outputs(246);
    outputs(1730) <= not(layer0_outputs(137)) or (layer0_outputs(75));
    outputs(1731) <= (layer0_outputs(2038)) and not (layer0_outputs(1385));
    outputs(1732) <= (layer0_outputs(1148)) and (layer0_outputs(1798));
    outputs(1733) <= (layer0_outputs(383)) and not (layer0_outputs(2416));
    outputs(1734) <= layer0_outputs(795);
    outputs(1735) <= not(layer0_outputs(2103));
    outputs(1736) <= not(layer0_outputs(2121));
    outputs(1737) <= not((layer0_outputs(661)) or (layer0_outputs(1439)));
    outputs(1738) <= not(layer0_outputs(2508));
    outputs(1739) <= (layer0_outputs(1316)) and not (layer0_outputs(2242));
    outputs(1740) <= not(layer0_outputs(1013));
    outputs(1741) <= not(layer0_outputs(446));
    outputs(1742) <= layer0_outputs(2384);
    outputs(1743) <= not(layer0_outputs(2092));
    outputs(1744) <= not((layer0_outputs(109)) and (layer0_outputs(749)));
    outputs(1745) <= (layer0_outputs(468)) and (layer0_outputs(2053));
    outputs(1746) <= not(layer0_outputs(1189));
    outputs(1747) <= layer0_outputs(1734);
    outputs(1748) <= not((layer0_outputs(2029)) or (layer0_outputs(1741)));
    outputs(1749) <= layer0_outputs(1158);
    outputs(1750) <= layer0_outputs(444);
    outputs(1751) <= (layer0_outputs(811)) and not (layer0_outputs(895));
    outputs(1752) <= not(layer0_outputs(740)) or (layer0_outputs(650));
    outputs(1753) <= not(layer0_outputs(545));
    outputs(1754) <= (layer0_outputs(1047)) and not (layer0_outputs(2482));
    outputs(1755) <= (layer0_outputs(1336)) or (layer0_outputs(974));
    outputs(1756) <= not(layer0_outputs(2256));
    outputs(1757) <= not((layer0_outputs(2185)) or (layer0_outputs(135)));
    outputs(1758) <= layer0_outputs(383);
    outputs(1759) <= not(layer0_outputs(429)) or (layer0_outputs(1084));
    outputs(1760) <= (layer0_outputs(1617)) and not (layer0_outputs(857));
    outputs(1761) <= layer0_outputs(1179);
    outputs(1762) <= (layer0_outputs(365)) and (layer0_outputs(1543));
    outputs(1763) <= (layer0_outputs(198)) and not (layer0_outputs(1098));
    outputs(1764) <= layer0_outputs(887);
    outputs(1765) <= not(layer0_outputs(121));
    outputs(1766) <= layer0_outputs(463);
    outputs(1767) <= (layer0_outputs(2074)) and not (layer0_outputs(944));
    outputs(1768) <= (layer0_outputs(1570)) and (layer0_outputs(1005));
    outputs(1769) <= not(layer0_outputs(752));
    outputs(1770) <= (layer0_outputs(1257)) and (layer0_outputs(961));
    outputs(1771) <= (layer0_outputs(1449)) and not (layer0_outputs(567));
    outputs(1772) <= not(layer0_outputs(2473));
    outputs(1773) <= not(layer0_outputs(1999));
    outputs(1774) <= (layer0_outputs(302)) xor (layer0_outputs(37));
    outputs(1775) <= (layer0_outputs(1946)) and not (layer0_outputs(519));
    outputs(1776) <= not((layer0_outputs(1533)) xor (layer0_outputs(68)));
    outputs(1777) <= (layer0_outputs(208)) and not (layer0_outputs(2311));
    outputs(1778) <= (layer0_outputs(144)) and not (layer0_outputs(2207));
    outputs(1779) <= not(layer0_outputs(381));
    outputs(1780) <= layer0_outputs(2039);
    outputs(1781) <= layer0_outputs(1553);
    outputs(1782) <= (layer0_outputs(346)) and not (layer0_outputs(1180));
    outputs(1783) <= layer0_outputs(1928);
    outputs(1784) <= not(layer0_outputs(1676)) or (layer0_outputs(340));
    outputs(1785) <= (layer0_outputs(1695)) and (layer0_outputs(110));
    outputs(1786) <= not(layer0_outputs(1811));
    outputs(1787) <= layer0_outputs(2175);
    outputs(1788) <= not(layer0_outputs(2433));
    outputs(1789) <= not((layer0_outputs(1482)) or (layer0_outputs(2486)));
    outputs(1790) <= (layer0_outputs(2177)) and (layer0_outputs(841));
    outputs(1791) <= not(layer0_outputs(2538));
    outputs(1792) <= (layer0_outputs(1255)) and not (layer0_outputs(786));
    outputs(1793) <= (layer0_outputs(1594)) and (layer0_outputs(1926));
    outputs(1794) <= not(layer0_outputs(1090)) or (layer0_outputs(100));
    outputs(1795) <= not(layer0_outputs(1820));
    outputs(1796) <= not((layer0_outputs(1432)) or (layer0_outputs(510)));
    outputs(1797) <= (layer0_outputs(1932)) and not (layer0_outputs(1322));
    outputs(1798) <= not(layer0_outputs(1493));
    outputs(1799) <= not(layer0_outputs(207));
    outputs(1800) <= not(layer0_outputs(1560));
    outputs(1801) <= not(layer0_outputs(671));
    outputs(1802) <= layer0_outputs(1912);
    outputs(1803) <= not(layer0_outputs(2222));
    outputs(1804) <= (layer0_outputs(1195)) and not (layer0_outputs(464));
    outputs(1805) <= (layer0_outputs(940)) and not (layer0_outputs(2364));
    outputs(1806) <= not((layer0_outputs(463)) or (layer0_outputs(1797)));
    outputs(1807) <= (layer0_outputs(487)) and not (layer0_outputs(1083));
    outputs(1808) <= not(layer0_outputs(888));
    outputs(1809) <= (layer0_outputs(1677)) or (layer0_outputs(1442));
    outputs(1810) <= not(layer0_outputs(271));
    outputs(1811) <= not(layer0_outputs(1458));
    outputs(1812) <= not(layer0_outputs(562));
    outputs(1813) <= (layer0_outputs(1747)) and not (layer0_outputs(1149));
    outputs(1814) <= not(layer0_outputs(693));
    outputs(1815) <= not(layer0_outputs(48));
    outputs(1816) <= not(layer0_outputs(1346)) or (layer0_outputs(78));
    outputs(1817) <= not((layer0_outputs(1462)) or (layer0_outputs(1035)));
    outputs(1818) <= (layer0_outputs(1325)) and (layer0_outputs(1078));
    outputs(1819) <= not(layer0_outputs(1466));
    outputs(1820) <= layer0_outputs(2082);
    outputs(1821) <= not((layer0_outputs(1229)) or (layer0_outputs(2331)));
    outputs(1822) <= not((layer0_outputs(2155)) or (layer0_outputs(636)));
    outputs(1823) <= not((layer0_outputs(1766)) or (layer0_outputs(2267)));
    outputs(1824) <= not((layer0_outputs(1655)) xor (layer0_outputs(2262)));
    outputs(1825) <= (layer0_outputs(1880)) and (layer0_outputs(77));
    outputs(1826) <= layer0_outputs(906);
    outputs(1827) <= (layer0_outputs(1160)) and not (layer0_outputs(982));
    outputs(1828) <= layer0_outputs(307);
    outputs(1829) <= layer0_outputs(2002);
    outputs(1830) <= not((layer0_outputs(2163)) xor (layer0_outputs(240)));
    outputs(1831) <= (layer0_outputs(1637)) and (layer0_outputs(1345));
    outputs(1832) <= (layer0_outputs(1539)) and not (layer0_outputs(430));
    outputs(1833) <= (layer0_outputs(66)) and not (layer0_outputs(2104));
    outputs(1834) <= (layer0_outputs(407)) and not (layer0_outputs(2187));
    outputs(1835) <= (layer0_outputs(2300)) and (layer0_outputs(681));
    outputs(1836) <= (layer0_outputs(1836)) and (layer0_outputs(875));
    outputs(1837) <= not(layer0_outputs(507));
    outputs(1838) <= not((layer0_outputs(1031)) or (layer0_outputs(1101)));
    outputs(1839) <= layer0_outputs(2083);
    outputs(1840) <= not(layer0_outputs(560));
    outputs(1841) <= (layer0_outputs(1404)) and (layer0_outputs(66));
    outputs(1842) <= (layer0_outputs(2473)) and not (layer0_outputs(2475));
    outputs(1843) <= (layer0_outputs(1967)) and not (layer0_outputs(2268));
    outputs(1844) <= layer0_outputs(2549);
    outputs(1845) <= layer0_outputs(2066);
    outputs(1846) <= not((layer0_outputs(968)) xor (layer0_outputs(1728)));
    outputs(1847) <= layer0_outputs(1650);
    outputs(1848) <= not((layer0_outputs(1642)) or (layer0_outputs(1854)));
    outputs(1849) <= not((layer0_outputs(1022)) or (layer0_outputs(540)));
    outputs(1850) <= not((layer0_outputs(395)) or (layer0_outputs(2475)));
    outputs(1851) <= (layer0_outputs(277)) or (layer0_outputs(205));
    outputs(1852) <= not((layer0_outputs(1313)) and (layer0_outputs(1332)));
    outputs(1853) <= not(layer0_outputs(14)) or (layer0_outputs(532));
    outputs(1854) <= not(layer0_outputs(1424));
    outputs(1855) <= (layer0_outputs(534)) and not (layer0_outputs(2483));
    outputs(1856) <= (layer0_outputs(206)) and not (layer0_outputs(195));
    outputs(1857) <= (layer0_outputs(787)) xor (layer0_outputs(220));
    outputs(1858) <= (layer0_outputs(38)) and (layer0_outputs(911));
    outputs(1859) <= (layer0_outputs(2464)) and not (layer0_outputs(1917));
    outputs(1860) <= (layer0_outputs(910)) and not (layer0_outputs(518));
    outputs(1861) <= (layer0_outputs(1892)) and (layer0_outputs(2047));
    outputs(1862) <= layer0_outputs(856);
    outputs(1863) <= not(layer0_outputs(2359));
    outputs(1864) <= layer0_outputs(1001);
    outputs(1865) <= (layer0_outputs(778)) and not (layer0_outputs(1448));
    outputs(1866) <= not(layer0_outputs(157));
    outputs(1867) <= layer0_outputs(414);
    outputs(1868) <= not((layer0_outputs(864)) and (layer0_outputs(2315)));
    outputs(1869) <= (layer0_outputs(765)) xor (layer0_outputs(1489));
    outputs(1870) <= layer0_outputs(1214);
    outputs(1871) <= (layer0_outputs(1183)) and not (layer0_outputs(2294));
    outputs(1872) <= not((layer0_outputs(82)) xor (layer0_outputs(2362)));
    outputs(1873) <= not((layer0_outputs(801)) xor (layer0_outputs(1827)));
    outputs(1874) <= (layer0_outputs(2242)) xor (layer0_outputs(179));
    outputs(1875) <= (layer0_outputs(1834)) or (layer0_outputs(2407));
    outputs(1876) <= not((layer0_outputs(457)) or (layer0_outputs(1785)));
    outputs(1877) <= layer0_outputs(376);
    outputs(1878) <= not((layer0_outputs(1561)) or (layer0_outputs(321)));
    outputs(1879) <= (layer0_outputs(2235)) xor (layer0_outputs(609));
    outputs(1880) <= (layer0_outputs(263)) and (layer0_outputs(119));
    outputs(1881) <= (layer0_outputs(1675)) and not (layer0_outputs(575));
    outputs(1882) <= (layer0_outputs(485)) or (layer0_outputs(1474));
    outputs(1883) <= (layer0_outputs(1268)) and not (layer0_outputs(1792));
    outputs(1884) <= layer0_outputs(2311);
    outputs(1885) <= layer0_outputs(2251);
    outputs(1886) <= layer0_outputs(1701);
    outputs(1887) <= (layer0_outputs(988)) and (layer0_outputs(1352));
    outputs(1888) <= (layer0_outputs(1682)) and not (layer0_outputs(2517));
    outputs(1889) <= not((layer0_outputs(2158)) or (layer0_outputs(2325)));
    outputs(1890) <= not(layer0_outputs(1217)) or (layer0_outputs(1911));
    outputs(1891) <= (layer0_outputs(525)) and (layer0_outputs(1923));
    outputs(1892) <= (layer0_outputs(1763)) and (layer0_outputs(194));
    outputs(1893) <= (layer0_outputs(291)) and not (layer0_outputs(809));
    outputs(1894) <= not(layer0_outputs(1988));
    outputs(1895) <= (layer0_outputs(2559)) and not (layer0_outputs(673));
    outputs(1896) <= (layer0_outputs(1202)) and (layer0_outputs(258));
    outputs(1897) <= (layer0_outputs(2355)) and not (layer0_outputs(1953));
    outputs(1898) <= (layer0_outputs(1848)) and not (layer0_outputs(1326));
    outputs(1899) <= layer0_outputs(1551);
    outputs(1900) <= not((layer0_outputs(1447)) or (layer0_outputs(510)));
    outputs(1901) <= layer0_outputs(1011);
    outputs(1902) <= (layer0_outputs(961)) and not (layer0_outputs(1132));
    outputs(1903) <= not(layer0_outputs(715));
    outputs(1904) <= (layer0_outputs(1954)) and not (layer0_outputs(1615));
    outputs(1905) <= not(layer0_outputs(1726));
    outputs(1906) <= not(layer0_outputs(551));
    outputs(1907) <= not(layer0_outputs(905));
    outputs(1908) <= (layer0_outputs(2348)) or (layer0_outputs(239));
    outputs(1909) <= not((layer0_outputs(2331)) or (layer0_outputs(299)));
    outputs(1910) <= (layer0_outputs(1738)) and not (layer0_outputs(1647));
    outputs(1911) <= (layer0_outputs(2265)) and not (layer0_outputs(688));
    outputs(1912) <= not((layer0_outputs(2553)) or (layer0_outputs(553)));
    outputs(1913) <= not((layer0_outputs(1434)) or (layer0_outputs(34)));
    outputs(1914) <= layer0_outputs(2370);
    outputs(1915) <= (layer0_outputs(1591)) and (layer0_outputs(1623));
    outputs(1916) <= (layer0_outputs(1033)) and (layer0_outputs(15));
    outputs(1917) <= layer0_outputs(702);
    outputs(1918) <= (layer0_outputs(913)) and not (layer0_outputs(1593));
    outputs(1919) <= not(layer0_outputs(951));
    outputs(1920) <= layer0_outputs(1144);
    outputs(1921) <= (layer0_outputs(232)) and (layer0_outputs(592));
    outputs(1922) <= (layer0_outputs(2159)) and not (layer0_outputs(694));
    outputs(1923) <= not((layer0_outputs(1534)) or (layer0_outputs(2359)));
    outputs(1924) <= not(layer0_outputs(965));
    outputs(1925) <= not((layer0_outputs(2354)) and (layer0_outputs(2406)));
    outputs(1926) <= (layer0_outputs(1093)) and not (layer0_outputs(321));
    outputs(1927) <= (layer0_outputs(1087)) and (layer0_outputs(2178));
    outputs(1928) <= not(layer0_outputs(1721));
    outputs(1929) <= not((layer0_outputs(1710)) or (layer0_outputs(2488)));
    outputs(1930) <= (layer0_outputs(973)) and not (layer0_outputs(1816));
    outputs(1931) <= not((layer0_outputs(63)) or (layer0_outputs(803)));
    outputs(1932) <= not(layer0_outputs(554));
    outputs(1933) <= not(layer0_outputs(1250)) or (layer0_outputs(1599));
    outputs(1934) <= (layer0_outputs(903)) and not (layer0_outputs(1485));
    outputs(1935) <= not((layer0_outputs(387)) and (layer0_outputs(18)));
    outputs(1936) <= (layer0_outputs(139)) xor (layer0_outputs(1476));
    outputs(1937) <= layer0_outputs(1992);
    outputs(1938) <= not(layer0_outputs(208));
    outputs(1939) <= layer0_outputs(1635);
    outputs(1940) <= layer0_outputs(1862);
    outputs(1941) <= not((layer0_outputs(357)) and (layer0_outputs(1928)));
    outputs(1942) <= (layer0_outputs(1363)) and not (layer0_outputs(74));
    outputs(1943) <= (layer0_outputs(1888)) and not (layer0_outputs(1389));
    outputs(1944) <= (layer0_outputs(418)) and not (layer0_outputs(331));
    outputs(1945) <= (layer0_outputs(1153)) and not (layer0_outputs(1736));
    outputs(1946) <= layer0_outputs(22);
    outputs(1947) <= not((layer0_outputs(883)) xor (layer0_outputs(1090)));
    outputs(1948) <= not((layer0_outputs(799)) or (layer0_outputs(776)));
    outputs(1949) <= not(layer0_outputs(767));
    outputs(1950) <= layer0_outputs(1968);
    outputs(1951) <= (layer0_outputs(1429)) or (layer0_outputs(2467));
    outputs(1952) <= layer0_outputs(1961);
    outputs(1953) <= layer0_outputs(2385);
    outputs(1954) <= not((layer0_outputs(1715)) xor (layer0_outputs(375)));
    outputs(1955) <= not((layer0_outputs(59)) xor (layer0_outputs(1802)));
    outputs(1956) <= not(layer0_outputs(1561));
    outputs(1957) <= (layer0_outputs(22)) and not (layer0_outputs(646));
    outputs(1958) <= not(layer0_outputs(1810));
    outputs(1959) <= not((layer0_outputs(144)) or (layer0_outputs(924)));
    outputs(1960) <= not(layer0_outputs(979)) or (layer0_outputs(1465));
    outputs(1961) <= (layer0_outputs(643)) and (layer0_outputs(1873));
    outputs(1962) <= layer0_outputs(448);
    outputs(1963) <= (layer0_outputs(796)) and not (layer0_outputs(2228));
    outputs(1964) <= not((layer0_outputs(2488)) and (layer0_outputs(1411)));
    outputs(1965) <= not(layer0_outputs(2201));
    outputs(1966) <= layer0_outputs(2093);
    outputs(1967) <= not(layer0_outputs(1004));
    outputs(1968) <= (layer0_outputs(64)) or (layer0_outputs(789));
    outputs(1969) <= (layer0_outputs(1422)) and not (layer0_outputs(2283));
    outputs(1970) <= not(layer0_outputs(1842));
    outputs(1971) <= (layer0_outputs(1253)) xor (layer0_outputs(2042));
    outputs(1972) <= (layer0_outputs(8)) and not (layer0_outputs(347));
    outputs(1973) <= (layer0_outputs(1382)) xor (layer0_outputs(484));
    outputs(1974) <= (layer0_outputs(1608)) and not (layer0_outputs(27));
    outputs(1975) <= (layer0_outputs(269)) and (layer0_outputs(449));
    outputs(1976) <= (layer0_outputs(1887)) and (layer0_outputs(1268));
    outputs(1977) <= not((layer0_outputs(1540)) or (layer0_outputs(947)));
    outputs(1978) <= layer0_outputs(1624);
    outputs(1979) <= (layer0_outputs(471)) and not (layer0_outputs(14));
    outputs(1980) <= layer0_outputs(2410);
    outputs(1981) <= (layer0_outputs(1665)) and not (layer0_outputs(74));
    outputs(1982) <= not((layer0_outputs(2225)) or (layer0_outputs(2090)));
    outputs(1983) <= (layer0_outputs(119)) and (layer0_outputs(2248));
    outputs(1984) <= not(layer0_outputs(898));
    outputs(1985) <= (layer0_outputs(290)) and not (layer0_outputs(918));
    outputs(1986) <= not((layer0_outputs(2196)) or (layer0_outputs(1048)));
    outputs(1987) <= not(layer0_outputs(401));
    outputs(1988) <= (layer0_outputs(913)) and not (layer0_outputs(524));
    outputs(1989) <= layer0_outputs(2552);
    outputs(1990) <= (layer0_outputs(231)) and not (layer0_outputs(261));
    outputs(1991) <= layer0_outputs(1529);
    outputs(1992) <= (layer0_outputs(2059)) and not (layer0_outputs(2520));
    outputs(1993) <= not(layer0_outputs(340));
    outputs(1994) <= layer0_outputs(257);
    outputs(1995) <= layer0_outputs(118);
    outputs(1996) <= not((layer0_outputs(409)) or (layer0_outputs(1085)));
    outputs(1997) <= layer0_outputs(1762);
    outputs(1998) <= (layer0_outputs(2254)) and not (layer0_outputs(1947));
    outputs(1999) <= not(layer0_outputs(500));
    outputs(2000) <= not((layer0_outputs(1156)) and (layer0_outputs(389)));
    outputs(2001) <= not(layer0_outputs(462));
    outputs(2002) <= not((layer0_outputs(2070)) and (layer0_outputs(1297)));
    outputs(2003) <= not((layer0_outputs(248)) and (layer0_outputs(1579)));
    outputs(2004) <= (layer0_outputs(5)) and (layer0_outputs(2451));
    outputs(2005) <= layer0_outputs(1583);
    outputs(2006) <= (layer0_outputs(2540)) and (layer0_outputs(2066));
    outputs(2007) <= not(layer0_outputs(481));
    outputs(2008) <= not(layer0_outputs(1095));
    outputs(2009) <= (layer0_outputs(338)) and (layer0_outputs(67));
    outputs(2010) <= not(layer0_outputs(367));
    outputs(2011) <= (layer0_outputs(1093)) and (layer0_outputs(1576));
    outputs(2012) <= not(layer0_outputs(1170)) or (layer0_outputs(1621));
    outputs(2013) <= (layer0_outputs(1651)) and not (layer0_outputs(703));
    outputs(2014) <= (layer0_outputs(1305)) and (layer0_outputs(1937));
    outputs(2015) <= (layer0_outputs(620)) and not (layer0_outputs(2215));
    outputs(2016) <= not(layer0_outputs(1884));
    outputs(2017) <= (layer0_outputs(234)) and (layer0_outputs(185));
    outputs(2018) <= not(layer0_outputs(1290)) or (layer0_outputs(1597));
    outputs(2019) <= (layer0_outputs(1787)) and not (layer0_outputs(2372));
    outputs(2020) <= not(layer0_outputs(2147));
    outputs(2021) <= (layer0_outputs(1431)) or (layer0_outputs(581));
    outputs(2022) <= not((layer0_outputs(2461)) or (layer0_outputs(1653)));
    outputs(2023) <= not((layer0_outputs(1646)) or (layer0_outputs(1499)));
    outputs(2024) <= (layer0_outputs(1323)) and (layer0_outputs(837));
    outputs(2025) <= (layer0_outputs(630)) and (layer0_outputs(114));
    outputs(2026) <= (layer0_outputs(1745)) xor (layer0_outputs(807));
    outputs(2027) <= (layer0_outputs(124)) and not (layer0_outputs(36));
    outputs(2028) <= layer0_outputs(2512);
    outputs(2029) <= (layer0_outputs(1552)) and not (layer0_outputs(1408));
    outputs(2030) <= (layer0_outputs(1602)) and (layer0_outputs(1554));
    outputs(2031) <= not(layer0_outputs(1743));
    outputs(2032) <= (layer0_outputs(21)) and not (layer0_outputs(2405));
    outputs(2033) <= (layer0_outputs(1552)) and (layer0_outputs(1003));
    outputs(2034) <= layer0_outputs(1555);
    outputs(2035) <= not(layer0_outputs(706));
    outputs(2036) <= not(layer0_outputs(477));
    outputs(2037) <= (layer0_outputs(1264)) and (layer0_outputs(935));
    outputs(2038) <= layer0_outputs(2197);
    outputs(2039) <= not(layer0_outputs(2375));
    outputs(2040) <= (layer0_outputs(1730)) and not (layer0_outputs(549));
    outputs(2041) <= (layer0_outputs(314)) and not (layer0_outputs(1015));
    outputs(2042) <= layer0_outputs(1191);
    outputs(2043) <= layer0_outputs(1287);
    outputs(2044) <= not(layer0_outputs(1368));
    outputs(2045) <= not((layer0_outputs(2543)) and (layer0_outputs(1495)));
    outputs(2046) <= not(layer0_outputs(1079));
    outputs(2047) <= layer0_outputs(1986);
    outputs(2048) <= (layer0_outputs(2238)) and not (layer0_outputs(351));
    outputs(2049) <= (layer0_outputs(1707)) and not (layer0_outputs(788));
    outputs(2050) <= not((layer0_outputs(93)) or (layer0_outputs(2153)));
    outputs(2051) <= (layer0_outputs(966)) and not (layer0_outputs(322));
    outputs(2052) <= not(layer0_outputs(1951));
    outputs(2053) <= not(layer0_outputs(2009)) or (layer0_outputs(682));
    outputs(2054) <= layer0_outputs(806);
    outputs(2055) <= (layer0_outputs(241)) xor (layer0_outputs(1831));
    outputs(2056) <= (layer0_outputs(628)) and not (layer0_outputs(639));
    outputs(2057) <= layer0_outputs(900);
    outputs(2058) <= not(layer0_outputs(561));
    outputs(2059) <= not(layer0_outputs(183)) or (layer0_outputs(1654));
    outputs(2060) <= (layer0_outputs(2297)) xor (layer0_outputs(335));
    outputs(2061) <= layer0_outputs(1284);
    outputs(2062) <= not((layer0_outputs(929)) or (layer0_outputs(2267)));
    outputs(2063) <= not(layer0_outputs(1062));
    outputs(2064) <= layer0_outputs(1376);
    outputs(2065) <= not(layer0_outputs(1238));
    outputs(2066) <= not(layer0_outputs(679));
    outputs(2067) <= not(layer0_outputs(54));
    outputs(2068) <= (layer0_outputs(1847)) and not (layer0_outputs(1023));
    outputs(2069) <= layer0_outputs(2095);
    outputs(2070) <= layer0_outputs(1275);
    outputs(2071) <= layer0_outputs(962);
    outputs(2072) <= (layer0_outputs(1704)) and (layer0_outputs(1616));
    outputs(2073) <= layer0_outputs(1840);
    outputs(2074) <= (layer0_outputs(1332)) and not (layer0_outputs(688));
    outputs(2075) <= (layer0_outputs(765)) and not (layer0_outputs(1051));
    outputs(2076) <= not(layer0_outputs(1809));
    outputs(2077) <= layer0_outputs(1853);
    outputs(2078) <= layer0_outputs(809);
    outputs(2079) <= (layer0_outputs(2534)) and not (layer0_outputs(1288));
    outputs(2080) <= layer0_outputs(2404);
    outputs(2081) <= not(layer0_outputs(1327));
    outputs(2082) <= (layer0_outputs(1559)) and not (layer0_outputs(2091));
    outputs(2083) <= not(layer0_outputs(2050));
    outputs(2084) <= not((layer0_outputs(2493)) and (layer0_outputs(1902)));
    outputs(2085) <= not(layer0_outputs(372));
    outputs(2086) <= not(layer0_outputs(1586)) or (layer0_outputs(2405));
    outputs(2087) <= (layer0_outputs(1296)) and (layer0_outputs(1075));
    outputs(2088) <= layer0_outputs(1403);
    outputs(2089) <= not(layer0_outputs(2031));
    outputs(2090) <= layer0_outputs(1428);
    outputs(2091) <= (layer0_outputs(692)) and not (layer0_outputs(1699));
    outputs(2092) <= layer0_outputs(69);
    outputs(2093) <= not((layer0_outputs(2363)) xor (layer0_outputs(2339)));
    outputs(2094) <= layer0_outputs(2197);
    outputs(2095) <= (layer0_outputs(1206)) and (layer0_outputs(1429));
    outputs(2096) <= (layer0_outputs(1591)) and (layer0_outputs(2141));
    outputs(2097) <= (layer0_outputs(1103)) xor (layer0_outputs(1881));
    outputs(2098) <= layer0_outputs(2138);
    outputs(2099) <= (layer0_outputs(859)) xor (layer0_outputs(337));
    outputs(2100) <= (layer0_outputs(949)) xor (layer0_outputs(1706));
    outputs(2101) <= (layer0_outputs(154)) and (layer0_outputs(2418));
    outputs(2102) <= layer0_outputs(2424);
    outputs(2103) <= (layer0_outputs(1005)) xor (layer0_outputs(25));
    outputs(2104) <= (layer0_outputs(1545)) and not (layer0_outputs(1575));
    outputs(2105) <= not((layer0_outputs(2295)) xor (layer0_outputs(760)));
    outputs(2106) <= layer0_outputs(2191);
    outputs(2107) <= (layer0_outputs(1538)) and (layer0_outputs(1584));
    outputs(2108) <= layer0_outputs(79);
    outputs(2109) <= not(layer0_outputs(1611));
    outputs(2110) <= not(layer0_outputs(632));
    outputs(2111) <= not(layer0_outputs(669));
    outputs(2112) <= layer0_outputs(482);
    outputs(2113) <= layer0_outputs(1399);
    outputs(2114) <= not(layer0_outputs(358)) or (layer0_outputs(1459));
    outputs(2115) <= not(layer0_outputs(1406));
    outputs(2116) <= not((layer0_outputs(2409)) or (layer0_outputs(1498)));
    outputs(2117) <= not((layer0_outputs(1942)) xor (layer0_outputs(71)));
    outputs(2118) <= not(layer0_outputs(288));
    outputs(2119) <= (layer0_outputs(352)) and not (layer0_outputs(565));
    outputs(2120) <= (layer0_outputs(1411)) and not (layer0_outputs(407));
    outputs(2121) <= (layer0_outputs(284)) or (layer0_outputs(1776));
    outputs(2122) <= not(layer0_outputs(403));
    outputs(2123) <= not(layer0_outputs(792));
    outputs(2124) <= layer0_outputs(1456);
    outputs(2125) <= (layer0_outputs(123)) and (layer0_outputs(1077));
    outputs(2126) <= not(layer0_outputs(303));
    outputs(2127) <= (layer0_outputs(2178)) and (layer0_outputs(101));
    outputs(2128) <= layer0_outputs(394);
    outputs(2129) <= layer0_outputs(2113);
    outputs(2130) <= not(layer0_outputs(410));
    outputs(2131) <= (layer0_outputs(865)) and (layer0_outputs(2415));
    outputs(2132) <= not(layer0_outputs(1118));
    outputs(2133) <= not(layer0_outputs(648));
    outputs(2134) <= not(layer0_outputs(2370));
    outputs(2135) <= not(layer0_outputs(129));
    outputs(2136) <= not(layer0_outputs(183)) or (layer0_outputs(1211));
    outputs(2137) <= layer0_outputs(2192);
    outputs(2138) <= (layer0_outputs(1421)) and not (layer0_outputs(440));
    outputs(2139) <= not((layer0_outputs(687)) and (layer0_outputs(1662)));
    outputs(2140) <= not(layer0_outputs(1845)) or (layer0_outputs(2413));
    outputs(2141) <= not(layer0_outputs(2388)) or (layer0_outputs(885));
    outputs(2142) <= layer0_outputs(218);
    outputs(2143) <= layer0_outputs(1150);
    outputs(2144) <= layer0_outputs(1446);
    outputs(2145) <= layer0_outputs(2529);
    outputs(2146) <= not(layer0_outputs(110)) or (layer0_outputs(1867));
    outputs(2147) <= (layer0_outputs(2173)) and not (layer0_outputs(300));
    outputs(2148) <= (layer0_outputs(1441)) or (layer0_outputs(195));
    outputs(2149) <= not((layer0_outputs(1562)) xor (layer0_outputs(1964)));
    outputs(2150) <= not((layer0_outputs(1824)) xor (layer0_outputs(742)));
    outputs(2151) <= layer0_outputs(519);
    outputs(2152) <= (layer0_outputs(2526)) and not (layer0_outputs(104));
    outputs(2153) <= layer0_outputs(188);
    outputs(2154) <= not(layer0_outputs(12));
    outputs(2155) <= not((layer0_outputs(1680)) or (layer0_outputs(2379)));
    outputs(2156) <= layer0_outputs(1243);
    outputs(2157) <= not((layer0_outputs(1916)) or (layer0_outputs(2356)));
    outputs(2158) <= (layer0_outputs(738)) xor (layer0_outputs(1019));
    outputs(2159) <= not(layer0_outputs(105));
    outputs(2160) <= not((layer0_outputs(742)) or (layer0_outputs(2018)));
    outputs(2161) <= not(layer0_outputs(1696)) or (layer0_outputs(1295));
    outputs(2162) <= not((layer0_outputs(886)) or (layer0_outputs(708)));
    outputs(2163) <= not(layer0_outputs(2007));
    outputs(2164) <= not((layer0_outputs(702)) or (layer0_outputs(1619)));
    outputs(2165) <= (layer0_outputs(1480)) or (layer0_outputs(2176));
    outputs(2166) <= (layer0_outputs(2334)) xor (layer0_outputs(1310));
    outputs(2167) <= not(layer0_outputs(1350));
    outputs(2168) <= (layer0_outputs(1109)) and (layer0_outputs(310));
    outputs(2169) <= not(layer0_outputs(1023));
    outputs(2170) <= (layer0_outputs(774)) and (layer0_outputs(2025));
    outputs(2171) <= not((layer0_outputs(472)) and (layer0_outputs(1898)));
    outputs(2172) <= not(layer0_outputs(812));
    outputs(2173) <= not(layer0_outputs(729));
    outputs(2174) <= not(layer0_outputs(304));
    outputs(2175) <= not((layer0_outputs(819)) or (layer0_outputs(1492)));
    outputs(2176) <= layer0_outputs(1930);
    outputs(2177) <= not(layer0_outputs(1777));
    outputs(2178) <= layer0_outputs(1634);
    outputs(2179) <= not(layer0_outputs(756));
    outputs(2180) <= layer0_outputs(296);
    outputs(2181) <= not(layer0_outputs(2004));
    outputs(2182) <= not(layer0_outputs(1781));
    outputs(2183) <= not(layer0_outputs(50));
    outputs(2184) <= not((layer0_outputs(2191)) xor (layer0_outputs(2076)));
    outputs(2185) <= (layer0_outputs(1068)) and not (layer0_outputs(1921));
    outputs(2186) <= not((layer0_outputs(1343)) or (layer0_outputs(1423)));
    outputs(2187) <= (layer0_outputs(853)) and not (layer0_outputs(571));
    outputs(2188) <= not(layer0_outputs(1407));
    outputs(2189) <= not(layer0_outputs(2001)) or (layer0_outputs(2476));
    outputs(2190) <= layer0_outputs(2238);
    outputs(2191) <= (layer0_outputs(1880)) and not (layer0_outputs(1002));
    outputs(2192) <= not(layer0_outputs(2206));
    outputs(2193) <= not((layer0_outputs(821)) or (layer0_outputs(427)));
    outputs(2194) <= not(layer0_outputs(696));
    outputs(2195) <= layer0_outputs(758);
    outputs(2196) <= (layer0_outputs(666)) and not (layer0_outputs(2356));
    outputs(2197) <= layer0_outputs(2184);
    outputs(2198) <= (layer0_outputs(876)) and not (layer0_outputs(129));
    outputs(2199) <= layer0_outputs(1691);
    outputs(2200) <= not((layer0_outputs(582)) and (layer0_outputs(1036)));
    outputs(2201) <= (layer0_outputs(2529)) and (layer0_outputs(2526));
    outputs(2202) <= not(layer0_outputs(302));
    outputs(2203) <= not(layer0_outputs(2032));
    outputs(2204) <= not(layer0_outputs(2442));
    outputs(2205) <= layer0_outputs(1145);
    outputs(2206) <= layer0_outputs(411);
    outputs(2207) <= layer0_outputs(431);
    outputs(2208) <= not(layer0_outputs(1177));
    outputs(2209) <= (layer0_outputs(1964)) xor (layer0_outputs(1066));
    outputs(2210) <= not(layer0_outputs(770)) or (layer0_outputs(952));
    outputs(2211) <= layer0_outputs(1101);
    outputs(2212) <= layer0_outputs(2299);
    outputs(2213) <= (layer0_outputs(719)) and not (layer0_outputs(2018));
    outputs(2214) <= layer0_outputs(1830);
    outputs(2215) <= not(layer0_outputs(654));
    outputs(2216) <= layer0_outputs(1796);
    outputs(2217) <= not((layer0_outputs(1378)) and (layer0_outputs(1700)));
    outputs(2218) <= not(layer0_outputs(152));
    outputs(2219) <= (layer0_outputs(870)) and not (layer0_outputs(2423));
    outputs(2220) <= not((layer0_outputs(1998)) or (layer0_outputs(1772)));
    outputs(2221) <= layer0_outputs(915);
    outputs(2222) <= layer0_outputs(1145);
    outputs(2223) <= not(layer0_outputs(1782));
    outputs(2224) <= layer0_outputs(293);
    outputs(2225) <= not((layer0_outputs(1954)) and (layer0_outputs(768)));
    outputs(2226) <= not(layer0_outputs(1401)) or (layer0_outputs(885));
    outputs(2227) <= not(layer0_outputs(1708));
    outputs(2228) <= not(layer0_outputs(665));
    outputs(2229) <= (layer0_outputs(1377)) and (layer0_outputs(578));
    outputs(2230) <= not((layer0_outputs(1933)) and (layer0_outputs(728)));
    outputs(2231) <= not(layer0_outputs(1032));
    outputs(2232) <= not(layer0_outputs(202));
    outputs(2233) <= not(layer0_outputs(193));
    outputs(2234) <= not(layer0_outputs(1959)) or (layer0_outputs(2123));
    outputs(2235) <= layer0_outputs(1623);
    outputs(2236) <= (layer0_outputs(1388)) and (layer0_outputs(1615));
    outputs(2237) <= not((layer0_outputs(277)) or (layer0_outputs(679)));
    outputs(2238) <= (layer0_outputs(999)) and not (layer0_outputs(1107));
    outputs(2239) <= layer0_outputs(2273);
    outputs(2240) <= layer0_outputs(1034);
    outputs(2241) <= (layer0_outputs(2107)) xor (layer0_outputs(2167));
    outputs(2242) <= (layer0_outputs(2260)) and not (layer0_outputs(892));
    outputs(2243) <= layer0_outputs(2115);
    outputs(2244) <= not(layer0_outputs(879));
    outputs(2245) <= (layer0_outputs(941)) or (layer0_outputs(2507));
    outputs(2246) <= not(layer0_outputs(2358)) or (layer0_outputs(2537));
    outputs(2247) <= not(layer0_outputs(791)) or (layer0_outputs(92));
    outputs(2248) <= layer0_outputs(827);
    outputs(2249) <= not(layer0_outputs(428)) or (layer0_outputs(2230));
    outputs(2250) <= layer0_outputs(1839);
    outputs(2251) <= not(layer0_outputs(93));
    outputs(2252) <= layer0_outputs(311);
    outputs(2253) <= not((layer0_outputs(1856)) xor (layer0_outputs(245)));
    outputs(2254) <= layer0_outputs(170);
    outputs(2255) <= not((layer0_outputs(1931)) or (layer0_outputs(1935)));
    outputs(2256) <= not((layer0_outputs(541)) xor (layer0_outputs(508)));
    outputs(2257) <= not((layer0_outputs(1293)) xor (layer0_outputs(1881)));
    outputs(2258) <= layer0_outputs(367);
    outputs(2259) <= (layer0_outputs(2135)) and not (layer0_outputs(756));
    outputs(2260) <= layer0_outputs(506);
    outputs(2261) <= not((layer0_outputs(2438)) and (layer0_outputs(1929)));
    outputs(2262) <= not((layer0_outputs(1663)) and (layer0_outputs(1070)));
    outputs(2263) <= layer0_outputs(972);
    outputs(2264) <= not(layer0_outputs(2164)) or (layer0_outputs(388));
    outputs(2265) <= layer0_outputs(816);
    outputs(2266) <= not((layer0_outputs(323)) xor (layer0_outputs(1088)));
    outputs(2267) <= layer0_outputs(1117);
    outputs(2268) <= layer0_outputs(2349);
    outputs(2269) <= layer0_outputs(1449);
    outputs(2270) <= (layer0_outputs(1322)) and (layer0_outputs(2361));
    outputs(2271) <= layer0_outputs(1996);
    outputs(2272) <= layer0_outputs(564);
    outputs(2273) <= layer0_outputs(2067);
    outputs(2274) <= layer0_outputs(1723);
    outputs(2275) <= layer0_outputs(1852);
    outputs(2276) <= (layer0_outputs(371)) and not (layer0_outputs(355));
    outputs(2277) <= not((layer0_outputs(2116)) or (layer0_outputs(2486)));
    outputs(2278) <= layer0_outputs(170);
    outputs(2279) <= (layer0_outputs(1209)) xor (layer0_outputs(2523));
    outputs(2280) <= (layer0_outputs(1053)) and not (layer0_outputs(78));
    outputs(2281) <= not(layer0_outputs(469));
    outputs(2282) <= not((layer0_outputs(1649)) xor (layer0_outputs(933)));
    outputs(2283) <= (layer0_outputs(2024)) and (layer0_outputs(1668));
    outputs(2284) <= (layer0_outputs(1889)) xor (layer0_outputs(1174));
    outputs(2285) <= (layer0_outputs(795)) and not (layer0_outputs(2243));
    outputs(2286) <= (layer0_outputs(689)) xor (layer0_outputs(306));
    outputs(2287) <= (layer0_outputs(166)) and not (layer0_outputs(96));
    outputs(2288) <= layer0_outputs(55);
    outputs(2289) <= layer0_outputs(2424);
    outputs(2290) <= layer0_outputs(955);
    outputs(2291) <= not((layer0_outputs(473)) or (layer0_outputs(192)));
    outputs(2292) <= not(layer0_outputs(1317));
    outputs(2293) <= not((layer0_outputs(2327)) xor (layer0_outputs(822)));
    outputs(2294) <= (layer0_outputs(1759)) or (layer0_outputs(1922));
    outputs(2295) <= not(layer0_outputs(660));
    outputs(2296) <= not(layer0_outputs(2308));
    outputs(2297) <= (layer0_outputs(1754)) or (layer0_outputs(1658));
    outputs(2298) <= (layer0_outputs(664)) and not (layer0_outputs(229));
    outputs(2299) <= not((layer0_outputs(1311)) xor (layer0_outputs(2332)));
    outputs(2300) <= not(layer0_outputs(2440));
    outputs(2301) <= not(layer0_outputs(565));
    outputs(2302) <= not(layer0_outputs(1537));
    outputs(2303) <= (layer0_outputs(343)) and (layer0_outputs(1221));
    outputs(2304) <= not(layer0_outputs(512));
    outputs(2305) <= (layer0_outputs(939)) and (layer0_outputs(298));
    outputs(2306) <= not((layer0_outputs(2521)) and (layer0_outputs(1321)));
    outputs(2307) <= layer0_outputs(924);
    outputs(2308) <= not(layer0_outputs(1237));
    outputs(2309) <= (layer0_outputs(650)) or (layer0_outputs(43));
    outputs(2310) <= (layer0_outputs(2556)) and (layer0_outputs(454));
    outputs(2311) <= not(layer0_outputs(1386));
    outputs(2312) <= not((layer0_outputs(65)) xor (layer0_outputs(2472)));
    outputs(2313) <= (layer0_outputs(1049)) and (layer0_outputs(1556));
    outputs(2314) <= (layer0_outputs(957)) and (layer0_outputs(876));
    outputs(2315) <= layer0_outputs(780);
    outputs(2316) <= not(layer0_outputs(231));
    outputs(2317) <= layer0_outputs(1772);
    outputs(2318) <= (layer0_outputs(1436)) and not (layer0_outputs(1416));
    outputs(2319) <= layer0_outputs(2458);
    outputs(2320) <= (layer0_outputs(588)) and (layer0_outputs(1846));
    outputs(2321) <= not(layer0_outputs(380));
    outputs(2322) <= not((layer0_outputs(817)) or (layer0_outputs(1172)));
    outputs(2323) <= (layer0_outputs(227)) and not (layer0_outputs(2149));
    outputs(2324) <= (layer0_outputs(2060)) and (layer0_outputs(1007));
    outputs(2325) <= (layer0_outputs(671)) and not (layer0_outputs(566));
    outputs(2326) <= layer0_outputs(1925);
    outputs(2327) <= not(layer0_outputs(165)) or (layer0_outputs(667));
    outputs(2328) <= layer0_outputs(1171);
    outputs(2329) <= not((layer0_outputs(1216)) or (layer0_outputs(840)));
    outputs(2330) <= not(layer0_outputs(1832));
    outputs(2331) <= not((layer0_outputs(781)) or (layer0_outputs(919)));
    outputs(2332) <= (layer0_outputs(2333)) and not (layer0_outputs(1453));
    outputs(2333) <= (layer0_outputs(2302)) and not (layer0_outputs(1500));
    outputs(2334) <= not((layer0_outputs(160)) or (layer0_outputs(2469)));
    outputs(2335) <= (layer0_outputs(1024)) xor (layer0_outputs(691));
    outputs(2336) <= not((layer0_outputs(6)) and (layer0_outputs(2322)));
    outputs(2337) <= not((layer0_outputs(1915)) and (layer0_outputs(386)));
    outputs(2338) <= layer0_outputs(2367);
    outputs(2339) <= layer0_outputs(1836);
    outputs(2340) <= not(layer0_outputs(1874));
    outputs(2341) <= layer0_outputs(1941);
    outputs(2342) <= (layer0_outputs(198)) and not (layer0_outputs(1058));
    outputs(2343) <= (layer0_outputs(2369)) and not (layer0_outputs(1673));
    outputs(2344) <= (layer0_outputs(1585)) and (layer0_outputs(2497));
    outputs(2345) <= (layer0_outputs(273)) xor (layer0_outputs(845));
    outputs(2346) <= (layer0_outputs(2556)) xor (layer0_outputs(1262));
    outputs(2347) <= (layer0_outputs(1241)) and (layer0_outputs(947));
    outputs(2348) <= (layer0_outputs(416)) and not (layer0_outputs(2112));
    outputs(2349) <= (layer0_outputs(1073)) and not (layer0_outputs(1269));
    outputs(2350) <= not(layer0_outputs(2168));
    outputs(2351) <= (layer0_outputs(103)) and (layer0_outputs(2492));
    outputs(2352) <= not(layer0_outputs(2113));
    outputs(2353) <= (layer0_outputs(147)) and not (layer0_outputs(2127));
    outputs(2354) <= (layer0_outputs(121)) and (layer0_outputs(2068));
    outputs(2355) <= not(layer0_outputs(1208));
    outputs(2356) <= (layer0_outputs(1727)) and not (layer0_outputs(2198));
    outputs(2357) <= layer0_outputs(1329);
    outputs(2358) <= layer0_outputs(1306);
    outputs(2359) <= layer0_outputs(1567);
    outputs(2360) <= not(layer0_outputs(479));
    outputs(2361) <= not((layer0_outputs(20)) and (layer0_outputs(2319)));
    outputs(2362) <= not(layer0_outputs(2383));
    outputs(2363) <= not((layer0_outputs(2284)) xor (layer0_outputs(1817)));
    outputs(2364) <= not((layer0_outputs(602)) or (layer0_outputs(587)));
    outputs(2365) <= (layer0_outputs(335)) xor (layer0_outputs(1505));
    outputs(2366) <= layer0_outputs(2339);
    outputs(2367) <= (layer0_outputs(996)) and (layer0_outputs(390));
    outputs(2368) <= not(layer0_outputs(1542));
    outputs(2369) <= layer0_outputs(2088);
    outputs(2370) <= not((layer0_outputs(1245)) or (layer0_outputs(1714)));
    outputs(2371) <= not(layer0_outputs(980));
    outputs(2372) <= layer0_outputs(1222);
    outputs(2373) <= layer0_outputs(235);
    outputs(2374) <= not(layer0_outputs(1805)) or (layer0_outputs(984));
    outputs(2375) <= layer0_outputs(622);
    outputs(2376) <= (layer0_outputs(585)) and not (layer0_outputs(150));
    outputs(2377) <= (layer0_outputs(2103)) and not (layer0_outputs(228));
    outputs(2378) <= (layer0_outputs(274)) and not (layer0_outputs(1742));
    outputs(2379) <= (layer0_outputs(167)) and not (layer0_outputs(2084));
    outputs(2380) <= layer0_outputs(2115);
    outputs(2381) <= not(layer0_outputs(636));
    outputs(2382) <= (layer0_outputs(1214)) and not (layer0_outputs(549));
    outputs(2383) <= not((layer0_outputs(186)) or (layer0_outputs(2387)));
    outputs(2384) <= not((layer0_outputs(1204)) or (layer0_outputs(834)));
    outputs(2385) <= layer0_outputs(2162);
    outputs(2386) <= not(layer0_outputs(2521));
    outputs(2387) <= not(layer0_outputs(1247));
    outputs(2388) <= (layer0_outputs(1586)) and not (layer0_outputs(453));
    outputs(2389) <= layer0_outputs(1076);
    outputs(2390) <= not(layer0_outputs(763));
    outputs(2391) <= (layer0_outputs(1512)) and (layer0_outputs(2557));
    outputs(2392) <= not(layer0_outputs(680));
    outputs(2393) <= (layer0_outputs(2100)) and not (layer0_outputs(1393));
    outputs(2394) <= (layer0_outputs(2555)) and (layer0_outputs(1977));
    outputs(2395) <= layer0_outputs(2068);
    outputs(2396) <= (layer0_outputs(888)) xor (layer0_outputs(1746));
    outputs(2397) <= (layer0_outputs(2327)) and (layer0_outputs(120));
    outputs(2398) <= (layer0_outputs(1285)) and not (layer0_outputs(2224));
    outputs(2399) <= not((layer0_outputs(649)) and (layer0_outputs(2536)));
    outputs(2400) <= not(layer0_outputs(343));
    outputs(2401) <= not(layer0_outputs(377));
    outputs(2402) <= (layer0_outputs(1171)) and not (layer0_outputs(157));
    outputs(2403) <= not((layer0_outputs(329)) xor (layer0_outputs(1690)));
    outputs(2404) <= not(layer0_outputs(989));
    outputs(2405) <= (layer0_outputs(1219)) and (layer0_outputs(1176));
    outputs(2406) <= not(layer0_outputs(364));
    outputs(2407) <= layer0_outputs(337);
    outputs(2408) <= layer0_outputs(1222);
    outputs(2409) <= (layer0_outputs(557)) and (layer0_outputs(1702));
    outputs(2410) <= layer0_outputs(1961);
    outputs(2411) <= (layer0_outputs(627)) and not (layer0_outputs(1795));
    outputs(2412) <= not((layer0_outputs(802)) or (layer0_outputs(878)));
    outputs(2413) <= not(layer0_outputs(846));
    outputs(2414) <= (layer0_outputs(1133)) and (layer0_outputs(242));
    outputs(2415) <= not((layer0_outputs(1938)) or (layer0_outputs(732)));
    outputs(2416) <= not(layer0_outputs(408));
    outputs(2417) <= layer0_outputs(238);
    outputs(2418) <= not((layer0_outputs(153)) xor (layer0_outputs(1291)));
    outputs(2419) <= layer0_outputs(2226);
    outputs(2420) <= (layer0_outputs(1972)) and not (layer0_outputs(923));
    outputs(2421) <= not((layer0_outputs(1261)) or (layer0_outputs(57)));
    outputs(2422) <= layer0_outputs(1821);
    outputs(2423) <= layer0_outputs(427);
    outputs(2424) <= not((layer0_outputs(1768)) and (layer0_outputs(2344)));
    outputs(2425) <= not(layer0_outputs(1046));
    outputs(2426) <= not(layer0_outputs(798));
    outputs(2427) <= layer0_outputs(896);
    outputs(2428) <= (layer0_outputs(140)) and not (layer0_outputs(638));
    outputs(2429) <= (layer0_outputs(1722)) and not (layer0_outputs(2222));
    outputs(2430) <= layer0_outputs(1796);
    outputs(2431) <= not((layer0_outputs(2307)) or (layer0_outputs(1203)));
    outputs(2432) <= not((layer0_outputs(262)) or (layer0_outputs(2440)));
    outputs(2433) <= (layer0_outputs(1918)) xor (layer0_outputs(589));
    outputs(2434) <= not(layer0_outputs(1946));
    outputs(2435) <= layer0_outputs(220);
    outputs(2436) <= not(layer0_outputs(1849));
    outputs(2437) <= (layer0_outputs(720)) and not (layer0_outputs(828));
    outputs(2438) <= (layer0_outputs(1705)) and (layer0_outputs(375));
    outputs(2439) <= (layer0_outputs(764)) and not (layer0_outputs(2503));
    outputs(2440) <= (layer0_outputs(861)) and (layer0_outputs(2378));
    outputs(2441) <= layer0_outputs(1737);
    outputs(2442) <= (layer0_outputs(1199)) and not (layer0_outputs(1681));
    outputs(2443) <= not((layer0_outputs(998)) xor (layer0_outputs(804)));
    outputs(2444) <= (layer0_outputs(2398)) and (layer0_outputs(1865));
    outputs(2445) <= not(layer0_outputs(46));
    outputs(2446) <= (layer0_outputs(2309)) and (layer0_outputs(2174));
    outputs(2447) <= not(layer0_outputs(740));
    outputs(2448) <= (layer0_outputs(1982)) and not (layer0_outputs(759));
    outputs(2449) <= not(layer0_outputs(1445));
    outputs(2450) <= (layer0_outputs(990)) and not (layer0_outputs(566));
    outputs(2451) <= not((layer0_outputs(1694)) or (layer0_outputs(139)));
    outputs(2452) <= not(layer0_outputs(550));
    outputs(2453) <= not((layer0_outputs(2199)) or (layer0_outputs(2422)));
    outputs(2454) <= layer0_outputs(850);
    outputs(2455) <= layer0_outputs(1180);
    outputs(2456) <= not(layer0_outputs(1124));
    outputs(2457) <= (layer0_outputs(1428)) and not (layer0_outputs(256));
    outputs(2458) <= not(layer0_outputs(2237));
    outputs(2459) <= not((layer0_outputs(1491)) and (layer0_outputs(1344)));
    outputs(2460) <= not(layer0_outputs(2186));
    outputs(2461) <= (layer0_outputs(1910)) and (layer0_outputs(232));
    outputs(2462) <= (layer0_outputs(1827)) and not (layer0_outputs(1152));
    outputs(2463) <= layer0_outputs(338);
    outputs(2464) <= (layer0_outputs(2373)) and (layer0_outputs(1320));
    outputs(2465) <= not(layer0_outputs(2520));
    outputs(2466) <= layer0_outputs(2436);
    outputs(2467) <= layer0_outputs(2003);
    outputs(2468) <= not(layer0_outputs(1099));
    outputs(2469) <= not((layer0_outputs(1124)) or (layer0_outputs(1310)));
    outputs(2470) <= (layer0_outputs(2086)) and (layer0_outputs(1233));
    outputs(2471) <= (layer0_outputs(1143)) and (layer0_outputs(1037));
    outputs(2472) <= not((layer0_outputs(363)) or (layer0_outputs(2032)));
    outputs(2473) <= layer0_outputs(1531);
    outputs(2474) <= layer0_outputs(1632);
    outputs(2475) <= not(layer0_outputs(1399));
    outputs(2476) <= layer0_outputs(1365);
    outputs(2477) <= (layer0_outputs(11)) and not (layer0_outputs(818));
    outputs(2478) <= (layer0_outputs(242)) and (layer0_outputs(1807));
    outputs(2479) <= (layer0_outputs(2230)) and (layer0_outputs(1655));
    outputs(2480) <= not(layer0_outputs(1627));
    outputs(2481) <= layer0_outputs(419);
    outputs(2482) <= not(layer0_outputs(2541));
    outputs(2483) <= not(layer0_outputs(1356));
    outputs(2484) <= not(layer0_outputs(1343));
    outputs(2485) <= (layer0_outputs(634)) and (layer0_outputs(431));
    outputs(2486) <= not(layer0_outputs(410));
    outputs(2487) <= layer0_outputs(1829);
    outputs(2488) <= not(layer0_outputs(2449));
    outputs(2489) <= not((layer0_outputs(596)) or (layer0_outputs(2245)));
    outputs(2490) <= layer0_outputs(725);
    outputs(2491) <= layer0_outputs(261);
    outputs(2492) <= not(layer0_outputs(75));
    outputs(2493) <= (layer0_outputs(249)) and not (layer0_outputs(2431));
    outputs(2494) <= not(layer0_outputs(1574));
    outputs(2495) <= not(layer0_outputs(1386));
    outputs(2496) <= not(layer0_outputs(158));
    outputs(2497) <= layer0_outputs(1573);
    outputs(2498) <= not((layer0_outputs(317)) or (layer0_outputs(2204)));
    outputs(2499) <= not(layer0_outputs(398));
    outputs(2500) <= (layer0_outputs(1398)) and (layer0_outputs(1116));
    outputs(2501) <= (layer0_outputs(490)) and not (layer0_outputs(112));
    outputs(2502) <= not((layer0_outputs(1541)) or (layer0_outputs(600)));
    outputs(2503) <= not(layer0_outputs(1906));
    outputs(2504) <= layer0_outputs(238);
    outputs(2505) <= (layer0_outputs(1692)) and not (layer0_outputs(862));
    outputs(2506) <= not((layer0_outputs(753)) and (layer0_outputs(2314)));
    outputs(2507) <= (layer0_outputs(2516)) and not (layer0_outputs(2202));
    outputs(2508) <= not((layer0_outputs(967)) xor (layer0_outputs(552)));
    outputs(2509) <= (layer0_outputs(2102)) xor (layer0_outputs(1084));
    outputs(2510) <= not(layer0_outputs(1484));
    outputs(2511) <= layer0_outputs(9);
    outputs(2512) <= (layer0_outputs(535)) and not (layer0_outputs(71));
    outputs(2513) <= (layer0_outputs(292)) and (layer0_outputs(274));
    outputs(2514) <= not(layer0_outputs(352));
    outputs(2515) <= (layer0_outputs(306)) and not (layer0_outputs(2506));
    outputs(2516) <= (layer0_outputs(414)) and (layer0_outputs(1860));
    outputs(2517) <= (layer0_outputs(1902)) and not (layer0_outputs(106));
    outputs(2518) <= layer0_outputs(2355);
    outputs(2519) <= not(layer0_outputs(1148));
    outputs(2520) <= not((layer0_outputs(1525)) or (layer0_outputs(1277)));
    outputs(2521) <= layer0_outputs(156);
    outputs(2522) <= not((layer0_outputs(320)) or (layer0_outputs(272)));
    outputs(2523) <= layer0_outputs(536);
    outputs(2524) <= (layer0_outputs(359)) and not (layer0_outputs(970));
    outputs(2525) <= (layer0_outputs(558)) xor (layer0_outputs(29));
    outputs(2526) <= layer0_outputs(511);
    outputs(2527) <= (layer0_outputs(2206)) and not (layer0_outputs(1250));
    outputs(2528) <= (layer0_outputs(523)) and not (layer0_outputs(2386));
    outputs(2529) <= (layer0_outputs(1318)) and not (layer0_outputs(776));
    outputs(2530) <= layer0_outputs(2216);
    outputs(2531) <= (layer0_outputs(39)) and not (layer0_outputs(1686));
    outputs(2532) <= not((layer0_outputs(2234)) or (layer0_outputs(1103)));
    outputs(2533) <= not(layer0_outputs(2449));
    outputs(2534) <= (layer0_outputs(1648)) and not (layer0_outputs(2040));
    outputs(2535) <= not((layer0_outputs(2445)) and (layer0_outputs(458)));
    outputs(2536) <= layer0_outputs(1712);
    outputs(2537) <= layer0_outputs(1821);
    outputs(2538) <= layer0_outputs(1104);
    outputs(2539) <= not((layer0_outputs(625)) or (layer0_outputs(2303)));
    outputs(2540) <= layer0_outputs(1927);
    outputs(2541) <= not(layer0_outputs(946));
    outputs(2542) <= not((layer0_outputs(1356)) or (layer0_outputs(1527)));
    outputs(2543) <= layer0_outputs(1169);
    outputs(2544) <= not(layer0_outputs(1984)) or (layer0_outputs(1328));
    outputs(2545) <= not(layer0_outputs(1379));
    outputs(2546) <= not((layer0_outputs(1906)) or (layer0_outputs(2336)));
    outputs(2547) <= (layer0_outputs(1545)) and (layer0_outputs(2092));
    outputs(2548) <= not((layer0_outputs(992)) or (layer0_outputs(2270)));
    outputs(2549) <= layer0_outputs(2286);
    outputs(2550) <= layer0_outputs(45);
    outputs(2551) <= not(layer0_outputs(966));
    outputs(2552) <= layer0_outputs(1894);
    outputs(2553) <= not(layer0_outputs(1401));
    outputs(2554) <= not((layer0_outputs(2346)) or (layer0_outputs(2157)));
    outputs(2555) <= (layer0_outputs(1433)) and (layer0_outputs(2142));
    outputs(2556) <= (layer0_outputs(1996)) and not (layer0_outputs(675));
    outputs(2557) <= not(layer0_outputs(1721)) or (layer0_outputs(1144));
    outputs(2558) <= (layer0_outputs(1563)) and not (layer0_outputs(1272));
    outputs(2559) <= (layer0_outputs(1891)) and not (layer0_outputs(1773));

end Behavioral;
