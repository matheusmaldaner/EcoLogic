module logic_network(
    input wire [1023:0] inputs,
    output wire [9:0] outputs
);

    wire [7679:0] layer0_outputs;

    assign layer0_outputs[0] = (inputs[781]) | (inputs[612]);
    assign layer0_outputs[1] = (inputs[266]) & ~(inputs[1006]);
    assign layer0_outputs[2] = (inputs[464]) & ~(inputs[164]);
    assign layer0_outputs[3] = inputs[182];
    assign layer0_outputs[4] = (inputs[443]) & ~(inputs[827]);
    assign layer0_outputs[5] = inputs[161];
    assign layer0_outputs[6] = ~(inputs[154]);
    assign layer0_outputs[7] = (inputs[261]) | (inputs[849]);
    assign layer0_outputs[8] = (inputs[217]) & (inputs[668]);
    assign layer0_outputs[9] = ~(inputs[815]) | (inputs[757]);
    assign layer0_outputs[10] = (inputs[261]) | (inputs[24]);
    assign layer0_outputs[11] = (inputs[653]) | (inputs[188]);
    assign layer0_outputs[12] = inputs[180];
    assign layer0_outputs[13] = ~((inputs[28]) | (inputs[943]));
    assign layer0_outputs[14] = inputs[271];
    assign layer0_outputs[15] = inputs[192];
    assign layer0_outputs[16] = ~(inputs[708]) | (inputs[537]);
    assign layer0_outputs[17] = ~((inputs[244]) ^ (inputs[23]));
    assign layer0_outputs[18] = 1'b0;
    assign layer0_outputs[19] = (inputs[45]) | (inputs[357]);
    assign layer0_outputs[20] = (inputs[715]) | (inputs[181]);
    assign layer0_outputs[21] = inputs[948];
    assign layer0_outputs[22] = ~((inputs[184]) | (inputs[537]));
    assign layer0_outputs[23] = ~(inputs[633]) | (inputs[736]);
    assign layer0_outputs[24] = inputs[421];
    assign layer0_outputs[25] = (inputs[457]) | (inputs[364]);
    assign layer0_outputs[26] = inputs[694];
    assign layer0_outputs[27] = (inputs[696]) & ~(inputs[517]);
    assign layer0_outputs[28] = inputs[500];
    assign layer0_outputs[29] = inputs[368];
    assign layer0_outputs[30] = inputs[758];
    assign layer0_outputs[31] = ~((inputs[361]) | (inputs[889]));
    assign layer0_outputs[32] = ~((inputs[941]) ^ (inputs[938]));
    assign layer0_outputs[33] = (inputs[316]) & ~(inputs[740]);
    assign layer0_outputs[34] = (inputs[722]) | (inputs[518]);
    assign layer0_outputs[35] = ~((inputs[534]) ^ (inputs[175]));
    assign layer0_outputs[36] = ~((inputs[570]) | (inputs[110]));
    assign layer0_outputs[37] = (inputs[231]) ^ (inputs[352]);
    assign layer0_outputs[38] = ~(inputs[726]);
    assign layer0_outputs[39] = ~((inputs[117]) ^ (inputs[128]));
    assign layer0_outputs[40] = ~(inputs[244]);
    assign layer0_outputs[41] = ~(inputs[397]) | (inputs[843]);
    assign layer0_outputs[42] = (inputs[543]) & ~(inputs[928]);
    assign layer0_outputs[43] = ~(inputs[238]);
    assign layer0_outputs[44] = (inputs[652]) | (inputs[664]);
    assign layer0_outputs[45] = ~((inputs[53]) & (inputs[78]));
    assign layer0_outputs[46] = ~((inputs[1008]) & (inputs[32]));
    assign layer0_outputs[47] = ~((inputs[250]) | (inputs[5]));
    assign layer0_outputs[48] = 1'b0;
    assign layer0_outputs[49] = ~(inputs[308]) | (inputs[517]);
    assign layer0_outputs[50] = inputs[809];
    assign layer0_outputs[51] = 1'b0;
    assign layer0_outputs[52] = (inputs[235]) | (inputs[789]);
    assign layer0_outputs[53] = ~((inputs[740]) ^ (inputs[761]));
    assign layer0_outputs[54] = ~(inputs[654]);
    assign layer0_outputs[55] = (inputs[167]) ^ (inputs[413]);
    assign layer0_outputs[56] = (inputs[472]) | (inputs[519]);
    assign layer0_outputs[57] = 1'b1;
    assign layer0_outputs[58] = (inputs[217]) & ~(inputs[196]);
    assign layer0_outputs[59] = ~(inputs[253]);
    assign layer0_outputs[60] = ~((inputs[514]) & (inputs[295]));
    assign layer0_outputs[61] = (inputs[472]) & ~(inputs[955]);
    assign layer0_outputs[62] = ~((inputs[825]) | (inputs[684]));
    assign layer0_outputs[63] = inputs[794];
    assign layer0_outputs[64] = (inputs[909]) | (inputs[533]);
    assign layer0_outputs[65] = ~((inputs[1001]) ^ (inputs[424]));
    assign layer0_outputs[66] = (inputs[545]) | (inputs[529]);
    assign layer0_outputs[67] = (inputs[418]) & ~(inputs[291]);
    assign layer0_outputs[68] = (inputs[146]) ^ (inputs[383]);
    assign layer0_outputs[69] = (inputs[701]) ^ (inputs[266]);
    assign layer0_outputs[70] = (inputs[294]) & ~(inputs[543]);
    assign layer0_outputs[71] = inputs[310];
    assign layer0_outputs[72] = ~((inputs[211]) | (inputs[730]));
    assign layer0_outputs[73] = ~(inputs[631]);
    assign layer0_outputs[74] = (inputs[263]) & ~(inputs[412]);
    assign layer0_outputs[75] = (inputs[217]) & ~(inputs[955]);
    assign layer0_outputs[76] = ~(inputs[99]) | (inputs[982]);
    assign layer0_outputs[77] = 1'b0;
    assign layer0_outputs[78] = ~(inputs[748]) | (inputs[838]);
    assign layer0_outputs[79] = (inputs[927]) | (inputs[681]);
    assign layer0_outputs[80] = (inputs[32]) ^ (inputs[714]);
    assign layer0_outputs[81] = (inputs[818]) | (inputs[1001]);
    assign layer0_outputs[82] = (inputs[653]) & ~(inputs[294]);
    assign layer0_outputs[83] = ~(inputs[467]);
    assign layer0_outputs[84] = ~((inputs[385]) | (inputs[314]));
    assign layer0_outputs[85] = ~(inputs[601]) | (inputs[417]);
    assign layer0_outputs[86] = ~((inputs[977]) | (inputs[649]));
    assign layer0_outputs[87] = ~(inputs[789]) | (inputs[896]);
    assign layer0_outputs[88] = inputs[416];
    assign layer0_outputs[89] = ~(inputs[171]);
    assign layer0_outputs[90] = (inputs[522]) & ~(inputs[507]);
    assign layer0_outputs[91] = ~((inputs[371]) | (inputs[644]));
    assign layer0_outputs[92] = ~((inputs[536]) ^ (inputs[42]));
    assign layer0_outputs[93] = ~(inputs[810]) | (inputs[48]);
    assign layer0_outputs[94] = ~(inputs[324]);
    assign layer0_outputs[95] = ~(inputs[283]);
    assign layer0_outputs[96] = inputs[202];
    assign layer0_outputs[97] = ~(inputs[750]) | (inputs[436]);
    assign layer0_outputs[98] = ~(inputs[283]);
    assign layer0_outputs[99] = 1'b0;
    assign layer0_outputs[100] = inputs[431];
    assign layer0_outputs[101] = inputs[584];
    assign layer0_outputs[102] = (inputs[811]) & ~(inputs[669]);
    assign layer0_outputs[103] = ~(inputs[242]);
    assign layer0_outputs[104] = 1'b1;
    assign layer0_outputs[105] = (inputs[403]) & ~(inputs[439]);
    assign layer0_outputs[106] = (inputs[334]) | (inputs[948]);
    assign layer0_outputs[107] = ~((inputs[219]) | (inputs[280]));
    assign layer0_outputs[108] = ~(inputs[473]);
    assign layer0_outputs[109] = (inputs[513]) | (inputs[142]);
    assign layer0_outputs[110] = ~((inputs[326]) | (inputs[300]));
    assign layer0_outputs[111] = ~((inputs[629]) & (inputs[756]));
    assign layer0_outputs[112] = (inputs[815]) | (inputs[81]);
    assign layer0_outputs[113] = ~((inputs[168]) ^ (inputs[353]));
    assign layer0_outputs[114] = (inputs[673]) | (inputs[236]);
    assign layer0_outputs[115] = (inputs[620]) ^ (inputs[771]);
    assign layer0_outputs[116] = (inputs[187]) | (inputs[687]);
    assign layer0_outputs[117] = (inputs[476]) ^ (inputs[10]);
    assign layer0_outputs[118] = 1'b1;
    assign layer0_outputs[119] = (inputs[818]) & ~(inputs[792]);
    assign layer0_outputs[120] = (inputs[887]) & (inputs[669]);
    assign layer0_outputs[121] = (inputs[511]) & ~(inputs[46]);
    assign layer0_outputs[122] = (inputs[787]) | (inputs[50]);
    assign layer0_outputs[123] = ~(inputs[40]) | (inputs[937]);
    assign layer0_outputs[124] = (inputs[35]) | (inputs[634]);
    assign layer0_outputs[125] = ~((inputs[658]) | (inputs[520]));
    assign layer0_outputs[126] = inputs[119];
    assign layer0_outputs[127] = inputs[86];
    assign layer0_outputs[128] = (inputs[102]) ^ (inputs[945]);
    assign layer0_outputs[129] = ~((inputs[924]) ^ (inputs[392]));
    assign layer0_outputs[130] = ~((inputs[465]) | (inputs[625]));
    assign layer0_outputs[131] = ~((inputs[670]) ^ (inputs[494]));
    assign layer0_outputs[132] = ~((inputs[874]) | (inputs[727]));
    assign layer0_outputs[133] = ~(inputs[133]) | (inputs[261]);
    assign layer0_outputs[134] = ~(inputs[704]);
    assign layer0_outputs[135] = ~((inputs[426]) & (inputs[276]));
    assign layer0_outputs[136] = 1'b1;
    assign layer0_outputs[137] = (inputs[378]) | (inputs[459]);
    assign layer0_outputs[138] = ~((inputs[790]) ^ (inputs[390]));
    assign layer0_outputs[139] = 1'b0;
    assign layer0_outputs[140] = ~(inputs[496]) | (inputs[231]);
    assign layer0_outputs[141] = inputs[718];
    assign layer0_outputs[142] = (inputs[599]) & ~(inputs[838]);
    assign layer0_outputs[143] = ~(inputs[620]);
    assign layer0_outputs[144] = inputs[400];
    assign layer0_outputs[145] = ~(inputs[227]) | (inputs[608]);
    assign layer0_outputs[146] = ~((inputs[563]) | (inputs[704]));
    assign layer0_outputs[147] = (inputs[645]) | (inputs[872]);
    assign layer0_outputs[148] = (inputs[775]) & ~(inputs[977]);
    assign layer0_outputs[149] = ~(inputs[208]);
    assign layer0_outputs[150] = ~((inputs[546]) ^ (inputs[209]));
    assign layer0_outputs[151] = inputs[844];
    assign layer0_outputs[152] = ~(inputs[292]) | (inputs[393]);
    assign layer0_outputs[153] = ~(inputs[524]) | (inputs[91]);
    assign layer0_outputs[154] = (inputs[929]) ^ (inputs[332]);
    assign layer0_outputs[155] = inputs[460];
    assign layer0_outputs[156] = ~((inputs[473]) | (inputs[104]));
    assign layer0_outputs[157] = inputs[247];
    assign layer0_outputs[158] = (inputs[145]) & ~(inputs[834]);
    assign layer0_outputs[159] = (inputs[31]) ^ (inputs[339]);
    assign layer0_outputs[160] = ~(inputs[747]);
    assign layer0_outputs[161] = inputs[511];
    assign layer0_outputs[162] = ~((inputs[544]) | (inputs[488]));
    assign layer0_outputs[163] = ~((inputs[535]) ^ (inputs[600]));
    assign layer0_outputs[164] = ~((inputs[884]) | (inputs[848]));
    assign layer0_outputs[165] = (inputs[112]) ^ (inputs[963]);
    assign layer0_outputs[166] = (inputs[374]) ^ (inputs[37]);
    assign layer0_outputs[167] = ~((inputs[763]) | (inputs[100]));
    assign layer0_outputs[168] = inputs[331];
    assign layer0_outputs[169] = (inputs[275]) & ~(inputs[288]);
    assign layer0_outputs[170] = ~((inputs[574]) ^ (inputs[792]));
    assign layer0_outputs[171] = inputs[620];
    assign layer0_outputs[172] = (inputs[810]) & ~(inputs[507]);
    assign layer0_outputs[173] = ~((inputs[314]) | (inputs[861]));
    assign layer0_outputs[174] = (inputs[565]) | (inputs[29]);
    assign layer0_outputs[175] = ~(inputs[962]) | (inputs[802]);
    assign layer0_outputs[176] = ~((inputs[619]) | (inputs[956]));
    assign layer0_outputs[177] = ~(inputs[224]);
    assign layer0_outputs[178] = inputs[514];
    assign layer0_outputs[179] = (inputs[556]) | (inputs[790]);
    assign layer0_outputs[180] = inputs[591];
    assign layer0_outputs[181] = 1'b0;
    assign layer0_outputs[182] = inputs[672];
    assign layer0_outputs[183] = ~((inputs[818]) | (inputs[290]));
    assign layer0_outputs[184] = (inputs[370]) & ~(inputs[647]);
    assign layer0_outputs[185] = (inputs[335]) | (inputs[57]);
    assign layer0_outputs[186] = (inputs[575]) & (inputs[291]);
    assign layer0_outputs[187] = ~(inputs[364]);
    assign layer0_outputs[188] = ~((inputs[76]) | (inputs[254]));
    assign layer0_outputs[189] = ~((inputs[12]) | (inputs[473]));
    assign layer0_outputs[190] = inputs[663];
    assign layer0_outputs[191] = (inputs[854]) & ~(inputs[163]);
    assign layer0_outputs[192] = ~((inputs[484]) & (inputs[182]));
    assign layer0_outputs[193] = (inputs[607]) & (inputs[153]);
    assign layer0_outputs[194] = (inputs[892]) & (inputs[857]);
    assign layer0_outputs[195] = inputs[490];
    assign layer0_outputs[196] = ~(inputs[491]) | (inputs[438]);
    assign layer0_outputs[197] = ~((inputs[234]) | (inputs[584]));
    assign layer0_outputs[198] = (inputs[974]) & (inputs[1017]);
    assign layer0_outputs[199] = (inputs[363]) & ~(inputs[293]);
    assign layer0_outputs[200] = (inputs[450]) | (inputs[171]);
    assign layer0_outputs[201] = ~(inputs[848]);
    assign layer0_outputs[202] = (inputs[805]) & (inputs[691]);
    assign layer0_outputs[203] = inputs[677];
    assign layer0_outputs[204] = (inputs[836]) | (inputs[228]);
    assign layer0_outputs[205] = (inputs[51]) & ~(inputs[123]);
    assign layer0_outputs[206] = ~((inputs[603]) | (inputs[437]));
    assign layer0_outputs[207] = 1'b1;
    assign layer0_outputs[208] = inputs[651];
    assign layer0_outputs[209] = (inputs[1018]) | (inputs[369]);
    assign layer0_outputs[210] = ~(inputs[664]) | (inputs[947]);
    assign layer0_outputs[211] = (inputs[462]) & ~(inputs[803]);
    assign layer0_outputs[212] = ~((inputs[776]) | (inputs[494]));
    assign layer0_outputs[213] = (inputs[600]) & ~(inputs[837]);
    assign layer0_outputs[214] = inputs[537];
    assign layer0_outputs[215] = ~((inputs[77]) ^ (inputs[119]));
    assign layer0_outputs[216] = ~((inputs[915]) ^ (inputs[317]));
    assign layer0_outputs[217] = inputs[509];
    assign layer0_outputs[218] = ~((inputs[748]) & (inputs[780]));
    assign layer0_outputs[219] = inputs[881];
    assign layer0_outputs[220] = inputs[591];
    assign layer0_outputs[221] = (inputs[789]) ^ (inputs[86]);
    assign layer0_outputs[222] = ~(inputs[392]);
    assign layer0_outputs[223] = ~(inputs[195]);
    assign layer0_outputs[224] = inputs[665];
    assign layer0_outputs[225] = (inputs[362]) & (inputs[30]);
    assign layer0_outputs[226] = inputs[926];
    assign layer0_outputs[227] = inputs[115];
    assign layer0_outputs[228] = ~(inputs[810]);
    assign layer0_outputs[229] = ~(inputs[523]) | (inputs[838]);
    assign layer0_outputs[230] = 1'b0;
    assign layer0_outputs[231] = ~((inputs[187]) | (inputs[880]));
    assign layer0_outputs[232] = ~(inputs[845]);
    assign layer0_outputs[233] = ~((inputs[773]) | (inputs[137]));
    assign layer0_outputs[234] = 1'b1;
    assign layer0_outputs[235] = (inputs[990]) | (inputs[989]);
    assign layer0_outputs[236] = (inputs[22]) | (inputs[807]);
    assign layer0_outputs[237] = (inputs[287]) & ~(inputs[887]);
    assign layer0_outputs[238] = ~(inputs[436]);
    assign layer0_outputs[239] = ~((inputs[337]) ^ (inputs[242]));
    assign layer0_outputs[240] = (inputs[506]) | (inputs[1008]);
    assign layer0_outputs[241] = ~((inputs[267]) | (inputs[482]));
    assign layer0_outputs[242] = ~((inputs[488]) | (inputs[361]));
    assign layer0_outputs[243] = (inputs[493]) & ~(inputs[869]);
    assign layer0_outputs[244] = inputs[141];
    assign layer0_outputs[245] = inputs[492];
    assign layer0_outputs[246] = ~((inputs[945]) ^ (inputs[691]));
    assign layer0_outputs[247] = ~(inputs[683]);
    assign layer0_outputs[248] = 1'b0;
    assign layer0_outputs[249] = (inputs[710]) ^ (inputs[469]);
    assign layer0_outputs[250] = ~((inputs[832]) ^ (inputs[402]));
    assign layer0_outputs[251] = ~((inputs[674]) | (inputs[686]));
    assign layer0_outputs[252] = ~(inputs[171]);
    assign layer0_outputs[253] = ~(inputs[546]);
    assign layer0_outputs[254] = ~((inputs[700]) | (inputs[108]));
    assign layer0_outputs[255] = ~(inputs[437]);
    assign layer0_outputs[256] = ~((inputs[103]) | (inputs[621]));
    assign layer0_outputs[257] = (inputs[296]) & ~(inputs[1]);
    assign layer0_outputs[258] = ~(inputs[571]);
    assign layer0_outputs[259] = inputs[140];
    assign layer0_outputs[260] = ~((inputs[682]) ^ (inputs[98]));
    assign layer0_outputs[261] = ~(inputs[522]);
    assign layer0_outputs[262] = ~(inputs[474]);
    assign layer0_outputs[263] = ~((inputs[666]) | (inputs[879]));
    assign layer0_outputs[264] = 1'b0;
    assign layer0_outputs[265] = ~((inputs[987]) | (inputs[201]));
    assign layer0_outputs[266] = ~((inputs[380]) | (inputs[693]));
    assign layer0_outputs[267] = (inputs[333]) ^ (inputs[932]);
    assign layer0_outputs[268] = ~((inputs[544]) & (inputs[657]));
    assign layer0_outputs[269] = ~((inputs[843]) | (inputs[553]));
    assign layer0_outputs[270] = (inputs[619]) | (inputs[140]);
    assign layer0_outputs[271] = ~((inputs[209]) | (inputs[819]));
    assign layer0_outputs[272] = inputs[557];
    assign layer0_outputs[273] = ~(inputs[519]);
    assign layer0_outputs[274] = ~(inputs[340]);
    assign layer0_outputs[275] = (inputs[256]) & ~(inputs[967]);
    assign layer0_outputs[276] = (inputs[985]) & ~(inputs[959]);
    assign layer0_outputs[277] = inputs[313];
    assign layer0_outputs[278] = inputs[172];
    assign layer0_outputs[279] = (inputs[801]) | (inputs[1012]);
    assign layer0_outputs[280] = (inputs[588]) & ~(inputs[76]);
    assign layer0_outputs[281] = (inputs[589]) & ~(inputs[515]);
    assign layer0_outputs[282] = (inputs[554]) & ~(inputs[643]);
    assign layer0_outputs[283] = ~(inputs[807]) | (inputs[322]);
    assign layer0_outputs[284] = ~(inputs[620]) | (inputs[941]);
    assign layer0_outputs[285] = ~((inputs[121]) ^ (inputs[804]));
    assign layer0_outputs[286] = ~((inputs[539]) | (inputs[323]));
    assign layer0_outputs[287] = ~(inputs[231]) | (inputs[548]);
    assign layer0_outputs[288] = inputs[782];
    assign layer0_outputs[289] = 1'b1;
    assign layer0_outputs[290] = (inputs[506]) & ~(inputs[296]);
    assign layer0_outputs[291] = ~((inputs[238]) | (inputs[203]));
    assign layer0_outputs[292] = inputs[275];
    assign layer0_outputs[293] = (inputs[584]) | (inputs[160]);
    assign layer0_outputs[294] = inputs[620];
    assign layer0_outputs[295] = ~((inputs[840]) | (inputs[880]));
    assign layer0_outputs[296] = (inputs[817]) ^ (inputs[612]);
    assign layer0_outputs[297] = ~(inputs[216]);
    assign layer0_outputs[298] = ~((inputs[797]) | (inputs[61]));
    assign layer0_outputs[299] = (inputs[626]) & ~(inputs[841]);
    assign layer0_outputs[300] = 1'b1;
    assign layer0_outputs[301] = (inputs[555]) ^ (inputs[230]);
    assign layer0_outputs[302] = (inputs[1000]) | (inputs[624]);
    assign layer0_outputs[303] = (inputs[376]) & ~(inputs[645]);
    assign layer0_outputs[304] = inputs[567];
    assign layer0_outputs[305] = (inputs[436]) | (inputs[306]);
    assign layer0_outputs[306] = inputs[427];
    assign layer0_outputs[307] = ~(inputs[758]);
    assign layer0_outputs[308] = (inputs[749]) ^ (inputs[755]);
    assign layer0_outputs[309] = ~((inputs[440]) | (inputs[613]));
    assign layer0_outputs[310] = 1'b1;
    assign layer0_outputs[311] = 1'b0;
    assign layer0_outputs[312] = (inputs[713]) | (inputs[647]);
    assign layer0_outputs[313] = (inputs[307]) | (inputs[577]);
    assign layer0_outputs[314] = (inputs[30]) & ~(inputs[190]);
    assign layer0_outputs[315] = (inputs[742]) & ~(inputs[966]);
    assign layer0_outputs[316] = (inputs[775]) & ~(inputs[157]);
    assign layer0_outputs[317] = (inputs[509]) & ~(inputs[669]);
    assign layer0_outputs[318] = 1'b1;
    assign layer0_outputs[319] = inputs[275];
    assign layer0_outputs[320] = ~((inputs[156]) | (inputs[6]));
    assign layer0_outputs[321] = (inputs[263]) | (inputs[302]);
    assign layer0_outputs[322] = ~(inputs[557]);
    assign layer0_outputs[323] = ~(inputs[534]);
    assign layer0_outputs[324] = ~((inputs[526]) | (inputs[494]));
    assign layer0_outputs[325] = ~((inputs[730]) | (inputs[261]));
    assign layer0_outputs[326] = (inputs[954]) ^ (inputs[491]);
    assign layer0_outputs[327] = (inputs[413]) ^ (inputs[344]);
    assign layer0_outputs[328] = ~((inputs[842]) ^ (inputs[992]));
    assign layer0_outputs[329] = ~(inputs[492]) | (inputs[547]);
    assign layer0_outputs[330] = ~((inputs[641]) | (inputs[968]));
    assign layer0_outputs[331] = inputs[810];
    assign layer0_outputs[332] = inputs[16];
    assign layer0_outputs[333] = ~(inputs[914]) | (inputs[39]);
    assign layer0_outputs[334] = ~(inputs[359]);
    assign layer0_outputs[335] = ~(inputs[69]);
    assign layer0_outputs[336] = (inputs[121]) & ~(inputs[994]);
    assign layer0_outputs[337] = (inputs[164]) ^ (inputs[356]);
    assign layer0_outputs[338] = (inputs[654]) | (inputs[803]);
    assign layer0_outputs[339] = (inputs[59]) & ~(inputs[701]);
    assign layer0_outputs[340] = (inputs[720]) | (inputs[515]);
    assign layer0_outputs[341] = (inputs[486]) & ~(inputs[1023]);
    assign layer0_outputs[342] = (inputs[336]) & (inputs[587]);
    assign layer0_outputs[343] = ~(inputs[588]);
    assign layer0_outputs[344] = ~((inputs[602]) | (inputs[733]));
    assign layer0_outputs[345] = (inputs[382]) & ~(inputs[10]);
    assign layer0_outputs[346] = ~((inputs[559]) ^ (inputs[707]));
    assign layer0_outputs[347] = (inputs[655]) ^ (inputs[51]);
    assign layer0_outputs[348] = ~((inputs[125]) ^ (inputs[387]));
    assign layer0_outputs[349] = (inputs[870]) ^ (inputs[511]);
    assign layer0_outputs[350] = ~((inputs[842]) ^ (inputs[784]));
    assign layer0_outputs[351] = ~(inputs[621]) | (inputs[701]);
    assign layer0_outputs[352] = (inputs[765]) & (inputs[99]);
    assign layer0_outputs[353] = (inputs[469]) ^ (inputs[599]);
    assign layer0_outputs[354] = ~((inputs[772]) | (inputs[341]));
    assign layer0_outputs[355] = (inputs[762]) & ~(inputs[25]);
    assign layer0_outputs[356] = ~(inputs[393]);
    assign layer0_outputs[357] = inputs[491];
    assign layer0_outputs[358] = (inputs[820]) & ~(inputs[68]);
    assign layer0_outputs[359] = (inputs[346]) ^ (inputs[23]);
    assign layer0_outputs[360] = ~((inputs[460]) ^ (inputs[354]));
    assign layer0_outputs[361] = ~((inputs[606]) & (inputs[768]));
    assign layer0_outputs[362] = (inputs[181]) | (inputs[505]);
    assign layer0_outputs[363] = ~(inputs[145]);
    assign layer0_outputs[364] = (inputs[97]) ^ (inputs[365]);
    assign layer0_outputs[365] = (inputs[821]) ^ (inputs[575]);
    assign layer0_outputs[366] = ~(inputs[820]);
    assign layer0_outputs[367] = ~(inputs[299]) | (inputs[99]);
    assign layer0_outputs[368] = (inputs[636]) | (inputs[985]);
    assign layer0_outputs[369] = inputs[786];
    assign layer0_outputs[370] = ~((inputs[653]) ^ (inputs[451]));
    assign layer0_outputs[371] = inputs[885];
    assign layer0_outputs[372] = (inputs[443]) | (inputs[696]);
    assign layer0_outputs[373] = ~(inputs[169]) | (inputs[386]);
    assign layer0_outputs[374] = ~((inputs[47]) ^ (inputs[1012]));
    assign layer0_outputs[375] = ~((inputs[517]) | (inputs[363]));
    assign layer0_outputs[376] = ~((inputs[480]) | (inputs[770]));
    assign layer0_outputs[377] = ~((inputs[527]) & (inputs[932]));
    assign layer0_outputs[378] = ~((inputs[303]) & (inputs[457]));
    assign layer0_outputs[379] = inputs[841];
    assign layer0_outputs[380] = inputs[812];
    assign layer0_outputs[381] = ~(inputs[900]);
    assign layer0_outputs[382] = (inputs[90]) | (inputs[384]);
    assign layer0_outputs[383] = ~((inputs[782]) & (inputs[273]));
    assign layer0_outputs[384] = (inputs[498]) & ~(inputs[56]);
    assign layer0_outputs[385] = inputs[891];
    assign layer0_outputs[386] = ~((inputs[532]) ^ (inputs[928]));
    assign layer0_outputs[387] = ~((inputs[158]) | (inputs[913]));
    assign layer0_outputs[388] = inputs[851];
    assign layer0_outputs[389] = ~((inputs[347]) | (inputs[422]));
    assign layer0_outputs[390] = inputs[401];
    assign layer0_outputs[391] = (inputs[968]) | (inputs[880]);
    assign layer0_outputs[392] = ~((inputs[595]) ^ (inputs[960]));
    assign layer0_outputs[393] = inputs[496];
    assign layer0_outputs[394] = (inputs[232]) & ~(inputs[386]);
    assign layer0_outputs[395] = (inputs[815]) & ~(inputs[976]);
    assign layer0_outputs[396] = (inputs[556]) & ~(inputs[190]);
    assign layer0_outputs[397] = ~(inputs[429]) | (inputs[842]);
    assign layer0_outputs[398] = ~((inputs[353]) | (inputs[365]));
    assign layer0_outputs[399] = (inputs[302]) & ~(inputs[811]);
    assign layer0_outputs[400] = (inputs[236]) ^ (inputs[599]);
    assign layer0_outputs[401] = ~(inputs[597]) | (inputs[530]);
    assign layer0_outputs[402] = (inputs[790]) & ~(inputs[47]);
    assign layer0_outputs[403] = (inputs[560]) & ~(inputs[761]);
    assign layer0_outputs[404] = ~(inputs[225]) | (inputs[159]);
    assign layer0_outputs[405] = 1'b1;
    assign layer0_outputs[406] = (inputs[886]) & ~(inputs[555]);
    assign layer0_outputs[407] = (inputs[777]) | (inputs[46]);
    assign layer0_outputs[408] = (inputs[125]) & (inputs[900]);
    assign layer0_outputs[409] = ~(inputs[970]);
    assign layer0_outputs[410] = inputs[617];
    assign layer0_outputs[411] = ~((inputs[636]) | (inputs[1022]));
    assign layer0_outputs[412] = inputs[473];
    assign layer0_outputs[413] = 1'b1;
    assign layer0_outputs[414] = inputs[32];
    assign layer0_outputs[415] = inputs[240];
    assign layer0_outputs[416] = (inputs[399]) | (inputs[661]);
    assign layer0_outputs[417] = (inputs[255]) & ~(inputs[498]);
    assign layer0_outputs[418] = inputs[228];
    assign layer0_outputs[419] = (inputs[562]) & ~(inputs[838]);
    assign layer0_outputs[420] = inputs[240];
    assign layer0_outputs[421] = ~(inputs[820]) | (inputs[186]);
    assign layer0_outputs[422] = ~(inputs[600]) | (inputs[309]);
    assign layer0_outputs[423] = ~((inputs[29]) | (inputs[80]));
    assign layer0_outputs[424] = ~((inputs[592]) | (inputs[638]));
    assign layer0_outputs[425] = inputs[178];
    assign layer0_outputs[426] = ~((inputs[56]) ^ (inputs[430]));
    assign layer0_outputs[427] = ~(inputs[707]);
    assign layer0_outputs[428] = ~((inputs[9]) | (inputs[532]));
    assign layer0_outputs[429] = (inputs[395]) | (inputs[127]);
    assign layer0_outputs[430] = ~((inputs[459]) ^ (inputs[831]));
    assign layer0_outputs[431] = ~((inputs[59]) | (inputs[64]));
    assign layer0_outputs[432] = (inputs[933]) & ~(inputs[187]);
    assign layer0_outputs[433] = ~((inputs[938]) | (inputs[241]));
    assign layer0_outputs[434] = ~(inputs[615]) | (inputs[317]);
    assign layer0_outputs[435] = (inputs[191]) ^ (inputs[126]);
    assign layer0_outputs[436] = ~((inputs[384]) | (inputs[272]));
    assign layer0_outputs[437] = (inputs[609]) & ~(inputs[970]);
    assign layer0_outputs[438] = ~(inputs[483]);
    assign layer0_outputs[439] = ~(inputs[257]) | (inputs[434]);
    assign layer0_outputs[440] = ~(inputs[503]);
    assign layer0_outputs[441] = (inputs[600]) & ~(inputs[114]);
    assign layer0_outputs[442] = ~(inputs[229]) | (inputs[15]);
    assign layer0_outputs[443] = (inputs[461]) | (inputs[867]);
    assign layer0_outputs[444] = (inputs[810]) & ~(inputs[405]);
    assign layer0_outputs[445] = ~(inputs[202]) | (inputs[124]);
    assign layer0_outputs[446] = (inputs[254]) ^ (inputs[504]);
    assign layer0_outputs[447] = inputs[924];
    assign layer0_outputs[448] = ~((inputs[191]) | (inputs[58]));
    assign layer0_outputs[449] = (inputs[524]) ^ (inputs[995]);
    assign layer0_outputs[450] = ~((inputs[846]) ^ (inputs[295]));
    assign layer0_outputs[451] = ~(inputs[472]);
    assign layer0_outputs[452] = ~((inputs[816]) ^ (inputs[1014]));
    assign layer0_outputs[453] = ~((inputs[518]) | (inputs[691]));
    assign layer0_outputs[454] = ~(inputs[742]);
    assign layer0_outputs[455] = ~(inputs[335]) | (inputs[482]);
    assign layer0_outputs[456] = (inputs[528]) & ~(inputs[1000]);
    assign layer0_outputs[457] = (inputs[268]) & ~(inputs[162]);
    assign layer0_outputs[458] = ~((inputs[172]) ^ (inputs[936]));
    assign layer0_outputs[459] = ~(inputs[683]) | (inputs[370]);
    assign layer0_outputs[460] = (inputs[435]) & ~(inputs[315]);
    assign layer0_outputs[461] = ~((inputs[984]) | (inputs[231]));
    assign layer0_outputs[462] = 1'b0;
    assign layer0_outputs[463] = ~(inputs[698]) | (inputs[880]);
    assign layer0_outputs[464] = 1'b0;
    assign layer0_outputs[465] = inputs[792];
    assign layer0_outputs[466] = (inputs[872]) | (inputs[219]);
    assign layer0_outputs[467] = (inputs[202]) & ~(inputs[876]);
    assign layer0_outputs[468] = (inputs[232]) ^ (inputs[85]);
    assign layer0_outputs[469] = (inputs[864]) | (inputs[440]);
    assign layer0_outputs[470] = ~(inputs[291]) | (inputs[221]);
    assign layer0_outputs[471] = inputs[416];
    assign layer0_outputs[472] = ~(inputs[463]);
    assign layer0_outputs[473] = (inputs[296]) | (inputs[759]);
    assign layer0_outputs[474] = ~((inputs[264]) ^ (inputs[647]));
    assign layer0_outputs[475] = ~((inputs[744]) | (inputs[83]));
    assign layer0_outputs[476] = (inputs[253]) | (inputs[377]);
    assign layer0_outputs[477] = ~((inputs[674]) & (inputs[676]));
    assign layer0_outputs[478] = (inputs[849]) & ~(inputs[139]);
    assign layer0_outputs[479] = ~(inputs[884]);
    assign layer0_outputs[480] = (inputs[658]) & ~(inputs[741]);
    assign layer0_outputs[481] = ~((inputs[213]) | (inputs[235]));
    assign layer0_outputs[482] = inputs[339];
    assign layer0_outputs[483] = (inputs[366]) & ~(inputs[420]);
    assign layer0_outputs[484] = inputs[728];
    assign layer0_outputs[485] = ~(inputs[939]);
    assign layer0_outputs[486] = (inputs[868]) ^ (inputs[984]);
    assign layer0_outputs[487] = (inputs[696]) & ~(inputs[627]);
    assign layer0_outputs[488] = ~(inputs[226]) | (inputs[294]);
    assign layer0_outputs[489] = ~(inputs[200]) | (inputs[1000]);
    assign layer0_outputs[490] = (inputs[468]) & ~(inputs[76]);
    assign layer0_outputs[491] = ~((inputs[768]) ^ (inputs[856]));
    assign layer0_outputs[492] = (inputs[763]) | (inputs[806]);
    assign layer0_outputs[493] = (inputs[710]) & ~(inputs[1005]);
    assign layer0_outputs[494] = (inputs[10]) & ~(inputs[733]);
    assign layer0_outputs[495] = (inputs[373]) & ~(inputs[24]);
    assign layer0_outputs[496] = ~((inputs[354]) | (inputs[503]));
    assign layer0_outputs[497] = (inputs[956]) ^ (inputs[329]);
    assign layer0_outputs[498] = inputs[502];
    assign layer0_outputs[499] = (inputs[682]) & ~(inputs[829]);
    assign layer0_outputs[500] = ~((inputs[262]) | (inputs[447]));
    assign layer0_outputs[501] = ~(inputs[759]) | (inputs[661]);
    assign layer0_outputs[502] = (inputs[275]) ^ (inputs[749]);
    assign layer0_outputs[503] = (inputs[460]) & ~(inputs[438]);
    assign layer0_outputs[504] = (inputs[920]) ^ (inputs[876]);
    assign layer0_outputs[505] = ~(inputs[434]) | (inputs[443]);
    assign layer0_outputs[506] = ~(inputs[565]) | (inputs[127]);
    assign layer0_outputs[507] = ~(inputs[358]) | (inputs[319]);
    assign layer0_outputs[508] = ~(inputs[173]) | (inputs[998]);
    assign layer0_outputs[509] = (inputs[746]) ^ (inputs[264]);
    assign layer0_outputs[510] = ~(inputs[95]) | (inputs[416]);
    assign layer0_outputs[511] = (inputs[12]) ^ (inputs[625]);
    assign layer0_outputs[512] = (inputs[907]) | (inputs[1006]);
    assign layer0_outputs[513] = ~((inputs[112]) ^ (inputs[180]));
    assign layer0_outputs[514] = inputs[71];
    assign layer0_outputs[515] = (inputs[940]) | (inputs[403]);
    assign layer0_outputs[516] = (inputs[283]) | (inputs[286]);
    assign layer0_outputs[517] = ~((inputs[286]) & (inputs[785]));
    assign layer0_outputs[518] = ~(inputs[456]);
    assign layer0_outputs[519] = (inputs[118]) ^ (inputs[734]);
    assign layer0_outputs[520] = ~((inputs[1001]) ^ (inputs[80]));
    assign layer0_outputs[521] = (inputs[911]) | (inputs[55]);
    assign layer0_outputs[522] = ~((inputs[823]) ^ (inputs[445]));
    assign layer0_outputs[523] = inputs[3];
    assign layer0_outputs[524] = inputs[248];
    assign layer0_outputs[525] = 1'b0;
    assign layer0_outputs[526] = ~((inputs[211]) ^ (inputs[766]));
    assign layer0_outputs[527] = (inputs[695]) ^ (inputs[900]);
    assign layer0_outputs[528] = ~(inputs[296]);
    assign layer0_outputs[529] = ~((inputs[130]) | (inputs[366]));
    assign layer0_outputs[530] = ~((inputs[813]) | (inputs[696]));
    assign layer0_outputs[531] = (inputs[344]) ^ (inputs[770]);
    assign layer0_outputs[532] = (inputs[935]) ^ (inputs[251]);
    assign layer0_outputs[533] = ~(inputs[778]) | (inputs[594]);
    assign layer0_outputs[534] = ~((inputs[256]) | (inputs[306]));
    assign layer0_outputs[535] = ~((inputs[145]) | (inputs[662]));
    assign layer0_outputs[536] = inputs[279];
    assign layer0_outputs[537] = (inputs[1002]) ^ (inputs[52]);
    assign layer0_outputs[538] = (inputs[39]) & (inputs[873]);
    assign layer0_outputs[539] = ~(inputs[754]);
    assign layer0_outputs[540] = inputs[715];
    assign layer0_outputs[541] = ~(inputs[218]) | (inputs[643]);
    assign layer0_outputs[542] = ~(inputs[163]);
    assign layer0_outputs[543] = (inputs[447]) | (inputs[599]);
    assign layer0_outputs[544] = (inputs[982]) | (inputs[500]);
    assign layer0_outputs[545] = (inputs[19]) ^ (inputs[661]);
    assign layer0_outputs[546] = ~(inputs[621]) | (inputs[829]);
    assign layer0_outputs[547] = inputs[782];
    assign layer0_outputs[548] = ~((inputs[540]) | (inputs[355]));
    assign layer0_outputs[549] = ~(inputs[278]);
    assign layer0_outputs[550] = ~((inputs[208]) | (inputs[176]));
    assign layer0_outputs[551] = (inputs[661]) & ~(inputs[285]);
    assign layer0_outputs[552] = (inputs[909]) & ~(inputs[999]);
    assign layer0_outputs[553] = ~(inputs[250]) | (inputs[607]);
    assign layer0_outputs[554] = (inputs[724]) & ~(inputs[898]);
    assign layer0_outputs[555] = (inputs[511]) & ~(inputs[166]);
    assign layer0_outputs[556] = (inputs[939]) ^ (inputs[157]);
    assign layer0_outputs[557] = (inputs[222]) ^ (inputs[455]);
    assign layer0_outputs[558] = (inputs[644]) ^ (inputs[856]);
    assign layer0_outputs[559] = 1'b0;
    assign layer0_outputs[560] = ~((inputs[172]) ^ (inputs[826]));
    assign layer0_outputs[561] = ~((inputs[992]) & (inputs[548]));
    assign layer0_outputs[562] = ~(inputs[167]);
    assign layer0_outputs[563] = ~((inputs[769]) ^ (inputs[616]));
    assign layer0_outputs[564] = ~(inputs[683]) | (inputs[1004]);
    assign layer0_outputs[565] = inputs[746];
    assign layer0_outputs[566] = ~(inputs[526]) | (inputs[46]);
    assign layer0_outputs[567] = (inputs[491]) & ~(inputs[263]);
    assign layer0_outputs[568] = ~(inputs[300]) | (inputs[136]);
    assign layer0_outputs[569] = (inputs[289]) | (inputs[433]);
    assign layer0_outputs[570] = ~((inputs[1005]) | (inputs[308]));
    assign layer0_outputs[571] = (inputs[317]) ^ (inputs[613]);
    assign layer0_outputs[572] = (inputs[327]) ^ (inputs[140]);
    assign layer0_outputs[573] = ~(inputs[647]) | (inputs[983]);
    assign layer0_outputs[574] = (inputs[216]) & ~(inputs[148]);
    assign layer0_outputs[575] = (inputs[269]) ^ (inputs[92]);
    assign layer0_outputs[576] = ~(inputs[366]);
    assign layer0_outputs[577] = ~((inputs[457]) | (inputs[54]));
    assign layer0_outputs[578] = ~((inputs[307]) | (inputs[909]));
    assign layer0_outputs[579] = ~((inputs[860]) ^ (inputs[913]));
    assign layer0_outputs[580] = (inputs[774]) & ~(inputs[839]);
    assign layer0_outputs[581] = 1'b0;
    assign layer0_outputs[582] = inputs[825];
    assign layer0_outputs[583] = (inputs[204]) & ~(inputs[802]);
    assign layer0_outputs[584] = (inputs[263]) ^ (inputs[671]);
    assign layer0_outputs[585] = (inputs[663]) | (inputs[898]);
    assign layer0_outputs[586] = (inputs[972]) | (inputs[555]);
    assign layer0_outputs[587] = inputs[203];
    assign layer0_outputs[588] = ~(inputs[56]) | (inputs[867]);
    assign layer0_outputs[589] = ~((inputs[28]) ^ (inputs[247]));
    assign layer0_outputs[590] = inputs[307];
    assign layer0_outputs[591] = ~((inputs[803]) ^ (inputs[727]));
    assign layer0_outputs[592] = (inputs[570]) | (inputs[52]);
    assign layer0_outputs[593] = ~((inputs[317]) | (inputs[306]));
    assign layer0_outputs[594] = ~(inputs[943]);
    assign layer0_outputs[595] = ~((inputs[596]) | (inputs[922]));
    assign layer0_outputs[596] = (inputs[407]) & ~(inputs[263]);
    assign layer0_outputs[597] = (inputs[657]) & ~(inputs[455]);
    assign layer0_outputs[598] = ~((inputs[753]) ^ (inputs[385]));
    assign layer0_outputs[599] = (inputs[817]) & ~(inputs[977]);
    assign layer0_outputs[600] = ~((inputs[955]) | (inputs[916]));
    assign layer0_outputs[601] = ~((inputs[135]) | (inputs[599]));
    assign layer0_outputs[602] = (inputs[478]) & ~(inputs[71]);
    assign layer0_outputs[603] = ~((inputs[806]) | (inputs[112]));
    assign layer0_outputs[604] = ~((inputs[799]) | (inputs[487]));
    assign layer0_outputs[605] = (inputs[692]) & ~(inputs[503]);
    assign layer0_outputs[606] = (inputs[402]) | (inputs[118]);
    assign layer0_outputs[607] = ~(inputs[500]);
    assign layer0_outputs[608] = (inputs[300]) | (inputs[5]);
    assign layer0_outputs[609] = ~((inputs[866]) | (inputs[53]));
    assign layer0_outputs[610] = (inputs[672]) & (inputs[999]);
    assign layer0_outputs[611] = ~(inputs[408]);
    assign layer0_outputs[612] = (inputs[418]) | (inputs[637]);
    assign layer0_outputs[613] = ~((inputs[644]) | (inputs[813]));
    assign layer0_outputs[614] = (inputs[54]) & ~(inputs[136]);
    assign layer0_outputs[615] = ~((inputs[951]) | (inputs[595]));
    assign layer0_outputs[616] = (inputs[289]) & (inputs[921]);
    assign layer0_outputs[617] = inputs[792];
    assign layer0_outputs[618] = ~(inputs[1011]) | (inputs[65]);
    assign layer0_outputs[619] = ~((inputs[981]) | (inputs[93]));
    assign layer0_outputs[620] = ~((inputs[868]) ^ (inputs[557]));
    assign layer0_outputs[621] = ~((inputs[342]) | (inputs[96]));
    assign layer0_outputs[622] = ~(inputs[846]);
    assign layer0_outputs[623] = ~(inputs[745]) | (inputs[479]);
    assign layer0_outputs[624] = ~((inputs[88]) | (inputs[485]));
    assign layer0_outputs[625] = (inputs[133]) | (inputs[39]);
    assign layer0_outputs[626] = ~(inputs[501]);
    assign layer0_outputs[627] = (inputs[558]) & ~(inputs[1021]);
    assign layer0_outputs[628] = (inputs[1005]) & ~(inputs[82]);
    assign layer0_outputs[629] = ~((inputs[804]) & (inputs[201]));
    assign layer0_outputs[630] = inputs[805];
    assign layer0_outputs[631] = (inputs[622]) & ~(inputs[505]);
    assign layer0_outputs[632] = inputs[474];
    assign layer0_outputs[633] = (inputs[500]) | (inputs[584]);
    assign layer0_outputs[634] = inputs[432];
    assign layer0_outputs[635] = (inputs[516]) & (inputs[628]);
    assign layer0_outputs[636] = ~(inputs[215]) | (inputs[376]);
    assign layer0_outputs[637] = ~((inputs[1019]) | (inputs[878]));
    assign layer0_outputs[638] = (inputs[170]) ^ (inputs[615]);
    assign layer0_outputs[639] = ~((inputs[566]) | (inputs[397]));
    assign layer0_outputs[640] = inputs[186];
    assign layer0_outputs[641] = ~(inputs[873]) | (inputs[168]);
    assign layer0_outputs[642] = inputs[133];
    assign layer0_outputs[643] = (inputs[509]) | (inputs[591]);
    assign layer0_outputs[644] = (inputs[582]) & ~(inputs[2]);
    assign layer0_outputs[645] = ~((inputs[711]) ^ (inputs[173]));
    assign layer0_outputs[646] = (inputs[627]) & ~(inputs[679]);
    assign layer0_outputs[647] = ~((inputs[952]) & (inputs[712]));
    assign layer0_outputs[648] = inputs[609];
    assign layer0_outputs[649] = inputs[151];
    assign layer0_outputs[650] = ~(inputs[355]) | (inputs[218]);
    assign layer0_outputs[651] = ~((inputs[429]) | (inputs[576]));
    assign layer0_outputs[652] = ~((inputs[794]) ^ (inputs[410]));
    assign layer0_outputs[653] = (inputs[588]) | (inputs[149]);
    assign layer0_outputs[654] = inputs[490];
    assign layer0_outputs[655] = (inputs[723]) | (inputs[257]);
    assign layer0_outputs[656] = ~(inputs[497]);
    assign layer0_outputs[657] = ~(inputs[499]);
    assign layer0_outputs[658] = (inputs[787]) | (inputs[552]);
    assign layer0_outputs[659] = (inputs[63]) | (inputs[742]);
    assign layer0_outputs[660] = 1'b1;
    assign layer0_outputs[661] = ~(inputs[121]);
    assign layer0_outputs[662] = ~(inputs[966]);
    assign layer0_outputs[663] = inputs[507];
    assign layer0_outputs[664] = ~((inputs[300]) | (inputs[827]));
    assign layer0_outputs[665] = (inputs[759]) ^ (inputs[521]);
    assign layer0_outputs[666] = (inputs[693]) & ~(inputs[769]);
    assign layer0_outputs[667] = (inputs[830]) ^ (inputs[247]);
    assign layer0_outputs[668] = ~(inputs[816]);
    assign layer0_outputs[669] = inputs[301];
    assign layer0_outputs[670] = inputs[16];
    assign layer0_outputs[671] = ~(inputs[830]) | (inputs[997]);
    assign layer0_outputs[672] = (inputs[373]) & ~(inputs[548]);
    assign layer0_outputs[673] = ~((inputs[1019]) | (inputs[36]));
    assign layer0_outputs[674] = ~((inputs[14]) | (inputs[806]));
    assign layer0_outputs[675] = ~((inputs[321]) ^ (inputs[941]));
    assign layer0_outputs[676] = (inputs[528]) & ~(inputs[698]);
    assign layer0_outputs[677] = ~(inputs[500]) | (inputs[571]);
    assign layer0_outputs[678] = (inputs[845]) & ~(inputs[190]);
    assign layer0_outputs[679] = ~(inputs[996]);
    assign layer0_outputs[680] = (inputs[217]) & ~(inputs[998]);
    assign layer0_outputs[681] = ~((inputs[940]) ^ (inputs[150]));
    assign layer0_outputs[682] = (inputs[539]) ^ (inputs[12]);
    assign layer0_outputs[683] = inputs[538];
    assign layer0_outputs[684] = (inputs[12]) ^ (inputs[172]);
    assign layer0_outputs[685] = ~((inputs[200]) | (inputs[818]));
    assign layer0_outputs[686] = inputs[306];
    assign layer0_outputs[687] = ~((inputs[869]) | (inputs[818]));
    assign layer0_outputs[688] = ~(inputs[338]) | (inputs[615]);
    assign layer0_outputs[689] = ~((inputs[368]) ^ (inputs[449]));
    assign layer0_outputs[690] = inputs[419];
    assign layer0_outputs[691] = ~((inputs[764]) | (inputs[619]));
    assign layer0_outputs[692] = ~(inputs[362]);
    assign layer0_outputs[693] = ~(inputs[728]) | (inputs[921]);
    assign layer0_outputs[694] = (inputs[692]) & (inputs[832]);
    assign layer0_outputs[695] = (inputs[179]) & ~(inputs[87]);
    assign layer0_outputs[696] = inputs[707];
    assign layer0_outputs[697] = inputs[550];
    assign layer0_outputs[698] = ~(inputs[846]) | (inputs[972]);
    assign layer0_outputs[699] = ~(inputs[181]);
    assign layer0_outputs[700] = inputs[533];
    assign layer0_outputs[701] = (inputs[312]) ^ (inputs[451]);
    assign layer0_outputs[702] = ~(inputs[382]) | (inputs[1002]);
    assign layer0_outputs[703] = (inputs[573]) | (inputs[559]);
    assign layer0_outputs[704] = ~(inputs[527]);
    assign layer0_outputs[705] = ~((inputs[627]) ^ (inputs[487]));
    assign layer0_outputs[706] = (inputs[742]) ^ (inputs[56]);
    assign layer0_outputs[707] = ~((inputs[284]) | (inputs[73]));
    assign layer0_outputs[708] = inputs[323];
    assign layer0_outputs[709] = (inputs[517]) & ~(inputs[80]);
    assign layer0_outputs[710] = (inputs[935]) | (inputs[894]);
    assign layer0_outputs[711] = (inputs[796]) & (inputs[18]);
    assign layer0_outputs[712] = ~((inputs[783]) | (inputs[171]));
    assign layer0_outputs[713] = (inputs[303]) ^ (inputs[778]);
    assign layer0_outputs[714] = ~(inputs[557]) | (inputs[418]);
    assign layer0_outputs[715] = inputs[558];
    assign layer0_outputs[716] = ~(inputs[698]);
    assign layer0_outputs[717] = ~(inputs[460]);
    assign layer0_outputs[718] = (inputs[918]) | (inputs[289]);
    assign layer0_outputs[719] = ~((inputs[574]) ^ (inputs[332]));
    assign layer0_outputs[720] = ~((inputs[444]) | (inputs[547]));
    assign layer0_outputs[721] = ~(inputs[241]) | (inputs[85]);
    assign layer0_outputs[722] = inputs[474];
    assign layer0_outputs[723] = inputs[370];
    assign layer0_outputs[724] = ~((inputs[740]) ^ (inputs[610]));
    assign layer0_outputs[725] = ~((inputs[1002]) ^ (inputs[820]));
    assign layer0_outputs[726] = (inputs[318]) | (inputs[678]);
    assign layer0_outputs[727] = (inputs[593]) & ~(inputs[836]);
    assign layer0_outputs[728] = (inputs[528]) & ~(inputs[973]);
    assign layer0_outputs[729] = ~(inputs[814]) | (inputs[796]);
    assign layer0_outputs[730] = inputs[876];
    assign layer0_outputs[731] = ~(inputs[496]) | (inputs[351]);
    assign layer0_outputs[732] = ~(inputs[528]) | (inputs[462]);
    assign layer0_outputs[733] = (inputs[878]) | (inputs[298]);
    assign layer0_outputs[734] = ~((inputs[150]) | (inputs[933]));
    assign layer0_outputs[735] = ~(inputs[503]) | (inputs[16]);
    assign layer0_outputs[736] = (inputs[101]) ^ (inputs[303]);
    assign layer0_outputs[737] = ~(inputs[542]) | (inputs[385]);
    assign layer0_outputs[738] = inputs[879];
    assign layer0_outputs[739] = inputs[423];
    assign layer0_outputs[740] = ~((inputs[457]) ^ (inputs[588]));
    assign layer0_outputs[741] = ~(inputs[805]) | (inputs[961]);
    assign layer0_outputs[742] = (inputs[388]) | (inputs[468]);
    assign layer0_outputs[743] = ~((inputs[532]) | (inputs[352]));
    assign layer0_outputs[744] = (inputs[583]) & ~(inputs[1006]);
    assign layer0_outputs[745] = ~(inputs[389]);
    assign layer0_outputs[746] = (inputs[18]) & (inputs[576]);
    assign layer0_outputs[747] = ~(inputs[505]);
    assign layer0_outputs[748] = ~(inputs[497]);
    assign layer0_outputs[749] = ~(inputs[51]) | (inputs[16]);
    assign layer0_outputs[750] = inputs[946];
    assign layer0_outputs[751] = (inputs[96]) & ~(inputs[709]);
    assign layer0_outputs[752] = ~((inputs[876]) ^ (inputs[162]));
    assign layer0_outputs[753] = (inputs[597]) ^ (inputs[55]);
    assign layer0_outputs[754] = ~(inputs[540]) | (inputs[769]);
    assign layer0_outputs[755] = ~(inputs[148]);
    assign layer0_outputs[756] = ~(inputs[81]);
    assign layer0_outputs[757] = ~(inputs[615]);
    assign layer0_outputs[758] = inputs[496];
    assign layer0_outputs[759] = inputs[407];
    assign layer0_outputs[760] = (inputs[868]) & (inputs[986]);
    assign layer0_outputs[761] = ~((inputs[720]) | (inputs[325]));
    assign layer0_outputs[762] = ~(inputs[616]);
    assign layer0_outputs[763] = (inputs[992]) & (inputs[234]);
    assign layer0_outputs[764] = ~(inputs[968]);
    assign layer0_outputs[765] = inputs[344];
    assign layer0_outputs[766] = ~(inputs[597]);
    assign layer0_outputs[767] = ~((inputs[233]) | (inputs[717]));
    assign layer0_outputs[768] = inputs[246];
    assign layer0_outputs[769] = ~((inputs[746]) ^ (inputs[996]));
    assign layer0_outputs[770] = ~((inputs[634]) & (inputs[1021]));
    assign layer0_outputs[771] = inputs[712];
    assign layer0_outputs[772] = (inputs[19]) | (inputs[600]);
    assign layer0_outputs[773] = (inputs[35]) | (inputs[491]);
    assign layer0_outputs[774] = (inputs[980]) & ~(inputs[760]);
    assign layer0_outputs[775] = ~(inputs[295]);
    assign layer0_outputs[776] = inputs[325];
    assign layer0_outputs[777] = (inputs[491]) & ~(inputs[174]);
    assign layer0_outputs[778] = ~(inputs[725]) | (inputs[977]);
    assign layer0_outputs[779] = (inputs[43]) | (inputs[545]);
    assign layer0_outputs[780] = (inputs[376]) ^ (inputs[767]);
    assign layer0_outputs[781] = inputs[969];
    assign layer0_outputs[782] = (inputs[121]) ^ (inputs[360]);
    assign layer0_outputs[783] = (inputs[853]) & ~(inputs[973]);
    assign layer0_outputs[784] = (inputs[207]) & ~(inputs[103]);
    assign layer0_outputs[785] = ~(inputs[374]) | (inputs[647]);
    assign layer0_outputs[786] = (inputs[484]) & ~(inputs[864]);
    assign layer0_outputs[787] = ~(inputs[324]);
    assign layer0_outputs[788] = ~(inputs[995]);
    assign layer0_outputs[789] = ~(inputs[714]);
    assign layer0_outputs[790] = ~(inputs[175]) | (inputs[978]);
    assign layer0_outputs[791] = (inputs[782]) & ~(inputs[473]);
    assign layer0_outputs[792] = ~((inputs[34]) ^ (inputs[81]));
    assign layer0_outputs[793] = inputs[614];
    assign layer0_outputs[794] = (inputs[91]) | (inputs[686]);
    assign layer0_outputs[795] = (inputs[204]) ^ (inputs[666]);
    assign layer0_outputs[796] = ~((inputs[636]) ^ (inputs[85]));
    assign layer0_outputs[797] = (inputs[940]) & ~(inputs[160]);
    assign layer0_outputs[798] = ~(inputs[651]);
    assign layer0_outputs[799] = inputs[243];
    assign layer0_outputs[800] = ~(inputs[202]) | (inputs[823]);
    assign layer0_outputs[801] = ~(inputs[783]) | (inputs[768]);
    assign layer0_outputs[802] = (inputs[238]) | (inputs[418]);
    assign layer0_outputs[803] = inputs[150];
    assign layer0_outputs[804] = ~(inputs[588]) | (inputs[193]);
    assign layer0_outputs[805] = ~((inputs[853]) | (inputs[953]));
    assign layer0_outputs[806] = (inputs[581]) ^ (inputs[798]);
    assign layer0_outputs[807] = inputs[143];
    assign layer0_outputs[808] = ~(inputs[143]) | (inputs[609]);
    assign layer0_outputs[809] = (inputs[108]) | (inputs[491]);
    assign layer0_outputs[810] = ~(inputs[398]);
    assign layer0_outputs[811] = ~(inputs[669]);
    assign layer0_outputs[812] = (inputs[18]) & ~(inputs[379]);
    assign layer0_outputs[813] = (inputs[777]) & ~(inputs[474]);
    assign layer0_outputs[814] = (inputs[319]) & (inputs[191]);
    assign layer0_outputs[815] = (inputs[819]) ^ (inputs[59]);
    assign layer0_outputs[816] = 1'b1;
    assign layer0_outputs[817] = ~(inputs[434]);
    assign layer0_outputs[818] = ~(inputs[523]) | (inputs[987]);
    assign layer0_outputs[819] = ~(inputs[100]) | (inputs[231]);
    assign layer0_outputs[820] = ~(inputs[288]);
    assign layer0_outputs[821] = (inputs[78]) & ~(inputs[988]);
    assign layer0_outputs[822] = ~((inputs[839]) | (inputs[823]));
    assign layer0_outputs[823] = ~(inputs[364]);
    assign layer0_outputs[824] = inputs[713];
    assign layer0_outputs[825] = ~(inputs[86]);
    assign layer0_outputs[826] = ~(inputs[538]);
    assign layer0_outputs[827] = ~((inputs[877]) | (inputs[838]));
    assign layer0_outputs[828] = 1'b0;
    assign layer0_outputs[829] = (inputs[810]) | (inputs[0]);
    assign layer0_outputs[830] = ~((inputs[860]) & (inputs[574]));
    assign layer0_outputs[831] = ~((inputs[448]) | (inputs[234]));
    assign layer0_outputs[832] = ~(inputs[809]) | (inputs[976]);
    assign layer0_outputs[833] = ~(inputs[332]);
    assign layer0_outputs[834] = ~(inputs[591]);
    assign layer0_outputs[835] = ~(inputs[956]) | (inputs[44]);
    assign layer0_outputs[836] = ~(inputs[659]);
    assign layer0_outputs[837] = ~(inputs[369]) | (inputs[756]);
    assign layer0_outputs[838] = ~((inputs[836]) ^ (inputs[215]));
    assign layer0_outputs[839] = ~((inputs[821]) | (inputs[481]));
    assign layer0_outputs[840] = ~((inputs[371]) ^ (inputs[866]));
    assign layer0_outputs[841] = inputs[251];
    assign layer0_outputs[842] = ~(inputs[330]);
    assign layer0_outputs[843] = ~(inputs[349]);
    assign layer0_outputs[844] = (inputs[0]) & ~(inputs[183]);
    assign layer0_outputs[845] = (inputs[21]) & (inputs[308]);
    assign layer0_outputs[846] = (inputs[706]) & ~(inputs[1009]);
    assign layer0_outputs[847] = (inputs[363]) & ~(inputs[678]);
    assign layer0_outputs[848] = ~((inputs[220]) | (inputs[834]));
    assign layer0_outputs[849] = (inputs[359]) | (inputs[291]);
    assign layer0_outputs[850] = ~(inputs[786]) | (inputs[125]);
    assign layer0_outputs[851] = (inputs[871]) & (inputs[894]);
    assign layer0_outputs[852] = (inputs[342]) & ~(inputs[257]);
    assign layer0_outputs[853] = ~((inputs[235]) ^ (inputs[556]));
    assign layer0_outputs[854] = ~(inputs[33]);
    assign layer0_outputs[855] = inputs[942];
    assign layer0_outputs[856] = ~(inputs[294]);
    assign layer0_outputs[857] = inputs[100];
    assign layer0_outputs[858] = (inputs[879]) & ~(inputs[697]);
    assign layer0_outputs[859] = ~(inputs[566]) | (inputs[432]);
    assign layer0_outputs[860] = (inputs[356]) & ~(inputs[856]);
    assign layer0_outputs[861] = (inputs[939]) & ~(inputs[614]);
    assign layer0_outputs[862] = ~(inputs[518]) | (inputs[482]);
    assign layer0_outputs[863] = ~(inputs[304]) | (inputs[93]);
    assign layer0_outputs[864] = (inputs[974]) | (inputs[355]);
    assign layer0_outputs[865] = (inputs[585]) | (inputs[405]);
    assign layer0_outputs[866] = inputs[369];
    assign layer0_outputs[867] = ~(inputs[303]);
    assign layer0_outputs[868] = ~((inputs[740]) ^ (inputs[544]));
    assign layer0_outputs[869] = inputs[462];
    assign layer0_outputs[870] = ~(inputs[178]) | (inputs[63]);
    assign layer0_outputs[871] = ~(inputs[895]) | (inputs[1013]);
    assign layer0_outputs[872] = inputs[586];
    assign layer0_outputs[873] = ~((inputs[917]) | (inputs[393]));
    assign layer0_outputs[874] = (inputs[451]) ^ (inputs[3]);
    assign layer0_outputs[875] = ~((inputs[869]) | (inputs[659]));
    assign layer0_outputs[876] = ~((inputs[37]) ^ (inputs[67]));
    assign layer0_outputs[877] = ~(inputs[519]) | (inputs[10]);
    assign layer0_outputs[878] = (inputs[328]) ^ (inputs[830]);
    assign layer0_outputs[879] = ~((inputs[746]) | (inputs[640]));
    assign layer0_outputs[880] = inputs[282];
    assign layer0_outputs[881] = (inputs[895]) | (inputs[581]);
    assign layer0_outputs[882] = ~((inputs[1000]) & (inputs[998]));
    assign layer0_outputs[883] = ~(inputs[496]) | (inputs[1017]);
    assign layer0_outputs[884] = (inputs[543]) | (inputs[622]);
    assign layer0_outputs[885] = ~((inputs[893]) | (inputs[733]));
    assign layer0_outputs[886] = (inputs[765]) | (inputs[650]);
    assign layer0_outputs[887] = inputs[507];
    assign layer0_outputs[888] = (inputs[242]) | (inputs[803]);
    assign layer0_outputs[889] = inputs[564];
    assign layer0_outputs[890] = (inputs[515]) ^ (inputs[659]);
    assign layer0_outputs[891] = ~((inputs[137]) | (inputs[144]));
    assign layer0_outputs[892] = ~((inputs[760]) ^ (inputs[809]));
    assign layer0_outputs[893] = ~(inputs[992]);
    assign layer0_outputs[894] = (inputs[453]) | (inputs[942]);
    assign layer0_outputs[895] = (inputs[303]) & (inputs[219]);
    assign layer0_outputs[896] = (inputs[760]) ^ (inputs[213]);
    assign layer0_outputs[897] = ~((inputs[198]) & (inputs[57]));
    assign layer0_outputs[898] = inputs[848];
    assign layer0_outputs[899] = ~((inputs[564]) | (inputs[312]));
    assign layer0_outputs[900] = ~((inputs[718]) | (inputs[743]));
    assign layer0_outputs[901] = (inputs[110]) & (inputs[35]);
    assign layer0_outputs[902] = ~((inputs[52]) ^ (inputs[252]));
    assign layer0_outputs[903] = ~((inputs[710]) | (inputs[912]));
    assign layer0_outputs[904] = ~(inputs[391]) | (inputs[671]);
    assign layer0_outputs[905] = ~((inputs[695]) & (inputs[395]));
    assign layer0_outputs[906] = ~((inputs[678]) & (inputs[971]));
    assign layer0_outputs[907] = ~(inputs[519]) | (inputs[815]);
    assign layer0_outputs[908] = ~((inputs[781]) | (inputs[7]));
    assign layer0_outputs[909] = ~(inputs[233]);
    assign layer0_outputs[910] = ~(inputs[375]);
    assign layer0_outputs[911] = (inputs[785]) & ~(inputs[827]);
    assign layer0_outputs[912] = inputs[280];
    assign layer0_outputs[913] = ~(inputs[680]);
    assign layer0_outputs[914] = ~((inputs[278]) | (inputs[360]));
    assign layer0_outputs[915] = ~(inputs[471]) | (inputs[605]);
    assign layer0_outputs[916] = (inputs[411]) & ~(inputs[112]);
    assign layer0_outputs[917] = 1'b0;
    assign layer0_outputs[918] = ~(inputs[915]) | (inputs[899]);
    assign layer0_outputs[919] = (inputs[541]) & ~(inputs[308]);
    assign layer0_outputs[920] = ~(inputs[338]);
    assign layer0_outputs[921] = ~(inputs[712]);
    assign layer0_outputs[922] = 1'b1;
    assign layer0_outputs[923] = (inputs[437]) & ~(inputs[538]);
    assign layer0_outputs[924] = ~((inputs[835]) ^ (inputs[378]));
    assign layer0_outputs[925] = ~(inputs[740]);
    assign layer0_outputs[926] = (inputs[1000]) | (inputs[6]);
    assign layer0_outputs[927] = (inputs[272]) & ~(inputs[610]);
    assign layer0_outputs[928] = (inputs[78]) & ~(inputs[228]);
    assign layer0_outputs[929] = ~(inputs[412]);
    assign layer0_outputs[930] = inputs[225];
    assign layer0_outputs[931] = ~(inputs[884]);
    assign layer0_outputs[932] = ~(inputs[561]);
    assign layer0_outputs[933] = inputs[839];
    assign layer0_outputs[934] = inputs[909];
    assign layer0_outputs[935] = ~(inputs[77]);
    assign layer0_outputs[936] = ~(inputs[401]);
    assign layer0_outputs[937] = inputs[245];
    assign layer0_outputs[938] = inputs[513];
    assign layer0_outputs[939] = inputs[907];
    assign layer0_outputs[940] = (inputs[654]) ^ (inputs[195]);
    assign layer0_outputs[941] = ~(inputs[927]) | (inputs[341]);
    assign layer0_outputs[942] = ~(inputs[103]) | (inputs[166]);
    assign layer0_outputs[943] = ~(inputs[531]);
    assign layer0_outputs[944] = (inputs[979]) | (inputs[532]);
    assign layer0_outputs[945] = ~((inputs[666]) | (inputs[797]));
    assign layer0_outputs[946] = ~((inputs[415]) ^ (inputs[968]));
    assign layer0_outputs[947] = ~(inputs[683]);
    assign layer0_outputs[948] = (inputs[501]) | (inputs[510]);
    assign layer0_outputs[949] = ~(inputs[533]) | (inputs[617]);
    assign layer0_outputs[950] = ~(inputs[313]);
    assign layer0_outputs[951] = ~((inputs[347]) ^ (inputs[134]));
    assign layer0_outputs[952] = ~((inputs[663]) | (inputs[994]));
    assign layer0_outputs[953] = (inputs[320]) & (inputs[263]);
    assign layer0_outputs[954] = 1'b0;
    assign layer0_outputs[955] = ~(inputs[687]) | (inputs[34]);
    assign layer0_outputs[956] = inputs[713];
    assign layer0_outputs[957] = (inputs[27]) ^ (inputs[749]);
    assign layer0_outputs[958] = (inputs[935]) ^ (inputs[398]);
    assign layer0_outputs[959] = (inputs[898]) ^ (inputs[842]);
    assign layer0_outputs[960] = ~(inputs[688]) | (inputs[443]);
    assign layer0_outputs[961] = (inputs[277]) & ~(inputs[185]);
    assign layer0_outputs[962] = ~(inputs[15]) | (inputs[1005]);
    assign layer0_outputs[963] = (inputs[209]) ^ (inputs[984]);
    assign layer0_outputs[964] = inputs[687];
    assign layer0_outputs[965] = ~(inputs[898]);
    assign layer0_outputs[966] = (inputs[311]) | (inputs[569]);
    assign layer0_outputs[967] = ~(inputs[702]);
    assign layer0_outputs[968] = inputs[846];
    assign layer0_outputs[969] = ~((inputs[352]) ^ (inputs[165]));
    assign layer0_outputs[970] = (inputs[343]) | (inputs[8]);
    assign layer0_outputs[971] = (inputs[775]) ^ (inputs[387]);
    assign layer0_outputs[972] = ~((inputs[643]) ^ (inputs[914]));
    assign layer0_outputs[973] = (inputs[786]) | (inputs[905]);
    assign layer0_outputs[974] = ~((inputs[36]) ^ (inputs[460]));
    assign layer0_outputs[975] = ~((inputs[188]) ^ (inputs[593]));
    assign layer0_outputs[976] = ~(inputs[126]);
    assign layer0_outputs[977] = ~(inputs[392]) | (inputs[886]);
    assign layer0_outputs[978] = 1'b1;
    assign layer0_outputs[979] = ~(inputs[158]);
    assign layer0_outputs[980] = ~((inputs[183]) ^ (inputs[546]));
    assign layer0_outputs[981] = (inputs[95]) & ~(inputs[611]);
    assign layer0_outputs[982] = ~((inputs[768]) | (inputs[307]));
    assign layer0_outputs[983] = (inputs[182]) ^ (inputs[836]);
    assign layer0_outputs[984] = ~((inputs[469]) | (inputs[45]));
    assign layer0_outputs[985] = (inputs[419]) & ~(inputs[965]);
    assign layer0_outputs[986] = ~((inputs[389]) ^ (inputs[878]));
    assign layer0_outputs[987] = ~((inputs[813]) | (inputs[594]));
    assign layer0_outputs[988] = 1'b1;
    assign layer0_outputs[989] = (inputs[185]) ^ (inputs[652]);
    assign layer0_outputs[990] = ~(inputs[850]);
    assign layer0_outputs[991] = ~((inputs[985]) & (inputs[259]));
    assign layer0_outputs[992] = ~(inputs[620]);
    assign layer0_outputs[993] = ~((inputs[56]) ^ (inputs[570]));
    assign layer0_outputs[994] = inputs[717];
    assign layer0_outputs[995] = ~(inputs[810]);
    assign layer0_outputs[996] = ~((inputs[610]) | (inputs[189]));
    assign layer0_outputs[997] = inputs[841];
    assign layer0_outputs[998] = (inputs[1001]) ^ (inputs[958]);
    assign layer0_outputs[999] = 1'b1;
    assign layer0_outputs[1000] = (inputs[555]) | (inputs[925]);
    assign layer0_outputs[1001] = ~(inputs[678]);
    assign layer0_outputs[1002] = ~((inputs[31]) & (inputs[416]));
    assign layer0_outputs[1003] = (inputs[510]) & ~(inputs[480]);
    assign layer0_outputs[1004] = ~(inputs[350]);
    assign layer0_outputs[1005] = ~((inputs[960]) | (inputs[951]));
    assign layer0_outputs[1006] = (inputs[457]) & (inputs[649]);
    assign layer0_outputs[1007] = ~((inputs[808]) | (inputs[910]));
    assign layer0_outputs[1008] = (inputs[1001]) ^ (inputs[748]);
    assign layer0_outputs[1009] = ~(inputs[381]) | (inputs[1013]);
    assign layer0_outputs[1010] = ~((inputs[320]) & (inputs[75]));
    assign layer0_outputs[1011] = ~(inputs[73]) | (inputs[116]);
    assign layer0_outputs[1012] = (inputs[670]) & ~(inputs[544]);
    assign layer0_outputs[1013] = (inputs[649]) & ~(inputs[224]);
    assign layer0_outputs[1014] = (inputs[527]) ^ (inputs[994]);
    assign layer0_outputs[1015] = (inputs[28]) | (inputs[116]);
    assign layer0_outputs[1016] = ~(inputs[302]);
    assign layer0_outputs[1017] = ~(inputs[605]) | (inputs[104]);
    assign layer0_outputs[1018] = (inputs[996]) & (inputs[448]);
    assign layer0_outputs[1019] = inputs[720];
    assign layer0_outputs[1020] = (inputs[530]) | (inputs[151]);
    assign layer0_outputs[1021] = ~((inputs[812]) | (inputs[666]));
    assign layer0_outputs[1022] = (inputs[189]) ^ (inputs[629]);
    assign layer0_outputs[1023] = (inputs[275]) & ~(inputs[573]);
    assign layer0_outputs[1024] = ~(inputs[85]);
    assign layer0_outputs[1025] = inputs[745];
    assign layer0_outputs[1026] = ~(inputs[39]);
    assign layer0_outputs[1027] = ~(inputs[130]);
    assign layer0_outputs[1028] = (inputs[472]) | (inputs[517]);
    assign layer0_outputs[1029] = ~((inputs[854]) ^ (inputs[844]));
    assign layer0_outputs[1030] = 1'b1;
    assign layer0_outputs[1031] = ~((inputs[23]) ^ (inputs[508]));
    assign layer0_outputs[1032] = (inputs[734]) | (inputs[371]);
    assign layer0_outputs[1033] = (inputs[510]) ^ (inputs[348]);
    assign layer0_outputs[1034] = (inputs[856]) | (inputs[859]);
    assign layer0_outputs[1035] = ~((inputs[847]) | (inputs[467]));
    assign layer0_outputs[1036] = (inputs[776]) | (inputs[323]);
    assign layer0_outputs[1037] = ~((inputs[252]) & (inputs[858]));
    assign layer0_outputs[1038] = (inputs[527]) & ~(inputs[288]);
    assign layer0_outputs[1039] = ~(inputs[492]);
    assign layer0_outputs[1040] = (inputs[747]) | (inputs[327]);
    assign layer0_outputs[1041] = (inputs[584]) ^ (inputs[143]);
    assign layer0_outputs[1042] = 1'b0;
    assign layer0_outputs[1043] = ~(inputs[202]) | (inputs[157]);
    assign layer0_outputs[1044] = (inputs[760]) | (inputs[68]);
    assign layer0_outputs[1045] = ~((inputs[642]) ^ (inputs[822]));
    assign layer0_outputs[1046] = (inputs[935]) ^ (inputs[461]);
    assign layer0_outputs[1047] = (inputs[1012]) & (inputs[972]);
    assign layer0_outputs[1048] = ~((inputs[627]) ^ (inputs[591]));
    assign layer0_outputs[1049] = (inputs[59]) | (inputs[234]);
    assign layer0_outputs[1050] = (inputs[183]) & (inputs[342]);
    assign layer0_outputs[1051] = (inputs[880]) & ~(inputs[79]);
    assign layer0_outputs[1052] = ~(inputs[4]);
    assign layer0_outputs[1053] = ~(inputs[408]);
    assign layer0_outputs[1054] = (inputs[514]) | (inputs[835]);
    assign layer0_outputs[1055] = inputs[968];
    assign layer0_outputs[1056] = (inputs[198]) & (inputs[90]);
    assign layer0_outputs[1057] = ~(inputs[140]);
    assign layer0_outputs[1058] = inputs[314];
    assign layer0_outputs[1059] = ~(inputs[495]);
    assign layer0_outputs[1060] = ~(inputs[660]) | (inputs[489]);
    assign layer0_outputs[1061] = (inputs[538]) ^ (inputs[322]);
    assign layer0_outputs[1062] = inputs[748];
    assign layer0_outputs[1063] = ~((inputs[911]) ^ (inputs[915]));
    assign layer0_outputs[1064] = ~((inputs[345]) | (inputs[446]));
    assign layer0_outputs[1065] = inputs[429];
    assign layer0_outputs[1066] = (inputs[307]) & ~(inputs[48]);
    assign layer0_outputs[1067] = ~(inputs[312]) | (inputs[108]);
    assign layer0_outputs[1068] = ~(inputs[859]);
    assign layer0_outputs[1069] = (inputs[404]) & ~(inputs[234]);
    assign layer0_outputs[1070] = ~((inputs[458]) | (inputs[289]));
    assign layer0_outputs[1071] = (inputs[434]) & ~(inputs[361]);
    assign layer0_outputs[1072] = (inputs[905]) | (inputs[759]);
    assign layer0_outputs[1073] = 1'b1;
    assign layer0_outputs[1074] = ~((inputs[216]) | (inputs[258]));
    assign layer0_outputs[1075] = inputs[311];
    assign layer0_outputs[1076] = ~(inputs[470]) | (inputs[993]);
    assign layer0_outputs[1077] = (inputs[27]) & ~(inputs[108]);
    assign layer0_outputs[1078] = (inputs[15]) & ~(inputs[356]);
    assign layer0_outputs[1079] = inputs[423];
    assign layer0_outputs[1080] = ~(inputs[348]) | (inputs[17]);
    assign layer0_outputs[1081] = ~(inputs[325]) | (inputs[13]);
    assign layer0_outputs[1082] = ~((inputs[459]) | (inputs[592]));
    assign layer0_outputs[1083] = ~((inputs[558]) | (inputs[130]));
    assign layer0_outputs[1084] = ~((inputs[468]) & (inputs[609]));
    assign layer0_outputs[1085] = inputs[214];
    assign layer0_outputs[1086] = ~(inputs[268]) | (inputs[980]);
    assign layer0_outputs[1087] = ~((inputs[988]) & (inputs[59]));
    assign layer0_outputs[1088] = 1'b0;
    assign layer0_outputs[1089] = (inputs[17]) | (inputs[508]);
    assign layer0_outputs[1090] = (inputs[267]) & ~(inputs[606]);
    assign layer0_outputs[1091] = inputs[436];
    assign layer0_outputs[1092] = (inputs[412]) & ~(inputs[929]);
    assign layer0_outputs[1093] = ~((inputs[475]) | (inputs[562]));
    assign layer0_outputs[1094] = ~((inputs[517]) | (inputs[271]));
    assign layer0_outputs[1095] = ~((inputs[774]) | (inputs[276]));
    assign layer0_outputs[1096] = inputs[247];
    assign layer0_outputs[1097] = inputs[216];
    assign layer0_outputs[1098] = ~(inputs[399]) | (inputs[553]);
    assign layer0_outputs[1099] = ~(inputs[70]) | (inputs[442]);
    assign layer0_outputs[1100] = (inputs[185]) | (inputs[636]);
    assign layer0_outputs[1101] = ~((inputs[142]) ^ (inputs[159]));
    assign layer0_outputs[1102] = (inputs[392]) & ~(inputs[413]);
    assign layer0_outputs[1103] = (inputs[46]) ^ (inputs[884]);
    assign layer0_outputs[1104] = ~((inputs[685]) | (inputs[418]));
    assign layer0_outputs[1105] = ~((inputs[10]) | (inputs[357]));
    assign layer0_outputs[1106] = ~((inputs[356]) ^ (inputs[580]));
    assign layer0_outputs[1107] = ~(inputs[531]);
    assign layer0_outputs[1108] = ~(inputs[318]);
    assign layer0_outputs[1109] = (inputs[977]) | (inputs[547]);
    assign layer0_outputs[1110] = ~(inputs[687]) | (inputs[414]);
    assign layer0_outputs[1111] = ~(inputs[561]) | (inputs[17]);
    assign layer0_outputs[1112] = (inputs[827]) & ~(inputs[609]);
    assign layer0_outputs[1113] = (inputs[684]) | (inputs[158]);
    assign layer0_outputs[1114] = ~((inputs[427]) | (inputs[646]));
    assign layer0_outputs[1115] = inputs[342];
    assign layer0_outputs[1116] = (inputs[186]) & (inputs[954]);
    assign layer0_outputs[1117] = (inputs[595]) | (inputs[132]);
    assign layer0_outputs[1118] = (inputs[885]) | (inputs[168]);
    assign layer0_outputs[1119] = ~(inputs[53]) | (inputs[624]);
    assign layer0_outputs[1120] = (inputs[262]) | (inputs[693]);
    assign layer0_outputs[1121] = ~((inputs[653]) ^ (inputs[241]));
    assign layer0_outputs[1122] = (inputs[617]) & ~(inputs[384]);
    assign layer0_outputs[1123] = ~((inputs[725]) | (inputs[497]));
    assign layer0_outputs[1124] = ~(inputs[392]) | (inputs[928]);
    assign layer0_outputs[1125] = ~(inputs[301]) | (inputs[689]);
    assign layer0_outputs[1126] = (inputs[426]) & ~(inputs[637]);
    assign layer0_outputs[1127] = ~(inputs[307]);
    assign layer0_outputs[1128] = ~(inputs[519]);
    assign layer0_outputs[1129] = ~(inputs[52]);
    assign layer0_outputs[1130] = (inputs[658]) ^ (inputs[802]);
    assign layer0_outputs[1131] = inputs[341];
    assign layer0_outputs[1132] = ~(inputs[415]) | (inputs[59]);
    assign layer0_outputs[1133] = ~((inputs[27]) | (inputs[606]));
    assign layer0_outputs[1134] = ~((inputs[469]) ^ (inputs[863]));
    assign layer0_outputs[1135] = ~(inputs[580]);
    assign layer0_outputs[1136] = (inputs[844]) ^ (inputs[155]);
    assign layer0_outputs[1137] = inputs[967];
    assign layer0_outputs[1138] = (inputs[88]) & (inputs[52]);
    assign layer0_outputs[1139] = ~(inputs[347]);
    assign layer0_outputs[1140] = ~(inputs[1003]);
    assign layer0_outputs[1141] = 1'b1;
    assign layer0_outputs[1142] = ~((inputs[338]) | (inputs[453]));
    assign layer0_outputs[1143] = (inputs[133]) ^ (inputs[698]);
    assign layer0_outputs[1144] = (inputs[210]) & ~(inputs[904]);
    assign layer0_outputs[1145] = ~((inputs[875]) | (inputs[245]));
    assign layer0_outputs[1146] = (inputs[556]) ^ (inputs[150]);
    assign layer0_outputs[1147] = ~(inputs[445]);
    assign layer0_outputs[1148] = ~(inputs[705]) | (inputs[958]);
    assign layer0_outputs[1149] = inputs[278];
    assign layer0_outputs[1150] = (inputs[367]) & ~(inputs[312]);
    assign layer0_outputs[1151] = ~((inputs[253]) & (inputs[632]));
    assign layer0_outputs[1152] = ~((inputs[630]) | (inputs[808]));
    assign layer0_outputs[1153] = ~((inputs[683]) ^ (inputs[479]));
    assign layer0_outputs[1154] = ~((inputs[62]) | (inputs[973]));
    assign layer0_outputs[1155] = ~((inputs[874]) ^ (inputs[128]));
    assign layer0_outputs[1156] = (inputs[393]) & ~(inputs[280]);
    assign layer0_outputs[1157] = ~(inputs[282]) | (inputs[53]);
    assign layer0_outputs[1158] = ~(inputs[1017]);
    assign layer0_outputs[1159] = ~(inputs[31]);
    assign layer0_outputs[1160] = (inputs[5]) & ~(inputs[351]);
    assign layer0_outputs[1161] = ~((inputs[465]) | (inputs[949]));
    assign layer0_outputs[1162] = ~(inputs[592]);
    assign layer0_outputs[1163] = (inputs[809]) | (inputs[645]);
    assign layer0_outputs[1164] = ~(inputs[529]);
    assign layer0_outputs[1165] = (inputs[627]) | (inputs[734]);
    assign layer0_outputs[1166] = inputs[850];
    assign layer0_outputs[1167] = ~(inputs[774]) | (inputs[647]);
    assign layer0_outputs[1168] = ~((inputs[284]) ^ (inputs[204]));
    assign layer0_outputs[1169] = ~(inputs[110]);
    assign layer0_outputs[1170] = ~(inputs[724]);
    assign layer0_outputs[1171] = (inputs[437]) | (inputs[880]);
    assign layer0_outputs[1172] = ~(inputs[611]) | (inputs[608]);
    assign layer0_outputs[1173] = ~(inputs[778]);
    assign layer0_outputs[1174] = ~((inputs[660]) ^ (inputs[610]));
    assign layer0_outputs[1175] = 1'b0;
    assign layer0_outputs[1176] = ~(inputs[286]) | (inputs[197]);
    assign layer0_outputs[1177] = (inputs[782]) | (inputs[806]);
    assign layer0_outputs[1178] = ~(inputs[544]) | (inputs[485]);
    assign layer0_outputs[1179] = ~((inputs[647]) | (inputs[722]));
    assign layer0_outputs[1180] = ~((inputs[460]) | (inputs[315]));
    assign layer0_outputs[1181] = (inputs[332]) ^ (inputs[218]);
    assign layer0_outputs[1182] = ~(inputs[501]);
    assign layer0_outputs[1183] = inputs[492];
    assign layer0_outputs[1184] = ~(inputs[498]);
    assign layer0_outputs[1185] = 1'b0;
    assign layer0_outputs[1186] = 1'b1;
    assign layer0_outputs[1187] = ~((inputs[11]) ^ (inputs[146]));
    assign layer0_outputs[1188] = ~(inputs[38]) | (inputs[829]);
    assign layer0_outputs[1189] = ~(inputs[654]) | (inputs[1006]);
    assign layer0_outputs[1190] = ~((inputs[728]) | (inputs[169]));
    assign layer0_outputs[1191] = (inputs[368]) | (inputs[96]);
    assign layer0_outputs[1192] = inputs[343];
    assign layer0_outputs[1193] = (inputs[934]) & ~(inputs[827]);
    assign layer0_outputs[1194] = (inputs[199]) ^ (inputs[120]);
    assign layer0_outputs[1195] = ~((inputs[659]) | (inputs[899]));
    assign layer0_outputs[1196] = (inputs[107]) | (inputs[917]);
    assign layer0_outputs[1197] = ~((inputs[886]) | (inputs[10]));
    assign layer0_outputs[1198] = (inputs[269]) & ~(inputs[877]);
    assign layer0_outputs[1199] = (inputs[708]) | (inputs[730]);
    assign layer0_outputs[1200] = 1'b0;
    assign layer0_outputs[1201] = ~((inputs[822]) ^ (inputs[831]));
    assign layer0_outputs[1202] = ~((inputs[610]) ^ (inputs[919]));
    assign layer0_outputs[1203] = (inputs[728]) & ~(inputs[983]);
    assign layer0_outputs[1204] = 1'b1;
    assign layer0_outputs[1205] = (inputs[801]) ^ (inputs[814]);
    assign layer0_outputs[1206] = ~((inputs[403]) | (inputs[229]));
    assign layer0_outputs[1207] = ~(inputs[765]) | (inputs[634]);
    assign layer0_outputs[1208] = inputs[528];
    assign layer0_outputs[1209] = ~((inputs[126]) | (inputs[514]));
    assign layer0_outputs[1210] = (inputs[873]) & ~(inputs[677]);
    assign layer0_outputs[1211] = (inputs[418]) | (inputs[934]);
    assign layer0_outputs[1212] = ~((inputs[426]) | (inputs[447]));
    assign layer0_outputs[1213] = ~(inputs[527]) | (inputs[575]);
    assign layer0_outputs[1214] = (inputs[16]) | (inputs[887]);
    assign layer0_outputs[1215] = ~(inputs[59]) | (inputs[195]);
    assign layer0_outputs[1216] = 1'b1;
    assign layer0_outputs[1217] = ~((inputs[542]) | (inputs[506]));
    assign layer0_outputs[1218] = ~((inputs[640]) & (inputs[540]));
    assign layer0_outputs[1219] = (inputs[817]) & ~(inputs[7]);
    assign layer0_outputs[1220] = ~(inputs[454]) | (inputs[219]);
    assign layer0_outputs[1221] = ~(inputs[600]) | (inputs[832]);
    assign layer0_outputs[1222] = inputs[717];
    assign layer0_outputs[1223] = (inputs[878]) ^ (inputs[1016]);
    assign layer0_outputs[1224] = inputs[365];
    assign layer0_outputs[1225] = inputs[553];
    assign layer0_outputs[1226] = ~(inputs[504]) | (inputs[969]);
    assign layer0_outputs[1227] = (inputs[494]) & ~(inputs[146]);
    assign layer0_outputs[1228] = ~((inputs[948]) | (inputs[296]));
    assign layer0_outputs[1229] = (inputs[965]) | (inputs[633]);
    assign layer0_outputs[1230] = ~(inputs[220]) | (inputs[316]);
    assign layer0_outputs[1231] = (inputs[1022]) ^ (inputs[456]);
    assign layer0_outputs[1232] = (inputs[317]) | (inputs[385]);
    assign layer0_outputs[1233] = ~((inputs[643]) ^ (inputs[798]));
    assign layer0_outputs[1234] = 1'b0;
    assign layer0_outputs[1235] = ~(inputs[681]);
    assign layer0_outputs[1236] = 1'b0;
    assign layer0_outputs[1237] = 1'b0;
    assign layer0_outputs[1238] = inputs[780];
    assign layer0_outputs[1239] = inputs[811];
    assign layer0_outputs[1240] = inputs[594];
    assign layer0_outputs[1241] = (inputs[877]) & ~(inputs[573]);
    assign layer0_outputs[1242] = ~(inputs[568]) | (inputs[860]);
    assign layer0_outputs[1243] = (inputs[232]) ^ (inputs[644]);
    assign layer0_outputs[1244] = (inputs[593]) & ~(inputs[185]);
    assign layer0_outputs[1245] = ~((inputs[0]) ^ (inputs[449]));
    assign layer0_outputs[1246] = inputs[164];
    assign layer0_outputs[1247] = ~(inputs[712]) | (inputs[152]);
    assign layer0_outputs[1248] = inputs[176];
    assign layer0_outputs[1249] = ~((inputs[440]) | (inputs[300]));
    assign layer0_outputs[1250] = inputs[776];
    assign layer0_outputs[1251] = ~(inputs[122]);
    assign layer0_outputs[1252] = inputs[69];
    assign layer0_outputs[1253] = ~(inputs[638]) | (inputs[616]);
    assign layer0_outputs[1254] = ~((inputs[119]) ^ (inputs[998]));
    assign layer0_outputs[1255] = inputs[521];
    assign layer0_outputs[1256] = ~(inputs[605]) | (inputs[138]);
    assign layer0_outputs[1257] = inputs[899];
    assign layer0_outputs[1258] = ~(inputs[47]) | (inputs[504]);
    assign layer0_outputs[1259] = (inputs[964]) & ~(inputs[162]);
    assign layer0_outputs[1260] = ~((inputs[813]) | (inputs[993]));
    assign layer0_outputs[1261] = (inputs[666]) & ~(inputs[44]);
    assign layer0_outputs[1262] = ~((inputs[578]) & (inputs[72]));
    assign layer0_outputs[1263] = inputs[141];
    assign layer0_outputs[1264] = ~((inputs[841]) | (inputs[664]));
    assign layer0_outputs[1265] = inputs[346];
    assign layer0_outputs[1266] = inputs[430];
    assign layer0_outputs[1267] = ~(inputs[636]);
    assign layer0_outputs[1268] = ~((inputs[699]) ^ (inputs[777]));
    assign layer0_outputs[1269] = ~(inputs[393]);
    assign layer0_outputs[1270] = inputs[913];
    assign layer0_outputs[1271] = (inputs[370]) ^ (inputs[257]);
    assign layer0_outputs[1272] = inputs[927];
    assign layer0_outputs[1273] = ~(inputs[631]) | (inputs[543]);
    assign layer0_outputs[1274] = ~(inputs[366]) | (inputs[477]);
    assign layer0_outputs[1275] = 1'b0;
    assign layer0_outputs[1276] = (inputs[594]) & ~(inputs[678]);
    assign layer0_outputs[1277] = ~(inputs[829]);
    assign layer0_outputs[1278] = (inputs[69]) ^ (inputs[894]);
    assign layer0_outputs[1279] = (inputs[807]) | (inputs[413]);
    assign layer0_outputs[1280] = ~(inputs[878]);
    assign layer0_outputs[1281] = (inputs[911]) ^ (inputs[774]);
    assign layer0_outputs[1282] = (inputs[429]) | (inputs[186]);
    assign layer0_outputs[1283] = ~(inputs[367]);
    assign layer0_outputs[1284] = (inputs[115]) ^ (inputs[357]);
    assign layer0_outputs[1285] = ~((inputs[513]) ^ (inputs[581]));
    assign layer0_outputs[1286] = ~(inputs[812]);
    assign layer0_outputs[1287] = 1'b1;
    assign layer0_outputs[1288] = ~(inputs[919]) | (inputs[252]);
    assign layer0_outputs[1289] = ~(inputs[51]);
    assign layer0_outputs[1290] = ~((inputs[916]) ^ (inputs[586]));
    assign layer0_outputs[1291] = (inputs[101]) | (inputs[422]);
    assign layer0_outputs[1292] = ~((inputs[443]) ^ (inputs[619]));
    assign layer0_outputs[1293] = inputs[707];
    assign layer0_outputs[1294] = inputs[712];
    assign layer0_outputs[1295] = ~(inputs[23]) | (inputs[971]);
    assign layer0_outputs[1296] = inputs[312];
    assign layer0_outputs[1297] = ~((inputs[147]) | (inputs[222]));
    assign layer0_outputs[1298] = ~(inputs[185]);
    assign layer0_outputs[1299] = ~(inputs[775]) | (inputs[946]);
    assign layer0_outputs[1300] = (inputs[662]) | (inputs[660]);
    assign layer0_outputs[1301] = inputs[752];
    assign layer0_outputs[1302] = (inputs[616]) | (inputs[266]);
    assign layer0_outputs[1303] = ~((inputs[283]) | (inputs[569]));
    assign layer0_outputs[1304] = (inputs[268]) & ~(inputs[218]);
    assign layer0_outputs[1305] = (inputs[529]) | (inputs[284]);
    assign layer0_outputs[1306] = (inputs[196]) | (inputs[632]);
    assign layer0_outputs[1307] = inputs[6];
    assign layer0_outputs[1308] = inputs[516];
    assign layer0_outputs[1309] = ~(inputs[1004]) | (inputs[524]);
    assign layer0_outputs[1310] = (inputs[395]) & ~(inputs[774]);
    assign layer0_outputs[1311] = (inputs[627]) & ~(inputs[951]);
    assign layer0_outputs[1312] = ~(inputs[238]);
    assign layer0_outputs[1313] = inputs[228];
    assign layer0_outputs[1314] = ~(inputs[739]) | (inputs[859]);
    assign layer0_outputs[1315] = ~(inputs[586]) | (inputs[105]);
    assign layer0_outputs[1316] = (inputs[448]) | (inputs[433]);
    assign layer0_outputs[1317] = 1'b1;
    assign layer0_outputs[1318] = (inputs[749]) | (inputs[126]);
    assign layer0_outputs[1319] = 1'b0;
    assign layer0_outputs[1320] = (inputs[533]) & ~(inputs[250]);
    assign layer0_outputs[1321] = ~(inputs[220]) | (inputs[770]);
    assign layer0_outputs[1322] = (inputs[420]) | (inputs[626]);
    assign layer0_outputs[1323] = (inputs[77]) | (inputs[914]);
    assign layer0_outputs[1324] = (inputs[342]) | (inputs[500]);
    assign layer0_outputs[1325] = ~(inputs[363]);
    assign layer0_outputs[1326] = ~(inputs[177]) | (inputs[960]);
    assign layer0_outputs[1327] = ~((inputs[731]) | (inputs[675]));
    assign layer0_outputs[1328] = inputs[765];
    assign layer0_outputs[1329] = ~((inputs[703]) ^ (inputs[764]));
    assign layer0_outputs[1330] = inputs[174];
    assign layer0_outputs[1331] = (inputs[760]) ^ (inputs[991]);
    assign layer0_outputs[1332] = (inputs[966]) ^ (inputs[483]);
    assign layer0_outputs[1333] = inputs[332];
    assign layer0_outputs[1334] = ~((inputs[306]) | (inputs[709]));
    assign layer0_outputs[1335] = inputs[631];
    assign layer0_outputs[1336] = (inputs[946]) | (inputs[13]);
    assign layer0_outputs[1337] = (inputs[897]) ^ (inputs[50]);
    assign layer0_outputs[1338] = ~((inputs[194]) & (inputs[155]));
    assign layer0_outputs[1339] = (inputs[587]) ^ (inputs[591]);
    assign layer0_outputs[1340] = inputs[582];
    assign layer0_outputs[1341] = inputs[102];
    assign layer0_outputs[1342] = ~(inputs[680]);
    assign layer0_outputs[1343] = ~((inputs[325]) | (inputs[985]));
    assign layer0_outputs[1344] = ~((inputs[244]) | (inputs[995]));
    assign layer0_outputs[1345] = ~(inputs[415]);
    assign layer0_outputs[1346] = inputs[208];
    assign layer0_outputs[1347] = (inputs[189]) | (inputs[837]);
    assign layer0_outputs[1348] = ~(inputs[662]);
    assign layer0_outputs[1349] = ~((inputs[15]) | (inputs[344]));
    assign layer0_outputs[1350] = ~((inputs[568]) & (inputs[509]));
    assign layer0_outputs[1351] = ~((inputs[990]) ^ (inputs[526]));
    assign layer0_outputs[1352] = ~(inputs[894]) | (inputs[220]);
    assign layer0_outputs[1353] = ~(inputs[836]) | (inputs[462]);
    assign layer0_outputs[1354] = ~(inputs[93]);
    assign layer0_outputs[1355] = inputs[394];
    assign layer0_outputs[1356] = (inputs[897]) ^ (inputs[559]);
    assign layer0_outputs[1357] = ~(inputs[121]) | (inputs[892]);
    assign layer0_outputs[1358] = (inputs[978]) & ~(inputs[907]);
    assign layer0_outputs[1359] = (inputs[683]) | (inputs[714]);
    assign layer0_outputs[1360] = ~(inputs[240]);
    assign layer0_outputs[1361] = ~((inputs[244]) | (inputs[108]));
    assign layer0_outputs[1362] = 1'b0;
    assign layer0_outputs[1363] = ~(inputs[114]) | (inputs[224]);
    assign layer0_outputs[1364] = (inputs[84]) & ~(inputs[704]);
    assign layer0_outputs[1365] = ~((inputs[621]) | (inputs[323]));
    assign layer0_outputs[1366] = ~(inputs[527]);
    assign layer0_outputs[1367] = (inputs[487]) ^ (inputs[656]);
    assign layer0_outputs[1368] = ~(inputs[813]);
    assign layer0_outputs[1369] = (inputs[26]) & ~(inputs[1023]);
    assign layer0_outputs[1370] = inputs[284];
    assign layer0_outputs[1371] = ~((inputs[441]) | (inputs[12]));
    assign layer0_outputs[1372] = ~(inputs[502]) | (inputs[291]);
    assign layer0_outputs[1373] = (inputs[689]) | (inputs[770]);
    assign layer0_outputs[1374] = (inputs[579]) ^ (inputs[620]);
    assign layer0_outputs[1375] = ~((inputs[854]) ^ (inputs[673]));
    assign layer0_outputs[1376] = (inputs[241]) & ~(inputs[797]);
    assign layer0_outputs[1377] = (inputs[524]) | (inputs[533]);
    assign layer0_outputs[1378] = inputs[980];
    assign layer0_outputs[1379] = ~((inputs[50]) & (inputs[357]));
    assign layer0_outputs[1380] = 1'b0;
    assign layer0_outputs[1381] = (inputs[972]) | (inputs[362]);
    assign layer0_outputs[1382] = ~((inputs[583]) ^ (inputs[667]));
    assign layer0_outputs[1383] = ~(inputs[91]) | (inputs[888]);
    assign layer0_outputs[1384] = ~(inputs[425]) | (inputs[142]);
    assign layer0_outputs[1385] = ~((inputs[608]) | (inputs[716]));
    assign layer0_outputs[1386] = ~(inputs[237]) | (inputs[118]);
    assign layer0_outputs[1387] = ~((inputs[705]) ^ (inputs[971]));
    assign layer0_outputs[1388] = ~((inputs[520]) | (inputs[473]));
    assign layer0_outputs[1389] = (inputs[769]) ^ (inputs[566]);
    assign layer0_outputs[1390] = (inputs[519]) | (inputs[390]);
    assign layer0_outputs[1391] = (inputs[32]) & (inputs[38]);
    assign layer0_outputs[1392] = ~(inputs[561]) | (inputs[379]);
    assign layer0_outputs[1393] = ~(inputs[186]) | (inputs[194]);
    assign layer0_outputs[1394] = (inputs[305]) & ~(inputs[380]);
    assign layer0_outputs[1395] = inputs[490];
    assign layer0_outputs[1396] = (inputs[567]) | (inputs[700]);
    assign layer0_outputs[1397] = ~((inputs[67]) | (inputs[953]));
    assign layer0_outputs[1398] = (inputs[591]) | (inputs[822]);
    assign layer0_outputs[1399] = inputs[732];
    assign layer0_outputs[1400] = ~(inputs[931]);
    assign layer0_outputs[1401] = ~(inputs[773]);
    assign layer0_outputs[1402] = (inputs[466]) ^ (inputs[529]);
    assign layer0_outputs[1403] = ~(inputs[787]) | (inputs[231]);
    assign layer0_outputs[1404] = (inputs[817]) & ~(inputs[731]);
    assign layer0_outputs[1405] = (inputs[632]) | (inputs[811]);
    assign layer0_outputs[1406] = ~(inputs[122]);
    assign layer0_outputs[1407] = (inputs[15]) & (inputs[1010]);
    assign layer0_outputs[1408] = ~((inputs[955]) ^ (inputs[874]));
    assign layer0_outputs[1409] = 1'b0;
    assign layer0_outputs[1410] = inputs[589];
    assign layer0_outputs[1411] = (inputs[326]) | (inputs[360]);
    assign layer0_outputs[1412] = inputs[538];
    assign layer0_outputs[1413] = (inputs[65]) ^ (inputs[685]);
    assign layer0_outputs[1414] = (inputs[206]) & ~(inputs[140]);
    assign layer0_outputs[1415] = (inputs[208]) | (inputs[698]);
    assign layer0_outputs[1416] = ~(inputs[965]);
    assign layer0_outputs[1417] = ~(inputs[507]);
    assign layer0_outputs[1418] = ~((inputs[321]) | (inputs[238]));
    assign layer0_outputs[1419] = 1'b0;
    assign layer0_outputs[1420] = inputs[952];
    assign layer0_outputs[1421] = (inputs[425]) ^ (inputs[1006]);
    assign layer0_outputs[1422] = ~(inputs[485]) | (inputs[25]);
    assign layer0_outputs[1423] = inputs[784];
    assign layer0_outputs[1424] = (inputs[656]) ^ (inputs[378]);
    assign layer0_outputs[1425] = ~((inputs[836]) | (inputs[565]));
    assign layer0_outputs[1426] = ~((inputs[771]) | (inputs[751]));
    assign layer0_outputs[1427] = ~(inputs[199]) | (inputs[549]);
    assign layer0_outputs[1428] = (inputs[872]) ^ (inputs[506]);
    assign layer0_outputs[1429] = ~((inputs[8]) ^ (inputs[578]));
    assign layer0_outputs[1430] = ~((inputs[153]) ^ (inputs[283]));
    assign layer0_outputs[1431] = ~(inputs[127]);
    assign layer0_outputs[1432] = (inputs[522]) & ~(inputs[1017]);
    assign layer0_outputs[1433] = inputs[357];
    assign layer0_outputs[1434] = (inputs[222]) & ~(inputs[363]);
    assign layer0_outputs[1435] = (inputs[151]) | (inputs[85]);
    assign layer0_outputs[1436] = inputs[883];
    assign layer0_outputs[1437] = (inputs[1003]) & ~(inputs[544]);
    assign layer0_outputs[1438] = inputs[788];
    assign layer0_outputs[1439] = ~(inputs[526]);
    assign layer0_outputs[1440] = ~(inputs[179]) | (inputs[406]);
    assign layer0_outputs[1441] = ~((inputs[400]) | (inputs[372]));
    assign layer0_outputs[1442] = ~((inputs[951]) | (inputs[587]));
    assign layer0_outputs[1443] = (inputs[774]) & ~(inputs[547]);
    assign layer0_outputs[1444] = (inputs[732]) | (inputs[391]);
    assign layer0_outputs[1445] = (inputs[651]) & ~(inputs[288]);
    assign layer0_outputs[1446] = ~((inputs[180]) ^ (inputs[94]));
    assign layer0_outputs[1447] = inputs[467];
    assign layer0_outputs[1448] = (inputs[515]) | (inputs[668]);
    assign layer0_outputs[1449] = ~(inputs[803]) | (inputs[91]);
    assign layer0_outputs[1450] = ~((inputs[981]) ^ (inputs[475]));
    assign layer0_outputs[1451] = ~(inputs[281]);
    assign layer0_outputs[1452] = ~(inputs[211]) | (inputs[58]);
    assign layer0_outputs[1453] = (inputs[780]) ^ (inputs[510]);
    assign layer0_outputs[1454] = ~(inputs[396]);
    assign layer0_outputs[1455] = (inputs[630]) ^ (inputs[857]);
    assign layer0_outputs[1456] = (inputs[970]) ^ (inputs[813]);
    assign layer0_outputs[1457] = ~(inputs[586]);
    assign layer0_outputs[1458] = (inputs[85]) | (inputs[858]);
    assign layer0_outputs[1459] = inputs[614];
    assign layer0_outputs[1460] = inputs[786];
    assign layer0_outputs[1461] = ~((inputs[164]) & (inputs[282]));
    assign layer0_outputs[1462] = inputs[434];
    assign layer0_outputs[1463] = inputs[791];
    assign layer0_outputs[1464] = (inputs[723]) & ~(inputs[37]);
    assign layer0_outputs[1465] = (inputs[664]) | (inputs[288]);
    assign layer0_outputs[1466] = ~(inputs[628]);
    assign layer0_outputs[1467] = inputs[944];
    assign layer0_outputs[1468] = ~((inputs[622]) | (inputs[227]));
    assign layer0_outputs[1469] = ~(inputs[521]) | (inputs[128]);
    assign layer0_outputs[1470] = ~((inputs[375]) | (inputs[176]));
    assign layer0_outputs[1471] = ~(inputs[218]) | (inputs[952]);
    assign layer0_outputs[1472] = 1'b1;
    assign layer0_outputs[1473] = ~(inputs[171]);
    assign layer0_outputs[1474] = inputs[660];
    assign layer0_outputs[1475] = (inputs[81]) & ~(inputs[178]);
    assign layer0_outputs[1476] = ~(inputs[237]) | (inputs[81]);
    assign layer0_outputs[1477] = (inputs[566]) | (inputs[397]);
    assign layer0_outputs[1478] = inputs[897];
    assign layer0_outputs[1479] = (inputs[78]) & ~(inputs[888]);
    assign layer0_outputs[1480] = ~(inputs[33]);
    assign layer0_outputs[1481] = (inputs[199]) | (inputs[792]);
    assign layer0_outputs[1482] = ~(inputs[282]) | (inputs[826]);
    assign layer0_outputs[1483] = (inputs[931]) | (inputs[982]);
    assign layer0_outputs[1484] = ~((inputs[979]) ^ (inputs[461]));
    assign layer0_outputs[1485] = ~(inputs[461]);
    assign layer0_outputs[1486] = inputs[902];
    assign layer0_outputs[1487] = (inputs[1016]) | (inputs[1020]);
    assign layer0_outputs[1488] = ~((inputs[4]) ^ (inputs[247]));
    assign layer0_outputs[1489] = ~((inputs[838]) | (inputs[863]));
    assign layer0_outputs[1490] = ~((inputs[607]) & (inputs[140]));
    assign layer0_outputs[1491] = (inputs[532]) & ~(inputs[844]);
    assign layer0_outputs[1492] = (inputs[624]) & ~(inputs[523]);
    assign layer0_outputs[1493] = ~(inputs[615]) | (inputs[479]);
    assign layer0_outputs[1494] = ~((inputs[116]) | (inputs[621]));
    assign layer0_outputs[1495] = ~(inputs[746]) | (inputs[685]);
    assign layer0_outputs[1496] = ~(inputs[187]) | (inputs[49]);
    assign layer0_outputs[1497] = ~(inputs[816]) | (inputs[766]);
    assign layer0_outputs[1498] = ~(inputs[535]);
    assign layer0_outputs[1499] = inputs[813];
    assign layer0_outputs[1500] = inputs[559];
    assign layer0_outputs[1501] = 1'b0;
    assign layer0_outputs[1502] = 1'b0;
    assign layer0_outputs[1503] = ~(inputs[159]) | (inputs[927]);
    assign layer0_outputs[1504] = (inputs[780]) & ~(inputs[642]);
    assign layer0_outputs[1505] = (inputs[1006]) & ~(inputs[735]);
    assign layer0_outputs[1506] = ~(inputs[49]);
    assign layer0_outputs[1507] = (inputs[587]) & ~(inputs[929]);
    assign layer0_outputs[1508] = (inputs[475]) ^ (inputs[918]);
    assign layer0_outputs[1509] = 1'b0;
    assign layer0_outputs[1510] = ~((inputs[73]) | (inputs[62]));
    assign layer0_outputs[1511] = ~((inputs[2]) | (inputs[89]));
    assign layer0_outputs[1512] = inputs[205];
    assign layer0_outputs[1513] = (inputs[925]) | (inputs[546]);
    assign layer0_outputs[1514] = inputs[582];
    assign layer0_outputs[1515] = ~(inputs[404]);
    assign layer0_outputs[1516] = ~((inputs[187]) | (inputs[498]));
    assign layer0_outputs[1517] = ~(inputs[881]);
    assign layer0_outputs[1518] = inputs[686];
    assign layer0_outputs[1519] = (inputs[720]) & ~(inputs[545]);
    assign layer0_outputs[1520] = ~((inputs[144]) | (inputs[606]));
    assign layer0_outputs[1521] = ~((inputs[710]) | (inputs[942]));
    assign layer0_outputs[1522] = ~((inputs[5]) & (inputs[997]));
    assign layer0_outputs[1523] = inputs[298];
    assign layer0_outputs[1524] = ~(inputs[882]);
    assign layer0_outputs[1525] = ~((inputs[900]) ^ (inputs[220]));
    assign layer0_outputs[1526] = ~(inputs[79]);
    assign layer0_outputs[1527] = ~(inputs[430]) | (inputs[140]);
    assign layer0_outputs[1528] = ~((inputs[711]) ^ (inputs[131]));
    assign layer0_outputs[1529] = ~((inputs[319]) | (inputs[800]));
    assign layer0_outputs[1530] = ~((inputs[141]) ^ (inputs[481]));
    assign layer0_outputs[1531] = ~((inputs[708]) & (inputs[415]));
    assign layer0_outputs[1532] = (inputs[35]) ^ (inputs[947]);
    assign layer0_outputs[1533] = ~(inputs[1009]);
    assign layer0_outputs[1534] = inputs[277];
    assign layer0_outputs[1535] = ~((inputs[68]) ^ (inputs[469]));
    assign layer0_outputs[1536] = (inputs[224]) & ~(inputs[859]);
    assign layer0_outputs[1537] = inputs[556];
    assign layer0_outputs[1538] = ~(inputs[722]) | (inputs[965]);
    assign layer0_outputs[1539] = 1'b1;
    assign layer0_outputs[1540] = inputs[950];
    assign layer0_outputs[1541] = ~(inputs[350]);
    assign layer0_outputs[1542] = (inputs[213]) & (inputs[0]);
    assign layer0_outputs[1543] = ~(inputs[718]) | (inputs[677]);
    assign layer0_outputs[1544] = ~(inputs[862]);
    assign layer0_outputs[1545] = (inputs[957]) & ~(inputs[298]);
    assign layer0_outputs[1546] = ~((inputs[68]) ^ (inputs[131]));
    assign layer0_outputs[1547] = (inputs[2]) & ~(inputs[613]);
    assign layer0_outputs[1548] = (inputs[916]) | (inputs[596]);
    assign layer0_outputs[1549] = 1'b0;
    assign layer0_outputs[1550] = ~(inputs[945]);
    assign layer0_outputs[1551] = inputs[754];
    assign layer0_outputs[1552] = inputs[105];
    assign layer0_outputs[1553] = ~(inputs[273]);
    assign layer0_outputs[1554] = ~(inputs[598]) | (inputs[414]);
    assign layer0_outputs[1555] = (inputs[795]) & (inputs[54]);
    assign layer0_outputs[1556] = ~((inputs[448]) ^ (inputs[70]));
    assign layer0_outputs[1557] = ~(inputs[206]);
    assign layer0_outputs[1558] = inputs[496];
    assign layer0_outputs[1559] = (inputs[775]) ^ (inputs[684]);
    assign layer0_outputs[1560] = (inputs[218]) ^ (inputs[750]);
    assign layer0_outputs[1561] = ~((inputs[817]) | (inputs[262]));
    assign layer0_outputs[1562] = ~(inputs[370]);
    assign layer0_outputs[1563] = ~((inputs[998]) | (inputs[390]));
    assign layer0_outputs[1564] = ~((inputs[45]) & (inputs[455]));
    assign layer0_outputs[1565] = ~((inputs[781]) ^ (inputs[892]));
    assign layer0_outputs[1566] = ~(inputs[321]);
    assign layer0_outputs[1567] = ~(inputs[173]) | (inputs[514]);
    assign layer0_outputs[1568] = ~(inputs[657]) | (inputs[538]);
    assign layer0_outputs[1569] = inputs[467];
    assign layer0_outputs[1570] = inputs[332];
    assign layer0_outputs[1571] = inputs[243];
    assign layer0_outputs[1572] = ~((inputs[241]) & (inputs[246]));
    assign layer0_outputs[1573] = (inputs[566]) | (inputs[256]);
    assign layer0_outputs[1574] = ~((inputs[129]) ^ (inputs[960]));
    assign layer0_outputs[1575] = ~((inputs[503]) | (inputs[165]));
    assign layer0_outputs[1576] = 1'b0;
    assign layer0_outputs[1577] = ~(inputs[614]);
    assign layer0_outputs[1578] = inputs[648];
    assign layer0_outputs[1579] = ~((inputs[494]) | (inputs[825]));
    assign layer0_outputs[1580] = (inputs[753]) & ~(inputs[772]);
    assign layer0_outputs[1581] = (inputs[312]) & (inputs[825]);
    assign layer0_outputs[1582] = ~((inputs[348]) ^ (inputs[909]));
    assign layer0_outputs[1583] = ~(inputs[153]);
    assign layer0_outputs[1584] = (inputs[205]) | (inputs[612]);
    assign layer0_outputs[1585] = (inputs[454]) | (inputs[298]);
    assign layer0_outputs[1586] = ~(inputs[336]) | (inputs[705]);
    assign layer0_outputs[1587] = (inputs[908]) & ~(inputs[1014]);
    assign layer0_outputs[1588] = inputs[663];
    assign layer0_outputs[1589] = ~((inputs[938]) & (inputs[133]));
    assign layer0_outputs[1590] = inputs[846];
    assign layer0_outputs[1591] = (inputs[196]) | (inputs[590]);
    assign layer0_outputs[1592] = ~((inputs[244]) ^ (inputs[273]));
    assign layer0_outputs[1593] = (inputs[279]) | (inputs[287]);
    assign layer0_outputs[1594] = inputs[716];
    assign layer0_outputs[1595] = ~(inputs[744]) | (inputs[55]);
    assign layer0_outputs[1596] = inputs[666];
    assign layer0_outputs[1597] = ~(inputs[779]) | (inputs[1011]);
    assign layer0_outputs[1598] = ~(inputs[318]) | (inputs[669]);
    assign layer0_outputs[1599] = ~(inputs[718]) | (inputs[440]);
    assign layer0_outputs[1600] = ~(inputs[497]);
    assign layer0_outputs[1601] = (inputs[602]) | (inputs[215]);
    assign layer0_outputs[1602] = ~(inputs[967]);
    assign layer0_outputs[1603] = inputs[591];
    assign layer0_outputs[1604] = ~(inputs[521]);
    assign layer0_outputs[1605] = (inputs[779]) ^ (inputs[869]);
    assign layer0_outputs[1606] = (inputs[490]) ^ (inputs[826]);
    assign layer0_outputs[1607] = (inputs[489]) | (inputs[390]);
    assign layer0_outputs[1608] = (inputs[283]) ^ (inputs[339]);
    assign layer0_outputs[1609] = inputs[682];
    assign layer0_outputs[1610] = ~(inputs[312]) | (inputs[733]);
    assign layer0_outputs[1611] = ~((inputs[476]) | (inputs[243]));
    assign layer0_outputs[1612] = (inputs[736]) ^ (inputs[810]);
    assign layer0_outputs[1613] = ~((inputs[566]) ^ (inputs[158]));
    assign layer0_outputs[1614] = ~((inputs[456]) ^ (inputs[62]));
    assign layer0_outputs[1615] = ~(inputs[633]);
    assign layer0_outputs[1616] = ~((inputs[616]) | (inputs[769]));
    assign layer0_outputs[1617] = (inputs[449]) & ~(inputs[505]);
    assign layer0_outputs[1618] = (inputs[424]) & ~(inputs[88]);
    assign layer0_outputs[1619] = ~(inputs[623]);
    assign layer0_outputs[1620] = ~(inputs[276]) | (inputs[999]);
    assign layer0_outputs[1621] = ~(inputs[285]) | (inputs[833]);
    assign layer0_outputs[1622] = ~(inputs[786]);
    assign layer0_outputs[1623] = (inputs[31]) | (inputs[555]);
    assign layer0_outputs[1624] = ~(inputs[1010]) | (inputs[360]);
    assign layer0_outputs[1625] = ~(inputs[378]);
    assign layer0_outputs[1626] = ~((inputs[666]) | (inputs[137]));
    assign layer0_outputs[1627] = ~((inputs[1000]) ^ (inputs[424]));
    assign layer0_outputs[1628] = inputs[134];
    assign layer0_outputs[1629] = ~((inputs[136]) & (inputs[882]));
    assign layer0_outputs[1630] = (inputs[680]) | (inputs[791]);
    assign layer0_outputs[1631] = ~((inputs[625]) & (inputs[83]));
    assign layer0_outputs[1632] = (inputs[688]) & ~(inputs[460]);
    assign layer0_outputs[1633] = (inputs[602]) & ~(inputs[69]);
    assign layer0_outputs[1634] = ~((inputs[371]) | (inputs[481]));
    assign layer0_outputs[1635] = 1'b1;
    assign layer0_outputs[1636] = ~(inputs[233]) | (inputs[6]);
    assign layer0_outputs[1637] = ~((inputs[288]) ^ (inputs[561]));
    assign layer0_outputs[1638] = ~((inputs[858]) ^ (inputs[179]));
    assign layer0_outputs[1639] = ~(inputs[338]);
    assign layer0_outputs[1640] = inputs[686];
    assign layer0_outputs[1641] = (inputs[369]) & ~(inputs[919]);
    assign layer0_outputs[1642] = ~(inputs[506]);
    assign layer0_outputs[1643] = ~(inputs[736]);
    assign layer0_outputs[1644] = ~((inputs[624]) | (inputs[1008]));
    assign layer0_outputs[1645] = inputs[464];
    assign layer0_outputs[1646] = (inputs[1015]) | (inputs[332]);
    assign layer0_outputs[1647] = ~(inputs[365]);
    assign layer0_outputs[1648] = ~((inputs[297]) | (inputs[40]));
    assign layer0_outputs[1649] = ~(inputs[758]) | (inputs[7]);
    assign layer0_outputs[1650] = inputs[241];
    assign layer0_outputs[1651] = inputs[988];
    assign layer0_outputs[1652] = ~(inputs[458]) | (inputs[255]);
    assign layer0_outputs[1653] = ~(inputs[409]) | (inputs[326]);
    assign layer0_outputs[1654] = inputs[211];
    assign layer0_outputs[1655] = (inputs[404]) & (inputs[563]);
    assign layer0_outputs[1656] = ~(inputs[888]) | (inputs[76]);
    assign layer0_outputs[1657] = inputs[225];
    assign layer0_outputs[1658] = ~((inputs[171]) ^ (inputs[97]));
    assign layer0_outputs[1659] = (inputs[21]) | (inputs[877]);
    assign layer0_outputs[1660] = ~((inputs[118]) ^ (inputs[453]));
    assign layer0_outputs[1661] = (inputs[292]) & (inputs[138]);
    assign layer0_outputs[1662] = (inputs[345]) | (inputs[191]);
    assign layer0_outputs[1663] = inputs[651];
    assign layer0_outputs[1664] = (inputs[808]) | (inputs[979]);
    assign layer0_outputs[1665] = ~((inputs[326]) | (inputs[264]));
    assign layer0_outputs[1666] = (inputs[201]) | (inputs[17]);
    assign layer0_outputs[1667] = ~(inputs[241]);
    assign layer0_outputs[1668] = inputs[846];
    assign layer0_outputs[1669] = (inputs[740]) | (inputs[466]);
    assign layer0_outputs[1670] = (inputs[800]) & ~(inputs[417]);
    assign layer0_outputs[1671] = (inputs[855]) & ~(inputs[48]);
    assign layer0_outputs[1672] = (inputs[642]) ^ (inputs[267]);
    assign layer0_outputs[1673] = (inputs[676]) | (inputs[306]);
    assign layer0_outputs[1674] = ~((inputs[526]) ^ (inputs[574]));
    assign layer0_outputs[1675] = ~(inputs[726]) | (inputs[282]);
    assign layer0_outputs[1676] = inputs[464];
    assign layer0_outputs[1677] = (inputs[888]) | (inputs[989]);
    assign layer0_outputs[1678] = (inputs[138]) | (inputs[602]);
    assign layer0_outputs[1679] = inputs[260];
    assign layer0_outputs[1680] = (inputs[643]) & (inputs[577]);
    assign layer0_outputs[1681] = ~((inputs[203]) ^ (inputs[343]));
    assign layer0_outputs[1682] = ~((inputs[880]) | (inputs[791]));
    assign layer0_outputs[1683] = 1'b1;
    assign layer0_outputs[1684] = ~(inputs[339]);
    assign layer0_outputs[1685] = (inputs[26]) ^ (inputs[171]);
    assign layer0_outputs[1686] = ~(inputs[528]);
    assign layer0_outputs[1687] = (inputs[974]) | (inputs[163]);
    assign layer0_outputs[1688] = ~(inputs[839]);
    assign layer0_outputs[1689] = ~(inputs[374]) | (inputs[472]);
    assign layer0_outputs[1690] = (inputs[128]) & (inputs[920]);
    assign layer0_outputs[1691] = 1'b0;
    assign layer0_outputs[1692] = ~((inputs[696]) | (inputs[743]));
    assign layer0_outputs[1693] = inputs[753];
    assign layer0_outputs[1694] = ~(inputs[524]);
    assign layer0_outputs[1695] = ~((inputs[654]) | (inputs[736]));
    assign layer0_outputs[1696] = ~((inputs[80]) | (inputs[509]));
    assign layer0_outputs[1697] = ~((inputs[553]) | (inputs[657]));
    assign layer0_outputs[1698] = ~(inputs[104]) | (inputs[408]);
    assign layer0_outputs[1699] = (inputs[37]) & (inputs[256]);
    assign layer0_outputs[1700] = inputs[264];
    assign layer0_outputs[1701] = (inputs[710]) | (inputs[876]);
    assign layer0_outputs[1702] = (inputs[74]) & ~(inputs[831]);
    assign layer0_outputs[1703] = inputs[858];
    assign layer0_outputs[1704] = ~(inputs[1007]);
    assign layer0_outputs[1705] = ~(inputs[401]);
    assign layer0_outputs[1706] = ~((inputs[181]) | (inputs[925]));
    assign layer0_outputs[1707] = (inputs[72]) ^ (inputs[1010]);
    assign layer0_outputs[1708] = (inputs[418]) & ~(inputs[115]);
    assign layer0_outputs[1709] = ~(inputs[457]);
    assign layer0_outputs[1710] = ~((inputs[695]) | (inputs[869]));
    assign layer0_outputs[1711] = (inputs[816]) & ~(inputs[144]);
    assign layer0_outputs[1712] = inputs[464];
    assign layer0_outputs[1713] = (inputs[475]) & (inputs[475]);
    assign layer0_outputs[1714] = (inputs[845]) | (inputs[518]);
    assign layer0_outputs[1715] = ~(inputs[61]);
    assign layer0_outputs[1716] = ~(inputs[474]);
    assign layer0_outputs[1717] = ~((inputs[940]) ^ (inputs[739]));
    assign layer0_outputs[1718] = (inputs[48]) ^ (inputs[616]);
    assign layer0_outputs[1719] = ~((inputs[869]) | (inputs[94]));
    assign layer0_outputs[1720] = ~(inputs[916]);
    assign layer0_outputs[1721] = ~((inputs[63]) | (inputs[971]));
    assign layer0_outputs[1722] = 1'b0;
    assign layer0_outputs[1723] = (inputs[284]) ^ (inputs[749]);
    assign layer0_outputs[1724] = ~(inputs[329]);
    assign layer0_outputs[1725] = ~((inputs[905]) ^ (inputs[323]));
    assign layer0_outputs[1726] = 1'b0;
    assign layer0_outputs[1727] = (inputs[719]) | (inputs[165]);
    assign layer0_outputs[1728] = ~((inputs[380]) & (inputs[164]));
    assign layer0_outputs[1729] = ~((inputs[488]) | (inputs[26]));
    assign layer0_outputs[1730] = ~(inputs[615]);
    assign layer0_outputs[1731] = inputs[925];
    assign layer0_outputs[1732] = (inputs[418]) ^ (inputs[140]);
    assign layer0_outputs[1733] = (inputs[176]) & ~(inputs[190]);
    assign layer0_outputs[1734] = ~(inputs[331]) | (inputs[94]);
    assign layer0_outputs[1735] = ~(inputs[433]);
    assign layer0_outputs[1736] = ~((inputs[714]) ^ (inputs[945]));
    assign layer0_outputs[1737] = ~(inputs[919]) | (inputs[861]);
    assign layer0_outputs[1738] = inputs[649];
    assign layer0_outputs[1739] = ~(inputs[293]) | (inputs[646]);
    assign layer0_outputs[1740] = ~((inputs[561]) | (inputs[743]));
    assign layer0_outputs[1741] = (inputs[108]) | (inputs[595]);
    assign layer0_outputs[1742] = (inputs[840]) & ~(inputs[18]);
    assign layer0_outputs[1743] = inputs[333];
    assign layer0_outputs[1744] = (inputs[662]) | (inputs[966]);
    assign layer0_outputs[1745] = ~(inputs[164]);
    assign layer0_outputs[1746] = (inputs[626]) & ~(inputs[896]);
    assign layer0_outputs[1747] = (inputs[12]) & ~(inputs[137]);
    assign layer0_outputs[1748] = inputs[132];
    assign layer0_outputs[1749] = ~((inputs[86]) | (inputs[153]));
    assign layer0_outputs[1750] = ~(inputs[632]) | (inputs[4]);
    assign layer0_outputs[1751] = (inputs[262]) | (inputs[113]);
    assign layer0_outputs[1752] = ~(inputs[914]);
    assign layer0_outputs[1753] = (inputs[1013]) | (inputs[436]);
    assign layer0_outputs[1754] = ~((inputs[166]) ^ (inputs[668]));
    assign layer0_outputs[1755] = ~(inputs[507]);
    assign layer0_outputs[1756] = ~((inputs[263]) & (inputs[793]));
    assign layer0_outputs[1757] = (inputs[188]) | (inputs[233]);
    assign layer0_outputs[1758] = inputs[999];
    assign layer0_outputs[1759] = ~(inputs[370]) | (inputs[422]);
    assign layer0_outputs[1760] = 1'b0;
    assign layer0_outputs[1761] = ~((inputs[745]) | (inputs[209]));
    assign layer0_outputs[1762] = ~(inputs[523]);
    assign layer0_outputs[1763] = ~(inputs[431]) | (inputs[1004]);
    assign layer0_outputs[1764] = (inputs[301]) & ~(inputs[433]);
    assign layer0_outputs[1765] = ~(inputs[235]);
    assign layer0_outputs[1766] = ~(inputs[239]) | (inputs[127]);
    assign layer0_outputs[1767] = (inputs[417]) ^ (inputs[298]);
    assign layer0_outputs[1768] = (inputs[57]) & (inputs[257]);
    assign layer0_outputs[1769] = ~((inputs[368]) | (inputs[1013]));
    assign layer0_outputs[1770] = ~((inputs[245]) ^ (inputs[631]));
    assign layer0_outputs[1771] = inputs[948];
    assign layer0_outputs[1772] = ~((inputs[594]) & (inputs[305]));
    assign layer0_outputs[1773] = (inputs[218]) & ~(inputs[468]);
    assign layer0_outputs[1774] = ~((inputs[972]) ^ (inputs[183]));
    assign layer0_outputs[1775] = inputs[428];
    assign layer0_outputs[1776] = ~(inputs[414]) | (inputs[989]);
    assign layer0_outputs[1777] = ~((inputs[889]) ^ (inputs[150]));
    assign layer0_outputs[1778] = (inputs[560]) & ~(inputs[969]);
    assign layer0_outputs[1779] = (inputs[764]) | (inputs[266]);
    assign layer0_outputs[1780] = ~((inputs[182]) | (inputs[776]));
    assign layer0_outputs[1781] = (inputs[291]) | (inputs[665]);
    assign layer0_outputs[1782] = ~((inputs[635]) | (inputs[268]));
    assign layer0_outputs[1783] = ~((inputs[461]) ^ (inputs[155]));
    assign layer0_outputs[1784] = inputs[875];
    assign layer0_outputs[1785] = ~(inputs[912]);
    assign layer0_outputs[1786] = ~(inputs[993]) | (inputs[999]);
    assign layer0_outputs[1787] = ~((inputs[68]) | (inputs[708]));
    assign layer0_outputs[1788] = inputs[36];
    assign layer0_outputs[1789] = inputs[118];
    assign layer0_outputs[1790] = ~((inputs[508]) ^ (inputs[181]));
    assign layer0_outputs[1791] = (inputs[787]) & ~(inputs[1023]);
    assign layer0_outputs[1792] = ~(inputs[271]) | (inputs[106]);
    assign layer0_outputs[1793] = ~(inputs[337]) | (inputs[317]);
    assign layer0_outputs[1794] = inputs[218];
    assign layer0_outputs[1795] = ~((inputs[741]) | (inputs[568]));
    assign layer0_outputs[1796] = inputs[896];
    assign layer0_outputs[1797] = (inputs[57]) ^ (inputs[498]);
    assign layer0_outputs[1798] = (inputs[633]) | (inputs[900]);
    assign layer0_outputs[1799] = (inputs[411]) | (inputs[394]);
    assign layer0_outputs[1800] = ~((inputs[663]) & (inputs[425]));
    assign layer0_outputs[1801] = (inputs[459]) & ~(inputs[903]);
    assign layer0_outputs[1802] = (inputs[467]) & ~(inputs[602]);
    assign layer0_outputs[1803] = (inputs[557]) & ~(inputs[70]);
    assign layer0_outputs[1804] = (inputs[341]) & ~(inputs[916]);
    assign layer0_outputs[1805] = ~(inputs[714]) | (inputs[710]);
    assign layer0_outputs[1806] = inputs[249];
    assign layer0_outputs[1807] = ~(inputs[521]);
    assign layer0_outputs[1808] = ~(inputs[842]) | (inputs[888]);
    assign layer0_outputs[1809] = ~(inputs[426]) | (inputs[908]);
    assign layer0_outputs[1810] = ~(inputs[350]);
    assign layer0_outputs[1811] = ~(inputs[847]);
    assign layer0_outputs[1812] = (inputs[789]) & ~(inputs[802]);
    assign layer0_outputs[1813] = ~((inputs[691]) | (inputs[725]));
    assign layer0_outputs[1814] = (inputs[847]) ^ (inputs[611]);
    assign layer0_outputs[1815] = inputs[691];
    assign layer0_outputs[1816] = ~((inputs[531]) | (inputs[372]));
    assign layer0_outputs[1817] = (inputs[262]) & ~(inputs[46]);
    assign layer0_outputs[1818] = inputs[42];
    assign layer0_outputs[1819] = ~(inputs[591]);
    assign layer0_outputs[1820] = (inputs[353]) | (inputs[856]);
    assign layer0_outputs[1821] = ~((inputs[236]) | (inputs[223]));
    assign layer0_outputs[1822] = (inputs[202]) & ~(inputs[1014]);
    assign layer0_outputs[1823] = (inputs[48]) | (inputs[477]);
    assign layer0_outputs[1824] = ~((inputs[263]) | (inputs[579]));
    assign layer0_outputs[1825] = (inputs[784]) & ~(inputs[281]);
    assign layer0_outputs[1826] = (inputs[193]) & ~(inputs[184]);
    assign layer0_outputs[1827] = ~(inputs[495]);
    assign layer0_outputs[1828] = (inputs[867]) | (inputs[314]);
    assign layer0_outputs[1829] = (inputs[589]) & ~(inputs[964]);
    assign layer0_outputs[1830] = ~(inputs[554]);
    assign layer0_outputs[1831] = ~(inputs[1020]);
    assign layer0_outputs[1832] = ~(inputs[606]) | (inputs[580]);
    assign layer0_outputs[1833] = ~(inputs[141]) | (inputs[14]);
    assign layer0_outputs[1834] = ~(inputs[306]);
    assign layer0_outputs[1835] = ~((inputs[53]) & (inputs[164]));
    assign layer0_outputs[1836] = ~(inputs[957]);
    assign layer0_outputs[1837] = (inputs[638]) ^ (inputs[704]);
    assign layer0_outputs[1838] = ~(inputs[637]);
    assign layer0_outputs[1839] = (inputs[689]) & ~(inputs[864]);
    assign layer0_outputs[1840] = (inputs[601]) & ~(inputs[384]);
    assign layer0_outputs[1841] = ~(inputs[662]) | (inputs[232]);
    assign layer0_outputs[1842] = (inputs[566]) & (inputs[245]);
    assign layer0_outputs[1843] = (inputs[150]) ^ (inputs[851]);
    assign layer0_outputs[1844] = 1'b1;
    assign layer0_outputs[1845] = (inputs[955]) & ~(inputs[935]);
    assign layer0_outputs[1846] = ~((inputs[142]) ^ (inputs[409]));
    assign layer0_outputs[1847] = ~(inputs[401]) | (inputs[335]);
    assign layer0_outputs[1848] = inputs[659];
    assign layer0_outputs[1849] = (inputs[816]) & ~(inputs[1022]);
    assign layer0_outputs[1850] = ~((inputs[890]) & (inputs[77]));
    assign layer0_outputs[1851] = ~(inputs[437]);
    assign layer0_outputs[1852] = ~((inputs[857]) ^ (inputs[59]));
    assign layer0_outputs[1853] = ~((inputs[1009]) | (inputs[7]));
    assign layer0_outputs[1854] = inputs[661];
    assign layer0_outputs[1855] = (inputs[910]) | (inputs[466]);
    assign layer0_outputs[1856] = (inputs[374]) & ~(inputs[538]);
    assign layer0_outputs[1857] = ~((inputs[250]) | (inputs[410]));
    assign layer0_outputs[1858] = (inputs[728]) & ~(inputs[293]);
    assign layer0_outputs[1859] = ~(inputs[522]);
    assign layer0_outputs[1860] = ~((inputs[664]) ^ (inputs[772]));
    assign layer0_outputs[1861] = ~(inputs[304]);
    assign layer0_outputs[1862] = ~((inputs[400]) | (inputs[540]));
    assign layer0_outputs[1863] = ~((inputs[64]) & (inputs[827]));
    assign layer0_outputs[1864] = (inputs[439]) | (inputs[728]);
    assign layer0_outputs[1865] = ~(inputs[478]);
    assign layer0_outputs[1866] = ~((inputs[365]) ^ (inputs[455]));
    assign layer0_outputs[1867] = ~(inputs[713]);
    assign layer0_outputs[1868] = inputs[615];
    assign layer0_outputs[1869] = inputs[365];
    assign layer0_outputs[1870] = ~(inputs[456]) | (inputs[228]);
    assign layer0_outputs[1871] = inputs[551];
    assign layer0_outputs[1872] = (inputs[35]) & ~(inputs[739]);
    assign layer0_outputs[1873] = (inputs[271]) | (inputs[171]);
    assign layer0_outputs[1874] = (inputs[24]) | (inputs[623]);
    assign layer0_outputs[1875] = inputs[939];
    assign layer0_outputs[1876] = ~(inputs[210]) | (inputs[182]);
    assign layer0_outputs[1877] = ~(inputs[685]);
    assign layer0_outputs[1878] = (inputs[648]) | (inputs[1005]);
    assign layer0_outputs[1879] = (inputs[817]) & ~(inputs[946]);
    assign layer0_outputs[1880] = ~((inputs[804]) ^ (inputs[832]));
    assign layer0_outputs[1881] = ~((inputs[771]) ^ (inputs[482]));
    assign layer0_outputs[1882] = (inputs[519]) & ~(inputs[736]);
    assign layer0_outputs[1883] = (inputs[697]) | (inputs[450]);
    assign layer0_outputs[1884] = ~((inputs[88]) ^ (inputs[557]));
    assign layer0_outputs[1885] = inputs[873];
    assign layer0_outputs[1886] = ~(inputs[500]);
    assign layer0_outputs[1887] = (inputs[962]) & (inputs[3]);
    assign layer0_outputs[1888] = ~((inputs[853]) | (inputs[391]));
    assign layer0_outputs[1889] = ~(inputs[535]);
    assign layer0_outputs[1890] = inputs[191];
    assign layer0_outputs[1891] = (inputs[308]) | (inputs[239]);
    assign layer0_outputs[1892] = (inputs[131]) & ~(inputs[603]);
    assign layer0_outputs[1893] = ~((inputs[430]) ^ (inputs[950]));
    assign layer0_outputs[1894] = ~(inputs[944]);
    assign layer0_outputs[1895] = ~(inputs[221]);
    assign layer0_outputs[1896] = ~((inputs[812]) | (inputs[340]));
    assign layer0_outputs[1897] = inputs[168];
    assign layer0_outputs[1898] = ~((inputs[429]) | (inputs[817]));
    assign layer0_outputs[1899] = (inputs[681]) & (inputs[843]);
    assign layer0_outputs[1900] = inputs[546];
    assign layer0_outputs[1901] = (inputs[667]) | (inputs[298]);
    assign layer0_outputs[1902] = ~((inputs[679]) | (inputs[835]));
    assign layer0_outputs[1903] = ~(inputs[312]);
    assign layer0_outputs[1904] = ~(inputs[382]) | (inputs[132]);
    assign layer0_outputs[1905] = (inputs[327]) & (inputs[22]);
    assign layer0_outputs[1906] = ~((inputs[789]) | (inputs[780]));
    assign layer0_outputs[1907] = ~((inputs[1]) & (inputs[709]));
    assign layer0_outputs[1908] = ~(inputs[209]);
    assign layer0_outputs[1909] = (inputs[821]) & (inputs[327]);
    assign layer0_outputs[1910] = ~(inputs[949]);
    assign layer0_outputs[1911] = inputs[632];
    assign layer0_outputs[1912] = ~(inputs[686]);
    assign layer0_outputs[1913] = 1'b0;
    assign layer0_outputs[1914] = (inputs[302]) | (inputs[868]);
    assign layer0_outputs[1915] = ~(inputs[242]) | (inputs[86]);
    assign layer0_outputs[1916] = ~(inputs[833]);
    assign layer0_outputs[1917] = (inputs[622]) | (inputs[992]);
    assign layer0_outputs[1918] = 1'b1;
    assign layer0_outputs[1919] = (inputs[502]) | (inputs[1010]);
    assign layer0_outputs[1920] = ~((inputs[929]) & (inputs[227]));
    assign layer0_outputs[1921] = ~((inputs[693]) ^ (inputs[908]));
    assign layer0_outputs[1922] = ~((inputs[1010]) ^ (inputs[618]));
    assign layer0_outputs[1923] = ~(inputs[652]) | (inputs[925]);
    assign layer0_outputs[1924] = (inputs[263]) & ~(inputs[1001]);
    assign layer0_outputs[1925] = (inputs[351]) & ~(inputs[993]);
    assign layer0_outputs[1926] = ~((inputs[321]) ^ (inputs[590]));
    assign layer0_outputs[1927] = (inputs[388]) | (inputs[406]);
    assign layer0_outputs[1928] = ~((inputs[85]) & (inputs[768]));
    assign layer0_outputs[1929] = (inputs[174]) ^ (inputs[468]);
    assign layer0_outputs[1930] = ~((inputs[821]) ^ (inputs[120]));
    assign layer0_outputs[1931] = ~(inputs[440]);
    assign layer0_outputs[1932] = ~((inputs[360]) | (inputs[617]));
    assign layer0_outputs[1933] = ~((inputs[369]) ^ (inputs[787]));
    assign layer0_outputs[1934] = inputs[142];
    assign layer0_outputs[1935] = ~((inputs[777]) & (inputs[617]));
    assign layer0_outputs[1936] = (inputs[890]) ^ (inputs[98]);
    assign layer0_outputs[1937] = ~(inputs[572]);
    assign layer0_outputs[1938] = (inputs[268]) | (inputs[919]);
    assign layer0_outputs[1939] = ~(inputs[725]) | (inputs[534]);
    assign layer0_outputs[1940] = ~((inputs[249]) | (inputs[956]));
    assign layer0_outputs[1941] = ~(inputs[907]) | (inputs[0]);
    assign layer0_outputs[1942] = (inputs[582]) & (inputs[359]);
    assign layer0_outputs[1943] = (inputs[299]) | (inputs[540]);
    assign layer0_outputs[1944] = inputs[652];
    assign layer0_outputs[1945] = (inputs[801]) | (inputs[964]);
    assign layer0_outputs[1946] = inputs[903];
    assign layer0_outputs[1947] = 1'b1;
    assign layer0_outputs[1948] = ~(inputs[333]) | (inputs[22]);
    assign layer0_outputs[1949] = (inputs[993]) & ~(inputs[774]);
    assign layer0_outputs[1950] = ~(inputs[783]);
    assign layer0_outputs[1951] = inputs[163];
    assign layer0_outputs[1952] = ~(inputs[733]) | (inputs[825]);
    assign layer0_outputs[1953] = 1'b0;
    assign layer0_outputs[1954] = (inputs[965]) & ~(inputs[73]);
    assign layer0_outputs[1955] = (inputs[137]) & ~(inputs[989]);
    assign layer0_outputs[1956] = (inputs[619]) & ~(inputs[46]);
    assign layer0_outputs[1957] = ~((inputs[886]) ^ (inputs[313]));
    assign layer0_outputs[1958] = ~(inputs[720]) | (inputs[322]);
    assign layer0_outputs[1959] = ~(inputs[890]) | (inputs[968]);
    assign layer0_outputs[1960] = (inputs[658]) & ~(inputs[1004]);
    assign layer0_outputs[1961] = inputs[712];
    assign layer0_outputs[1962] = ~((inputs[699]) ^ (inputs[41]));
    assign layer0_outputs[1963] = inputs[624];
    assign layer0_outputs[1964] = (inputs[997]) & ~(inputs[403]);
    assign layer0_outputs[1965] = (inputs[855]) ^ (inputs[892]);
    assign layer0_outputs[1966] = inputs[952];
    assign layer0_outputs[1967] = (inputs[1008]) | (inputs[411]);
    assign layer0_outputs[1968] = (inputs[225]) ^ (inputs[127]);
    assign layer0_outputs[1969] = ~((inputs[152]) | (inputs[434]));
    assign layer0_outputs[1970] = ~(inputs[872]);
    assign layer0_outputs[1971] = (inputs[591]) & ~(inputs[503]);
    assign layer0_outputs[1972] = 1'b1;
    assign layer0_outputs[1973] = ~(inputs[201]) | (inputs[899]);
    assign layer0_outputs[1974] = ~(inputs[363]);
    assign layer0_outputs[1975] = (inputs[382]) ^ (inputs[372]);
    assign layer0_outputs[1976] = (inputs[290]) ^ (inputs[978]);
    assign layer0_outputs[1977] = inputs[346];
    assign layer0_outputs[1978] = inputs[377];
    assign layer0_outputs[1979] = ~((inputs[354]) | (inputs[725]));
    assign layer0_outputs[1980] = ~((inputs[156]) | (inputs[272]));
    assign layer0_outputs[1981] = inputs[994];
    assign layer0_outputs[1982] = inputs[74];
    assign layer0_outputs[1983] = ~((inputs[593]) ^ (inputs[961]));
    assign layer0_outputs[1984] = inputs[489];
    assign layer0_outputs[1985] = (inputs[367]) & ~(inputs[586]);
    assign layer0_outputs[1986] = ~((inputs[653]) | (inputs[192]));
    assign layer0_outputs[1987] = ~((inputs[445]) & (inputs[61]));
    assign layer0_outputs[1988] = ~((inputs[399]) ^ (inputs[1011]));
    assign layer0_outputs[1989] = inputs[249];
    assign layer0_outputs[1990] = inputs[536];
    assign layer0_outputs[1991] = inputs[688];
    assign layer0_outputs[1992] = (inputs[236]) ^ (inputs[246]);
    assign layer0_outputs[1993] = (inputs[946]) | (inputs[162]);
    assign layer0_outputs[1994] = ~((inputs[987]) | (inputs[523]));
    assign layer0_outputs[1995] = (inputs[315]) & ~(inputs[428]);
    assign layer0_outputs[1996] = ~((inputs[975]) | (inputs[629]));
    assign layer0_outputs[1997] = inputs[503];
    assign layer0_outputs[1998] = ~((inputs[955]) ^ (inputs[694]));
    assign layer0_outputs[1999] = (inputs[752]) | (inputs[805]);
    assign layer0_outputs[2000] = (inputs[943]) ^ (inputs[882]);
    assign layer0_outputs[2001] = (inputs[386]) ^ (inputs[9]);
    assign layer0_outputs[2002] = ~((inputs[394]) | (inputs[182]));
    assign layer0_outputs[2003] = inputs[549];
    assign layer0_outputs[2004] = ~(inputs[604]);
    assign layer0_outputs[2005] = ~((inputs[234]) | (inputs[906]));
    assign layer0_outputs[2006] = ~(inputs[275]);
    assign layer0_outputs[2007] = (inputs[231]) | (inputs[48]);
    assign layer0_outputs[2008] = (inputs[456]) & ~(inputs[180]);
    assign layer0_outputs[2009] = inputs[754];
    assign layer0_outputs[2010] = (inputs[353]) ^ (inputs[781]);
    assign layer0_outputs[2011] = (inputs[875]) | (inputs[315]);
    assign layer0_outputs[2012] = (inputs[48]) & (inputs[259]);
    assign layer0_outputs[2013] = (inputs[1020]) & (inputs[412]);
    assign layer0_outputs[2014] = inputs[822];
    assign layer0_outputs[2015] = (inputs[207]) | (inputs[566]);
    assign layer0_outputs[2016] = ~(inputs[750]) | (inputs[407]);
    assign layer0_outputs[2017] = (inputs[577]) | (inputs[199]);
    assign layer0_outputs[2018] = ~((inputs[85]) | (inputs[660]));
    assign layer0_outputs[2019] = 1'b0;
    assign layer0_outputs[2020] = (inputs[885]) | (inputs[678]);
    assign layer0_outputs[2021] = ~(inputs[716]);
    assign layer0_outputs[2022] = ~(inputs[1008]);
    assign layer0_outputs[2023] = 1'b1;
    assign layer0_outputs[2024] = ~((inputs[508]) ^ (inputs[567]));
    assign layer0_outputs[2025] = (inputs[397]) | (inputs[909]);
    assign layer0_outputs[2026] = 1'b0;
    assign layer0_outputs[2027] = (inputs[1013]) ^ (inputs[272]);
    assign layer0_outputs[2028] = ~(inputs[270]) | (inputs[917]);
    assign layer0_outputs[2029] = ~((inputs[258]) ^ (inputs[532]));
    assign layer0_outputs[2030] = ~(inputs[584]) | (inputs[889]);
    assign layer0_outputs[2031] = ~((inputs[958]) ^ (inputs[742]));
    assign layer0_outputs[2032] = ~(inputs[570]) | (inputs[611]);
    assign layer0_outputs[2033] = ~(inputs[91]);
    assign layer0_outputs[2034] = (inputs[688]) & ~(inputs[705]);
    assign layer0_outputs[2035] = (inputs[313]) & ~(inputs[612]);
    assign layer0_outputs[2036] = (inputs[795]) | (inputs[180]);
    assign layer0_outputs[2037] = 1'b0;
    assign layer0_outputs[2038] = (inputs[111]) & ~(inputs[388]);
    assign layer0_outputs[2039] = ~((inputs[145]) | (inputs[561]));
    assign layer0_outputs[2040] = ~(inputs[211]) | (inputs[831]);
    assign layer0_outputs[2041] = ~((inputs[65]) | (inputs[982]));
    assign layer0_outputs[2042] = (inputs[603]) ^ (inputs[707]);
    assign layer0_outputs[2043] = ~(inputs[423]) | (inputs[126]);
    assign layer0_outputs[2044] = ~((inputs[725]) ^ (inputs[358]));
    assign layer0_outputs[2045] = inputs[943];
    assign layer0_outputs[2046] = inputs[914];
    assign layer0_outputs[2047] = (inputs[581]) & ~(inputs[491]);
    assign layer0_outputs[2048] = ~((inputs[721]) & (inputs[69]));
    assign layer0_outputs[2049] = ~(inputs[955]) | (inputs[106]);
    assign layer0_outputs[2050] = inputs[212];
    assign layer0_outputs[2051] = (inputs[583]) ^ (inputs[74]);
    assign layer0_outputs[2052] = ~(inputs[59]) | (inputs[108]);
    assign layer0_outputs[2053] = ~((inputs[599]) | (inputs[368]));
    assign layer0_outputs[2054] = inputs[604];
    assign layer0_outputs[2055] = ~(inputs[498]);
    assign layer0_outputs[2056] = ~((inputs[944]) | (inputs[970]));
    assign layer0_outputs[2057] = ~(inputs[658]);
    assign layer0_outputs[2058] = (inputs[475]) ^ (inputs[316]);
    assign layer0_outputs[2059] = 1'b1;
    assign layer0_outputs[2060] = ~(inputs[436]);
    assign layer0_outputs[2061] = ~(inputs[110]);
    assign layer0_outputs[2062] = ~((inputs[925]) | (inputs[80]));
    assign layer0_outputs[2063] = inputs[366];
    assign layer0_outputs[2064] = inputs[461];
    assign layer0_outputs[2065] = inputs[139];
    assign layer0_outputs[2066] = ~((inputs[511]) ^ (inputs[536]));
    assign layer0_outputs[2067] = ~(inputs[401]) | (inputs[40]);
    assign layer0_outputs[2068] = 1'b0;
    assign layer0_outputs[2069] = inputs[206];
    assign layer0_outputs[2070] = ~((inputs[680]) | (inputs[698]));
    assign layer0_outputs[2071] = (inputs[0]) | (inputs[214]);
    assign layer0_outputs[2072] = ~(inputs[765]) | (inputs[574]);
    assign layer0_outputs[2073] = (inputs[662]) & ~(inputs[607]);
    assign layer0_outputs[2074] = (inputs[891]) ^ (inputs[243]);
    assign layer0_outputs[2075] = ~((inputs[290]) ^ (inputs[399]));
    assign layer0_outputs[2076] = inputs[551];
    assign layer0_outputs[2077] = 1'b1;
    assign layer0_outputs[2078] = ~(inputs[544]);
    assign layer0_outputs[2079] = inputs[649];
    assign layer0_outputs[2080] = (inputs[629]) ^ (inputs[455]);
    assign layer0_outputs[2081] = (inputs[735]) & ~(inputs[928]);
    assign layer0_outputs[2082] = ~(inputs[114]) | (inputs[505]);
    assign layer0_outputs[2083] = ~(inputs[593]);
    assign layer0_outputs[2084] = (inputs[121]) & ~(inputs[1022]);
    assign layer0_outputs[2085] = 1'b1;
    assign layer0_outputs[2086] = inputs[538];
    assign layer0_outputs[2087] = (inputs[572]) & ~(inputs[135]);
    assign layer0_outputs[2088] = (inputs[211]) ^ (inputs[759]);
    assign layer0_outputs[2089] = ~((inputs[494]) ^ (inputs[867]));
    assign layer0_outputs[2090] = ~((inputs[560]) ^ (inputs[481]));
    assign layer0_outputs[2091] = (inputs[448]) ^ (inputs[987]);
    assign layer0_outputs[2092] = (inputs[411]) ^ (inputs[350]);
    assign layer0_outputs[2093] = inputs[848];
    assign layer0_outputs[2094] = (inputs[848]) ^ (inputs[141]);
    assign layer0_outputs[2095] = ~(inputs[901]) | (inputs[486]);
    assign layer0_outputs[2096] = ~((inputs[33]) ^ (inputs[149]));
    assign layer0_outputs[2097] = ~(inputs[26]);
    assign layer0_outputs[2098] = (inputs[413]) ^ (inputs[260]);
    assign layer0_outputs[2099] = ~((inputs[165]) & (inputs[449]));
    assign layer0_outputs[2100] = inputs[556];
    assign layer0_outputs[2101] = ~((inputs[162]) & (inputs[513]));
    assign layer0_outputs[2102] = 1'b0;
    assign layer0_outputs[2103] = ~((inputs[17]) | (inputs[337]));
    assign layer0_outputs[2104] = (inputs[333]) & ~(inputs[74]);
    assign layer0_outputs[2105] = ~(inputs[784]);
    assign layer0_outputs[2106] = ~(inputs[876]);
    assign layer0_outputs[2107] = ~(inputs[166]) | (inputs[412]);
    assign layer0_outputs[2108] = ~(inputs[254]);
    assign layer0_outputs[2109] = (inputs[396]) & ~(inputs[613]);
    assign layer0_outputs[2110] = (inputs[444]) | (inputs[448]);
    assign layer0_outputs[2111] = ~(inputs[876]);
    assign layer0_outputs[2112] = ~(inputs[740]);
    assign layer0_outputs[2113] = ~((inputs[976]) ^ (inputs[548]));
    assign layer0_outputs[2114] = 1'b0;
    assign layer0_outputs[2115] = ~(inputs[513]);
    assign layer0_outputs[2116] = ~((inputs[429]) ^ (inputs[485]));
    assign layer0_outputs[2117] = inputs[969];
    assign layer0_outputs[2118] = ~((inputs[985]) & (inputs[999]));
    assign layer0_outputs[2119] = ~((inputs[93]) & (inputs[867]));
    assign layer0_outputs[2120] = ~((inputs[110]) | (inputs[1006]));
    assign layer0_outputs[2121] = (inputs[750]) | (inputs[381]);
    assign layer0_outputs[2122] = ~((inputs[338]) | (inputs[357]));
    assign layer0_outputs[2123] = (inputs[769]) | (inputs[583]);
    assign layer0_outputs[2124] = inputs[330];
    assign layer0_outputs[2125] = ~((inputs[905]) | (inputs[824]));
    assign layer0_outputs[2126] = inputs[776];
    assign layer0_outputs[2127] = ~(inputs[680]) | (inputs[257]);
    assign layer0_outputs[2128] = ~((inputs[63]) ^ (inputs[201]));
    assign layer0_outputs[2129] = inputs[507];
    assign layer0_outputs[2130] = ~((inputs[598]) ^ (inputs[361]));
    assign layer0_outputs[2131] = (inputs[49]) & ~(inputs[923]);
    assign layer0_outputs[2132] = ~(inputs[1006]) | (inputs[34]);
    assign layer0_outputs[2133] = (inputs[227]) | (inputs[501]);
    assign layer0_outputs[2134] = (inputs[169]) | (inputs[980]);
    assign layer0_outputs[2135] = ~((inputs[942]) | (inputs[639]));
    assign layer0_outputs[2136] = (inputs[551]) & ~(inputs[139]);
    assign layer0_outputs[2137] = ~(inputs[850]);
    assign layer0_outputs[2138] = ~((inputs[731]) ^ (inputs[416]));
    assign layer0_outputs[2139] = ~(inputs[67]);
    assign layer0_outputs[2140] = ~(inputs[590]);
    assign layer0_outputs[2141] = ~((inputs[242]) ^ (inputs[731]));
    assign layer0_outputs[2142] = ~((inputs[47]) | (inputs[599]));
    assign layer0_outputs[2143] = inputs[340];
    assign layer0_outputs[2144] = (inputs[524]) & ~(inputs[870]);
    assign layer0_outputs[2145] = inputs[859];
    assign layer0_outputs[2146] = ~(inputs[318]) | (inputs[990]);
    assign layer0_outputs[2147] = ~(inputs[63]) | (inputs[98]);
    assign layer0_outputs[2148] = ~(inputs[480]) | (inputs[544]);
    assign layer0_outputs[2149] = inputs[340];
    assign layer0_outputs[2150] = ~(inputs[523]);
    assign layer0_outputs[2151] = ~(inputs[116]);
    assign layer0_outputs[2152] = ~(inputs[361]) | (inputs[573]);
    assign layer0_outputs[2153] = (inputs[206]) & ~(inputs[36]);
    assign layer0_outputs[2154] = ~(inputs[278]);
    assign layer0_outputs[2155] = 1'b1;
    assign layer0_outputs[2156] = inputs[111];
    assign layer0_outputs[2157] = ~((inputs[9]) | (inputs[885]));
    assign layer0_outputs[2158] = (inputs[170]) & ~(inputs[286]);
    assign layer0_outputs[2159] = ~(inputs[176]);
    assign layer0_outputs[2160] = (inputs[365]) | (inputs[388]);
    assign layer0_outputs[2161] = ~(inputs[592]);
    assign layer0_outputs[2162] = inputs[451];
    assign layer0_outputs[2163] = 1'b1;
    assign layer0_outputs[2164] = (inputs[753]) ^ (inputs[579]);
    assign layer0_outputs[2165] = inputs[561];
    assign layer0_outputs[2166] = (inputs[78]) | (inputs[474]);
    assign layer0_outputs[2167] = ~((inputs[312]) ^ (inputs[70]));
    assign layer0_outputs[2168] = (inputs[0]) & ~(inputs[905]);
    assign layer0_outputs[2169] = (inputs[11]) & ~(inputs[6]);
    assign layer0_outputs[2170] = (inputs[188]) & ~(inputs[570]);
    assign layer0_outputs[2171] = (inputs[562]) ^ (inputs[486]);
    assign layer0_outputs[2172] = (inputs[254]) ^ (inputs[911]);
    assign layer0_outputs[2173] = (inputs[725]) & ~(inputs[970]);
    assign layer0_outputs[2174] = ~((inputs[759]) | (inputs[170]));
    assign layer0_outputs[2175] = ~(inputs[1009]) | (inputs[382]);
    assign layer0_outputs[2176] = ~(inputs[700]) | (inputs[638]);
    assign layer0_outputs[2177] = ~((inputs[341]) | (inputs[18]));
    assign layer0_outputs[2178] = ~(inputs[615]);
    assign layer0_outputs[2179] = (inputs[616]) | (inputs[490]);
    assign layer0_outputs[2180] = ~(inputs[274]);
    assign layer0_outputs[2181] = ~((inputs[488]) | (inputs[879]));
    assign layer0_outputs[2182] = ~((inputs[724]) ^ (inputs[867]));
    assign layer0_outputs[2183] = inputs[890];
    assign layer0_outputs[2184] = ~((inputs[539]) ^ (inputs[465]));
    assign layer0_outputs[2185] = ~((inputs[531]) | (inputs[859]));
    assign layer0_outputs[2186] = (inputs[812]) ^ (inputs[881]);
    assign layer0_outputs[2187] = (inputs[756]) | (inputs[287]);
    assign layer0_outputs[2188] = ~((inputs[556]) ^ (inputs[994]));
    assign layer0_outputs[2189] = inputs[432];
    assign layer0_outputs[2190] = ~((inputs[246]) | (inputs[832]));
    assign layer0_outputs[2191] = ~(inputs[747]);
    assign layer0_outputs[2192] = ~(inputs[540]) | (inputs[1016]);
    assign layer0_outputs[2193] = inputs[329];
    assign layer0_outputs[2194] = ~(inputs[959]);
    assign layer0_outputs[2195] = ~((inputs[213]) | (inputs[67]));
    assign layer0_outputs[2196] = ~((inputs[743]) | (inputs[977]));
    assign layer0_outputs[2197] = 1'b0;
    assign layer0_outputs[2198] = (inputs[840]) & ~(inputs[107]);
    assign layer0_outputs[2199] = (inputs[251]) | (inputs[314]);
    assign layer0_outputs[2200] = (inputs[227]) | (inputs[874]);
    assign layer0_outputs[2201] = (inputs[633]) | (inputs[435]);
    assign layer0_outputs[2202] = ~((inputs[938]) ^ (inputs[428]));
    assign layer0_outputs[2203] = 1'b0;
    assign layer0_outputs[2204] = inputs[322];
    assign layer0_outputs[2205] = 1'b0;
    assign layer0_outputs[2206] = (inputs[769]) & (inputs[202]);
    assign layer0_outputs[2207] = inputs[234];
    assign layer0_outputs[2208] = ~((inputs[951]) | (inputs[202]));
    assign layer0_outputs[2209] = inputs[937];
    assign layer0_outputs[2210] = ~(inputs[643]);
    assign layer0_outputs[2211] = ~((inputs[864]) ^ (inputs[403]));
    assign layer0_outputs[2212] = (inputs[549]) | (inputs[135]);
    assign layer0_outputs[2213] = ~(inputs[684]);
    assign layer0_outputs[2214] = inputs[136];
    assign layer0_outputs[2215] = (inputs[421]) | (inputs[166]);
    assign layer0_outputs[2216] = ~(inputs[743]) | (inputs[988]);
    assign layer0_outputs[2217] = ~((inputs[9]) | (inputs[267]));
    assign layer0_outputs[2218] = (inputs[813]) & ~(inputs[471]);
    assign layer0_outputs[2219] = ~(inputs[454]);
    assign layer0_outputs[2220] = ~(inputs[290]) | (inputs[58]);
    assign layer0_outputs[2221] = 1'b0;
    assign layer0_outputs[2222] = ~((inputs[139]) & (inputs[574]));
    assign layer0_outputs[2223] = (inputs[809]) & ~(inputs[278]);
    assign layer0_outputs[2224] = ~(inputs[469]) | (inputs[213]);
    assign layer0_outputs[2225] = (inputs[394]) & ~(inputs[783]);
    assign layer0_outputs[2226] = (inputs[617]) | (inputs[570]);
    assign layer0_outputs[2227] = ~((inputs[58]) ^ (inputs[936]));
    assign layer0_outputs[2228] = (inputs[287]) & ~(inputs[378]);
    assign layer0_outputs[2229] = ~((inputs[749]) ^ (inputs[737]));
    assign layer0_outputs[2230] = ~(inputs[190]);
    assign layer0_outputs[2231] = ~((inputs[168]) | (inputs[866]));
    assign layer0_outputs[2232] = (inputs[287]) ^ (inputs[32]);
    assign layer0_outputs[2233] = ~(inputs[399]) | (inputs[699]);
    assign layer0_outputs[2234] = ~(inputs[76]);
    assign layer0_outputs[2235] = ~((inputs[956]) ^ (inputs[794]));
    assign layer0_outputs[2236] = ~(inputs[595]) | (inputs[27]);
    assign layer0_outputs[2237] = (inputs[453]) ^ (inputs[851]);
    assign layer0_outputs[2238] = ~((inputs[880]) | (inputs[393]));
    assign layer0_outputs[2239] = (inputs[124]) ^ (inputs[682]);
    assign layer0_outputs[2240] = (inputs[206]) ^ (inputs[161]);
    assign layer0_outputs[2241] = inputs[773];
    assign layer0_outputs[2242] = ~((inputs[552]) | (inputs[335]));
    assign layer0_outputs[2243] = (inputs[724]) & ~(inputs[976]);
    assign layer0_outputs[2244] = ~((inputs[418]) | (inputs[828]));
    assign layer0_outputs[2245] = ~((inputs[702]) | (inputs[817]));
    assign layer0_outputs[2246] = ~((inputs[739]) & (inputs[134]));
    assign layer0_outputs[2247] = (inputs[898]) ^ (inputs[870]);
    assign layer0_outputs[2248] = (inputs[978]) | (inputs[129]);
    assign layer0_outputs[2249] = (inputs[310]) ^ (inputs[849]);
    assign layer0_outputs[2250] = (inputs[920]) | (inputs[727]);
    assign layer0_outputs[2251] = (inputs[229]) & ~(inputs[289]);
    assign layer0_outputs[2252] = (inputs[545]) | (inputs[400]);
    assign layer0_outputs[2253] = 1'b0;
    assign layer0_outputs[2254] = ~(inputs[495]) | (inputs[640]);
    assign layer0_outputs[2255] = ~((inputs[77]) | (inputs[707]));
    assign layer0_outputs[2256] = inputs[363];
    assign layer0_outputs[2257] = inputs[657];
    assign layer0_outputs[2258] = inputs[816];
    assign layer0_outputs[2259] = (inputs[652]) & (inputs[45]);
    assign layer0_outputs[2260] = 1'b1;
    assign layer0_outputs[2261] = ~((inputs[123]) ^ (inputs[676]));
    assign layer0_outputs[2262] = ~((inputs[441]) ^ (inputs[577]));
    assign layer0_outputs[2263] = (inputs[66]) ^ (inputs[860]);
    assign layer0_outputs[2264] = (inputs[278]) | (inputs[730]);
    assign layer0_outputs[2265] = ~(inputs[487]);
    assign layer0_outputs[2266] = ~((inputs[512]) | (inputs[146]));
    assign layer0_outputs[2267] = ~(inputs[177]);
    assign layer0_outputs[2268] = ~(inputs[618]);
    assign layer0_outputs[2269] = ~((inputs[903]) | (inputs[230]));
    assign layer0_outputs[2270] = (inputs[433]) | (inputs[680]);
    assign layer0_outputs[2271] = (inputs[334]) & (inputs[398]);
    assign layer0_outputs[2272] = inputs[492];
    assign layer0_outputs[2273] = (inputs[494]) & ~(inputs[325]);
    assign layer0_outputs[2274] = inputs[85];
    assign layer0_outputs[2275] = ~(inputs[916]) | (inputs[738]);
    assign layer0_outputs[2276] = ~(inputs[983]) | (inputs[40]);
    assign layer0_outputs[2277] = (inputs[711]) | (inputs[559]);
    assign layer0_outputs[2278] = (inputs[62]) & ~(inputs[228]);
    assign layer0_outputs[2279] = ~(inputs[724]) | (inputs[503]);
    assign layer0_outputs[2280] = inputs[399];
    assign layer0_outputs[2281] = ~((inputs[446]) | (inputs[623]));
    assign layer0_outputs[2282] = 1'b0;
    assign layer0_outputs[2283] = ~((inputs[335]) | (inputs[1005]));
    assign layer0_outputs[2284] = (inputs[819]) | (inputs[267]);
    assign layer0_outputs[2285] = ~(inputs[552]);
    assign layer0_outputs[2286] = inputs[938];
    assign layer0_outputs[2287] = (inputs[512]) ^ (inputs[341]);
    assign layer0_outputs[2288] = ~((inputs[277]) & (inputs[285]));
    assign layer0_outputs[2289] = ~(inputs[381]);
    assign layer0_outputs[2290] = (inputs[732]) & ~(inputs[3]);
    assign layer0_outputs[2291] = (inputs[464]) ^ (inputs[323]);
    assign layer0_outputs[2292] = ~(inputs[656]);
    assign layer0_outputs[2293] = ~((inputs[394]) | (inputs[678]));
    assign layer0_outputs[2294] = (inputs[14]) ^ (inputs[178]);
    assign layer0_outputs[2295] = ~(inputs[537]);
    assign layer0_outputs[2296] = (inputs[876]) & (inputs[972]);
    assign layer0_outputs[2297] = ~(inputs[851]) | (inputs[760]);
    assign layer0_outputs[2298] = (inputs[684]) & ~(inputs[167]);
    assign layer0_outputs[2299] = ~(inputs[567]) | (inputs[952]);
    assign layer0_outputs[2300] = (inputs[649]) | (inputs[448]);
    assign layer0_outputs[2301] = ~(inputs[431]);
    assign layer0_outputs[2302] = (inputs[596]) ^ (inputs[729]);
    assign layer0_outputs[2303] = ~(inputs[77]);
    assign layer0_outputs[2304] = 1'b1;
    assign layer0_outputs[2305] = ~(inputs[860]) | (inputs[863]);
    assign layer0_outputs[2306] = (inputs[81]) & ~(inputs[229]);
    assign layer0_outputs[2307] = (inputs[929]) ^ (inputs[917]);
    assign layer0_outputs[2308] = ~(inputs[564]);
    assign layer0_outputs[2309] = (inputs[73]) & ~(inputs[264]);
    assign layer0_outputs[2310] = ~(inputs[696]) | (inputs[814]);
    assign layer0_outputs[2311] = (inputs[983]) ^ (inputs[973]);
    assign layer0_outputs[2312] = ~(inputs[199]) | (inputs[896]);
    assign layer0_outputs[2313] = ~(inputs[637]) | (inputs[25]);
    assign layer0_outputs[2314] = ~((inputs[703]) & (inputs[308]));
    assign layer0_outputs[2315] = ~(inputs[353]);
    assign layer0_outputs[2316] = ~(inputs[439]) | (inputs[120]);
    assign layer0_outputs[2317] = inputs[414];
    assign layer0_outputs[2318] = (inputs[660]) & ~(inputs[82]);
    assign layer0_outputs[2319] = (inputs[74]) & ~(inputs[219]);
    assign layer0_outputs[2320] = (inputs[424]) & ~(inputs[101]);
    assign layer0_outputs[2321] = (inputs[564]) ^ (inputs[125]);
    assign layer0_outputs[2322] = ~(inputs[405]) | (inputs[572]);
    assign layer0_outputs[2323] = (inputs[270]) | (inputs[161]);
    assign layer0_outputs[2324] = inputs[717];
    assign layer0_outputs[2325] = ~(inputs[621]);
    assign layer0_outputs[2326] = ~(inputs[225]) | (inputs[107]);
    assign layer0_outputs[2327] = (inputs[671]) & ~(inputs[112]);
    assign layer0_outputs[2328] = inputs[661];
    assign layer0_outputs[2329] = 1'b0;
    assign layer0_outputs[2330] = 1'b1;
    assign layer0_outputs[2331] = ~(inputs[390]);
    assign layer0_outputs[2332] = inputs[460];
    assign layer0_outputs[2333] = (inputs[984]) ^ (inputs[660]);
    assign layer0_outputs[2334] = ~(inputs[246]);
    assign layer0_outputs[2335] = ~(inputs[536]) | (inputs[1015]);
    assign layer0_outputs[2336] = (inputs[343]) & ~(inputs[390]);
    assign layer0_outputs[2337] = inputs[609];
    assign layer0_outputs[2338] = ~(inputs[297]);
    assign layer0_outputs[2339] = inputs[685];
    assign layer0_outputs[2340] = (inputs[202]) | (inputs[475]);
    assign layer0_outputs[2341] = ~((inputs[422]) | (inputs[969]));
    assign layer0_outputs[2342] = (inputs[13]) | (inputs[1013]);
    assign layer0_outputs[2343] = ~(inputs[685]);
    assign layer0_outputs[2344] = ~((inputs[726]) ^ (inputs[342]));
    assign layer0_outputs[2345] = (inputs[111]) | (inputs[944]);
    assign layer0_outputs[2346] = 1'b0;
    assign layer0_outputs[2347] = (inputs[817]) | (inputs[879]);
    assign layer0_outputs[2348] = ~((inputs[67]) & (inputs[512]));
    assign layer0_outputs[2349] = (inputs[243]) | (inputs[939]);
    assign layer0_outputs[2350] = ~((inputs[76]) | (inputs[267]));
    assign layer0_outputs[2351] = (inputs[172]) ^ (inputs[384]);
    assign layer0_outputs[2352] = ~(inputs[346]) | (inputs[991]);
    assign layer0_outputs[2353] = inputs[432];
    assign layer0_outputs[2354] = ~((inputs[732]) | (inputs[840]));
    assign layer0_outputs[2355] = ~((inputs[537]) | (inputs[64]));
    assign layer0_outputs[2356] = (inputs[654]) ^ (inputs[800]);
    assign layer0_outputs[2357] = (inputs[526]) & ~(inputs[861]);
    assign layer0_outputs[2358] = ~(inputs[994]);
    assign layer0_outputs[2359] = (inputs[25]) & ~(inputs[888]);
    assign layer0_outputs[2360] = inputs[234];
    assign layer0_outputs[2361] = ~((inputs[522]) ^ (inputs[454]));
    assign layer0_outputs[2362] = inputs[294];
    assign layer0_outputs[2363] = inputs[43];
    assign layer0_outputs[2364] = 1'b1;
    assign layer0_outputs[2365] = inputs[240];
    assign layer0_outputs[2366] = ~((inputs[19]) | (inputs[143]));
    assign layer0_outputs[2367] = inputs[272];
    assign layer0_outputs[2368] = (inputs[286]) | (inputs[786]);
    assign layer0_outputs[2369] = ~((inputs[22]) | (inputs[250]));
    assign layer0_outputs[2370] = (inputs[787]) | (inputs[793]);
    assign layer0_outputs[2371] = ~(inputs[464]) | (inputs[419]);
    assign layer0_outputs[2372] = ~((inputs[1003]) | (inputs[692]));
    assign layer0_outputs[2373] = (inputs[860]) & ~(inputs[278]);
    assign layer0_outputs[2374] = ~((inputs[188]) | (inputs[441]));
    assign layer0_outputs[2375] = ~(inputs[1011]) | (inputs[940]);
    assign layer0_outputs[2376] = ~(inputs[245]);
    assign layer0_outputs[2377] = (inputs[696]) | (inputs[278]);
    assign layer0_outputs[2378] = ~(inputs[927]);
    assign layer0_outputs[2379] = ~(inputs[4]);
    assign layer0_outputs[2380] = (inputs[523]) & ~(inputs[585]);
    assign layer0_outputs[2381] = (inputs[284]) & ~(inputs[759]);
    assign layer0_outputs[2382] = ~(inputs[211]);
    assign layer0_outputs[2383] = inputs[679];
    assign layer0_outputs[2384] = (inputs[760]) ^ (inputs[699]);
    assign layer0_outputs[2385] = (inputs[598]) & ~(inputs[743]);
    assign layer0_outputs[2386] = ~(inputs[957]) | (inputs[741]);
    assign layer0_outputs[2387] = (inputs[182]) & ~(inputs[346]);
    assign layer0_outputs[2388] = ~((inputs[730]) ^ (inputs[469]));
    assign layer0_outputs[2389] = ~(inputs[874]);
    assign layer0_outputs[2390] = inputs[522];
    assign layer0_outputs[2391] = inputs[593];
    assign layer0_outputs[2392] = (inputs[634]) ^ (inputs[298]);
    assign layer0_outputs[2393] = ~((inputs[652]) | (inputs[377]));
    assign layer0_outputs[2394] = 1'b1;
    assign layer0_outputs[2395] = (inputs[596]) & ~(inputs[237]);
    assign layer0_outputs[2396] = inputs[627];
    assign layer0_outputs[2397] = (inputs[662]) ^ (inputs[223]);
    assign layer0_outputs[2398] = ~((inputs[295]) | (inputs[292]));
    assign layer0_outputs[2399] = (inputs[11]) ^ (inputs[836]);
    assign layer0_outputs[2400] = ~(inputs[14]) | (inputs[799]);
    assign layer0_outputs[2401] = ~(inputs[114]);
    assign layer0_outputs[2402] = ~(inputs[114]) | (inputs[1016]);
    assign layer0_outputs[2403] = (inputs[684]) & ~(inputs[897]);
    assign layer0_outputs[2404] = ~(inputs[992]);
    assign layer0_outputs[2405] = ~((inputs[250]) | (inputs[187]));
    assign layer0_outputs[2406] = (inputs[464]) & ~(inputs[132]);
    assign layer0_outputs[2407] = ~((inputs[762]) ^ (inputs[510]));
    assign layer0_outputs[2408] = ~(inputs[555]) | (inputs[143]);
    assign layer0_outputs[2409] = ~(inputs[146]) | (inputs[984]);
    assign layer0_outputs[2410] = 1'b1;
    assign layer0_outputs[2411] = ~(inputs[1011]) | (inputs[301]);
    assign layer0_outputs[2412] = (inputs[435]) & ~(inputs[541]);
    assign layer0_outputs[2413] = inputs[834];
    assign layer0_outputs[2414] = ~((inputs[900]) | (inputs[329]));
    assign layer0_outputs[2415] = inputs[719];
    assign layer0_outputs[2416] = inputs[365];
    assign layer0_outputs[2417] = ~(inputs[806]);
    assign layer0_outputs[2418] = ~((inputs[729]) | (inputs[974]));
    assign layer0_outputs[2419] = ~((inputs[259]) | (inputs[121]));
    assign layer0_outputs[2420] = (inputs[645]) ^ (inputs[56]);
    assign layer0_outputs[2421] = ~((inputs[989]) | (inputs[1015]));
    assign layer0_outputs[2422] = ~(inputs[795]);
    assign layer0_outputs[2423] = (inputs[765]) | (inputs[32]);
    assign layer0_outputs[2424] = 1'b1;
    assign layer0_outputs[2425] = ~((inputs[258]) & (inputs[937]));
    assign layer0_outputs[2426] = ~((inputs[167]) ^ (inputs[127]));
    assign layer0_outputs[2427] = ~((inputs[975]) ^ (inputs[73]));
    assign layer0_outputs[2428] = ~((inputs[663]) | (inputs[492]));
    assign layer0_outputs[2429] = ~(inputs[671]);
    assign layer0_outputs[2430] = (inputs[530]) & ~(inputs[744]);
    assign layer0_outputs[2431] = ~(inputs[1018]);
    assign layer0_outputs[2432] = ~((inputs[115]) & (inputs[168]));
    assign layer0_outputs[2433] = ~(inputs[550]);
    assign layer0_outputs[2434] = ~((inputs[343]) | (inputs[294]));
    assign layer0_outputs[2435] = ~(inputs[70]);
    assign layer0_outputs[2436] = ~((inputs[151]) ^ (inputs[962]));
    assign layer0_outputs[2437] = inputs[173];
    assign layer0_outputs[2438] = (inputs[697]) | (inputs[723]);
    assign layer0_outputs[2439] = (inputs[759]) | (inputs[273]);
    assign layer0_outputs[2440] = (inputs[988]) | (inputs[323]);
    assign layer0_outputs[2441] = ~((inputs[253]) ^ (inputs[151]));
    assign layer0_outputs[2442] = (inputs[455]) & ~(inputs[763]);
    assign layer0_outputs[2443] = (inputs[410]) | (inputs[890]);
    assign layer0_outputs[2444] = (inputs[936]) | (inputs[336]);
    assign layer0_outputs[2445] = inputs[754];
    assign layer0_outputs[2446] = ~(inputs[918]) | (inputs[992]);
    assign layer0_outputs[2447] = ~((inputs[909]) | (inputs[395]));
    assign layer0_outputs[2448] = ~(inputs[859]);
    assign layer0_outputs[2449] = inputs[682];
    assign layer0_outputs[2450] = (inputs[428]) & ~(inputs[452]);
    assign layer0_outputs[2451] = ~(inputs[679]);
    assign layer0_outputs[2452] = ~((inputs[674]) ^ (inputs[539]));
    assign layer0_outputs[2453] = ~(inputs[639]) | (inputs[165]);
    assign layer0_outputs[2454] = ~((inputs[248]) & (inputs[1021]));
    assign layer0_outputs[2455] = ~(inputs[837]);
    assign layer0_outputs[2456] = ~(inputs[304]) | (inputs[727]);
    assign layer0_outputs[2457] = ~(inputs[1002]);
    assign layer0_outputs[2458] = inputs[628];
    assign layer0_outputs[2459] = ~((inputs[1015]) ^ (inputs[551]));
    assign layer0_outputs[2460] = ~((inputs[478]) | (inputs[352]));
    assign layer0_outputs[2461] = inputs[330];
    assign layer0_outputs[2462] = 1'b1;
    assign layer0_outputs[2463] = (inputs[268]) ^ (inputs[342]);
    assign layer0_outputs[2464] = inputs[776];
    assign layer0_outputs[2465] = (inputs[200]) | (inputs[83]);
    assign layer0_outputs[2466] = ~(inputs[366]) | (inputs[924]);
    assign layer0_outputs[2467] = inputs[115];
    assign layer0_outputs[2468] = inputs[640];
    assign layer0_outputs[2469] = ~((inputs[203]) & (inputs[96]));
    assign layer0_outputs[2470] = inputs[432];
    assign layer0_outputs[2471] = ~((inputs[590]) ^ (inputs[923]));
    assign layer0_outputs[2472] = (inputs[175]) & (inputs[831]);
    assign layer0_outputs[2473] = (inputs[542]) & ~(inputs[41]);
    assign layer0_outputs[2474] = ~((inputs[553]) | (inputs[717]));
    assign layer0_outputs[2475] = (inputs[171]) ^ (inputs[86]);
    assign layer0_outputs[2476] = inputs[294];
    assign layer0_outputs[2477] = ~(inputs[365]);
    assign layer0_outputs[2478] = ~(inputs[686]) | (inputs[156]);
    assign layer0_outputs[2479] = (inputs[358]) | (inputs[504]);
    assign layer0_outputs[2480] = ~((inputs[329]) & (inputs[553]));
    assign layer0_outputs[2481] = ~(inputs[648]) | (inputs[2]);
    assign layer0_outputs[2482] = (inputs[592]) & ~(inputs[301]);
    assign layer0_outputs[2483] = ~((inputs[363]) | (inputs[550]));
    assign layer0_outputs[2484] = (inputs[289]) | (inputs[417]);
    assign layer0_outputs[2485] = ~(inputs[876]);
    assign layer0_outputs[2486] = ~(inputs[592]) | (inputs[583]);
    assign layer0_outputs[2487] = ~((inputs[625]) | (inputs[220]));
    assign layer0_outputs[2488] = (inputs[446]) | (inputs[729]);
    assign layer0_outputs[2489] = (inputs[401]) ^ (inputs[278]);
    assign layer0_outputs[2490] = ~((inputs[442]) ^ (inputs[29]));
    assign layer0_outputs[2491] = ~(inputs[66]);
    assign layer0_outputs[2492] = ~(inputs[300]) | (inputs[516]);
    assign layer0_outputs[2493] = ~(inputs[458]);
    assign layer0_outputs[2494] = ~((inputs[619]) | (inputs[589]));
    assign layer0_outputs[2495] = ~(inputs[435]);
    assign layer0_outputs[2496] = (inputs[748]) & ~(inputs[877]);
    assign layer0_outputs[2497] = (inputs[404]) & ~(inputs[345]);
    assign layer0_outputs[2498] = (inputs[982]) | (inputs[954]);
    assign layer0_outputs[2499] = inputs[379];
    assign layer0_outputs[2500] = ~(inputs[125]);
    assign layer0_outputs[2501] = ~((inputs[829]) | (inputs[824]));
    assign layer0_outputs[2502] = (inputs[236]) & ~(inputs[838]);
    assign layer0_outputs[2503] = inputs[467];
    assign layer0_outputs[2504] = ~((inputs[601]) ^ (inputs[759]));
    assign layer0_outputs[2505] = (inputs[335]) & (inputs[778]);
    assign layer0_outputs[2506] = ~((inputs[392]) & (inputs[649]));
    assign layer0_outputs[2507] = ~(inputs[707]);
    assign layer0_outputs[2508] = ~(inputs[150]);
    assign layer0_outputs[2509] = inputs[245];
    assign layer0_outputs[2510] = (inputs[851]) & (inputs[44]);
    assign layer0_outputs[2511] = ~(inputs[558]);
    assign layer0_outputs[2512] = 1'b1;
    assign layer0_outputs[2513] = ~(inputs[885]) | (inputs[142]);
    assign layer0_outputs[2514] = ~(inputs[249]) | (inputs[543]);
    assign layer0_outputs[2515] = ~(inputs[313]);
    assign layer0_outputs[2516] = inputs[856];
    assign layer0_outputs[2517] = ~((inputs[107]) | (inputs[608]));
    assign layer0_outputs[2518] = (inputs[959]) & (inputs[800]);
    assign layer0_outputs[2519] = ~(inputs[480]) | (inputs[452]);
    assign layer0_outputs[2520] = (inputs[184]) & ~(inputs[358]);
    assign layer0_outputs[2521] = inputs[177];
    assign layer0_outputs[2522] = ~((inputs[47]) ^ (inputs[170]));
    assign layer0_outputs[2523] = (inputs[963]) & ~(inputs[885]);
    assign layer0_outputs[2524] = ~((inputs[383]) & (inputs[642]));
    assign layer0_outputs[2525] = ~((inputs[953]) | (inputs[932]));
    assign layer0_outputs[2526] = (inputs[943]) | (inputs[270]);
    assign layer0_outputs[2527] = 1'b1;
    assign layer0_outputs[2528] = ~((inputs[156]) | (inputs[84]));
    assign layer0_outputs[2529] = inputs[369];
    assign layer0_outputs[2530] = ~(inputs[595]) | (inputs[665]);
    assign layer0_outputs[2531] = (inputs[336]) & ~(inputs[727]);
    assign layer0_outputs[2532] = ~((inputs[473]) ^ (inputs[328]));
    assign layer0_outputs[2533] = 1'b0;
    assign layer0_outputs[2534] = ~(inputs[928]);
    assign layer0_outputs[2535] = (inputs[496]) | (inputs[444]);
    assign layer0_outputs[2536] = (inputs[244]) | (inputs[34]);
    assign layer0_outputs[2537] = 1'b0;
    assign layer0_outputs[2538] = (inputs[38]) ^ (inputs[688]);
    assign layer0_outputs[2539] = (inputs[537]) | (inputs[989]);
    assign layer0_outputs[2540] = ~((inputs[626]) ^ (inputs[984]));
    assign layer0_outputs[2541] = ~((inputs[177]) | (inputs[196]));
    assign layer0_outputs[2542] = inputs[45];
    assign layer0_outputs[2543] = ~((inputs[862]) ^ (inputs[888]));
    assign layer0_outputs[2544] = ~((inputs[444]) & (inputs[865]));
    assign layer0_outputs[2545] = ~(inputs[773]) | (inputs[127]);
    assign layer0_outputs[2546] = ~(inputs[823]) | (inputs[95]);
    assign layer0_outputs[2547] = ~(inputs[569]) | (inputs[596]);
    assign layer0_outputs[2548] = inputs[243];
    assign layer0_outputs[2549] = ~((inputs[612]) & (inputs[829]));
    assign layer0_outputs[2550] = (inputs[303]) & ~(inputs[1010]);
    assign layer0_outputs[2551] = (inputs[954]) | (inputs[284]);
    assign layer0_outputs[2552] = (inputs[396]) & ~(inputs[171]);
    assign layer0_outputs[2553] = ~((inputs[410]) | (inputs[164]));
    assign layer0_outputs[2554] = ~(inputs[315]) | (inputs[704]);
    assign layer0_outputs[2555] = ~(inputs[586]);
    assign layer0_outputs[2556] = inputs[701];
    assign layer0_outputs[2557] = (inputs[728]) | (inputs[571]);
    assign layer0_outputs[2558] = inputs[260];
    assign layer0_outputs[2559] = (inputs[584]) & (inputs[509]);
    assign layer0_outputs[2560] = ~((inputs[586]) ^ (inputs[122]));
    assign layer0_outputs[2561] = inputs[344];
    assign layer0_outputs[2562] = ~((inputs[911]) & (inputs[873]));
    assign layer0_outputs[2563] = (inputs[1010]) & (inputs[187]);
    assign layer0_outputs[2564] = ~(inputs[320]) | (inputs[674]);
    assign layer0_outputs[2565] = inputs[364];
    assign layer0_outputs[2566] = 1'b1;
    assign layer0_outputs[2567] = inputs[715];
    assign layer0_outputs[2568] = ~((inputs[567]) | (inputs[68]));
    assign layer0_outputs[2569] = (inputs[128]) | (inputs[796]);
    assign layer0_outputs[2570] = inputs[106];
    assign layer0_outputs[2571] = ~((inputs[903]) ^ (inputs[612]));
    assign layer0_outputs[2572] = ~(inputs[772]) | (inputs[671]);
    assign layer0_outputs[2573] = (inputs[568]) | (inputs[110]);
    assign layer0_outputs[2574] = (inputs[103]) | (inputs[260]);
    assign layer0_outputs[2575] = (inputs[151]) ^ (inputs[796]);
    assign layer0_outputs[2576] = (inputs[545]) ^ (inputs[570]);
    assign layer0_outputs[2577] = (inputs[1011]) ^ (inputs[552]);
    assign layer0_outputs[2578] = inputs[519];
    assign layer0_outputs[2579] = 1'b0;
    assign layer0_outputs[2580] = ~(inputs[880]) | (inputs[175]);
    assign layer0_outputs[2581] = ~((inputs[729]) ^ (inputs[614]));
    assign layer0_outputs[2582] = (inputs[152]) & ~(inputs[1023]);
    assign layer0_outputs[2583] = ~(inputs[766]) | (inputs[827]);
    assign layer0_outputs[2584] = (inputs[428]) | (inputs[698]);
    assign layer0_outputs[2585] = ~((inputs[203]) ^ (inputs[678]));
    assign layer0_outputs[2586] = (inputs[364]) | (inputs[5]);
    assign layer0_outputs[2587] = inputs[653];
    assign layer0_outputs[2588] = inputs[182];
    assign layer0_outputs[2589] = (inputs[692]) | (inputs[248]);
    assign layer0_outputs[2590] = ~((inputs[702]) ^ (inputs[797]));
    assign layer0_outputs[2591] = ~(inputs[753]) | (inputs[276]);
    assign layer0_outputs[2592] = ~(inputs[567]) | (inputs[827]);
    assign layer0_outputs[2593] = ~(inputs[398]) | (inputs[227]);
    assign layer0_outputs[2594] = ~(inputs[205]);
    assign layer0_outputs[2595] = (inputs[309]) & ~(inputs[137]);
    assign layer0_outputs[2596] = inputs[59];
    assign layer0_outputs[2597] = ~(inputs[250]) | (inputs[672]);
    assign layer0_outputs[2598] = ~(inputs[585]) | (inputs[446]);
    assign layer0_outputs[2599] = ~(inputs[687]);
    assign layer0_outputs[2600] = 1'b1;
    assign layer0_outputs[2601] = (inputs[284]) & ~(inputs[258]);
    assign layer0_outputs[2602] = ~(inputs[623]) | (inputs[130]);
    assign layer0_outputs[2603] = (inputs[7]) ^ (inputs[873]);
    assign layer0_outputs[2604] = (inputs[441]) & ~(inputs[383]);
    assign layer0_outputs[2605] = ~((inputs[608]) ^ (inputs[776]));
    assign layer0_outputs[2606] = (inputs[110]) ^ (inputs[70]);
    assign layer0_outputs[2607] = ~(inputs[143]);
    assign layer0_outputs[2608] = ~((inputs[36]) | (inputs[71]));
    assign layer0_outputs[2609] = ~(inputs[125]);
    assign layer0_outputs[2610] = ~(inputs[87]);
    assign layer0_outputs[2611] = (inputs[28]) & ~(inputs[104]);
    assign layer0_outputs[2612] = ~((inputs[321]) | (inputs[764]));
    assign layer0_outputs[2613] = ~((inputs[732]) | (inputs[381]));
    assign layer0_outputs[2614] = 1'b1;
    assign layer0_outputs[2615] = (inputs[5]) | (inputs[359]);
    assign layer0_outputs[2616] = ~((inputs[1015]) ^ (inputs[636]));
    assign layer0_outputs[2617] = ~(inputs[877]);
    assign layer0_outputs[2618] = ~((inputs[663]) ^ (inputs[596]));
    assign layer0_outputs[2619] = ~(inputs[401]);
    assign layer0_outputs[2620] = 1'b1;
    assign layer0_outputs[2621] = (inputs[383]) | (inputs[171]);
    assign layer0_outputs[2622] = (inputs[606]) ^ (inputs[325]);
    assign layer0_outputs[2623] = ~((inputs[216]) ^ (inputs[576]));
    assign layer0_outputs[2624] = ~(inputs[457]) | (inputs[451]);
    assign layer0_outputs[2625] = (inputs[1012]) ^ (inputs[608]);
    assign layer0_outputs[2626] = ~((inputs[424]) | (inputs[46]));
    assign layer0_outputs[2627] = ~((inputs[234]) | (inputs[299]));
    assign layer0_outputs[2628] = ~(inputs[612]);
    assign layer0_outputs[2629] = (inputs[620]) & ~(inputs[759]);
    assign layer0_outputs[2630] = (inputs[309]) & ~(inputs[434]);
    assign layer0_outputs[2631] = (inputs[365]) & ~(inputs[232]);
    assign layer0_outputs[2632] = ~(inputs[531]);
    assign layer0_outputs[2633] = ~(inputs[459]);
    assign layer0_outputs[2634] = ~(inputs[487]);
    assign layer0_outputs[2635] = (inputs[481]) & (inputs[124]);
    assign layer0_outputs[2636] = (inputs[720]) ^ (inputs[1017]);
    assign layer0_outputs[2637] = ~(inputs[592]) | (inputs[985]);
    assign layer0_outputs[2638] = (inputs[603]) & ~(inputs[87]);
    assign layer0_outputs[2639] = ~(inputs[459]);
    assign layer0_outputs[2640] = ~((inputs[19]) | (inputs[554]));
    assign layer0_outputs[2641] = (inputs[569]) ^ (inputs[630]);
    assign layer0_outputs[2642] = ~((inputs[355]) | (inputs[738]));
    assign layer0_outputs[2643] = inputs[185];
    assign layer0_outputs[2644] = inputs[517];
    assign layer0_outputs[2645] = ~(inputs[328]);
    assign layer0_outputs[2646] = (inputs[375]) & ~(inputs[629]);
    assign layer0_outputs[2647] = (inputs[780]) | (inputs[698]);
    assign layer0_outputs[2648] = ~(inputs[942]);
    assign layer0_outputs[2649] = (inputs[149]) | (inputs[30]);
    assign layer0_outputs[2650] = (inputs[463]) ^ (inputs[804]);
    assign layer0_outputs[2651] = (inputs[157]) & ~(inputs[976]);
    assign layer0_outputs[2652] = inputs[746];
    assign layer0_outputs[2653] = inputs[309];
    assign layer0_outputs[2654] = inputs[784];
    assign layer0_outputs[2655] = (inputs[1000]) & (inputs[197]);
    assign layer0_outputs[2656] = ~((inputs[962]) ^ (inputs[192]));
    assign layer0_outputs[2657] = (inputs[427]) ^ (inputs[577]);
    assign layer0_outputs[2658] = ~((inputs[824]) | (inputs[711]));
    assign layer0_outputs[2659] = 1'b0;
    assign layer0_outputs[2660] = ~((inputs[270]) | (inputs[319]));
    assign layer0_outputs[2661] = (inputs[562]) & ~(inputs[649]);
    assign layer0_outputs[2662] = (inputs[635]) ^ (inputs[504]);
    assign layer0_outputs[2663] = inputs[3];
    assign layer0_outputs[2664] = inputs[149];
    assign layer0_outputs[2665] = ~((inputs[2]) ^ (inputs[754]));
    assign layer0_outputs[2666] = 1'b0;
    assign layer0_outputs[2667] = (inputs[580]) | (inputs[980]);
    assign layer0_outputs[2668] = ~(inputs[412]) | (inputs[833]);
    assign layer0_outputs[2669] = (inputs[629]) & ~(inputs[794]);
    assign layer0_outputs[2670] = ~(inputs[273]);
    assign layer0_outputs[2671] = (inputs[541]) ^ (inputs[823]);
    assign layer0_outputs[2672] = ~(inputs[503]);
    assign layer0_outputs[2673] = (inputs[489]) & ~(inputs[940]);
    assign layer0_outputs[2674] = (inputs[197]) & ~(inputs[104]);
    assign layer0_outputs[2675] = ~(inputs[622]) | (inputs[316]);
    assign layer0_outputs[2676] = ~(inputs[206]);
    assign layer0_outputs[2677] = inputs[402];
    assign layer0_outputs[2678] = ~(inputs[607]);
    assign layer0_outputs[2679] = (inputs[921]) | (inputs[631]);
    assign layer0_outputs[2680] = (inputs[884]) | (inputs[190]);
    assign layer0_outputs[2681] = ~(inputs[587]);
    assign layer0_outputs[2682] = ~((inputs[442]) | (inputs[777]));
    assign layer0_outputs[2683] = (inputs[257]) | (inputs[795]);
    assign layer0_outputs[2684] = (inputs[838]) ^ (inputs[744]);
    assign layer0_outputs[2685] = (inputs[1018]) & ~(inputs[20]);
    assign layer0_outputs[2686] = ~(inputs[24]);
    assign layer0_outputs[2687] = (inputs[827]) | (inputs[698]);
    assign layer0_outputs[2688] = (inputs[212]) & ~(inputs[339]);
    assign layer0_outputs[2689] = (inputs[967]) ^ (inputs[672]);
    assign layer0_outputs[2690] = (inputs[254]) | (inputs[326]);
    assign layer0_outputs[2691] = (inputs[318]) & (inputs[484]);
    assign layer0_outputs[2692] = ~((inputs[558]) & (inputs[715]));
    assign layer0_outputs[2693] = ~(inputs[539]);
    assign layer0_outputs[2694] = ~(inputs[728]);
    assign layer0_outputs[2695] = 1'b0;
    assign layer0_outputs[2696] = ~(inputs[535]) | (inputs[233]);
    assign layer0_outputs[2697] = ~((inputs[717]) | (inputs[174]));
    assign layer0_outputs[2698] = ~(inputs[647]);
    assign layer0_outputs[2699] = ~((inputs[524]) | (inputs[988]));
    assign layer0_outputs[2700] = (inputs[1023]) | (inputs[716]);
    assign layer0_outputs[2701] = 1'b1;
    assign layer0_outputs[2702] = ~(inputs[559]);
    assign layer0_outputs[2703] = (inputs[144]) ^ (inputs[120]);
    assign layer0_outputs[2704] = inputs[149];
    assign layer0_outputs[2705] = inputs[924];
    assign layer0_outputs[2706] = (inputs[86]) & (inputs[671]);
    assign layer0_outputs[2707] = (inputs[305]) & ~(inputs[545]);
    assign layer0_outputs[2708] = inputs[96];
    assign layer0_outputs[2709] = (inputs[532]) & ~(inputs[414]);
    assign layer0_outputs[2710] = (inputs[465]) & ~(inputs[219]);
    assign layer0_outputs[2711] = (inputs[631]) & (inputs[748]);
    assign layer0_outputs[2712] = ~(inputs[436]) | (inputs[91]);
    assign layer0_outputs[2713] = ~(inputs[839]) | (inputs[852]);
    assign layer0_outputs[2714] = ~((inputs[709]) ^ (inputs[714]));
    assign layer0_outputs[2715] = ~(inputs[665]);
    assign layer0_outputs[2716] = ~(inputs[679]);
    assign layer0_outputs[2717] = ~(inputs[509]) | (inputs[1011]);
    assign layer0_outputs[2718] = ~(inputs[536]) | (inputs[874]);
    assign layer0_outputs[2719] = (inputs[765]) | (inputs[205]);
    assign layer0_outputs[2720] = (inputs[739]) | (inputs[676]);
    assign layer0_outputs[2721] = ~((inputs[425]) ^ (inputs[96]));
    assign layer0_outputs[2722] = ~(inputs[554]) | (inputs[637]);
    assign layer0_outputs[2723] = (inputs[822]) | (inputs[794]);
    assign layer0_outputs[2724] = (inputs[676]) | (inputs[551]);
    assign layer0_outputs[2725] = (inputs[757]) | (inputs[699]);
    assign layer0_outputs[2726] = inputs[619];
    assign layer0_outputs[2727] = ~(inputs[70]);
    assign layer0_outputs[2728] = (inputs[470]) & (inputs[258]);
    assign layer0_outputs[2729] = ~(inputs[261]);
    assign layer0_outputs[2730] = ~((inputs[852]) | (inputs[323]));
    assign layer0_outputs[2731] = ~(inputs[457]);
    assign layer0_outputs[2732] = ~(inputs[402]) | (inputs[65]);
    assign layer0_outputs[2733] = ~(inputs[226]) | (inputs[622]);
    assign layer0_outputs[2734] = (inputs[730]) | (inputs[692]);
    assign layer0_outputs[2735] = ~(inputs[701]);
    assign layer0_outputs[2736] = inputs[464];
    assign layer0_outputs[2737] = ~((inputs[189]) | (inputs[553]));
    assign layer0_outputs[2738] = (inputs[790]) & ~(inputs[621]);
    assign layer0_outputs[2739] = (inputs[31]) ^ (inputs[187]);
    assign layer0_outputs[2740] = ~(inputs[177]);
    assign layer0_outputs[2741] = (inputs[987]) & (inputs[75]);
    assign layer0_outputs[2742] = (inputs[439]) & ~(inputs[914]);
    assign layer0_outputs[2743] = ~(inputs[757]) | (inputs[517]);
    assign layer0_outputs[2744] = (inputs[435]) | (inputs[62]);
    assign layer0_outputs[2745] = ~(inputs[811]);
    assign layer0_outputs[2746] = ~(inputs[302]);
    assign layer0_outputs[2747] = ~((inputs[951]) | (inputs[884]));
    assign layer0_outputs[2748] = ~(inputs[832]) | (inputs[452]);
    assign layer0_outputs[2749] = ~(inputs[650]) | (inputs[834]);
    assign layer0_outputs[2750] = (inputs[732]) | (inputs[2]);
    assign layer0_outputs[2751] = ~(inputs[302]) | (inputs[137]);
    assign layer0_outputs[2752] = ~((inputs[65]) | (inputs[613]));
    assign layer0_outputs[2753] = (inputs[265]) & ~(inputs[994]);
    assign layer0_outputs[2754] = ~(inputs[444]);
    assign layer0_outputs[2755] = (inputs[519]) ^ (inputs[969]);
    assign layer0_outputs[2756] = (inputs[16]) ^ (inputs[84]);
    assign layer0_outputs[2757] = 1'b1;
    assign layer0_outputs[2758] = 1'b0;
    assign layer0_outputs[2759] = inputs[473];
    assign layer0_outputs[2760] = ~(inputs[412]);
    assign layer0_outputs[2761] = ~(inputs[717]);
    assign layer0_outputs[2762] = inputs[446];
    assign layer0_outputs[2763] = ~(inputs[971]) | (inputs[153]);
    assign layer0_outputs[2764] = inputs[346];
    assign layer0_outputs[2765] = (inputs[593]) | (inputs[156]);
    assign layer0_outputs[2766] = ~((inputs[276]) | (inputs[859]));
    assign layer0_outputs[2767] = (inputs[619]) & ~(inputs[996]);
    assign layer0_outputs[2768] = ~(inputs[686]);
    assign layer0_outputs[2769] = inputs[749];
    assign layer0_outputs[2770] = (inputs[821]) & ~(inputs[833]);
    assign layer0_outputs[2771] = ~(inputs[213]) | (inputs[544]);
    assign layer0_outputs[2772] = ~(inputs[616]);
    assign layer0_outputs[2773] = (inputs[134]) | (inputs[249]);
    assign layer0_outputs[2774] = inputs[396];
    assign layer0_outputs[2775] = ~(inputs[245]);
    assign layer0_outputs[2776] = (inputs[369]) | (inputs[770]);
    assign layer0_outputs[2777] = (inputs[565]) & ~(inputs[443]);
    assign layer0_outputs[2778] = inputs[503];
    assign layer0_outputs[2779] = (inputs[100]) ^ (inputs[796]);
    assign layer0_outputs[2780] = ~((inputs[571]) | (inputs[195]));
    assign layer0_outputs[2781] = ~((inputs[893]) ^ (inputs[778]));
    assign layer0_outputs[2782] = inputs[887];
    assign layer0_outputs[2783] = inputs[330];
    assign layer0_outputs[2784] = (inputs[359]) | (inputs[227]);
    assign layer0_outputs[2785] = ~(inputs[16]) | (inputs[23]);
    assign layer0_outputs[2786] = ~((inputs[280]) | (inputs[251]));
    assign layer0_outputs[2787] = ~((inputs[285]) | (inputs[215]));
    assign layer0_outputs[2788] = (inputs[850]) ^ (inputs[815]);
    assign layer0_outputs[2789] = (inputs[817]) | (inputs[163]);
    assign layer0_outputs[2790] = ~(inputs[516]) | (inputs[291]);
    assign layer0_outputs[2791] = ~(inputs[427]) | (inputs[130]);
    assign layer0_outputs[2792] = ~(inputs[204]);
    assign layer0_outputs[2793] = inputs[325];
    assign layer0_outputs[2794] = inputs[531];
    assign layer0_outputs[2795] = inputs[760];
    assign layer0_outputs[2796] = (inputs[416]) | (inputs[676]);
    assign layer0_outputs[2797] = inputs[843];
    assign layer0_outputs[2798] = inputs[457];
    assign layer0_outputs[2799] = (inputs[808]) | (inputs[761]);
    assign layer0_outputs[2800] = ~(inputs[871]);
    assign layer0_outputs[2801] = (inputs[354]) & ~(inputs[806]);
    assign layer0_outputs[2802] = ~((inputs[657]) | (inputs[655]));
    assign layer0_outputs[2803] = (inputs[993]) & (inputs[1019]);
    assign layer0_outputs[2804] = (inputs[371]) | (inputs[147]);
    assign layer0_outputs[2805] = ~(inputs[786]) | (inputs[871]);
    assign layer0_outputs[2806] = ~((inputs[734]) | (inputs[3]));
    assign layer0_outputs[2807] = (inputs[49]) | (inputs[340]);
    assign layer0_outputs[2808] = (inputs[79]) | (inputs[591]);
    assign layer0_outputs[2809] = (inputs[273]) & ~(inputs[681]);
    assign layer0_outputs[2810] = (inputs[756]) & ~(inputs[538]);
    assign layer0_outputs[2811] = inputs[857];
    assign layer0_outputs[2812] = inputs[784];
    assign layer0_outputs[2813] = 1'b1;
    assign layer0_outputs[2814] = (inputs[149]) & ~(inputs[741]);
    assign layer0_outputs[2815] = (inputs[765]) & (inputs[319]);
    assign layer0_outputs[2816] = ~((inputs[63]) ^ (inputs[476]));
    assign layer0_outputs[2817] = (inputs[352]) & (inputs[979]);
    assign layer0_outputs[2818] = ~(inputs[762]) | (inputs[79]);
    assign layer0_outputs[2819] = inputs[936];
    assign layer0_outputs[2820] = ~((inputs[27]) ^ (inputs[436]));
    assign layer0_outputs[2821] = (inputs[200]) ^ (inputs[719]);
    assign layer0_outputs[2822] = (inputs[170]) & ~(inputs[674]);
    assign layer0_outputs[2823] = (inputs[65]) ^ (inputs[436]);
    assign layer0_outputs[2824] = (inputs[782]) | (inputs[218]);
    assign layer0_outputs[2825] = inputs[43];
    assign layer0_outputs[2826] = inputs[142];
    assign layer0_outputs[2827] = (inputs[896]) ^ (inputs[106]);
    assign layer0_outputs[2828] = (inputs[446]) | (inputs[432]);
    assign layer0_outputs[2829] = ~(inputs[2]);
    assign layer0_outputs[2830] = (inputs[617]) & ~(inputs[814]);
    assign layer0_outputs[2831] = ~((inputs[828]) ^ (inputs[907]));
    assign layer0_outputs[2832] = (inputs[504]) & ~(inputs[355]);
    assign layer0_outputs[2833] = ~((inputs[174]) | (inputs[84]));
    assign layer0_outputs[2834] = (inputs[50]) & ~(inputs[117]);
    assign layer0_outputs[2835] = (inputs[738]) | (inputs[685]);
    assign layer0_outputs[2836] = (inputs[834]) & ~(inputs[804]);
    assign layer0_outputs[2837] = (inputs[334]) ^ (inputs[226]);
    assign layer0_outputs[2838] = inputs[642];
    assign layer0_outputs[2839] = (inputs[723]) & ~(inputs[572]);
    assign layer0_outputs[2840] = (inputs[565]) | (inputs[80]);
    assign layer0_outputs[2841] = (inputs[364]) & ~(inputs[33]);
    assign layer0_outputs[2842] = (inputs[392]) ^ (inputs[510]);
    assign layer0_outputs[2843] = (inputs[524]) ^ (inputs[999]);
    assign layer0_outputs[2844] = (inputs[469]) & ~(inputs[849]);
    assign layer0_outputs[2845] = ~(inputs[287]) | (inputs[129]);
    assign layer0_outputs[2846] = ~((inputs[371]) | (inputs[852]));
    assign layer0_outputs[2847] = ~((inputs[738]) ^ (inputs[349]));
    assign layer0_outputs[2848] = inputs[371];
    assign layer0_outputs[2849] = 1'b1;
    assign layer0_outputs[2850] = (inputs[536]) | (inputs[228]);
    assign layer0_outputs[2851] = (inputs[295]) | (inputs[515]);
    assign layer0_outputs[2852] = ~(inputs[602]) | (inputs[130]);
    assign layer0_outputs[2853] = ~(inputs[441]);
    assign layer0_outputs[2854] = ~((inputs[79]) ^ (inputs[167]));
    assign layer0_outputs[2855] = ~(inputs[131]) | (inputs[124]);
    assign layer0_outputs[2856] = (inputs[623]) | (inputs[557]);
    assign layer0_outputs[2857] = 1'b0;
    assign layer0_outputs[2858] = (inputs[378]) | (inputs[160]);
    assign layer0_outputs[2859] = inputs[1005];
    assign layer0_outputs[2860] = (inputs[897]) | (inputs[528]);
    assign layer0_outputs[2861] = inputs[685];
    assign layer0_outputs[2862] = (inputs[328]) & ~(inputs[959]);
    assign layer0_outputs[2863] = 1'b1;
    assign layer0_outputs[2864] = ~((inputs[755]) | (inputs[179]));
    assign layer0_outputs[2865] = ~((inputs[961]) | (inputs[328]));
    assign layer0_outputs[2866] = ~((inputs[342]) ^ (inputs[348]));
    assign layer0_outputs[2867] = (inputs[33]) & ~(inputs[576]);
    assign layer0_outputs[2868] = (inputs[23]) & ~(inputs[542]);
    assign layer0_outputs[2869] = 1'b1;
    assign layer0_outputs[2870] = ~(inputs[804]);
    assign layer0_outputs[2871] = ~(inputs[120]) | (inputs[352]);
    assign layer0_outputs[2872] = ~(inputs[360]);
    assign layer0_outputs[2873] = ~(inputs[760]) | (inputs[71]);
    assign layer0_outputs[2874] = (inputs[751]) & ~(inputs[175]);
    assign layer0_outputs[2875] = (inputs[826]) ^ (inputs[693]);
    assign layer0_outputs[2876] = ~(inputs[771]);
    assign layer0_outputs[2877] = ~(inputs[1000]);
    assign layer0_outputs[2878] = (inputs[769]) & ~(inputs[650]);
    assign layer0_outputs[2879] = (inputs[837]) | (inputs[809]);
    assign layer0_outputs[2880] = ~(inputs[242]) | (inputs[894]);
    assign layer0_outputs[2881] = (inputs[164]) & ~(inputs[155]);
    assign layer0_outputs[2882] = (inputs[23]) | (inputs[625]);
    assign layer0_outputs[2883] = (inputs[301]) | (inputs[923]);
    assign layer0_outputs[2884] = ~(inputs[816]);
    assign layer0_outputs[2885] = ~(inputs[934]);
    assign layer0_outputs[2886] = ~((inputs[440]) & (inputs[289]));
    assign layer0_outputs[2887] = (inputs[284]) | (inputs[236]);
    assign layer0_outputs[2888] = ~(inputs[642]) | (inputs[72]);
    assign layer0_outputs[2889] = ~(inputs[234]);
    assign layer0_outputs[2890] = ~((inputs[211]) | (inputs[745]));
    assign layer0_outputs[2891] = inputs[193];
    assign layer0_outputs[2892] = 1'b1;
    assign layer0_outputs[2893] = 1'b1;
    assign layer0_outputs[2894] = ~(inputs[624]) | (inputs[839]);
    assign layer0_outputs[2895] = ~(inputs[72]) | (inputs[209]);
    assign layer0_outputs[2896] = (inputs[925]) & ~(inputs[232]);
    assign layer0_outputs[2897] = (inputs[75]) | (inputs[904]);
    assign layer0_outputs[2898] = inputs[498];
    assign layer0_outputs[2899] = ~(inputs[309]);
    assign layer0_outputs[2900] = (inputs[551]) ^ (inputs[643]);
    assign layer0_outputs[2901] = (inputs[845]) | (inputs[417]);
    assign layer0_outputs[2902] = (inputs[262]) | (inputs[349]);
    assign layer0_outputs[2903] = ~((inputs[13]) | (inputs[64]));
    assign layer0_outputs[2904] = ~(inputs[616]) | (inputs[942]);
    assign layer0_outputs[2905] = (inputs[344]) | (inputs[933]);
    assign layer0_outputs[2906] = ~(inputs[168]) | (inputs[163]);
    assign layer0_outputs[2907] = ~(inputs[376]);
    assign layer0_outputs[2908] = inputs[300];
    assign layer0_outputs[2909] = ~(inputs[977]);
    assign layer0_outputs[2910] = ~(inputs[590]);
    assign layer0_outputs[2911] = (inputs[552]) & ~(inputs[163]);
    assign layer0_outputs[2912] = (inputs[522]) | (inputs[412]);
    assign layer0_outputs[2913] = inputs[554];
    assign layer0_outputs[2914] = ~((inputs[720]) ^ (inputs[292]));
    assign layer0_outputs[2915] = ~((inputs[248]) | (inputs[645]));
    assign layer0_outputs[2916] = ~((inputs[1018]) & (inputs[1021]));
    assign layer0_outputs[2917] = (inputs[366]) | (inputs[387]);
    assign layer0_outputs[2918] = inputs[334];
    assign layer0_outputs[2919] = (inputs[827]) | (inputs[882]);
    assign layer0_outputs[2920] = (inputs[699]) ^ (inputs[744]);
    assign layer0_outputs[2921] = (inputs[901]) | (inputs[562]);
    assign layer0_outputs[2922] = ~((inputs[1007]) ^ (inputs[216]));
    assign layer0_outputs[2923] = (inputs[1004]) & (inputs[828]);
    assign layer0_outputs[2924] = (inputs[1018]) & ~(inputs[28]);
    assign layer0_outputs[2925] = (inputs[54]) & ~(inputs[642]);
    assign layer0_outputs[2926] = (inputs[792]) ^ (inputs[147]);
    assign layer0_outputs[2927] = (inputs[381]) ^ (inputs[406]);
    assign layer0_outputs[2928] = ~((inputs[78]) | (inputs[123]));
    assign layer0_outputs[2929] = ~(inputs[528]);
    assign layer0_outputs[2930] = ~(inputs[920]) | (inputs[256]);
    assign layer0_outputs[2931] = ~(inputs[692]) | (inputs[859]);
    assign layer0_outputs[2932] = (inputs[85]) | (inputs[191]);
    assign layer0_outputs[2933] = 1'b0;
    assign layer0_outputs[2934] = (inputs[395]) & ~(inputs[795]);
    assign layer0_outputs[2935] = inputs[490];
    assign layer0_outputs[2936] = ~(inputs[566]);
    assign layer0_outputs[2937] = (inputs[72]) & ~(inputs[131]);
    assign layer0_outputs[2938] = (inputs[833]) & ~(inputs[897]);
    assign layer0_outputs[2939] = ~((inputs[923]) | (inputs[916]));
    assign layer0_outputs[2940] = ~(inputs[538]);
    assign layer0_outputs[2941] = 1'b0;
    assign layer0_outputs[2942] = (inputs[251]) & ~(inputs[963]);
    assign layer0_outputs[2943] = ~(inputs[808]) | (inputs[315]);
    assign layer0_outputs[2944] = 1'b1;
    assign layer0_outputs[2945] = ~(inputs[789]) | (inputs[800]);
    assign layer0_outputs[2946] = ~((inputs[792]) | (inputs[858]));
    assign layer0_outputs[2947] = 1'b1;
    assign layer0_outputs[2948] = ~((inputs[94]) ^ (inputs[600]));
    assign layer0_outputs[2949] = inputs[335];
    assign layer0_outputs[2950] = ~(inputs[53]);
    assign layer0_outputs[2951] = (inputs[783]) & (inputs[470]);
    assign layer0_outputs[2952] = ~((inputs[957]) | (inputs[372]));
    assign layer0_outputs[2953] = ~(inputs[498]) | (inputs[382]);
    assign layer0_outputs[2954] = ~((inputs[486]) & (inputs[11]));
    assign layer0_outputs[2955] = 1'b0;
    assign layer0_outputs[2956] = ~((inputs[796]) ^ (inputs[343]));
    assign layer0_outputs[2957] = ~((inputs[204]) | (inputs[725]));
    assign layer0_outputs[2958] = (inputs[35]) & ~(inputs[395]);
    assign layer0_outputs[2959] = ~(inputs[780]) | (inputs[487]);
    assign layer0_outputs[2960] = (inputs[205]) | (inputs[727]);
    assign layer0_outputs[2961] = (inputs[354]) | (inputs[875]);
    assign layer0_outputs[2962] = ~((inputs[259]) | (inputs[340]));
    assign layer0_outputs[2963] = (inputs[117]) ^ (inputs[286]);
    assign layer0_outputs[2964] = (inputs[731]) & (inputs[35]);
    assign layer0_outputs[2965] = (inputs[462]) & ~(inputs[443]);
    assign layer0_outputs[2966] = ~((inputs[755]) | (inputs[873]));
    assign layer0_outputs[2967] = ~(inputs[718]);
    assign layer0_outputs[2968] = (inputs[968]) | (inputs[546]);
    assign layer0_outputs[2969] = ~(inputs[214]) | (inputs[139]);
    assign layer0_outputs[2970] = (inputs[354]) & ~(inputs[994]);
    assign layer0_outputs[2971] = ~(inputs[426]);
    assign layer0_outputs[2972] = (inputs[405]) & ~(inputs[480]);
    assign layer0_outputs[2973] = ~(inputs[567]);
    assign layer0_outputs[2974] = ~((inputs[223]) | (inputs[24]));
    assign layer0_outputs[2975] = (inputs[902]) | (inputs[327]);
    assign layer0_outputs[2976] = (inputs[531]) & ~(inputs[46]);
    assign layer0_outputs[2977] = (inputs[346]) ^ (inputs[605]);
    assign layer0_outputs[2978] = ~((inputs[80]) & (inputs[466]));
    assign layer0_outputs[2979] = (inputs[380]) & ~(inputs[904]);
    assign layer0_outputs[2980] = 1'b1;
    assign layer0_outputs[2981] = ~((inputs[26]) | (inputs[594]));
    assign layer0_outputs[2982] = ~((inputs[687]) | (inputs[756]));
    assign layer0_outputs[2983] = ~(inputs[791]);
    assign layer0_outputs[2984] = ~((inputs[902]) ^ (inputs[281]));
    assign layer0_outputs[2985] = inputs[895];
    assign layer0_outputs[2986] = ~((inputs[650]) | (inputs[759]));
    assign layer0_outputs[2987] = (inputs[760]) & ~(inputs[101]);
    assign layer0_outputs[2988] = (inputs[84]) & (inputs[727]);
    assign layer0_outputs[2989] = (inputs[906]) & ~(inputs[149]);
    assign layer0_outputs[2990] = ~((inputs[250]) & (inputs[484]));
    assign layer0_outputs[2991] = ~(inputs[594]) | (inputs[101]);
    assign layer0_outputs[2992] = (inputs[468]) | (inputs[1006]);
    assign layer0_outputs[2993] = 1'b1;
    assign layer0_outputs[2994] = ~((inputs[388]) ^ (inputs[201]));
    assign layer0_outputs[2995] = ~(inputs[238]);
    assign layer0_outputs[2996] = (inputs[967]) | (inputs[465]);
    assign layer0_outputs[2997] = ~((inputs[766]) & (inputs[423]));
    assign layer0_outputs[2998] = (inputs[404]) & ~(inputs[158]);
    assign layer0_outputs[2999] = (inputs[953]) & ~(inputs[700]);
    assign layer0_outputs[3000] = ~((inputs[660]) ^ (inputs[132]));
    assign layer0_outputs[3001] = ~(inputs[528]);
    assign layer0_outputs[3002] = (inputs[7]) | (inputs[616]);
    assign layer0_outputs[3003] = (inputs[758]) ^ (inputs[623]);
    assign layer0_outputs[3004] = ~(inputs[546]) | (inputs[189]);
    assign layer0_outputs[3005] = ~((inputs[750]) ^ (inputs[367]));
    assign layer0_outputs[3006] = ~(inputs[309]) | (inputs[660]);
    assign layer0_outputs[3007] = ~(inputs[721]);
    assign layer0_outputs[3008] = ~((inputs[295]) | (inputs[906]));
    assign layer0_outputs[3009] = ~((inputs[159]) ^ (inputs[607]));
    assign layer0_outputs[3010] = (inputs[470]) & ~(inputs[448]);
    assign layer0_outputs[3011] = (inputs[161]) | (inputs[184]);
    assign layer0_outputs[3012] = ~((inputs[934]) | (inputs[268]));
    assign layer0_outputs[3013] = (inputs[922]) | (inputs[697]);
    assign layer0_outputs[3014] = ~((inputs[963]) | (inputs[881]));
    assign layer0_outputs[3015] = (inputs[447]) & ~(inputs[73]);
    assign layer0_outputs[3016] = (inputs[526]) & ~(inputs[197]);
    assign layer0_outputs[3017] = ~(inputs[178]) | (inputs[834]);
    assign layer0_outputs[3018] = ~(inputs[811]) | (inputs[1008]);
    assign layer0_outputs[3019] = inputs[808];
    assign layer0_outputs[3020] = ~((inputs[329]) | (inputs[193]));
    assign layer0_outputs[3021] = (inputs[198]) & ~(inputs[56]);
    assign layer0_outputs[3022] = ~(inputs[881]) | (inputs[142]);
    assign layer0_outputs[3023] = ~((inputs[995]) & (inputs[1005]));
    assign layer0_outputs[3024] = (inputs[8]) | (inputs[163]);
    assign layer0_outputs[3025] = (inputs[371]) ^ (inputs[247]);
    assign layer0_outputs[3026] = (inputs[609]) | (inputs[50]);
    assign layer0_outputs[3027] = 1'b1;
    assign layer0_outputs[3028] = (inputs[744]) & ~(inputs[930]);
    assign layer0_outputs[3029] = (inputs[823]) ^ (inputs[225]);
    assign layer0_outputs[3030] = ~((inputs[185]) ^ (inputs[448]));
    assign layer0_outputs[3031] = ~((inputs[892]) ^ (inputs[938]));
    assign layer0_outputs[3032] = inputs[23];
    assign layer0_outputs[3033] = (inputs[436]) ^ (inputs[642]);
    assign layer0_outputs[3034] = (inputs[908]) & ~(inputs[191]);
    assign layer0_outputs[3035] = ~(inputs[363]);
    assign layer0_outputs[3036] = ~((inputs[507]) ^ (inputs[219]));
    assign layer0_outputs[3037] = ~(inputs[333]) | (inputs[1009]);
    assign layer0_outputs[3038] = ~((inputs[185]) ^ (inputs[228]));
    assign layer0_outputs[3039] = ~(inputs[154]);
    assign layer0_outputs[3040] = (inputs[716]) | (inputs[727]);
    assign layer0_outputs[3041] = (inputs[49]) | (inputs[776]);
    assign layer0_outputs[3042] = inputs[623];
    assign layer0_outputs[3043] = ~(inputs[181]);
    assign layer0_outputs[3044] = (inputs[122]) ^ (inputs[249]);
    assign layer0_outputs[3045] = ~((inputs[883]) | (inputs[619]));
    assign layer0_outputs[3046] = (inputs[917]) | (inputs[927]);
    assign layer0_outputs[3047] = (inputs[645]) | (inputs[826]);
    assign layer0_outputs[3048] = inputs[362];
    assign layer0_outputs[3049] = ~((inputs[636]) | (inputs[171]));
    assign layer0_outputs[3050] = inputs[131];
    assign layer0_outputs[3051] = ~(inputs[928]);
    assign layer0_outputs[3052] = ~(inputs[745]);
    assign layer0_outputs[3053] = inputs[520];
    assign layer0_outputs[3054] = (inputs[956]) ^ (inputs[560]);
    assign layer0_outputs[3055] = (inputs[377]) | (inputs[825]);
    assign layer0_outputs[3056] = ~((inputs[653]) | (inputs[1009]));
    assign layer0_outputs[3057] = inputs[615];
    assign layer0_outputs[3058] = (inputs[85]) | (inputs[506]);
    assign layer0_outputs[3059] = (inputs[730]) | (inputs[386]);
    assign layer0_outputs[3060] = ~(inputs[785]);
    assign layer0_outputs[3061] = ~((inputs[732]) ^ (inputs[758]));
    assign layer0_outputs[3062] = ~((inputs[1002]) | (inputs[950]));
    assign layer0_outputs[3063] = inputs[78];
    assign layer0_outputs[3064] = (inputs[144]) | (inputs[728]);
    assign layer0_outputs[3065] = (inputs[654]) & ~(inputs[940]);
    assign layer0_outputs[3066] = ~(inputs[208]);
    assign layer0_outputs[3067] = (inputs[609]) ^ (inputs[182]);
    assign layer0_outputs[3068] = (inputs[826]) & ~(inputs[252]);
    assign layer0_outputs[3069] = (inputs[552]) & ~(inputs[191]);
    assign layer0_outputs[3070] = ~((inputs[499]) | (inputs[441]));
    assign layer0_outputs[3071] = ~(inputs[720]) | (inputs[483]);
    assign layer0_outputs[3072] = ~(inputs[43]);
    assign layer0_outputs[3073] = (inputs[959]) & ~(inputs[64]);
    assign layer0_outputs[3074] = (inputs[588]) & ~(inputs[250]);
    assign layer0_outputs[3075] = ~((inputs[121]) & (inputs[208]));
    assign layer0_outputs[3076] = (inputs[408]) ^ (inputs[448]);
    assign layer0_outputs[3077] = (inputs[814]) & ~(inputs[508]);
    assign layer0_outputs[3078] = inputs[785];
    assign layer0_outputs[3079] = ~((inputs[119]) ^ (inputs[598]));
    assign layer0_outputs[3080] = inputs[417];
    assign layer0_outputs[3081] = inputs[664];
    assign layer0_outputs[3082] = ~((inputs[648]) | (inputs[170]));
    assign layer0_outputs[3083] = (inputs[742]) ^ (inputs[2]);
    assign layer0_outputs[3084] = ~(inputs[553]) | (inputs[769]);
    assign layer0_outputs[3085] = inputs[298];
    assign layer0_outputs[3086] = (inputs[890]) & ~(inputs[955]);
    assign layer0_outputs[3087] = (inputs[181]) ^ (inputs[1004]);
    assign layer0_outputs[3088] = ~(inputs[417]);
    assign layer0_outputs[3089] = ~(inputs[265]) | (inputs[154]);
    assign layer0_outputs[3090] = ~(inputs[332]);
    assign layer0_outputs[3091] = inputs[644];
    assign layer0_outputs[3092] = inputs[586];
    assign layer0_outputs[3093] = (inputs[172]) & ~(inputs[128]);
    assign layer0_outputs[3094] = (inputs[822]) & ~(inputs[987]);
    assign layer0_outputs[3095] = (inputs[924]) | (inputs[256]);
    assign layer0_outputs[3096] = (inputs[84]) ^ (inputs[1005]);
    assign layer0_outputs[3097] = ~(inputs[146]);
    assign layer0_outputs[3098] = inputs[148];
    assign layer0_outputs[3099] = inputs[661];
    assign layer0_outputs[3100] = inputs[135];
    assign layer0_outputs[3101] = (inputs[596]) | (inputs[510]);
    assign layer0_outputs[3102] = ~((inputs[297]) | (inputs[242]));
    assign layer0_outputs[3103] = ~(inputs[469]) | (inputs[111]);
    assign layer0_outputs[3104] = (inputs[443]) | (inputs[684]);
    assign layer0_outputs[3105] = 1'b1;
    assign layer0_outputs[3106] = ~((inputs[984]) | (inputs[558]));
    assign layer0_outputs[3107] = ~(inputs[1022]);
    assign layer0_outputs[3108] = (inputs[842]) | (inputs[317]);
    assign layer0_outputs[3109] = ~((inputs[1007]) | (inputs[541]));
    assign layer0_outputs[3110] = 1'b1;
    assign layer0_outputs[3111] = (inputs[318]) | (inputs[571]);
    assign layer0_outputs[3112] = ~(inputs[1018]);
    assign layer0_outputs[3113] = ~(inputs[936]);
    assign layer0_outputs[3114] = inputs[442];
    assign layer0_outputs[3115] = ~(inputs[501]) | (inputs[13]);
    assign layer0_outputs[3116] = ~(inputs[623]) | (inputs[120]);
    assign layer0_outputs[3117] = ~((inputs[733]) | (inputs[275]));
    assign layer0_outputs[3118] = ~((inputs[377]) | (inputs[389]));
    assign layer0_outputs[3119] = (inputs[485]) | (inputs[239]);
    assign layer0_outputs[3120] = (inputs[697]) ^ (inputs[442]);
    assign layer0_outputs[3121] = ~(inputs[362]) | (inputs[14]);
    assign layer0_outputs[3122] = ~((inputs[875]) | (inputs[285]));
    assign layer0_outputs[3123] = ~(inputs[340]) | (inputs[550]);
    assign layer0_outputs[3124] = ~((inputs[405]) & (inputs[756]));
    assign layer0_outputs[3125] = (inputs[993]) & ~(inputs[962]);
    assign layer0_outputs[3126] = ~(inputs[188]) | (inputs[412]);
    assign layer0_outputs[3127] = ~((inputs[681]) ^ (inputs[928]));
    assign layer0_outputs[3128] = ~((inputs[855]) ^ (inputs[158]));
    assign layer0_outputs[3129] = ~(inputs[209]);
    assign layer0_outputs[3130] = ~((inputs[5]) | (inputs[855]));
    assign layer0_outputs[3131] = inputs[946];
    assign layer0_outputs[3132] = (inputs[868]) ^ (inputs[226]);
    assign layer0_outputs[3133] = (inputs[534]) & ~(inputs[837]);
    assign layer0_outputs[3134] = ~(inputs[307]);
    assign layer0_outputs[3135] = ~((inputs[14]) ^ (inputs[644]));
    assign layer0_outputs[3136] = (inputs[318]) & ~(inputs[158]);
    assign layer0_outputs[3137] = (inputs[669]) & ~(inputs[83]);
    assign layer0_outputs[3138] = ~(inputs[819]) | (inputs[119]);
    assign layer0_outputs[3139] = ~(inputs[628]);
    assign layer0_outputs[3140] = (inputs[213]) | (inputs[636]);
    assign layer0_outputs[3141] = ~((inputs[766]) ^ (inputs[826]));
    assign layer0_outputs[3142] = ~((inputs[254]) | (inputs[871]));
    assign layer0_outputs[3143] = ~(inputs[763]);
    assign layer0_outputs[3144] = ~((inputs[120]) ^ (inputs[167]));
    assign layer0_outputs[3145] = 1'b1;
    assign layer0_outputs[3146] = (inputs[464]) & ~(inputs[414]);
    assign layer0_outputs[3147] = (inputs[667]) & ~(inputs[830]);
    assign layer0_outputs[3148] = (inputs[93]) ^ (inputs[745]);
    assign layer0_outputs[3149] = inputs[191];
    assign layer0_outputs[3150] = (inputs[449]) ^ (inputs[900]);
    assign layer0_outputs[3151] = ~((inputs[545]) ^ (inputs[889]));
    assign layer0_outputs[3152] = (inputs[863]) ^ (inputs[683]);
    assign layer0_outputs[3153] = 1'b0;
    assign layer0_outputs[3154] = ~((inputs[501]) | (inputs[512]));
    assign layer0_outputs[3155] = ~((inputs[319]) & (inputs[751]));
    assign layer0_outputs[3156] = (inputs[857]) | (inputs[690]);
    assign layer0_outputs[3157] = ~(inputs[473]);
    assign layer0_outputs[3158] = inputs[221];
    assign layer0_outputs[3159] = ~((inputs[718]) | (inputs[82]));
    assign layer0_outputs[3160] = ~(inputs[592]) | (inputs[15]);
    assign layer0_outputs[3161] = (inputs[795]) | (inputs[377]);
    assign layer0_outputs[3162] = (inputs[369]) | (inputs[764]);
    assign layer0_outputs[3163] = ~((inputs[618]) ^ (inputs[93]));
    assign layer0_outputs[3164] = (inputs[873]) & ~(inputs[220]);
    assign layer0_outputs[3165] = (inputs[829]) & (inputs[115]);
    assign layer0_outputs[3166] = ~((inputs[493]) ^ (inputs[606]));
    assign layer0_outputs[3167] = ~((inputs[444]) ^ (inputs[450]));
    assign layer0_outputs[3168] = ~(inputs[694]) | (inputs[433]);
    assign layer0_outputs[3169] = inputs[623];
    assign layer0_outputs[3170] = (inputs[747]) & ~(inputs[623]);
    assign layer0_outputs[3171] = (inputs[610]) & ~(inputs[674]);
    assign layer0_outputs[3172] = (inputs[466]) & ~(inputs[846]);
    assign layer0_outputs[3173] = ~((inputs[110]) ^ (inputs[0]));
    assign layer0_outputs[3174] = 1'b1;
    assign layer0_outputs[3175] = (inputs[635]) | (inputs[723]);
    assign layer0_outputs[3176] = inputs[110];
    assign layer0_outputs[3177] = inputs[430];
    assign layer0_outputs[3178] = (inputs[117]) & (inputs[944]);
    assign layer0_outputs[3179] = inputs[724];
    assign layer0_outputs[3180] = inputs[333];
    assign layer0_outputs[3181] = (inputs[521]) & ~(inputs[43]);
    assign layer0_outputs[3182] = ~((inputs[650]) | (inputs[627]));
    assign layer0_outputs[3183] = ~(inputs[756]) | (inputs[990]);
    assign layer0_outputs[3184] = (inputs[790]) & ~(inputs[104]);
    assign layer0_outputs[3185] = inputs[757];
    assign layer0_outputs[3186] = (inputs[16]) | (inputs[407]);
    assign layer0_outputs[3187] = ~(inputs[614]) | (inputs[13]);
    assign layer0_outputs[3188] = 1'b0;
    assign layer0_outputs[3189] = inputs[684];
    assign layer0_outputs[3190] = (inputs[983]) | (inputs[204]);
    assign layer0_outputs[3191] = (inputs[89]) & (inputs[581]);
    assign layer0_outputs[3192] = ~((inputs[216]) ^ (inputs[1008]));
    assign layer0_outputs[3193] = ~(inputs[313]);
    assign layer0_outputs[3194] = inputs[315];
    assign layer0_outputs[3195] = ~((inputs[282]) | (inputs[856]));
    assign layer0_outputs[3196] = inputs[233];
    assign layer0_outputs[3197] = ~((inputs[426]) ^ (inputs[335]));
    assign layer0_outputs[3198] = ~((inputs[346]) | (inputs[622]));
    assign layer0_outputs[3199] = ~(inputs[973]) | (inputs[672]);
    assign layer0_outputs[3200] = ~(inputs[526]);
    assign layer0_outputs[3201] = inputs[615];
    assign layer0_outputs[3202] = ~(inputs[888]) | (inputs[73]);
    assign layer0_outputs[3203] = ~((inputs[760]) | (inputs[618]));
    assign layer0_outputs[3204] = (inputs[72]) & (inputs[330]);
    assign layer0_outputs[3205] = (inputs[668]) & (inputs[798]);
    assign layer0_outputs[3206] = (inputs[564]) & ~(inputs[899]);
    assign layer0_outputs[3207] = (inputs[233]) & ~(inputs[106]);
    assign layer0_outputs[3208] = ~((inputs[1007]) & (inputs[482]));
    assign layer0_outputs[3209] = ~(inputs[235]);
    assign layer0_outputs[3210] = 1'b1;
    assign layer0_outputs[3211] = (inputs[10]) | (inputs[319]);
    assign layer0_outputs[3212] = inputs[23];
    assign layer0_outputs[3213] = inputs[1006];
    assign layer0_outputs[3214] = inputs[274];
    assign layer0_outputs[3215] = (inputs[739]) ^ (inputs[1015]);
    assign layer0_outputs[3216] = ~(inputs[558]);
    assign layer0_outputs[3217] = (inputs[210]) | (inputs[812]);
    assign layer0_outputs[3218] = ~(inputs[728]);
    assign layer0_outputs[3219] = (inputs[388]) & ~(inputs[706]);
    assign layer0_outputs[3220] = 1'b1;
    assign layer0_outputs[3221] = inputs[496];
    assign layer0_outputs[3222] = (inputs[689]) | (inputs[160]);
    assign layer0_outputs[3223] = ~(inputs[946]);
    assign layer0_outputs[3224] = ~(inputs[789]) | (inputs[160]);
    assign layer0_outputs[3225] = (inputs[184]) & ~(inputs[850]);
    assign layer0_outputs[3226] = 1'b1;
    assign layer0_outputs[3227] = ~((inputs[367]) | (inputs[384]));
    assign layer0_outputs[3228] = (inputs[553]) & ~(inputs[994]);
    assign layer0_outputs[3229] = ~(inputs[593]) | (inputs[890]);
    assign layer0_outputs[3230] = (inputs[331]) & ~(inputs[727]);
    assign layer0_outputs[3231] = inputs[301];
    assign layer0_outputs[3232] = ~((inputs[438]) | (inputs[223]));
    assign layer0_outputs[3233] = ~((inputs[933]) & (inputs[848]));
    assign layer0_outputs[3234] = (inputs[656]) & ~(inputs[608]);
    assign layer0_outputs[3235] = (inputs[421]) | (inputs[594]);
    assign layer0_outputs[3236] = (inputs[468]) | (inputs[598]);
    assign layer0_outputs[3237] = ~(inputs[113]);
    assign layer0_outputs[3238] = ~(inputs[274]);
    assign layer0_outputs[3239] = (inputs[551]) | (inputs[1021]);
    assign layer0_outputs[3240] = ~(inputs[408]) | (inputs[539]);
    assign layer0_outputs[3241] = ~((inputs[790]) ^ (inputs[609]));
    assign layer0_outputs[3242] = (inputs[25]) ^ (inputs[493]);
    assign layer0_outputs[3243] = (inputs[957]) ^ (inputs[813]);
    assign layer0_outputs[3244] = ~((inputs[44]) | (inputs[188]));
    assign layer0_outputs[3245] = (inputs[966]) & ~(inputs[111]);
    assign layer0_outputs[3246] = (inputs[554]) | (inputs[194]);
    assign layer0_outputs[3247] = ~(inputs[73]);
    assign layer0_outputs[3248] = 1'b1;
    assign layer0_outputs[3249] = (inputs[154]) | (inputs[131]);
    assign layer0_outputs[3250] = ~(inputs[155]);
    assign layer0_outputs[3251] = ~((inputs[113]) | (inputs[718]));
    assign layer0_outputs[3252] = ~((inputs[356]) & (inputs[517]));
    assign layer0_outputs[3253] = (inputs[901]) ^ (inputs[559]);
    assign layer0_outputs[3254] = ~((inputs[333]) ^ (inputs[102]));
    assign layer0_outputs[3255] = ~(inputs[907]);
    assign layer0_outputs[3256] = 1'b0;
    assign layer0_outputs[3257] = ~(inputs[655]) | (inputs[924]);
    assign layer0_outputs[3258] = (inputs[490]) & ~(inputs[408]);
    assign layer0_outputs[3259] = (inputs[555]) & ~(inputs[12]);
    assign layer0_outputs[3260] = ~(inputs[440]);
    assign layer0_outputs[3261] = ~((inputs[88]) ^ (inputs[76]));
    assign layer0_outputs[3262] = ~((inputs[173]) | (inputs[825]));
    assign layer0_outputs[3263] = ~(inputs[274]);
    assign layer0_outputs[3264] = ~(inputs[398]) | (inputs[1019]);
    assign layer0_outputs[3265] = (inputs[392]) | (inputs[269]);
    assign layer0_outputs[3266] = ~((inputs[740]) | (inputs[678]));
    assign layer0_outputs[3267] = ~((inputs[897]) & (inputs[383]));
    assign layer0_outputs[3268] = 1'b0;
    assign layer0_outputs[3269] = (inputs[285]) | (inputs[913]);
    assign layer0_outputs[3270] = (inputs[924]) ^ (inputs[767]);
    assign layer0_outputs[3271] = ~(inputs[529]) | (inputs[871]);
    assign layer0_outputs[3272] = ~((inputs[506]) ^ (inputs[916]));
    assign layer0_outputs[3273] = (inputs[431]) | (inputs[904]);
    assign layer0_outputs[3274] = (inputs[520]) ^ (inputs[287]);
    assign layer0_outputs[3275] = 1'b1;
    assign layer0_outputs[3276] = ~(inputs[680]) | (inputs[986]);
    assign layer0_outputs[3277] = 1'b1;
    assign layer0_outputs[3278] = ~(inputs[860]) | (inputs[573]);
    assign layer0_outputs[3279] = ~(inputs[626]) | (inputs[381]);
    assign layer0_outputs[3280] = (inputs[855]) & ~(inputs[898]);
    assign layer0_outputs[3281] = inputs[92];
    assign layer0_outputs[3282] = inputs[253];
    assign layer0_outputs[3283] = ~((inputs[80]) ^ (inputs[41]));
    assign layer0_outputs[3284] = (inputs[391]) & ~(inputs[543]);
    assign layer0_outputs[3285] = (inputs[801]) ^ (inputs[463]);
    assign layer0_outputs[3286] = ~(inputs[209]) | (inputs[442]);
    assign layer0_outputs[3287] = (inputs[214]) & ~(inputs[191]);
    assign layer0_outputs[3288] = ~(inputs[652]);
    assign layer0_outputs[3289] = ~(inputs[917]);
    assign layer0_outputs[3290] = ~(inputs[821]) | (inputs[542]);
    assign layer0_outputs[3291] = ~((inputs[47]) ^ (inputs[433]));
    assign layer0_outputs[3292] = inputs[792];
    assign layer0_outputs[3293] = 1'b1;
    assign layer0_outputs[3294] = ~((inputs[441]) ^ (inputs[986]));
    assign layer0_outputs[3295] = ~(inputs[654]) | (inputs[439]);
    assign layer0_outputs[3296] = (inputs[259]) | (inputs[167]);
    assign layer0_outputs[3297] = inputs[777];
    assign layer0_outputs[3298] = (inputs[823]) & ~(inputs[968]);
    assign layer0_outputs[3299] = ~((inputs[409]) ^ (inputs[981]));
    assign layer0_outputs[3300] = ~(inputs[680]);
    assign layer0_outputs[3301] = ~((inputs[371]) | (inputs[948]));
    assign layer0_outputs[3302] = 1'b0;
    assign layer0_outputs[3303] = 1'b1;
    assign layer0_outputs[3304] = (inputs[889]) ^ (inputs[877]);
    assign layer0_outputs[3305] = ~((inputs[310]) | (inputs[264]));
    assign layer0_outputs[3306] = inputs[372];
    assign layer0_outputs[3307] = (inputs[342]) & ~(inputs[489]);
    assign layer0_outputs[3308] = (inputs[6]) & ~(inputs[514]);
    assign layer0_outputs[3309] = (inputs[268]) ^ (inputs[690]);
    assign layer0_outputs[3310] = (inputs[36]) ^ (inputs[645]);
    assign layer0_outputs[3311] = ~((inputs[863]) | (inputs[921]));
    assign layer0_outputs[3312] = (inputs[534]) | (inputs[878]);
    assign layer0_outputs[3313] = 1'b1;
    assign layer0_outputs[3314] = 1'b1;
    assign layer0_outputs[3315] = ~(inputs[851]);
    assign layer0_outputs[3316] = (inputs[164]) | (inputs[853]);
    assign layer0_outputs[3317] = inputs[584];
    assign layer0_outputs[3318] = ~(inputs[718]) | (inputs[270]);
    assign layer0_outputs[3319] = ~(inputs[584]) | (inputs[863]);
    assign layer0_outputs[3320] = ~((inputs[965]) | (inputs[594]));
    assign layer0_outputs[3321] = (inputs[764]) & (inputs[72]);
    assign layer0_outputs[3322] = ~((inputs[348]) | (inputs[284]));
    assign layer0_outputs[3323] = inputs[433];
    assign layer0_outputs[3324] = ~(inputs[428]) | (inputs[348]);
    assign layer0_outputs[3325] = (inputs[726]) & ~(inputs[505]);
    assign layer0_outputs[3326] = ~((inputs[928]) ^ (inputs[704]));
    assign layer0_outputs[3327] = ~(inputs[705]) | (inputs[911]);
    assign layer0_outputs[3328] = ~((inputs[45]) | (inputs[233]));
    assign layer0_outputs[3329] = inputs[883];
    assign layer0_outputs[3330] = ~((inputs[145]) | (inputs[626]));
    assign layer0_outputs[3331] = ~(inputs[682]) | (inputs[9]);
    assign layer0_outputs[3332] = ~(inputs[231]);
    assign layer0_outputs[3333] = inputs[619];
    assign layer0_outputs[3334] = (inputs[513]) ^ (inputs[363]);
    assign layer0_outputs[3335] = (inputs[601]) & ~(inputs[16]);
    assign layer0_outputs[3336] = ~(inputs[848]) | (inputs[763]);
    assign layer0_outputs[3337] = inputs[442];
    assign layer0_outputs[3338] = (inputs[919]) | (inputs[418]);
    assign layer0_outputs[3339] = (inputs[464]) & ~(inputs[391]);
    assign layer0_outputs[3340] = 1'b1;
    assign layer0_outputs[3341] = ~(inputs[914]);
    assign layer0_outputs[3342] = ~(inputs[240]) | (inputs[704]);
    assign layer0_outputs[3343] = (inputs[182]) ^ (inputs[248]);
    assign layer0_outputs[3344] = inputs[658];
    assign layer0_outputs[3345] = ~((inputs[701]) | (inputs[504]));
    assign layer0_outputs[3346] = (inputs[352]) & (inputs[145]);
    assign layer0_outputs[3347] = (inputs[586]) | (inputs[210]);
    assign layer0_outputs[3348] = inputs[716];
    assign layer0_outputs[3349] = (inputs[240]) ^ (inputs[244]);
    assign layer0_outputs[3350] = (inputs[290]) ^ (inputs[733]);
    assign layer0_outputs[3351] = inputs[403];
    assign layer0_outputs[3352] = (inputs[423]) & (inputs[37]);
    assign layer0_outputs[3353] = ~((inputs[262]) ^ (inputs[364]));
    assign layer0_outputs[3354] = inputs[273];
    assign layer0_outputs[3355] = inputs[506];
    assign layer0_outputs[3356] = ~(inputs[628]);
    assign layer0_outputs[3357] = (inputs[26]) & (inputs[734]);
    assign layer0_outputs[3358] = inputs[205];
    assign layer0_outputs[3359] = ~((inputs[980]) | (inputs[185]));
    assign layer0_outputs[3360] = (inputs[679]) ^ (inputs[975]);
    assign layer0_outputs[3361] = ~((inputs[750]) | (inputs[139]));
    assign layer0_outputs[3362] = (inputs[381]) ^ (inputs[912]);
    assign layer0_outputs[3363] = (inputs[739]) | (inputs[45]);
    assign layer0_outputs[3364] = ~((inputs[405]) ^ (inputs[576]));
    assign layer0_outputs[3365] = inputs[778];
    assign layer0_outputs[3366] = ~((inputs[472]) | (inputs[965]));
    assign layer0_outputs[3367] = inputs[489];
    assign layer0_outputs[3368] = ~((inputs[452]) & (inputs[188]));
    assign layer0_outputs[3369] = ~((inputs[64]) | (inputs[881]));
    assign layer0_outputs[3370] = ~(inputs[949]) | (inputs[79]);
    assign layer0_outputs[3371] = (inputs[175]) & ~(inputs[868]);
    assign layer0_outputs[3372] = (inputs[429]) & ~(inputs[935]);
    assign layer0_outputs[3373] = (inputs[688]) & ~(inputs[920]);
    assign layer0_outputs[3374] = (inputs[592]) | (inputs[501]);
    assign layer0_outputs[3375] = (inputs[252]) | (inputs[316]);
    assign layer0_outputs[3376] = (inputs[67]) & ~(inputs[97]);
    assign layer0_outputs[3377] = ~(inputs[133]) | (inputs[514]);
    assign layer0_outputs[3378] = ~(inputs[519]) | (inputs[960]);
    assign layer0_outputs[3379] = inputs[605];
    assign layer0_outputs[3380] = ~((inputs[852]) ^ (inputs[930]));
    assign layer0_outputs[3381] = ~(inputs[801]);
    assign layer0_outputs[3382] = ~(inputs[107]);
    assign layer0_outputs[3383] = inputs[395];
    assign layer0_outputs[3384] = inputs[239];
    assign layer0_outputs[3385] = inputs[707];
    assign layer0_outputs[3386] = (inputs[509]) ^ (inputs[659]);
    assign layer0_outputs[3387] = inputs[287];
    assign layer0_outputs[3388] = ~(inputs[838]) | (inputs[992]);
    assign layer0_outputs[3389] = (inputs[525]) | (inputs[235]);
    assign layer0_outputs[3390] = ~((inputs[913]) | (inputs[356]));
    assign layer0_outputs[3391] = ~(inputs[843]) | (inputs[99]);
    assign layer0_outputs[3392] = ~(inputs[275]);
    assign layer0_outputs[3393] = inputs[119];
    assign layer0_outputs[3394] = ~((inputs[546]) ^ (inputs[310]));
    assign layer0_outputs[3395] = inputs[490];
    assign layer0_outputs[3396] = ~(inputs[878]) | (inputs[990]);
    assign layer0_outputs[3397] = (inputs[714]) & ~(inputs[526]);
    assign layer0_outputs[3398] = (inputs[757]) ^ (inputs[126]);
    assign layer0_outputs[3399] = ~((inputs[508]) | (inputs[438]));
    assign layer0_outputs[3400] = ~((inputs[177]) | (inputs[638]));
    assign layer0_outputs[3401] = (inputs[567]) & (inputs[713]);
    assign layer0_outputs[3402] = ~(inputs[361]) | (inputs[832]);
    assign layer0_outputs[3403] = ~(inputs[954]) | (inputs[565]);
    assign layer0_outputs[3404] = (inputs[420]) ^ (inputs[323]);
    assign layer0_outputs[3405] = ~((inputs[874]) & (inputs[35]));
    assign layer0_outputs[3406] = (inputs[396]) & ~(inputs[718]);
    assign layer0_outputs[3407] = ~(inputs[518]) | (inputs[889]);
    assign layer0_outputs[3408] = ~((inputs[344]) | (inputs[339]));
    assign layer0_outputs[3409] = ~((inputs[1016]) & (inputs[277]));
    assign layer0_outputs[3410] = inputs[702];
    assign layer0_outputs[3411] = ~(inputs[901]);
    assign layer0_outputs[3412] = ~(inputs[735]);
    assign layer0_outputs[3413] = (inputs[54]) & ~(inputs[0]);
    assign layer0_outputs[3414] = (inputs[828]) | (inputs[724]);
    assign layer0_outputs[3415] = inputs[886];
    assign layer0_outputs[3416] = ~((inputs[630]) | (inputs[892]));
    assign layer0_outputs[3417] = ~((inputs[562]) | (inputs[836]));
    assign layer0_outputs[3418] = ~((inputs[254]) | (inputs[497]));
    assign layer0_outputs[3419] = ~((inputs[761]) ^ (inputs[505]));
    assign layer0_outputs[3420] = ~(inputs[376]);
    assign layer0_outputs[3421] = ~(inputs[653]);
    assign layer0_outputs[3422] = ~((inputs[372]) | (inputs[457]));
    assign layer0_outputs[3423] = ~((inputs[259]) | (inputs[277]));
    assign layer0_outputs[3424] = (inputs[956]) | (inputs[25]);
    assign layer0_outputs[3425] = (inputs[473]) ^ (inputs[60]);
    assign layer0_outputs[3426] = ~((inputs[873]) | (inputs[788]));
    assign layer0_outputs[3427] = (inputs[738]) | (inputs[458]);
    assign layer0_outputs[3428] = (inputs[988]) & ~(inputs[178]);
    assign layer0_outputs[3429] = (inputs[854]) & ~(inputs[38]);
    assign layer0_outputs[3430] = (inputs[548]) & ~(inputs[40]);
    assign layer0_outputs[3431] = (inputs[1003]) & (inputs[194]);
    assign layer0_outputs[3432] = ~(inputs[772]) | (inputs[935]);
    assign layer0_outputs[3433] = (inputs[457]) & ~(inputs[835]);
    assign layer0_outputs[3434] = (inputs[904]) | (inputs[481]);
    assign layer0_outputs[3435] = (inputs[359]) & ~(inputs[9]);
    assign layer0_outputs[3436] = (inputs[130]) & (inputs[289]);
    assign layer0_outputs[3437] = inputs[181];
    assign layer0_outputs[3438] = inputs[712];
    assign layer0_outputs[3439] = (inputs[1]) ^ (inputs[458]);
    assign layer0_outputs[3440] = ~(inputs[933]) | (inputs[898]);
    assign layer0_outputs[3441] = (inputs[628]) & ~(inputs[633]);
    assign layer0_outputs[3442] = inputs[702];
    assign layer0_outputs[3443] = (inputs[953]) & ~(inputs[477]);
    assign layer0_outputs[3444] = (inputs[582]) | (inputs[569]);
    assign layer0_outputs[3445] = inputs[746];
    assign layer0_outputs[3446] = ~(inputs[308]) | (inputs[445]);
    assign layer0_outputs[3447] = inputs[130];
    assign layer0_outputs[3448] = ~(inputs[961]);
    assign layer0_outputs[3449] = ~((inputs[756]) & (inputs[547]));
    assign layer0_outputs[3450] = (inputs[313]) | (inputs[396]);
    assign layer0_outputs[3451] = inputs[488];
    assign layer0_outputs[3452] = ~(inputs[408]);
    assign layer0_outputs[3453] = ~((inputs[650]) ^ (inputs[655]));
    assign layer0_outputs[3454] = inputs[291];
    assign layer0_outputs[3455] = (inputs[929]) & (inputs[836]);
    assign layer0_outputs[3456] = (inputs[413]) & (inputs[24]);
    assign layer0_outputs[3457] = ~(inputs[672]);
    assign layer0_outputs[3458] = ~((inputs[942]) | (inputs[33]));
    assign layer0_outputs[3459] = (inputs[923]) | (inputs[366]);
    assign layer0_outputs[3460] = (inputs[587]) & ~(inputs[935]);
    assign layer0_outputs[3461] = inputs[575];
    assign layer0_outputs[3462] = ~(inputs[707]) | (inputs[450]);
    assign layer0_outputs[3463] = ~((inputs[456]) | (inputs[102]));
    assign layer0_outputs[3464] = ~(inputs[276]);
    assign layer0_outputs[3465] = inputs[771];
    assign layer0_outputs[3466] = (inputs[93]) ^ (inputs[973]);
    assign layer0_outputs[3467] = ~(inputs[814]);
    assign layer0_outputs[3468] = (inputs[852]) & ~(inputs[907]);
    assign layer0_outputs[3469] = inputs[605];
    assign layer0_outputs[3470] = (inputs[932]) & ~(inputs[351]);
    assign layer0_outputs[3471] = (inputs[74]) & (inputs[943]);
    assign layer0_outputs[3472] = inputs[87];
    assign layer0_outputs[3473] = 1'b0;
    assign layer0_outputs[3474] = 1'b1;
    assign layer0_outputs[3475] = (inputs[728]) & ~(inputs[219]);
    assign layer0_outputs[3476] = ~((inputs[1]) | (inputs[664]));
    assign layer0_outputs[3477] = 1'b0;
    assign layer0_outputs[3478] = inputs[136];
    assign layer0_outputs[3479] = ~(inputs[13]);
    assign layer0_outputs[3480] = (inputs[884]) & ~(inputs[107]);
    assign layer0_outputs[3481] = ~((inputs[374]) ^ (inputs[340]));
    assign layer0_outputs[3482] = ~(inputs[90]);
    assign layer0_outputs[3483] = ~(inputs[721]) | (inputs[361]);
    assign layer0_outputs[3484] = ~(inputs[625]);
    assign layer0_outputs[3485] = (inputs[157]) | (inputs[597]);
    assign layer0_outputs[3486] = (inputs[813]) & ~(inputs[869]);
    assign layer0_outputs[3487] = 1'b1;
    assign layer0_outputs[3488] = ~((inputs[805]) | (inputs[205]));
    assign layer0_outputs[3489] = ~((inputs[173]) ^ (inputs[927]));
    assign layer0_outputs[3490] = inputs[520];
    assign layer0_outputs[3491] = ~((inputs[487]) | (inputs[479]));
    assign layer0_outputs[3492] = (inputs[548]) | (inputs[192]);
    assign layer0_outputs[3493] = (inputs[237]) | (inputs[950]);
    assign layer0_outputs[3494] = (inputs[315]) & ~(inputs[61]);
    assign layer0_outputs[3495] = ~(inputs[212]) | (inputs[1021]);
    assign layer0_outputs[3496] = (inputs[11]) ^ (inputs[471]);
    assign layer0_outputs[3497] = 1'b1;
    assign layer0_outputs[3498] = (inputs[950]) | (inputs[390]);
    assign layer0_outputs[3499] = ~((inputs[397]) ^ (inputs[578]));
    assign layer0_outputs[3500] = inputs[776];
    assign layer0_outputs[3501] = (inputs[411]) ^ (inputs[918]);
    assign layer0_outputs[3502] = (inputs[459]) | (inputs[748]);
    assign layer0_outputs[3503] = ~(inputs[175]) | (inputs[131]);
    assign layer0_outputs[3504] = (inputs[341]) | (inputs[857]);
    assign layer0_outputs[3505] = ~(inputs[427]);
    assign layer0_outputs[3506] = ~(inputs[686]) | (inputs[256]);
    assign layer0_outputs[3507] = inputs[933];
    assign layer0_outputs[3508] = (inputs[505]) & ~(inputs[34]);
    assign layer0_outputs[3509] = ~((inputs[760]) ^ (inputs[813]));
    assign layer0_outputs[3510] = ~(inputs[203]) | (inputs[984]);
    assign layer0_outputs[3511] = inputs[115];
    assign layer0_outputs[3512] = (inputs[429]) & ~(inputs[158]);
    assign layer0_outputs[3513] = inputs[315];
    assign layer0_outputs[3514] = inputs[256];
    assign layer0_outputs[3515] = (inputs[226]) ^ (inputs[777]);
    assign layer0_outputs[3516] = 1'b1;
    assign layer0_outputs[3517] = ~((inputs[327]) | (inputs[515]));
    assign layer0_outputs[3518] = (inputs[439]) | (inputs[589]);
    assign layer0_outputs[3519] = ~(inputs[843]) | (inputs[995]);
    assign layer0_outputs[3520] = ~((inputs[368]) | (inputs[740]));
    assign layer0_outputs[3521] = ~((inputs[533]) | (inputs[372]));
    assign layer0_outputs[3522] = (inputs[79]) & ~(inputs[227]);
    assign layer0_outputs[3523] = ~(inputs[870]);
    assign layer0_outputs[3524] = ~((inputs[62]) ^ (inputs[709]));
    assign layer0_outputs[3525] = ~(inputs[93]);
    assign layer0_outputs[3526] = ~((inputs[1003]) & (inputs[614]));
    assign layer0_outputs[3527] = (inputs[404]) | (inputs[588]);
    assign layer0_outputs[3528] = ~((inputs[146]) | (inputs[515]));
    assign layer0_outputs[3529] = ~(inputs[791]) | (inputs[832]);
    assign layer0_outputs[3530] = ~((inputs[782]) & (inputs[700]));
    assign layer0_outputs[3531] = (inputs[353]) & ~(inputs[929]);
    assign layer0_outputs[3532] = inputs[648];
    assign layer0_outputs[3533] = ~((inputs[754]) ^ (inputs[850]));
    assign layer0_outputs[3534] = ~((inputs[170]) | (inputs[1023]));
    assign layer0_outputs[3535] = ~((inputs[71]) ^ (inputs[322]));
    assign layer0_outputs[3536] = (inputs[486]) ^ (inputs[147]);
    assign layer0_outputs[3537] = (inputs[508]) & (inputs[510]);
    assign layer0_outputs[3538] = ~(inputs[85]) | (inputs[162]);
    assign layer0_outputs[3539] = ~(inputs[398]) | (inputs[822]);
    assign layer0_outputs[3540] = (inputs[206]) & ~(inputs[634]);
    assign layer0_outputs[3541] = (inputs[945]) & ~(inputs[56]);
    assign layer0_outputs[3542] = ~(inputs[470]);
    assign layer0_outputs[3543] = (inputs[114]) | (inputs[134]);
    assign layer0_outputs[3544] = ~((inputs[842]) | (inputs[410]));
    assign layer0_outputs[3545] = ~(inputs[561]) | (inputs[172]);
    assign layer0_outputs[3546] = ~(inputs[216]);
    assign layer0_outputs[3547] = (inputs[675]) & ~(inputs[961]);
    assign layer0_outputs[3548] = (inputs[363]) & ~(inputs[726]);
    assign layer0_outputs[3549] = ~((inputs[571]) ^ (inputs[273]));
    assign layer0_outputs[3550] = (inputs[561]) & ~(inputs[199]);
    assign layer0_outputs[3551] = ~(inputs[919]);
    assign layer0_outputs[3552] = ~(inputs[361]);
    assign layer0_outputs[3553] = ~((inputs[799]) | (inputs[716]));
    assign layer0_outputs[3554] = inputs[657];
    assign layer0_outputs[3555] = ~(inputs[664]);
    assign layer0_outputs[3556] = ~((inputs[966]) ^ (inputs[908]));
    assign layer0_outputs[3557] = ~(inputs[674]) | (inputs[265]);
    assign layer0_outputs[3558] = ~((inputs[532]) & (inputs[993]));
    assign layer0_outputs[3559] = ~(inputs[795]);
    assign layer0_outputs[3560] = ~((inputs[690]) ^ (inputs[15]));
    assign layer0_outputs[3561] = inputs[419];
    assign layer0_outputs[3562] = ~((inputs[812]) | (inputs[409]));
    assign layer0_outputs[3563] = ~((inputs[752]) | (inputs[141]));
    assign layer0_outputs[3564] = (inputs[210]) & ~(inputs[703]);
    assign layer0_outputs[3565] = (inputs[393]) | (inputs[532]);
    assign layer0_outputs[3566] = ~((inputs[930]) | (inputs[887]));
    assign layer0_outputs[3567] = (inputs[1]) | (inputs[656]);
    assign layer0_outputs[3568] = (inputs[43]) & ~(inputs[920]);
    assign layer0_outputs[3569] = inputs[550];
    assign layer0_outputs[3570] = (inputs[272]) & ~(inputs[709]);
    assign layer0_outputs[3571] = (inputs[538]) | (inputs[450]);
    assign layer0_outputs[3572] = ~((inputs[447]) & (inputs[226]));
    assign layer0_outputs[3573] = ~(inputs[613]) | (inputs[966]);
    assign layer0_outputs[3574] = ~(inputs[558]);
    assign layer0_outputs[3575] = ~((inputs[26]) | (inputs[62]));
    assign layer0_outputs[3576] = inputs[471];
    assign layer0_outputs[3577] = ~(inputs[589]) | (inputs[386]);
    assign layer0_outputs[3578] = (inputs[379]) | (inputs[311]);
    assign layer0_outputs[3579] = ~((inputs[865]) ^ (inputs[1]));
    assign layer0_outputs[3580] = inputs[187];
    assign layer0_outputs[3581] = ~(inputs[50]) | (inputs[65]);
    assign layer0_outputs[3582] = ~(inputs[369]);
    assign layer0_outputs[3583] = inputs[100];
    assign layer0_outputs[3584] = inputs[787];
    assign layer0_outputs[3585] = (inputs[316]) & ~(inputs[766]);
    assign layer0_outputs[3586] = ~(inputs[874]) | (inputs[669]);
    assign layer0_outputs[3587] = (inputs[462]) | (inputs[492]);
    assign layer0_outputs[3588] = ~((inputs[158]) ^ (inputs[1006]));
    assign layer0_outputs[3589] = ~(inputs[52]);
    assign layer0_outputs[3590] = ~(inputs[660]) | (inputs[453]);
    assign layer0_outputs[3591] = ~(inputs[196]);
    assign layer0_outputs[3592] = ~((inputs[289]) | (inputs[10]));
    assign layer0_outputs[3593] = inputs[344];
    assign layer0_outputs[3594] = ~(inputs[847]);
    assign layer0_outputs[3595] = inputs[46];
    assign layer0_outputs[3596] = (inputs[983]) & (inputs[737]);
    assign layer0_outputs[3597] = inputs[990];
    assign layer0_outputs[3598] = inputs[442];
    assign layer0_outputs[3599] = (inputs[324]) ^ (inputs[710]);
    assign layer0_outputs[3600] = ~(inputs[526]);
    assign layer0_outputs[3601] = (inputs[162]) | (inputs[589]);
    assign layer0_outputs[3602] = ~((inputs[390]) & (inputs[960]));
    assign layer0_outputs[3603] = inputs[1014];
    assign layer0_outputs[3604] = ~((inputs[929]) ^ (inputs[56]));
    assign layer0_outputs[3605] = ~(inputs[893]);
    assign layer0_outputs[3606] = ~(inputs[986]) | (inputs[482]);
    assign layer0_outputs[3607] = (inputs[502]) ^ (inputs[373]);
    assign layer0_outputs[3608] = ~(inputs[536]);
    assign layer0_outputs[3609] = (inputs[849]) & ~(inputs[902]);
    assign layer0_outputs[3610] = ~((inputs[57]) ^ (inputs[583]));
    assign layer0_outputs[3611] = (inputs[337]) | (inputs[275]);
    assign layer0_outputs[3612] = ~(inputs[229]);
    assign layer0_outputs[3613] = (inputs[1015]) | (inputs[870]);
    assign layer0_outputs[3614] = (inputs[934]) | (inputs[545]);
    assign layer0_outputs[3615] = (inputs[588]) | (inputs[153]);
    assign layer0_outputs[3616] = ~((inputs[831]) | (inputs[305]));
    assign layer0_outputs[3617] = ~((inputs[998]) | (inputs[396]));
    assign layer0_outputs[3618] = ~(inputs[566]) | (inputs[747]);
    assign layer0_outputs[3619] = 1'b1;
    assign layer0_outputs[3620] = 1'b1;
    assign layer0_outputs[3621] = ~((inputs[770]) | (inputs[352]));
    assign layer0_outputs[3622] = 1'b0;
    assign layer0_outputs[3623] = ~((inputs[983]) ^ (inputs[761]));
    assign layer0_outputs[3624] = (inputs[1011]) | (inputs[715]);
    assign layer0_outputs[3625] = inputs[333];
    assign layer0_outputs[3626] = inputs[946];
    assign layer0_outputs[3627] = ~((inputs[91]) ^ (inputs[265]));
    assign layer0_outputs[3628] = (inputs[95]) | (inputs[212]);
    assign layer0_outputs[3629] = (inputs[750]) ^ (inputs[492]);
    assign layer0_outputs[3630] = ~(inputs[449]) | (inputs[1022]);
    assign layer0_outputs[3631] = ~((inputs[169]) ^ (inputs[584]));
    assign layer0_outputs[3632] = ~(inputs[678]);
    assign layer0_outputs[3633] = ~((inputs[475]) & (inputs[847]));
    assign layer0_outputs[3634] = ~(inputs[773]);
    assign layer0_outputs[3635] = inputs[180];
    assign layer0_outputs[3636] = inputs[142];
    assign layer0_outputs[3637] = (inputs[788]) ^ (inputs[18]);
    assign layer0_outputs[3638] = ~((inputs[461]) ^ (inputs[671]));
    assign layer0_outputs[3639] = (inputs[365]) | (inputs[97]);
    assign layer0_outputs[3640] = ~(inputs[495]) | (inputs[734]);
    assign layer0_outputs[3641] = ~((inputs[811]) ^ (inputs[132]));
    assign layer0_outputs[3642] = (inputs[899]) | (inputs[443]);
    assign layer0_outputs[3643] = inputs[674];
    assign layer0_outputs[3644] = ~((inputs[506]) ^ (inputs[805]));
    assign layer0_outputs[3645] = (inputs[370]) ^ (inputs[480]);
    assign layer0_outputs[3646] = ~((inputs[894]) ^ (inputs[751]));
    assign layer0_outputs[3647] = 1'b0;
    assign layer0_outputs[3648] = (inputs[729]) ^ (inputs[613]);
    assign layer0_outputs[3649] = ~(inputs[496]) | (inputs[451]);
    assign layer0_outputs[3650] = (inputs[530]) & ~(inputs[387]);
    assign layer0_outputs[3651] = (inputs[919]) | (inputs[549]);
    assign layer0_outputs[3652] = (inputs[326]) | (inputs[592]);
    assign layer0_outputs[3653] = ~(inputs[241]);
    assign layer0_outputs[3654] = (inputs[646]) & ~(inputs[707]);
    assign layer0_outputs[3655] = ~(inputs[510]) | (inputs[991]);
    assign layer0_outputs[3656] = ~(inputs[401]) | (inputs[327]);
    assign layer0_outputs[3657] = inputs[413];
    assign layer0_outputs[3658] = (inputs[338]) & ~(inputs[131]);
    assign layer0_outputs[3659] = ~((inputs[260]) ^ (inputs[627]));
    assign layer0_outputs[3660] = ~((inputs[962]) & (inputs[412]));
    assign layer0_outputs[3661] = ~(inputs[673]) | (inputs[382]);
    assign layer0_outputs[3662] = ~((inputs[1021]) ^ (inputs[206]));
    assign layer0_outputs[3663] = (inputs[198]) | (inputs[589]);
    assign layer0_outputs[3664] = ~(inputs[864]) | (inputs[267]);
    assign layer0_outputs[3665] = (inputs[216]) | (inputs[358]);
    assign layer0_outputs[3666] = (inputs[567]) & ~(inputs[93]);
    assign layer0_outputs[3667] = ~(inputs[214]) | (inputs[160]);
    assign layer0_outputs[3668] = 1'b1;
    assign layer0_outputs[3669] = inputs[791];
    assign layer0_outputs[3670] = ~(inputs[363]);
    assign layer0_outputs[3671] = (inputs[208]) ^ (inputs[932]);
    assign layer0_outputs[3672] = ~((inputs[912]) ^ (inputs[7]));
    assign layer0_outputs[3673] = (inputs[39]) ^ (inputs[716]);
    assign layer0_outputs[3674] = ~(inputs[835]) | (inputs[1019]);
    assign layer0_outputs[3675] = ~((inputs[337]) | (inputs[1016]));
    assign layer0_outputs[3676] = (inputs[255]) & ~(inputs[133]);
    assign layer0_outputs[3677] = 1'b0;
    assign layer0_outputs[3678] = ~(inputs[441]) | (inputs[610]);
    assign layer0_outputs[3679] = (inputs[307]) & ~(inputs[587]);
    assign layer0_outputs[3680] = inputs[331];
    assign layer0_outputs[3681] = ~((inputs[634]) | (inputs[147]));
    assign layer0_outputs[3682] = ~(inputs[207]);
    assign layer0_outputs[3683] = (inputs[727]) & ~(inputs[89]);
    assign layer0_outputs[3684] = (inputs[319]) ^ (inputs[507]);
    assign layer0_outputs[3685] = ~((inputs[418]) ^ (inputs[398]));
    assign layer0_outputs[3686] = (inputs[606]) ^ (inputs[345]);
    assign layer0_outputs[3687] = (inputs[336]) & ~(inputs[356]);
    assign layer0_outputs[3688] = inputs[337];
    assign layer0_outputs[3689] = (inputs[603]) ^ (inputs[1002]);
    assign layer0_outputs[3690] = ~((inputs[563]) | (inputs[451]));
    assign layer0_outputs[3691] = (inputs[490]) & ~(inputs[699]);
    assign layer0_outputs[3692] = (inputs[873]) ^ (inputs[749]);
    assign layer0_outputs[3693] = (inputs[127]) | (inputs[906]);
    assign layer0_outputs[3694] = 1'b0;
    assign layer0_outputs[3695] = ~(inputs[845]) | (inputs[867]);
    assign layer0_outputs[3696] = (inputs[620]) & ~(inputs[932]);
    assign layer0_outputs[3697] = (inputs[1001]) | (inputs[647]);
    assign layer0_outputs[3698] = inputs[521];
    assign layer0_outputs[3699] = inputs[524];
    assign layer0_outputs[3700] = ~(inputs[372]) | (inputs[708]);
    assign layer0_outputs[3701] = ~((inputs[462]) ^ (inputs[830]));
    assign layer0_outputs[3702] = inputs[247];
    assign layer0_outputs[3703] = ~((inputs[736]) & (inputs[521]));
    assign layer0_outputs[3704] = (inputs[525]) | (inputs[719]);
    assign layer0_outputs[3705] = ~(inputs[502]) | (inputs[217]);
    assign layer0_outputs[3706] = (inputs[415]) ^ (inputs[855]);
    assign layer0_outputs[3707] = ~((inputs[208]) | (inputs[616]));
    assign layer0_outputs[3708] = (inputs[759]) & ~(inputs[92]);
    assign layer0_outputs[3709] = (inputs[881]) | (inputs[768]);
    assign layer0_outputs[3710] = ~(inputs[691]) | (inputs[673]);
    assign layer0_outputs[3711] = (inputs[66]) ^ (inputs[360]);
    assign layer0_outputs[3712] = ~((inputs[124]) ^ (inputs[421]));
    assign layer0_outputs[3713] = inputs[853];
    assign layer0_outputs[3714] = inputs[627];
    assign layer0_outputs[3715] = ~(inputs[226]);
    assign layer0_outputs[3716] = ~((inputs[81]) ^ (inputs[893]));
    assign layer0_outputs[3717] = ~(inputs[986]);
    assign layer0_outputs[3718] = ~(inputs[815]);
    assign layer0_outputs[3719] = ~(inputs[691]) | (inputs[349]);
    assign layer0_outputs[3720] = (inputs[939]) & (inputs[360]);
    assign layer0_outputs[3721] = inputs[661];
    assign layer0_outputs[3722] = (inputs[293]) & ~(inputs[932]);
    assign layer0_outputs[3723] = ~((inputs[423]) | (inputs[907]));
    assign layer0_outputs[3724] = (inputs[373]) & ~(inputs[868]);
    assign layer0_outputs[3725] = ~((inputs[375]) | (inputs[950]));
    assign layer0_outputs[3726] = 1'b1;
    assign layer0_outputs[3727] = ~((inputs[931]) | (inputs[561]));
    assign layer0_outputs[3728] = (inputs[207]) & ~(inputs[428]);
    assign layer0_outputs[3729] = inputs[1012];
    assign layer0_outputs[3730] = ~(inputs[499]);
    assign layer0_outputs[3731] = ~((inputs[150]) ^ (inputs[973]));
    assign layer0_outputs[3732] = (inputs[509]) ^ (inputs[915]);
    assign layer0_outputs[3733] = (inputs[367]) & ~(inputs[230]);
    assign layer0_outputs[3734] = ~(inputs[27]) | (inputs[477]);
    assign layer0_outputs[3735] = (inputs[691]) & ~(inputs[972]);
    assign layer0_outputs[3736] = ~((inputs[899]) ^ (inputs[854]));
    assign layer0_outputs[3737] = (inputs[584]) ^ (inputs[51]);
    assign layer0_outputs[3738] = ~(inputs[279]);
    assign layer0_outputs[3739] = (inputs[543]) & ~(inputs[283]);
    assign layer0_outputs[3740] = ~(inputs[553]);
    assign layer0_outputs[3741] = ~((inputs[966]) | (inputs[468]));
    assign layer0_outputs[3742] = ~(inputs[679]);
    assign layer0_outputs[3743] = (inputs[431]) | (inputs[303]);
    assign layer0_outputs[3744] = (inputs[856]) | (inputs[80]);
    assign layer0_outputs[3745] = (inputs[98]) & (inputs[767]);
    assign layer0_outputs[3746] = ~(inputs[387]) | (inputs[53]);
    assign layer0_outputs[3747] = ~((inputs[38]) ^ (inputs[741]));
    assign layer0_outputs[3748] = (inputs[713]) & ~(inputs[66]);
    assign layer0_outputs[3749] = 1'b0;
    assign layer0_outputs[3750] = ~((inputs[783]) & (inputs[290]));
    assign layer0_outputs[3751] = (inputs[551]) & ~(inputs[293]);
    assign layer0_outputs[3752] = ~(inputs[318]) | (inputs[762]);
    assign layer0_outputs[3753] = ~(inputs[695]);
    assign layer0_outputs[3754] = ~(inputs[69]) | (inputs[477]);
    assign layer0_outputs[3755] = ~(inputs[823]) | (inputs[125]);
    assign layer0_outputs[3756] = ~((inputs[742]) | (inputs[971]));
    assign layer0_outputs[3757] = ~(inputs[442]);
    assign layer0_outputs[3758] = (inputs[68]) | (inputs[971]);
    assign layer0_outputs[3759] = ~((inputs[235]) | (inputs[605]));
    assign layer0_outputs[3760] = ~((inputs[751]) ^ (inputs[217]));
    assign layer0_outputs[3761] = (inputs[53]) & (inputs[77]);
    assign layer0_outputs[3762] = ~(inputs[975]);
    assign layer0_outputs[3763] = (inputs[954]) & ~(inputs[767]);
    assign layer0_outputs[3764] = 1'b1;
    assign layer0_outputs[3765] = ~((inputs[236]) | (inputs[664]));
    assign layer0_outputs[3766] = (inputs[434]) | (inputs[654]);
    assign layer0_outputs[3767] = ~((inputs[680]) & (inputs[634]));
    assign layer0_outputs[3768] = ~(inputs[51]);
    assign layer0_outputs[3769] = ~((inputs[972]) | (inputs[729]));
    assign layer0_outputs[3770] = inputs[683];
    assign layer0_outputs[3771] = ~(inputs[770]) | (inputs[925]);
    assign layer0_outputs[3772] = ~(inputs[462]) | (inputs[655]);
    assign layer0_outputs[3773] = (inputs[932]) & ~(inputs[111]);
    assign layer0_outputs[3774] = (inputs[334]) | (inputs[393]);
    assign layer0_outputs[3775] = ~((inputs[9]) ^ (inputs[684]));
    assign layer0_outputs[3776] = ~((inputs[947]) ^ (inputs[808]));
    assign layer0_outputs[3777] = ~(inputs[748]);
    assign layer0_outputs[3778] = ~((inputs[821]) | (inputs[729]));
    assign layer0_outputs[3779] = inputs[26];
    assign layer0_outputs[3780] = (inputs[264]) | (inputs[889]);
    assign layer0_outputs[3781] = (inputs[324]) & (inputs[312]);
    assign layer0_outputs[3782] = ~((inputs[820]) | (inputs[232]));
    assign layer0_outputs[3783] = (inputs[998]) & ~(inputs[217]);
    assign layer0_outputs[3784] = ~(inputs[464]);
    assign layer0_outputs[3785] = ~(inputs[562]) | (inputs[329]);
    assign layer0_outputs[3786] = (inputs[951]) | (inputs[751]);
    assign layer0_outputs[3787] = ~((inputs[357]) ^ (inputs[805]));
    assign layer0_outputs[3788] = inputs[854];
    assign layer0_outputs[3789] = ~((inputs[749]) | (inputs[539]));
    assign layer0_outputs[3790] = inputs[721];
    assign layer0_outputs[3791] = (inputs[812]) & (inputs[471]);
    assign layer0_outputs[3792] = ~(inputs[1019]);
    assign layer0_outputs[3793] = (inputs[662]) & ~(inputs[1009]);
    assign layer0_outputs[3794] = ~(inputs[377]);
    assign layer0_outputs[3795] = (inputs[555]) | (inputs[255]);
    assign layer0_outputs[3796] = ~(inputs[788]) | (inputs[732]);
    assign layer0_outputs[3797] = inputs[493];
    assign layer0_outputs[3798] = (inputs[213]) | (inputs[91]);
    assign layer0_outputs[3799] = ~(inputs[709]);
    assign layer0_outputs[3800] = inputs[479];
    assign layer0_outputs[3801] = ~((inputs[394]) | (inputs[547]));
    assign layer0_outputs[3802] = (inputs[763]) | (inputs[799]);
    assign layer0_outputs[3803] = inputs[98];
    assign layer0_outputs[3804] = ~((inputs[116]) & (inputs[735]));
    assign layer0_outputs[3805] = (inputs[123]) ^ (inputs[388]);
    assign layer0_outputs[3806] = ~(inputs[798]) | (inputs[923]);
    assign layer0_outputs[3807] = ~((inputs[316]) | (inputs[732]));
    assign layer0_outputs[3808] = (inputs[77]) | (inputs[571]);
    assign layer0_outputs[3809] = ~(inputs[621]) | (inputs[327]);
    assign layer0_outputs[3810] = ~(inputs[430]);
    assign layer0_outputs[3811] = (inputs[514]) | (inputs[476]);
    assign layer0_outputs[3812] = inputs[281];
    assign layer0_outputs[3813] = inputs[61];
    assign layer0_outputs[3814] = inputs[558];
    assign layer0_outputs[3815] = 1'b0;
    assign layer0_outputs[3816] = ~(inputs[618]) | (inputs[920]);
    assign layer0_outputs[3817] = (inputs[404]) | (inputs[147]);
    assign layer0_outputs[3818] = ~((inputs[351]) | (inputs[334]));
    assign layer0_outputs[3819] = (inputs[177]) | (inputs[795]);
    assign layer0_outputs[3820] = ~((inputs[631]) ^ (inputs[297]));
    assign layer0_outputs[3821] = ~((inputs[223]) ^ (inputs[234]));
    assign layer0_outputs[3822] = (inputs[311]) | (inputs[332]);
    assign layer0_outputs[3823] = (inputs[131]) ^ (inputs[351]);
    assign layer0_outputs[3824] = (inputs[785]) & ~(inputs[902]);
    assign layer0_outputs[3825] = inputs[142];
    assign layer0_outputs[3826] = ~((inputs[824]) ^ (inputs[13]));
    assign layer0_outputs[3827] = inputs[155];
    assign layer0_outputs[3828] = (inputs[309]) ^ (inputs[701]);
    assign layer0_outputs[3829] = ~(inputs[532]);
    assign layer0_outputs[3830] = ~(inputs[601]) | (inputs[366]);
    assign layer0_outputs[3831] = ~((inputs[44]) | (inputs[432]));
    assign layer0_outputs[3832] = (inputs[292]) & ~(inputs[667]);
    assign layer0_outputs[3833] = ~((inputs[311]) | (inputs[860]));
    assign layer0_outputs[3834] = ~((inputs[655]) & (inputs[104]));
    assign layer0_outputs[3835] = (inputs[166]) & ~(inputs[840]);
    assign layer0_outputs[3836] = ~((inputs[818]) ^ (inputs[190]));
    assign layer0_outputs[3837] = ~((inputs[2]) ^ (inputs[667]));
    assign layer0_outputs[3838] = inputs[882];
    assign layer0_outputs[3839] = (inputs[400]) & ~(inputs[330]);
    assign layer0_outputs[3840] = inputs[941];
    assign layer0_outputs[3841] = (inputs[232]) | (inputs[790]);
    assign layer0_outputs[3842] = (inputs[34]) | (inputs[513]);
    assign layer0_outputs[3843] = ~((inputs[50]) | (inputs[274]));
    assign layer0_outputs[3844] = ~(inputs[724]);
    assign layer0_outputs[3845] = ~((inputs[730]) | (inputs[745]));
    assign layer0_outputs[3846] = ~(inputs[694]);
    assign layer0_outputs[3847] = ~(inputs[412]);
    assign layer0_outputs[3848] = (inputs[553]) & ~(inputs[916]);
    assign layer0_outputs[3849] = inputs[598];
    assign layer0_outputs[3850] = ~(inputs[520]) | (inputs[545]);
    assign layer0_outputs[3851] = 1'b1;
    assign layer0_outputs[3852] = inputs[528];
    assign layer0_outputs[3853] = ~(inputs[945]) | (inputs[576]);
    assign layer0_outputs[3854] = (inputs[476]) & (inputs[228]);
    assign layer0_outputs[3855] = ~((inputs[175]) | (inputs[9]));
    assign layer0_outputs[3856] = (inputs[781]) & ~(inputs[94]);
    assign layer0_outputs[3857] = ~((inputs[872]) | (inputs[365]));
    assign layer0_outputs[3858] = (inputs[746]) ^ (inputs[122]);
    assign layer0_outputs[3859] = ~(inputs[826]) | (inputs[254]);
    assign layer0_outputs[3860] = 1'b0;
    assign layer0_outputs[3861] = inputs[683];
    assign layer0_outputs[3862] = ~(inputs[623]);
    assign layer0_outputs[3863] = ~((inputs[817]) ^ (inputs[247]));
    assign layer0_outputs[3864] = (inputs[230]) ^ (inputs[471]);
    assign layer0_outputs[3865] = ~((inputs[996]) | (inputs[419]));
    assign layer0_outputs[3866] = ~((inputs[975]) ^ (inputs[470]));
    assign layer0_outputs[3867] = 1'b0;
    assign layer0_outputs[3868] = ~(inputs[615]);
    assign layer0_outputs[3869] = ~((inputs[745]) | (inputs[312]));
    assign layer0_outputs[3870] = (inputs[283]) & ~(inputs[604]);
    assign layer0_outputs[3871] = ~(inputs[857]) | (inputs[703]);
    assign layer0_outputs[3872] = ~((inputs[94]) | (inputs[904]));
    assign layer0_outputs[3873] = ~(inputs[269]);
    assign layer0_outputs[3874] = (inputs[763]) & ~(inputs[974]);
    assign layer0_outputs[3875] = inputs[360];
    assign layer0_outputs[3876] = (inputs[9]) | (inputs[235]);
    assign layer0_outputs[3877] = ~((inputs[548]) | (inputs[314]));
    assign layer0_outputs[3878] = ~(inputs[683]);
    assign layer0_outputs[3879] = inputs[828];
    assign layer0_outputs[3880] = ~(inputs[237]);
    assign layer0_outputs[3881] = ~((inputs[18]) ^ (inputs[469]));
    assign layer0_outputs[3882] = (inputs[687]) | (inputs[870]);
    assign layer0_outputs[3883] = (inputs[817]) ^ (inputs[466]);
    assign layer0_outputs[3884] = inputs[997];
    assign layer0_outputs[3885] = ~((inputs[933]) ^ (inputs[270]));
    assign layer0_outputs[3886] = ~((inputs[847]) | (inputs[165]));
    assign layer0_outputs[3887] = ~((inputs[888]) | (inputs[510]));
    assign layer0_outputs[3888] = (inputs[399]) & ~(inputs[385]);
    assign layer0_outputs[3889] = ~((inputs[379]) | (inputs[866]));
    assign layer0_outputs[3890] = (inputs[279]) | (inputs[851]);
    assign layer0_outputs[3891] = (inputs[563]) | (inputs[919]);
    assign layer0_outputs[3892] = ~(inputs[720]) | (inputs[644]);
    assign layer0_outputs[3893] = (inputs[384]) ^ (inputs[525]);
    assign layer0_outputs[3894] = ~(inputs[600]);
    assign layer0_outputs[3895] = inputs[173];
    assign layer0_outputs[3896] = (inputs[1002]) & (inputs[221]);
    assign layer0_outputs[3897] = (inputs[606]) & ~(inputs[482]);
    assign layer0_outputs[3898] = ~((inputs[11]) | (inputs[862]));
    assign layer0_outputs[3899] = (inputs[90]) | (inputs[61]);
    assign layer0_outputs[3900] = (inputs[498]) & ~(inputs[736]);
    assign layer0_outputs[3901] = (inputs[850]) | (inputs[253]);
    assign layer0_outputs[3902] = inputs[722];
    assign layer0_outputs[3903] = (inputs[249]) ^ (inputs[83]);
    assign layer0_outputs[3904] = ~((inputs[670]) & (inputs[485]));
    assign layer0_outputs[3905] = (inputs[25]) ^ (inputs[509]);
    assign layer0_outputs[3906] = ~((inputs[295]) | (inputs[33]));
    assign layer0_outputs[3907] = ~(inputs[395]) | (inputs[699]);
    assign layer0_outputs[3908] = ~(inputs[709]) | (inputs[260]);
    assign layer0_outputs[3909] = inputs[427];
    assign layer0_outputs[3910] = inputs[282];
    assign layer0_outputs[3911] = (inputs[637]) ^ (inputs[443]);
    assign layer0_outputs[3912] = ~(inputs[787]) | (inputs[198]);
    assign layer0_outputs[3913] = (inputs[236]) | (inputs[453]);
    assign layer0_outputs[3914] = ~(inputs[525]) | (inputs[989]);
    assign layer0_outputs[3915] = ~((inputs[322]) | (inputs[562]));
    assign layer0_outputs[3916] = (inputs[327]) & ~(inputs[892]);
    assign layer0_outputs[3917] = ~(inputs[512]);
    assign layer0_outputs[3918] = ~(inputs[331]) | (inputs[602]);
    assign layer0_outputs[3919] = ~((inputs[880]) ^ (inputs[771]));
    assign layer0_outputs[3920] = ~((inputs[243]) | (inputs[306]));
    assign layer0_outputs[3921] = (inputs[686]) & ~(inputs[380]);
    assign layer0_outputs[3922] = ~((inputs[217]) | (inputs[522]));
    assign layer0_outputs[3923] = (inputs[593]) & ~(inputs[246]);
    assign layer0_outputs[3924] = (inputs[862]) | (inputs[790]);
    assign layer0_outputs[3925] = ~((inputs[135]) | (inputs[786]));
    assign layer0_outputs[3926] = ~(inputs[563]);
    assign layer0_outputs[3927] = ~((inputs[850]) | (inputs[669]));
    assign layer0_outputs[3928] = ~(inputs[862]);
    assign layer0_outputs[3929] = 1'b1;
    assign layer0_outputs[3930] = (inputs[192]) | (inputs[207]);
    assign layer0_outputs[3931] = inputs[348];
    assign layer0_outputs[3932] = (inputs[621]) ^ (inputs[354]);
    assign layer0_outputs[3933] = inputs[310];
    assign layer0_outputs[3934] = ~(inputs[592]);
    assign layer0_outputs[3935] = inputs[818];
    assign layer0_outputs[3936] = ~((inputs[866]) ^ (inputs[906]));
    assign layer0_outputs[3937] = ~(inputs[313]);
    assign layer0_outputs[3938] = ~(inputs[601]) | (inputs[451]);
    assign layer0_outputs[3939] = inputs[35];
    assign layer0_outputs[3940] = 1'b1;
    assign layer0_outputs[3941] = (inputs[829]) | (inputs[688]);
    assign layer0_outputs[3942] = ~((inputs[160]) ^ (inputs[611]));
    assign layer0_outputs[3943] = ~(inputs[588]) | (inputs[774]);
    assign layer0_outputs[3944] = ~(inputs[345]);
    assign layer0_outputs[3945] = (inputs[178]) ^ (inputs[788]);
    assign layer0_outputs[3946] = ~((inputs[845]) | (inputs[917]));
    assign layer0_outputs[3947] = (inputs[161]) & ~(inputs[542]);
    assign layer0_outputs[3948] = (inputs[271]) ^ (inputs[657]);
    assign layer0_outputs[3949] = inputs[772];
    assign layer0_outputs[3950] = (inputs[551]) & ~(inputs[902]);
    assign layer0_outputs[3951] = (inputs[335]) ^ (inputs[602]);
    assign layer0_outputs[3952] = ~(inputs[852]) | (inputs[1008]);
    assign layer0_outputs[3953] = (inputs[430]) | (inputs[854]);
    assign layer0_outputs[3954] = inputs[193];
    assign layer0_outputs[3955] = (inputs[63]) ^ (inputs[594]);
    assign layer0_outputs[3956] = inputs[83];
    assign layer0_outputs[3957] = inputs[972];
    assign layer0_outputs[3958] = ~((inputs[74]) & (inputs[225]));
    assign layer0_outputs[3959] = inputs[194];
    assign layer0_outputs[3960] = ~((inputs[1014]) & (inputs[921]));
    assign layer0_outputs[3961] = (inputs[586]) & ~(inputs[948]);
    assign layer0_outputs[3962] = (inputs[800]) | (inputs[847]);
    assign layer0_outputs[3963] = ~(inputs[251]);
    assign layer0_outputs[3964] = (inputs[141]) | (inputs[841]);
    assign layer0_outputs[3965] = ~((inputs[140]) | (inputs[862]));
    assign layer0_outputs[3966] = ~((inputs[939]) ^ (inputs[961]));
    assign layer0_outputs[3967] = (inputs[792]) | (inputs[649]);
    assign layer0_outputs[3968] = inputs[909];
    assign layer0_outputs[3969] = ~((inputs[417]) & (inputs[258]));
    assign layer0_outputs[3970] = ~(inputs[490]) | (inputs[324]);
    assign layer0_outputs[3971] = ~((inputs[773]) | (inputs[267]));
    assign layer0_outputs[3972] = inputs[346];
    assign layer0_outputs[3973] = inputs[941];
    assign layer0_outputs[3974] = ~((inputs[967]) | (inputs[174]));
    assign layer0_outputs[3975] = ~((inputs[95]) ^ (inputs[314]));
    assign layer0_outputs[3976] = ~(inputs[565]) | (inputs[977]);
    assign layer0_outputs[3977] = ~((inputs[106]) | (inputs[855]));
    assign layer0_outputs[3978] = ~((inputs[405]) | (inputs[189]));
    assign layer0_outputs[3979] = ~((inputs[646]) | (inputs[304]));
    assign layer0_outputs[3980] = ~((inputs[288]) & (inputs[982]));
    assign layer0_outputs[3981] = (inputs[841]) | (inputs[1010]);
    assign layer0_outputs[3982] = ~(inputs[770]);
    assign layer0_outputs[3983] = ~(inputs[937]);
    assign layer0_outputs[3984] = (inputs[435]) ^ (inputs[78]);
    assign layer0_outputs[3985] = inputs[497];
    assign layer0_outputs[3986] = ~((inputs[329]) ^ (inputs[952]));
    assign layer0_outputs[3987] = ~(inputs[789]) | (inputs[84]);
    assign layer0_outputs[3988] = ~(inputs[799]);
    assign layer0_outputs[3989] = ~(inputs[713]);
    assign layer0_outputs[3990] = (inputs[737]) ^ (inputs[277]);
    assign layer0_outputs[3991] = inputs[341];
    assign layer0_outputs[3992] = ~((inputs[4]) ^ (inputs[347]));
    assign layer0_outputs[3993] = ~((inputs[271]) ^ (inputs[676]));
    assign layer0_outputs[3994] = inputs[839];
    assign layer0_outputs[3995] = inputs[588];
    assign layer0_outputs[3996] = (inputs[466]) & ~(inputs[217]);
    assign layer0_outputs[3997] = ~(inputs[596]);
    assign layer0_outputs[3998] = (inputs[89]) & ~(inputs[386]);
    assign layer0_outputs[3999] = (inputs[207]) & ~(inputs[484]);
    assign layer0_outputs[4000] = ~((inputs[172]) ^ (inputs[269]));
    assign layer0_outputs[4001] = ~(inputs[112]);
    assign layer0_outputs[4002] = ~(inputs[741]) | (inputs[930]);
    assign layer0_outputs[4003] = ~((inputs[536]) ^ (inputs[967]));
    assign layer0_outputs[4004] = (inputs[646]) & (inputs[108]);
    assign layer0_outputs[4005] = (inputs[981]) & ~(inputs[232]);
    assign layer0_outputs[4006] = ~((inputs[154]) | (inputs[798]));
    assign layer0_outputs[4007] = (inputs[478]) | (inputs[339]);
    assign layer0_outputs[4008] = (inputs[667]) ^ (inputs[296]);
    assign layer0_outputs[4009] = ~(inputs[349]);
    assign layer0_outputs[4010] = (inputs[254]) ^ (inputs[743]);
    assign layer0_outputs[4011] = ~((inputs[918]) | (inputs[568]));
    assign layer0_outputs[4012] = (inputs[331]) | (inputs[638]);
    assign layer0_outputs[4013] = ~(inputs[405]);
    assign layer0_outputs[4014] = ~(inputs[757]) | (inputs[515]);
    assign layer0_outputs[4015] = (inputs[409]) & ~(inputs[109]);
    assign layer0_outputs[4016] = ~((inputs[208]) | (inputs[765]));
    assign layer0_outputs[4017] = ~(inputs[114]) | (inputs[950]);
    assign layer0_outputs[4018] = ~((inputs[889]) & (inputs[88]));
    assign layer0_outputs[4019] = ~((inputs[637]) | (inputs[766]));
    assign layer0_outputs[4020] = (inputs[488]) | (inputs[216]);
    assign layer0_outputs[4021] = inputs[300];
    assign layer0_outputs[4022] = (inputs[8]) ^ (inputs[178]);
    assign layer0_outputs[4023] = (inputs[47]) | (inputs[468]);
    assign layer0_outputs[4024] = (inputs[765]) | (inputs[364]);
    assign layer0_outputs[4025] = ~(inputs[396]) | (inputs[27]);
    assign layer0_outputs[4026] = (inputs[975]) ^ (inputs[1005]);
    assign layer0_outputs[4027] = ~(inputs[242]);
    assign layer0_outputs[4028] = 1'b0;
    assign layer0_outputs[4029] = inputs[909];
    assign layer0_outputs[4030] = ~(inputs[836]) | (inputs[184]);
    assign layer0_outputs[4031] = ~((inputs[152]) ^ (inputs[513]));
    assign layer0_outputs[4032] = ~((inputs[102]) & (inputs[982]));
    assign layer0_outputs[4033] = ~(inputs[401]);
    assign layer0_outputs[4034] = inputs[843];
    assign layer0_outputs[4035] = (inputs[270]) & ~(inputs[796]);
    assign layer0_outputs[4036] = 1'b0;
    assign layer0_outputs[4037] = ~((inputs[704]) | (inputs[578]));
    assign layer0_outputs[4038] = inputs[424];
    assign layer0_outputs[4039] = ~(inputs[282]);
    assign layer0_outputs[4040] = ~((inputs[49]) ^ (inputs[329]));
    assign layer0_outputs[4041] = ~((inputs[269]) | (inputs[432]));
    assign layer0_outputs[4042] = ~((inputs[783]) | (inputs[30]));
    assign layer0_outputs[4043] = ~((inputs[675]) ^ (inputs[872]));
    assign layer0_outputs[4044] = ~(inputs[251]);
    assign layer0_outputs[4045] = (inputs[723]) & ~(inputs[975]);
    assign layer0_outputs[4046] = (inputs[487]) | (inputs[108]);
    assign layer0_outputs[4047] = (inputs[422]) | (inputs[293]);
    assign layer0_outputs[4048] = (inputs[620]) ^ (inputs[705]);
    assign layer0_outputs[4049] = (inputs[567]) & (inputs[489]);
    assign layer0_outputs[4050] = (inputs[122]) ^ (inputs[904]);
    assign layer0_outputs[4051] = ~((inputs[361]) ^ (inputs[554]));
    assign layer0_outputs[4052] = (inputs[251]) & ~(inputs[485]);
    assign layer0_outputs[4053] = (inputs[107]) | (inputs[569]);
    assign layer0_outputs[4054] = 1'b0;
    assign layer0_outputs[4055] = inputs[283];
    assign layer0_outputs[4056] = (inputs[952]) | (inputs[488]);
    assign layer0_outputs[4057] = ~(inputs[815]);
    assign layer0_outputs[4058] = (inputs[984]) & (inputs[155]);
    assign layer0_outputs[4059] = inputs[711];
    assign layer0_outputs[4060] = ~(inputs[982]) | (inputs[639]);
    assign layer0_outputs[4061] = (inputs[677]) & ~(inputs[122]);
    assign layer0_outputs[4062] = (inputs[713]) & ~(inputs[629]);
    assign layer0_outputs[4063] = (inputs[706]) ^ (inputs[389]);
    assign layer0_outputs[4064] = ~((inputs[562]) | (inputs[120]));
    assign layer0_outputs[4065] = ~(inputs[134]) | (inputs[738]);
    assign layer0_outputs[4066] = ~(inputs[175]) | (inputs[256]);
    assign layer0_outputs[4067] = ~((inputs[167]) ^ (inputs[51]));
    assign layer0_outputs[4068] = (inputs[867]) ^ (inputs[586]);
    assign layer0_outputs[4069] = ~(inputs[697]);
    assign layer0_outputs[4070] = ~(inputs[522]) | (inputs[54]);
    assign layer0_outputs[4071] = (inputs[890]) | (inputs[504]);
    assign layer0_outputs[4072] = ~(inputs[648]);
    assign layer0_outputs[4073] = (inputs[582]) | (inputs[921]);
    assign layer0_outputs[4074] = (inputs[915]) & ~(inputs[218]);
    assign layer0_outputs[4075] = ~(inputs[407]);
    assign layer0_outputs[4076] = ~(inputs[518]);
    assign layer0_outputs[4077] = ~((inputs[77]) | (inputs[426]));
    assign layer0_outputs[4078] = (inputs[696]) | (inputs[458]);
    assign layer0_outputs[4079] = (inputs[187]) ^ (inputs[449]);
    assign layer0_outputs[4080] = ~(inputs[1013]);
    assign layer0_outputs[4081] = (inputs[674]) & ~(inputs[544]);
    assign layer0_outputs[4082] = ~((inputs[116]) ^ (inputs[123]));
    assign layer0_outputs[4083] = ~((inputs[466]) | (inputs[382]));
    assign layer0_outputs[4084] = ~((inputs[539]) | (inputs[833]));
    assign layer0_outputs[4085] = ~(inputs[944]) | (inputs[286]);
    assign layer0_outputs[4086] = ~((inputs[42]) ^ (inputs[313]));
    assign layer0_outputs[4087] = (inputs[572]) & ~(inputs[997]);
    assign layer0_outputs[4088] = ~((inputs[339]) ^ (inputs[329]));
    assign layer0_outputs[4089] = ~(inputs[690]);
    assign layer0_outputs[4090] = ~(inputs[458]) | (inputs[782]);
    assign layer0_outputs[4091] = ~(inputs[771]) | (inputs[1020]);
    assign layer0_outputs[4092] = ~((inputs[694]) & (inputs[601]));
    assign layer0_outputs[4093] = (inputs[287]) | (inputs[631]);
    assign layer0_outputs[4094] = (inputs[193]) | (inputs[702]);
    assign layer0_outputs[4095] = ~((inputs[52]) | (inputs[290]));
    assign layer0_outputs[4096] = (inputs[255]) | (inputs[660]);
    assign layer0_outputs[4097] = ~((inputs[754]) | (inputs[976]));
    assign layer0_outputs[4098] = inputs[159];
    assign layer0_outputs[4099] = (inputs[88]) ^ (inputs[281]);
    assign layer0_outputs[4100] = ~(inputs[949]) | (inputs[383]);
    assign layer0_outputs[4101] = ~((inputs[643]) ^ (inputs[912]));
    assign layer0_outputs[4102] = inputs[265];
    assign layer0_outputs[4103] = ~((inputs[393]) ^ (inputs[648]));
    assign layer0_outputs[4104] = ~(inputs[493]);
    assign layer0_outputs[4105] = inputs[441];
    assign layer0_outputs[4106] = (inputs[775]) & ~(inputs[705]);
    assign layer0_outputs[4107] = (inputs[316]) | (inputs[698]);
    assign layer0_outputs[4108] = ~(inputs[302]);
    assign layer0_outputs[4109] = ~(inputs[783]) | (inputs[218]);
    assign layer0_outputs[4110] = ~(inputs[938]);
    assign layer0_outputs[4111] = inputs[590];
    assign layer0_outputs[4112] = ~(inputs[524]);
    assign layer0_outputs[4113] = ~(inputs[297]) | (inputs[771]);
    assign layer0_outputs[4114] = inputs[714];
    assign layer0_outputs[4115] = ~(inputs[498]) | (inputs[179]);
    assign layer0_outputs[4116] = (inputs[904]) | (inputs[151]);
    assign layer0_outputs[4117] = inputs[31];
    assign layer0_outputs[4118] = (inputs[538]) ^ (inputs[477]);
    assign layer0_outputs[4119] = (inputs[525]) | (inputs[544]);
    assign layer0_outputs[4120] = ~(inputs[645]);
    assign layer0_outputs[4121] = ~((inputs[455]) | (inputs[572]));
    assign layer0_outputs[4122] = 1'b1;
    assign layer0_outputs[4123] = ~(inputs[677]) | (inputs[858]);
    assign layer0_outputs[4124] = ~((inputs[739]) ^ (inputs[19]));
    assign layer0_outputs[4125] = ~((inputs[974]) & (inputs[711]));
    assign layer0_outputs[4126] = ~((inputs[539]) | (inputs[288]));
    assign layer0_outputs[4127] = (inputs[745]) | (inputs[755]);
    assign layer0_outputs[4128] = (inputs[373]) ^ (inputs[391]);
    assign layer0_outputs[4129] = (inputs[1017]) ^ (inputs[476]);
    assign layer0_outputs[4130] = ~(inputs[503]);
    assign layer0_outputs[4131] = inputs[425];
    assign layer0_outputs[4132] = (inputs[570]) ^ (inputs[264]);
    assign layer0_outputs[4133] = ~((inputs[809]) | (inputs[894]));
    assign layer0_outputs[4134] = (inputs[693]) & ~(inputs[97]);
    assign layer0_outputs[4135] = ~((inputs[165]) | (inputs[614]));
    assign layer0_outputs[4136] = 1'b0;
    assign layer0_outputs[4137] = (inputs[305]) & ~(inputs[693]);
    assign layer0_outputs[4138] = (inputs[777]) & ~(inputs[470]);
    assign layer0_outputs[4139] = (inputs[505]) ^ (inputs[194]);
    assign layer0_outputs[4140] = inputs[395];
    assign layer0_outputs[4141] = ~((inputs[399]) | (inputs[350]));
    assign layer0_outputs[4142] = ~(inputs[528]);
    assign layer0_outputs[4143] = ~((inputs[541]) | (inputs[272]));
    assign layer0_outputs[4144] = (inputs[395]) & ~(inputs[281]);
    assign layer0_outputs[4145] = (inputs[699]) & ~(inputs[908]);
    assign layer0_outputs[4146] = (inputs[475]) & ~(inputs[199]);
    assign layer0_outputs[4147] = ~((inputs[635]) | (inputs[921]));
    assign layer0_outputs[4148] = (inputs[842]) ^ (inputs[96]);
    assign layer0_outputs[4149] = (inputs[3]) | (inputs[846]);
    assign layer0_outputs[4150] = ~((inputs[947]) | (inputs[907]));
    assign layer0_outputs[4151] = (inputs[685]) & ~(inputs[581]);
    assign layer0_outputs[4152] = ~(inputs[536]);
    assign layer0_outputs[4153] = (inputs[721]) & ~(inputs[326]);
    assign layer0_outputs[4154] = inputs[747];
    assign layer0_outputs[4155] = (inputs[903]) & ~(inputs[223]);
    assign layer0_outputs[4156] = ~(inputs[516]);
    assign layer0_outputs[4157] = ~(inputs[857]) | (inputs[973]);
    assign layer0_outputs[4158] = ~(inputs[923]) | (inputs[892]);
    assign layer0_outputs[4159] = (inputs[578]) ^ (inputs[976]);
    assign layer0_outputs[4160] = (inputs[877]) | (inputs[977]);
    assign layer0_outputs[4161] = (inputs[501]) & ~(inputs[184]);
    assign layer0_outputs[4162] = (inputs[71]) & (inputs[783]);
    assign layer0_outputs[4163] = (inputs[858]) ^ (inputs[350]);
    assign layer0_outputs[4164] = ~((inputs[272]) | (inputs[743]));
    assign layer0_outputs[4165] = (inputs[339]) | (inputs[263]);
    assign layer0_outputs[4166] = (inputs[283]) & ~(inputs[475]);
    assign layer0_outputs[4167] = ~(inputs[585]);
    assign layer0_outputs[4168] = ~((inputs[271]) | (inputs[191]));
    assign layer0_outputs[4169] = ~(inputs[333]);
    assign layer0_outputs[4170] = ~((inputs[588]) | (inputs[231]));
    assign layer0_outputs[4171] = (inputs[232]) | (inputs[812]);
    assign layer0_outputs[4172] = ~(inputs[377]);
    assign layer0_outputs[4173] = ~((inputs[914]) & (inputs[128]));
    assign layer0_outputs[4174] = ~(inputs[383]);
    assign layer0_outputs[4175] = (inputs[789]) ^ (inputs[256]);
    assign layer0_outputs[4176] = (inputs[609]) | (inputs[602]);
    assign layer0_outputs[4177] = ~((inputs[712]) ^ (inputs[705]));
    assign layer0_outputs[4178] = (inputs[439]) & ~(inputs[95]);
    assign layer0_outputs[4179] = 1'b1;
    assign layer0_outputs[4180] = ~((inputs[801]) ^ (inputs[896]));
    assign layer0_outputs[4181] = ~((inputs[369]) ^ (inputs[238]));
    assign layer0_outputs[4182] = ~(inputs[679]);
    assign layer0_outputs[4183] = ~((inputs[999]) ^ (inputs[127]));
    assign layer0_outputs[4184] = ~(inputs[697]);
    assign layer0_outputs[4185] = ~((inputs[112]) | (inputs[151]));
    assign layer0_outputs[4186] = (inputs[8]) & (inputs[806]);
    assign layer0_outputs[4187] = ~((inputs[151]) | (inputs[717]));
    assign layer0_outputs[4188] = 1'b1;
    assign layer0_outputs[4189] = ~((inputs[495]) ^ (inputs[24]));
    assign layer0_outputs[4190] = ~(inputs[282]);
    assign layer0_outputs[4191] = (inputs[72]) ^ (inputs[768]);
    assign layer0_outputs[4192] = ~(inputs[305]) | (inputs[133]);
    assign layer0_outputs[4193] = (inputs[102]) | (inputs[677]);
    assign layer0_outputs[4194] = (inputs[837]) & (inputs[164]);
    assign layer0_outputs[4195] = ~((inputs[161]) ^ (inputs[529]));
    assign layer0_outputs[4196] = (inputs[258]) & ~(inputs[971]);
    assign layer0_outputs[4197] = 1'b0;
    assign layer0_outputs[4198] = inputs[196];
    assign layer0_outputs[4199] = ~(inputs[556]);
    assign layer0_outputs[4200] = ~((inputs[755]) ^ (inputs[766]));
    assign layer0_outputs[4201] = ~((inputs[274]) ^ (inputs[987]));
    assign layer0_outputs[4202] = ~(inputs[14]);
    assign layer0_outputs[4203] = ~((inputs[22]) ^ (inputs[255]));
    assign layer0_outputs[4204] = (inputs[688]) | (inputs[974]);
    assign layer0_outputs[4205] = ~((inputs[980]) | (inputs[907]));
    assign layer0_outputs[4206] = ~((inputs[335]) | (inputs[120]));
    assign layer0_outputs[4207] = inputs[555];
    assign layer0_outputs[4208] = (inputs[87]) & (inputs[421]);
    assign layer0_outputs[4209] = ~((inputs[377]) | (inputs[331]));
    assign layer0_outputs[4210] = inputs[912];
    assign layer0_outputs[4211] = ~((inputs[966]) | (inputs[878]));
    assign layer0_outputs[4212] = (inputs[245]) & (inputs[281]);
    assign layer0_outputs[4213] = ~(inputs[140]);
    assign layer0_outputs[4214] = (inputs[776]) | (inputs[91]);
    assign layer0_outputs[4215] = ~((inputs[976]) | (inputs[402]));
    assign layer0_outputs[4216] = (inputs[242]) & ~(inputs[9]);
    assign layer0_outputs[4217] = (inputs[303]) & ~(inputs[902]);
    assign layer0_outputs[4218] = 1'b0;
    assign layer0_outputs[4219] = ~((inputs[28]) ^ (inputs[569]));
    assign layer0_outputs[4220] = (inputs[793]) & ~(inputs[284]);
    assign layer0_outputs[4221] = ~((inputs[1020]) | (inputs[622]));
    assign layer0_outputs[4222] = ~(inputs[656]);
    assign layer0_outputs[4223] = inputs[360];
    assign layer0_outputs[4224] = ~((inputs[610]) & (inputs[362]));
    assign layer0_outputs[4225] = (inputs[958]) & ~(inputs[33]);
    assign layer0_outputs[4226] = (inputs[365]) & ~(inputs[202]);
    assign layer0_outputs[4227] = (inputs[331]) & ~(inputs[122]);
    assign layer0_outputs[4228] = inputs[877];
    assign layer0_outputs[4229] = ~(inputs[477]) | (inputs[92]);
    assign layer0_outputs[4230] = (inputs[216]) & (inputs[200]);
    assign layer0_outputs[4231] = ~((inputs[351]) | (inputs[243]));
    assign layer0_outputs[4232] = 1'b0;
    assign layer0_outputs[4233] = ~(inputs[657]) | (inputs[632]);
    assign layer0_outputs[4234] = (inputs[133]) | (inputs[743]);
    assign layer0_outputs[4235] = (inputs[682]) | (inputs[573]);
    assign layer0_outputs[4236] = (inputs[194]) ^ (inputs[617]);
    assign layer0_outputs[4237] = (inputs[714]) & ~(inputs[435]);
    assign layer0_outputs[4238] = ~((inputs[275]) | (inputs[310]));
    assign layer0_outputs[4239] = ~(inputs[273]);
    assign layer0_outputs[4240] = ~(inputs[920]);
    assign layer0_outputs[4241] = ~((inputs[267]) ^ (inputs[726]));
    assign layer0_outputs[4242] = (inputs[546]) ^ (inputs[750]);
    assign layer0_outputs[4243] = (inputs[623]) ^ (inputs[580]);
    assign layer0_outputs[4244] = ~(inputs[810]);
    assign layer0_outputs[4245] = ~(inputs[650]);
    assign layer0_outputs[4246] = ~((inputs[852]) | (inputs[249]));
    assign layer0_outputs[4247] = (inputs[374]) | (inputs[373]);
    assign layer0_outputs[4248] = ~((inputs[739]) & (inputs[100]));
    assign layer0_outputs[4249] = (inputs[114]) & ~(inputs[541]);
    assign layer0_outputs[4250] = ~(inputs[492]);
    assign layer0_outputs[4251] = (inputs[274]) | (inputs[732]);
    assign layer0_outputs[4252] = (inputs[555]) & ~(inputs[178]);
    assign layer0_outputs[4253] = ~(inputs[699]) | (inputs[265]);
    assign layer0_outputs[4254] = ~((inputs[98]) ^ (inputs[628]));
    assign layer0_outputs[4255] = 1'b0;
    assign layer0_outputs[4256] = (inputs[310]) ^ (inputs[700]);
    assign layer0_outputs[4257] = ~(inputs[194]) | (inputs[978]);
    assign layer0_outputs[4258] = inputs[560];
    assign layer0_outputs[4259] = inputs[681];
    assign layer0_outputs[4260] = ~(inputs[501]);
    assign layer0_outputs[4261] = inputs[468];
    assign layer0_outputs[4262] = ~(inputs[692]) | (inputs[370]);
    assign layer0_outputs[4263] = (inputs[520]) & ~(inputs[163]);
    assign layer0_outputs[4264] = ~(inputs[269]) | (inputs[1004]);
    assign layer0_outputs[4265] = ~((inputs[83]) ^ (inputs[675]));
    assign layer0_outputs[4266] = ~((inputs[343]) | (inputs[368]));
    assign layer0_outputs[4267] = ~(inputs[715]) | (inputs[934]);
    assign layer0_outputs[4268] = inputs[148];
    assign layer0_outputs[4269] = (inputs[557]) & ~(inputs[670]);
    assign layer0_outputs[4270] = ~((inputs[931]) | (inputs[324]));
    assign layer0_outputs[4271] = (inputs[963]) & ~(inputs[294]);
    assign layer0_outputs[4272] = (inputs[844]) & ~(inputs[75]);
    assign layer0_outputs[4273] = (inputs[495]) & ~(inputs[388]);
    assign layer0_outputs[4274] = (inputs[293]) ^ (inputs[546]);
    assign layer0_outputs[4275] = ~((inputs[381]) | (inputs[814]));
    assign layer0_outputs[4276] = ~((inputs[623]) | (inputs[225]));
    assign layer0_outputs[4277] = ~(inputs[401]);
    assign layer0_outputs[4278] = inputs[754];
    assign layer0_outputs[4279] = inputs[55];
    assign layer0_outputs[4280] = ~(inputs[129]);
    assign layer0_outputs[4281] = ~((inputs[505]) | (inputs[555]));
    assign layer0_outputs[4282] = (inputs[910]) | (inputs[214]);
    assign layer0_outputs[4283] = inputs[293];
    assign layer0_outputs[4284] = ~(inputs[338]);
    assign layer0_outputs[4285] = (inputs[755]) & ~(inputs[641]);
    assign layer0_outputs[4286] = ~((inputs[31]) & (inputs[510]));
    assign layer0_outputs[4287] = (inputs[486]) & ~(inputs[233]);
    assign layer0_outputs[4288] = inputs[520];
    assign layer0_outputs[4289] = (inputs[853]) & ~(inputs[41]);
    assign layer0_outputs[4290] = (inputs[1020]) & ~(inputs[932]);
    assign layer0_outputs[4291] = inputs[84];
    assign layer0_outputs[4292] = (inputs[935]) & ~(inputs[151]);
    assign layer0_outputs[4293] = inputs[557];
    assign layer0_outputs[4294] = 1'b0;
    assign layer0_outputs[4295] = (inputs[554]) & ~(inputs[199]);
    assign layer0_outputs[4296] = ~((inputs[42]) | (inputs[111]));
    assign layer0_outputs[4297] = ~((inputs[465]) | (inputs[943]));
    assign layer0_outputs[4298] = ~(inputs[663]) | (inputs[63]);
    assign layer0_outputs[4299] = ~(inputs[215]) | (inputs[225]);
    assign layer0_outputs[4300] = (inputs[672]) & ~(inputs[896]);
    assign layer0_outputs[4301] = ~(inputs[201]) | (inputs[283]);
    assign layer0_outputs[4302] = (inputs[910]) ^ (inputs[12]);
    assign layer0_outputs[4303] = ~((inputs[694]) | (inputs[295]));
    assign layer0_outputs[4304] = (inputs[405]) | (inputs[104]);
    assign layer0_outputs[4305] = (inputs[904]) & ~(inputs[252]);
    assign layer0_outputs[4306] = ~((inputs[373]) | (inputs[709]));
    assign layer0_outputs[4307] = ~(inputs[86]) | (inputs[327]);
    assign layer0_outputs[4308] = ~((inputs[367]) | (inputs[864]));
    assign layer0_outputs[4309] = ~(inputs[964]) | (inputs[1020]);
    assign layer0_outputs[4310] = (inputs[402]) | (inputs[965]);
    assign layer0_outputs[4311] = 1'b0;
    assign layer0_outputs[4312] = ~((inputs[116]) | (inputs[30]));
    assign layer0_outputs[4313] = ~(inputs[246]);
    assign layer0_outputs[4314] = ~(inputs[110]);
    assign layer0_outputs[4315] = (inputs[423]) & ~(inputs[954]);
    assign layer0_outputs[4316] = inputs[266];
    assign layer0_outputs[4317] = (inputs[779]) ^ (inputs[910]);
    assign layer0_outputs[4318] = (inputs[162]) | (inputs[523]);
    assign layer0_outputs[4319] = ~(inputs[37]);
    assign layer0_outputs[4320] = (inputs[525]) & ~(inputs[336]);
    assign layer0_outputs[4321] = inputs[690];
    assign layer0_outputs[4322] = ~((inputs[254]) ^ (inputs[450]));
    assign layer0_outputs[4323] = (inputs[960]) ^ (inputs[476]);
    assign layer0_outputs[4324] = ~(inputs[82]);
    assign layer0_outputs[4325] = (inputs[62]) & (inputs[22]);
    assign layer0_outputs[4326] = ~(inputs[980]);
    assign layer0_outputs[4327] = (inputs[662]) ^ (inputs[702]);
    assign layer0_outputs[4328] = ~(inputs[320]) | (inputs[174]);
    assign layer0_outputs[4329] = ~((inputs[855]) | (inputs[712]));
    assign layer0_outputs[4330] = inputs[819];
    assign layer0_outputs[4331] = (inputs[174]) & ~(inputs[261]);
    assign layer0_outputs[4332] = ~((inputs[850]) & (inputs[332]));
    assign layer0_outputs[4333] = ~((inputs[920]) | (inputs[557]));
    assign layer0_outputs[4334] = ~((inputs[346]) | (inputs[207]));
    assign layer0_outputs[4335] = inputs[493];
    assign layer0_outputs[4336] = ~((inputs[411]) | (inputs[665]));
    assign layer0_outputs[4337] = inputs[493];
    assign layer0_outputs[4338] = inputs[143];
    assign layer0_outputs[4339] = ~((inputs[628]) ^ (inputs[787]));
    assign layer0_outputs[4340] = ~(inputs[340]) | (inputs[984]);
    assign layer0_outputs[4341] = inputs[840];
    assign layer0_outputs[4342] = ~((inputs[492]) | (inputs[679]));
    assign layer0_outputs[4343] = ~(inputs[205]);
    assign layer0_outputs[4344] = ~((inputs[217]) | (inputs[975]));
    assign layer0_outputs[4345] = ~(inputs[42]) | (inputs[57]);
    assign layer0_outputs[4346] = inputs[203];
    assign layer0_outputs[4347] = ~(inputs[703]) | (inputs[18]);
    assign layer0_outputs[4348] = (inputs[399]) ^ (inputs[134]);
    assign layer0_outputs[4349] = (inputs[961]) ^ (inputs[695]);
    assign layer0_outputs[4350] = ~(inputs[275]) | (inputs[779]);
    assign layer0_outputs[4351] = (inputs[341]) ^ (inputs[215]);
    assign layer0_outputs[4352] = ~(inputs[698]);
    assign layer0_outputs[4353] = ~(inputs[163]) | (inputs[666]);
    assign layer0_outputs[4354] = inputs[78];
    assign layer0_outputs[4355] = ~(inputs[583]) | (inputs[345]);
    assign layer0_outputs[4356] = (inputs[757]) ^ (inputs[274]);
    assign layer0_outputs[4357] = inputs[112];
    assign layer0_outputs[4358] = ~((inputs[149]) ^ (inputs[750]));
    assign layer0_outputs[4359] = ~(inputs[744]) | (inputs[550]);
    assign layer0_outputs[4360] = ~((inputs[906]) | (inputs[116]));
    assign layer0_outputs[4361] = ~((inputs[802]) | (inputs[656]));
    assign layer0_outputs[4362] = ~(inputs[303]) | (inputs[524]);
    assign layer0_outputs[4363] = inputs[1006];
    assign layer0_outputs[4364] = ~(inputs[571]) | (inputs[517]);
    assign layer0_outputs[4365] = ~(inputs[1018]) | (inputs[75]);
    assign layer0_outputs[4366] = (inputs[349]) | (inputs[790]);
    assign layer0_outputs[4367] = (inputs[798]) ^ (inputs[600]);
    assign layer0_outputs[4368] = (inputs[831]) & ~(inputs[81]);
    assign layer0_outputs[4369] = ~((inputs[402]) | (inputs[564]));
    assign layer0_outputs[4370] = ~(inputs[844]) | (inputs[419]);
    assign layer0_outputs[4371] = (inputs[79]) & ~(inputs[869]);
    assign layer0_outputs[4372] = inputs[438];
    assign layer0_outputs[4373] = ~((inputs[165]) | (inputs[404]));
    assign layer0_outputs[4374] = ~(inputs[424]) | (inputs[382]);
    assign layer0_outputs[4375] = ~(inputs[711]) | (inputs[904]);
    assign layer0_outputs[4376] = ~(inputs[390]);
    assign layer0_outputs[4377] = inputs[578];
    assign layer0_outputs[4378] = inputs[63];
    assign layer0_outputs[4379] = (inputs[203]) | (inputs[292]);
    assign layer0_outputs[4380] = ~(inputs[881]);
    assign layer0_outputs[4381] = (inputs[523]) & ~(inputs[45]);
    assign layer0_outputs[4382] = 1'b1;
    assign layer0_outputs[4383] = ~((inputs[510]) ^ (inputs[23]));
    assign layer0_outputs[4384] = ~((inputs[568]) | (inputs[598]));
    assign layer0_outputs[4385] = inputs[69];
    assign layer0_outputs[4386] = (inputs[471]) & ~(inputs[963]);
    assign layer0_outputs[4387] = ~((inputs[505]) | (inputs[101]));
    assign layer0_outputs[4388] = ~((inputs[947]) | (inputs[376]));
    assign layer0_outputs[4389] = ~((inputs[809]) | (inputs[238]));
    assign layer0_outputs[4390] = ~(inputs[425]);
    assign layer0_outputs[4391] = inputs[113];
    assign layer0_outputs[4392] = (inputs[809]) | (inputs[839]);
    assign layer0_outputs[4393] = inputs[179];
    assign layer0_outputs[4394] = ~(inputs[746]);
    assign layer0_outputs[4395] = ~((inputs[207]) | (inputs[969]));
    assign layer0_outputs[4396] = ~(inputs[721]);
    assign layer0_outputs[4397] = 1'b1;
    assign layer0_outputs[4398] = ~(inputs[374]);
    assign layer0_outputs[4399] = (inputs[529]) & ~(inputs[773]);
    assign layer0_outputs[4400] = inputs[244];
    assign layer0_outputs[4401] = (inputs[284]) & ~(inputs[70]);
    assign layer0_outputs[4402] = (inputs[852]) | (inputs[747]);
    assign layer0_outputs[4403] = (inputs[674]) | (inputs[405]);
    assign layer0_outputs[4404] = (inputs[670]) ^ (inputs[540]);
    assign layer0_outputs[4405] = ~(inputs[425]);
    assign layer0_outputs[4406] = inputs[682];
    assign layer0_outputs[4407] = ~(inputs[36]);
    assign layer0_outputs[4408] = ~(inputs[307]);
    assign layer0_outputs[4409] = inputs[695];
    assign layer0_outputs[4410] = (inputs[58]) & ~(inputs[987]);
    assign layer0_outputs[4411] = (inputs[623]) & ~(inputs[51]);
    assign layer0_outputs[4412] = ~(inputs[964]) | (inputs[67]);
    assign layer0_outputs[4413] = ~((inputs[938]) ^ (inputs[1012]));
    assign layer0_outputs[4414] = ~((inputs[839]) ^ (inputs[338]));
    assign layer0_outputs[4415] = ~(inputs[119]);
    assign layer0_outputs[4416] = ~(inputs[429]) | (inputs[600]);
    assign layer0_outputs[4417] = 1'b1;
    assign layer0_outputs[4418] = (inputs[434]) | (inputs[644]);
    assign layer0_outputs[4419] = ~((inputs[842]) | (inputs[729]));
    assign layer0_outputs[4420] = (inputs[188]) | (inputs[19]);
    assign layer0_outputs[4421] = ~((inputs[336]) ^ (inputs[359]));
    assign layer0_outputs[4422] = inputs[731];
    assign layer0_outputs[4423] = ~((inputs[150]) ^ (inputs[500]));
    assign layer0_outputs[4424] = ~(inputs[655]);
    assign layer0_outputs[4425] = ~(inputs[470]);
    assign layer0_outputs[4426] = 1'b0;
    assign layer0_outputs[4427] = ~(inputs[890]) | (inputs[1021]);
    assign layer0_outputs[4428] = ~(inputs[560]) | (inputs[163]);
    assign layer0_outputs[4429] = (inputs[906]) | (inputs[403]);
    assign layer0_outputs[4430] = ~(inputs[765]) | (inputs[135]);
    assign layer0_outputs[4431] = (inputs[887]) & (inputs[73]);
    assign layer0_outputs[4432] = ~(inputs[661]) | (inputs[577]);
    assign layer0_outputs[4433] = inputs[297];
    assign layer0_outputs[4434] = ~((inputs[1012]) | (inputs[866]));
    assign layer0_outputs[4435] = ~(inputs[626]);
    assign layer0_outputs[4436] = (inputs[789]) | (inputs[328]);
    assign layer0_outputs[4437] = inputs[397];
    assign layer0_outputs[4438] = (inputs[507]) | (inputs[419]);
    assign layer0_outputs[4439] = ~(inputs[531]);
    assign layer0_outputs[4440] = ~((inputs[822]) ^ (inputs[98]));
    assign layer0_outputs[4441] = 1'b0;
    assign layer0_outputs[4442] = (inputs[602]) | (inputs[803]);
    assign layer0_outputs[4443] = ~(inputs[375]);
    assign layer0_outputs[4444] = ~((inputs[779]) | (inputs[830]));
    assign layer0_outputs[4445] = (inputs[840]) | (inputs[987]);
    assign layer0_outputs[4446] = inputs[763];
    assign layer0_outputs[4447] = ~((inputs[599]) ^ (inputs[202]));
    assign layer0_outputs[4448] = ~((inputs[368]) | (inputs[22]));
    assign layer0_outputs[4449] = inputs[169];
    assign layer0_outputs[4450] = (inputs[88]) | (inputs[461]);
    assign layer0_outputs[4451] = ~(inputs[425]);
    assign layer0_outputs[4452] = (inputs[301]) & ~(inputs[866]);
    assign layer0_outputs[4453] = (inputs[901]) & (inputs[947]);
    assign layer0_outputs[4454] = (inputs[828]) ^ (inputs[800]);
    assign layer0_outputs[4455] = ~(inputs[214]);
    assign layer0_outputs[4456] = ~(inputs[491]) | (inputs[99]);
    assign layer0_outputs[4457] = ~(inputs[757]);
    assign layer0_outputs[4458] = ~(inputs[870]) | (inputs[554]);
    assign layer0_outputs[4459] = (inputs[292]) ^ (inputs[953]);
    assign layer0_outputs[4460] = ~(inputs[577]);
    assign layer0_outputs[4461] = ~((inputs[79]) | (inputs[377]));
    assign layer0_outputs[4462] = 1'b0;
    assign layer0_outputs[4463] = ~((inputs[536]) | (inputs[34]));
    assign layer0_outputs[4464] = (inputs[964]) & (inputs[1015]);
    assign layer0_outputs[4465] = ~((inputs[366]) ^ (inputs[867]));
    assign layer0_outputs[4466] = inputs[463];
    assign layer0_outputs[4467] = (inputs[467]) & ~(inputs[746]);
    assign layer0_outputs[4468] = ~(inputs[34]);
    assign layer0_outputs[4469] = (inputs[843]) & ~(inputs[136]);
    assign layer0_outputs[4470] = ~((inputs[374]) & (inputs[240]));
    assign layer0_outputs[4471] = ~(inputs[371]);
    assign layer0_outputs[4472] = inputs[542];
    assign layer0_outputs[4473] = ~(inputs[431]);
    assign layer0_outputs[4474] = (inputs[1009]) & (inputs[702]);
    assign layer0_outputs[4475] = (inputs[537]) | (inputs[721]);
    assign layer0_outputs[4476] = inputs[690];
    assign layer0_outputs[4477] = (inputs[617]) & ~(inputs[641]);
    assign layer0_outputs[4478] = (inputs[305]) & ~(inputs[5]);
    assign layer0_outputs[4479] = ~((inputs[556]) | (inputs[334]));
    assign layer0_outputs[4480] = ~((inputs[931]) | (inputs[779]));
    assign layer0_outputs[4481] = (inputs[997]) & ~(inputs[864]);
    assign layer0_outputs[4482] = (inputs[846]) ^ (inputs[743]);
    assign layer0_outputs[4483] = ~(inputs[310]);
    assign layer0_outputs[4484] = ~(inputs[443]);
    assign layer0_outputs[4485] = (inputs[95]) | (inputs[129]);
    assign layer0_outputs[4486] = (inputs[406]) & (inputs[273]);
    assign layer0_outputs[4487] = ~((inputs[501]) ^ (inputs[732]));
    assign layer0_outputs[4488] = (inputs[1016]) & (inputs[930]);
    assign layer0_outputs[4489] = (inputs[517]) & ~(inputs[936]);
    assign layer0_outputs[4490] = ~(inputs[720]) | (inputs[831]);
    assign layer0_outputs[4491] = ~((inputs[449]) | (inputs[671]));
    assign layer0_outputs[4492] = (inputs[533]) | (inputs[789]);
    assign layer0_outputs[4493] = ~((inputs[498]) | (inputs[547]));
    assign layer0_outputs[4494] = ~((inputs[90]) & (inputs[81]));
    assign layer0_outputs[4495] = (inputs[437]) & ~(inputs[519]);
    assign layer0_outputs[4496] = ~(inputs[431]) | (inputs[508]);
    assign layer0_outputs[4497] = ~((inputs[835]) ^ (inputs[367]));
    assign layer0_outputs[4498] = (inputs[766]) & ~(inputs[162]);
    assign layer0_outputs[4499] = ~((inputs[560]) | (inputs[152]));
    assign layer0_outputs[4500] = ~(inputs[376]);
    assign layer0_outputs[4501] = inputs[315];
    assign layer0_outputs[4502] = (inputs[502]) & ~(inputs[573]);
    assign layer0_outputs[4503] = (inputs[758]) & ~(inputs[36]);
    assign layer0_outputs[4504] = ~((inputs[706]) | (inputs[612]));
    assign layer0_outputs[4505] = ~((inputs[847]) ^ (inputs[973]));
    assign layer0_outputs[4506] = (inputs[868]) & ~(inputs[349]);
    assign layer0_outputs[4507] = ~((inputs[709]) | (inputs[214]));
    assign layer0_outputs[4508] = ~(inputs[661]);
    assign layer0_outputs[4509] = (inputs[896]) & ~(inputs[867]);
    assign layer0_outputs[4510] = inputs[626];
    assign layer0_outputs[4511] = ~(inputs[379]);
    assign layer0_outputs[4512] = ~(inputs[741]);
    assign layer0_outputs[4513] = (inputs[475]) | (inputs[630]);
    assign layer0_outputs[4514] = inputs[337];
    assign layer0_outputs[4515] = ~((inputs[664]) | (inputs[644]));
    assign layer0_outputs[4516] = ~(inputs[570]) | (inputs[924]);
    assign layer0_outputs[4517] = inputs[140];
    assign layer0_outputs[4518] = ~((inputs[347]) ^ (inputs[66]));
    assign layer0_outputs[4519] = ~((inputs[574]) | (inputs[294]));
    assign layer0_outputs[4520] = ~(inputs[550]) | (inputs[268]);
    assign layer0_outputs[4521] = ~(inputs[745]) | (inputs[708]);
    assign layer0_outputs[4522] = ~(inputs[179]);
    assign layer0_outputs[4523] = ~(inputs[942]);
    assign layer0_outputs[4524] = (inputs[499]) ^ (inputs[745]);
    assign layer0_outputs[4525] = (inputs[217]) ^ (inputs[956]);
    assign layer0_outputs[4526] = ~((inputs[799]) | (inputs[269]));
    assign layer0_outputs[4527] = ~(inputs[986]) | (inputs[420]);
    assign layer0_outputs[4528] = inputs[665];
    assign layer0_outputs[4529] = (inputs[679]) & (inputs[90]);
    assign layer0_outputs[4530] = ~(inputs[470]);
    assign layer0_outputs[4531] = ~((inputs[562]) | (inputs[947]));
    assign layer0_outputs[4532] = ~(inputs[305]) | (inputs[181]);
    assign layer0_outputs[4533] = (inputs[752]) | (inputs[737]);
    assign layer0_outputs[4534] = (inputs[280]) | (inputs[663]);
    assign layer0_outputs[4535] = (inputs[396]) & ~(inputs[767]);
    assign layer0_outputs[4536] = (inputs[138]) & ~(inputs[991]);
    assign layer0_outputs[4537] = ~(inputs[433]) | (inputs[117]);
    assign layer0_outputs[4538] = ~((inputs[903]) | (inputs[386]));
    assign layer0_outputs[4539] = ~(inputs[715]);
    assign layer0_outputs[4540] = (inputs[562]) & ~(inputs[613]);
    assign layer0_outputs[4541] = inputs[400];
    assign layer0_outputs[4542] = 1'b1;
    assign layer0_outputs[4543] = (inputs[184]) | (inputs[845]);
    assign layer0_outputs[4544] = (inputs[103]) & ~(inputs[837]);
    assign layer0_outputs[4545] = inputs[587];
    assign layer0_outputs[4546] = ~((inputs[741]) & (inputs[738]));
    assign layer0_outputs[4547] = ~((inputs[922]) ^ (inputs[218]));
    assign layer0_outputs[4548] = (inputs[948]) & ~(inputs[176]);
    assign layer0_outputs[4549] = ~(inputs[329]) | (inputs[14]);
    assign layer0_outputs[4550] = inputs[375];
    assign layer0_outputs[4551] = ~(inputs[28]) | (inputs[541]);
    assign layer0_outputs[4552] = (inputs[422]) & ~(inputs[21]);
    assign layer0_outputs[4553] = ~((inputs[1008]) ^ (inputs[298]));
    assign layer0_outputs[4554] = (inputs[293]) ^ (inputs[501]);
    assign layer0_outputs[4555] = ~((inputs[433]) | (inputs[466]));
    assign layer0_outputs[4556] = inputs[495];
    assign layer0_outputs[4557] = ~((inputs[407]) | (inputs[269]));
    assign layer0_outputs[4558] = ~(inputs[403]);
    assign layer0_outputs[4559] = ~(inputs[657]);
    assign layer0_outputs[4560] = (inputs[267]) | (inputs[781]);
    assign layer0_outputs[4561] = (inputs[372]) | (inputs[574]);
    assign layer0_outputs[4562] = ~(inputs[176]);
    assign layer0_outputs[4563] = ~(inputs[715]) | (inputs[96]);
    assign layer0_outputs[4564] = ~(inputs[245]);
    assign layer0_outputs[4565] = inputs[907];
    assign layer0_outputs[4566] = ~(inputs[403]);
    assign layer0_outputs[4567] = ~((inputs[355]) | (inputs[322]));
    assign layer0_outputs[4568] = (inputs[200]) ^ (inputs[265]);
    assign layer0_outputs[4569] = ~((inputs[971]) | (inputs[196]));
    assign layer0_outputs[4570] = ~((inputs[91]) | (inputs[157]));
    assign layer0_outputs[4571] = ~((inputs[991]) | (inputs[317]));
    assign layer0_outputs[4572] = ~((inputs[794]) | (inputs[54]));
    assign layer0_outputs[4573] = ~(inputs[417]) | (inputs[447]);
    assign layer0_outputs[4574] = (inputs[663]) & ~(inputs[859]);
    assign layer0_outputs[4575] = ~((inputs[765]) ^ (inputs[456]));
    assign layer0_outputs[4576] = ~((inputs[397]) | (inputs[21]));
    assign layer0_outputs[4577] = (inputs[29]) & ~(inputs[931]);
    assign layer0_outputs[4578] = 1'b1;
    assign layer0_outputs[4579] = (inputs[996]) | (inputs[683]);
    assign layer0_outputs[4580] = inputs[551];
    assign layer0_outputs[4581] = ~((inputs[710]) | (inputs[105]));
    assign layer0_outputs[4582] = (inputs[149]) | (inputs[694]);
    assign layer0_outputs[4583] = ~(inputs[4]);
    assign layer0_outputs[4584] = (inputs[876]) ^ (inputs[866]);
    assign layer0_outputs[4585] = (inputs[73]) | (inputs[549]);
    assign layer0_outputs[4586] = ~(inputs[811]);
    assign layer0_outputs[4587] = inputs[347];
    assign layer0_outputs[4588] = ~(inputs[834]) | (inputs[929]);
    assign layer0_outputs[4589] = inputs[548];
    assign layer0_outputs[4590] = ~(inputs[427]);
    assign layer0_outputs[4591] = (inputs[617]) ^ (inputs[92]);
    assign layer0_outputs[4592] = inputs[584];
    assign layer0_outputs[4593] = ~((inputs[169]) | (inputs[784]));
    assign layer0_outputs[4594] = (inputs[878]) | (inputs[304]);
    assign layer0_outputs[4595] = (inputs[423]) & ~(inputs[449]);
    assign layer0_outputs[4596] = (inputs[90]) ^ (inputs[94]);
    assign layer0_outputs[4597] = ~(inputs[678]);
    assign layer0_outputs[4598] = (inputs[496]) & (inputs[249]);
    assign layer0_outputs[4599] = ~((inputs[168]) & (inputs[37]));
    assign layer0_outputs[4600] = ~(inputs[266]);
    assign layer0_outputs[4601] = (inputs[355]) ^ (inputs[506]);
    assign layer0_outputs[4602] = ~(inputs[237]);
    assign layer0_outputs[4603] = (inputs[175]) ^ (inputs[81]);
    assign layer0_outputs[4604] = inputs[211];
    assign layer0_outputs[4605] = (inputs[240]) ^ (inputs[776]);
    assign layer0_outputs[4606] = inputs[494];
    assign layer0_outputs[4607] = (inputs[136]) | (inputs[498]);
    assign layer0_outputs[4608] = (inputs[779]) | (inputs[502]);
    assign layer0_outputs[4609] = ~(inputs[398]);
    assign layer0_outputs[4610] = ~(inputs[866]) | (inputs[477]);
    assign layer0_outputs[4611] = ~(inputs[439]) | (inputs[771]);
    assign layer0_outputs[4612] = (inputs[843]) | (inputs[231]);
    assign layer0_outputs[4613] = ~((inputs[564]) & (inputs[270]));
    assign layer0_outputs[4614] = (inputs[490]) ^ (inputs[396]);
    assign layer0_outputs[4615] = ~((inputs[358]) ^ (inputs[707]));
    assign layer0_outputs[4616] = (inputs[811]) ^ (inputs[443]);
    assign layer0_outputs[4617] = (inputs[820]) & ~(inputs[192]);
    assign layer0_outputs[4618] = (inputs[624]) & ~(inputs[50]);
    assign layer0_outputs[4619] = ~(inputs[878]) | (inputs[539]);
    assign layer0_outputs[4620] = inputs[335];
    assign layer0_outputs[4621] = inputs[861];
    assign layer0_outputs[4622] = ~(inputs[930]) | (inputs[123]);
    assign layer0_outputs[4623] = (inputs[483]) & ~(inputs[925]);
    assign layer0_outputs[4624] = ~(inputs[674]) | (inputs[731]);
    assign layer0_outputs[4625] = ~((inputs[708]) | (inputs[306]));
    assign layer0_outputs[4626] = inputs[427];
    assign layer0_outputs[4627] = (inputs[193]) & (inputs[641]);
    assign layer0_outputs[4628] = ~(inputs[106]) | (inputs[670]);
    assign layer0_outputs[4629] = ~(inputs[852]);
    assign layer0_outputs[4630] = ~((inputs[560]) ^ (inputs[227]));
    assign layer0_outputs[4631] = ~(inputs[976]);
    assign layer0_outputs[4632] = ~(inputs[45]);
    assign layer0_outputs[4633] = ~((inputs[122]) | (inputs[495]));
    assign layer0_outputs[4634] = ~((inputs[911]) | (inputs[152]));
    assign layer0_outputs[4635] = (inputs[228]) & (inputs[735]);
    assign layer0_outputs[4636] = ~(inputs[658]) | (inputs[839]);
    assign layer0_outputs[4637] = inputs[304];
    assign layer0_outputs[4638] = inputs[270];
    assign layer0_outputs[4639] = (inputs[801]) | (inputs[458]);
    assign layer0_outputs[4640] = ~(inputs[901]);
    assign layer0_outputs[4641] = ~((inputs[931]) | (inputs[654]));
    assign layer0_outputs[4642] = ~((inputs[906]) | (inputs[431]));
    assign layer0_outputs[4643] = inputs[737];
    assign layer0_outputs[4644] = (inputs[192]) ^ (inputs[555]);
    assign layer0_outputs[4645] = ~(inputs[406]) | (inputs[861]);
    assign layer0_outputs[4646] = (inputs[586]) & ~(inputs[600]);
    assign layer0_outputs[4647] = (inputs[931]) & (inputs[162]);
    assign layer0_outputs[4648] = (inputs[788]) & ~(inputs[671]);
    assign layer0_outputs[4649] = ~((inputs[841]) | (inputs[95]));
    assign layer0_outputs[4650] = (inputs[790]) & ~(inputs[1018]);
    assign layer0_outputs[4651] = ~(inputs[696]) | (inputs[833]);
    assign layer0_outputs[4652] = ~((inputs[876]) & (inputs[752]));
    assign layer0_outputs[4653] = ~((inputs[687]) ^ (inputs[767]));
    assign layer0_outputs[4654] = (inputs[411]) | (inputs[227]);
    assign layer0_outputs[4655] = ~(inputs[559]) | (inputs[76]);
    assign layer0_outputs[4656] = (inputs[332]) | (inputs[487]);
    assign layer0_outputs[4657] = (inputs[207]) & ~(inputs[835]);
    assign layer0_outputs[4658] = (inputs[147]) & ~(inputs[764]);
    assign layer0_outputs[4659] = 1'b0;
    assign layer0_outputs[4660] = inputs[444];
    assign layer0_outputs[4661] = (inputs[176]) | (inputs[770]);
    assign layer0_outputs[4662] = ~(inputs[459]) | (inputs[807]);
    assign layer0_outputs[4663] = ~(inputs[625]) | (inputs[538]);
    assign layer0_outputs[4664] = ~((inputs[758]) ^ (inputs[552]));
    assign layer0_outputs[4665] = ~((inputs[19]) ^ (inputs[93]));
    assign layer0_outputs[4666] = (inputs[272]) | (inputs[649]);
    assign layer0_outputs[4667] = ~((inputs[820]) | (inputs[374]));
    assign layer0_outputs[4668] = ~(inputs[316]) | (inputs[326]);
    assign layer0_outputs[4669] = (inputs[123]) ^ (inputs[807]);
    assign layer0_outputs[4670] = (inputs[728]) | (inputs[765]);
    assign layer0_outputs[4671] = ~((inputs[458]) | (inputs[926]));
    assign layer0_outputs[4672] = (inputs[586]) & ~(inputs[912]);
    assign layer0_outputs[4673] = ~(inputs[768]);
    assign layer0_outputs[4674] = (inputs[310]) | (inputs[193]);
    assign layer0_outputs[4675] = ~((inputs[392]) | (inputs[499]));
    assign layer0_outputs[4676] = ~(inputs[487]) | (inputs[858]);
    assign layer0_outputs[4677] = (inputs[881]) & (inputs[570]);
    assign layer0_outputs[4678] = ~(inputs[95]) | (inputs[292]);
    assign layer0_outputs[4679] = inputs[472];
    assign layer0_outputs[4680] = (inputs[850]) | (inputs[598]);
    assign layer0_outputs[4681] = ~((inputs[676]) | (inputs[8]));
    assign layer0_outputs[4682] = ~(inputs[1008]);
    assign layer0_outputs[4683] = (inputs[239]) ^ (inputs[176]);
    assign layer0_outputs[4684] = ~((inputs[611]) ^ (inputs[6]));
    assign layer0_outputs[4685] = ~(inputs[407]);
    assign layer0_outputs[4686] = (inputs[344]) & ~(inputs[804]);
    assign layer0_outputs[4687] = (inputs[1008]) ^ (inputs[187]);
    assign layer0_outputs[4688] = inputs[902];
    assign layer0_outputs[4689] = ~(inputs[427]);
    assign layer0_outputs[4690] = (inputs[220]) & ~(inputs[236]);
    assign layer0_outputs[4691] = ~((inputs[756]) | (inputs[113]));
    assign layer0_outputs[4692] = ~(inputs[814]) | (inputs[109]);
    assign layer0_outputs[4693] = ~((inputs[265]) | (inputs[817]));
    assign layer0_outputs[4694] = (inputs[808]) | (inputs[483]);
    assign layer0_outputs[4695] = ~(inputs[302]) | (inputs[868]);
    assign layer0_outputs[4696] = ~((inputs[701]) | (inputs[274]));
    assign layer0_outputs[4697] = inputs[771];
    assign layer0_outputs[4698] = ~((inputs[351]) ^ (inputs[595]));
    assign layer0_outputs[4699] = ~(inputs[899]);
    assign layer0_outputs[4700] = (inputs[468]) | (inputs[901]);
    assign layer0_outputs[4701] = ~(inputs[1010]) | (inputs[727]);
    assign layer0_outputs[4702] = (inputs[96]) & (inputs[964]);
    assign layer0_outputs[4703] = inputs[245];
    assign layer0_outputs[4704] = (inputs[723]) | (inputs[252]);
    assign layer0_outputs[4705] = ~(inputs[836]);
    assign layer0_outputs[4706] = inputs[144];
    assign layer0_outputs[4707] = (inputs[133]) & (inputs[537]);
    assign layer0_outputs[4708] = (inputs[930]) ^ (inputs[986]);
    assign layer0_outputs[4709] = ~(inputs[308]) | (inputs[325]);
    assign layer0_outputs[4710] = ~(inputs[435]);
    assign layer0_outputs[4711] = (inputs[222]) & ~(inputs[514]);
    assign layer0_outputs[4712] = ~((inputs[846]) | (inputs[697]));
    assign layer0_outputs[4713] = ~(inputs[817]);
    assign layer0_outputs[4714] = (inputs[801]) & (inputs[506]);
    assign layer0_outputs[4715] = 1'b1;
    assign layer0_outputs[4716] = ~(inputs[154]) | (inputs[512]);
    assign layer0_outputs[4717] = 1'b0;
    assign layer0_outputs[4718] = (inputs[271]) & ~(inputs[603]);
    assign layer0_outputs[4719] = ~((inputs[54]) | (inputs[306]));
    assign layer0_outputs[4720] = 1'b1;
    assign layer0_outputs[4721] = ~(inputs[360]) | (inputs[920]);
    assign layer0_outputs[4722] = (inputs[142]) | (inputs[481]);
    assign layer0_outputs[4723] = (inputs[655]) | (inputs[456]);
    assign layer0_outputs[4724] = ~((inputs[799]) ^ (inputs[777]));
    assign layer0_outputs[4725] = ~((inputs[199]) | (inputs[370]));
    assign layer0_outputs[4726] = ~(inputs[507]) | (inputs[165]);
    assign layer0_outputs[4727] = ~((inputs[458]) ^ (inputs[417]));
    assign layer0_outputs[4728] = ~((inputs[444]) ^ (inputs[734]));
    assign layer0_outputs[4729] = (inputs[19]) & ~(inputs[574]);
    assign layer0_outputs[4730] = inputs[39];
    assign layer0_outputs[4731] = (inputs[988]) ^ (inputs[899]);
    assign layer0_outputs[4732] = inputs[993];
    assign layer0_outputs[4733] = ~(inputs[972]) | (inputs[143]);
    assign layer0_outputs[4734] = (inputs[556]) ^ (inputs[84]);
    assign layer0_outputs[4735] = (inputs[183]) | (inputs[875]);
    assign layer0_outputs[4736] = (inputs[716]) | (inputs[857]);
    assign layer0_outputs[4737] = (inputs[233]) | (inputs[757]);
    assign layer0_outputs[4738] = ~(inputs[560]);
    assign layer0_outputs[4739] = 1'b0;
    assign layer0_outputs[4740] = ~((inputs[420]) & (inputs[927]));
    assign layer0_outputs[4741] = (inputs[668]) | (inputs[717]);
    assign layer0_outputs[4742] = (inputs[368]) & ~(inputs[18]);
    assign layer0_outputs[4743] = inputs[38];
    assign layer0_outputs[4744] = ~((inputs[527]) ^ (inputs[53]));
    assign layer0_outputs[4745] = ~((inputs[776]) ^ (inputs[69]));
    assign layer0_outputs[4746] = inputs[301];
    assign layer0_outputs[4747] = inputs[148];
    assign layer0_outputs[4748] = ~(inputs[521]) | (inputs[293]);
    assign layer0_outputs[4749] = (inputs[773]) & (inputs[861]);
    assign layer0_outputs[4750] = (inputs[867]) | (inputs[8]);
    assign layer0_outputs[4751] = (inputs[345]) | (inputs[629]);
    assign layer0_outputs[4752] = ~((inputs[646]) ^ (inputs[573]));
    assign layer0_outputs[4753] = (inputs[409]) | (inputs[261]);
    assign layer0_outputs[4754] = 1'b1;
    assign layer0_outputs[4755] = ~(inputs[819]);
    assign layer0_outputs[4756] = (inputs[337]) & ~(inputs[450]);
    assign layer0_outputs[4757] = (inputs[92]) | (inputs[659]);
    assign layer0_outputs[4758] = ~((inputs[846]) | (inputs[1003]));
    assign layer0_outputs[4759] = ~(inputs[908]);
    assign layer0_outputs[4760] = ~((inputs[653]) ^ (inputs[479]));
    assign layer0_outputs[4761] = ~(inputs[113]) | (inputs[102]);
    assign layer0_outputs[4762] = (inputs[306]) & ~(inputs[696]);
    assign layer0_outputs[4763] = (inputs[473]) ^ (inputs[240]);
    assign layer0_outputs[4764] = (inputs[180]) & ~(inputs[423]);
    assign layer0_outputs[4765] = (inputs[424]) | (inputs[362]);
    assign layer0_outputs[4766] = ~((inputs[915]) | (inputs[266]));
    assign layer0_outputs[4767] = ~(inputs[440]);
    assign layer0_outputs[4768] = ~((inputs[864]) ^ (inputs[133]));
    assign layer0_outputs[4769] = 1'b0;
    assign layer0_outputs[4770] = (inputs[775]) ^ (inputs[6]);
    assign layer0_outputs[4771] = (inputs[215]) | (inputs[634]);
    assign layer0_outputs[4772] = (inputs[366]) & ~(inputs[105]);
    assign layer0_outputs[4773] = inputs[979];
    assign layer0_outputs[4774] = ~(inputs[940]);
    assign layer0_outputs[4775] = 1'b1;
    assign layer0_outputs[4776] = ~(inputs[529]) | (inputs[12]);
    assign layer0_outputs[4777] = ~(inputs[41]);
    assign layer0_outputs[4778] = (inputs[479]) | (inputs[582]);
    assign layer0_outputs[4779] = (inputs[322]) & ~(inputs[321]);
    assign layer0_outputs[4780] = (inputs[753]) & ~(inputs[749]);
    assign layer0_outputs[4781] = (inputs[345]) | (inputs[276]);
    assign layer0_outputs[4782] = ~((inputs[146]) ^ (inputs[103]));
    assign layer0_outputs[4783] = ~(inputs[906]);
    assign layer0_outputs[4784] = (inputs[877]) & ~(inputs[987]);
    assign layer0_outputs[4785] = inputs[814];
    assign layer0_outputs[4786] = (inputs[922]) & (inputs[956]);
    assign layer0_outputs[4787] = (inputs[698]) ^ (inputs[762]);
    assign layer0_outputs[4788] = ~((inputs[530]) | (inputs[316]));
    assign layer0_outputs[4789] = ~(inputs[840]) | (inputs[504]);
    assign layer0_outputs[4790] = (inputs[851]) ^ (inputs[923]);
    assign layer0_outputs[4791] = (inputs[604]) | (inputs[264]);
    assign layer0_outputs[4792] = (inputs[890]) & (inputs[870]);
    assign layer0_outputs[4793] = ~(inputs[630]);
    assign layer0_outputs[4794] = inputs[743];
    assign layer0_outputs[4795] = (inputs[314]) ^ (inputs[512]);
    assign layer0_outputs[4796] = (inputs[515]) & (inputs[797]);
    assign layer0_outputs[4797] = ~((inputs[375]) ^ (inputs[379]));
    assign layer0_outputs[4798] = (inputs[331]) ^ (inputs[937]);
    assign layer0_outputs[4799] = (inputs[595]) & ~(inputs[756]);
    assign layer0_outputs[4800] = ~(inputs[631]) | (inputs[393]);
    assign layer0_outputs[4801] = ~((inputs[56]) ^ (inputs[735]));
    assign layer0_outputs[4802] = (inputs[535]) | (inputs[250]);
    assign layer0_outputs[4803] = ~((inputs[973]) ^ (inputs[114]));
    assign layer0_outputs[4804] = ~(inputs[469]);
    assign layer0_outputs[4805] = ~((inputs[142]) | (inputs[539]));
    assign layer0_outputs[4806] = inputs[706];
    assign layer0_outputs[4807] = (inputs[805]) ^ (inputs[705]);
    assign layer0_outputs[4808] = ~(inputs[345]) | (inputs[355]);
    assign layer0_outputs[4809] = inputs[277];
    assign layer0_outputs[4810] = (inputs[974]) | (inputs[599]);
    assign layer0_outputs[4811] = (inputs[659]) & (inputs[275]);
    assign layer0_outputs[4812] = ~((inputs[159]) | (inputs[10]));
    assign layer0_outputs[4813] = ~(inputs[434]) | (inputs[4]);
    assign layer0_outputs[4814] = (inputs[499]) & ~(inputs[283]);
    assign layer0_outputs[4815] = ~(inputs[361]);
    assign layer0_outputs[4816] = ~(inputs[1007]) | (inputs[983]);
    assign layer0_outputs[4817] = inputs[139];
    assign layer0_outputs[4818] = (inputs[105]) & (inputs[926]);
    assign layer0_outputs[4819] = (inputs[429]) & ~(inputs[89]);
    assign layer0_outputs[4820] = ~((inputs[445]) ^ (inputs[429]));
    assign layer0_outputs[4821] = ~(inputs[719]);
    assign layer0_outputs[4822] = (inputs[334]) | (inputs[1012]);
    assign layer0_outputs[4823] = inputs[736];
    assign layer0_outputs[4824] = (inputs[353]) ^ (inputs[492]);
    assign layer0_outputs[4825] = ~((inputs[903]) ^ (inputs[892]));
    assign layer0_outputs[4826] = ~((inputs[199]) ^ (inputs[703]));
    assign layer0_outputs[4827] = ~(inputs[430]);
    assign layer0_outputs[4828] = (inputs[450]) & ~(inputs[890]);
    assign layer0_outputs[4829] = 1'b1;
    assign layer0_outputs[4830] = ~(inputs[941]);
    assign layer0_outputs[4831] = (inputs[989]) ^ (inputs[349]);
    assign layer0_outputs[4832] = (inputs[105]) & ~(inputs[67]);
    assign layer0_outputs[4833] = (inputs[906]) | (inputs[203]);
    assign layer0_outputs[4834] = (inputs[165]) & (inputs[116]);
    assign layer0_outputs[4835] = ~(inputs[476]);
    assign layer0_outputs[4836] = ~(inputs[12]) | (inputs[923]);
    assign layer0_outputs[4837] = ~((inputs[771]) | (inputs[376]));
    assign layer0_outputs[4838] = (inputs[650]) | (inputs[486]);
    assign layer0_outputs[4839] = inputs[585];
    assign layer0_outputs[4840] = ~(inputs[4]);
    assign layer0_outputs[4841] = (inputs[386]) ^ (inputs[375]);
    assign layer0_outputs[4842] = ~(inputs[855]);
    assign layer0_outputs[4843] = ~(inputs[221]);
    assign layer0_outputs[4844] = ~(inputs[847]);
    assign layer0_outputs[4845] = 1'b1;
    assign layer0_outputs[4846] = ~(inputs[938]);
    assign layer0_outputs[4847] = 1'b1;
    assign layer0_outputs[4848] = ~(inputs[729]);
    assign layer0_outputs[4849] = 1'b0;
    assign layer0_outputs[4850] = ~((inputs[151]) | (inputs[752]));
    assign layer0_outputs[4851] = ~(inputs[898]);
    assign layer0_outputs[4852] = ~((inputs[730]) ^ (inputs[304]));
    assign layer0_outputs[4853] = ~((inputs[100]) | (inputs[738]));
    assign layer0_outputs[4854] = (inputs[883]) & (inputs[10]);
    assign layer0_outputs[4855] = ~(inputs[980]);
    assign layer0_outputs[4856] = inputs[532];
    assign layer0_outputs[4857] = ~((inputs[364]) | (inputs[629]));
    assign layer0_outputs[4858] = ~(inputs[409]) | (inputs[259]);
    assign layer0_outputs[4859] = 1'b1;
    assign layer0_outputs[4860] = inputs[911];
    assign layer0_outputs[4861] = (inputs[635]) | (inputs[777]);
    assign layer0_outputs[4862] = inputs[564];
    assign layer0_outputs[4863] = inputs[717];
    assign layer0_outputs[4864] = (inputs[521]) & ~(inputs[872]);
    assign layer0_outputs[4865] = inputs[138];
    assign layer0_outputs[4866] = ~(inputs[500]);
    assign layer0_outputs[4867] = ~(inputs[473]) | (inputs[630]);
    assign layer0_outputs[4868] = ~((inputs[730]) | (inputs[109]));
    assign layer0_outputs[4869] = ~((inputs[377]) ^ (inputs[803]));
    assign layer0_outputs[4870] = (inputs[535]) ^ (inputs[813]);
    assign layer0_outputs[4871] = (inputs[20]) & ~(inputs[99]);
    assign layer0_outputs[4872] = ~(inputs[231]);
    assign layer0_outputs[4873] = ~((inputs[793]) | (inputs[646]));
    assign layer0_outputs[4874] = inputs[667];
    assign layer0_outputs[4875] = ~(inputs[488]);
    assign layer0_outputs[4876] = ~(inputs[818]);
    assign layer0_outputs[4877] = (inputs[479]) | (inputs[958]);
    assign layer0_outputs[4878] = (inputs[86]) | (inputs[146]);
    assign layer0_outputs[4879] = ~(inputs[355]) | (inputs[157]);
    assign layer0_outputs[4880] = (inputs[745]) ^ (inputs[800]);
    assign layer0_outputs[4881] = ~((inputs[397]) | (inputs[891]));
    assign layer0_outputs[4882] = (inputs[375]) | (inputs[874]);
    assign layer0_outputs[4883] = ~(inputs[411]) | (inputs[478]);
    assign layer0_outputs[4884] = inputs[467];
    assign layer0_outputs[4885] = (inputs[900]) | (inputs[716]);
    assign layer0_outputs[4886] = ~(inputs[549]);
    assign layer0_outputs[4887] = ~(inputs[98]);
    assign layer0_outputs[4888] = ~(inputs[492]);
    assign layer0_outputs[4889] = (inputs[1005]) & ~(inputs[666]);
    assign layer0_outputs[4890] = ~(inputs[888]) | (inputs[378]);
    assign layer0_outputs[4891] = ~(inputs[689]);
    assign layer0_outputs[4892] = ~(inputs[651]);
    assign layer0_outputs[4893] = ~((inputs[959]) ^ (inputs[780]));
    assign layer0_outputs[4894] = (inputs[514]) | (inputs[500]);
    assign layer0_outputs[4895] = inputs[248];
    assign layer0_outputs[4896] = 1'b1;
    assign layer0_outputs[4897] = ~(inputs[382]);
    assign layer0_outputs[4898] = (inputs[137]) & ~(inputs[925]);
    assign layer0_outputs[4899] = (inputs[751]) ^ (inputs[225]);
    assign layer0_outputs[4900] = ~(inputs[805]) | (inputs[455]);
    assign layer0_outputs[4901] = inputs[883];
    assign layer0_outputs[4902] = ~((inputs[779]) | (inputs[349]));
    assign layer0_outputs[4903] = inputs[495];
    assign layer0_outputs[4904] = ~((inputs[1015]) ^ (inputs[74]));
    assign layer0_outputs[4905] = (inputs[207]) | (inputs[722]);
    assign layer0_outputs[4906] = (inputs[671]) ^ (inputs[571]);
    assign layer0_outputs[4907] = inputs[844];
    assign layer0_outputs[4908] = ~(inputs[28]);
    assign layer0_outputs[4909] = 1'b0;
    assign layer0_outputs[4910] = inputs[838];
    assign layer0_outputs[4911] = ~(inputs[533]) | (inputs[27]);
    assign layer0_outputs[4912] = inputs[495];
    assign layer0_outputs[4913] = ~((inputs[965]) ^ (inputs[122]));
    assign layer0_outputs[4914] = ~((inputs[819]) ^ (inputs[754]));
    assign layer0_outputs[4915] = inputs[514];
    assign layer0_outputs[4916] = (inputs[865]) ^ (inputs[834]);
    assign layer0_outputs[4917] = ~(inputs[816]) | (inputs[70]);
    assign layer0_outputs[4918] = ~(inputs[818]) | (inputs[260]);
    assign layer0_outputs[4919] = ~(inputs[524]) | (inputs[402]);
    assign layer0_outputs[4920] = 1'b0;
    assign layer0_outputs[4921] = ~(inputs[435]);
    assign layer0_outputs[4922] = ~(inputs[949]) | (inputs[996]);
    assign layer0_outputs[4923] = inputs[953];
    assign layer0_outputs[4924] = 1'b1;
    assign layer0_outputs[4925] = (inputs[815]) & ~(inputs[568]);
    assign layer0_outputs[4926] = ~((inputs[372]) ^ (inputs[864]));
    assign layer0_outputs[4927] = ~(inputs[963]);
    assign layer0_outputs[4928] = (inputs[437]) ^ (inputs[37]);
    assign layer0_outputs[4929] = inputs[596];
    assign layer0_outputs[4930] = ~((inputs[440]) ^ (inputs[863]));
    assign layer0_outputs[4931] = 1'b0;
    assign layer0_outputs[4932] = (inputs[154]) | (inputs[742]);
    assign layer0_outputs[4933] = ~(inputs[179]) | (inputs[792]);
    assign layer0_outputs[4934] = ~((inputs[958]) | (inputs[431]));
    assign layer0_outputs[4935] = ~(inputs[10]) | (inputs[988]);
    assign layer0_outputs[4936] = (inputs[345]) | (inputs[907]);
    assign layer0_outputs[4937] = ~(inputs[371]) | (inputs[948]);
    assign layer0_outputs[4938] = ~((inputs[643]) | (inputs[969]));
    assign layer0_outputs[4939] = ~((inputs[966]) ^ (inputs[885]));
    assign layer0_outputs[4940] = 1'b1;
    assign layer0_outputs[4941] = ~((inputs[95]) | (inputs[389]));
    assign layer0_outputs[4942] = (inputs[158]) | (inputs[378]);
    assign layer0_outputs[4943] = inputs[780];
    assign layer0_outputs[4944] = ~(inputs[949]) | (inputs[80]);
    assign layer0_outputs[4945] = (inputs[726]) & ~(inputs[616]);
    assign layer0_outputs[4946] = inputs[687];
    assign layer0_outputs[4947] = (inputs[783]) ^ (inputs[625]);
    assign layer0_outputs[4948] = (inputs[138]) ^ (inputs[461]);
    assign layer0_outputs[4949] = (inputs[495]) | (inputs[726]);
    assign layer0_outputs[4950] = ~(inputs[676]);
    assign layer0_outputs[4951] = ~((inputs[111]) | (inputs[202]));
    assign layer0_outputs[4952] = ~((inputs[610]) | (inputs[726]));
    assign layer0_outputs[4953] = (inputs[531]) ^ (inputs[597]);
    assign layer0_outputs[4954] = ~((inputs[868]) ^ (inputs[15]));
    assign layer0_outputs[4955] = ~((inputs[601]) ^ (inputs[659]));
    assign layer0_outputs[4956] = inputs[453];
    assign layer0_outputs[4957] = ~(inputs[966]) | (inputs[796]);
    assign layer0_outputs[4958] = ~((inputs[68]) & (inputs[924]));
    assign layer0_outputs[4959] = (inputs[679]) ^ (inputs[542]);
    assign layer0_outputs[4960] = (inputs[75]) & (inputs[544]);
    assign layer0_outputs[4961] = (inputs[766]) | (inputs[239]);
    assign layer0_outputs[4962] = ~(inputs[531]) | (inputs[279]);
    assign layer0_outputs[4963] = inputs[431];
    assign layer0_outputs[4964] = (inputs[297]) ^ (inputs[876]);
    assign layer0_outputs[4965] = ~(inputs[537]) | (inputs[266]);
    assign layer0_outputs[4966] = ~(inputs[951]) | (inputs[766]);
    assign layer0_outputs[4967] = ~((inputs[196]) | (inputs[262]));
    assign layer0_outputs[4968] = inputs[909];
    assign layer0_outputs[4969] = 1'b1;
    assign layer0_outputs[4970] = ~((inputs[985]) | (inputs[357]));
    assign layer0_outputs[4971] = ~((inputs[723]) | (inputs[212]));
    assign layer0_outputs[4972] = ~(inputs[119]) | (inputs[643]);
    assign layer0_outputs[4973] = (inputs[841]) & ~(inputs[221]);
    assign layer0_outputs[4974] = (inputs[402]) | (inputs[937]);
    assign layer0_outputs[4975] = (inputs[853]) | (inputs[870]);
    assign layer0_outputs[4976] = ~(inputs[534]);
    assign layer0_outputs[4977] = ~(inputs[721]) | (inputs[21]);
    assign layer0_outputs[4978] = inputs[204];
    assign layer0_outputs[4979] = inputs[495];
    assign layer0_outputs[4980] = ~(inputs[540]) | (inputs[55]);
    assign layer0_outputs[4981] = ~(inputs[220]);
    assign layer0_outputs[4982] = (inputs[190]) ^ (inputs[930]);
    assign layer0_outputs[4983] = ~(inputs[374]) | (inputs[580]);
    assign layer0_outputs[4984] = ~(inputs[292]);
    assign layer0_outputs[4985] = ~(inputs[83]) | (inputs[910]);
    assign layer0_outputs[4986] = ~((inputs[998]) | (inputs[601]));
    assign layer0_outputs[4987] = ~((inputs[554]) ^ (inputs[259]));
    assign layer0_outputs[4988] = inputs[549];
    assign layer0_outputs[4989] = (inputs[973]) | (inputs[310]);
    assign layer0_outputs[4990] = inputs[860];
    assign layer0_outputs[4991] = ~(inputs[794]);
    assign layer0_outputs[4992] = (inputs[150]) | (inputs[170]);
    assign layer0_outputs[4993] = 1'b0;
    assign layer0_outputs[4994] = (inputs[884]) & ~(inputs[710]);
    assign layer0_outputs[4995] = ~(inputs[757]);
    assign layer0_outputs[4996] = (inputs[732]) | (inputs[815]);
    assign layer0_outputs[4997] = inputs[612];
    assign layer0_outputs[4998] = (inputs[585]) & ~(inputs[967]);
    assign layer0_outputs[4999] = 1'b1;
    assign layer0_outputs[5000] = (inputs[64]) & (inputs[580]);
    assign layer0_outputs[5001] = (inputs[665]) & ~(inputs[995]);
    assign layer0_outputs[5002] = ~(inputs[587]);
    assign layer0_outputs[5003] = (inputs[585]) & ~(inputs[330]);
    assign layer0_outputs[5004] = (inputs[816]) | (inputs[325]);
    assign layer0_outputs[5005] = (inputs[499]) ^ (inputs[7]);
    assign layer0_outputs[5006] = (inputs[694]) & ~(inputs[1]);
    assign layer0_outputs[5007] = ~((inputs[551]) ^ (inputs[1020]));
    assign layer0_outputs[5008] = ~((inputs[183]) | (inputs[49]));
    assign layer0_outputs[5009] = inputs[877];
    assign layer0_outputs[5010] = (inputs[983]) & (inputs[953]);
    assign layer0_outputs[5011] = (inputs[57]) & ~(inputs[75]);
    assign layer0_outputs[5012] = (inputs[325]) | (inputs[795]);
    assign layer0_outputs[5013] = ~((inputs[182]) ^ (inputs[1005]));
    assign layer0_outputs[5014] = (inputs[780]) | (inputs[79]);
    assign layer0_outputs[5015] = ~(inputs[921]);
    assign layer0_outputs[5016] = ~(inputs[784]) | (inputs[844]);
    assign layer0_outputs[5017] = 1'b1;
    assign layer0_outputs[5018] = (inputs[328]) ^ (inputs[316]);
    assign layer0_outputs[5019] = ~(inputs[420]);
    assign layer0_outputs[5020] = ~(inputs[856]);
    assign layer0_outputs[5021] = ~(inputs[20]) | (inputs[768]);
    assign layer0_outputs[5022] = 1'b1;
    assign layer0_outputs[5023] = (inputs[243]) & ~(inputs[285]);
    assign layer0_outputs[5024] = ~(inputs[844]);
    assign layer0_outputs[5025] = ~(inputs[810]) | (inputs[572]);
    assign layer0_outputs[5026] = 1'b0;
    assign layer0_outputs[5027] = 1'b1;
    assign layer0_outputs[5028] = ~(inputs[436]);
    assign layer0_outputs[5029] = ~((inputs[697]) | (inputs[183]));
    assign layer0_outputs[5030] = (inputs[236]) & (inputs[512]);
    assign layer0_outputs[5031] = (inputs[474]) ^ (inputs[336]);
    assign layer0_outputs[5032] = (inputs[543]) | (inputs[812]);
    assign layer0_outputs[5033] = (inputs[21]) ^ (inputs[178]);
    assign layer0_outputs[5034] = (inputs[379]) | (inputs[691]);
    assign layer0_outputs[5035] = (inputs[94]) | (inputs[321]);
    assign layer0_outputs[5036] = ~(inputs[604]) | (inputs[995]);
    assign layer0_outputs[5037] = ~(inputs[624]);
    assign layer0_outputs[5038] = (inputs[825]) & ~(inputs[867]);
    assign layer0_outputs[5039] = inputs[682];
    assign layer0_outputs[5040] = (inputs[824]) | (inputs[399]);
    assign layer0_outputs[5041] = inputs[374];
    assign layer0_outputs[5042] = ~((inputs[341]) | (inputs[933]));
    assign layer0_outputs[5043] = ~((inputs[739]) ^ (inputs[811]));
    assign layer0_outputs[5044] = inputs[293];
    assign layer0_outputs[5045] = inputs[274];
    assign layer0_outputs[5046] = (inputs[717]) & ~(inputs[280]);
    assign layer0_outputs[5047] = (inputs[161]) & ~(inputs[966]);
    assign layer0_outputs[5048] = ~(inputs[651]) | (inputs[704]);
    assign layer0_outputs[5049] = (inputs[529]) & ~(inputs[233]);
    assign layer0_outputs[5050] = ~(inputs[881]);
    assign layer0_outputs[5051] = ~((inputs[842]) | (inputs[934]));
    assign layer0_outputs[5052] = ~(inputs[267]);
    assign layer0_outputs[5053] = ~(inputs[329]);
    assign layer0_outputs[5054] = ~(inputs[25]);
    assign layer0_outputs[5055] = ~((inputs[857]) & (inputs[190]));
    assign layer0_outputs[5056] = (inputs[160]) ^ (inputs[645]);
    assign layer0_outputs[5057] = ~((inputs[812]) | (inputs[796]));
    assign layer0_outputs[5058] = (inputs[536]) | (inputs[79]);
    assign layer0_outputs[5059] = (inputs[128]) ^ (inputs[344]);
    assign layer0_outputs[5060] = ~(inputs[338]) | (inputs[476]);
    assign layer0_outputs[5061] = ~(inputs[116]);
    assign layer0_outputs[5062] = (inputs[998]) & ~(inputs[105]);
    assign layer0_outputs[5063] = ~(inputs[492]);
    assign layer0_outputs[5064] = (inputs[41]) & (inputs[582]);
    assign layer0_outputs[5065] = 1'b1;
    assign layer0_outputs[5066] = ~((inputs[654]) | (inputs[793]));
    assign layer0_outputs[5067] = (inputs[373]) & ~(inputs[511]);
    assign layer0_outputs[5068] = ~(inputs[72]) | (inputs[511]);
    assign layer0_outputs[5069] = inputs[779];
    assign layer0_outputs[5070] = ~((inputs[940]) ^ (inputs[608]));
    assign layer0_outputs[5071] = ~(inputs[834]) | (inputs[219]);
    assign layer0_outputs[5072] = inputs[955];
    assign layer0_outputs[5073] = ~((inputs[787]) ^ (inputs[992]));
    assign layer0_outputs[5074] = ~(inputs[522]);
    assign layer0_outputs[5075] = (inputs[398]) | (inputs[476]);
    assign layer0_outputs[5076] = ~(inputs[473]);
    assign layer0_outputs[5077] = (inputs[204]) | (inputs[687]);
    assign layer0_outputs[5078] = (inputs[88]) ^ (inputs[72]);
    assign layer0_outputs[5079] = ~(inputs[115]);
    assign layer0_outputs[5080] = 1'b0;
    assign layer0_outputs[5081] = inputs[215];
    assign layer0_outputs[5082] = ~(inputs[583]) | (inputs[778]);
    assign layer0_outputs[5083] = ~((inputs[963]) | (inputs[655]));
    assign layer0_outputs[5084] = ~((inputs[65]) | (inputs[697]));
    assign layer0_outputs[5085] = (inputs[686]) & ~(inputs[410]);
    assign layer0_outputs[5086] = ~(inputs[622]);
    assign layer0_outputs[5087] = (inputs[30]) | (inputs[549]);
    assign layer0_outputs[5088] = (inputs[8]) ^ (inputs[420]);
    assign layer0_outputs[5089] = ~((inputs[836]) | (inputs[892]));
    assign layer0_outputs[5090] = ~(inputs[117]);
    assign layer0_outputs[5091] = ~(inputs[688]);
    assign layer0_outputs[5092] = (inputs[542]) & (inputs[866]);
    assign layer0_outputs[5093] = ~(inputs[404]);
    assign layer0_outputs[5094] = (inputs[708]) ^ (inputs[176]);
    assign layer0_outputs[5095] = ~((inputs[637]) | (inputs[176]));
    assign layer0_outputs[5096] = ~((inputs[66]) ^ (inputs[429]));
    assign layer0_outputs[5097] = ~((inputs[79]) | (inputs[691]));
    assign layer0_outputs[5098] = inputs[421];
    assign layer0_outputs[5099] = ~((inputs[806]) | (inputs[46]));
    assign layer0_outputs[5100] = ~(inputs[432]) | (inputs[735]);
    assign layer0_outputs[5101] = ~(inputs[597]) | (inputs[619]);
    assign layer0_outputs[5102] = (inputs[520]) | (inputs[904]);
    assign layer0_outputs[5103] = ~(inputs[498]);
    assign layer0_outputs[5104] = 1'b0;
    assign layer0_outputs[5105] = ~(inputs[107]) | (inputs[967]);
    assign layer0_outputs[5106] = (inputs[974]) | (inputs[157]);
    assign layer0_outputs[5107] = ~((inputs[653]) | (inputs[692]));
    assign layer0_outputs[5108] = ~(inputs[818]) | (inputs[148]);
    assign layer0_outputs[5109] = (inputs[721]) | (inputs[797]);
    assign layer0_outputs[5110] = ~((inputs[648]) ^ (inputs[478]));
    assign layer0_outputs[5111] = ~((inputs[51]) | (inputs[177]));
    assign layer0_outputs[5112] = ~(inputs[813]);
    assign layer0_outputs[5113] = inputs[416];
    assign layer0_outputs[5114] = ~((inputs[697]) | (inputs[795]));
    assign layer0_outputs[5115] = ~(inputs[849]);
    assign layer0_outputs[5116] = 1'b1;
    assign layer0_outputs[5117] = ~((inputs[60]) & (inputs[829]));
    assign layer0_outputs[5118] = (inputs[139]) | (inputs[845]);
    assign layer0_outputs[5119] = ~(inputs[200]) | (inputs[147]);
    assign layer0_outputs[5120] = 1'b0;
    assign layer0_outputs[5121] = (inputs[779]) & ~(inputs[254]);
    assign layer0_outputs[5122] = ~(inputs[363]) | (inputs[205]);
    assign layer0_outputs[5123] = ~((inputs[369]) ^ (inputs[269]));
    assign layer0_outputs[5124] = inputs[213];
    assign layer0_outputs[5125] = ~((inputs[640]) ^ (inputs[20]));
    assign layer0_outputs[5126] = (inputs[881]) & ~(inputs[987]);
    assign layer0_outputs[5127] = ~(inputs[900]) | (inputs[909]);
    assign layer0_outputs[5128] = (inputs[59]) | (inputs[874]);
    assign layer0_outputs[5129] = ~((inputs[540]) ^ (inputs[782]));
    assign layer0_outputs[5130] = ~((inputs[389]) ^ (inputs[633]));
    assign layer0_outputs[5131] = (inputs[936]) | (inputs[503]);
    assign layer0_outputs[5132] = (inputs[554]) & ~(inputs[420]);
    assign layer0_outputs[5133] = (inputs[407]) ^ (inputs[201]);
    assign layer0_outputs[5134] = inputs[783];
    assign layer0_outputs[5135] = inputs[879];
    assign layer0_outputs[5136] = inputs[334];
    assign layer0_outputs[5137] = inputs[737];
    assign layer0_outputs[5138] = (inputs[585]) ^ (inputs[448]);
    assign layer0_outputs[5139] = ~(inputs[212]);
    assign layer0_outputs[5140] = 1'b0;
    assign layer0_outputs[5141] = (inputs[62]) & ~(inputs[169]);
    assign layer0_outputs[5142] = ~((inputs[800]) ^ (inputs[965]));
    assign layer0_outputs[5143] = (inputs[577]) & (inputs[953]);
    assign layer0_outputs[5144] = (inputs[823]) & ~(inputs[344]);
    assign layer0_outputs[5145] = ~((inputs[703]) | (inputs[875]));
    assign layer0_outputs[5146] = ~((inputs[367]) ^ (inputs[334]));
    assign layer0_outputs[5147] = 1'b1;
    assign layer0_outputs[5148] = (inputs[305]) | (inputs[287]);
    assign layer0_outputs[5149] = (inputs[792]) ^ (inputs[663]);
    assign layer0_outputs[5150] = ~((inputs[63]) | (inputs[224]));
    assign layer0_outputs[5151] = ~(inputs[313]);
    assign layer0_outputs[5152] = (inputs[311]) | (inputs[30]);
    assign layer0_outputs[5153] = inputs[432];
    assign layer0_outputs[5154] = (inputs[916]) ^ (inputs[199]);
    assign layer0_outputs[5155] = ~((inputs[150]) ^ (inputs[751]));
    assign layer0_outputs[5156] = ~(inputs[436]);
    assign layer0_outputs[5157] = ~((inputs[480]) ^ (inputs[245]));
    assign layer0_outputs[5158] = ~(inputs[122]);
    assign layer0_outputs[5159] = 1'b1;
    assign layer0_outputs[5160] = (inputs[1021]) | (inputs[550]);
    assign layer0_outputs[5161] = ~((inputs[912]) ^ (inputs[559]));
    assign layer0_outputs[5162] = (inputs[553]) & ~(inputs[991]);
    assign layer0_outputs[5163] = ~((inputs[598]) ^ (inputs[821]));
    assign layer0_outputs[5164] = ~((inputs[136]) | (inputs[40]));
    assign layer0_outputs[5165] = (inputs[493]) ^ (inputs[806]);
    assign layer0_outputs[5166] = ~(inputs[844]);
    assign layer0_outputs[5167] = inputs[66];
    assign layer0_outputs[5168] = ~(inputs[594]);
    assign layer0_outputs[5169] = ~(inputs[703]);
    assign layer0_outputs[5170] = ~(inputs[489]) | (inputs[384]);
    assign layer0_outputs[5171] = (inputs[858]) ^ (inputs[30]);
    assign layer0_outputs[5172] = ~(inputs[749]);
    assign layer0_outputs[5173] = ~((inputs[87]) ^ (inputs[692]));
    assign layer0_outputs[5174] = ~(inputs[726]) | (inputs[883]);
    assign layer0_outputs[5175] = (inputs[465]) & ~(inputs[426]);
    assign layer0_outputs[5176] = ~((inputs[474]) | (inputs[428]));
    assign layer0_outputs[5177] = (inputs[200]) & ~(inputs[858]);
    assign layer0_outputs[5178] = (inputs[357]) & (inputs[132]);
    assign layer0_outputs[5179] = inputs[428];
    assign layer0_outputs[5180] = 1'b0;
    assign layer0_outputs[5181] = ~((inputs[258]) ^ (inputs[710]));
    assign layer0_outputs[5182] = (inputs[589]) | (inputs[668]);
    assign layer0_outputs[5183] = ~(inputs[153]);
    assign layer0_outputs[5184] = (inputs[617]) ^ (inputs[997]);
    assign layer0_outputs[5185] = ~((inputs[214]) & (inputs[832]));
    assign layer0_outputs[5186] = (inputs[189]) & ~(inputs[14]);
    assign layer0_outputs[5187] = ~(inputs[534]) | (inputs[87]);
    assign layer0_outputs[5188] = (inputs[35]) ^ (inputs[605]);
    assign layer0_outputs[5189] = inputs[314];
    assign layer0_outputs[5190] = ~((inputs[690]) | (inputs[118]));
    assign layer0_outputs[5191] = (inputs[385]) & ~(inputs[573]);
    assign layer0_outputs[5192] = inputs[307];
    assign layer0_outputs[5193] = ~(inputs[717]) | (inputs[277]);
    assign layer0_outputs[5194] = ~(inputs[472]) | (inputs[201]);
    assign layer0_outputs[5195] = ~(inputs[731]);
    assign layer0_outputs[5196] = inputs[780];
    assign layer0_outputs[5197] = ~(inputs[756]) | (inputs[510]);
    assign layer0_outputs[5198] = 1'b0;
    assign layer0_outputs[5199] = (inputs[927]) | (inputs[724]);
    assign layer0_outputs[5200] = (inputs[380]) | (inputs[143]);
    assign layer0_outputs[5201] = 1'b1;
    assign layer0_outputs[5202] = ~(inputs[395]) | (inputs[355]);
    assign layer0_outputs[5203] = ~(inputs[913]);
    assign layer0_outputs[5204] = ~(inputs[237]);
    assign layer0_outputs[5205] = ~(inputs[454]) | (inputs[796]);
    assign layer0_outputs[5206] = ~((inputs[469]) ^ (inputs[670]));
    assign layer0_outputs[5207] = inputs[653];
    assign layer0_outputs[5208] = (inputs[453]) & ~(inputs[197]);
    assign layer0_outputs[5209] = ~((inputs[844]) | (inputs[213]));
    assign layer0_outputs[5210] = inputs[615];
    assign layer0_outputs[5211] = inputs[571];
    assign layer0_outputs[5212] = inputs[308];
    assign layer0_outputs[5213] = ~(inputs[70]) | (inputs[871]);
    assign layer0_outputs[5214] = ~((inputs[368]) & (inputs[337]));
    assign layer0_outputs[5215] = ~((inputs[520]) | (inputs[879]));
    assign layer0_outputs[5216] = (inputs[437]) & ~(inputs[667]);
    assign layer0_outputs[5217] = ~((inputs[222]) | (inputs[854]));
    assign layer0_outputs[5218] = (inputs[273]) ^ (inputs[131]);
    assign layer0_outputs[5219] = (inputs[376]) ^ (inputs[406]);
    assign layer0_outputs[5220] = ~(inputs[294]);
    assign layer0_outputs[5221] = inputs[617];
    assign layer0_outputs[5222] = 1'b1;
    assign layer0_outputs[5223] = ~(inputs[792]);
    assign layer0_outputs[5224] = (inputs[3]) ^ (inputs[400]);
    assign layer0_outputs[5225] = (inputs[481]) ^ (inputs[276]);
    assign layer0_outputs[5226] = ~(inputs[807]);
    assign layer0_outputs[5227] = (inputs[719]) & ~(inputs[518]);
    assign layer0_outputs[5228] = (inputs[380]) ^ (inputs[712]);
    assign layer0_outputs[5229] = ~(inputs[743]);
    assign layer0_outputs[5230] = 1'b0;
    assign layer0_outputs[5231] = (inputs[195]) ^ (inputs[494]);
    assign layer0_outputs[5232] = ~(inputs[241]);
    assign layer0_outputs[5233] = ~(inputs[798]);
    assign layer0_outputs[5234] = ~(inputs[511]);
    assign layer0_outputs[5235] = ~(inputs[348]) | (inputs[769]);
    assign layer0_outputs[5236] = (inputs[508]) & ~(inputs[324]);
    assign layer0_outputs[5237] = inputs[242];
    assign layer0_outputs[5238] = ~((inputs[566]) ^ (inputs[479]));
    assign layer0_outputs[5239] = inputs[556];
    assign layer0_outputs[5240] = (inputs[1013]) | (inputs[981]);
    assign layer0_outputs[5241] = (inputs[351]) ^ (inputs[651]);
    assign layer0_outputs[5242] = (inputs[261]) ^ (inputs[480]);
    assign layer0_outputs[5243] = (inputs[1021]) | (inputs[289]);
    assign layer0_outputs[5244] = (inputs[870]) | (inputs[328]);
    assign layer0_outputs[5245] = (inputs[145]) ^ (inputs[610]);
    assign layer0_outputs[5246] = (inputs[496]) | (inputs[871]);
    assign layer0_outputs[5247] = ~(inputs[911]) | (inputs[797]);
    assign layer0_outputs[5248] = inputs[338];
    assign layer0_outputs[5249] = (inputs[166]) ^ (inputs[948]);
    assign layer0_outputs[5250] = (inputs[935]) | (inputs[690]);
    assign layer0_outputs[5251] = ~((inputs[946]) ^ (inputs[739]));
    assign layer0_outputs[5252] = (inputs[522]) | (inputs[725]);
    assign layer0_outputs[5253] = ~(inputs[389]);
    assign layer0_outputs[5254] = ~(inputs[475]);
    assign layer0_outputs[5255] = ~((inputs[750]) | (inputs[420]));
    assign layer0_outputs[5256] = (inputs[525]) & ~(inputs[860]);
    assign layer0_outputs[5257] = ~((inputs[543]) ^ (inputs[319]));
    assign layer0_outputs[5258] = ~(inputs[367]);
    assign layer0_outputs[5259] = ~(inputs[97]) | (inputs[931]);
    assign layer0_outputs[5260] = (inputs[876]) & ~(inputs[640]);
    assign layer0_outputs[5261] = ~((inputs[192]) ^ (inputs[533]));
    assign layer0_outputs[5262] = ~((inputs[150]) | (inputs[94]));
    assign layer0_outputs[5263] = 1'b0;
    assign layer0_outputs[5264] = (inputs[13]) ^ (inputs[805]);
    assign layer0_outputs[5265] = (inputs[708]) | (inputs[266]);
    assign layer0_outputs[5266] = 1'b0;
    assign layer0_outputs[5267] = ~((inputs[444]) ^ (inputs[632]));
    assign layer0_outputs[5268] = ~((inputs[62]) & (inputs[936]));
    assign layer0_outputs[5269] = 1'b0;
    assign layer0_outputs[5270] = ~((inputs[819]) | (inputs[330]));
    assign layer0_outputs[5271] = (inputs[377]) ^ (inputs[371]);
    assign layer0_outputs[5272] = (inputs[720]) ^ (inputs[607]);
    assign layer0_outputs[5273] = 1'b0;
    assign layer0_outputs[5274] = (inputs[985]) & ~(inputs[967]);
    assign layer0_outputs[5275] = (inputs[751]) ^ (inputs[946]);
    assign layer0_outputs[5276] = ~(inputs[503]);
    assign layer0_outputs[5277] = (inputs[298]) | (inputs[768]);
    assign layer0_outputs[5278] = ~(inputs[568]) | (inputs[251]);
    assign layer0_outputs[5279] = (inputs[30]) ^ (inputs[115]);
    assign layer0_outputs[5280] = inputs[329];
    assign layer0_outputs[5281] = ~((inputs[608]) & (inputs[980]));
    assign layer0_outputs[5282] = (inputs[811]) & ~(inputs[415]);
    assign layer0_outputs[5283] = ~(inputs[213]);
    assign layer0_outputs[5284] = ~(inputs[118]);
    assign layer0_outputs[5285] = ~(inputs[551]);
    assign layer0_outputs[5286] = ~((inputs[513]) & (inputs[320]));
    assign layer0_outputs[5287] = inputs[253];
    assign layer0_outputs[5288] = inputs[272];
    assign layer0_outputs[5289] = ~(inputs[444]) | (inputs[449]);
    assign layer0_outputs[5290] = ~(inputs[331]);
    assign layer0_outputs[5291] = ~(inputs[282]);
    assign layer0_outputs[5292] = ~((inputs[353]) ^ (inputs[1010]));
    assign layer0_outputs[5293] = (inputs[989]) & (inputs[453]);
    assign layer0_outputs[5294] = ~(inputs[827]);
    assign layer0_outputs[5295] = ~(inputs[996]);
    assign layer0_outputs[5296] = (inputs[109]) ^ (inputs[618]);
    assign layer0_outputs[5297] = (inputs[599]) | (inputs[630]);
    assign layer0_outputs[5298] = ~(inputs[27]) | (inputs[803]);
    assign layer0_outputs[5299] = (inputs[883]) & ~(inputs[75]);
    assign layer0_outputs[5300] = ~(inputs[666]) | (inputs[892]);
    assign layer0_outputs[5301] = (inputs[441]) ^ (inputs[597]);
    assign layer0_outputs[5302] = ~((inputs[153]) & (inputs[735]));
    assign layer0_outputs[5303] = ~((inputs[747]) | (inputs[775]));
    assign layer0_outputs[5304] = ~((inputs[680]) ^ (inputs[362]));
    assign layer0_outputs[5305] = (inputs[415]) | (inputs[214]);
    assign layer0_outputs[5306] = 1'b1;
    assign layer0_outputs[5307] = ~(inputs[781]) | (inputs[901]);
    assign layer0_outputs[5308] = ~(inputs[124]);
    assign layer0_outputs[5309] = ~(inputs[23]) | (inputs[118]);
    assign layer0_outputs[5310] = ~(inputs[390]) | (inputs[137]);
    assign layer0_outputs[5311] = ~(inputs[641]) | (inputs[952]);
    assign layer0_outputs[5312] = (inputs[564]) | (inputs[764]);
    assign layer0_outputs[5313] = inputs[172];
    assign layer0_outputs[5314] = (inputs[119]) | (inputs[634]);
    assign layer0_outputs[5315] = (inputs[843]) & ~(inputs[109]);
    assign layer0_outputs[5316] = (inputs[863]) | (inputs[238]);
    assign layer0_outputs[5317] = ~(inputs[656]);
    assign layer0_outputs[5318] = inputs[879];
    assign layer0_outputs[5319] = (inputs[139]) & ~(inputs[66]);
    assign layer0_outputs[5320] = ~((inputs[26]) ^ (inputs[918]));
    assign layer0_outputs[5321] = (inputs[944]) | (inputs[394]);
    assign layer0_outputs[5322] = ~(inputs[584]) | (inputs[144]);
    assign layer0_outputs[5323] = (inputs[908]) | (inputs[257]);
    assign layer0_outputs[5324] = 1'b1;
    assign layer0_outputs[5325] = ~((inputs[243]) | (inputs[117]));
    assign layer0_outputs[5326] = (inputs[467]) | (inputs[517]);
    assign layer0_outputs[5327] = (inputs[823]) | (inputs[965]);
    assign layer0_outputs[5328] = ~(inputs[498]) | (inputs[118]);
    assign layer0_outputs[5329] = (inputs[109]) ^ (inputs[607]);
    assign layer0_outputs[5330] = ~(inputs[559]);
    assign layer0_outputs[5331] = ~((inputs[770]) & (inputs[951]));
    assign layer0_outputs[5332] = 1'b0;
    assign layer0_outputs[5333] = inputs[795];
    assign layer0_outputs[5334] = ~((inputs[876]) ^ (inputs[579]));
    assign layer0_outputs[5335] = (inputs[618]) ^ (inputs[106]);
    assign layer0_outputs[5336] = (inputs[250]) ^ (inputs[379]);
    assign layer0_outputs[5337] = (inputs[203]) & ~(inputs[248]);
    assign layer0_outputs[5338] = ~(inputs[631]) | (inputs[283]);
    assign layer0_outputs[5339] = inputs[398];
    assign layer0_outputs[5340] = (inputs[730]) | (inputs[280]);
    assign layer0_outputs[5341] = (inputs[761]) | (inputs[477]);
    assign layer0_outputs[5342] = (inputs[993]) | (inputs[219]);
    assign layer0_outputs[5343] = ~(inputs[352]);
    assign layer0_outputs[5344] = inputs[747];
    assign layer0_outputs[5345] = ~((inputs[736]) | (inputs[748]));
    assign layer0_outputs[5346] = (inputs[189]) & (inputs[675]);
    assign layer0_outputs[5347] = ~((inputs[346]) ^ (inputs[996]));
    assign layer0_outputs[5348] = ~(inputs[793]) | (inputs[121]);
    assign layer0_outputs[5349] = (inputs[376]) & ~(inputs[44]);
    assign layer0_outputs[5350] = inputs[998];
    assign layer0_outputs[5351] = 1'b0;
    assign layer0_outputs[5352] = (inputs[642]) & ~(inputs[800]);
    assign layer0_outputs[5353] = ~(inputs[731]) | (inputs[102]);
    assign layer0_outputs[5354] = ~(inputs[546]);
    assign layer0_outputs[5355] = (inputs[537]) & ~(inputs[639]);
    assign layer0_outputs[5356] = ~(inputs[725]);
    assign layer0_outputs[5357] = inputs[753];
    assign layer0_outputs[5358] = ~((inputs[882]) | (inputs[827]));
    assign layer0_outputs[5359] = inputs[208];
    assign layer0_outputs[5360] = (inputs[323]) | (inputs[377]);
    assign layer0_outputs[5361] = ~(inputs[132]);
    assign layer0_outputs[5362] = inputs[813];
    assign layer0_outputs[5363] = (inputs[603]) & ~(inputs[798]);
    assign layer0_outputs[5364] = (inputs[118]) | (inputs[621]);
    assign layer0_outputs[5365] = ~(inputs[144]);
    assign layer0_outputs[5366] = ~(inputs[157]);
    assign layer0_outputs[5367] = ~(inputs[723]);
    assign layer0_outputs[5368] = (inputs[42]) ^ (inputs[810]);
    assign layer0_outputs[5369] = 1'b1;
    assign layer0_outputs[5370] = inputs[729];
    assign layer0_outputs[5371] = ~((inputs[478]) | (inputs[910]));
    assign layer0_outputs[5372] = inputs[314];
    assign layer0_outputs[5373] = (inputs[349]) | (inputs[781]);
    assign layer0_outputs[5374] = (inputs[840]) | (inputs[754]);
    assign layer0_outputs[5375] = ~(inputs[667]) | (inputs[83]);
    assign layer0_outputs[5376] = (inputs[574]) | (inputs[391]);
    assign layer0_outputs[5377] = ~((inputs[366]) ^ (inputs[1019]));
    assign layer0_outputs[5378] = (inputs[967]) ^ (inputs[343]);
    assign layer0_outputs[5379] = (inputs[226]) & ~(inputs[984]);
    assign layer0_outputs[5380] = (inputs[900]) ^ (inputs[326]);
    assign layer0_outputs[5381] = ~(inputs[186]) | (inputs[144]);
    assign layer0_outputs[5382] = inputs[673];
    assign layer0_outputs[5383] = ~(inputs[376]);
    assign layer0_outputs[5384] = (inputs[968]) ^ (inputs[289]);
    assign layer0_outputs[5385] = ~(inputs[742]);
    assign layer0_outputs[5386] = inputs[531];
    assign layer0_outputs[5387] = ~((inputs[199]) | (inputs[588]));
    assign layer0_outputs[5388] = inputs[974];
    assign layer0_outputs[5389] = ~((inputs[332]) | (inputs[730]));
    assign layer0_outputs[5390] = ~((inputs[803]) | (inputs[614]));
    assign layer0_outputs[5391] = ~((inputs[229]) & (inputs[632]));
    assign layer0_outputs[5392] = inputs[463];
    assign layer0_outputs[5393] = inputs[589];
    assign layer0_outputs[5394] = ~((inputs[385]) ^ (inputs[584]));
    assign layer0_outputs[5395] = ~((inputs[749]) | (inputs[137]));
    assign layer0_outputs[5396] = (inputs[245]) & ~(inputs[567]);
    assign layer0_outputs[5397] = (inputs[939]) | (inputs[942]);
    assign layer0_outputs[5398] = (inputs[733]) ^ (inputs[38]);
    assign layer0_outputs[5399] = inputs[662];
    assign layer0_outputs[5400] = ~((inputs[948]) | (inputs[566]));
    assign layer0_outputs[5401] = (inputs[1016]) & ~(inputs[515]);
    assign layer0_outputs[5402] = ~(inputs[430]);
    assign layer0_outputs[5403] = inputs[449];
    assign layer0_outputs[5404] = (inputs[174]) & ~(inputs[976]);
    assign layer0_outputs[5405] = ~((inputs[201]) | (inputs[747]));
    assign layer0_outputs[5406] = (inputs[69]) & (inputs[735]);
    assign layer0_outputs[5407] = ~((inputs[294]) | (inputs[595]));
    assign layer0_outputs[5408] = (inputs[39]) ^ (inputs[887]);
    assign layer0_outputs[5409] = (inputs[820]) & ~(inputs[1004]);
    assign layer0_outputs[5410] = (inputs[395]) ^ (inputs[1015]);
    assign layer0_outputs[5411] = ~((inputs[790]) | (inputs[352]));
    assign layer0_outputs[5412] = ~(inputs[493]);
    assign layer0_outputs[5413] = (inputs[212]) | (inputs[351]);
    assign layer0_outputs[5414] = ~(inputs[804]);
    assign layer0_outputs[5415] = inputs[721];
    assign layer0_outputs[5416] = ~(inputs[587]) | (inputs[859]);
    assign layer0_outputs[5417] = ~(inputs[430]) | (inputs[734]);
    assign layer0_outputs[5418] = (inputs[886]) ^ (inputs[982]);
    assign layer0_outputs[5419] = (inputs[345]) & ~(inputs[140]);
    assign layer0_outputs[5420] = (inputs[297]) & ~(inputs[180]);
    assign layer0_outputs[5421] = (inputs[234]) | (inputs[772]);
    assign layer0_outputs[5422] = ~(inputs[362]) | (inputs[668]);
    assign layer0_outputs[5423] = (inputs[18]) & ~(inputs[19]);
    assign layer0_outputs[5424] = (inputs[685]) | (inputs[80]);
    assign layer0_outputs[5425] = inputs[627];
    assign layer0_outputs[5426] = ~((inputs[724]) ^ (inputs[75]));
    assign layer0_outputs[5427] = ~((inputs[21]) ^ (inputs[480]));
    assign layer0_outputs[5428] = ~(inputs[785]) | (inputs[764]);
    assign layer0_outputs[5429] = (inputs[659]) & ~(inputs[362]);
    assign layer0_outputs[5430] = (inputs[152]) | (inputs[461]);
    assign layer0_outputs[5431] = ~((inputs[90]) ^ (inputs[656]));
    assign layer0_outputs[5432] = ~(inputs[242]);
    assign layer0_outputs[5433] = inputs[375];
    assign layer0_outputs[5434] = inputs[339];
    assign layer0_outputs[5435] = (inputs[472]) ^ (inputs[82]);
    assign layer0_outputs[5436] = (inputs[334]) & ~(inputs[670]);
    assign layer0_outputs[5437] = ~(inputs[1022]);
    assign layer0_outputs[5438] = ~((inputs[625]) | (inputs[795]));
    assign layer0_outputs[5439] = ~(inputs[432]);
    assign layer0_outputs[5440] = ~(inputs[906]);
    assign layer0_outputs[5441] = ~(inputs[553]) | (inputs[793]);
    assign layer0_outputs[5442] = ~((inputs[48]) ^ (inputs[708]));
    assign layer0_outputs[5443] = (inputs[568]) | (inputs[792]);
    assign layer0_outputs[5444] = ~(inputs[471]);
    assign layer0_outputs[5445] = (inputs[454]) | (inputs[939]);
    assign layer0_outputs[5446] = inputs[163];
    assign layer0_outputs[5447] = ~((inputs[950]) ^ (inputs[161]));
    assign layer0_outputs[5448] = ~(inputs[363]);
    assign layer0_outputs[5449] = ~(inputs[706]);
    assign layer0_outputs[5450] = (inputs[676]) | (inputs[534]);
    assign layer0_outputs[5451] = (inputs[649]) & ~(inputs[677]);
    assign layer0_outputs[5452] = ~((inputs[147]) | (inputs[372]));
    assign layer0_outputs[5453] = (inputs[190]) | (inputs[678]);
    assign layer0_outputs[5454] = (inputs[638]) & (inputs[967]);
    assign layer0_outputs[5455] = (inputs[138]) & ~(inputs[581]);
    assign layer0_outputs[5456] = (inputs[288]) ^ (inputs[993]);
    assign layer0_outputs[5457] = ~(inputs[465]);
    assign layer0_outputs[5458] = (inputs[52]) & (inputs[161]);
    assign layer0_outputs[5459] = (inputs[290]) ^ (inputs[380]);
    assign layer0_outputs[5460] = ~(inputs[498]);
    assign layer0_outputs[5461] = (inputs[192]) & ~(inputs[41]);
    assign layer0_outputs[5462] = ~((inputs[534]) | (inputs[576]));
    assign layer0_outputs[5463] = ~(inputs[272]) | (inputs[219]);
    assign layer0_outputs[5464] = inputs[556];
    assign layer0_outputs[5465] = (inputs[800]) ^ (inputs[370]);
    assign layer0_outputs[5466] = inputs[715];
    assign layer0_outputs[5467] = ~(inputs[779]) | (inputs[282]);
    assign layer0_outputs[5468] = 1'b0;
    assign layer0_outputs[5469] = ~(inputs[882]);
    assign layer0_outputs[5470] = (inputs[75]) ^ (inputs[332]);
    assign layer0_outputs[5471] = inputs[462];
    assign layer0_outputs[5472] = ~(inputs[568]);
    assign layer0_outputs[5473] = inputs[716];
    assign layer0_outputs[5474] = ~((inputs[863]) & (inputs[541]));
    assign layer0_outputs[5475] = 1'b0;
    assign layer0_outputs[5476] = ~(inputs[546]);
    assign layer0_outputs[5477] = ~((inputs[881]) ^ (inputs[646]));
    assign layer0_outputs[5478] = ~(inputs[523]) | (inputs[272]);
    assign layer0_outputs[5479] = (inputs[84]) ^ (inputs[44]);
    assign layer0_outputs[5480] = (inputs[814]) & ~(inputs[60]);
    assign layer0_outputs[5481] = inputs[583];
    assign layer0_outputs[5482] = (inputs[196]) & ~(inputs[825]);
    assign layer0_outputs[5483] = ~(inputs[652]);
    assign layer0_outputs[5484] = (inputs[978]) | (inputs[7]);
    assign layer0_outputs[5485] = 1'b0;
    assign layer0_outputs[5486] = ~(inputs[883]) | (inputs[705]);
    assign layer0_outputs[5487] = (inputs[675]) | (inputs[615]);
    assign layer0_outputs[5488] = (inputs[287]) & ~(inputs[2]);
    assign layer0_outputs[5489] = ~((inputs[402]) ^ (inputs[723]));
    assign layer0_outputs[5490] = ~((inputs[483]) | (inputs[610]));
    assign layer0_outputs[5491] = ~((inputs[541]) | (inputs[57]));
    assign layer0_outputs[5492] = (inputs[431]) & ~(inputs[898]);
    assign layer0_outputs[5493] = ~(inputs[153]) | (inputs[385]);
    assign layer0_outputs[5494] = ~(inputs[521]) | (inputs[913]);
    assign layer0_outputs[5495] = (inputs[204]) & ~(inputs[801]);
    assign layer0_outputs[5496] = inputs[842];
    assign layer0_outputs[5497] = ~((inputs[229]) ^ (inputs[92]));
    assign layer0_outputs[5498] = ~((inputs[118]) | (inputs[651]));
    assign layer0_outputs[5499] = ~((inputs[963]) | (inputs[919]));
    assign layer0_outputs[5500] = ~((inputs[178]) | (inputs[345]));
    assign layer0_outputs[5501] = (inputs[609]) & (inputs[160]);
    assign layer0_outputs[5502] = ~((inputs[266]) | (inputs[373]));
    assign layer0_outputs[5503] = ~(inputs[197]) | (inputs[321]);
    assign layer0_outputs[5504] = ~(inputs[649]) | (inputs[917]);
    assign layer0_outputs[5505] = 1'b1;
    assign layer0_outputs[5506] = (inputs[166]) | (inputs[980]);
    assign layer0_outputs[5507] = ~(inputs[272]);
    assign layer0_outputs[5508] = ~(inputs[442]);
    assign layer0_outputs[5509] = 1'b0;
    assign layer0_outputs[5510] = (inputs[399]) & ~(inputs[944]);
    assign layer0_outputs[5511] = ~((inputs[321]) ^ (inputs[703]));
    assign layer0_outputs[5512] = ~((inputs[1]) ^ (inputs[792]));
    assign layer0_outputs[5513] = (inputs[658]) ^ (inputs[802]);
    assign layer0_outputs[5514] = (inputs[918]) | (inputs[209]);
    assign layer0_outputs[5515] = 1'b1;
    assign layer0_outputs[5516] = (inputs[1016]) & ~(inputs[737]);
    assign layer0_outputs[5517] = 1'b1;
    assign layer0_outputs[5518] = ~((inputs[438]) ^ (inputs[530]));
    assign layer0_outputs[5519] = ~(inputs[599]) | (inputs[481]);
    assign layer0_outputs[5520] = ~((inputs[313]) | (inputs[268]));
    assign layer0_outputs[5521] = 1'b1;
    assign layer0_outputs[5522] = inputs[529];
    assign layer0_outputs[5523] = ~((inputs[99]) | (inputs[946]));
    assign layer0_outputs[5524] = (inputs[369]) | (inputs[580]);
    assign layer0_outputs[5525] = (inputs[57]) ^ (inputs[960]);
    assign layer0_outputs[5526] = ~((inputs[347]) ^ (inputs[728]));
    assign layer0_outputs[5527] = ~((inputs[420]) | (inputs[186]));
    assign layer0_outputs[5528] = ~((inputs[316]) | (inputs[409]));
    assign layer0_outputs[5529] = inputs[597];
    assign layer0_outputs[5530] = ~(inputs[656]);
    assign layer0_outputs[5531] = (inputs[17]) ^ (inputs[189]);
    assign layer0_outputs[5532] = ~((inputs[383]) ^ (inputs[334]));
    assign layer0_outputs[5533] = inputs[522];
    assign layer0_outputs[5534] = inputs[426];
    assign layer0_outputs[5535] = ~((inputs[300]) ^ (inputs[103]));
    assign layer0_outputs[5536] = ~(inputs[650]) | (inputs[155]);
    assign layer0_outputs[5537] = inputs[399];
    assign layer0_outputs[5538] = inputs[90];
    assign layer0_outputs[5539] = 1'b1;
    assign layer0_outputs[5540] = (inputs[237]) & ~(inputs[176]);
    assign layer0_outputs[5541] = inputs[174];
    assign layer0_outputs[5542] = (inputs[602]) & ~(inputs[895]);
    assign layer0_outputs[5543] = inputs[932];
    assign layer0_outputs[5544] = ~(inputs[945]);
    assign layer0_outputs[5545] = ~(inputs[296]);
    assign layer0_outputs[5546] = (inputs[299]) | (inputs[210]);
    assign layer0_outputs[5547] = inputs[715];
    assign layer0_outputs[5548] = ~(inputs[224]);
    assign layer0_outputs[5549] = inputs[246];
    assign layer0_outputs[5550] = (inputs[112]) ^ (inputs[48]);
    assign layer0_outputs[5551] = (inputs[109]) ^ (inputs[734]);
    assign layer0_outputs[5552] = ~((inputs[696]) ^ (inputs[312]));
    assign layer0_outputs[5553] = (inputs[433]) & ~(inputs[881]);
    assign layer0_outputs[5554] = ~(inputs[123]) | (inputs[155]);
    assign layer0_outputs[5555] = (inputs[41]) ^ (inputs[704]);
    assign layer0_outputs[5556] = ~((inputs[914]) | (inputs[423]));
    assign layer0_outputs[5557] = ~(inputs[277]);
    assign layer0_outputs[5558] = ~(inputs[209]) | (inputs[486]);
    assign layer0_outputs[5559] = ~(inputs[779]) | (inputs[827]);
    assign layer0_outputs[5560] = (inputs[87]) ^ (inputs[146]);
    assign layer0_outputs[5561] = ~(inputs[162]);
    assign layer0_outputs[5562] = (inputs[992]) & ~(inputs[579]);
    assign layer0_outputs[5563] = (inputs[148]) & ~(inputs[644]);
    assign layer0_outputs[5564] = inputs[648];
    assign layer0_outputs[5565] = (inputs[121]) & ~(inputs[546]);
    assign layer0_outputs[5566] = inputs[308];
    assign layer0_outputs[5567] = (inputs[21]) & ~(inputs[974]);
    assign layer0_outputs[5568] = ~((inputs[916]) ^ (inputs[771]));
    assign layer0_outputs[5569] = ~(inputs[435]);
    assign layer0_outputs[5570] = 1'b0;
    assign layer0_outputs[5571] = inputs[552];
    assign layer0_outputs[5572] = ~((inputs[451]) ^ (inputs[425]));
    assign layer0_outputs[5573] = ~(inputs[979]);
    assign layer0_outputs[5574] = (inputs[561]) & ~(inputs[137]);
    assign layer0_outputs[5575] = (inputs[654]) & ~(inputs[953]);
    assign layer0_outputs[5576] = 1'b0;
    assign layer0_outputs[5577] = (inputs[778]) ^ (inputs[905]);
    assign layer0_outputs[5578] = (inputs[968]) | (inputs[841]);
    assign layer0_outputs[5579] = ~((inputs[317]) & (inputs[895]));
    assign layer0_outputs[5580] = ~(inputs[523]) | (inputs[30]);
    assign layer0_outputs[5581] = ~((inputs[622]) | (inputs[265]));
    assign layer0_outputs[5582] = ~(inputs[911]);
    assign layer0_outputs[5583] = inputs[398];
    assign layer0_outputs[5584] = (inputs[42]) ^ (inputs[447]);
    assign layer0_outputs[5585] = (inputs[472]) ^ (inputs[31]);
    assign layer0_outputs[5586] = ~((inputs[212]) | (inputs[653]));
    assign layer0_outputs[5587] = inputs[627];
    assign layer0_outputs[5588] = ~(inputs[419]);
    assign layer0_outputs[5589] = ~(inputs[658]) | (inputs[837]);
    assign layer0_outputs[5590] = (inputs[302]) | (inputs[73]);
    assign layer0_outputs[5591] = inputs[805];
    assign layer0_outputs[5592] = ~(inputs[228]);
    assign layer0_outputs[5593] = (inputs[686]) & (inputs[719]);
    assign layer0_outputs[5594] = ~((inputs[554]) | (inputs[58]));
    assign layer0_outputs[5595] = ~(inputs[330]);
    assign layer0_outputs[5596] = (inputs[814]) | (inputs[873]);
    assign layer0_outputs[5597] = ~((inputs[436]) ^ (inputs[612]));
    assign layer0_outputs[5598] = (inputs[143]) | (inputs[121]);
    assign layer0_outputs[5599] = ~((inputs[295]) | (inputs[991]));
    assign layer0_outputs[5600] = ~((inputs[611]) | (inputs[651]));
    assign layer0_outputs[5601] = inputs[141];
    assign layer0_outputs[5602] = ~(inputs[401]) | (inputs[708]);
    assign layer0_outputs[5603] = inputs[355];
    assign layer0_outputs[5604] = ~(inputs[359]) | (inputs[1023]);
    assign layer0_outputs[5605] = ~(inputs[710]);
    assign layer0_outputs[5606] = (inputs[397]) ^ (inputs[72]);
    assign layer0_outputs[5607] = ~((inputs[428]) ^ (inputs[487]));
    assign layer0_outputs[5608] = inputs[402];
    assign layer0_outputs[5609] = inputs[845];
    assign layer0_outputs[5610] = ~((inputs[214]) | (inputs[576]));
    assign layer0_outputs[5611] = (inputs[24]) | (inputs[569]);
    assign layer0_outputs[5612] = ~((inputs[141]) | (inputs[6]));
    assign layer0_outputs[5613] = ~(inputs[208]);
    assign layer0_outputs[5614] = (inputs[960]) ^ (inputs[545]);
    assign layer0_outputs[5615] = ~(inputs[852]);
    assign layer0_outputs[5616] = ~(inputs[146]) | (inputs[346]);
    assign layer0_outputs[5617] = ~((inputs[393]) | (inputs[212]));
    assign layer0_outputs[5618] = ~((inputs[469]) | (inputs[612]));
    assign layer0_outputs[5619] = ~(inputs[247]);
    assign layer0_outputs[5620] = ~((inputs[1017]) ^ (inputs[61]));
    assign layer0_outputs[5621] = ~(inputs[175]);
    assign layer0_outputs[5622] = ~(inputs[926]);
    assign layer0_outputs[5623] = ~((inputs[689]) | (inputs[714]));
    assign layer0_outputs[5624] = (inputs[97]) & (inputs[1015]);
    assign layer0_outputs[5625] = ~(inputs[970]) | (inputs[25]);
    assign layer0_outputs[5626] = ~(inputs[622]);
    assign layer0_outputs[5627] = ~((inputs[655]) | (inputs[17]));
    assign layer0_outputs[5628] = inputs[979];
    assign layer0_outputs[5629] = (inputs[84]) ^ (inputs[519]);
    assign layer0_outputs[5630] = inputs[941];
    assign layer0_outputs[5631] = (inputs[670]) & ~(inputs[223]);
    assign layer0_outputs[5632] = ~(inputs[669]);
    assign layer0_outputs[5633] = (inputs[17]) | (inputs[661]);
    assign layer0_outputs[5634] = ~((inputs[169]) | (inputs[238]));
    assign layer0_outputs[5635] = ~(inputs[214]);
    assign layer0_outputs[5636] = (inputs[50]) ^ (inputs[848]);
    assign layer0_outputs[5637] = ~((inputs[417]) | (inputs[97]));
    assign layer0_outputs[5638] = (inputs[340]) & ~(inputs[788]);
    assign layer0_outputs[5639] = inputs[75];
    assign layer0_outputs[5640] = ~(inputs[688]) | (inputs[695]);
    assign layer0_outputs[5641] = inputs[636];
    assign layer0_outputs[5642] = inputs[895];
    assign layer0_outputs[5643] = inputs[818];
    assign layer0_outputs[5644] = (inputs[949]) | (inputs[918]);
    assign layer0_outputs[5645] = ~(inputs[188]);
    assign layer0_outputs[5646] = (inputs[633]) | (inputs[810]);
    assign layer0_outputs[5647] = inputs[950];
    assign layer0_outputs[5648] = ~(inputs[681]);
    assign layer0_outputs[5649] = (inputs[125]) | (inputs[811]);
    assign layer0_outputs[5650] = (inputs[843]) & ~(inputs[140]);
    assign layer0_outputs[5651] = (inputs[1015]) ^ (inputs[905]);
    assign layer0_outputs[5652] = ~((inputs[801]) | (inputs[455]));
    assign layer0_outputs[5653] = 1'b1;
    assign layer0_outputs[5654] = ~(inputs[397]);
    assign layer0_outputs[5655] = ~((inputs[603]) | (inputs[776]));
    assign layer0_outputs[5656] = ~((inputs[44]) | (inputs[862]));
    assign layer0_outputs[5657] = (inputs[863]) & ~(inputs[852]);
    assign layer0_outputs[5658] = ~(inputs[54]) | (inputs[126]);
    assign layer0_outputs[5659] = inputs[682];
    assign layer0_outputs[5660] = inputs[436];
    assign layer0_outputs[5661] = (inputs[114]) | (inputs[729]);
    assign layer0_outputs[5662] = (inputs[1011]) ^ (inputs[435]);
    assign layer0_outputs[5663] = ~((inputs[237]) ^ (inputs[535]));
    assign layer0_outputs[5664] = (inputs[958]) ^ (inputs[434]);
    assign layer0_outputs[5665] = ~(inputs[527]);
    assign layer0_outputs[5666] = ~((inputs[789]) ^ (inputs[834]));
    assign layer0_outputs[5667] = (inputs[632]) | (inputs[838]);
    assign layer0_outputs[5668] = (inputs[379]) | (inputs[252]);
    assign layer0_outputs[5669] = ~((inputs[804]) ^ (inputs[115]));
    assign layer0_outputs[5670] = 1'b1;
    assign layer0_outputs[5671] = ~(inputs[950]);
    assign layer0_outputs[5672] = ~((inputs[850]) | (inputs[347]));
    assign layer0_outputs[5673] = 1'b1;
    assign layer0_outputs[5674] = 1'b0;
    assign layer0_outputs[5675] = inputs[429];
    assign layer0_outputs[5676] = ~(inputs[564]) | (inputs[961]);
    assign layer0_outputs[5677] = 1'b0;
    assign layer0_outputs[5678] = ~((inputs[63]) ^ (inputs[918]));
    assign layer0_outputs[5679] = (inputs[822]) & ~(inputs[516]);
    assign layer0_outputs[5680] = ~((inputs[879]) ^ (inputs[251]));
    assign layer0_outputs[5681] = ~(inputs[723]) | (inputs[319]);
    assign layer0_outputs[5682] = (inputs[825]) ^ (inputs[338]);
    assign layer0_outputs[5683] = ~((inputs[148]) | (inputs[146]));
    assign layer0_outputs[5684] = ~((inputs[675]) & (inputs[67]));
    assign layer0_outputs[5685] = ~((inputs[508]) ^ (inputs[677]));
    assign layer0_outputs[5686] = inputs[825];
    assign layer0_outputs[5687] = ~((inputs[20]) ^ (inputs[479]));
    assign layer0_outputs[5688] = ~(inputs[880]);
    assign layer0_outputs[5689] = (inputs[68]) | (inputs[887]);
    assign layer0_outputs[5690] = (inputs[537]) & ~(inputs[924]);
    assign layer0_outputs[5691] = (inputs[1018]) & ~(inputs[192]);
    assign layer0_outputs[5692] = (inputs[240]) ^ (inputs[107]);
    assign layer0_outputs[5693] = (inputs[718]) & ~(inputs[947]);
    assign layer0_outputs[5694] = ~((inputs[236]) | (inputs[441]));
    assign layer0_outputs[5695] = (inputs[688]) | (inputs[781]);
    assign layer0_outputs[5696] = (inputs[751]) | (inputs[633]);
    assign layer0_outputs[5697] = ~((inputs[917]) ^ (inputs[809]));
    assign layer0_outputs[5698] = ~(inputs[685]);
    assign layer0_outputs[5699] = ~((inputs[402]) | (inputs[49]));
    assign layer0_outputs[5700] = ~(inputs[394]);
    assign layer0_outputs[5701] = ~(inputs[755]);
    assign layer0_outputs[5702] = ~((inputs[640]) | (inputs[374]));
    assign layer0_outputs[5703] = (inputs[593]) & ~(inputs[451]);
    assign layer0_outputs[5704] = ~((inputs[875]) | (inputs[65]));
    assign layer0_outputs[5705] = ~((inputs[773]) | (inputs[905]));
    assign layer0_outputs[5706] = ~(inputs[184]) | (inputs[123]);
    assign layer0_outputs[5707] = ~((inputs[486]) & (inputs[27]));
    assign layer0_outputs[5708] = (inputs[665]) ^ (inputs[497]);
    assign layer0_outputs[5709] = (inputs[284]) ^ (inputs[230]);
    assign layer0_outputs[5710] = (inputs[32]) ^ (inputs[569]);
    assign layer0_outputs[5711] = ~(inputs[743]);
    assign layer0_outputs[5712] = ~((inputs[1014]) | (inputs[27]));
    assign layer0_outputs[5713] = ~(inputs[560]) | (inputs[52]);
    assign layer0_outputs[5714] = (inputs[594]) | (inputs[992]);
    assign layer0_outputs[5715] = (inputs[822]) | (inputs[221]);
    assign layer0_outputs[5716] = inputs[525];
    assign layer0_outputs[5717] = inputs[32];
    assign layer0_outputs[5718] = ~((inputs[916]) ^ (inputs[172]));
    assign layer0_outputs[5719] = (inputs[524]) & ~(inputs[344]);
    assign layer0_outputs[5720] = inputs[351];
    assign layer0_outputs[5721] = ~(inputs[677]) | (inputs[886]);
    assign layer0_outputs[5722] = (inputs[823]) & ~(inputs[198]);
    assign layer0_outputs[5723] = 1'b1;
    assign layer0_outputs[5724] = ~(inputs[701]);
    assign layer0_outputs[5725] = ~(inputs[438]);
    assign layer0_outputs[5726] = ~(inputs[571]) | (inputs[380]);
    assign layer0_outputs[5727] = inputs[56];
    assign layer0_outputs[5728] = inputs[923];
    assign layer0_outputs[5729] = ~(inputs[527]) | (inputs[262]);
    assign layer0_outputs[5730] = (inputs[403]) & ~(inputs[951]);
    assign layer0_outputs[5731] = (inputs[521]) ^ (inputs[193]);
    assign layer0_outputs[5732] = ~(inputs[594]);
    assign layer0_outputs[5733] = inputs[241];
    assign layer0_outputs[5734] = (inputs[590]) & ~(inputs[202]);
    assign layer0_outputs[5735] = inputs[656];
    assign layer0_outputs[5736] = inputs[750];
    assign layer0_outputs[5737] = ~(inputs[832]) | (inputs[862]);
    assign layer0_outputs[5738] = ~((inputs[533]) | (inputs[912]));
    assign layer0_outputs[5739] = (inputs[720]) ^ (inputs[238]);
    assign layer0_outputs[5740] = ~((inputs[770]) ^ (inputs[97]));
    assign layer0_outputs[5741] = ~((inputs[1003]) | (inputs[575]));
    assign layer0_outputs[5742] = ~((inputs[418]) & (inputs[976]));
    assign layer0_outputs[5743] = ~((inputs[443]) | (inputs[107]));
    assign layer0_outputs[5744] = ~((inputs[625]) | (inputs[413]));
    assign layer0_outputs[5745] = (inputs[643]) & ~(inputs[349]);
    assign layer0_outputs[5746] = ~((inputs[772]) | (inputs[148]));
    assign layer0_outputs[5747] = ~((inputs[208]) & (inputs[720]));
    assign layer0_outputs[5748] = (inputs[592]) & ~(inputs[148]);
    assign layer0_outputs[5749] = ~(inputs[401]);
    assign layer0_outputs[5750] = ~(inputs[41]);
    assign layer0_outputs[5751] = (inputs[904]) | (inputs[478]);
    assign layer0_outputs[5752] = ~(inputs[104]);
    assign layer0_outputs[5753] = ~(inputs[951]);
    assign layer0_outputs[5754] = inputs[248];
    assign layer0_outputs[5755] = (inputs[200]) & ~(inputs[24]);
    assign layer0_outputs[5756] = (inputs[774]) | (inputs[107]);
    assign layer0_outputs[5757] = (inputs[1]) & ~(inputs[643]);
    assign layer0_outputs[5758] = ~(inputs[815]);
    assign layer0_outputs[5759] = ~(inputs[695]);
    assign layer0_outputs[5760] = ~(inputs[234]) | (inputs[426]);
    assign layer0_outputs[5761] = ~(inputs[441]);
    assign layer0_outputs[5762] = (inputs[204]) ^ (inputs[296]);
    assign layer0_outputs[5763] = (inputs[138]) & ~(inputs[451]);
    assign layer0_outputs[5764] = inputs[656];
    assign layer0_outputs[5765] = (inputs[619]) & ~(inputs[77]);
    assign layer0_outputs[5766] = 1'b1;
    assign layer0_outputs[5767] = ~((inputs[130]) ^ (inputs[80]));
    assign layer0_outputs[5768] = (inputs[657]) | (inputs[440]);
    assign layer0_outputs[5769] = ~(inputs[755]);
    assign layer0_outputs[5770] = ~(inputs[657]);
    assign layer0_outputs[5771] = (inputs[611]) ^ (inputs[275]);
    assign layer0_outputs[5772] = ~((inputs[463]) | (inputs[366]));
    assign layer0_outputs[5773] = (inputs[83]) | (inputs[205]);
    assign layer0_outputs[5774] = (inputs[276]) | (inputs[857]);
    assign layer0_outputs[5775] = ~((inputs[744]) ^ (inputs[749]));
    assign layer0_outputs[5776] = ~((inputs[378]) | (inputs[189]));
    assign layer0_outputs[5777] = ~(inputs[729]);
    assign layer0_outputs[5778] = ~(inputs[31]);
    assign layer0_outputs[5779] = (inputs[864]) ^ (inputs[314]);
    assign layer0_outputs[5780] = (inputs[76]) | (inputs[437]);
    assign layer0_outputs[5781] = (inputs[1017]) | (inputs[868]);
    assign layer0_outputs[5782] = ~(inputs[340]) | (inputs[391]);
    assign layer0_outputs[5783] = ~(inputs[635]) | (inputs[485]);
    assign layer0_outputs[5784] = 1'b1;
    assign layer0_outputs[5785] = ~((inputs[359]) & (inputs[898]));
    assign layer0_outputs[5786] = ~(inputs[403]) | (inputs[823]);
    assign layer0_outputs[5787] = 1'b0;
    assign layer0_outputs[5788] = (inputs[674]) ^ (inputs[988]);
    assign layer0_outputs[5789] = ~((inputs[596]) | (inputs[170]));
    assign layer0_outputs[5790] = ~(inputs[425]);
    assign layer0_outputs[5791] = ~((inputs[882]) | (inputs[413]));
    assign layer0_outputs[5792] = ~(inputs[226]) | (inputs[543]);
    assign layer0_outputs[5793] = ~(inputs[917]);
    assign layer0_outputs[5794] = (inputs[306]) & ~(inputs[334]);
    assign layer0_outputs[5795] = ~(inputs[933]) | (inputs[89]);
    assign layer0_outputs[5796] = inputs[531];
    assign layer0_outputs[5797] = ~(inputs[139]) | (inputs[60]);
    assign layer0_outputs[5798] = ~((inputs[381]) | (inputs[484]));
    assign layer0_outputs[5799] = (inputs[149]) | (inputs[127]);
    assign layer0_outputs[5800] = ~(inputs[333]);
    assign layer0_outputs[5801] = (inputs[489]) & ~(inputs[936]);
    assign layer0_outputs[5802] = (inputs[714]) | (inputs[699]);
    assign layer0_outputs[5803] = (inputs[494]) & ~(inputs[235]);
    assign layer0_outputs[5804] = ~(inputs[147]) | (inputs[937]);
    assign layer0_outputs[5805] = ~((inputs[941]) ^ (inputs[951]));
    assign layer0_outputs[5806] = ~((inputs[310]) ^ (inputs[50]));
    assign layer0_outputs[5807] = ~(inputs[410]) | (inputs[98]);
    assign layer0_outputs[5808] = (inputs[621]) & ~(inputs[896]);
    assign layer0_outputs[5809] = (inputs[179]) & ~(inputs[359]);
    assign layer0_outputs[5810] = (inputs[111]) | (inputs[438]);
    assign layer0_outputs[5811] = ~((inputs[534]) ^ (inputs[225]));
    assign layer0_outputs[5812] = ~(inputs[69]);
    assign layer0_outputs[5813] = ~((inputs[895]) | (inputs[821]));
    assign layer0_outputs[5814] = ~((inputs[943]) | (inputs[370]));
    assign layer0_outputs[5815] = ~(inputs[907]) | (inputs[639]);
    assign layer0_outputs[5816] = (inputs[381]) & (inputs[569]);
    assign layer0_outputs[5817] = ~(inputs[942]);
    assign layer0_outputs[5818] = (inputs[285]) | (inputs[276]);
    assign layer0_outputs[5819] = (inputs[695]) | (inputs[299]);
    assign layer0_outputs[5820] = ~(inputs[939]) | (inputs[412]);
    assign layer0_outputs[5821] = (inputs[837]) & ~(inputs[16]);
    assign layer0_outputs[5822] = (inputs[762]) & ~(inputs[447]);
    assign layer0_outputs[5823] = (inputs[457]) & (inputs[813]);
    assign layer0_outputs[5824] = inputs[149];
    assign layer0_outputs[5825] = (inputs[284]) | (inputs[365]);
    assign layer0_outputs[5826] = ~((inputs[644]) & (inputs[823]));
    assign layer0_outputs[5827] = (inputs[259]) | (inputs[129]);
    assign layer0_outputs[5828] = 1'b1;
    assign layer0_outputs[5829] = (inputs[398]) | (inputs[432]);
    assign layer0_outputs[5830] = (inputs[683]) & ~(inputs[1010]);
    assign layer0_outputs[5831] = ~(inputs[932]);
    assign layer0_outputs[5832] = ~(inputs[269]);
    assign layer0_outputs[5833] = (inputs[244]) | (inputs[938]);
    assign layer0_outputs[5834] = ~(inputs[619]);
    assign layer0_outputs[5835] = (inputs[957]) | (inputs[658]);
    assign layer0_outputs[5836] = ~(inputs[410]) | (inputs[152]);
    assign layer0_outputs[5837] = (inputs[561]) & ~(inputs[324]);
    assign layer0_outputs[5838] = (inputs[325]) | (inputs[206]);
    assign layer0_outputs[5839] = ~((inputs[439]) | (inputs[362]));
    assign layer0_outputs[5840] = ~(inputs[420]) | (inputs[414]);
    assign layer0_outputs[5841] = ~((inputs[695]) | (inputs[13]));
    assign layer0_outputs[5842] = (inputs[475]) & ~(inputs[553]);
    assign layer0_outputs[5843] = (inputs[824]) & (inputs[169]);
    assign layer0_outputs[5844] = ~(inputs[550]);
    assign layer0_outputs[5845] = ~(inputs[279]);
    assign layer0_outputs[5846] = inputs[878];
    assign layer0_outputs[5847] = ~(inputs[833]);
    assign layer0_outputs[5848] = ~(inputs[947]) | (inputs[921]);
    assign layer0_outputs[5849] = inputs[940];
    assign layer0_outputs[5850] = (inputs[422]) & ~(inputs[443]);
    assign layer0_outputs[5851] = ~(inputs[388]) | (inputs[169]);
    assign layer0_outputs[5852] = (inputs[524]) & ~(inputs[60]);
    assign layer0_outputs[5853] = ~((inputs[871]) | (inputs[538]));
    assign layer0_outputs[5854] = (inputs[565]) | (inputs[304]);
    assign layer0_outputs[5855] = ~((inputs[910]) | (inputs[264]));
    assign layer0_outputs[5856] = ~((inputs[700]) | (inputs[550]));
    assign layer0_outputs[5857] = (inputs[627]) & ~(inputs[919]);
    assign layer0_outputs[5858] = ~(inputs[405]);
    assign layer0_outputs[5859] = inputs[406];
    assign layer0_outputs[5860] = ~(inputs[301]);
    assign layer0_outputs[5861] = (inputs[758]) | (inputs[168]);
    assign layer0_outputs[5862] = ~((inputs[790]) ^ (inputs[600]));
    assign layer0_outputs[5863] = ~((inputs[926]) & (inputs[8]));
    assign layer0_outputs[5864] = ~((inputs[312]) | (inputs[246]));
    assign layer0_outputs[5865] = ~((inputs[976]) ^ (inputs[973]));
    assign layer0_outputs[5866] = ~(inputs[719]);
    assign layer0_outputs[5867] = inputs[654];
    assign layer0_outputs[5868] = (inputs[61]) & ~(inputs[134]);
    assign layer0_outputs[5869] = ~(inputs[408]) | (inputs[43]);
    assign layer0_outputs[5870] = ~(inputs[211]);
    assign layer0_outputs[5871] = ~(inputs[714]) | (inputs[917]);
    assign layer0_outputs[5872] = ~(inputs[339]);
    assign layer0_outputs[5873] = inputs[212];
    assign layer0_outputs[5874] = (inputs[541]) & ~(inputs[331]);
    assign layer0_outputs[5875] = ~(inputs[858]) | (inputs[386]);
    assign layer0_outputs[5876] = (inputs[681]) & ~(inputs[914]);
    assign layer0_outputs[5877] = (inputs[881]) | (inputs[148]);
    assign layer0_outputs[5878] = ~((inputs[400]) | (inputs[814]));
    assign layer0_outputs[5879] = (inputs[205]) ^ (inputs[470]);
    assign layer0_outputs[5880] = inputs[654];
    assign layer0_outputs[5881] = ~((inputs[225]) | (inputs[379]));
    assign layer0_outputs[5882] = ~(inputs[840]);
    assign layer0_outputs[5883] = (inputs[1019]) & (inputs[631]);
    assign layer0_outputs[5884] = ~((inputs[385]) | (inputs[597]));
    assign layer0_outputs[5885] = (inputs[421]) | (inputs[721]);
    assign layer0_outputs[5886] = (inputs[333]) & ~(inputs[481]);
    assign layer0_outputs[5887] = ~(inputs[372]) | (inputs[886]);
    assign layer0_outputs[5888] = (inputs[396]) & ~(inputs[672]);
    assign layer0_outputs[5889] = ~((inputs[928]) ^ (inputs[336]));
    assign layer0_outputs[5890] = inputs[321];
    assign layer0_outputs[5891] = inputs[713];
    assign layer0_outputs[5892] = ~((inputs[354]) | (inputs[380]));
    assign layer0_outputs[5893] = inputs[347];
    assign layer0_outputs[5894] = ~((inputs[317]) | (inputs[887]));
    assign layer0_outputs[5895] = (inputs[930]) & ~(inputs[995]);
    assign layer0_outputs[5896] = (inputs[189]) & ~(inputs[349]);
    assign layer0_outputs[5897] = ~((inputs[383]) & (inputs[1]));
    assign layer0_outputs[5898] = (inputs[758]) | (inputs[174]);
    assign layer0_outputs[5899] = inputs[99];
    assign layer0_outputs[5900] = ~(inputs[971]) | (inputs[158]);
    assign layer0_outputs[5901] = ~(inputs[402]);
    assign layer0_outputs[5902] = ~((inputs[390]) ^ (inputs[767]));
    assign layer0_outputs[5903] = ~((inputs[155]) | (inputs[350]));
    assign layer0_outputs[5904] = (inputs[488]) & ~(inputs[742]);
    assign layer0_outputs[5905] = (inputs[14]) & ~(inputs[635]);
    assign layer0_outputs[5906] = inputs[326];
    assign layer0_outputs[5907] = ~((inputs[152]) ^ (inputs[936]));
    assign layer0_outputs[5908] = ~(inputs[205]) | (inputs[120]);
    assign layer0_outputs[5909] = ~(inputs[336]);
    assign layer0_outputs[5910] = ~((inputs[344]) | (inputs[807]));
    assign layer0_outputs[5911] = (inputs[445]) & ~(inputs[222]);
    assign layer0_outputs[5912] = ~(inputs[336]);
    assign layer0_outputs[5913] = ~((inputs[49]) | (inputs[983]));
    assign layer0_outputs[5914] = (inputs[431]) & ~(inputs[580]);
    assign layer0_outputs[5915] = ~((inputs[124]) | (inputs[124]));
    assign layer0_outputs[5916] = ~((inputs[937]) | (inputs[478]));
    assign layer0_outputs[5917] = 1'b0;
    assign layer0_outputs[5918] = ~(inputs[465]);
    assign layer0_outputs[5919] = ~((inputs[117]) | (inputs[419]));
    assign layer0_outputs[5920] = (inputs[747]) | (inputs[853]);
    assign layer0_outputs[5921] = ~((inputs[217]) | (inputs[990]));
    assign layer0_outputs[5922] = ~(inputs[848]);
    assign layer0_outputs[5923] = inputs[396];
    assign layer0_outputs[5924] = ~((inputs[232]) | (inputs[320]));
    assign layer0_outputs[5925] = (inputs[883]) & ~(inputs[255]);
    assign layer0_outputs[5926] = (inputs[141]) & (inputs[739]);
    assign layer0_outputs[5927] = inputs[437];
    assign layer0_outputs[5928] = inputs[780];
    assign layer0_outputs[5929] = ~((inputs[672]) ^ (inputs[793]));
    assign layer0_outputs[5930] = (inputs[363]) | (inputs[484]);
    assign layer0_outputs[5931] = ~((inputs[787]) & (inputs[801]));
    assign layer0_outputs[5932] = ~(inputs[14]) | (inputs[59]);
    assign layer0_outputs[5933] = inputs[970];
    assign layer0_outputs[5934] = ~(inputs[392]);
    assign layer0_outputs[5935] = (inputs[815]) | (inputs[535]);
    assign layer0_outputs[5936] = ~((inputs[894]) | (inputs[523]));
    assign layer0_outputs[5937] = ~((inputs[43]) | (inputs[747]));
    assign layer0_outputs[5938] = (inputs[888]) | (inputs[710]);
    assign layer0_outputs[5939] = ~(inputs[145]);
    assign layer0_outputs[5940] = 1'b1;
    assign layer0_outputs[5941] = ~(inputs[410]);
    assign layer0_outputs[5942] = (inputs[438]) & ~(inputs[747]);
    assign layer0_outputs[5943] = inputs[239];
    assign layer0_outputs[5944] = ~(inputs[373]) | (inputs[82]);
    assign layer0_outputs[5945] = ~(inputs[368]) | (inputs[434]);
    assign layer0_outputs[5946] = (inputs[134]) | (inputs[113]);
    assign layer0_outputs[5947] = ~(inputs[885]) | (inputs[937]);
    assign layer0_outputs[5948] = inputs[618];
    assign layer0_outputs[5949] = inputs[504];
    assign layer0_outputs[5950] = ~((inputs[223]) ^ (inputs[940]));
    assign layer0_outputs[5951] = (inputs[807]) | (inputs[711]);
    assign layer0_outputs[5952] = (inputs[919]) & ~(inputs[257]);
    assign layer0_outputs[5953] = ~(inputs[117]);
    assign layer0_outputs[5954] = (inputs[736]) & ~(inputs[496]);
    assign layer0_outputs[5955] = ~(inputs[684]);
    assign layer0_outputs[5956] = ~((inputs[649]) | (inputs[459]));
    assign layer0_outputs[5957] = ~((inputs[462]) ^ (inputs[34]));
    assign layer0_outputs[5958] = inputs[278];
    assign layer0_outputs[5959] = (inputs[764]) & ~(inputs[543]);
    assign layer0_outputs[5960] = ~((inputs[891]) | (inputs[628]));
    assign layer0_outputs[5961] = (inputs[66]) & (inputs[197]);
    assign layer0_outputs[5962] = (inputs[664]) & ~(inputs[525]);
    assign layer0_outputs[5963] = (inputs[991]) & (inputs[412]);
    assign layer0_outputs[5964] = ~((inputs[337]) | (inputs[690]));
    assign layer0_outputs[5965] = ~(inputs[702]) | (inputs[196]);
    assign layer0_outputs[5966] = ~((inputs[863]) ^ (inputs[336]));
    assign layer0_outputs[5967] = 1'b1;
    assign layer0_outputs[5968] = (inputs[287]) | (inputs[915]);
    assign layer0_outputs[5969] = (inputs[504]) ^ (inputs[1022]);
    assign layer0_outputs[5970] = (inputs[187]) & ~(inputs[981]);
    assign layer0_outputs[5971] = (inputs[29]) ^ (inputs[662]);
    assign layer0_outputs[5972] = (inputs[738]) ^ (inputs[218]);
    assign layer0_outputs[5973] = 1'b0;
    assign layer0_outputs[5974] = inputs[693];
    assign layer0_outputs[5975] = ~((inputs[655]) ^ (inputs[383]));
    assign layer0_outputs[5976] = ~(inputs[398]) | (inputs[40]);
    assign layer0_outputs[5977] = ~(inputs[362]);
    assign layer0_outputs[5978] = ~(inputs[17]);
    assign layer0_outputs[5979] = (inputs[173]) & ~(inputs[767]);
    assign layer0_outputs[5980] = (inputs[37]) & ~(inputs[902]);
    assign layer0_outputs[5981] = ~(inputs[560]) | (inputs[55]);
    assign layer0_outputs[5982] = (inputs[756]) | (inputs[572]);
    assign layer0_outputs[5983] = ~((inputs[502]) & (inputs[262]));
    assign layer0_outputs[5984] = (inputs[477]) | (inputs[879]);
    assign layer0_outputs[5985] = ~(inputs[309]) | (inputs[604]);
    assign layer0_outputs[5986] = ~(inputs[684]) | (inputs[706]);
    assign layer0_outputs[5987] = ~((inputs[587]) | (inputs[890]));
    assign layer0_outputs[5988] = ~(inputs[772]) | (inputs[262]);
    assign layer0_outputs[5989] = ~(inputs[527]) | (inputs[612]);
    assign layer0_outputs[5990] = (inputs[302]) ^ (inputs[449]);
    assign layer0_outputs[5991] = ~((inputs[513]) ^ (inputs[416]));
    assign layer0_outputs[5992] = ~((inputs[223]) | (inputs[42]));
    assign layer0_outputs[5993] = ~(inputs[515]) | (inputs[897]);
    assign layer0_outputs[5994] = inputs[359];
    assign layer0_outputs[5995] = ~(inputs[910]);
    assign layer0_outputs[5996] = (inputs[843]) ^ (inputs[835]);
    assign layer0_outputs[5997] = ~(inputs[460]) | (inputs[286]);
    assign layer0_outputs[5998] = (inputs[888]) | (inputs[82]);
    assign layer0_outputs[5999] = ~(inputs[597]);
    assign layer0_outputs[6000] = (inputs[312]) ^ (inputs[575]);
    assign layer0_outputs[6001] = inputs[895];
    assign layer0_outputs[6002] = (inputs[319]) | (inputs[460]);
    assign layer0_outputs[6003] = ~(inputs[405]);
    assign layer0_outputs[6004] = (inputs[132]) | (inputs[885]);
    assign layer0_outputs[6005] = (inputs[838]) & ~(inputs[107]);
    assign layer0_outputs[6006] = inputs[719];
    assign layer0_outputs[6007] = ~(inputs[882]) | (inputs[763]);
    assign layer0_outputs[6008] = inputs[650];
    assign layer0_outputs[6009] = ~((inputs[457]) | (inputs[875]));
    assign layer0_outputs[6010] = ~((inputs[45]) | (inputs[973]));
    assign layer0_outputs[6011] = ~(inputs[1]) | (inputs[827]);
    assign layer0_outputs[6012] = ~((inputs[744]) | (inputs[265]));
    assign layer0_outputs[6013] = ~((inputs[951]) ^ (inputs[923]));
    assign layer0_outputs[6014] = ~(inputs[726]) | (inputs[865]);
    assign layer0_outputs[6015] = (inputs[696]) & ~(inputs[384]);
    assign layer0_outputs[6016] = inputs[129];
    assign layer0_outputs[6017] = ~(inputs[370]);
    assign layer0_outputs[6018] = (inputs[270]) & ~(inputs[129]);
    assign layer0_outputs[6019] = ~(inputs[592]) | (inputs[196]);
    assign layer0_outputs[6020] = (inputs[400]) | (inputs[466]);
    assign layer0_outputs[6021] = ~(inputs[581]) | (inputs[579]);
    assign layer0_outputs[6022] = ~(inputs[782]) | (inputs[231]);
    assign layer0_outputs[6023] = ~(inputs[889]);
    assign layer0_outputs[6024] = (inputs[601]) | (inputs[138]);
    assign layer0_outputs[6025] = ~((inputs[628]) | (inputs[972]));
    assign layer0_outputs[6026] = ~(inputs[981]) | (inputs[581]);
    assign layer0_outputs[6027] = inputs[488];
    assign layer0_outputs[6028] = ~((inputs[635]) & (inputs[332]));
    assign layer0_outputs[6029] = ~((inputs[119]) | (inputs[496]));
    assign layer0_outputs[6030] = 1'b1;
    assign layer0_outputs[6031] = (inputs[135]) ^ (inputs[295]);
    assign layer0_outputs[6032] = ~((inputs[753]) ^ (inputs[1021]));
    assign layer0_outputs[6033] = (inputs[174]) | (inputs[32]);
    assign layer0_outputs[6034] = (inputs[44]) ^ (inputs[185]);
    assign layer0_outputs[6035] = (inputs[170]) & ~(inputs[475]);
    assign layer0_outputs[6036] = ~((inputs[508]) | (inputs[980]));
    assign layer0_outputs[6037] = inputs[744];
    assign layer0_outputs[6038] = ~(inputs[628]);
    assign layer0_outputs[6039] = 1'b1;
    assign layer0_outputs[6040] = ~(inputs[528]);
    assign layer0_outputs[6041] = ~(inputs[108]);
    assign layer0_outputs[6042] = ~((inputs[964]) | (inputs[124]));
    assign layer0_outputs[6043] = ~(inputs[785]) | (inputs[855]);
    assign layer0_outputs[6044] = ~(inputs[347]);
    assign layer0_outputs[6045] = ~(inputs[797]) | (inputs[90]);
    assign layer0_outputs[6046] = (inputs[458]) & ~(inputs[773]);
    assign layer0_outputs[6047] = (inputs[555]) & ~(inputs[1007]);
    assign layer0_outputs[6048] = 1'b0;
    assign layer0_outputs[6049] = (inputs[660]) | (inputs[391]);
    assign layer0_outputs[6050] = (inputs[603]) | (inputs[706]);
    assign layer0_outputs[6051] = (inputs[497]) | (inputs[430]);
    assign layer0_outputs[6052] = ~(inputs[746]);
    assign layer0_outputs[6053] = ~(inputs[613]);
    assign layer0_outputs[6054] = (inputs[725]) ^ (inputs[566]);
    assign layer0_outputs[6055] = (inputs[215]) & ~(inputs[577]);
    assign layer0_outputs[6056] = ~((inputs[726]) | (inputs[271]));
    assign layer0_outputs[6057] = (inputs[437]) | (inputs[705]);
    assign layer0_outputs[6058] = inputs[685];
    assign layer0_outputs[6059] = inputs[166];
    assign layer0_outputs[6060] = ~(inputs[299]) | (inputs[143]);
    assign layer0_outputs[6061] = (inputs[299]) ^ (inputs[214]);
    assign layer0_outputs[6062] = (inputs[459]) & ~(inputs[422]);
    assign layer0_outputs[6063] = (inputs[85]) ^ (inputs[203]);
    assign layer0_outputs[6064] = ~((inputs[328]) ^ (inputs[737]));
    assign layer0_outputs[6065] = (inputs[618]) & ~(inputs[356]);
    assign layer0_outputs[6066] = ~((inputs[467]) & (inputs[778]));
    assign layer0_outputs[6067] = ~(inputs[847]) | (inputs[762]);
    assign layer0_outputs[6068] = ~(inputs[424]) | (inputs[215]);
    assign layer0_outputs[6069] = (inputs[191]) | (inputs[90]);
    assign layer0_outputs[6070] = ~(inputs[107]);
    assign layer0_outputs[6071] = ~((inputs[529]) | (inputs[51]));
    assign layer0_outputs[6072] = 1'b1;
    assign layer0_outputs[6073] = ~(inputs[374]) | (inputs[315]);
    assign layer0_outputs[6074] = ~((inputs[643]) | (inputs[15]));
    assign layer0_outputs[6075] = inputs[741];
    assign layer0_outputs[6076] = ~(inputs[128]);
    assign layer0_outputs[6077] = (inputs[216]) | (inputs[582]);
    assign layer0_outputs[6078] = (inputs[765]) ^ (inputs[539]);
    assign layer0_outputs[6079] = (inputs[558]) ^ (inputs[681]);
    assign layer0_outputs[6080] = (inputs[271]) ^ (inputs[665]);
    assign layer0_outputs[6081] = ~(inputs[20]) | (inputs[987]);
    assign layer0_outputs[6082] = ~(inputs[585]) | (inputs[663]);
    assign layer0_outputs[6083] = (inputs[100]) | (inputs[581]);
    assign layer0_outputs[6084] = (inputs[723]) & ~(inputs[123]);
    assign layer0_outputs[6085] = ~((inputs[393]) | (inputs[1016]));
    assign layer0_outputs[6086] = ~(inputs[602]) | (inputs[60]);
    assign layer0_outputs[6087] = ~((inputs[378]) | (inputs[320]));
    assign layer0_outputs[6088] = inputs[609];
    assign layer0_outputs[6089] = (inputs[428]) | (inputs[457]);
    assign layer0_outputs[6090] = inputs[237];
    assign layer0_outputs[6091] = ~((inputs[860]) ^ (inputs[599]));
    assign layer0_outputs[6092] = ~(inputs[718]) | (inputs[471]);
    assign layer0_outputs[6093] = ~(inputs[995]) | (inputs[955]);
    assign layer0_outputs[6094] = (inputs[686]) ^ (inputs[373]);
    assign layer0_outputs[6095] = (inputs[820]) & (inputs[848]);
    assign layer0_outputs[6096] = (inputs[159]) & (inputs[590]);
    assign layer0_outputs[6097] = ~((inputs[620]) | (inputs[558]));
    assign layer0_outputs[6098] = (inputs[410]) & ~(inputs[922]);
    assign layer0_outputs[6099] = ~((inputs[725]) | (inputs[711]));
    assign layer0_outputs[6100] = ~(inputs[995]) | (inputs[924]);
    assign layer0_outputs[6101] = (inputs[222]) & ~(inputs[30]);
    assign layer0_outputs[6102] = (inputs[824]) & ~(inputs[931]);
    assign layer0_outputs[6103] = ~((inputs[830]) | (inputs[945]));
    assign layer0_outputs[6104] = ~(inputs[694]);
    assign layer0_outputs[6105] = ~((inputs[272]) | (inputs[1006]));
    assign layer0_outputs[6106] = 1'b1;
    assign layer0_outputs[6107] = inputs[466];
    assign layer0_outputs[6108] = (inputs[512]) | (inputs[405]);
    assign layer0_outputs[6109] = (inputs[530]) & ~(inputs[1022]);
    assign layer0_outputs[6110] = (inputs[495]) & ~(inputs[173]);
    assign layer0_outputs[6111] = inputs[1019];
    assign layer0_outputs[6112] = (inputs[763]) | (inputs[791]);
    assign layer0_outputs[6113] = (inputs[737]) & ~(inputs[221]);
    assign layer0_outputs[6114] = inputs[6];
    assign layer0_outputs[6115] = ~(inputs[499]);
    assign layer0_outputs[6116] = 1'b0;
    assign layer0_outputs[6117] = inputs[138];
    assign layer0_outputs[6118] = 1'b0;
    assign layer0_outputs[6119] = (inputs[68]) ^ (inputs[246]);
    assign layer0_outputs[6120] = 1'b0;
    assign layer0_outputs[6121] = (inputs[471]) | (inputs[550]);
    assign layer0_outputs[6122] = (inputs[715]) ^ (inputs[250]);
    assign layer0_outputs[6123] = ~(inputs[944]) | (inputs[549]);
    assign layer0_outputs[6124] = ~((inputs[751]) | (inputs[799]));
    assign layer0_outputs[6125] = ~((inputs[7]) | (inputs[143]));
    assign layer0_outputs[6126] = (inputs[975]) ^ (inputs[476]);
    assign layer0_outputs[6127] = ~(inputs[414]) | (inputs[212]);
    assign layer0_outputs[6128] = ~((inputs[668]) & (inputs[60]));
    assign layer0_outputs[6129] = (inputs[657]) | (inputs[52]);
    assign layer0_outputs[6130] = ~(inputs[456]) | (inputs[66]);
    assign layer0_outputs[6131] = (inputs[748]) & ~(inputs[120]);
    assign layer0_outputs[6132] = (inputs[77]) ^ (inputs[741]);
    assign layer0_outputs[6133] = ~(inputs[425]);
    assign layer0_outputs[6134] = 1'b0;
    assign layer0_outputs[6135] = (inputs[454]) | (inputs[173]);
    assign layer0_outputs[6136] = inputs[301];
    assign layer0_outputs[6137] = ~(inputs[40]) | (inputs[933]);
    assign layer0_outputs[6138] = (inputs[79]) | (inputs[214]);
    assign layer0_outputs[6139] = (inputs[891]) | (inputs[851]);
    assign layer0_outputs[6140] = inputs[929];
    assign layer0_outputs[6141] = ~(inputs[636]) | (inputs[85]);
    assign layer0_outputs[6142] = (inputs[618]) & ~(inputs[128]);
    assign layer0_outputs[6143] = (inputs[469]) & ~(inputs[569]);
    assign layer0_outputs[6144] = (inputs[513]) ^ (inputs[896]);
    assign layer0_outputs[6145] = (inputs[975]) & ~(inputs[103]);
    assign layer0_outputs[6146] = (inputs[945]) & ~(inputs[722]);
    assign layer0_outputs[6147] = ~(inputs[905]);
    assign layer0_outputs[6148] = (inputs[896]) | (inputs[540]);
    assign layer0_outputs[6149] = ~(inputs[238]) | (inputs[548]);
    assign layer0_outputs[6150] = inputs[754];
    assign layer0_outputs[6151] = (inputs[149]) ^ (inputs[465]);
    assign layer0_outputs[6152] = (inputs[504]) ^ (inputs[525]);
    assign layer0_outputs[6153] = 1'b0;
    assign layer0_outputs[6154] = ~((inputs[948]) | (inputs[791]));
    assign layer0_outputs[6155] = ~((inputs[509]) & (inputs[350]));
    assign layer0_outputs[6156] = ~((inputs[388]) | (inputs[684]));
    assign layer0_outputs[6157] = (inputs[687]) | (inputs[440]);
    assign layer0_outputs[6158] = inputs[423];
    assign layer0_outputs[6159] = (inputs[215]) & ~(inputs[853]);
    assign layer0_outputs[6160] = ~(inputs[789]) | (inputs[260]);
    assign layer0_outputs[6161] = (inputs[895]) & ~(inputs[516]);
    assign layer0_outputs[6162] = (inputs[36]) & ~(inputs[613]);
    assign layer0_outputs[6163] = inputs[358];
    assign layer0_outputs[6164] = (inputs[672]) | (inputs[540]);
    assign layer0_outputs[6165] = 1'b0;
    assign layer0_outputs[6166] = ~((inputs[269]) | (inputs[908]));
    assign layer0_outputs[6167] = ~(inputs[295]);
    assign layer0_outputs[6168] = 1'b0;
    assign layer0_outputs[6169] = inputs[562];
    assign layer0_outputs[6170] = ~((inputs[655]) | (inputs[995]));
    assign layer0_outputs[6171] = ~(inputs[644]) | (inputs[154]);
    assign layer0_outputs[6172] = inputs[744];
    assign layer0_outputs[6173] = ~(inputs[490]) | (inputs[706]);
    assign layer0_outputs[6174] = (inputs[587]) | (inputs[161]);
    assign layer0_outputs[6175] = ~(inputs[974]);
    assign layer0_outputs[6176] = ~(inputs[619]);
    assign layer0_outputs[6177] = (inputs[983]) & ~(inputs[63]);
    assign layer0_outputs[6178] = 1'b1;
    assign layer0_outputs[6179] = ~(inputs[533]);
    assign layer0_outputs[6180] = (inputs[851]) & ~(inputs[922]);
    assign layer0_outputs[6181] = ~(inputs[491]);
    assign layer0_outputs[6182] = ~(inputs[591]) | (inputs[413]);
    assign layer0_outputs[6183] = (inputs[266]) ^ (inputs[397]);
    assign layer0_outputs[6184] = (inputs[663]) & (inputs[418]);
    assign layer0_outputs[6185] = ~((inputs[163]) | (inputs[333]));
    assign layer0_outputs[6186] = inputs[459];
    assign layer0_outputs[6187] = 1'b0;
    assign layer0_outputs[6188] = ~((inputs[497]) | (inputs[313]));
    assign layer0_outputs[6189] = (inputs[670]) | (inputs[727]);
    assign layer0_outputs[6190] = inputs[461];
    assign layer0_outputs[6191] = inputs[884];
    assign layer0_outputs[6192] = 1'b1;
    assign layer0_outputs[6193] = ~(inputs[377]) | (inputs[959]);
    assign layer0_outputs[6194] = (inputs[113]) & ~(inputs[642]);
    assign layer0_outputs[6195] = inputs[266];
    assign layer0_outputs[6196] = (inputs[407]) ^ (inputs[259]);
    assign layer0_outputs[6197] = 1'b1;
    assign layer0_outputs[6198] = (inputs[203]) & ~(inputs[46]);
    assign layer0_outputs[6199] = (inputs[266]) ^ (inputs[125]);
    assign layer0_outputs[6200] = ~((inputs[38]) ^ (inputs[63]));
    assign layer0_outputs[6201] = (inputs[385]) | (inputs[402]);
    assign layer0_outputs[6202] = inputs[186];
    assign layer0_outputs[6203] = ~((inputs[1010]) ^ (inputs[777]));
    assign layer0_outputs[6204] = ~(inputs[855]);
    assign layer0_outputs[6205] = ~(inputs[578]) | (inputs[271]);
    assign layer0_outputs[6206] = (inputs[691]) & ~(inputs[518]);
    assign layer0_outputs[6207] = inputs[299];
    assign layer0_outputs[6208] = (inputs[861]) | (inputs[83]);
    assign layer0_outputs[6209] = ~((inputs[702]) & (inputs[64]));
    assign layer0_outputs[6210] = 1'b1;
    assign layer0_outputs[6211] = inputs[574];
    assign layer0_outputs[6212] = (inputs[977]) & ~(inputs[401]);
    assign layer0_outputs[6213] = (inputs[858]) ^ (inputs[537]);
    assign layer0_outputs[6214] = ~((inputs[955]) | (inputs[329]));
    assign layer0_outputs[6215] = ~(inputs[560]);
    assign layer0_outputs[6216] = (inputs[327]) | (inputs[112]);
    assign layer0_outputs[6217] = ~((inputs[702]) ^ (inputs[1009]));
    assign layer0_outputs[6218] = ~(inputs[297]);
    assign layer0_outputs[6219] = ~(inputs[580]);
    assign layer0_outputs[6220] = inputs[315];
    assign layer0_outputs[6221] = (inputs[379]) & ~(inputs[493]);
    assign layer0_outputs[6222] = (inputs[877]) | (inputs[317]);
    assign layer0_outputs[6223] = (inputs[1011]) | (inputs[179]);
    assign layer0_outputs[6224] = inputs[894];
    assign layer0_outputs[6225] = inputs[775];
    assign layer0_outputs[6226] = (inputs[757]) | (inputs[681]);
    assign layer0_outputs[6227] = ~((inputs[381]) | (inputs[426]));
    assign layer0_outputs[6228] = 1'b1;
    assign layer0_outputs[6229] = (inputs[985]) | (inputs[689]);
    assign layer0_outputs[6230] = ~(inputs[127]);
    assign layer0_outputs[6231] = (inputs[446]) & (inputs[147]);
    assign layer0_outputs[6232] = ~(inputs[594]) | (inputs[387]);
    assign layer0_outputs[6233] = (inputs[778]) | (inputs[812]);
    assign layer0_outputs[6234] = inputs[243];
    assign layer0_outputs[6235] = (inputs[82]) | (inputs[171]);
    assign layer0_outputs[6236] = inputs[433];
    assign layer0_outputs[6237] = (inputs[461]) & ~(inputs[945]);
    assign layer0_outputs[6238] = ~(inputs[581]);
    assign layer0_outputs[6239] = 1'b1;
    assign layer0_outputs[6240] = ~(inputs[445]);
    assign layer0_outputs[6241] = (inputs[203]) & ~(inputs[948]);
    assign layer0_outputs[6242] = (inputs[824]) | (inputs[17]);
    assign layer0_outputs[6243] = inputs[836];
    assign layer0_outputs[6244] = inputs[499];
    assign layer0_outputs[6245] = inputs[372];
    assign layer0_outputs[6246] = inputs[428];
    assign layer0_outputs[6247] = (inputs[100]) | (inputs[587]);
    assign layer0_outputs[6248] = (inputs[404]) & ~(inputs[788]);
    assign layer0_outputs[6249] = (inputs[980]) ^ (inputs[984]);
    assign layer0_outputs[6250] = ~(inputs[887]);
    assign layer0_outputs[6251] = ~(inputs[428]) | (inputs[474]);
    assign layer0_outputs[6252] = (inputs[241]) | (inputs[249]);
    assign layer0_outputs[6253] = (inputs[324]) | (inputs[99]);
    assign layer0_outputs[6254] = ~((inputs[466]) | (inputs[500]));
    assign layer0_outputs[6255] = ~(inputs[358]) | (inputs[1001]);
    assign layer0_outputs[6256] = ~((inputs[378]) | (inputs[493]));
    assign layer0_outputs[6257] = ~(inputs[460]);
    assign layer0_outputs[6258] = (inputs[697]) | (inputs[911]);
    assign layer0_outputs[6259] = 1'b1;
    assign layer0_outputs[6260] = (inputs[166]) | (inputs[669]);
    assign layer0_outputs[6261] = (inputs[617]) | (inputs[406]);
    assign layer0_outputs[6262] = ~((inputs[559]) | (inputs[713]));
    assign layer0_outputs[6263] = ~(inputs[753]) | (inputs[21]);
    assign layer0_outputs[6264] = ~((inputs[1000]) & (inputs[82]));
    assign layer0_outputs[6265] = (inputs[986]) ^ (inputs[206]);
    assign layer0_outputs[6266] = (inputs[305]) & ~(inputs[90]);
    assign layer0_outputs[6267] = 1'b1;
    assign layer0_outputs[6268] = (inputs[1012]) | (inputs[300]);
    assign layer0_outputs[6269] = ~(inputs[81]) | (inputs[542]);
    assign layer0_outputs[6270] = (inputs[441]) & ~(inputs[802]);
    assign layer0_outputs[6271] = (inputs[120]) & ~(inputs[1004]);
    assign layer0_outputs[6272] = inputs[497];
    assign layer0_outputs[6273] = 1'b0;
    assign layer0_outputs[6274] = ~((inputs[422]) | (inputs[53]));
    assign layer0_outputs[6275] = inputs[997];
    assign layer0_outputs[6276] = (inputs[383]) & (inputs[961]);
    assign layer0_outputs[6277] = ~(inputs[245]) | (inputs[448]);
    assign layer0_outputs[6278] = ~((inputs[943]) | (inputs[20]));
    assign layer0_outputs[6279] = (inputs[407]) | (inputs[165]);
    assign layer0_outputs[6280] = ~((inputs[889]) | (inputs[1004]));
    assign layer0_outputs[6281] = ~((inputs[964]) ^ (inputs[773]));
    assign layer0_outputs[6282] = (inputs[590]) | (inputs[230]);
    assign layer0_outputs[6283] = (inputs[798]) | (inputs[724]);
    assign layer0_outputs[6284] = (inputs[639]) & (inputs[446]);
    assign layer0_outputs[6285] = ~(inputs[409]);
    assign layer0_outputs[6286] = ~(inputs[808]) | (inputs[868]);
    assign layer0_outputs[6287] = (inputs[496]) & ~(inputs[739]);
    assign layer0_outputs[6288] = ~((inputs[933]) ^ (inputs[234]));
    assign layer0_outputs[6289] = ~((inputs[0]) ^ (inputs[26]));
    assign layer0_outputs[6290] = (inputs[961]) & ~(inputs[20]);
    assign layer0_outputs[6291] = ~((inputs[342]) | (inputs[810]));
    assign layer0_outputs[6292] = (inputs[780]) & ~(inputs[974]);
    assign layer0_outputs[6293] = inputs[638];
    assign layer0_outputs[6294] = ~((inputs[253]) ^ (inputs[462]));
    assign layer0_outputs[6295] = ~((inputs[818]) | (inputs[424]));
    assign layer0_outputs[6296] = inputs[311];
    assign layer0_outputs[6297] = ~((inputs[134]) & (inputs[734]));
    assign layer0_outputs[6298] = 1'b0;
    assign layer0_outputs[6299] = ~((inputs[780]) ^ (inputs[830]));
    assign layer0_outputs[6300] = (inputs[483]) | (inputs[467]);
    assign layer0_outputs[6301] = ~(inputs[529]) | (inputs[100]);
    assign layer0_outputs[6302] = (inputs[648]) & ~(inputs[926]);
    assign layer0_outputs[6303] = ~((inputs[353]) | (inputs[525]));
    assign layer0_outputs[6304] = ~(inputs[897]);
    assign layer0_outputs[6305] = ~(inputs[301]);
    assign layer0_outputs[6306] = ~(inputs[201]);
    assign layer0_outputs[6307] = ~(inputs[337]);
    assign layer0_outputs[6308] = ~(inputs[533]) | (inputs[871]);
    assign layer0_outputs[6309] = ~((inputs[540]) | (inputs[757]));
    assign layer0_outputs[6310] = (inputs[694]) & (inputs[720]);
    assign layer0_outputs[6311] = (inputs[857]) ^ (inputs[651]);
    assign layer0_outputs[6312] = ~(inputs[46]) | (inputs[13]);
    assign layer0_outputs[6313] = ~(inputs[815]);
    assign layer0_outputs[6314] = ~((inputs[382]) & (inputs[292]));
    assign layer0_outputs[6315] = inputs[639];
    assign layer0_outputs[6316] = ~((inputs[153]) ^ (inputs[219]));
    assign layer0_outputs[6317] = ~((inputs[960]) | (inputs[962]));
    assign layer0_outputs[6318] = ~(inputs[717]);
    assign layer0_outputs[6319] = (inputs[335]) | (inputs[923]);
    assign layer0_outputs[6320] = inputs[422];
    assign layer0_outputs[6321] = (inputs[489]) | (inputs[255]);
    assign layer0_outputs[6322] = ~((inputs[273]) ^ (inputs[975]));
    assign layer0_outputs[6323] = ~((inputs[361]) | (inputs[313]));
    assign layer0_outputs[6324] = (inputs[803]) ^ (inputs[506]);
    assign layer0_outputs[6325] = inputs[539];
    assign layer0_outputs[6326] = inputs[280];
    assign layer0_outputs[6327] = ~(inputs[106]);
    assign layer0_outputs[6328] = ~(inputs[338]) | (inputs[378]);
    assign layer0_outputs[6329] = (inputs[241]) & ~(inputs[452]);
    assign layer0_outputs[6330] = (inputs[596]) & ~(inputs[41]);
    assign layer0_outputs[6331] = ~((inputs[356]) | (inputs[43]));
    assign layer0_outputs[6332] = ~(inputs[146]);
    assign layer0_outputs[6333] = (inputs[539]) & ~(inputs[257]);
    assign layer0_outputs[6334] = 1'b1;
    assign layer0_outputs[6335] = ~(inputs[740]) | (inputs[39]);
    assign layer0_outputs[6336] = ~((inputs[420]) ^ (inputs[912]));
    assign layer0_outputs[6337] = ~(inputs[468]);
    assign layer0_outputs[6338] = (inputs[274]) & (inputs[193]);
    assign layer0_outputs[6339] = ~(inputs[505]);
    assign layer0_outputs[6340] = ~(inputs[519]);
    assign layer0_outputs[6341] = (inputs[476]) | (inputs[563]);
    assign layer0_outputs[6342] = 1'b0;
    assign layer0_outputs[6343] = (inputs[547]) ^ (inputs[578]);
    assign layer0_outputs[6344] = 1'b1;
    assign layer0_outputs[6345] = ~(inputs[151]);
    assign layer0_outputs[6346] = ~((inputs[968]) | (inputs[345]));
    assign layer0_outputs[6347] = ~((inputs[434]) & (inputs[1014]));
    assign layer0_outputs[6348] = ~(inputs[607]) | (inputs[762]);
    assign layer0_outputs[6349] = ~(inputs[264]);
    assign layer0_outputs[6350] = (inputs[580]) | (inputs[884]);
    assign layer0_outputs[6351] = inputs[786];
    assign layer0_outputs[6352] = ~(inputs[154]) | (inputs[9]);
    assign layer0_outputs[6353] = ~((inputs[917]) & (inputs[348]));
    assign layer0_outputs[6354] = ~((inputs[13]) ^ (inputs[251]));
    assign layer0_outputs[6355] = ~((inputs[724]) | (inputs[201]));
    assign layer0_outputs[6356] = ~((inputs[509]) | (inputs[396]));
    assign layer0_outputs[6357] = 1'b1;
    assign layer0_outputs[6358] = ~((inputs[207]) | (inputs[156]));
    assign layer0_outputs[6359] = 1'b1;
    assign layer0_outputs[6360] = inputs[661];
    assign layer0_outputs[6361] = (inputs[43]) ^ (inputs[937]);
    assign layer0_outputs[6362] = (inputs[701]) | (inputs[389]);
    assign layer0_outputs[6363] = ~((inputs[774]) | (inputs[695]));
    assign layer0_outputs[6364] = ~(inputs[800]);
    assign layer0_outputs[6365] = ~(inputs[522]) | (inputs[343]);
    assign layer0_outputs[6366] = 1'b0;
    assign layer0_outputs[6367] = (inputs[195]) ^ (inputs[442]);
    assign layer0_outputs[6368] = ~((inputs[667]) ^ (inputs[886]));
    assign layer0_outputs[6369] = ~((inputs[767]) | (inputs[449]));
    assign layer0_outputs[6370] = ~(inputs[849]);
    assign layer0_outputs[6371] = inputs[812];
    assign layer0_outputs[6372] = (inputs[624]) | (inputs[590]);
    assign layer0_outputs[6373] = (inputs[958]) ^ (inputs[816]);
    assign layer0_outputs[6374] = 1'b0;
    assign layer0_outputs[6375] = ~(inputs[986]);
    assign layer0_outputs[6376] = (inputs[87]) & ~(inputs[610]);
    assign layer0_outputs[6377] = ~((inputs[89]) ^ (inputs[157]));
    assign layer0_outputs[6378] = ~(inputs[347]) | (inputs[638]);
    assign layer0_outputs[6379] = ~((inputs[678]) ^ (inputs[604]));
    assign layer0_outputs[6380] = ~(inputs[56]);
    assign layer0_outputs[6381] = inputs[492];
    assign layer0_outputs[6382] = (inputs[583]) & ~(inputs[939]);
    assign layer0_outputs[6383] = ~(inputs[913]);
    assign layer0_outputs[6384] = ~(inputs[727]);
    assign layer0_outputs[6385] = (inputs[220]) & ~(inputs[387]);
    assign layer0_outputs[6386] = (inputs[507]) & ~(inputs[942]);
    assign layer0_outputs[6387] = (inputs[884]) | (inputs[136]);
    assign layer0_outputs[6388] = ~((inputs[307]) | (inputs[680]));
    assign layer0_outputs[6389] = (inputs[1014]) & ~(inputs[635]);
    assign layer0_outputs[6390] = inputs[15];
    assign layer0_outputs[6391] = ~((inputs[682]) | (inputs[52]));
    assign layer0_outputs[6392] = ~((inputs[261]) | (inputs[294]));
    assign layer0_outputs[6393] = (inputs[597]) & ~(inputs[835]);
    assign layer0_outputs[6394] = inputs[585];
    assign layer0_outputs[6395] = ~(inputs[264]) | (inputs[713]);
    assign layer0_outputs[6396] = (inputs[650]) & ~(inputs[912]);
    assign layer0_outputs[6397] = (inputs[806]) ^ (inputs[453]);
    assign layer0_outputs[6398] = (inputs[462]) & ~(inputs[24]);
    assign layer0_outputs[6399] = ~(inputs[695]);
    assign layer0_outputs[6400] = ~((inputs[772]) & (inputs[1004]));
    assign layer0_outputs[6401] = (inputs[681]) ^ (inputs[789]);
    assign layer0_outputs[6402] = 1'b1;
    assign layer0_outputs[6403] = inputs[879];
    assign layer0_outputs[6404] = 1'b1;
    assign layer0_outputs[6405] = (inputs[117]) ^ (inputs[402]);
    assign layer0_outputs[6406] = (inputs[718]) & ~(inputs[728]);
    assign layer0_outputs[6407] = (inputs[196]) ^ (inputs[552]);
    assign layer0_outputs[6408] = ~(inputs[242]);
    assign layer0_outputs[6409] = inputs[885];
    assign layer0_outputs[6410] = (inputs[561]) | (inputs[186]);
    assign layer0_outputs[6411] = ~(inputs[335]) | (inputs[100]);
    assign layer0_outputs[6412] = (inputs[684]) ^ (inputs[445]);
    assign layer0_outputs[6413] = (inputs[434]) | (inputs[198]);
    assign layer0_outputs[6414] = 1'b1;
    assign layer0_outputs[6415] = (inputs[109]) & (inputs[950]);
    assign layer0_outputs[6416] = (inputs[49]) ^ (inputs[119]);
    assign layer0_outputs[6417] = ~(inputs[186]);
    assign layer0_outputs[6418] = (inputs[568]) & ~(inputs[285]);
    assign layer0_outputs[6419] = inputs[124];
    assign layer0_outputs[6420] = ~(inputs[844]);
    assign layer0_outputs[6421] = (inputs[824]) ^ (inputs[1001]);
    assign layer0_outputs[6422] = ~(inputs[264]);
    assign layer0_outputs[6423] = ~(inputs[84]);
    assign layer0_outputs[6424] = (inputs[851]) | (inputs[433]);
    assign layer0_outputs[6425] = (inputs[29]) | (inputs[567]);
    assign layer0_outputs[6426] = ~((inputs[114]) ^ (inputs[715]));
    assign layer0_outputs[6427] = ~((inputs[61]) ^ (inputs[274]));
    assign layer0_outputs[6428] = ~(inputs[364]) | (inputs[279]);
    assign layer0_outputs[6429] = (inputs[479]) & ~(inputs[181]);
    assign layer0_outputs[6430] = ~(inputs[71]) | (inputs[1012]);
    assign layer0_outputs[6431] = ~((inputs[28]) | (inputs[150]));
    assign layer0_outputs[6432] = (inputs[650]) | (inputs[142]);
    assign layer0_outputs[6433] = ~((inputs[184]) ^ (inputs[746]));
    assign layer0_outputs[6434] = (inputs[754]) | (inputs[1002]);
    assign layer0_outputs[6435] = (inputs[913]) & ~(inputs[55]);
    assign layer0_outputs[6436] = (inputs[265]) | (inputs[201]);
    assign layer0_outputs[6437] = ~((inputs[280]) ^ (inputs[411]));
    assign layer0_outputs[6438] = (inputs[686]) | (inputs[704]);
    assign layer0_outputs[6439] = ~(inputs[726]);
    assign layer0_outputs[6440] = ~(inputs[946]);
    assign layer0_outputs[6441] = (inputs[431]) & ~(inputs[444]);
    assign layer0_outputs[6442] = (inputs[34]) ^ (inputs[487]);
    assign layer0_outputs[6443] = ~((inputs[92]) | (inputs[95]));
    assign layer0_outputs[6444] = (inputs[640]) | (inputs[877]);
    assign layer0_outputs[6445] = ~(inputs[1022]);
    assign layer0_outputs[6446] = (inputs[830]) & ~(inputs[540]);
    assign layer0_outputs[6447] = ~((inputs[152]) | (inputs[41]));
    assign layer0_outputs[6448] = ~((inputs[977]) | (inputs[979]));
    assign layer0_outputs[6449] = inputs[651];
    assign layer0_outputs[6450] = ~(inputs[241]);
    assign layer0_outputs[6451] = ~((inputs[129]) & (inputs[257]));
    assign layer0_outputs[6452] = inputs[527];
    assign layer0_outputs[6453] = (inputs[1014]) & ~(inputs[801]);
    assign layer0_outputs[6454] = inputs[331];
    assign layer0_outputs[6455] = (inputs[588]) | (inputs[688]);
    assign layer0_outputs[6456] = (inputs[409]) ^ (inputs[323]);
    assign layer0_outputs[6457] = (inputs[144]) & ~(inputs[930]);
    assign layer0_outputs[6458] = (inputs[716]) | (inputs[147]);
    assign layer0_outputs[6459] = ~(inputs[853]) | (inputs[42]);
    assign layer0_outputs[6460] = (inputs[899]) | (inputs[444]);
    assign layer0_outputs[6461] = ~(inputs[5]) | (inputs[145]);
    assign layer0_outputs[6462] = inputs[777];
    assign layer0_outputs[6463] = ~(inputs[624]);
    assign layer0_outputs[6464] = (inputs[328]) & ~(inputs[1008]);
    assign layer0_outputs[6465] = ~(inputs[704]) | (inputs[1006]);
    assign layer0_outputs[6466] = ~(inputs[194]);
    assign layer0_outputs[6467] = (inputs[885]) & ~(inputs[165]);
    assign layer0_outputs[6468] = (inputs[109]) & ~(inputs[1013]);
    assign layer0_outputs[6469] = ~((inputs[865]) & (inputs[362]));
    assign layer0_outputs[6470] = inputs[820];
    assign layer0_outputs[6471] = ~((inputs[791]) | (inputs[127]));
    assign layer0_outputs[6472] = (inputs[1003]) & ~(inputs[797]);
    assign layer0_outputs[6473] = ~((inputs[705]) ^ (inputs[791]));
    assign layer0_outputs[6474] = ~(inputs[6]);
    assign layer0_outputs[6475] = ~(inputs[423]) | (inputs[320]);
    assign layer0_outputs[6476] = (inputs[185]) & ~(inputs[738]);
    assign layer0_outputs[6477] = ~(inputs[909]);
    assign layer0_outputs[6478] = ~(inputs[871]) | (inputs[194]);
    assign layer0_outputs[6479] = (inputs[981]) & ~(inputs[101]);
    assign layer0_outputs[6480] = (inputs[276]) ^ (inputs[724]);
    assign layer0_outputs[6481] = ~((inputs[991]) ^ (inputs[842]));
    assign layer0_outputs[6482] = ~((inputs[21]) ^ (inputs[935]));
    assign layer0_outputs[6483] = ~(inputs[807]);
    assign layer0_outputs[6484] = inputs[325];
    assign layer0_outputs[6485] = (inputs[171]) & ~(inputs[408]);
    assign layer0_outputs[6486] = ~(inputs[752]);
    assign layer0_outputs[6487] = (inputs[505]) & ~(inputs[957]);
    assign layer0_outputs[6488] = 1'b1;
    assign layer0_outputs[6489] = ~(inputs[676]);
    assign layer0_outputs[6490] = ~((inputs[338]) ^ (inputs[213]));
    assign layer0_outputs[6491] = ~(inputs[156]);
    assign layer0_outputs[6492] = ~(inputs[527]);
    assign layer0_outputs[6493] = ~((inputs[649]) | (inputs[438]));
    assign layer0_outputs[6494] = inputs[256];
    assign layer0_outputs[6495] = inputs[808];
    assign layer0_outputs[6496] = ~(inputs[77]);
    assign layer0_outputs[6497] = ~((inputs[978]) ^ (inputs[815]));
    assign layer0_outputs[6498] = ~((inputs[468]) | (inputs[675]));
    assign layer0_outputs[6499] = 1'b0;
    assign layer0_outputs[6500] = inputs[999];
    assign layer0_outputs[6501] = ~(inputs[497]);
    assign layer0_outputs[6502] = ~((inputs[247]) | (inputs[511]));
    assign layer0_outputs[6503] = ~(inputs[979]) | (inputs[955]);
    assign layer0_outputs[6504] = ~(inputs[902]);
    assign layer0_outputs[6505] = ~(inputs[681]);
    assign layer0_outputs[6506] = (inputs[926]) & ~(inputs[971]);
    assign layer0_outputs[6507] = ~(inputs[865]) | (inputs[55]);
    assign layer0_outputs[6508] = ~((inputs[141]) | (inputs[49]));
    assign layer0_outputs[6509] = ~((inputs[404]) | (inputs[659]));
    assign layer0_outputs[6510] = 1'b1;
    assign layer0_outputs[6511] = ~(inputs[198]) | (inputs[840]);
    assign layer0_outputs[6512] = (inputs[96]) | (inputs[943]);
    assign layer0_outputs[6513] = ~((inputs[616]) | (inputs[545]));
    assign layer0_outputs[6514] = ~(inputs[99]) | (inputs[635]);
    assign layer0_outputs[6515] = ~(inputs[36]) | (inputs[285]);
    assign layer0_outputs[6516] = inputs[870];
    assign layer0_outputs[6517] = ~(inputs[677]) | (inputs[116]);
    assign layer0_outputs[6518] = (inputs[437]) & ~(inputs[941]);
    assign layer0_outputs[6519] = ~((inputs[180]) ^ (inputs[795]));
    assign layer0_outputs[6520] = ~(inputs[210]) | (inputs[262]);
    assign layer0_outputs[6521] = (inputs[914]) & ~(inputs[665]);
    assign layer0_outputs[6522] = inputs[47];
    assign layer0_outputs[6523] = (inputs[929]) | (inputs[221]);
    assign layer0_outputs[6524] = ~((inputs[174]) | (inputs[844]));
    assign layer0_outputs[6525] = (inputs[370]) & ~(inputs[354]);
    assign layer0_outputs[6526] = (inputs[521]) & ~(inputs[855]);
    assign layer0_outputs[6527] = ~(inputs[285]) | (inputs[290]);
    assign layer0_outputs[6528] = ~((inputs[64]) ^ (inputs[409]));
    assign layer0_outputs[6529] = ~(inputs[458]) | (inputs[686]);
    assign layer0_outputs[6530] = (inputs[96]) | (inputs[558]);
    assign layer0_outputs[6531] = ~(inputs[604]) | (inputs[350]);
    assign layer0_outputs[6532] = ~(inputs[246]);
    assign layer0_outputs[6533] = (inputs[912]) | (inputs[485]);
    assign layer0_outputs[6534] = ~((inputs[112]) | (inputs[248]));
    assign layer0_outputs[6535] = ~(inputs[915]);
    assign layer0_outputs[6536] = ~((inputs[537]) & (inputs[952]));
    assign layer0_outputs[6537] = (inputs[374]) & ~(inputs[324]);
    assign layer0_outputs[6538] = ~(inputs[251]);
    assign layer0_outputs[6539] = inputs[454];
    assign layer0_outputs[6540] = (inputs[775]) ^ (inputs[400]);
    assign layer0_outputs[6541] = inputs[299];
    assign layer0_outputs[6542] = ~(inputs[557]) | (inputs[905]);
    assign layer0_outputs[6543] = ~((inputs[1000]) & (inputs[630]));
    assign layer0_outputs[6544] = ~((inputs[378]) ^ (inputs[894]));
    assign layer0_outputs[6545] = ~((inputs[207]) | (inputs[288]));
    assign layer0_outputs[6546] = ~((inputs[534]) | (inputs[424]));
    assign layer0_outputs[6547] = 1'b1;
    assign layer0_outputs[6548] = inputs[711];
    assign layer0_outputs[6549] = ~((inputs[482]) & (inputs[136]));
    assign layer0_outputs[6550] = (inputs[774]) | (inputs[440]);
    assign layer0_outputs[6551] = inputs[960];
    assign layer0_outputs[6552] = ~((inputs[688]) ^ (inputs[989]));
    assign layer0_outputs[6553] = (inputs[368]) | (inputs[700]);
    assign layer0_outputs[6554] = ~((inputs[244]) ^ (inputs[483]));
    assign layer0_outputs[6555] = inputs[618];
    assign layer0_outputs[6556] = ~(inputs[155]);
    assign layer0_outputs[6557] = ~((inputs[711]) & (inputs[173]));
    assign layer0_outputs[6558] = ~(inputs[341]);
    assign layer0_outputs[6559] = (inputs[702]) | (inputs[115]);
    assign layer0_outputs[6560] = (inputs[334]) & ~(inputs[16]);
    assign layer0_outputs[6561] = (inputs[144]) ^ (inputs[733]);
    assign layer0_outputs[6562] = ~((inputs[631]) | (inputs[173]));
    assign layer0_outputs[6563] = inputs[224];
    assign layer0_outputs[6564] = ~(inputs[926]) | (inputs[169]);
    assign layer0_outputs[6565] = ~((inputs[1006]) | (inputs[129]));
    assign layer0_outputs[6566] = ~((inputs[435]) | (inputs[340]));
    assign layer0_outputs[6567] = inputs[525];
    assign layer0_outputs[6568] = (inputs[247]) & ~(inputs[507]);
    assign layer0_outputs[6569] = ~(inputs[139]) | (inputs[860]);
    assign layer0_outputs[6570] = inputs[485];
    assign layer0_outputs[6571] = ~(inputs[777]);
    assign layer0_outputs[6572] = (inputs[480]) ^ (inputs[930]);
    assign layer0_outputs[6573] = inputs[522];
    assign layer0_outputs[6574] = ~(inputs[239]) | (inputs[321]);
    assign layer0_outputs[6575] = 1'b0;
    assign layer0_outputs[6576] = (inputs[496]) & ~(inputs[905]);
    assign layer0_outputs[6577] = (inputs[690]) & ~(inputs[34]);
    assign layer0_outputs[6578] = ~(inputs[13]) | (inputs[60]);
    assign layer0_outputs[6579] = ~(inputs[994]) | (inputs[971]);
    assign layer0_outputs[6580] = (inputs[358]) ^ (inputs[422]);
    assign layer0_outputs[6581] = ~(inputs[280]);
    assign layer0_outputs[6582] = inputs[831];
    assign layer0_outputs[6583] = (inputs[350]) & ~(inputs[702]);
    assign layer0_outputs[6584] = ~(inputs[523]);
    assign layer0_outputs[6585] = ~((inputs[840]) & (inputs[982]));
    assign layer0_outputs[6586] = ~((inputs[862]) ^ (inputs[925]));
    assign layer0_outputs[6587] = (inputs[103]) & ~(inputs[734]);
    assign layer0_outputs[6588] = ~(inputs[58]) | (inputs[376]);
    assign layer0_outputs[6589] = ~((inputs[870]) | (inputs[719]));
    assign layer0_outputs[6590] = ~(inputs[89]);
    assign layer0_outputs[6591] = ~((inputs[391]) ^ (inputs[201]));
    assign layer0_outputs[6592] = ~(inputs[713]) | (inputs[826]);
    assign layer0_outputs[6593] = ~((inputs[964]) | (inputs[240]));
    assign layer0_outputs[6594] = ~(inputs[282]) | (inputs[1022]);
    assign layer0_outputs[6595] = ~((inputs[868]) | (inputs[802]));
    assign layer0_outputs[6596] = ~((inputs[568]) | (inputs[572]));
    assign layer0_outputs[6597] = (inputs[942]) ^ (inputs[821]);
    assign layer0_outputs[6598] = (inputs[934]) & ~(inputs[92]);
    assign layer0_outputs[6599] = ~(inputs[407]) | (inputs[420]);
    assign layer0_outputs[6600] = (inputs[882]) ^ (inputs[260]);
    assign layer0_outputs[6601] = (inputs[274]) & ~(inputs[287]);
    assign layer0_outputs[6602] = 1'b0;
    assign layer0_outputs[6603] = ~(inputs[560]);
    assign layer0_outputs[6604] = 1'b0;
    assign layer0_outputs[6605] = ~(inputs[573]);
    assign layer0_outputs[6606] = (inputs[847]) ^ (inputs[382]);
    assign layer0_outputs[6607] = (inputs[172]) & ~(inputs[937]);
    assign layer0_outputs[6608] = ~((inputs[922]) & (inputs[580]));
    assign layer0_outputs[6609] = inputs[279];
    assign layer0_outputs[6610] = (inputs[437]) & ~(inputs[778]);
    assign layer0_outputs[6611] = (inputs[1010]) | (inputs[880]);
    assign layer0_outputs[6612] = inputs[494];
    assign layer0_outputs[6613] = ~(inputs[812]);
    assign layer0_outputs[6614] = (inputs[145]) | (inputs[491]);
    assign layer0_outputs[6615] = 1'b0;
    assign layer0_outputs[6616] = ~(inputs[364]);
    assign layer0_outputs[6617] = inputs[239];
    assign layer0_outputs[6618] = (inputs[714]) & ~(inputs[925]);
    assign layer0_outputs[6619] = (inputs[98]) ^ (inputs[673]);
    assign layer0_outputs[6620] = ~(inputs[780]);
    assign layer0_outputs[6621] = 1'b0;
    assign layer0_outputs[6622] = inputs[439];
    assign layer0_outputs[6623] = inputs[471];
    assign layer0_outputs[6624] = ~((inputs[288]) | (inputs[247]));
    assign layer0_outputs[6625] = inputs[462];
    assign layer0_outputs[6626] = inputs[452];
    assign layer0_outputs[6627] = ~((inputs[605]) & (inputs[29]));
    assign layer0_outputs[6628] = 1'b1;
    assign layer0_outputs[6629] = ~(inputs[740]) | (inputs[485]);
    assign layer0_outputs[6630] = ~(inputs[501]);
    assign layer0_outputs[6631] = ~(inputs[692]) | (inputs[324]);
    assign layer0_outputs[6632] = (inputs[327]) ^ (inputs[710]);
    assign layer0_outputs[6633] = ~((inputs[565]) | (inputs[600]));
    assign layer0_outputs[6634] = ~((inputs[513]) ^ (inputs[432]));
    assign layer0_outputs[6635] = ~((inputs[152]) ^ (inputs[547]));
    assign layer0_outputs[6636] = (inputs[902]) & ~(inputs[222]);
    assign layer0_outputs[6637] = ~(inputs[459]) | (inputs[400]);
    assign layer0_outputs[6638] = (inputs[618]) & ~(inputs[947]);
    assign layer0_outputs[6639] = (inputs[69]) & ~(inputs[16]);
    assign layer0_outputs[6640] = ~((inputs[803]) | (inputs[464]));
    assign layer0_outputs[6641] = (inputs[257]) | (inputs[265]);
    assign layer0_outputs[6642] = inputs[263];
    assign layer0_outputs[6643] = ~((inputs[502]) ^ (inputs[217]));
    assign layer0_outputs[6644] = ~((inputs[321]) ^ (inputs[230]));
    assign layer0_outputs[6645] = (inputs[1000]) & (inputs[12]);
    assign layer0_outputs[6646] = (inputs[232]) & ~(inputs[86]);
    assign layer0_outputs[6647] = ~((inputs[189]) ^ (inputs[427]));
    assign layer0_outputs[6648] = 1'b0;
    assign layer0_outputs[6649] = ~(inputs[339]);
    assign layer0_outputs[6650] = (inputs[144]) | (inputs[446]);
    assign layer0_outputs[6651] = ~(inputs[403]) | (inputs[55]);
    assign layer0_outputs[6652] = ~((inputs[441]) & (inputs[95]));
    assign layer0_outputs[6653] = ~((inputs[375]) | (inputs[981]));
    assign layer0_outputs[6654] = ~(inputs[466]) | (inputs[279]);
    assign layer0_outputs[6655] = ~((inputs[204]) | (inputs[882]));
    assign layer0_outputs[6656] = (inputs[603]) & ~(inputs[132]);
    assign layer0_outputs[6657] = (inputs[171]) & ~(inputs[12]);
    assign layer0_outputs[6658] = inputs[42];
    assign layer0_outputs[6659] = (inputs[384]) & (inputs[926]);
    assign layer0_outputs[6660] = ~(inputs[896]);
    assign layer0_outputs[6661] = (inputs[535]) ^ (inputs[875]);
    assign layer0_outputs[6662] = ~(inputs[22]);
    assign layer0_outputs[6663] = (inputs[52]) | (inputs[853]);
    assign layer0_outputs[6664] = ~((inputs[378]) | (inputs[662]));
    assign layer0_outputs[6665] = ~((inputs[32]) | (inputs[235]));
    assign layer0_outputs[6666] = ~(inputs[468]);
    assign layer0_outputs[6667] = ~((inputs[236]) ^ (inputs[101]));
    assign layer0_outputs[6668] = 1'b1;
    assign layer0_outputs[6669] = ~((inputs[925]) | (inputs[869]));
    assign layer0_outputs[6670] = ~(inputs[358]);
    assign layer0_outputs[6671] = ~(inputs[626]) | (inputs[683]);
    assign layer0_outputs[6672] = inputs[157];
    assign layer0_outputs[6673] = ~((inputs[594]) ^ (inputs[4]));
    assign layer0_outputs[6674] = ~((inputs[279]) | (inputs[19]));
    assign layer0_outputs[6675] = (inputs[60]) & ~(inputs[447]);
    assign layer0_outputs[6676] = ~((inputs[72]) ^ (inputs[427]));
    assign layer0_outputs[6677] = ~((inputs[595]) | (inputs[407]));
    assign layer0_outputs[6678] = (inputs[104]) ^ (inputs[324]);
    assign layer0_outputs[6679] = ~(inputs[880]);
    assign layer0_outputs[6680] = ~((inputs[601]) | (inputs[28]));
    assign layer0_outputs[6681] = ~((inputs[934]) | (inputs[400]));
    assign layer0_outputs[6682] = inputs[362];
    assign layer0_outputs[6683] = ~((inputs[857]) | (inputs[227]));
    assign layer0_outputs[6684] = (inputs[535]) & ~(inputs[93]);
    assign layer0_outputs[6685] = 1'b0;
    assign layer0_outputs[6686] = ~((inputs[579]) | (inputs[238]));
    assign layer0_outputs[6687] = ~(inputs[988]);
    assign layer0_outputs[6688] = ~((inputs[928]) & (inputs[474]));
    assign layer0_outputs[6689] = ~(inputs[170]) | (inputs[572]);
    assign layer0_outputs[6690] = (inputs[229]) & ~(inputs[484]);
    assign layer0_outputs[6691] = ~((inputs[280]) ^ (inputs[181]));
    assign layer0_outputs[6692] = ~(inputs[426]);
    assign layer0_outputs[6693] = ~((inputs[58]) | (inputs[450]));
    assign layer0_outputs[6694] = ~(inputs[352]) | (inputs[43]);
    assign layer0_outputs[6695] = ~((inputs[22]) & (inputs[136]));
    assign layer0_outputs[6696] = (inputs[1001]) | (inputs[297]);
    assign layer0_outputs[6697] = 1'b0;
    assign layer0_outputs[6698] = (inputs[106]) ^ (inputs[755]);
    assign layer0_outputs[6699] = ~(inputs[682]);
    assign layer0_outputs[6700] = ~(inputs[534]) | (inputs[112]);
    assign layer0_outputs[6701] = (inputs[57]) | (inputs[845]);
    assign layer0_outputs[6702] = 1'b1;
    assign layer0_outputs[6703] = (inputs[493]) & ~(inputs[861]);
    assign layer0_outputs[6704] = (inputs[699]) ^ (inputs[387]);
    assign layer0_outputs[6705] = ~(inputs[732]);
    assign layer0_outputs[6706] = ~(inputs[753]) | (inputs[883]);
    assign layer0_outputs[6707] = ~((inputs[478]) ^ (inputs[954]));
    assign layer0_outputs[6708] = inputs[317];
    assign layer0_outputs[6709] = ~(inputs[660]) | (inputs[421]);
    assign layer0_outputs[6710] = (inputs[882]) & ~(inputs[544]);
    assign layer0_outputs[6711] = (inputs[799]) | (inputs[723]);
    assign layer0_outputs[6712] = 1'b0;
    assign layer0_outputs[6713] = inputs[645];
    assign layer0_outputs[6714] = ~(inputs[530]);
    assign layer0_outputs[6715] = inputs[894];
    assign layer0_outputs[6716] = (inputs[723]) | (inputs[45]);
    assign layer0_outputs[6717] = ~((inputs[427]) ^ (inputs[29]));
    assign layer0_outputs[6718] = ~((inputs[989]) | (inputs[101]));
    assign layer0_outputs[6719] = ~((inputs[382]) | (inputs[97]));
    assign layer0_outputs[6720] = (inputs[511]) | (inputs[200]);
    assign layer0_outputs[6721] = ~((inputs[828]) | (inputs[763]));
    assign layer0_outputs[6722] = (inputs[782]) & ~(inputs[76]);
    assign layer0_outputs[6723] = (inputs[268]) | (inputs[950]);
    assign layer0_outputs[6724] = (inputs[657]) | (inputs[711]);
    assign layer0_outputs[6725] = ~((inputs[696]) | (inputs[752]));
    assign layer0_outputs[6726] = ~(inputs[243]);
    assign layer0_outputs[6727] = ~((inputs[478]) & (inputs[573]));
    assign layer0_outputs[6728] = ~(inputs[309]);
    assign layer0_outputs[6729] = ~(inputs[548]);
    assign layer0_outputs[6730] = ~(inputs[839]) | (inputs[640]);
    assign layer0_outputs[6731] = (inputs[966]) | (inputs[483]);
    assign layer0_outputs[6732] = (inputs[1002]) & ~(inputs[422]);
    assign layer0_outputs[6733] = ~((inputs[381]) ^ (inputs[875]));
    assign layer0_outputs[6734] = (inputs[530]) & ~(inputs[906]);
    assign layer0_outputs[6735] = ~(inputs[614]);
    assign layer0_outputs[6736] = (inputs[459]) & ~(inputs[58]);
    assign layer0_outputs[6737] = inputs[992];
    assign layer0_outputs[6738] = ~((inputs[385]) & (inputs[611]));
    assign layer0_outputs[6739] = (inputs[337]) ^ (inputs[485]);
    assign layer0_outputs[6740] = (inputs[563]) & ~(inputs[748]);
    assign layer0_outputs[6741] = ~((inputs[215]) ^ (inputs[577]));
    assign layer0_outputs[6742] = ~(inputs[209]);
    assign layer0_outputs[6743] = (inputs[806]) & ~(inputs[775]);
    assign layer0_outputs[6744] = ~((inputs[316]) | (inputs[74]));
    assign layer0_outputs[6745] = inputs[92];
    assign layer0_outputs[6746] = inputs[330];
    assign layer0_outputs[6747] = inputs[917];
    assign layer0_outputs[6748] = inputs[651];
    assign layer0_outputs[6749] = ~((inputs[226]) | (inputs[737]));
    assign layer0_outputs[6750] = ~((inputs[900]) ^ (inputs[230]));
    assign layer0_outputs[6751] = ~((inputs[181]) | (inputs[98]));
    assign layer0_outputs[6752] = ~(inputs[713]) | (inputs[877]);
    assign layer0_outputs[6753] = ~(inputs[1015]);
    assign layer0_outputs[6754] = (inputs[401]) & ~(inputs[665]);
    assign layer0_outputs[6755] = ~((inputs[406]) ^ (inputs[639]));
    assign layer0_outputs[6756] = (inputs[288]) & ~(inputs[982]);
    assign layer0_outputs[6757] = (inputs[763]) & (inputs[7]);
    assign layer0_outputs[6758] = ~((inputs[240]) ^ (inputs[824]));
    assign layer0_outputs[6759] = ~(inputs[945]);
    assign layer0_outputs[6760] = (inputs[830]) & (inputs[936]);
    assign layer0_outputs[6761] = ~((inputs[337]) | (inputs[195]));
    assign layer0_outputs[6762] = ~(inputs[956]);
    assign layer0_outputs[6763] = ~(inputs[1023]);
    assign layer0_outputs[6764] = ~(inputs[620]);
    assign layer0_outputs[6765] = ~(inputs[506]) | (inputs[99]);
    assign layer0_outputs[6766] = ~((inputs[511]) ^ (inputs[439]));
    assign layer0_outputs[6767] = inputs[37];
    assign layer0_outputs[6768] = 1'b1;
    assign layer0_outputs[6769] = (inputs[0]) | (inputs[704]);
    assign layer0_outputs[6770] = ~((inputs[679]) ^ (inputs[921]));
    assign layer0_outputs[6771] = 1'b0;
    assign layer0_outputs[6772] = (inputs[233]) & ~(inputs[545]);
    assign layer0_outputs[6773] = (inputs[68]) | (inputs[463]);
    assign layer0_outputs[6774] = ~(inputs[653]);
    assign layer0_outputs[6775] = (inputs[413]) & (inputs[39]);
    assign layer0_outputs[6776] = inputs[622];
    assign layer0_outputs[6777] = ~(inputs[851]);
    assign layer0_outputs[6778] = (inputs[935]) ^ (inputs[91]);
    assign layer0_outputs[6779] = ~(inputs[617]) | (inputs[434]);
    assign layer0_outputs[6780] = ~(inputs[314]);
    assign layer0_outputs[6781] = 1'b1;
    assign layer0_outputs[6782] = ~(inputs[395]) | (inputs[294]);
    assign layer0_outputs[6783] = (inputs[972]) | (inputs[89]);
    assign layer0_outputs[6784] = (inputs[690]) & ~(inputs[335]);
    assign layer0_outputs[6785] = ~((inputs[166]) | (inputs[621]));
    assign layer0_outputs[6786] = (inputs[291]) & (inputs[515]);
    assign layer0_outputs[6787] = ~(inputs[1020]) | (inputs[299]);
    assign layer0_outputs[6788] = (inputs[433]) | (inputs[197]);
    assign layer0_outputs[6789] = (inputs[796]) | (inputs[408]);
    assign layer0_outputs[6790] = inputs[610];
    assign layer0_outputs[6791] = 1'b0;
    assign layer0_outputs[6792] = ~(inputs[949]);
    assign layer0_outputs[6793] = ~((inputs[605]) ^ (inputs[759]));
    assign layer0_outputs[6794] = inputs[215];
    assign layer0_outputs[6795] = (inputs[947]) ^ (inputs[893]);
    assign layer0_outputs[6796] = (inputs[834]) & (inputs[107]);
    assign layer0_outputs[6797] = ~((inputs[179]) | (inputs[217]));
    assign layer0_outputs[6798] = ~((inputs[397]) ^ (inputs[389]));
    assign layer0_outputs[6799] = ~(inputs[129]) | (inputs[602]);
    assign layer0_outputs[6800] = (inputs[646]) | (inputs[906]);
    assign layer0_outputs[6801] = (inputs[174]) ^ (inputs[501]);
    assign layer0_outputs[6802] = ~((inputs[960]) | (inputs[793]));
    assign layer0_outputs[6803] = (inputs[504]) | (inputs[583]);
    assign layer0_outputs[6804] = (inputs[331]) | (inputs[854]);
    assign layer0_outputs[6805] = (inputs[679]) & ~(inputs[997]);
    assign layer0_outputs[6806] = (inputs[356]) & ~(inputs[559]);
    assign layer0_outputs[6807] = ~((inputs[262]) | (inputs[565]));
    assign layer0_outputs[6808] = inputs[360];
    assign layer0_outputs[6809] = ~((inputs[216]) | (inputs[455]));
    assign layer0_outputs[6810] = (inputs[110]) | (inputs[293]);
    assign layer0_outputs[6811] = ~((inputs[388]) ^ (inputs[500]));
    assign layer0_outputs[6812] = ~((inputs[716]) | (inputs[200]));
    assign layer0_outputs[6813] = (inputs[403]) | (inputs[236]);
    assign layer0_outputs[6814] = (inputs[198]) | (inputs[341]);
    assign layer0_outputs[6815] = ~(inputs[494]) | (inputs[226]);
    assign layer0_outputs[6816] = ~((inputs[230]) ^ (inputs[404]));
    assign layer0_outputs[6817] = ~(inputs[137]) | (inputs[676]);
    assign layer0_outputs[6818] = inputs[641];
    assign layer0_outputs[6819] = ~((inputs[224]) ^ (inputs[64]));
    assign layer0_outputs[6820] = ~(inputs[128]);
    assign layer0_outputs[6821] = ~(inputs[948]);
    assign layer0_outputs[6822] = ~((inputs[621]) ^ (inputs[222]));
    assign layer0_outputs[6823] = (inputs[552]) ^ (inputs[894]);
    assign layer0_outputs[6824] = (inputs[38]) & (inputs[482]);
    assign layer0_outputs[6825] = ~((inputs[821]) ^ (inputs[614]));
    assign layer0_outputs[6826] = ~((inputs[435]) | (inputs[391]));
    assign layer0_outputs[6827] = inputs[530];
    assign layer0_outputs[6828] = (inputs[567]) & (inputs[324]);
    assign layer0_outputs[6829] = ~((inputs[235]) | (inputs[115]));
    assign layer0_outputs[6830] = ~((inputs[862]) ^ (inputs[833]));
    assign layer0_outputs[6831] = ~((inputs[138]) | (inputs[763]));
    assign layer0_outputs[6832] = inputs[651];
    assign layer0_outputs[6833] = inputs[957];
    assign layer0_outputs[6834] = ~((inputs[230]) | (inputs[740]));
    assign layer0_outputs[6835] = (inputs[718]) & ~(inputs[516]);
    assign layer0_outputs[6836] = (inputs[334]) | (inputs[837]);
    assign layer0_outputs[6837] = ~((inputs[567]) | (inputs[447]));
    assign layer0_outputs[6838] = (inputs[305]) & ~(inputs[85]);
    assign layer0_outputs[6839] = inputs[443];
    assign layer0_outputs[6840] = ~(inputs[685]) | (inputs[49]);
    assign layer0_outputs[6841] = ~((inputs[198]) | (inputs[371]));
    assign layer0_outputs[6842] = ~((inputs[788]) | (inputs[708]));
    assign layer0_outputs[6843] = (inputs[500]) | (inputs[530]);
    assign layer0_outputs[6844] = ~(inputs[755]) | (inputs[392]);
    assign layer0_outputs[6845] = (inputs[634]) & ~(inputs[102]);
    assign layer0_outputs[6846] = (inputs[376]) | (inputs[205]);
    assign layer0_outputs[6847] = (inputs[941]) ^ (inputs[970]);
    assign layer0_outputs[6848] = ~(inputs[591]);
    assign layer0_outputs[6849] = (inputs[105]) ^ (inputs[438]);
    assign layer0_outputs[6850] = ~((inputs[872]) ^ (inputs[520]));
    assign layer0_outputs[6851] = (inputs[46]) & (inputs[574]);
    assign layer0_outputs[6852] = ~(inputs[114]) | (inputs[383]);
    assign layer0_outputs[6853] = ~((inputs[688]) | (inputs[101]));
    assign layer0_outputs[6854] = (inputs[270]) | (inputs[337]);
    assign layer0_outputs[6855] = ~((inputs[681]) | (inputs[906]));
    assign layer0_outputs[6856] = (inputs[344]) ^ (inputs[802]);
    assign layer0_outputs[6857] = ~(inputs[206]) | (inputs[1000]);
    assign layer0_outputs[6858] = (inputs[213]) & (inputs[777]);
    assign layer0_outputs[6859] = (inputs[683]) | (inputs[8]);
    assign layer0_outputs[6860] = ~((inputs[71]) ^ (inputs[89]));
    assign layer0_outputs[6861] = ~((inputs[127]) | (inputs[809]));
    assign layer0_outputs[6862] = ~((inputs[395]) ^ (inputs[970]));
    assign layer0_outputs[6863] = ~(inputs[563]);
    assign layer0_outputs[6864] = ~(inputs[325]);
    assign layer0_outputs[6865] = inputs[650];
    assign layer0_outputs[6866] = 1'b1;
    assign layer0_outputs[6867] = ~((inputs[113]) ^ (inputs[429]));
    assign layer0_outputs[6868] = (inputs[105]) & (inputs[1018]);
    assign layer0_outputs[6869] = (inputs[281]) ^ (inputs[144]);
    assign layer0_outputs[6870] = (inputs[869]) & (inputs[219]);
    assign layer0_outputs[6871] = (inputs[38]) & (inputs[2]);
    assign layer0_outputs[6872] = inputs[527];
    assign layer0_outputs[6873] = (inputs[591]) | (inputs[738]);
    assign layer0_outputs[6874] = inputs[255];
    assign layer0_outputs[6875] = inputs[304];
    assign layer0_outputs[6876] = inputs[441];
    assign layer0_outputs[6877] = ~(inputs[820]);
    assign layer0_outputs[6878] = 1'b0;
    assign layer0_outputs[6879] = 1'b1;
    assign layer0_outputs[6880] = inputs[698];
    assign layer0_outputs[6881] = ~(inputs[416]) | (inputs[421]);
    assign layer0_outputs[6882] = ~((inputs[952]) ^ (inputs[542]));
    assign layer0_outputs[6883] = (inputs[946]) & ~(inputs[83]);
    assign layer0_outputs[6884] = ~(inputs[595]) | (inputs[519]);
    assign layer0_outputs[6885] = ~(inputs[668]) | (inputs[415]);
    assign layer0_outputs[6886] = (inputs[687]) & ~(inputs[571]);
    assign layer0_outputs[6887] = (inputs[70]) | (inputs[302]);
    assign layer0_outputs[6888] = (inputs[158]) & ~(inputs[647]);
    assign layer0_outputs[6889] = ~((inputs[833]) | (inputs[812]));
    assign layer0_outputs[6890] = ~((inputs[670]) ^ (inputs[754]));
    assign layer0_outputs[6891] = (inputs[167]) ^ (inputs[530]);
    assign layer0_outputs[6892] = inputs[717];
    assign layer0_outputs[6893] = ~((inputs[828]) ^ (inputs[356]));
    assign layer0_outputs[6894] = ~(inputs[870]) | (inputs[349]);
    assign layer0_outputs[6895] = inputs[871];
    assign layer0_outputs[6896] = inputs[694];
    assign layer0_outputs[6897] = (inputs[307]) & ~(inputs[74]);
    assign layer0_outputs[6898] = ~((inputs[223]) | (inputs[938]));
    assign layer0_outputs[6899] = 1'b0;
    assign layer0_outputs[6900] = ~(inputs[622]) | (inputs[614]);
    assign layer0_outputs[6901] = ~(inputs[194]);
    assign layer0_outputs[6902] = ~((inputs[278]) | (inputs[66]));
    assign layer0_outputs[6903] = (inputs[306]) | (inputs[378]);
    assign layer0_outputs[6904] = inputs[516];
    assign layer0_outputs[6905] = (inputs[629]) & ~(inputs[783]);
    assign layer0_outputs[6906] = inputs[835];
    assign layer0_outputs[6907] = (inputs[664]) ^ (inputs[762]);
    assign layer0_outputs[6908] = ~(inputs[705]);
    assign layer0_outputs[6909] = inputs[366];
    assign layer0_outputs[6910] = (inputs[369]) | (inputs[806]);
    assign layer0_outputs[6911] = ~((inputs[135]) | (inputs[570]));
    assign layer0_outputs[6912] = (inputs[301]) & ~(inputs[136]);
    assign layer0_outputs[6913] = (inputs[627]) ^ (inputs[449]);
    assign layer0_outputs[6914] = ~(inputs[699]) | (inputs[675]);
    assign layer0_outputs[6915] = ~((inputs[74]) & (inputs[978]));
    assign layer0_outputs[6916] = (inputs[985]) | (inputs[304]);
    assign layer0_outputs[6917] = (inputs[465]) ^ (inputs[589]);
    assign layer0_outputs[6918] = ~((inputs[84]) ^ (inputs[620]));
    assign layer0_outputs[6919] = ~(inputs[149]);
    assign layer0_outputs[6920] = ~(inputs[426]) | (inputs[758]);
    assign layer0_outputs[6921] = ~(inputs[430]);
    assign layer0_outputs[6922] = ~(inputs[231]) | (inputs[897]);
    assign layer0_outputs[6923] = ~(inputs[725]) | (inputs[67]);
    assign layer0_outputs[6924] = ~((inputs[650]) ^ (inputs[243]));
    assign layer0_outputs[6925] = ~((inputs[223]) | (inputs[44]));
    assign layer0_outputs[6926] = ~((inputs[195]) & (inputs[88]));
    assign layer0_outputs[6927] = ~(inputs[246]);
    assign layer0_outputs[6928] = (inputs[458]) & ~(inputs[733]);
    assign layer0_outputs[6929] = ~((inputs[798]) | (inputs[652]));
    assign layer0_outputs[6930] = 1'b0;
    assign layer0_outputs[6931] = ~((inputs[949]) | (inputs[310]));
    assign layer0_outputs[6932] = (inputs[198]) ^ (inputs[474]);
    assign layer0_outputs[6933] = ~(inputs[816]) | (inputs[985]);
    assign layer0_outputs[6934] = ~((inputs[452]) & (inputs[73]));
    assign layer0_outputs[6935] = ~((inputs[732]) ^ (inputs[291]));
    assign layer0_outputs[6936] = ~(inputs[848]) | (inputs[319]);
    assign layer0_outputs[6937] = inputs[412];
    assign layer0_outputs[6938] = (inputs[911]) | (inputs[411]);
    assign layer0_outputs[6939] = inputs[148];
    assign layer0_outputs[6940] = (inputs[179]) | (inputs[779]);
    assign layer0_outputs[6941] = ~((inputs[802]) | (inputs[375]));
    assign layer0_outputs[6942] = 1'b1;
    assign layer0_outputs[6943] = ~(inputs[405]);
    assign layer0_outputs[6944] = (inputs[467]) & ~(inputs[348]);
    assign layer0_outputs[6945] = (inputs[386]) ^ (inputs[556]);
    assign layer0_outputs[6946] = (inputs[515]) | (inputs[438]);
    assign layer0_outputs[6947] = ~(inputs[358]) | (inputs[887]);
    assign layer0_outputs[6948] = ~(inputs[719]);
    assign layer0_outputs[6949] = ~(inputs[853]);
    assign layer0_outputs[6950] = (inputs[563]) & ~(inputs[645]);
    assign layer0_outputs[6951] = ~((inputs[0]) ^ (inputs[530]));
    assign layer0_outputs[6952] = ~(inputs[941]) | (inputs[72]);
    assign layer0_outputs[6953] = ~(inputs[598]);
    assign layer0_outputs[6954] = ~((inputs[985]) | (inputs[473]));
    assign layer0_outputs[6955] = ~(inputs[926]) | (inputs[135]);
    assign layer0_outputs[6956] = ~((inputs[606]) ^ (inputs[290]));
    assign layer0_outputs[6957] = ~((inputs[616]) ^ (inputs[381]));
    assign layer0_outputs[6958] = (inputs[178]) ^ (inputs[351]);
    assign layer0_outputs[6959] = ~(inputs[621]);
    assign layer0_outputs[6960] = ~((inputs[975]) | (inputs[949]));
    assign layer0_outputs[6961] = ~(inputs[266]) | (inputs[551]);
    assign layer0_outputs[6962] = inputs[520];
    assign layer0_outputs[6963] = (inputs[891]) | (inputs[936]);
    assign layer0_outputs[6964] = 1'b1;
    assign layer0_outputs[6965] = inputs[175];
    assign layer0_outputs[6966] = (inputs[227]) | (inputs[708]);
    assign layer0_outputs[6967] = (inputs[389]) | (inputs[712]);
    assign layer0_outputs[6968] = ~((inputs[974]) | (inputs[668]));
    assign layer0_outputs[6969] = (inputs[446]) ^ (inputs[273]);
    assign layer0_outputs[6970] = ~(inputs[652]);
    assign layer0_outputs[6971] = ~((inputs[565]) | (inputs[672]));
    assign layer0_outputs[6972] = ~(inputs[589]) | (inputs[58]);
    assign layer0_outputs[6973] = inputs[755];
    assign layer0_outputs[6974] = ~((inputs[408]) | (inputs[627]));
    assign layer0_outputs[6975] = ~((inputs[111]) ^ (inputs[197]));
    assign layer0_outputs[6976] = ~(inputs[581]) | (inputs[639]);
    assign layer0_outputs[6977] = inputs[395];
    assign layer0_outputs[6978] = ~((inputs[922]) | (inputs[489]));
    assign layer0_outputs[6979] = ~(inputs[772]) | (inputs[161]);
    assign layer0_outputs[6980] = ~((inputs[808]) & (inputs[468]));
    assign layer0_outputs[6981] = ~((inputs[491]) | (inputs[283]));
    assign layer0_outputs[6982] = ~(inputs[614]);
    assign layer0_outputs[6983] = ~(inputs[242]) | (inputs[13]);
    assign layer0_outputs[6984] = ~(inputs[86]) | (inputs[549]);
    assign layer0_outputs[6985] = ~(inputs[169]) | (inputs[700]);
    assign layer0_outputs[6986] = ~((inputs[183]) | (inputs[647]));
    assign layer0_outputs[6987] = ~((inputs[169]) ^ (inputs[891]));
    assign layer0_outputs[6988] = 1'b0;
    assign layer0_outputs[6989] = (inputs[179]) | (inputs[196]);
    assign layer0_outputs[6990] = ~(inputs[166]);
    assign layer0_outputs[6991] = (inputs[283]) | (inputs[130]);
    assign layer0_outputs[6992] = ~((inputs[445]) | (inputs[34]));
    assign layer0_outputs[6993] = (inputs[795]) ^ (inputs[818]);
    assign layer0_outputs[6994] = ~((inputs[255]) & (inputs[651]));
    assign layer0_outputs[6995] = ~(inputs[274]) | (inputs[903]);
    assign layer0_outputs[6996] = 1'b1;
    assign layer0_outputs[6997] = ~((inputs[761]) | (inputs[762]));
    assign layer0_outputs[6998] = ~(inputs[695]) | (inputs[981]);
    assign layer0_outputs[6999] = 1'b0;
    assign layer0_outputs[7000] = (inputs[252]) & ~(inputs[146]);
    assign layer0_outputs[7001] = (inputs[737]) | (inputs[660]);
    assign layer0_outputs[7002] = ~((inputs[679]) | (inputs[585]));
    assign layer0_outputs[7003] = ~(inputs[411]);
    assign layer0_outputs[7004] = ~(inputs[624]) | (inputs[668]);
    assign layer0_outputs[7005] = ~((inputs[332]) ^ (inputs[335]));
    assign layer0_outputs[7006] = ~((inputs[421]) | (inputs[326]));
    assign layer0_outputs[7007] = inputs[430];
    assign layer0_outputs[7008] = ~(inputs[185]) | (inputs[110]);
    assign layer0_outputs[7009] = (inputs[922]) ^ (inputs[180]);
    assign layer0_outputs[7010] = ~(inputs[364]) | (inputs[86]);
    assign layer0_outputs[7011] = (inputs[617]) & ~(inputs[175]);
    assign layer0_outputs[7012] = ~(inputs[386]);
    assign layer0_outputs[7013] = (inputs[976]) & ~(inputs[587]);
    assign layer0_outputs[7014] = inputs[403];
    assign layer0_outputs[7015] = inputs[550];
    assign layer0_outputs[7016] = ~((inputs[358]) ^ (inputs[576]));
    assign layer0_outputs[7017] = ~((inputs[697]) ^ (inputs[604]));
    assign layer0_outputs[7018] = (inputs[928]) ^ (inputs[490]);
    assign layer0_outputs[7019] = inputs[762];
    assign layer0_outputs[7020] = (inputs[582]) ^ (inputs[195]);
    assign layer0_outputs[7021] = ~(inputs[882]) | (inputs[531]);
    assign layer0_outputs[7022] = 1'b1;
    assign layer0_outputs[7023] = ~((inputs[147]) & (inputs[899]));
    assign layer0_outputs[7024] = inputs[648];
    assign layer0_outputs[7025] = (inputs[278]) & ~(inputs[874]);
    assign layer0_outputs[7026] = ~((inputs[240]) | (inputs[490]));
    assign layer0_outputs[7027] = ~(inputs[712]);
    assign layer0_outputs[7028] = ~(inputs[590]) | (inputs[237]);
    assign layer0_outputs[7029] = ~(inputs[300]);
    assign layer0_outputs[7030] = (inputs[318]) | (inputs[744]);
    assign layer0_outputs[7031] = ~(inputs[563]);
    assign layer0_outputs[7032] = ~((inputs[595]) | (inputs[414]));
    assign layer0_outputs[7033] = ~((inputs[400]) ^ (inputs[697]));
    assign layer0_outputs[7034] = inputs[308];
    assign layer0_outputs[7035] = ~(inputs[251]);
    assign layer0_outputs[7036] = ~(inputs[634]) | (inputs[351]);
    assign layer0_outputs[7037] = ~(inputs[302]) | (inputs[680]);
    assign layer0_outputs[7038] = (inputs[791]) ^ (inputs[48]);
    assign layer0_outputs[7039] = (inputs[755]) & ~(inputs[768]);
    assign layer0_outputs[7040] = (inputs[160]) ^ (inputs[149]);
    assign layer0_outputs[7041] = (inputs[847]) & ~(inputs[636]);
    assign layer0_outputs[7042] = (inputs[934]) & (inputs[324]);
    assign layer0_outputs[7043] = inputs[71];
    assign layer0_outputs[7044] = (inputs[761]) ^ (inputs[489]);
    assign layer0_outputs[7045] = (inputs[442]) & ~(inputs[1021]);
    assign layer0_outputs[7046] = ~(inputs[699]) | (inputs[996]);
    assign layer0_outputs[7047] = ~((inputs[973]) | (inputs[711]));
    assign layer0_outputs[7048] = inputs[346];
    assign layer0_outputs[7049] = inputs[520];
    assign layer0_outputs[7050] = ~((inputs[793]) ^ (inputs[3]));
    assign layer0_outputs[7051] = ~(inputs[209]) | (inputs[157]);
    assign layer0_outputs[7052] = (inputs[98]) & ~(inputs[738]);
    assign layer0_outputs[7053] = (inputs[315]) ^ (inputs[60]);
    assign layer0_outputs[7054] = inputs[707];
    assign layer0_outputs[7055] = ~((inputs[963]) | (inputs[866]));
    assign layer0_outputs[7056] = ~(inputs[913]) | (inputs[46]);
    assign layer0_outputs[7057] = ~((inputs[867]) ^ (inputs[168]));
    assign layer0_outputs[7058] = ~((inputs[114]) & (inputs[79]));
    assign layer0_outputs[7059] = ~(inputs[56]) | (inputs[923]);
    assign layer0_outputs[7060] = ~(inputs[493]);
    assign layer0_outputs[7061] = (inputs[839]) & ~(inputs[889]);
    assign layer0_outputs[7062] = ~((inputs[755]) | (inputs[258]));
    assign layer0_outputs[7063] = (inputs[49]) ^ (inputs[694]);
    assign layer0_outputs[7064] = ~((inputs[222]) ^ (inputs[384]));
    assign layer0_outputs[7065] = ~((inputs[723]) & (inputs[751]));
    assign layer0_outputs[7066] = (inputs[129]) ^ (inputs[1003]);
    assign layer0_outputs[7067] = (inputs[943]) & ~(inputs[646]);
    assign layer0_outputs[7068] = ~((inputs[185]) | (inputs[474]));
    assign layer0_outputs[7069] = (inputs[822]) | (inputs[601]);
    assign layer0_outputs[7070] = (inputs[470]) | (inputs[25]);
    assign layer0_outputs[7071] = (inputs[956]) & (inputs[897]);
    assign layer0_outputs[7072] = ~(inputs[577]);
    assign layer0_outputs[7073] = ~((inputs[426]) ^ (inputs[168]));
    assign layer0_outputs[7074] = (inputs[356]) | (inputs[399]);
    assign layer0_outputs[7075] = inputs[244];
    assign layer0_outputs[7076] = ~((inputs[72]) ^ (inputs[942]));
    assign layer0_outputs[7077] = (inputs[691]) | (inputs[988]);
    assign layer0_outputs[7078] = ~(inputs[268]) | (inputs[906]);
    assign layer0_outputs[7079] = (inputs[1009]) | (inputs[250]);
    assign layer0_outputs[7080] = (inputs[831]) ^ (inputs[424]);
    assign layer0_outputs[7081] = (inputs[889]) & ~(inputs[965]);
    assign layer0_outputs[7082] = (inputs[886]) & (inputs[166]);
    assign layer0_outputs[7083] = inputs[433];
    assign layer0_outputs[7084] = (inputs[570]) ^ (inputs[482]);
    assign layer0_outputs[7085] = (inputs[854]) & ~(inputs[979]);
    assign layer0_outputs[7086] = inputs[749];
    assign layer0_outputs[7087] = ~((inputs[31]) & (inputs[261]));
    assign layer0_outputs[7088] = ~(inputs[513]) | (inputs[677]);
    assign layer0_outputs[7089] = 1'b0;
    assign layer0_outputs[7090] = inputs[808];
    assign layer0_outputs[7091] = ~((inputs[565]) ^ (inputs[764]));
    assign layer0_outputs[7092] = (inputs[208]) & ~(inputs[197]);
    assign layer0_outputs[7093] = (inputs[347]) | (inputs[930]);
    assign layer0_outputs[7094] = ~(inputs[120]) | (inputs[931]);
    assign layer0_outputs[7095] = ~(inputs[1012]);
    assign layer0_outputs[7096] = ~((inputs[808]) ^ (inputs[954]));
    assign layer0_outputs[7097] = ~((inputs[654]) | (inputs[548]));
    assign layer0_outputs[7098] = 1'b1;
    assign layer0_outputs[7099] = inputs[261];
    assign layer0_outputs[7100] = (inputs[566]) & ~(inputs[406]);
    assign layer0_outputs[7101] = ~((inputs[40]) | (inputs[289]));
    assign layer0_outputs[7102] = ~(inputs[463]) | (inputs[893]);
    assign layer0_outputs[7103] = (inputs[339]) & ~(inputs[700]);
    assign layer0_outputs[7104] = 1'b1;
    assign layer0_outputs[7105] = (inputs[471]) ^ (inputs[703]);
    assign layer0_outputs[7106] = ~(inputs[282]);
    assign layer0_outputs[7107] = (inputs[421]) & ~(inputs[262]);
    assign layer0_outputs[7108] = ~((inputs[491]) ^ (inputs[37]));
    assign layer0_outputs[7109] = (inputs[782]) & ~(inputs[873]);
    assign layer0_outputs[7110] = ~(inputs[472]) | (inputs[54]);
    assign layer0_outputs[7111] = (inputs[223]) ^ (inputs[837]);
    assign layer0_outputs[7112] = ~(inputs[646]);
    assign layer0_outputs[7113] = (inputs[320]) ^ (inputs[742]);
    assign layer0_outputs[7114] = ~((inputs[5]) ^ (inputs[982]));
    assign layer0_outputs[7115] = ~(inputs[418]) | (inputs[994]);
    assign layer0_outputs[7116] = ~(inputs[336]) | (inputs[143]);
    assign layer0_outputs[7117] = ~((inputs[249]) | (inputs[208]));
    assign layer0_outputs[7118] = ~(inputs[454]);
    assign layer0_outputs[7119] = (inputs[710]) & ~(inputs[159]);
    assign layer0_outputs[7120] = ~((inputs[208]) | (inputs[17]));
    assign layer0_outputs[7121] = (inputs[632]) | (inputs[692]);
    assign layer0_outputs[7122] = inputs[119];
    assign layer0_outputs[7123] = (inputs[873]) | (inputs[350]);
    assign layer0_outputs[7124] = ~((inputs[211]) ^ (inputs[51]));
    assign layer0_outputs[7125] = ~(inputs[758]) | (inputs[996]);
    assign layer0_outputs[7126] = (inputs[416]) & ~(inputs[786]);
    assign layer0_outputs[7127] = ~((inputs[97]) ^ (inputs[962]));
    assign layer0_outputs[7128] = ~((inputs[646]) | (inputs[552]));
    assign layer0_outputs[7129] = ~((inputs[912]) | (inputs[482]));
    assign layer0_outputs[7130] = ~((inputs[313]) | (inputs[605]));
    assign layer0_outputs[7131] = 1'b1;
    assign layer0_outputs[7132] = (inputs[880]) ^ (inputs[310]);
    assign layer0_outputs[7133] = inputs[962];
    assign layer0_outputs[7134] = ~(inputs[248]);
    assign layer0_outputs[7135] = ~((inputs[308]) | (inputs[3]));
    assign layer0_outputs[7136] = inputs[749];
    assign layer0_outputs[7137] = ~(inputs[915]);
    assign layer0_outputs[7138] = 1'b1;
    assign layer0_outputs[7139] = ~(inputs[258]);
    assign layer0_outputs[7140] = ~((inputs[1004]) ^ (inputs[248]));
    assign layer0_outputs[7141] = ~((inputs[269]) ^ (inputs[722]));
    assign layer0_outputs[7142] = ~(inputs[265]);
    assign layer0_outputs[7143] = (inputs[15]) ^ (inputs[308]);
    assign layer0_outputs[7144] = inputs[824];
    assign layer0_outputs[7145] = ~(inputs[683]) | (inputs[554]);
    assign layer0_outputs[7146] = ~((inputs[9]) ^ (inputs[666]));
    assign layer0_outputs[7147] = inputs[253];
    assign layer0_outputs[7148] = (inputs[644]) & (inputs[708]);
    assign layer0_outputs[7149] = ~(inputs[69]);
    assign layer0_outputs[7150] = ~(inputs[914]) | (inputs[604]);
    assign layer0_outputs[7151] = ~(inputs[309]) | (inputs[796]);
    assign layer0_outputs[7152] = ~(inputs[905]) | (inputs[576]);
    assign layer0_outputs[7153] = (inputs[796]) | (inputs[959]);
    assign layer0_outputs[7154] = (inputs[615]) ^ (inputs[93]);
    assign layer0_outputs[7155] = ~((inputs[167]) ^ (inputs[942]));
    assign layer0_outputs[7156] = ~((inputs[797]) ^ (inputs[517]));
    assign layer0_outputs[7157] = (inputs[786]) ^ (inputs[788]);
    assign layer0_outputs[7158] = (inputs[526]) | (inputs[204]);
    assign layer0_outputs[7159] = ~(inputs[1009]);
    assign layer0_outputs[7160] = ~((inputs[228]) ^ (inputs[625]));
    assign layer0_outputs[7161] = ~((inputs[5]) ^ (inputs[931]));
    assign layer0_outputs[7162] = (inputs[460]) ^ (inputs[425]);
    assign layer0_outputs[7163] = 1'b1;
    assign layer0_outputs[7164] = (inputs[630]) | (inputs[263]);
    assign layer0_outputs[7165] = ~((inputs[455]) ^ (inputs[255]));
    assign layer0_outputs[7166] = ~((inputs[173]) & (inputs[39]));
    assign layer0_outputs[7167] = 1'b0;
    assign layer0_outputs[7168] = ~(inputs[852]) | (inputs[106]);
    assign layer0_outputs[7169] = ~(inputs[458]) | (inputs[633]);
    assign layer0_outputs[7170] = (inputs[297]) & ~(inputs[182]);
    assign layer0_outputs[7171] = ~((inputs[406]) | (inputs[973]));
    assign layer0_outputs[7172] = (inputs[252]) | (inputs[883]);
    assign layer0_outputs[7173] = inputs[404];
    assign layer0_outputs[7174] = inputs[438];
    assign layer0_outputs[7175] = (inputs[239]) ^ (inputs[993]);
    assign layer0_outputs[7176] = ~((inputs[652]) | (inputs[186]));
    assign layer0_outputs[7177] = ~((inputs[439]) | (inputs[127]));
    assign layer0_outputs[7178] = ~(inputs[279]);
    assign layer0_outputs[7179] = (inputs[536]) | (inputs[136]);
    assign layer0_outputs[7180] = 1'b0;
    assign layer0_outputs[7181] = ~(inputs[908]);
    assign layer0_outputs[7182] = ~((inputs[286]) ^ (inputs[141]));
    assign layer0_outputs[7183] = (inputs[626]) ^ (inputs[67]);
    assign layer0_outputs[7184] = ~((inputs[472]) | (inputs[471]));
    assign layer0_outputs[7185] = ~((inputs[750]) | (inputs[357]));
    assign layer0_outputs[7186] = (inputs[653]) | (inputs[611]);
    assign layer0_outputs[7187] = ~((inputs[914]) | (inputs[689]));
    assign layer0_outputs[7188] = (inputs[690]) | (inputs[501]);
    assign layer0_outputs[7189] = ~(inputs[672]);
    assign layer0_outputs[7190] = (inputs[499]) | (inputs[669]);
    assign layer0_outputs[7191] = ~(inputs[806]);
    assign layer0_outputs[7192] = 1'b0;
    assign layer0_outputs[7193] = ~(inputs[431]);
    assign layer0_outputs[7194] = ~((inputs[1019]) ^ (inputs[367]));
    assign layer0_outputs[7195] = (inputs[632]) | (inputs[289]);
    assign layer0_outputs[7196] = ~((inputs[681]) ^ (inputs[354]));
    assign layer0_outputs[7197] = ~(inputs[41]);
    assign layer0_outputs[7198] = ~((inputs[735]) & (inputs[944]));
    assign layer0_outputs[7199] = ~(inputs[871]) | (inputs[253]);
    assign layer0_outputs[7200] = ~((inputs[843]) | (inputs[177]));
    assign layer0_outputs[7201] = (inputs[841]) & ~(inputs[76]);
    assign layer0_outputs[7202] = ~(inputs[32]);
    assign layer0_outputs[7203] = (inputs[486]) | (inputs[743]);
    assign layer0_outputs[7204] = (inputs[938]) ^ (inputs[1007]);
    assign layer0_outputs[7205] = ~((inputs[162]) | (inputs[435]));
    assign layer0_outputs[7206] = ~((inputs[24]) | (inputs[992]));
    assign layer0_outputs[7207] = ~(inputs[413]);
    assign layer0_outputs[7208] = ~(inputs[101]) | (inputs[792]);
    assign layer0_outputs[7209] = inputs[969];
    assign layer0_outputs[7210] = (inputs[700]) & (inputs[71]);
    assign layer0_outputs[7211] = (inputs[306]) & (inputs[631]);
    assign layer0_outputs[7212] = inputs[489];
    assign layer0_outputs[7213] = ~(inputs[645]) | (inputs[674]);
    assign layer0_outputs[7214] = ~((inputs[212]) | (inputs[694]));
    assign layer0_outputs[7215] = (inputs[671]) & ~(inputs[10]);
    assign layer0_outputs[7216] = (inputs[642]) | (inputs[788]);
    assign layer0_outputs[7217] = (inputs[711]) | (inputs[788]);
    assign layer0_outputs[7218] = ~((inputs[825]) | (inputs[118]));
    assign layer0_outputs[7219] = inputs[921];
    assign layer0_outputs[7220] = (inputs[234]) | (inputs[162]);
    assign layer0_outputs[7221] = ~((inputs[687]) | (inputs[357]));
    assign layer0_outputs[7222] = (inputs[206]) & ~(inputs[11]);
    assign layer0_outputs[7223] = ~(inputs[554]);
    assign layer0_outputs[7224] = ~((inputs[645]) | (inputs[963]));
    assign layer0_outputs[7225] = (inputs[693]) | (inputs[242]);
    assign layer0_outputs[7226] = ~(inputs[861]);
    assign layer0_outputs[7227] = ~(inputs[195]);
    assign layer0_outputs[7228] = ~((inputs[893]) ^ (inputs[770]));
    assign layer0_outputs[7229] = (inputs[210]) | (inputs[48]);
    assign layer0_outputs[7230] = (inputs[841]) ^ (inputs[534]);
    assign layer0_outputs[7231] = (inputs[117]) ^ (inputs[922]);
    assign layer0_outputs[7232] = (inputs[221]) & (inputs[891]);
    assign layer0_outputs[7233] = (inputs[758]) ^ (inputs[328]);
    assign layer0_outputs[7234] = 1'b0;
    assign layer0_outputs[7235] = ~(inputs[829]) | (inputs[998]);
    assign layer0_outputs[7236] = (inputs[227]) ^ (inputs[499]);
    assign layer0_outputs[7237] = ~(inputs[685]);
    assign layer0_outputs[7238] = (inputs[410]) ^ (inputs[757]);
    assign layer0_outputs[7239] = (inputs[130]) | (inputs[327]);
    assign layer0_outputs[7240] = (inputs[649]) | (inputs[105]);
    assign layer0_outputs[7241] = (inputs[229]) | (inputs[293]);
    assign layer0_outputs[7242] = (inputs[805]) ^ (inputs[502]);
    assign layer0_outputs[7243] = (inputs[693]) ^ (inputs[769]);
    assign layer0_outputs[7244] = ~(inputs[693]) | (inputs[407]);
    assign layer0_outputs[7245] = ~((inputs[782]) | (inputs[761]));
    assign layer0_outputs[7246] = ~((inputs[34]) | (inputs[77]));
    assign layer0_outputs[7247] = (inputs[795]) & ~(inputs[893]);
    assign layer0_outputs[7248] = ~(inputs[731]);
    assign layer0_outputs[7249] = (inputs[640]) & ~(inputs[194]);
    assign layer0_outputs[7250] = ~(inputs[218]);
    assign layer0_outputs[7251] = ~((inputs[845]) | (inputs[39]));
    assign layer0_outputs[7252] = (inputs[216]) | (inputs[582]);
    assign layer0_outputs[7253] = ~((inputs[447]) & (inputs[18]));
    assign layer0_outputs[7254] = (inputs[603]) ^ (inputs[179]);
    assign layer0_outputs[7255] = (inputs[491]) ^ (inputs[160]);
    assign layer0_outputs[7256] = (inputs[864]) | (inputs[944]);
    assign layer0_outputs[7257] = (inputs[664]) & ~(inputs[928]);
    assign layer0_outputs[7258] = ~(inputs[607]) | (inputs[380]);
    assign layer0_outputs[7259] = (inputs[626]) & ~(inputs[922]);
    assign layer0_outputs[7260] = inputs[467];
    assign layer0_outputs[7261] = ~((inputs[50]) ^ (inputs[585]));
    assign layer0_outputs[7262] = (inputs[642]) ^ (inputs[195]);
    assign layer0_outputs[7263] = ~((inputs[512]) ^ (inputs[722]));
    assign layer0_outputs[7264] = ~(inputs[94]);
    assign layer0_outputs[7265] = ~((inputs[888]) ^ (inputs[910]));
    assign layer0_outputs[7266] = ~(inputs[461]);
    assign layer0_outputs[7267] = ~(inputs[211]) | (inputs[869]);
    assign layer0_outputs[7268] = ~(inputs[1003]) | (inputs[768]);
    assign layer0_outputs[7269] = (inputs[198]) | (inputs[818]);
    assign layer0_outputs[7270] = ~(inputs[550]);
    assign layer0_outputs[7271] = ~(inputs[280]) | (inputs[981]);
    assign layer0_outputs[7272] = ~(inputs[396]);
    assign layer0_outputs[7273] = (inputs[117]) ^ (inputs[781]);
    assign layer0_outputs[7274] = ~(inputs[314]) | (inputs[1004]);
    assign layer0_outputs[7275] = (inputs[552]) & ~(inputs[939]);
    assign layer0_outputs[7276] = ~(inputs[585]);
    assign layer0_outputs[7277] = (inputs[745]) & (inputs[352]);
    assign layer0_outputs[7278] = ~(inputs[927]);
    assign layer0_outputs[7279] = (inputs[298]) & ~(inputs[411]);
    assign layer0_outputs[7280] = (inputs[29]) | (inputs[58]);
    assign layer0_outputs[7281] = (inputs[915]) | (inputs[419]);
    assign layer0_outputs[7282] = ~((inputs[407]) ^ (inputs[139]));
    assign layer0_outputs[7283] = ~((inputs[846]) & (inputs[700]));
    assign layer0_outputs[7284] = (inputs[636]) | (inputs[744]);
    assign layer0_outputs[7285] = (inputs[898]) & ~(inputs[103]);
    assign layer0_outputs[7286] = (inputs[783]) ^ (inputs[761]);
    assign layer0_outputs[7287] = (inputs[419]) & ~(inputs[994]);
    assign layer0_outputs[7288] = ~(inputs[811]);
    assign layer0_outputs[7289] = (inputs[189]) & ~(inputs[451]);
    assign layer0_outputs[7290] = ~(inputs[717]);
    assign layer0_outputs[7291] = ~((inputs[239]) | (inputs[929]));
    assign layer0_outputs[7292] = (inputs[829]) ^ (inputs[1016]);
    assign layer0_outputs[7293] = (inputs[633]) & ~(inputs[456]);
    assign layer0_outputs[7294] = ~(inputs[253]) | (inputs[132]);
    assign layer0_outputs[7295] = ~(inputs[606]);
    assign layer0_outputs[7296] = ~((inputs[64]) ^ (inputs[1007]));
    assign layer0_outputs[7297] = (inputs[582]) & ~(inputs[898]);
    assign layer0_outputs[7298] = (inputs[561]) & ~(inputs[11]);
    assign layer0_outputs[7299] = ~(inputs[251]);
    assign layer0_outputs[7300] = ~(inputs[596]);
    assign layer0_outputs[7301] = ~((inputs[369]) & (inputs[593]));
    assign layer0_outputs[7302] = ~((inputs[549]) | (inputs[596]));
    assign layer0_outputs[7303] = inputs[9];
    assign layer0_outputs[7304] = ~(inputs[826]);
    assign layer0_outputs[7305] = ~((inputs[524]) ^ (inputs[533]));
    assign layer0_outputs[7306] = (inputs[408]) | (inputs[916]);
    assign layer0_outputs[7307] = ~(inputs[684]);
    assign layer0_outputs[7308] = (inputs[1011]) | (inputs[360]);
    assign layer0_outputs[7309] = inputs[424];
    assign layer0_outputs[7310] = ~((inputs[30]) | (inputs[582]));
    assign layer0_outputs[7311] = (inputs[354]) & (inputs[1020]);
    assign layer0_outputs[7312] = (inputs[692]) | (inputs[488]);
    assign layer0_outputs[7313] = inputs[774];
    assign layer0_outputs[7314] = (inputs[375]) ^ (inputs[311]);
    assign layer0_outputs[7315] = inputs[788];
    assign layer0_outputs[7316] = ~(inputs[552]);
    assign layer0_outputs[7317] = inputs[387];
    assign layer0_outputs[7318] = ~((inputs[734]) & (inputs[330]));
    assign layer0_outputs[7319] = (inputs[452]) & ~(inputs[193]);
    assign layer0_outputs[7320] = ~(inputs[303]);
    assign layer0_outputs[7321] = inputs[390];
    assign layer0_outputs[7322] = (inputs[295]) & ~(inputs[193]);
    assign layer0_outputs[7323] = inputs[467];
    assign layer0_outputs[7324] = ~(inputs[314]) | (inputs[552]);
    assign layer0_outputs[7325] = inputs[916];
    assign layer0_outputs[7326] = (inputs[734]) ^ (inputs[134]);
    assign layer0_outputs[7327] = inputs[255];
    assign layer0_outputs[7328] = (inputs[941]) | (inputs[271]);
    assign layer0_outputs[7329] = ~(inputs[425]);
    assign layer0_outputs[7330] = ~((inputs[837]) ^ (inputs[568]));
    assign layer0_outputs[7331] = (inputs[409]) ^ (inputs[862]);
    assign layer0_outputs[7332] = ~((inputs[516]) | (inputs[889]));
    assign layer0_outputs[7333] = (inputs[557]) ^ (inputs[835]);
    assign layer0_outputs[7334] = (inputs[182]) & (inputs[178]);
    assign layer0_outputs[7335] = (inputs[787]) & ~(inputs[547]);
    assign layer0_outputs[7336] = (inputs[740]) ^ (inputs[353]);
    assign layer0_outputs[7337] = ~(inputs[176]);
    assign layer0_outputs[7338] = inputs[183];
    assign layer0_outputs[7339] = ~((inputs[748]) | (inputs[644]));
    assign layer0_outputs[7340] = ~(inputs[2]) | (inputs[518]);
    assign layer0_outputs[7341] = (inputs[254]) | (inputs[522]);
    assign layer0_outputs[7342] = ~(inputs[456]) | (inputs[195]);
    assign layer0_outputs[7343] = ~((inputs[411]) | (inputs[778]));
    assign layer0_outputs[7344] = (inputs[997]) & ~(inputs[799]);
    assign layer0_outputs[7345] = ~(inputs[97]);
    assign layer0_outputs[7346] = (inputs[228]) ^ (inputs[685]);
    assign layer0_outputs[7347] = ~(inputs[819]) | (inputs[918]);
    assign layer0_outputs[7348] = (inputs[196]) | (inputs[111]);
    assign layer0_outputs[7349] = (inputs[33]) ^ (inputs[1002]);
    assign layer0_outputs[7350] = ~((inputs[188]) ^ (inputs[263]));
    assign layer0_outputs[7351] = ~((inputs[36]) & (inputs[275]));
    assign layer0_outputs[7352] = ~((inputs[58]) | (inputs[842]));
    assign layer0_outputs[7353] = (inputs[817]) | (inputs[798]);
    assign layer0_outputs[7354] = (inputs[526]) & ~(inputs[11]);
    assign layer0_outputs[7355] = ~(inputs[610]);
    assign layer0_outputs[7356] = (inputs[170]) | (inputs[364]);
    assign layer0_outputs[7357] = 1'b1;
    assign layer0_outputs[7358] = (inputs[464]) & ~(inputs[865]);
    assign layer0_outputs[7359] = (inputs[760]) & ~(inputs[618]);
    assign layer0_outputs[7360] = ~(inputs[47]) | (inputs[1007]);
    assign layer0_outputs[7361] = (inputs[943]) & ~(inputs[666]);
    assign layer0_outputs[7362] = (inputs[856]) ^ (inputs[1011]);
    assign layer0_outputs[7363] = (inputs[652]) | (inputs[759]);
    assign layer0_outputs[7364] = ~(inputs[924]) | (inputs[861]);
    assign layer0_outputs[7365] = ~(inputs[248]) | (inputs[58]);
    assign layer0_outputs[7366] = ~(inputs[715]);
    assign layer0_outputs[7367] = (inputs[462]) & ~(inputs[580]);
    assign layer0_outputs[7368] = ~(inputs[746]) | (inputs[978]);
    assign layer0_outputs[7369] = ~((inputs[677]) ^ (inputs[40]));
    assign layer0_outputs[7370] = (inputs[669]) & (inputs[292]);
    assign layer0_outputs[7371] = 1'b1;
    assign layer0_outputs[7372] = ~(inputs[500]);
    assign layer0_outputs[7373] = inputs[598];
    assign layer0_outputs[7374] = ~(inputs[926]) | (inputs[964]);
    assign layer0_outputs[7375] = (inputs[145]) & ~(inputs[838]);
    assign layer0_outputs[7376] = ~(inputs[595]) | (inputs[725]);
    assign layer0_outputs[7377] = (inputs[322]) & ~(inputs[164]);
    assign layer0_outputs[7378] = inputs[509];
    assign layer0_outputs[7379] = ~(inputs[113]);
    assign layer0_outputs[7380] = inputs[638];
    assign layer0_outputs[7381] = (inputs[494]) & ~(inputs[539]);
    assign layer0_outputs[7382] = inputs[222];
    assign layer0_outputs[7383] = (inputs[684]) & ~(inputs[297]);
    assign layer0_outputs[7384] = ~((inputs[864]) | (inputs[528]));
    assign layer0_outputs[7385] = ~(inputs[237]);
    assign layer0_outputs[7386] = ~((inputs[761]) ^ (inputs[820]));
    assign layer0_outputs[7387] = ~(inputs[455]);
    assign layer0_outputs[7388] = ~((inputs[612]) & (inputs[95]));
    assign layer0_outputs[7389] = (inputs[794]) ^ (inputs[231]);
    assign layer0_outputs[7390] = ~(inputs[682]) | (inputs[135]);
    assign layer0_outputs[7391] = (inputs[258]) ^ (inputs[592]);
    assign layer0_outputs[7392] = (inputs[855]) & ~(inputs[150]);
    assign layer0_outputs[7393] = ~((inputs[937]) | (inputs[412]));
    assign layer0_outputs[7394] = ~(inputs[680]);
    assign layer0_outputs[7395] = ~(inputs[52]);
    assign layer0_outputs[7396] = ~((inputs[712]) ^ (inputs[68]));
    assign layer0_outputs[7397] = ~(inputs[632]);
    assign layer0_outputs[7398] = ~(inputs[489]) | (inputs[543]);
    assign layer0_outputs[7399] = (inputs[830]) & ~(inputs[1014]);
    assign layer0_outputs[7400] = (inputs[655]) | (inputs[330]);
    assign layer0_outputs[7401] = (inputs[993]) & ~(inputs[62]);
    assign layer0_outputs[7402] = (inputs[439]) | (inputs[144]);
    assign layer0_outputs[7403] = (inputs[563]) | (inputs[804]);
    assign layer0_outputs[7404] = ~(inputs[547]);
    assign layer0_outputs[7405] = ~((inputs[134]) | (inputs[147]));
    assign layer0_outputs[7406] = inputs[73];
    assign layer0_outputs[7407] = ~(inputs[726]) | (inputs[219]);
    assign layer0_outputs[7408] = (inputs[318]) & ~(inputs[92]);
    assign layer0_outputs[7409] = ~(inputs[629]) | (inputs[282]);
    assign layer0_outputs[7410] = (inputs[451]) & ~(inputs[484]);
    assign layer0_outputs[7411] = (inputs[585]) & ~(inputs[23]);
    assign layer0_outputs[7412] = (inputs[828]) | (inputs[918]);
    assign layer0_outputs[7413] = (inputs[457]) ^ (inputs[582]);
    assign layer0_outputs[7414] = (inputs[407]) & ~(inputs[609]);
    assign layer0_outputs[7415] = (inputs[345]) | (inputs[135]);
    assign layer0_outputs[7416] = inputs[125];
    assign layer0_outputs[7417] = (inputs[1009]) | (inputs[782]);
    assign layer0_outputs[7418] = ~((inputs[952]) & (inputs[320]));
    assign layer0_outputs[7419] = ~((inputs[807]) & (inputs[1019]));
    assign layer0_outputs[7420] = ~((inputs[458]) | (inputs[687]));
    assign layer0_outputs[7421] = inputs[746];
    assign layer0_outputs[7422] = (inputs[840]) & ~(inputs[753]);
    assign layer0_outputs[7423] = inputs[362];
    assign layer0_outputs[7424] = ~(inputs[773]);
    assign layer0_outputs[7425] = ~(inputs[367]) | (inputs[864]);
    assign layer0_outputs[7426] = (inputs[779]) & ~(inputs[422]);
    assign layer0_outputs[7427] = ~(inputs[511]) | (inputs[156]);
    assign layer0_outputs[7428] = ~((inputs[831]) | (inputs[106]));
    assign layer0_outputs[7429] = ~(inputs[990]) | (inputs[195]);
    assign layer0_outputs[7430] = (inputs[187]) ^ (inputs[652]);
    assign layer0_outputs[7431] = (inputs[461]) & ~(inputs[803]);
    assign layer0_outputs[7432] = (inputs[151]) ^ (inputs[865]);
    assign layer0_outputs[7433] = ~(inputs[436]) | (inputs[82]);
    assign layer0_outputs[7434] = 1'b1;
    assign layer0_outputs[7435] = inputs[625];
    assign layer0_outputs[7436] = (inputs[293]) | (inputs[248]);
    assign layer0_outputs[7437] = ~((inputs[459]) ^ (inputs[29]));
    assign layer0_outputs[7438] = 1'b0;
    assign layer0_outputs[7439] = 1'b1;
    assign layer0_outputs[7440] = ~(inputs[61]);
    assign layer0_outputs[7441] = inputs[30];
    assign layer0_outputs[7442] = 1'b0;
    assign layer0_outputs[7443] = ~((inputs[336]) | (inputs[570]));
    assign layer0_outputs[7444] = ~((inputs[256]) | (inputs[470]));
    assign layer0_outputs[7445] = (inputs[923]) & ~(inputs[950]);
    assign layer0_outputs[7446] = ~((inputs[858]) ^ (inputs[306]));
    assign layer0_outputs[7447] = ~(inputs[532]) | (inputs[838]);
    assign layer0_outputs[7448] = inputs[652];
    assign layer0_outputs[7449] = (inputs[583]) | (inputs[651]);
    assign layer0_outputs[7450] = ~((inputs[87]) | (inputs[947]));
    assign layer0_outputs[7451] = ~(inputs[914]) | (inputs[793]);
    assign layer0_outputs[7452] = ~((inputs[581]) ^ (inputs[638]));
    assign layer0_outputs[7453] = ~(inputs[882]) | (inputs[825]);
    assign layer0_outputs[7454] = ~((inputs[876]) | (inputs[202]));
    assign layer0_outputs[7455] = (inputs[707]) ^ (inputs[202]);
    assign layer0_outputs[7456] = ~(inputs[212]) | (inputs[733]);
    assign layer0_outputs[7457] = (inputs[487]) & ~(inputs[751]);
    assign layer0_outputs[7458] = ~(inputs[117]);
    assign layer0_outputs[7459] = (inputs[804]) | (inputs[249]);
    assign layer0_outputs[7460] = ~(inputs[368]);
    assign layer0_outputs[7461] = ~(inputs[860]);
    assign layer0_outputs[7462] = ~(inputs[529]) | (inputs[110]);
    assign layer0_outputs[7463] = ~(inputs[532]) | (inputs[538]);
    assign layer0_outputs[7464] = 1'b0;
    assign layer0_outputs[7465] = ~(inputs[877]);
    assign layer0_outputs[7466] = (inputs[732]) | (inputs[143]);
    assign layer0_outputs[7467] = 1'b0;
    assign layer0_outputs[7468] = (inputs[689]) | (inputs[677]);
    assign layer0_outputs[7469] = (inputs[944]) ^ (inputs[159]);
    assign layer0_outputs[7470] = (inputs[643]) | (inputs[669]);
    assign layer0_outputs[7471] = (inputs[34]) & (inputs[156]);
    assign layer0_outputs[7472] = ~((inputs[206]) ^ (inputs[625]));
    assign layer0_outputs[7473] = ~((inputs[764]) & (inputs[972]));
    assign layer0_outputs[7474] = inputs[90];
    assign layer0_outputs[7475] = (inputs[307]) & ~(inputs[356]);
    assign layer0_outputs[7476] = ~(inputs[972]);
    assign layer0_outputs[7477] = ~((inputs[804]) ^ (inputs[1021]));
    assign layer0_outputs[7478] = ~(inputs[673]) | (inputs[677]);
    assign layer0_outputs[7479] = (inputs[348]) & ~(inputs[894]);
    assign layer0_outputs[7480] = (inputs[960]) | (inputs[536]);
    assign layer0_outputs[7481] = ~((inputs[191]) ^ (inputs[936]));
    assign layer0_outputs[7482] = inputs[239];
    assign layer0_outputs[7483] = ~((inputs[887]) | (inputs[707]));
    assign layer0_outputs[7484] = ~((inputs[474]) ^ (inputs[148]));
    assign layer0_outputs[7485] = ~(inputs[591]) | (inputs[793]);
    assign layer0_outputs[7486] = inputs[891];
    assign layer0_outputs[7487] = ~(inputs[848]);
    assign layer0_outputs[7488] = (inputs[356]) | (inputs[901]);
    assign layer0_outputs[7489] = ~(inputs[290]) | (inputs[589]);
    assign layer0_outputs[7490] = (inputs[4]) ^ (inputs[156]);
    assign layer0_outputs[7491] = inputs[827];
    assign layer0_outputs[7492] = inputs[943];
    assign layer0_outputs[7493] = ~((inputs[230]) ^ (inputs[463]));
    assign layer0_outputs[7494] = inputs[22];
    assign layer0_outputs[7495] = 1'b0;
    assign layer0_outputs[7496] = (inputs[51]) ^ (inputs[252]);
    assign layer0_outputs[7497] = (inputs[307]) & ~(inputs[388]);
    assign layer0_outputs[7498] = inputs[394];
    assign layer0_outputs[7499] = ~(inputs[389]);
    assign layer0_outputs[7500] = inputs[518];
    assign layer0_outputs[7501] = inputs[775];
    assign layer0_outputs[7502] = inputs[775];
    assign layer0_outputs[7503] = (inputs[818]) & ~(inputs[969]);
    assign layer0_outputs[7504] = ~(inputs[396]) | (inputs[938]);
    assign layer0_outputs[7505] = ~((inputs[248]) ^ (inputs[642]));
    assign layer0_outputs[7506] = ~((inputs[694]) | (inputs[601]));
    assign layer0_outputs[7507] = (inputs[893]) ^ (inputs[845]);
    assign layer0_outputs[7508] = (inputs[387]) & ~(inputs[932]);
    assign layer0_outputs[7509] = ~((inputs[500]) | (inputs[956]));
    assign layer0_outputs[7510] = (inputs[530]) & ~(inputs[207]);
    assign layer0_outputs[7511] = (inputs[675]) | (inputs[1010]);
    assign layer0_outputs[7512] = 1'b0;
    assign layer0_outputs[7513] = ~(inputs[527]) | (inputs[474]);
    assign layer0_outputs[7514] = (inputs[742]) | (inputs[755]);
    assign layer0_outputs[7515] = ~((inputs[459]) | (inputs[564]));
    assign layer0_outputs[7516] = ~(inputs[119]);
    assign layer0_outputs[7517] = ~(inputs[886]);
    assign layer0_outputs[7518] = ~(inputs[521]);
    assign layer0_outputs[7519] = (inputs[87]) ^ (inputs[984]);
    assign layer0_outputs[7520] = ~(inputs[540]) | (inputs[1017]);
    assign layer0_outputs[7521] = ~((inputs[308]) ^ (inputs[484]));
    assign layer0_outputs[7522] = ~(inputs[299]) | (inputs[43]);
    assign layer0_outputs[7523] = ~((inputs[543]) | (inputs[722]));
    assign layer0_outputs[7524] = (inputs[413]) & (inputs[239]);
    assign layer0_outputs[7525] = ~(inputs[601]) | (inputs[989]);
    assign layer0_outputs[7526] = (inputs[408]) & ~(inputs[83]);
    assign layer0_outputs[7527] = (inputs[190]) & (inputs[210]);
    assign layer0_outputs[7528] = ~((inputs[23]) ^ (inputs[565]));
    assign layer0_outputs[7529] = (inputs[104]) ^ (inputs[488]);
    assign layer0_outputs[7530] = inputs[598];
    assign layer0_outputs[7531] = ~((inputs[261]) | (inputs[490]));
    assign layer0_outputs[7532] = ~((inputs[178]) | (inputs[953]));
    assign layer0_outputs[7533] = inputs[879];
    assign layer0_outputs[7534] = ~((inputs[751]) ^ (inputs[1008]));
    assign layer0_outputs[7535] = ~(inputs[865]) | (inputs[977]);
    assign layer0_outputs[7536] = inputs[367];
    assign layer0_outputs[7537] = (inputs[427]) | (inputs[648]);
    assign layer0_outputs[7538] = (inputs[432]) ^ (inputs[866]);
    assign layer0_outputs[7539] = ~((inputs[691]) ^ (inputs[5]));
    assign layer0_outputs[7540] = (inputs[209]) ^ (inputs[49]);
    assign layer0_outputs[7541] = (inputs[263]) | (inputs[11]);
    assign layer0_outputs[7542] = ~((inputs[508]) & (inputs[802]));
    assign layer0_outputs[7543] = ~(inputs[658]) | (inputs[742]);
    assign layer0_outputs[7544] = (inputs[861]) & (inputs[482]);
    assign layer0_outputs[7545] = (inputs[836]) | (inputs[262]);
    assign layer0_outputs[7546] = inputs[464];
    assign layer0_outputs[7547] = (inputs[949]) & ~(inputs[604]);
    assign layer0_outputs[7548] = ~((inputs[733]) | (inputs[535]));
    assign layer0_outputs[7549] = (inputs[987]) & ~(inputs[609]);
    assign layer0_outputs[7550] = (inputs[115]) ^ (inputs[940]);
    assign layer0_outputs[7551] = ~(inputs[504]) | (inputs[927]);
    assign layer0_outputs[7552] = (inputs[129]) ^ (inputs[480]);
    assign layer0_outputs[7553] = (inputs[268]) ^ (inputs[360]);
    assign layer0_outputs[7554] = ~((inputs[261]) | (inputs[744]));
    assign layer0_outputs[7555] = ~((inputs[161]) & (inputs[187]));
    assign layer0_outputs[7556] = ~(inputs[558]) | (inputs[808]);
    assign layer0_outputs[7557] = ~(inputs[692]);
    assign layer0_outputs[7558] = ~(inputs[237]) | (inputs[154]);
    assign layer0_outputs[7559] = ~(inputs[317]) | (inputs[101]);
    assign layer0_outputs[7560] = (inputs[807]) ^ (inputs[958]);
    assign layer0_outputs[7561] = ~(inputs[945]) | (inputs[491]);
    assign layer0_outputs[7562] = ~((inputs[212]) | (inputs[637]));
    assign layer0_outputs[7563] = ~((inputs[348]) & (inputs[415]));
    assign layer0_outputs[7564] = ~((inputs[833]) | (inputs[586]));
    assign layer0_outputs[7565] = ~(inputs[518]) | (inputs[442]);
    assign layer0_outputs[7566] = (inputs[493]) & ~(inputs[948]);
    assign layer0_outputs[7567] = ~((inputs[738]) | (inputs[196]));
    assign layer0_outputs[7568] = ~((inputs[670]) ^ (inputs[259]));
    assign layer0_outputs[7569] = ~(inputs[858]);
    assign layer0_outputs[7570] = (inputs[403]) | (inputs[901]);
    assign layer0_outputs[7571] = (inputs[736]) ^ (inputs[445]);
    assign layer0_outputs[7572] = (inputs[446]) | (inputs[247]);
    assign layer0_outputs[7573] = ~((inputs[849]) & (inputs[898]));
    assign layer0_outputs[7574] = ~(inputs[142]) | (inputs[879]);
    assign layer0_outputs[7575] = (inputs[590]) & ~(inputs[870]);
    assign layer0_outputs[7576] = (inputs[957]) & ~(inputs[798]);
    assign layer0_outputs[7577] = (inputs[462]) & ~(inputs[321]);
    assign layer0_outputs[7578] = ~((inputs[671]) | (inputs[232]));
    assign layer0_outputs[7579] = (inputs[535]) | (inputs[470]);
    assign layer0_outputs[7580] = (inputs[919]) ^ (inputs[946]);
    assign layer0_outputs[7581] = (inputs[173]) & ~(inputs[969]);
    assign layer0_outputs[7582] = ~(inputs[951]);
    assign layer0_outputs[7583] = inputs[177];
    assign layer0_outputs[7584] = inputs[421];
    assign layer0_outputs[7585] = (inputs[339]) & ~(inputs[742]);
    assign layer0_outputs[7586] = (inputs[442]) & ~(inputs[986]);
    assign layer0_outputs[7587] = (inputs[774]) ^ (inputs[243]);
    assign layer0_outputs[7588] = ~((inputs[486]) ^ (inputs[238]));
    assign layer0_outputs[7589] = ~(inputs[463]);
    assign layer0_outputs[7590] = (inputs[658]) & (inputs[658]);
    assign layer0_outputs[7591] = inputs[576];
    assign layer0_outputs[7592] = (inputs[585]) ^ (inputs[995]);
    assign layer0_outputs[7593] = (inputs[12]) ^ (inputs[958]);
    assign layer0_outputs[7594] = (inputs[294]) & (inputs[639]);
    assign layer0_outputs[7595] = 1'b0;
    assign layer0_outputs[7596] = (inputs[277]) & ~(inputs[701]);
    assign layer0_outputs[7597] = inputs[373];
    assign layer0_outputs[7598] = (inputs[170]) | (inputs[212]);
    assign layer0_outputs[7599] = ~(inputs[220]) | (inputs[671]);
    assign layer0_outputs[7600] = 1'b0;
    assign layer0_outputs[7601] = ~(inputs[361]);
    assign layer0_outputs[7602] = ~((inputs[798]) | (inputs[424]));
    assign layer0_outputs[7603] = ~((inputs[277]) | (inputs[305]));
    assign layer0_outputs[7604] = (inputs[961]) | (inputs[816]);
    assign layer0_outputs[7605] = (inputs[324]) | (inputs[849]);
    assign layer0_outputs[7606] = (inputs[463]) | (inputs[738]);
    assign layer0_outputs[7607] = ~((inputs[465]) | (inputs[147]));
    assign layer0_outputs[7608] = inputs[210];
    assign layer0_outputs[7609] = inputs[747];
    assign layer0_outputs[7610] = ~(inputs[848]);
    assign layer0_outputs[7611] = ~(inputs[592]) | (inputs[469]);
    assign layer0_outputs[7612] = ~(inputs[477]);
    assign layer0_outputs[7613] = ~(inputs[236]);
    assign layer0_outputs[7614] = ~(inputs[811]);
    assign layer0_outputs[7615] = (inputs[165]) ^ (inputs[674]);
    assign layer0_outputs[7616] = ~(inputs[820]) | (inputs[25]);
    assign layer0_outputs[7617] = (inputs[343]) | (inputs[562]);
    assign layer0_outputs[7618] = ~((inputs[265]) | (inputs[289]));
    assign layer0_outputs[7619] = ~(inputs[494]) | (inputs[68]);
    assign layer0_outputs[7620] = ~(inputs[962]) | (inputs[57]);
    assign layer0_outputs[7621] = inputs[653];
    assign layer0_outputs[7622] = inputs[851];
    assign layer0_outputs[7623] = (inputs[915]) ^ (inputs[117]);
    assign layer0_outputs[7624] = ~(inputs[325]) | (inputs[35]);
    assign layer0_outputs[7625] = 1'b0;
    assign layer0_outputs[7626] = inputs[623];
    assign layer0_outputs[7627] = inputs[325];
    assign layer0_outputs[7628] = ~(inputs[797]);
    assign layer0_outputs[7629] = ~((inputs[21]) | (inputs[145]));
    assign layer0_outputs[7630] = inputs[886];
    assign layer0_outputs[7631] = ~(inputs[711]) | (inputs[518]);
    assign layer0_outputs[7632] = inputs[528];
    assign layer0_outputs[7633] = ~((inputs[1001]) | (inputs[526]));
    assign layer0_outputs[7634] = inputs[180];
    assign layer0_outputs[7635] = (inputs[606]) & ~(inputs[862]);
    assign layer0_outputs[7636] = ~(inputs[493]);
    assign layer0_outputs[7637] = (inputs[460]) ^ (inputs[210]);
    assign layer0_outputs[7638] = (inputs[536]) | (inputs[661]);
    assign layer0_outputs[7639] = (inputs[427]) & ~(inputs[721]);
    assign layer0_outputs[7640] = (inputs[597]) ^ (inputs[575]);
    assign layer0_outputs[7641] = ~(inputs[277]) | (inputs[495]);
    assign layer0_outputs[7642] = (inputs[552]) & ~(inputs[108]);
    assign layer0_outputs[7643] = (inputs[781]) & ~(inputs[983]);
    assign layer0_outputs[7644] = ~((inputs[898]) & (inputs[340]));
    assign layer0_outputs[7645] = ~(inputs[692]) | (inputs[580]);
    assign layer0_outputs[7646] = ~(inputs[897]) | (inputs[832]);
    assign layer0_outputs[7647] = ~(inputs[33]) | (inputs[966]);
    assign layer0_outputs[7648] = inputs[661];
    assign layer0_outputs[7649] = ~((inputs[453]) | (inputs[19]));
    assign layer0_outputs[7650] = ~((inputs[616]) ^ (inputs[624]));
    assign layer0_outputs[7651] = (inputs[251]) & ~(inputs[668]);
    assign layer0_outputs[7652] = (inputs[484]) ^ (inputs[956]);
    assign layer0_outputs[7653] = (inputs[889]) | (inputs[330]);
    assign layer0_outputs[7654] = ~((inputs[355]) ^ (inputs[809]));
    assign layer0_outputs[7655] = (inputs[849]) & ~(inputs[715]);
    assign layer0_outputs[7656] = ~((inputs[697]) & (inputs[675]));
    assign layer0_outputs[7657] = ~((inputs[525]) | (inputs[662]));
    assign layer0_outputs[7658] = ~((inputs[825]) | (inputs[590]));
    assign layer0_outputs[7659] = ~(inputs[111]) | (inputs[35]);
    assign layer0_outputs[7660] = ~((inputs[33]) | (inputs[588]));
    assign layer0_outputs[7661] = (inputs[446]) | (inputs[636]);
    assign layer0_outputs[7662] = (inputs[348]) | (inputs[205]);
    assign layer0_outputs[7663] = (inputs[201]) ^ (inputs[990]);
    assign layer0_outputs[7664] = (inputs[783]) ^ (inputs[845]);
    assign layer0_outputs[7665] = ~(inputs[1017]);
    assign layer0_outputs[7666] = ~((inputs[601]) | (inputs[483]));
    assign layer0_outputs[7667] = ~(inputs[624]);
    assign layer0_outputs[7668] = (inputs[872]) & ~(inputs[774]);
    assign layer0_outputs[7669] = inputs[394];
    assign layer0_outputs[7670] = inputs[648];
    assign layer0_outputs[7671] = (inputs[747]) & ~(inputs[96]);
    assign layer0_outputs[7672] = ~(inputs[510]);
    assign layer0_outputs[7673] = ~((inputs[390]) | (inputs[682]));
    assign layer0_outputs[7674] = 1'b1;
    assign layer0_outputs[7675] = ~(inputs[348]);
    assign layer0_outputs[7676] = (inputs[709]) | (inputs[761]);
    assign layer0_outputs[7677] = (inputs[845]) & ~(inputs[452]);
    assign layer0_outputs[7678] = (inputs[26]) & ~(inputs[232]);
    assign layer0_outputs[7679] = inputs[622];
    assign outputs[0] = (layer0_outputs[4064]) & ~(layer0_outputs[2045]);
    assign outputs[1] = ~(layer0_outputs[5137]);
    assign outputs[2] = ~(layer0_outputs[573]);
    assign outputs[3] = ~((layer0_outputs[6695]) & (layer0_outputs[5057]));
    assign outputs[4] = layer0_outputs[5378];
    assign outputs[5] = (layer0_outputs[5972]) ^ (layer0_outputs[7461]);
    assign outputs[6] = layer0_outputs[137];
    assign outputs[7] = layer0_outputs[392];
    assign outputs[8] = ~(layer0_outputs[7355]) | (layer0_outputs[1136]);
    assign outputs[9] = ~((layer0_outputs[6178]) & (layer0_outputs[3235]));
    assign outputs[10] = layer0_outputs[7080];
    assign outputs[11] = ~(layer0_outputs[5521]) | (layer0_outputs[3359]);
    assign outputs[12] = ~((layer0_outputs[5511]) ^ (layer0_outputs[3113]));
    assign outputs[13] = ~(layer0_outputs[4109]);
    assign outputs[14] = ~(layer0_outputs[5648]) | (layer0_outputs[4251]);
    assign outputs[15] = ~(layer0_outputs[3235]);
    assign outputs[16] = (layer0_outputs[3556]) | (layer0_outputs[4199]);
    assign outputs[17] = (layer0_outputs[7389]) ^ (layer0_outputs[3672]);
    assign outputs[18] = layer0_outputs[6589];
    assign outputs[19] = ~(layer0_outputs[3870]);
    assign outputs[20] = (layer0_outputs[1584]) ^ (layer0_outputs[3497]);
    assign outputs[21] = layer0_outputs[505];
    assign outputs[22] = ~(layer0_outputs[621]);
    assign outputs[23] = ~(layer0_outputs[5007]);
    assign outputs[24] = layer0_outputs[1302];
    assign outputs[25] = ~(layer0_outputs[5709]);
    assign outputs[26] = ~(layer0_outputs[189]) | (layer0_outputs[7587]);
    assign outputs[27] = ~((layer0_outputs[186]) ^ (layer0_outputs[5701]));
    assign outputs[28] = (layer0_outputs[2301]) & ~(layer0_outputs[7403]);
    assign outputs[29] = (layer0_outputs[6683]) & (layer0_outputs[6367]);
    assign outputs[30] = ~((layer0_outputs[254]) ^ (layer0_outputs[2642]));
    assign outputs[31] = ~(layer0_outputs[1388]) | (layer0_outputs[5488]);
    assign outputs[32] = (layer0_outputs[242]) ^ (layer0_outputs[3710]);
    assign outputs[33] = (layer0_outputs[3821]) ^ (layer0_outputs[1378]);
    assign outputs[34] = (layer0_outputs[3030]) & (layer0_outputs[5086]);
    assign outputs[35] = layer0_outputs[2910];
    assign outputs[36] = ~(layer0_outputs[7455]);
    assign outputs[37] = layer0_outputs[7411];
    assign outputs[38] = layer0_outputs[3384];
    assign outputs[39] = ~(layer0_outputs[913]);
    assign outputs[40] = ~(layer0_outputs[4204]);
    assign outputs[41] = (layer0_outputs[6603]) & ~(layer0_outputs[4658]);
    assign outputs[42] = ~(layer0_outputs[2307]);
    assign outputs[43] = ~(layer0_outputs[2248]);
    assign outputs[44] = ~(layer0_outputs[2714]);
    assign outputs[45] = ~(layer0_outputs[5240]) | (layer0_outputs[2617]);
    assign outputs[46] = ~(layer0_outputs[3399]);
    assign outputs[47] = ~((layer0_outputs[4904]) ^ (layer0_outputs[4567]));
    assign outputs[48] = (layer0_outputs[1758]) ^ (layer0_outputs[1506]);
    assign outputs[49] = ~(layer0_outputs[5226]) | (layer0_outputs[471]);
    assign outputs[50] = (layer0_outputs[2134]) & (layer0_outputs[7268]);
    assign outputs[51] = ~((layer0_outputs[6184]) | (layer0_outputs[718]));
    assign outputs[52] = ~(layer0_outputs[5761]);
    assign outputs[53] = layer0_outputs[1131];
    assign outputs[54] = ~((layer0_outputs[6760]) ^ (layer0_outputs[7545]));
    assign outputs[55] = (layer0_outputs[6471]) & ~(layer0_outputs[623]);
    assign outputs[56] = ~(layer0_outputs[2384]);
    assign outputs[57] = (layer0_outputs[553]) & (layer0_outputs[1972]);
    assign outputs[58] = (layer0_outputs[4257]) & (layer0_outputs[1314]);
    assign outputs[59] = ~(layer0_outputs[2316]) | (layer0_outputs[5710]);
    assign outputs[60] = ~((layer0_outputs[2209]) | (layer0_outputs[4767]));
    assign outputs[61] = (layer0_outputs[4100]) ^ (layer0_outputs[3134]);
    assign outputs[62] = (layer0_outputs[2072]) & (layer0_outputs[3487]);
    assign outputs[63] = ~((layer0_outputs[4689]) & (layer0_outputs[7553]));
    assign outputs[64] = ~(layer0_outputs[1021]) | (layer0_outputs[2801]);
    assign outputs[65] = ~(layer0_outputs[1373]);
    assign outputs[66] = ~(layer0_outputs[6441]);
    assign outputs[67] = layer0_outputs[1455];
    assign outputs[68] = layer0_outputs[6451];
    assign outputs[69] = (layer0_outputs[5447]) ^ (layer0_outputs[6963]);
    assign outputs[70] = (layer0_outputs[6839]) | (layer0_outputs[2951]);
    assign outputs[71] = ~(layer0_outputs[1165]);
    assign outputs[72] = ~(layer0_outputs[1495]);
    assign outputs[73] = layer0_outputs[4105];
    assign outputs[74] = (layer0_outputs[3041]) | (layer0_outputs[2767]);
    assign outputs[75] = ~(layer0_outputs[463]) | (layer0_outputs[560]);
    assign outputs[76] = ~((layer0_outputs[6032]) ^ (layer0_outputs[2825]));
    assign outputs[77] = ~((layer0_outputs[4210]) ^ (layer0_outputs[4831]));
    assign outputs[78] = layer0_outputs[3291];
    assign outputs[79] = ~((layer0_outputs[703]) ^ (layer0_outputs[5398]));
    assign outputs[80] = layer0_outputs[5962];
    assign outputs[81] = ~((layer0_outputs[3074]) ^ (layer0_outputs[5783]));
    assign outputs[82] = ~((layer0_outputs[1910]) ^ (layer0_outputs[704]));
    assign outputs[83] = ~(layer0_outputs[2400]) | (layer0_outputs[575]);
    assign outputs[84] = (layer0_outputs[2225]) ^ (layer0_outputs[3460]);
    assign outputs[85] = ~(layer0_outputs[5077]);
    assign outputs[86] = ~(layer0_outputs[2884]) | (layer0_outputs[4015]);
    assign outputs[87] = ~(layer0_outputs[1497]);
    assign outputs[88] = layer0_outputs[834];
    assign outputs[89] = (layer0_outputs[6447]) & ~(layer0_outputs[4401]);
    assign outputs[90] = (layer0_outputs[1027]) ^ (layer0_outputs[740]);
    assign outputs[91] = ~(layer0_outputs[2714]);
    assign outputs[92] = layer0_outputs[2912];
    assign outputs[93] = ~(layer0_outputs[3825]);
    assign outputs[94] = layer0_outputs[4236];
    assign outputs[95] = ~(layer0_outputs[466]);
    assign outputs[96] = 1'b1;
    assign outputs[97] = (layer0_outputs[4425]) ^ (layer0_outputs[5331]);
    assign outputs[98] = (layer0_outputs[7406]) ^ (layer0_outputs[4684]);
    assign outputs[99] = ~(layer0_outputs[3718]);
    assign outputs[100] = ~(layer0_outputs[6235]);
    assign outputs[101] = layer0_outputs[5133];
    assign outputs[102] = layer0_outputs[566];
    assign outputs[103] = ~((layer0_outputs[2643]) ^ (layer0_outputs[2965]));
    assign outputs[104] = ~(layer0_outputs[165]) | (layer0_outputs[3749]);
    assign outputs[105] = layer0_outputs[2179];
    assign outputs[106] = ~((layer0_outputs[7322]) | (layer0_outputs[6130]));
    assign outputs[107] = 1'b1;
    assign outputs[108] = ~(layer0_outputs[460]);
    assign outputs[109] = ~(layer0_outputs[2]);
    assign outputs[110] = (layer0_outputs[4970]) & (layer0_outputs[5993]);
    assign outputs[111] = ~(layer0_outputs[534]);
    assign outputs[112] = ~(layer0_outputs[3423]);
    assign outputs[113] = (layer0_outputs[2785]) ^ (layer0_outputs[6583]);
    assign outputs[114] = ~((layer0_outputs[6829]) ^ (layer0_outputs[4044]));
    assign outputs[115] = layer0_outputs[2450];
    assign outputs[116] = ~((layer0_outputs[5019]) ^ (layer0_outputs[6744]));
    assign outputs[117] = (layer0_outputs[98]) & (layer0_outputs[1619]);
    assign outputs[118] = layer0_outputs[2143];
    assign outputs[119] = (layer0_outputs[3372]) ^ (layer0_outputs[3029]);
    assign outputs[120] = ~(layer0_outputs[259]) | (layer0_outputs[6907]);
    assign outputs[121] = ~(layer0_outputs[6309]);
    assign outputs[122] = layer0_outputs[5037];
    assign outputs[123] = ~(layer0_outputs[1931]);
    assign outputs[124] = ~(layer0_outputs[1841]) | (layer0_outputs[2449]);
    assign outputs[125] = ~((layer0_outputs[3183]) ^ (layer0_outputs[4476]));
    assign outputs[126] = layer0_outputs[1206];
    assign outputs[127] = ~(layer0_outputs[5096]);
    assign outputs[128] = layer0_outputs[4252];
    assign outputs[129] = ~(layer0_outputs[467]);
    assign outputs[130] = layer0_outputs[1195];
    assign outputs[131] = ~(layer0_outputs[6063]);
    assign outputs[132] = (layer0_outputs[5053]) | (layer0_outputs[4038]);
    assign outputs[133] = ~(layer0_outputs[4510]);
    assign outputs[134] = layer0_outputs[4486];
    assign outputs[135] = ~(layer0_outputs[7200]) | (layer0_outputs[683]);
    assign outputs[136] = ~((layer0_outputs[6169]) ^ (layer0_outputs[7336]));
    assign outputs[137] = ~(layer0_outputs[3260]) | (layer0_outputs[4592]);
    assign outputs[138] = ~(layer0_outputs[6607]);
    assign outputs[139] = ~((layer0_outputs[4742]) ^ (layer0_outputs[1850]));
    assign outputs[140] = ~(layer0_outputs[6413]);
    assign outputs[141] = ~((layer0_outputs[4129]) ^ (layer0_outputs[5536]));
    assign outputs[142] = layer0_outputs[2438];
    assign outputs[143] = ~(layer0_outputs[1807]);
    assign outputs[144] = layer0_outputs[1879];
    assign outputs[145] = layer0_outputs[681];
    assign outputs[146] = layer0_outputs[1884];
    assign outputs[147] = layer0_outputs[6858];
    assign outputs[148] = layer0_outputs[2595];
    assign outputs[149] = ~(layer0_outputs[3408]);
    assign outputs[150] = ~((layer0_outputs[1070]) | (layer0_outputs[2223]));
    assign outputs[151] = layer0_outputs[7121];
    assign outputs[152] = layer0_outputs[5442];
    assign outputs[153] = layer0_outputs[2505];
    assign outputs[154] = layer0_outputs[6854];
    assign outputs[155] = (layer0_outputs[1134]) & ~(layer0_outputs[3176]);
    assign outputs[156] = (layer0_outputs[346]) ^ (layer0_outputs[2215]);
    assign outputs[157] = ~(layer0_outputs[5871]);
    assign outputs[158] = ~(layer0_outputs[4930]) | (layer0_outputs[632]);
    assign outputs[159] = layer0_outputs[7031];
    assign outputs[160] = ~((layer0_outputs[4900]) ^ (layer0_outputs[2980]));
    assign outputs[161] = layer0_outputs[608];
    assign outputs[162] = ~((layer0_outputs[2259]) ^ (layer0_outputs[4157]));
    assign outputs[163] = layer0_outputs[1041];
    assign outputs[164] = (layer0_outputs[3411]) & ~(layer0_outputs[7151]);
    assign outputs[165] = (layer0_outputs[2599]) | (layer0_outputs[3956]);
    assign outputs[166] = layer0_outputs[3829];
    assign outputs[167] = layer0_outputs[6853];
    assign outputs[168] = (layer0_outputs[4973]) ^ (layer0_outputs[1203]);
    assign outputs[169] = ~((layer0_outputs[767]) ^ (layer0_outputs[2799]));
    assign outputs[170] = (layer0_outputs[2056]) & ~(layer0_outputs[7010]);
    assign outputs[171] = ~(layer0_outputs[4958]) | (layer0_outputs[1115]);
    assign outputs[172] = ~(layer0_outputs[719]);
    assign outputs[173] = ~((layer0_outputs[3269]) | (layer0_outputs[2618]));
    assign outputs[174] = ~((layer0_outputs[2038]) | (layer0_outputs[4869]));
    assign outputs[175] = ~((layer0_outputs[4175]) ^ (layer0_outputs[2461]));
    assign outputs[176] = ~(layer0_outputs[1800]) | (layer0_outputs[1796]);
    assign outputs[177] = ~(layer0_outputs[6982]);
    assign outputs[178] = (layer0_outputs[135]) ^ (layer0_outputs[5387]);
    assign outputs[179] = ~(layer0_outputs[5375]) | (layer0_outputs[5305]);
    assign outputs[180] = layer0_outputs[748];
    assign outputs[181] = (layer0_outputs[6630]) ^ (layer0_outputs[2777]);
    assign outputs[182] = ~(layer0_outputs[108]);
    assign outputs[183] = (layer0_outputs[1118]) ^ (layer0_outputs[7332]);
    assign outputs[184] = (layer0_outputs[5295]) & ~(layer0_outputs[2782]);
    assign outputs[185] = ~(layer0_outputs[5662]);
    assign outputs[186] = (layer0_outputs[5242]) ^ (layer0_outputs[5612]);
    assign outputs[187] = layer0_outputs[3170];
    assign outputs[188] = ~((layer0_outputs[5269]) ^ (layer0_outputs[1500]));
    assign outputs[189] = layer0_outputs[771];
    assign outputs[190] = ~(layer0_outputs[4334]) | (layer0_outputs[1842]);
    assign outputs[191] = layer0_outputs[5451];
    assign outputs[192] = ~((layer0_outputs[5106]) ^ (layer0_outputs[109]));
    assign outputs[193] = ~(layer0_outputs[5880]);
    assign outputs[194] = ~((layer0_outputs[6867]) ^ (layer0_outputs[1442]));
    assign outputs[195] = (layer0_outputs[2112]) ^ (layer0_outputs[1671]);
    assign outputs[196] = ~((layer0_outputs[2367]) ^ (layer0_outputs[2096]));
    assign outputs[197] = layer0_outputs[322];
    assign outputs[198] = (layer0_outputs[2400]) ^ (layer0_outputs[1308]);
    assign outputs[199] = ~(layer0_outputs[2853]);
    assign outputs[200] = (layer0_outputs[4734]) ^ (layer0_outputs[2377]);
    assign outputs[201] = ~(layer0_outputs[4597]);
    assign outputs[202] = ~(layer0_outputs[6554]) | (layer0_outputs[815]);
    assign outputs[203] = ~((layer0_outputs[6102]) ^ (layer0_outputs[3941]));
    assign outputs[204] = ~(layer0_outputs[4088]);
    assign outputs[205] = ~(layer0_outputs[3804]) | (layer0_outputs[5801]);
    assign outputs[206] = ~(layer0_outputs[4239]) | (layer0_outputs[3521]);
    assign outputs[207] = layer0_outputs[1225];
    assign outputs[208] = ~(layer0_outputs[281]);
    assign outputs[209] = ~(layer0_outputs[2361]);
    assign outputs[210] = ~((layer0_outputs[6865]) ^ (layer0_outputs[6053]));
    assign outputs[211] = ~(layer0_outputs[6983]);
    assign outputs[212] = ~(layer0_outputs[3920]);
    assign outputs[213] = layer0_outputs[5037];
    assign outputs[214] = 1'b1;
    assign outputs[215] = layer0_outputs[4838];
    assign outputs[216] = (layer0_outputs[5967]) & (layer0_outputs[5411]);
    assign outputs[217] = 1'b1;
    assign outputs[218] = ~(layer0_outputs[757]);
    assign outputs[219] = (layer0_outputs[2336]) & ~(layer0_outputs[332]);
    assign outputs[220] = (layer0_outputs[142]) & (layer0_outputs[6171]);
    assign outputs[221] = ~(layer0_outputs[3207]);
    assign outputs[222] = (layer0_outputs[754]) ^ (layer0_outputs[6380]);
    assign outputs[223] = (layer0_outputs[6174]) & ~(layer0_outputs[2773]);
    assign outputs[224] = ~((layer0_outputs[4624]) ^ (layer0_outputs[4435]));
    assign outputs[225] = ~(layer0_outputs[606]);
    assign outputs[226] = layer0_outputs[256];
    assign outputs[227] = layer0_outputs[449];
    assign outputs[228] = ~(layer0_outputs[2682]);
    assign outputs[229] = ~(layer0_outputs[6827]);
    assign outputs[230] = layer0_outputs[5650];
    assign outputs[231] = (layer0_outputs[6894]) & (layer0_outputs[316]);
    assign outputs[232] = ~(layer0_outputs[1356]);
    assign outputs[233] = (layer0_outputs[507]) & ~(layer0_outputs[2924]);
    assign outputs[234] = ~(layer0_outputs[2329]) | (layer0_outputs[2468]);
    assign outputs[235] = layer0_outputs[5995];
    assign outputs[236] = layer0_outputs[3598];
    assign outputs[237] = layer0_outputs[7607];
    assign outputs[238] = ~(layer0_outputs[7108]);
    assign outputs[239] = (layer0_outputs[3450]) ^ (layer0_outputs[841]);
    assign outputs[240] = ~(layer0_outputs[6244]);
    assign outputs[241] = layer0_outputs[4905];
    assign outputs[242] = ~(layer0_outputs[7468]);
    assign outputs[243] = (layer0_outputs[6237]) & ~(layer0_outputs[494]);
    assign outputs[244] = ~(layer0_outputs[1754]);
    assign outputs[245] = ~((layer0_outputs[6141]) & (layer0_outputs[4570]));
    assign outputs[246] = ~(layer0_outputs[4398]);
    assign outputs[247] = layer0_outputs[4591];
    assign outputs[248] = (layer0_outputs[3149]) ^ (layer0_outputs[61]);
    assign outputs[249] = (layer0_outputs[6299]) ^ (layer0_outputs[2564]);
    assign outputs[250] = ~(layer0_outputs[2555]);
    assign outputs[251] = ~((layer0_outputs[3734]) ^ (layer0_outputs[7555]));
    assign outputs[252] = ~((layer0_outputs[6628]) & (layer0_outputs[5745]));
    assign outputs[253] = layer0_outputs[3587];
    assign outputs[254] = (layer0_outputs[994]) ^ (layer0_outputs[4034]);
    assign outputs[255] = ~(layer0_outputs[2191]);
    assign outputs[256] = 1'b1;
    assign outputs[257] = ~(layer0_outputs[7062]);
    assign outputs[258] = layer0_outputs[1465];
    assign outputs[259] = ~(layer0_outputs[6586]);
    assign outputs[260] = (layer0_outputs[4009]) & ~(layer0_outputs[5484]);
    assign outputs[261] = (layer0_outputs[5570]) ^ (layer0_outputs[44]);
    assign outputs[262] = ~(layer0_outputs[7358]);
    assign outputs[263] = layer0_outputs[5460];
    assign outputs[264] = ~(layer0_outputs[4258]);
    assign outputs[265] = layer0_outputs[4435];
    assign outputs[266] = (layer0_outputs[1228]) & (layer0_outputs[7529]);
    assign outputs[267] = layer0_outputs[6852];
    assign outputs[268] = (layer0_outputs[4644]) ^ (layer0_outputs[1306]);
    assign outputs[269] = layer0_outputs[7605];
    assign outputs[270] = (layer0_outputs[3866]) ^ (layer0_outputs[7224]);
    assign outputs[271] = ~(layer0_outputs[2672]);
    assign outputs[272] = layer0_outputs[3417];
    assign outputs[273] = (layer0_outputs[4839]) | (layer0_outputs[4128]);
    assign outputs[274] = (layer0_outputs[1516]) & ~(layer0_outputs[1378]);
    assign outputs[275] = layer0_outputs[898];
    assign outputs[276] = (layer0_outputs[6969]) | (layer0_outputs[7025]);
    assign outputs[277] = (layer0_outputs[5075]) | (layer0_outputs[5104]);
    assign outputs[278] = (layer0_outputs[6128]) & (layer0_outputs[2119]);
    assign outputs[279] = (layer0_outputs[2857]) | (layer0_outputs[7090]);
    assign outputs[280] = (layer0_outputs[618]) ^ (layer0_outputs[6723]);
    assign outputs[281] = ~((layer0_outputs[7623]) | (layer0_outputs[4325]));
    assign outputs[282] = layer0_outputs[3730];
    assign outputs[283] = ~(layer0_outputs[3955]);
    assign outputs[284] = 1'b1;
    assign outputs[285] = layer0_outputs[4866];
    assign outputs[286] = layer0_outputs[5659];
    assign outputs[287] = ~(layer0_outputs[5390]);
    assign outputs[288] = ~((layer0_outputs[5128]) & (layer0_outputs[3782]));
    assign outputs[289] = ~((layer0_outputs[3997]) ^ (layer0_outputs[4170]));
    assign outputs[290] = layer0_outputs[71];
    assign outputs[291] = ~(layer0_outputs[5941]);
    assign outputs[292] = layer0_outputs[3360];
    assign outputs[293] = layer0_outputs[2653];
    assign outputs[294] = layer0_outputs[5023];
    assign outputs[295] = (layer0_outputs[4222]) & ~(layer0_outputs[3802]);
    assign outputs[296] = (layer0_outputs[3444]) & ~(layer0_outputs[5393]);
    assign outputs[297] = ~(layer0_outputs[4429]);
    assign outputs[298] = (layer0_outputs[4857]) ^ (layer0_outputs[2217]);
    assign outputs[299] = ~((layer0_outputs[4201]) ^ (layer0_outputs[7066]));
    assign outputs[300] = (layer0_outputs[3784]) & ~(layer0_outputs[1917]);
    assign outputs[301] = ~((layer0_outputs[7173]) ^ (layer0_outputs[295]));
    assign outputs[302] = ~(layer0_outputs[5532]);
    assign outputs[303] = (layer0_outputs[6714]) & (layer0_outputs[4962]);
    assign outputs[304] = (layer0_outputs[338]) ^ (layer0_outputs[3377]);
    assign outputs[305] = layer0_outputs[4636];
    assign outputs[306] = (layer0_outputs[551]) ^ (layer0_outputs[7257]);
    assign outputs[307] = ~(layer0_outputs[5176]);
    assign outputs[308] = ~((layer0_outputs[7354]) ^ (layer0_outputs[985]));
    assign outputs[309] = layer0_outputs[4591];
    assign outputs[310] = ~(layer0_outputs[92]);
    assign outputs[311] = layer0_outputs[5199];
    assign outputs[312] = ~(layer0_outputs[6530]);
    assign outputs[313] = layer0_outputs[4572];
    assign outputs[314] = (layer0_outputs[4099]) ^ (layer0_outputs[7405]);
    assign outputs[315] = layer0_outputs[6367];
    assign outputs[316] = ~((layer0_outputs[3061]) & (layer0_outputs[5376]));
    assign outputs[317] = layer0_outputs[6047];
    assign outputs[318] = ~((layer0_outputs[5072]) | (layer0_outputs[6248]));
    assign outputs[319] = ~(layer0_outputs[6843]);
    assign outputs[320] = (layer0_outputs[4874]) & ~(layer0_outputs[1358]);
    assign outputs[321] = (layer0_outputs[216]) & ~(layer0_outputs[1951]);
    assign outputs[322] = layer0_outputs[7050];
    assign outputs[323] = (layer0_outputs[3823]) ^ (layer0_outputs[3135]);
    assign outputs[324] = ~((layer0_outputs[5195]) & (layer0_outputs[3562]));
    assign outputs[325] = ~((layer0_outputs[948]) ^ (layer0_outputs[1091]));
    assign outputs[326] = (layer0_outputs[6997]) ^ (layer0_outputs[2834]);
    assign outputs[327] = ~(layer0_outputs[286]);
    assign outputs[328] = ~(layer0_outputs[903]);
    assign outputs[329] = layer0_outputs[1514];
    assign outputs[330] = ~((layer0_outputs[4341]) ^ (layer0_outputs[2199]));
    assign outputs[331] = (layer0_outputs[1687]) ^ (layer0_outputs[7182]);
    assign outputs[332] = layer0_outputs[4222];
    assign outputs[333] = ~((layer0_outputs[3599]) ^ (layer0_outputs[3981]));
    assign outputs[334] = ~(layer0_outputs[1643]) | (layer0_outputs[1346]);
    assign outputs[335] = ~((layer0_outputs[7305]) ^ (layer0_outputs[2422]));
    assign outputs[336] = (layer0_outputs[6454]) & (layer0_outputs[6335]);
    assign outputs[337] = (layer0_outputs[381]) & ~(layer0_outputs[3676]);
    assign outputs[338] = ~(layer0_outputs[6107]);
    assign outputs[339] = (layer0_outputs[4072]) ^ (layer0_outputs[7115]);
    assign outputs[340] = layer0_outputs[3784];
    assign outputs[341] = ~((layer0_outputs[5416]) | (layer0_outputs[139]));
    assign outputs[342] = ~(layer0_outputs[4293]);
    assign outputs[343] = layer0_outputs[1535];
    assign outputs[344] = ~(layer0_outputs[5194]) | (layer0_outputs[6221]);
    assign outputs[345] = layer0_outputs[5160];
    assign outputs[346] = (layer0_outputs[2638]) & ~(layer0_outputs[6134]);
    assign outputs[347] = layer0_outputs[3627];
    assign outputs[348] = (layer0_outputs[5592]) ^ (layer0_outputs[7541]);
    assign outputs[349] = ~((layer0_outputs[6941]) | (layer0_outputs[3435]));
    assign outputs[350] = layer0_outputs[2055];
    assign outputs[351] = layer0_outputs[3583];
    assign outputs[352] = ~(layer0_outputs[6861]);
    assign outputs[353] = (layer0_outputs[214]) ^ (layer0_outputs[7370]);
    assign outputs[354] = ~(layer0_outputs[2683]);
    assign outputs[355] = (layer0_outputs[7055]) ^ (layer0_outputs[2757]);
    assign outputs[356] = ~(layer0_outputs[5508]);
    assign outputs[357] = ~(layer0_outputs[4647]);
    assign outputs[358] = layer0_outputs[2807];
    assign outputs[359] = layer0_outputs[500];
    assign outputs[360] = (layer0_outputs[4843]) & ~(layer0_outputs[355]);
    assign outputs[361] = layer0_outputs[3642];
    assign outputs[362] = layer0_outputs[2254];
    assign outputs[363] = ~((layer0_outputs[2547]) ^ (layer0_outputs[2131]));
    assign outputs[364] = layer0_outputs[4630];
    assign outputs[365] = ~(layer0_outputs[7577]);
    assign outputs[366] = ~((layer0_outputs[6481]) | (layer0_outputs[1893]));
    assign outputs[367] = ~(layer0_outputs[5559]);
    assign outputs[368] = layer0_outputs[4369];
    assign outputs[369] = ~(layer0_outputs[183]);
    assign outputs[370] = layer0_outputs[6897];
    assign outputs[371] = ~((layer0_outputs[2231]) ^ (layer0_outputs[3862]));
    assign outputs[372] = layer0_outputs[5939];
    assign outputs[373] = ~(layer0_outputs[729]);
    assign outputs[374] = (layer0_outputs[3424]) ^ (layer0_outputs[2129]);
    assign outputs[375] = (layer0_outputs[5079]) & ~(layer0_outputs[5250]);
    assign outputs[376] = (layer0_outputs[2297]) & ~(layer0_outputs[1284]);
    assign outputs[377] = ~((layer0_outputs[2817]) ^ (layer0_outputs[7274]));
    assign outputs[378] = ~((layer0_outputs[3101]) | (layer0_outputs[6512]));
    assign outputs[379] = ~(layer0_outputs[2808]);
    assign outputs[380] = ~((layer0_outputs[2022]) & (layer0_outputs[7290]));
    assign outputs[381] = (layer0_outputs[1055]) ^ (layer0_outputs[4569]);
    assign outputs[382] = ~((layer0_outputs[1268]) ^ (layer0_outputs[5927]));
    assign outputs[383] = (layer0_outputs[7566]) ^ (layer0_outputs[7476]);
    assign outputs[384] = ~((layer0_outputs[2454]) & (layer0_outputs[3616]));
    assign outputs[385] = layer0_outputs[6325];
    assign outputs[386] = layer0_outputs[6337];
    assign outputs[387] = (layer0_outputs[3515]) ^ (layer0_outputs[1661]);
    assign outputs[388] = layer0_outputs[1120];
    assign outputs[389] = (layer0_outputs[1966]) | (layer0_outputs[3746]);
    assign outputs[390] = ~((layer0_outputs[7323]) | (layer0_outputs[5200]));
    assign outputs[391] = ~((layer0_outputs[3105]) ^ (layer0_outputs[5616]));
    assign outputs[392] = layer0_outputs[1827];
    assign outputs[393] = ~(layer0_outputs[2040]) | (layer0_outputs[3397]);
    assign outputs[394] = ~(layer0_outputs[4986]);
    assign outputs[395] = layer0_outputs[4666];
    assign outputs[396] = ~((layer0_outputs[6432]) ^ (layer0_outputs[965]));
    assign outputs[397] = ~(layer0_outputs[2311]);
    assign outputs[398] = layer0_outputs[2083];
    assign outputs[399] = ~((layer0_outputs[5509]) & (layer0_outputs[3630]));
    assign outputs[400] = ~((layer0_outputs[7435]) | (layer0_outputs[4094]));
    assign outputs[401] = ~(layer0_outputs[2044]);
    assign outputs[402] = ~(layer0_outputs[627]);
    assign outputs[403] = (layer0_outputs[6573]) | (layer0_outputs[1370]);
    assign outputs[404] = ~((layer0_outputs[43]) ^ (layer0_outputs[997]));
    assign outputs[405] = (layer0_outputs[5218]) & ~(layer0_outputs[1283]);
    assign outputs[406] = (layer0_outputs[1355]) ^ (layer0_outputs[2366]);
    assign outputs[407] = ~(layer0_outputs[6631]);
    assign outputs[408] = (layer0_outputs[4756]) & ~(layer0_outputs[7054]);
    assign outputs[409] = layer0_outputs[3291];
    assign outputs[410] = ~((layer0_outputs[3738]) ^ (layer0_outputs[4247]));
    assign outputs[411] = (layer0_outputs[2649]) ^ (layer0_outputs[540]);
    assign outputs[412] = layer0_outputs[7542];
    assign outputs[413] = ~(layer0_outputs[1640]);
    assign outputs[414] = (layer0_outputs[3615]) ^ (layer0_outputs[7155]);
    assign outputs[415] = (layer0_outputs[4615]) & ~(layer0_outputs[278]);
    assign outputs[416] = layer0_outputs[3791];
    assign outputs[417] = ~(layer0_outputs[1709]);
    assign outputs[418] = (layer0_outputs[1025]) & ~(layer0_outputs[6476]);
    assign outputs[419] = layer0_outputs[6875];
    assign outputs[420] = ~((layer0_outputs[6632]) ^ (layer0_outputs[4588]));
    assign outputs[421] = ~((layer0_outputs[6791]) ^ (layer0_outputs[5536]));
    assign outputs[422] = ~((layer0_outputs[1329]) & (layer0_outputs[6149]));
    assign outputs[423] = (layer0_outputs[4150]) & ~(layer0_outputs[3897]);
    assign outputs[424] = ~(layer0_outputs[1548]);
    assign outputs[425] = ~(layer0_outputs[4339]);
    assign outputs[426] = ~(layer0_outputs[6438]);
    assign outputs[427] = ~(layer0_outputs[6891]);
    assign outputs[428] = ~(layer0_outputs[5694]);
    assign outputs[429] = layer0_outputs[415];
    assign outputs[430] = ~(layer0_outputs[526]);
    assign outputs[431] = ~(layer0_outputs[1716]) | (layer0_outputs[1900]);
    assign outputs[432] = ~((layer0_outputs[7123]) ^ (layer0_outputs[7593]));
    assign outputs[433] = ~(layer0_outputs[1736]);
    assign outputs[434] = layer0_outputs[7045];
    assign outputs[435] = layer0_outputs[1869];
    assign outputs[436] = ~(layer0_outputs[3187]);
    assign outputs[437] = ~(layer0_outputs[7653]) | (layer0_outputs[1319]);
    assign outputs[438] = ~(layer0_outputs[5322]);
    assign outputs[439] = ~(layer0_outputs[262]);
    assign outputs[440] = ~(layer0_outputs[4922]) | (layer0_outputs[1376]);
    assign outputs[441] = layer0_outputs[458];
    assign outputs[442] = (layer0_outputs[2069]) | (layer0_outputs[7084]);
    assign outputs[443] = ~(layer0_outputs[4370]);
    assign outputs[444] = ~((layer0_outputs[6153]) ^ (layer0_outputs[1768]));
    assign outputs[445] = ~(layer0_outputs[2542]) | (layer0_outputs[2313]);
    assign outputs[446] = layer0_outputs[6526];
    assign outputs[447] = ~(layer0_outputs[6350]);
    assign outputs[448] = layer0_outputs[6422];
    assign outputs[449] = ~(layer0_outputs[1357]) | (layer0_outputs[3811]);
    assign outputs[450] = (layer0_outputs[4034]) | (layer0_outputs[4871]);
    assign outputs[451] = ~((layer0_outputs[2681]) & (layer0_outputs[5885]));
    assign outputs[452] = (layer0_outputs[2395]) | (layer0_outputs[970]);
    assign outputs[453] = (layer0_outputs[3555]) ^ (layer0_outputs[6812]);
    assign outputs[454] = (layer0_outputs[1878]) & ~(layer0_outputs[684]);
    assign outputs[455] = ~((layer0_outputs[4336]) & (layer0_outputs[6090]));
    assign outputs[456] = (layer0_outputs[4152]) ^ (layer0_outputs[4940]);
    assign outputs[457] = (layer0_outputs[1105]) & ~(layer0_outputs[4975]);
    assign outputs[458] = (layer0_outputs[7232]) ^ (layer0_outputs[312]);
    assign outputs[459] = ~(layer0_outputs[1527]);
    assign outputs[460] = ~((layer0_outputs[5522]) | (layer0_outputs[3882]));
    assign outputs[461] = (layer0_outputs[5618]) & ~(layer0_outputs[6755]);
    assign outputs[462] = ~((layer0_outputs[2876]) ^ (layer0_outputs[5440]));
    assign outputs[463] = ~((layer0_outputs[2831]) ^ (layer0_outputs[2078]));
    assign outputs[464] = ~(layer0_outputs[6889]);
    assign outputs[465] = layer0_outputs[5316];
    assign outputs[466] = ~((layer0_outputs[5686]) | (layer0_outputs[3011]));
    assign outputs[467] = layer0_outputs[793];
    assign outputs[468] = (layer0_outputs[2383]) | (layer0_outputs[4579]);
    assign outputs[469] = (layer0_outputs[7539]) ^ (layer0_outputs[6259]);
    assign outputs[470] = ~(layer0_outputs[570]);
    assign outputs[471] = layer0_outputs[7677];
    assign outputs[472] = ~(layer0_outputs[1903]) | (layer0_outputs[5926]);
    assign outputs[473] = ~(layer0_outputs[5647]) | (layer0_outputs[4595]);
    assign outputs[474] = ~((layer0_outputs[5867]) | (layer0_outputs[7220]));
    assign outputs[475] = ~((layer0_outputs[7188]) & (layer0_outputs[4342]));
    assign outputs[476] = (layer0_outputs[3105]) & ~(layer0_outputs[7002]);
    assign outputs[477] = ~(layer0_outputs[3533]);
    assign outputs[478] = layer0_outputs[1023];
    assign outputs[479] = ~(layer0_outputs[2469]) | (layer0_outputs[4520]);
    assign outputs[480] = ~(layer0_outputs[2765]);
    assign outputs[481] = layer0_outputs[1184];
    assign outputs[482] = ~(layer0_outputs[1417]);
    assign outputs[483] = (layer0_outputs[6682]) & ~(layer0_outputs[7081]);
    assign outputs[484] = ~(layer0_outputs[2356]);
    assign outputs[485] = layer0_outputs[911];
    assign outputs[486] = ~((layer0_outputs[660]) ^ (layer0_outputs[6743]));
    assign outputs[487] = (layer0_outputs[5014]) & (layer0_outputs[6903]);
    assign outputs[488] = (layer0_outputs[5596]) & ~(layer0_outputs[5664]);
    assign outputs[489] = ~(layer0_outputs[5163]);
    assign outputs[490] = ~(layer0_outputs[5519]);
    assign outputs[491] = (layer0_outputs[6722]) & ~(layer0_outputs[7099]);
    assign outputs[492] = ~(layer0_outputs[356]) | (layer0_outputs[5419]);
    assign outputs[493] = layer0_outputs[6785];
    assign outputs[494] = ~((layer0_outputs[4069]) & (layer0_outputs[2354]));
    assign outputs[495] = (layer0_outputs[2188]) ^ (layer0_outputs[4229]);
    assign outputs[496] = (layer0_outputs[6940]) & ~(layer0_outputs[1316]);
    assign outputs[497] = ~(layer0_outputs[1795]);
    assign outputs[498] = ~(layer0_outputs[1780]);
    assign outputs[499] = layer0_outputs[1840];
    assign outputs[500] = ~(layer0_outputs[2698]);
    assign outputs[501] = ~(layer0_outputs[990]);
    assign outputs[502] = ~((layer0_outputs[1669]) | (layer0_outputs[6771]));
    assign outputs[503] = ~((layer0_outputs[4724]) & (layer0_outputs[3836]));
    assign outputs[504] = ~(layer0_outputs[1264]);
    assign outputs[505] = layer0_outputs[6774];
    assign outputs[506] = (layer0_outputs[3490]) & ~(layer0_outputs[995]);
    assign outputs[507] = (layer0_outputs[1505]) ^ (layer0_outputs[6245]);
    assign outputs[508] = (layer0_outputs[6294]) & (layer0_outputs[5950]);
    assign outputs[509] = layer0_outputs[722];
    assign outputs[510] = layer0_outputs[6669];
    assign outputs[511] = (layer0_outputs[2711]) ^ (layer0_outputs[1056]);
    assign outputs[512] = (layer0_outputs[5627]) & ~(layer0_outputs[204]);
    assign outputs[513] = layer0_outputs[3997];
    assign outputs[514] = (layer0_outputs[5604]) & ~(layer0_outputs[7615]);
    assign outputs[515] = layer0_outputs[7596];
    assign outputs[516] = 1'b0;
    assign outputs[517] = layer0_outputs[632];
    assign outputs[518] = layer0_outputs[2802];
    assign outputs[519] = (layer0_outputs[4396]) & ~(layer0_outputs[7330]);
    assign outputs[520] = ~(layer0_outputs[1410]);
    assign outputs[521] = layer0_outputs[1296];
    assign outputs[522] = ~((layer0_outputs[3434]) ^ (layer0_outputs[3670]));
    assign outputs[523] = (layer0_outputs[5260]) ^ (layer0_outputs[1215]);
    assign outputs[524] = ~((layer0_outputs[4806]) ^ (layer0_outputs[4196]));
    assign outputs[525] = (layer0_outputs[307]) ^ (layer0_outputs[6704]);
    assign outputs[526] = ~(layer0_outputs[5215]);
    assign outputs[527] = layer0_outputs[5678];
    assign outputs[528] = layer0_outputs[2778];
    assign outputs[529] = layer0_outputs[5823];
    assign outputs[530] = layer0_outputs[5581];
    assign outputs[531] = (layer0_outputs[4496]) | (layer0_outputs[1715]);
    assign outputs[532] = ~(layer0_outputs[5393]);
    assign outputs[533] = ~(layer0_outputs[4258]);
    assign outputs[534] = ~(layer0_outputs[5213]) | (layer0_outputs[6698]);
    assign outputs[535] = (layer0_outputs[2779]) | (layer0_outputs[657]);
    assign outputs[536] = ~(layer0_outputs[1447]);
    assign outputs[537] = ~(layer0_outputs[6433]);
    assign outputs[538] = ~((layer0_outputs[7563]) ^ (layer0_outputs[2312]));
    assign outputs[539] = ~((layer0_outputs[1452]) & (layer0_outputs[6735]));
    assign outputs[540] = ~((layer0_outputs[2130]) ^ (layer0_outputs[2955]));
    assign outputs[541] = layer0_outputs[3751];
    assign outputs[542] = ~((layer0_outputs[2541]) ^ (layer0_outputs[2960]));
    assign outputs[543] = layer0_outputs[7497];
    assign outputs[544] = (layer0_outputs[5733]) & ~(layer0_outputs[490]);
    assign outputs[545] = ~(layer0_outputs[6193]) | (layer0_outputs[3243]);
    assign outputs[546] = (layer0_outputs[2869]) & (layer0_outputs[6029]);
    assign outputs[547] = ~(layer0_outputs[127]);
    assign outputs[548] = layer0_outputs[2858];
    assign outputs[549] = layer0_outputs[7132];
    assign outputs[550] = (layer0_outputs[4424]) ^ (layer0_outputs[6675]);
    assign outputs[551] = layer0_outputs[4256];
    assign outputs[552] = layer0_outputs[1535];
    assign outputs[553] = (layer0_outputs[4347]) & ~(layer0_outputs[2538]);
    assign outputs[554] = layer0_outputs[636];
    assign outputs[555] = layer0_outputs[4776];
    assign outputs[556] = (layer0_outputs[640]) ^ (layer0_outputs[4156]);
    assign outputs[557] = ~((layer0_outputs[3805]) ^ (layer0_outputs[3903]));
    assign outputs[558] = layer0_outputs[5629];
    assign outputs[559] = layer0_outputs[5438];
    assign outputs[560] = (layer0_outputs[1719]) & ~(layer0_outputs[2428]);
    assign outputs[561] = layer0_outputs[4559];
    assign outputs[562] = ~(layer0_outputs[6104]);
    assign outputs[563] = ~(layer0_outputs[4219]) | (layer0_outputs[5876]);
    assign outputs[564] = ~((layer0_outputs[1935]) & (layer0_outputs[1290]));
    assign outputs[565] = ~(layer0_outputs[4790]) | (layer0_outputs[6331]);
    assign outputs[566] = ~(layer0_outputs[4204]);
    assign outputs[567] = ~(layer0_outputs[3789]) | (layer0_outputs[3475]);
    assign outputs[568] = (layer0_outputs[3613]) ^ (layer0_outputs[6018]);
    assign outputs[569] = ~(layer0_outputs[6889]);
    assign outputs[570] = (layer0_outputs[4594]) & (layer0_outputs[6980]);
    assign outputs[571] = layer0_outputs[2920];
    assign outputs[572] = ~((layer0_outputs[1933]) ^ (layer0_outputs[2197]));
    assign outputs[573] = ~(layer0_outputs[2139]) | (layer0_outputs[1967]);
    assign outputs[574] = layer0_outputs[1847];
    assign outputs[575] = ~((layer0_outputs[1909]) ^ (layer0_outputs[5385]));
    assign outputs[576] = layer0_outputs[1714];
    assign outputs[577] = ~(layer0_outputs[2575]);
    assign outputs[578] = layer0_outputs[7421];
    assign outputs[579] = layer0_outputs[672];
    assign outputs[580] = ~(layer0_outputs[4346]);
    assign outputs[581] = (layer0_outputs[2676]) ^ (layer0_outputs[4001]);
    assign outputs[582] = layer0_outputs[6459];
    assign outputs[583] = ~(layer0_outputs[3868]);
    assign outputs[584] = ~(layer0_outputs[1437]);
    assign outputs[585] = ~((layer0_outputs[6668]) & (layer0_outputs[4500]));
    assign outputs[586] = (layer0_outputs[466]) ^ (layer0_outputs[6819]);
    assign outputs[587] = (layer0_outputs[6102]) ^ (layer0_outputs[2101]);
    assign outputs[588] = layer0_outputs[6805];
    assign outputs[589] = 1'b1;
    assign outputs[590] = ~((layer0_outputs[5715]) ^ (layer0_outputs[2472]));
    assign outputs[591] = ~((layer0_outputs[538]) ^ (layer0_outputs[3498]));
    assign outputs[592] = ~((layer0_outputs[634]) ^ (layer0_outputs[6479]));
    assign outputs[593] = layer0_outputs[4477];
    assign outputs[594] = layer0_outputs[1255];
    assign outputs[595] = layer0_outputs[159];
    assign outputs[596] = layer0_outputs[1089];
    assign outputs[597] = ~(layer0_outputs[1349]);
    assign outputs[598] = ~((layer0_outputs[1259]) ^ (layer0_outputs[1809]));
    assign outputs[599] = ~(layer0_outputs[1898]);
    assign outputs[600] = ~(layer0_outputs[1410]);
    assign outputs[601] = layer0_outputs[6845];
    assign outputs[602] = ~((layer0_outputs[2998]) ^ (layer0_outputs[2195]));
    assign outputs[603] = ~((layer0_outputs[1595]) & (layer0_outputs[6820]));
    assign outputs[604] = ~(layer0_outputs[3617]) | (layer0_outputs[620]);
    assign outputs[605] = (layer0_outputs[5363]) | (layer0_outputs[4553]);
    assign outputs[606] = ~(layer0_outputs[6203]);
    assign outputs[607] = layer0_outputs[6254];
    assign outputs[608] = layer0_outputs[6303];
    assign outputs[609] = ~(layer0_outputs[2553]);
    assign outputs[610] = ~(layer0_outputs[4929]);
    assign outputs[611] = ~(layer0_outputs[1876]) | (layer0_outputs[567]);
    assign outputs[612] = layer0_outputs[2552];
    assign outputs[613] = ~((layer0_outputs[3296]) | (layer0_outputs[1757]));
    assign outputs[614] = ~(layer0_outputs[2766]);
    assign outputs[615] = ~((layer0_outputs[3493]) ^ (layer0_outputs[4702]));
    assign outputs[616] = ~(layer0_outputs[4709]);
    assign outputs[617] = (layer0_outputs[4717]) ^ (layer0_outputs[6908]);
    assign outputs[618] = ~(layer0_outputs[6837]);
    assign outputs[619] = ~(layer0_outputs[6757]) | (layer0_outputs[203]);
    assign outputs[620] = ~((layer0_outputs[5414]) ^ (layer0_outputs[1266]));
    assign outputs[621] = layer0_outputs[5815];
    assign outputs[622] = (layer0_outputs[6952]) & ~(layer0_outputs[6450]);
    assign outputs[623] = ~(layer0_outputs[515]);
    assign outputs[624] = layer0_outputs[2742];
    assign outputs[625] = ~(layer0_outputs[7068]);
    assign outputs[626] = ~(layer0_outputs[5997]);
    assign outputs[627] = ~(layer0_outputs[6201]);
    assign outputs[628] = layer0_outputs[1665];
    assign outputs[629] = ~((layer0_outputs[4162]) ^ (layer0_outputs[729]));
    assign outputs[630] = (layer0_outputs[6073]) ^ (layer0_outputs[2115]);
    assign outputs[631] = layer0_outputs[2450];
    assign outputs[632] = ~(layer0_outputs[3539]);
    assign outputs[633] = (layer0_outputs[1713]) | (layer0_outputs[2789]);
    assign outputs[634] = ~((layer0_outputs[2019]) ^ (layer0_outputs[5715]));
    assign outputs[635] = (layer0_outputs[5958]) & ~(layer0_outputs[4480]);
    assign outputs[636] = (layer0_outputs[6003]) ^ (layer0_outputs[4017]);
    assign outputs[637] = layer0_outputs[3418];
    assign outputs[638] = (layer0_outputs[5817]) & ~(layer0_outputs[5165]);
    assign outputs[639] = ~(layer0_outputs[7343]);
    assign outputs[640] = ~((layer0_outputs[6514]) ^ (layer0_outputs[5465]));
    assign outputs[641] = layer0_outputs[6718];
    assign outputs[642] = (layer0_outputs[7493]) ^ (layer0_outputs[2342]);
    assign outputs[643] = layer0_outputs[677];
    assign outputs[644] = layer0_outputs[5690];
    assign outputs[645] = layer0_outputs[3890];
    assign outputs[646] = (layer0_outputs[3177]) & (layer0_outputs[959]);
    assign outputs[647] = ~(layer0_outputs[1247]) | (layer0_outputs[3962]);
    assign outputs[648] = ~(layer0_outputs[4510]);
    assign outputs[649] = ~(layer0_outputs[4607]);
    assign outputs[650] = ~(layer0_outputs[2316]);
    assign outputs[651] = layer0_outputs[765];
    assign outputs[652] = ~(layer0_outputs[4692]);
    assign outputs[653] = ~(layer0_outputs[7443]) | (layer0_outputs[3957]);
    assign outputs[654] = ~(layer0_outputs[908]);
    assign outputs[655] = (layer0_outputs[6712]) | (layer0_outputs[4499]);
    assign outputs[656] = (layer0_outputs[3239]) & (layer0_outputs[322]);
    assign outputs[657] = ~((layer0_outputs[7307]) ^ (layer0_outputs[5677]));
    assign outputs[658] = layer0_outputs[2755];
    assign outputs[659] = layer0_outputs[6498];
    assign outputs[660] = ~(layer0_outputs[3275]) | (layer0_outputs[6951]);
    assign outputs[661] = (layer0_outputs[5482]) ^ (layer0_outputs[6382]);
    assign outputs[662] = ~((layer0_outputs[4908]) ^ (layer0_outputs[1366]));
    assign outputs[663] = ~((layer0_outputs[2043]) ^ (layer0_outputs[241]));
    assign outputs[664] = layer0_outputs[1774];
    assign outputs[665] = ~(layer0_outputs[3366]);
    assign outputs[666] = ~(layer0_outputs[4470]);
    assign outputs[667] = (layer0_outputs[4107]) ^ (layer0_outputs[5121]);
    assign outputs[668] = layer0_outputs[4471];
    assign outputs[669] = ~((layer0_outputs[4750]) ^ (layer0_outputs[1470]));
    assign outputs[670] = (layer0_outputs[6689]) ^ (layer0_outputs[3941]);
    assign outputs[671] = ~((layer0_outputs[2501]) ^ (layer0_outputs[7618]));
    assign outputs[672] = (layer0_outputs[3517]) & ~(layer0_outputs[5557]);
    assign outputs[673] = (layer0_outputs[2844]) ^ (layer0_outputs[2733]);
    assign outputs[674] = ~(layer0_outputs[3944]) | (layer0_outputs[1453]);
    assign outputs[675] = layer0_outputs[3450];
    assign outputs[676] = layer0_outputs[47];
    assign outputs[677] = ~((layer0_outputs[3646]) ^ (layer0_outputs[738]));
    assign outputs[678] = ~((layer0_outputs[1043]) ^ (layer0_outputs[4966]));
    assign outputs[679] = layer0_outputs[1414];
    assign outputs[680] = layer0_outputs[102];
    assign outputs[681] = ~(layer0_outputs[6637]);
    assign outputs[682] = ~(layer0_outputs[6517]);
    assign outputs[683] = ~((layer0_outputs[2436]) ^ (layer0_outputs[6638]));
    assign outputs[684] = ~(layer0_outputs[1991]);
    assign outputs[685] = (layer0_outputs[6439]) ^ (layer0_outputs[4976]);
    assign outputs[686] = ~((layer0_outputs[492]) ^ (layer0_outputs[6767]));
    assign outputs[687] = ~((layer0_outputs[4390]) | (layer0_outputs[7623]));
    assign outputs[688] = layer0_outputs[932];
    assign outputs[689] = (layer0_outputs[3142]) ^ (layer0_outputs[7474]);
    assign outputs[690] = ~((layer0_outputs[5222]) ^ (layer0_outputs[6422]));
    assign outputs[691] = layer0_outputs[482];
    assign outputs[692] = ~((layer0_outputs[1537]) ^ (layer0_outputs[298]));
    assign outputs[693] = ~((layer0_outputs[4018]) & (layer0_outputs[2608]));
    assign outputs[694] = layer0_outputs[3007];
    assign outputs[695] = ~(layer0_outputs[1069]) | (layer0_outputs[1582]);
    assign outputs[696] = (layer0_outputs[5065]) & ~(layer0_outputs[4320]);
    assign outputs[697] = ~(layer0_outputs[4955]);
    assign outputs[698] = ~(layer0_outputs[2097]) | (layer0_outputs[3798]);
    assign outputs[699] = layer0_outputs[2872];
    assign outputs[700] = layer0_outputs[130];
    assign outputs[701] = layer0_outputs[7526];
    assign outputs[702] = ~(layer0_outputs[305]);
    assign outputs[703] = (layer0_outputs[3790]) ^ (layer0_outputs[5982]);
    assign outputs[704] = layer0_outputs[1412];
    assign outputs[705] = ~(layer0_outputs[6872]) | (layer0_outputs[1670]);
    assign outputs[706] = ~((layer0_outputs[4529]) | (layer0_outputs[1793]));
    assign outputs[707] = ~((layer0_outputs[5191]) ^ (layer0_outputs[4420]));
    assign outputs[708] = layer0_outputs[3702];
    assign outputs[709] = ~((layer0_outputs[3999]) ^ (layer0_outputs[3804]));
    assign outputs[710] = layer0_outputs[4605];
    assign outputs[711] = ~((layer0_outputs[5372]) ^ (layer0_outputs[3385]));
    assign outputs[712] = layer0_outputs[6863];
    assign outputs[713] = (layer0_outputs[3084]) ^ (layer0_outputs[2265]);
    assign outputs[714] = layer0_outputs[2088];
    assign outputs[715] = ~((layer0_outputs[2103]) & (layer0_outputs[2477]));
    assign outputs[716] = (layer0_outputs[5544]) & (layer0_outputs[5828]);
    assign outputs[717] = (layer0_outputs[7212]) & ~(layer0_outputs[6190]);
    assign outputs[718] = ~(layer0_outputs[3519]);
    assign outputs[719] = (layer0_outputs[6284]) | (layer0_outputs[6858]);
    assign outputs[720] = (layer0_outputs[2227]) & ~(layer0_outputs[4081]);
    assign outputs[721] = 1'b1;
    assign outputs[722] = ~(layer0_outputs[4757]);
    assign outputs[723] = layer0_outputs[6489];
    assign outputs[724] = (layer0_outputs[6359]) & ~(layer0_outputs[2247]);
    assign outputs[725] = ~((layer0_outputs[3013]) ^ (layer0_outputs[6918]));
    assign outputs[726] = layer0_outputs[4486];
    assign outputs[727] = ~((layer0_outputs[2970]) ^ (layer0_outputs[5880]));
    assign outputs[728] = (layer0_outputs[2062]) & (layer0_outputs[5927]);
    assign outputs[729] = ~((layer0_outputs[4218]) | (layer0_outputs[2190]));
    assign outputs[730] = ~(layer0_outputs[6599]);
    assign outputs[731] = ~((layer0_outputs[967]) ^ (layer0_outputs[5637]));
    assign outputs[732] = ~((layer0_outputs[6553]) ^ (layer0_outputs[4395]));
    assign outputs[733] = ~(layer0_outputs[5043]);
    assign outputs[734] = layer0_outputs[5371];
    assign outputs[735] = (layer0_outputs[7351]) ^ (layer0_outputs[4852]);
    assign outputs[736] = (layer0_outputs[5234]) & ~(layer0_outputs[7570]);
    assign outputs[737] = layer0_outputs[2157];
    assign outputs[738] = ~(layer0_outputs[3675]) | (layer0_outputs[2502]);
    assign outputs[739] = layer0_outputs[1983];
    assign outputs[740] = ~(layer0_outputs[6983]);
    assign outputs[741] = ~(layer0_outputs[180]);
    assign outputs[742] = (layer0_outputs[3887]) & (layer0_outputs[2444]);
    assign outputs[743] = ~(layer0_outputs[2452]);
    assign outputs[744] = (layer0_outputs[4583]) ^ (layer0_outputs[2145]);
    assign outputs[745] = (layer0_outputs[5793]) ^ (layer0_outputs[3636]);
    assign outputs[746] = ~(layer0_outputs[4609]);
    assign outputs[747] = ~((layer0_outputs[1808]) & (layer0_outputs[7657]));
    assign outputs[748] = ~(layer0_outputs[3042]);
    assign outputs[749] = ~((layer0_outputs[6094]) ^ (layer0_outputs[3398]));
    assign outputs[750] = (layer0_outputs[3679]) ^ (layer0_outputs[2946]);
    assign outputs[751] = ~(layer0_outputs[3704]);
    assign outputs[752] = ~(layer0_outputs[5807]);
    assign outputs[753] = layer0_outputs[1219];
    assign outputs[754] = ~((layer0_outputs[4801]) ^ (layer0_outputs[6510]));
    assign outputs[755] = layer0_outputs[5206];
    assign outputs[756] = layer0_outputs[6693];
    assign outputs[757] = layer0_outputs[1340];
    assign outputs[758] = ~(layer0_outputs[4676]);
    assign outputs[759] = layer0_outputs[5003];
    assign outputs[760] = layer0_outputs[5466];
    assign outputs[761] = layer0_outputs[3170];
    assign outputs[762] = ~(layer0_outputs[2283]);
    assign outputs[763] = (layer0_outputs[7597]) & ~(layer0_outputs[6173]);
    assign outputs[764] = ~((layer0_outputs[5501]) ^ (layer0_outputs[2201]));
    assign outputs[765] = layer0_outputs[592];
    assign outputs[766] = layer0_outputs[6537];
    assign outputs[767] = layer0_outputs[1149];
    assign outputs[768] = ~(layer0_outputs[2883]);
    assign outputs[769] = (layer0_outputs[4185]) & ~(layer0_outputs[1324]);
    assign outputs[770] = (layer0_outputs[4405]) & ~(layer0_outputs[419]);
    assign outputs[771] = (layer0_outputs[4123]) & ~(layer0_outputs[4992]);
    assign outputs[772] = (layer0_outputs[6257]) & (layer0_outputs[3765]);
    assign outputs[773] = (layer0_outputs[1430]) & ~(layer0_outputs[1583]);
    assign outputs[774] = ~((layer0_outputs[6061]) | (layer0_outputs[4414]));
    assign outputs[775] = (layer0_outputs[3985]) & (layer0_outputs[5834]);
    assign outputs[776] = (layer0_outputs[5941]) & ~(layer0_outputs[7356]);
    assign outputs[777] = (layer0_outputs[6017]) ^ (layer0_outputs[6292]);
    assign outputs[778] = (layer0_outputs[3843]) & (layer0_outputs[819]);
    assign outputs[779] = (layer0_outputs[7073]) & ~(layer0_outputs[1322]);
    assign outputs[780] = ~((layer0_outputs[3498]) | (layer0_outputs[4366]));
    assign outputs[781] = (layer0_outputs[5692]) & ~(layer0_outputs[4733]);
    assign outputs[782] = ~(layer0_outputs[5857]);
    assign outputs[783] = (layer0_outputs[5402]) & ~(layer0_outputs[3133]);
    assign outputs[784] = (layer0_outputs[1894]) & ~(layer0_outputs[3360]);
    assign outputs[785] = ~(layer0_outputs[3649]);
    assign outputs[786] = (layer0_outputs[1063]) & ~(layer0_outputs[7421]);
    assign outputs[787] = (layer0_outputs[1915]) & (layer0_outputs[2818]);
    assign outputs[788] = (layer0_outputs[3796]) ^ (layer0_outputs[564]);
    assign outputs[789] = (layer0_outputs[2317]) & ~(layer0_outputs[3655]);
    assign outputs[790] = (layer0_outputs[6596]) & (layer0_outputs[7390]);
    assign outputs[791] = (layer0_outputs[2003]) & ~(layer0_outputs[2647]);
    assign outputs[792] = ~((layer0_outputs[1031]) ^ (layer0_outputs[5725]));
    assign outputs[793] = (layer0_outputs[4759]) & ~(layer0_outputs[6570]);
    assign outputs[794] = ~((layer0_outputs[6682]) | (layer0_outputs[2051]));
    assign outputs[795] = ~(layer0_outputs[5825]);
    assign outputs[796] = ~((layer0_outputs[2887]) | (layer0_outputs[1281]));
    assign outputs[797] = layer0_outputs[6639];
    assign outputs[798] = ~((layer0_outputs[5571]) | (layer0_outputs[191]));
    assign outputs[799] = ~((layer0_outputs[2725]) ^ (layer0_outputs[1282]));
    assign outputs[800] = (layer0_outputs[3948]) ^ (layer0_outputs[1129]);
    assign outputs[801] = (layer0_outputs[5176]) & ~(layer0_outputs[341]);
    assign outputs[802] = layer0_outputs[144];
    assign outputs[803] = (layer0_outputs[5447]) & (layer0_outputs[7412]);
    assign outputs[804] = (layer0_outputs[1492]) & ~(layer0_outputs[1744]);
    assign outputs[805] = ~((layer0_outputs[3640]) | (layer0_outputs[6226]));
    assign outputs[806] = ~((layer0_outputs[5709]) | (layer0_outputs[6977]));
    assign outputs[807] = ~((layer0_outputs[2951]) | (layer0_outputs[7460]));
    assign outputs[808] = ~(layer0_outputs[4322]) | (layer0_outputs[1016]);
    assign outputs[809] = (layer0_outputs[3025]) ^ (layer0_outputs[548]);
    assign outputs[810] = (layer0_outputs[3137]) & ~(layer0_outputs[5408]);
    assign outputs[811] = ~(layer0_outputs[3085]);
    assign outputs[812] = ~(layer0_outputs[2841]);
    assign outputs[813] = ~(layer0_outputs[1416]);
    assign outputs[814] = ~(layer0_outputs[2505]);
    assign outputs[815] = ~((layer0_outputs[5419]) | (layer0_outputs[2534]));
    assign outputs[816] = ~((layer0_outputs[6215]) ^ (layer0_outputs[928]));
    assign outputs[817] = ~((layer0_outputs[2080]) | (layer0_outputs[1819]));
    assign outputs[818] = (layer0_outputs[6807]) & (layer0_outputs[2853]);
    assign outputs[819] = ~(layer0_outputs[6066]);
    assign outputs[820] = (layer0_outputs[3436]) & ~(layer0_outputs[1295]);
    assign outputs[821] = (layer0_outputs[1137]) & ~(layer0_outputs[1786]);
    assign outputs[822] = ~((layer0_outputs[6131]) ^ (layer0_outputs[4532]));
    assign outputs[823] = ~(layer0_outputs[2424]);
    assign outputs[824] = ~(layer0_outputs[1421]);
    assign outputs[825] = (layer0_outputs[163]) & ~(layer0_outputs[1475]);
    assign outputs[826] = ~((layer0_outputs[3727]) | (layer0_outputs[2921]));
    assign outputs[827] = 1'b0;
    assign outputs[828] = (layer0_outputs[520]) & ~(layer0_outputs[1984]);
    assign outputs[829] = layer0_outputs[3037];
    assign outputs[830] = 1'b0;
    assign outputs[831] = layer0_outputs[4112];
    assign outputs[832] = ~(layer0_outputs[2004]);
    assign outputs[833] = ~(layer0_outputs[60]);
    assign outputs[834] = layer0_outputs[1932];
    assign outputs[835] = (layer0_outputs[6576]) & (layer0_outputs[2984]);
    assign outputs[836] = (layer0_outputs[3588]) & (layer0_outputs[2983]);
    assign outputs[837] = ~((layer0_outputs[3048]) | (layer0_outputs[1714]));
    assign outputs[838] = layer0_outputs[2174];
    assign outputs[839] = (layer0_outputs[1613]) & ~(layer0_outputs[584]);
    assign outputs[840] = layer0_outputs[7298];
    assign outputs[841] = ~((layer0_outputs[5729]) | (layer0_outputs[3749]));
    assign outputs[842] = (layer0_outputs[3245]) & ~(layer0_outputs[6240]);
    assign outputs[843] = ~(layer0_outputs[3009]);
    assign outputs[844] = ~(layer0_outputs[1864]);
    assign outputs[845] = (layer0_outputs[7148]) & ~(layer0_outputs[3391]);
    assign outputs[846] = layer0_outputs[3778];
    assign outputs[847] = ~(layer0_outputs[5826]);
    assign outputs[848] = (layer0_outputs[1996]) & ~(layer0_outputs[2073]);
    assign outputs[849] = (layer0_outputs[3707]) & ~(layer0_outputs[101]);
    assign outputs[850] = ~(layer0_outputs[5083]);
    assign outputs[851] = (layer0_outputs[6705]) & ~(layer0_outputs[4400]);
    assign outputs[852] = (layer0_outputs[5146]) & ~(layer0_outputs[5822]);
    assign outputs[853] = ~((layer0_outputs[3451]) | (layer0_outputs[3184]));
    assign outputs[854] = (layer0_outputs[5220]) & (layer0_outputs[1275]);
    assign outputs[855] = layer0_outputs[5215];
    assign outputs[856] = ~(layer0_outputs[1468]);
    assign outputs[857] = ~(layer0_outputs[7656]);
    assign outputs[858] = ~(layer0_outputs[6950]);
    assign outputs[859] = (layer0_outputs[4593]) ^ (layer0_outputs[2919]);
    assign outputs[860] = ~((layer0_outputs[2144]) | (layer0_outputs[3131]));
    assign outputs[861] = (layer0_outputs[1246]) & ~(layer0_outputs[1882]);
    assign outputs[862] = ~(layer0_outputs[5819]);
    assign outputs[863] = (layer0_outputs[7481]) & ~(layer0_outputs[975]);
    assign outputs[864] = ~((layer0_outputs[2819]) | (layer0_outputs[5275]));
    assign outputs[865] = (layer0_outputs[747]) & ~(layer0_outputs[4532]);
    assign outputs[866] = (layer0_outputs[6855]) & (layer0_outputs[734]);
    assign outputs[867] = (layer0_outputs[4896]) & (layer0_outputs[3701]);
    assign outputs[868] = layer0_outputs[4487];
    assign outputs[869] = layer0_outputs[7029];
    assign outputs[870] = ~((layer0_outputs[4331]) | (layer0_outputs[6718]));
    assign outputs[871] = (layer0_outputs[1697]) & ~(layer0_outputs[2095]);
    assign outputs[872] = (layer0_outputs[775]) & ~(layer0_outputs[7331]);
    assign outputs[873] = ~((layer0_outputs[4476]) | (layer0_outputs[7093]));
    assign outputs[874] = (layer0_outputs[7019]) ^ (layer0_outputs[4857]);
    assign outputs[875] = ~(layer0_outputs[7243]);
    assign outputs[876] = (layer0_outputs[5863]) & ~(layer0_outputs[2917]);
    assign outputs[877] = (layer0_outputs[4662]) & (layer0_outputs[7129]);
    assign outputs[878] = (layer0_outputs[5618]) & (layer0_outputs[4888]);
    assign outputs[879] = ~(layer0_outputs[1446]);
    assign outputs[880] = ~((layer0_outputs[3129]) ^ (layer0_outputs[2298]));
    assign outputs[881] = (layer0_outputs[428]) & ~(layer0_outputs[3228]);
    assign outputs[882] = ~((layer0_outputs[7617]) | (layer0_outputs[7625]));
    assign outputs[883] = ~((layer0_outputs[6541]) & (layer0_outputs[5117]));
    assign outputs[884] = (layer0_outputs[4169]) | (layer0_outputs[3188]);
    assign outputs[885] = (layer0_outputs[5892]) & ~(layer0_outputs[1028]);
    assign outputs[886] = ~((layer0_outputs[6790]) ^ (layer0_outputs[1224]));
    assign outputs[887] = (layer0_outputs[5884]) & (layer0_outputs[3373]);
    assign outputs[888] = (layer0_outputs[4565]) ^ (layer0_outputs[4816]);
    assign outputs[889] = (layer0_outputs[4821]) ^ (layer0_outputs[3776]);
    assign outputs[890] = (layer0_outputs[2114]) & ~(layer0_outputs[4462]);
    assign outputs[891] = (layer0_outputs[3949]) & ~(layer0_outputs[6649]);
    assign outputs[892] = ~((layer0_outputs[5337]) | (layer0_outputs[5846]));
    assign outputs[893] = ~(layer0_outputs[5373]);
    assign outputs[894] = ~(layer0_outputs[5179]);
    assign outputs[895] = (layer0_outputs[2693]) & ~(layer0_outputs[7507]);
    assign outputs[896] = 1'b0;
    assign outputs[897] = (layer0_outputs[4788]) & (layer0_outputs[4782]);
    assign outputs[898] = (layer0_outputs[4117]) & (layer0_outputs[7519]);
    assign outputs[899] = (layer0_outputs[967]) & ~(layer0_outputs[1079]);
    assign outputs[900] = (layer0_outputs[2580]) & (layer0_outputs[7666]);
    assign outputs[901] = (layer0_outputs[2700]) & ~(layer0_outputs[3684]);
    assign outputs[902] = (layer0_outputs[5032]) ^ (layer0_outputs[5040]);
    assign outputs[903] = layer0_outputs[2689];
    assign outputs[904] = 1'b0;
    assign outputs[905] = ~((layer0_outputs[5485]) ^ (layer0_outputs[6610]));
    assign outputs[906] = (layer0_outputs[2125]) & ~(layer0_outputs[1066]);
    assign outputs[907] = (layer0_outputs[3874]) & ~(layer0_outputs[6021]);
    assign outputs[908] = (layer0_outputs[7035]) & ~(layer0_outputs[813]);
    assign outputs[909] = ~(layer0_outputs[837]);
    assign outputs[910] = (layer0_outputs[1930]) & ~(layer0_outputs[4776]);
    assign outputs[911] = (layer0_outputs[3773]) & (layer0_outputs[4253]);
    assign outputs[912] = (layer0_outputs[6293]) & ~(layer0_outputs[2826]);
    assign outputs[913] = (layer0_outputs[983]) & ~(layer0_outputs[879]);
    assign outputs[914] = ~(layer0_outputs[3496]);
    assign outputs[915] = (layer0_outputs[7557]) & ~(layer0_outputs[3094]);
    assign outputs[916] = layer0_outputs[6957];
    assign outputs[917] = (layer0_outputs[6811]) & ~(layer0_outputs[6790]);
    assign outputs[918] = layer0_outputs[3232];
    assign outputs[919] = ~((layer0_outputs[4678]) | (layer0_outputs[3463]));
    assign outputs[920] = (layer0_outputs[4727]) & ~(layer0_outputs[1121]);
    assign outputs[921] = ~((layer0_outputs[7238]) | (layer0_outputs[2926]));
    assign outputs[922] = (layer0_outputs[899]) & ~(layer0_outputs[4195]);
    assign outputs[923] = ~(layer0_outputs[2877]);
    assign outputs[924] = (layer0_outputs[5290]) & ~(layer0_outputs[6661]);
    assign outputs[925] = ~((layer0_outputs[529]) ^ (layer0_outputs[1627]));
    assign outputs[926] = layer0_outputs[7445];
    assign outputs[927] = layer0_outputs[6971];
    assign outputs[928] = ~((layer0_outputs[638]) | (layer0_outputs[1284]));
    assign outputs[929] = (layer0_outputs[266]) & (layer0_outputs[5090]);
    assign outputs[930] = ~((layer0_outputs[7365]) ^ (layer0_outputs[1494]));
    assign outputs[931] = (layer0_outputs[2031]) & ~(layer0_outputs[5446]);
    assign outputs[932] = layer0_outputs[1905];
    assign outputs[933] = ~((layer0_outputs[327]) | (layer0_outputs[1797]));
    assign outputs[934] = ~((layer0_outputs[5092]) | (layer0_outputs[1873]));
    assign outputs[935] = (layer0_outputs[1484]) & (layer0_outputs[5574]);
    assign outputs[936] = (layer0_outputs[2344]) & ~(layer0_outputs[6330]);
    assign outputs[937] = layer0_outputs[3045];
    assign outputs[938] = layer0_outputs[1398];
    assign outputs[939] = (layer0_outputs[4384]) & ~(layer0_outputs[4193]);
    assign outputs[940] = (layer0_outputs[539]) & ~(layer0_outputs[2047]);
    assign outputs[941] = (layer0_outputs[6935]) & ~(layer0_outputs[4791]);
    assign outputs[942] = (layer0_outputs[3143]) ^ (layer0_outputs[2067]);
    assign outputs[943] = ~(layer0_outputs[905]);
    assign outputs[944] = ~(layer0_outputs[6109]);
    assign outputs[945] = (layer0_outputs[223]) & (layer0_outputs[2721]);
    assign outputs[946] = (layer0_outputs[6055]) & ~(layer0_outputs[7277]);
    assign outputs[947] = ~(layer0_outputs[1499]);
    assign outputs[948] = (layer0_outputs[7552]) & ~(layer0_outputs[5397]);
    assign outputs[949] = (layer0_outputs[6323]) & ~(layer0_outputs[1013]);
    assign outputs[950] = (layer0_outputs[4496]) ^ (layer0_outputs[1344]);
    assign outputs[951] = (layer0_outputs[3328]) & ~(layer0_outputs[4874]);
    assign outputs[952] = (layer0_outputs[5760]) & ~(layer0_outputs[3565]);
    assign outputs[953] = (layer0_outputs[5486]) & ~(layer0_outputs[4770]);
    assign outputs[954] = 1'b0;
    assign outputs[955] = (layer0_outputs[5769]) ^ (layer0_outputs[7617]);
    assign outputs[956] = (layer0_outputs[6822]) & (layer0_outputs[3452]);
    assign outputs[957] = (layer0_outputs[382]) & ~(layer0_outputs[5688]);
    assign outputs[958] = ~(layer0_outputs[5882]);
    assign outputs[959] = (layer0_outputs[2024]) & ~(layer0_outputs[6463]);
    assign outputs[960] = ~((layer0_outputs[6106]) | (layer0_outputs[6644]));
    assign outputs[961] = ~((layer0_outputs[6031]) | (layer0_outputs[4288]));
    assign outputs[962] = layer0_outputs[6941];
    assign outputs[963] = ~((layer0_outputs[4337]) | (layer0_outputs[7413]));
    assign outputs[964] = ~(layer0_outputs[4700]);
    assign outputs[965] = ~(layer0_outputs[1507]);
    assign outputs[966] = (layer0_outputs[5592]) & ~(layer0_outputs[1878]);
    assign outputs[967] = ~(layer0_outputs[6469]);
    assign outputs[968] = ~((layer0_outputs[2429]) | (layer0_outputs[3602]));
    assign outputs[969] = layer0_outputs[2531];
    assign outputs[970] = (layer0_outputs[639]) & ~(layer0_outputs[6723]);
    assign outputs[971] = layer0_outputs[454];
    assign outputs[972] = ~((layer0_outputs[2211]) ^ (layer0_outputs[7176]));
    assign outputs[973] = ~((layer0_outputs[3930]) | (layer0_outputs[7665]));
    assign outputs[974] = (layer0_outputs[3082]) & (layer0_outputs[2986]);
    assign outputs[975] = (layer0_outputs[3856]) ^ (layer0_outputs[5024]);
    assign outputs[976] = (layer0_outputs[6055]) & (layer0_outputs[7350]);
    assign outputs[977] = ~((layer0_outputs[3791]) | (layer0_outputs[6849]));
    assign outputs[978] = (layer0_outputs[6140]) & ~(layer0_outputs[2576]);
    assign outputs[979] = ~((layer0_outputs[4251]) | (layer0_outputs[359]));
    assign outputs[980] = ~(layer0_outputs[7188]);
    assign outputs[981] = (layer0_outputs[1669]) & ~(layer0_outputs[5606]);
    assign outputs[982] = ~(layer0_outputs[2109]);
    assign outputs[983] = (layer0_outputs[2715]) ^ (layer0_outputs[2875]);
    assign outputs[984] = (layer0_outputs[5625]) & ~(layer0_outputs[2226]);
    assign outputs[985] = ~(layer0_outputs[4436]);
    assign outputs[986] = (layer0_outputs[6039]) ^ (layer0_outputs[6934]);
    assign outputs[987] = layer0_outputs[5522];
    assign outputs[988] = (layer0_outputs[4736]) & ~(layer0_outputs[1343]);
    assign outputs[989] = (layer0_outputs[6978]) & ~(layer0_outputs[4802]);
    assign outputs[990] = ~(layer0_outputs[2243]);
    assign outputs[991] = (layer0_outputs[1554]) & ~(layer0_outputs[3152]);
    assign outputs[992] = (layer0_outputs[320]) & (layer0_outputs[2741]);
    assign outputs[993] = ~(layer0_outputs[3831]);
    assign outputs[994] = ~((layer0_outputs[509]) ^ (layer0_outputs[1181]));
    assign outputs[995] = ~((layer0_outputs[7041]) | (layer0_outputs[6775]));
    assign outputs[996] = layer0_outputs[2538];
    assign outputs[997] = (layer0_outputs[3106]) & ~(layer0_outputs[3267]);
    assign outputs[998] = layer0_outputs[7636];
    assign outputs[999] = ~((layer0_outputs[4592]) | (layer0_outputs[6390]));
    assign outputs[1000] = (layer0_outputs[3547]) ^ (layer0_outputs[2308]);
    assign outputs[1001] = ~(layer0_outputs[3099]);
    assign outputs[1002] = ~((layer0_outputs[6042]) | (layer0_outputs[5816]));
    assign outputs[1003] = ~(layer0_outputs[5935]);
    assign outputs[1004] = 1'b0;
    assign outputs[1005] = ~(layer0_outputs[253]);
    assign outputs[1006] = layer0_outputs[4089];
    assign outputs[1007] = ~((layer0_outputs[5233]) | (layer0_outputs[4202]));
    assign outputs[1008] = ~((layer0_outputs[3265]) | (layer0_outputs[1738]));
    assign outputs[1009] = (layer0_outputs[36]) & (layer0_outputs[6159]);
    assign outputs[1010] = 1'b0;
    assign outputs[1011] = ~((layer0_outputs[7505]) | (layer0_outputs[4433]));
    assign outputs[1012] = (layer0_outputs[4245]) & ~(layer0_outputs[7162]);
    assign outputs[1013] = ~((layer0_outputs[2584]) | (layer0_outputs[2171]));
    assign outputs[1014] = (layer0_outputs[4983]) & (layer0_outputs[1560]);
    assign outputs[1015] = layer0_outputs[2127];
    assign outputs[1016] = (layer0_outputs[6970]) & (layer0_outputs[6959]);
    assign outputs[1017] = (layer0_outputs[2251]) & ~(layer0_outputs[4504]);
    assign outputs[1018] = (layer0_outputs[2373]) & (layer0_outputs[7576]);
    assign outputs[1019] = ~(layer0_outputs[6286]);
    assign outputs[1020] = (layer0_outputs[1906]) & ~(layer0_outputs[5184]);
    assign outputs[1021] = ~((layer0_outputs[1043]) ^ (layer0_outputs[2632]));
    assign outputs[1022] = ~((layer0_outputs[7088]) | (layer0_outputs[7375]));
    assign outputs[1023] = (layer0_outputs[4330]) & ~(layer0_outputs[2468]);
    assign outputs[1024] = ~((layer0_outputs[5491]) | (layer0_outputs[7182]));
    assign outputs[1025] = (layer0_outputs[6771]) & ~(layer0_outputs[2417]);
    assign outputs[1026] = (layer0_outputs[6493]) & (layer0_outputs[4551]);
    assign outputs[1027] = (layer0_outputs[6756]) & ~(layer0_outputs[6932]);
    assign outputs[1028] = (layer0_outputs[942]) & ~(layer0_outputs[3231]);
    assign outputs[1029] = (layer0_outputs[3303]) & ~(layer0_outputs[6541]);
    assign outputs[1030] = ~((layer0_outputs[4010]) | (layer0_outputs[364]));
    assign outputs[1031] = (layer0_outputs[1220]) & ~(layer0_outputs[7174]);
    assign outputs[1032] = (layer0_outputs[7404]) & ~(layer0_outputs[400]);
    assign outputs[1033] = ~(layer0_outputs[4180]);
    assign outputs[1034] = (layer0_outputs[4273]) & ~(layer0_outputs[1864]);
    assign outputs[1035] = (layer0_outputs[3631]) & ~(layer0_outputs[1678]);
    assign outputs[1036] = ~(layer0_outputs[470]);
    assign outputs[1037] = (layer0_outputs[4318]) ^ (layer0_outputs[2994]);
    assign outputs[1038] = (layer0_outputs[2244]) & ~(layer0_outputs[543]);
    assign outputs[1039] = (layer0_outputs[1778]) & (layer0_outputs[4873]);
    assign outputs[1040] = (layer0_outputs[7575]) & (layer0_outputs[175]);
    assign outputs[1041] = (layer0_outputs[4097]) & (layer0_outputs[2634]);
    assign outputs[1042] = (layer0_outputs[712]) & ~(layer0_outputs[7195]);
    assign outputs[1043] = ~((layer0_outputs[5795]) ^ (layer0_outputs[2447]));
    assign outputs[1044] = ~((layer0_outputs[6828]) ^ (layer0_outputs[3414]));
    assign outputs[1045] = (layer0_outputs[779]) | (layer0_outputs[1462]);
    assign outputs[1046] = layer0_outputs[1425];
    assign outputs[1047] = (layer0_outputs[5743]) & (layer0_outputs[2466]);
    assign outputs[1048] = ~(layer0_outputs[3913]);
    assign outputs[1049] = ~(layer0_outputs[2471]);
    assign outputs[1050] = layer0_outputs[1035];
    assign outputs[1051] = (layer0_outputs[5302]) ^ (layer0_outputs[1258]);
    assign outputs[1052] = ~(layer0_outputs[1164]);
    assign outputs[1053] = (layer0_outputs[2645]) & (layer0_outputs[3866]);
    assign outputs[1054] = (layer0_outputs[976]) ^ (layer0_outputs[3138]);
    assign outputs[1055] = (layer0_outputs[4324]) & ~(layer0_outputs[194]);
    assign outputs[1056] = ~((layer0_outputs[3236]) | (layer0_outputs[989]));
    assign outputs[1057] = (layer0_outputs[1974]) & (layer0_outputs[3946]);
    assign outputs[1058] = (layer0_outputs[611]) & ~(layer0_outputs[5670]);
    assign outputs[1059] = ~(layer0_outputs[5951]);
    assign outputs[1060] = layer0_outputs[5238];
    assign outputs[1061] = ~((layer0_outputs[5236]) ^ (layer0_outputs[424]));
    assign outputs[1062] = (layer0_outputs[5069]) & ~(layer0_outputs[1243]);
    assign outputs[1063] = (layer0_outputs[1114]) & ~(layer0_outputs[3190]);
    assign outputs[1064] = ~((layer0_outputs[982]) ^ (layer0_outputs[103]));
    assign outputs[1065] = (layer0_outputs[6719]) & ~(layer0_outputs[6371]);
    assign outputs[1066] = (layer0_outputs[6978]) & (layer0_outputs[5289]);
    assign outputs[1067] = (layer0_outputs[2353]) & (layer0_outputs[1895]);
    assign outputs[1068] = (layer0_outputs[5081]) & (layer0_outputs[6346]);
    assign outputs[1069] = 1'b0;
    assign outputs[1070] = layer0_outputs[574];
    assign outputs[1071] = (layer0_outputs[4186]) & ~(layer0_outputs[1463]);
    assign outputs[1072] = ~((layer0_outputs[5730]) ^ (layer0_outputs[3286]));
    assign outputs[1073] = (layer0_outputs[2866]) ^ (layer0_outputs[7193]);
    assign outputs[1074] = layer0_outputs[4815];
    assign outputs[1075] = ~((layer0_outputs[214]) | (layer0_outputs[1599]));
    assign outputs[1076] = (layer0_outputs[2699]) & ~(layer0_outputs[3309]);
    assign outputs[1077] = ~((layer0_outputs[5059]) | (layer0_outputs[147]));
    assign outputs[1078] = ~(layer0_outputs[3504]);
    assign outputs[1079] = ~((layer0_outputs[6296]) | (layer0_outputs[3161]));
    assign outputs[1080] = ~(layer0_outputs[3714]);
    assign outputs[1081] = 1'b0;
    assign outputs[1082] = ~(layer0_outputs[7197]);
    assign outputs[1083] = ~((layer0_outputs[3397]) | (layer0_outputs[5330]));
    assign outputs[1084] = 1'b0;
    assign outputs[1085] = ~((layer0_outputs[5877]) | (layer0_outputs[353]));
    assign outputs[1086] = (layer0_outputs[6009]) & (layer0_outputs[3753]);
    assign outputs[1087] = ~(layer0_outputs[656]);
    assign outputs[1088] = ~((layer0_outputs[1070]) ^ (layer0_outputs[6894]));
    assign outputs[1089] = layer0_outputs[7394];
    assign outputs[1090] = 1'b0;
    assign outputs[1091] = ~(layer0_outputs[3120]);
    assign outputs[1092] = (layer0_outputs[6438]) & ~(layer0_outputs[4073]);
    assign outputs[1093] = (layer0_outputs[7317]) & ~(layer0_outputs[1544]);
    assign outputs[1094] = (layer0_outputs[7444]) & (layer0_outputs[7141]);
    assign outputs[1095] = 1'b0;
    assign outputs[1096] = ~(layer0_outputs[3004]) | (layer0_outputs[2598]);
    assign outputs[1097] = (layer0_outputs[1503]) & (layer0_outputs[5357]);
    assign outputs[1098] = ~((layer0_outputs[6602]) | (layer0_outputs[6436]));
    assign outputs[1099] = layer0_outputs[450];
    assign outputs[1100] = 1'b0;
    assign outputs[1101] = ~(layer0_outputs[4203]) | (layer0_outputs[3087]);
    assign outputs[1102] = 1'b0;
    assign outputs[1103] = (layer0_outputs[6402]) ^ (layer0_outputs[2424]);
    assign outputs[1104] = ~((layer0_outputs[2629]) ^ (layer0_outputs[6245]));
    assign outputs[1105] = (layer0_outputs[5767]) & ~(layer0_outputs[1156]);
    assign outputs[1106] = (layer0_outputs[2393]) & (layer0_outputs[6497]);
    assign outputs[1107] = (layer0_outputs[3417]) & ~(layer0_outputs[6449]);
    assign outputs[1108] = (layer0_outputs[5262]) & ~(layer0_outputs[973]);
    assign outputs[1109] = (layer0_outputs[5572]) & ~(layer0_outputs[7154]);
    assign outputs[1110] = (layer0_outputs[4387]) & (layer0_outputs[1092]);
    assign outputs[1111] = (layer0_outputs[657]) & ~(layer0_outputs[1606]);
    assign outputs[1112] = ~(layer0_outputs[572]);
    assign outputs[1113] = (layer0_outputs[6443]) & ~(layer0_outputs[2241]);
    assign outputs[1114] = layer0_outputs[3416];
    assign outputs[1115] = (layer0_outputs[6954]) & ~(layer0_outputs[3246]);
    assign outputs[1116] = ~(layer0_outputs[3156]);
    assign outputs[1117] = layer0_outputs[7422];
    assign outputs[1118] = (layer0_outputs[1431]) & ~(layer0_outputs[1223]);
    assign outputs[1119] = (layer0_outputs[3573]) & ~(layer0_outputs[4971]);
    assign outputs[1120] = layer0_outputs[5181];
    assign outputs[1121] = ~((layer0_outputs[7266]) ^ (layer0_outputs[2863]));
    assign outputs[1122] = ~((layer0_outputs[1094]) ^ (layer0_outputs[884]));
    assign outputs[1123] = ~(layer0_outputs[2390]);
    assign outputs[1124] = (layer0_outputs[4914]) & ~(layer0_outputs[4237]);
    assign outputs[1125] = ~((layer0_outputs[7225]) | (layer0_outputs[7203]));
    assign outputs[1126] = layer0_outputs[5917];
    assign outputs[1127] = (layer0_outputs[4147]) & ~(layer0_outputs[6183]);
    assign outputs[1128] = (layer0_outputs[1985]) & ~(layer0_outputs[64]);
    assign outputs[1129] = (layer0_outputs[1489]) & ~(layer0_outputs[6380]);
    assign outputs[1130] = ~((layer0_outputs[1631]) ^ (layer0_outputs[6099]));
    assign outputs[1131] = ~((layer0_outputs[3038]) & (layer0_outputs[2684]));
    assign outputs[1132] = ~(layer0_outputs[5749]);
    assign outputs[1133] = (layer0_outputs[5334]) & ~(layer0_outputs[2850]);
    assign outputs[1134] = layer0_outputs[393];
    assign outputs[1135] = ~((layer0_outputs[181]) ^ (layer0_outputs[6152]));
    assign outputs[1136] = (layer0_outputs[4216]) ^ (layer0_outputs[2403]);
    assign outputs[1137] = ~((layer0_outputs[6783]) | (layer0_outputs[849]));
    assign outputs[1138] = 1'b0;
    assign outputs[1139] = layer0_outputs[6918];
    assign outputs[1140] = ~(layer0_outputs[3312]);
    assign outputs[1141] = layer0_outputs[184];
    assign outputs[1142] = (layer0_outputs[4726]) & ~(layer0_outputs[6803]);
    assign outputs[1143] = layer0_outputs[2162];
    assign outputs[1144] = ~((layer0_outputs[3797]) | (layer0_outputs[5450]));
    assign outputs[1145] = (layer0_outputs[7047]) & ~(layer0_outputs[3570]);
    assign outputs[1146] = ~(layer0_outputs[4160]);
    assign outputs[1147] = (layer0_outputs[3827]) & (layer0_outputs[4005]);
    assign outputs[1148] = (layer0_outputs[2318]) ^ (layer0_outputs[4067]);
    assign outputs[1149] = (layer0_outputs[4022]) & ~(layer0_outputs[4003]);
    assign outputs[1150] = (layer0_outputs[4388]) & ~(layer0_outputs[3180]);
    assign outputs[1151] = (layer0_outputs[631]) ^ (layer0_outputs[3371]);
    assign outputs[1152] = ~((layer0_outputs[2117]) | (layer0_outputs[7157]));
    assign outputs[1153] = ~(layer0_outputs[115]);
    assign outputs[1154] = (layer0_outputs[1237]) & ~(layer0_outputs[6559]);
    assign outputs[1155] = (layer0_outputs[2023]) & ~(layer0_outputs[4798]);
    assign outputs[1156] = (layer0_outputs[7251]) & (layer0_outputs[977]);
    assign outputs[1157] = (layer0_outputs[5334]) & ~(layer0_outputs[4448]);
    assign outputs[1158] = (layer0_outputs[4720]) & ~(layer0_outputs[2349]);
    assign outputs[1159] = ~((layer0_outputs[2782]) | (layer0_outputs[5116]));
    assign outputs[1160] = (layer0_outputs[740]) & (layer0_outputs[5995]);
    assign outputs[1161] = ~(layer0_outputs[3967]);
    assign outputs[1162] = layer0_outputs[1272];
    assign outputs[1163] = ~(layer0_outputs[7102]) | (layer0_outputs[5972]);
    assign outputs[1164] = ~((layer0_outputs[7053]) | (layer0_outputs[3281]));
    assign outputs[1165] = (layer0_outputs[206]) & ~(layer0_outputs[6078]);
    assign outputs[1166] = (layer0_outputs[5251]) & ~(layer0_outputs[208]);
    assign outputs[1167] = layer0_outputs[2238];
    assign outputs[1168] = (layer0_outputs[85]) & ~(layer0_outputs[5861]);
    assign outputs[1169] = (layer0_outputs[4759]) & ~(layer0_outputs[1540]);
    assign outputs[1170] = ~(layer0_outputs[6507]);
    assign outputs[1171] = (layer0_outputs[1575]) & (layer0_outputs[3082]);
    assign outputs[1172] = ~(layer0_outputs[4513]);
    assign outputs[1173] = ~((layer0_outputs[616]) ^ (layer0_outputs[2475]));
    assign outputs[1174] = layer0_outputs[3356];
    assign outputs[1175] = ~((layer0_outputs[14]) ^ (layer0_outputs[4408]));
    assign outputs[1176] = (layer0_outputs[1677]) & (layer0_outputs[1318]);
    assign outputs[1177] = layer0_outputs[5290];
    assign outputs[1178] = ~(layer0_outputs[6945]);
    assign outputs[1179] = (layer0_outputs[1341]) & ~(layer0_outputs[4271]);
    assign outputs[1180] = (layer0_outputs[3937]) & ~(layer0_outputs[1199]);
    assign outputs[1181] = (layer0_outputs[4025]) & ~(layer0_outputs[243]);
    assign outputs[1182] = ~((layer0_outputs[4492]) | (layer0_outputs[7024]));
    assign outputs[1183] = ~(layer0_outputs[6074]);
    assign outputs[1184] = (layer0_outputs[6032]) & ~(layer0_outputs[3298]);
    assign outputs[1185] = (layer0_outputs[5745]) & ~(layer0_outputs[4747]);
    assign outputs[1186] = (layer0_outputs[6506]) | (layer0_outputs[4399]);
    assign outputs[1187] = (layer0_outputs[5580]) & ~(layer0_outputs[4909]);
    assign outputs[1188] = layer0_outputs[7305];
    assign outputs[1189] = layer0_outputs[2068];
    assign outputs[1190] = ~((layer0_outputs[1066]) ^ (layer0_outputs[5507]));
    assign outputs[1191] = ~(layer0_outputs[6784]);
    assign outputs[1192] = (layer0_outputs[4690]) & ~(layer0_outputs[5061]);
    assign outputs[1193] = ~((layer0_outputs[3389]) | (layer0_outputs[4655]));
    assign outputs[1194] = ~((layer0_outputs[2376]) ^ (layer0_outputs[6252]));
    assign outputs[1195] = ~((layer0_outputs[790]) | (layer0_outputs[3940]));
    assign outputs[1196] = ~(layer0_outputs[5360]);
    assign outputs[1197] = (layer0_outputs[5337]) ^ (layer0_outputs[702]);
    assign outputs[1198] = ~((layer0_outputs[7341]) | (layer0_outputs[2007]));
    assign outputs[1199] = ~(layer0_outputs[1960]);
    assign outputs[1200] = ~(layer0_outputs[7395]);
    assign outputs[1201] = layer0_outputs[5085];
    assign outputs[1202] = ~(layer0_outputs[883]);
    assign outputs[1203] = (layer0_outputs[1242]) & ~(layer0_outputs[7258]);
    assign outputs[1204] = ~(layer0_outputs[5590]);
    assign outputs[1205] = ~(layer0_outputs[2457]);
    assign outputs[1206] = (layer0_outputs[1615]) & ~(layer0_outputs[985]);
    assign outputs[1207] = (layer0_outputs[4170]) & ~(layer0_outputs[7362]);
    assign outputs[1208] = (layer0_outputs[2527]) & (layer0_outputs[2481]);
    assign outputs[1209] = ~((layer0_outputs[2967]) ^ (layer0_outputs[5516]));
    assign outputs[1210] = (layer0_outputs[5448]) & (layer0_outputs[6130]);
    assign outputs[1211] = ~(layer0_outputs[7637]);
    assign outputs[1212] = (layer0_outputs[3976]) & (layer0_outputs[5708]);
    assign outputs[1213] = ~((layer0_outputs[6914]) | (layer0_outputs[7582]));
    assign outputs[1214] = ~((layer0_outputs[5391]) & (layer0_outputs[5747]));
    assign outputs[1215] = (layer0_outputs[5452]) & (layer0_outputs[4675]);
    assign outputs[1216] = layer0_outputs[6886];
    assign outputs[1217] = (layer0_outputs[5648]) & ~(layer0_outputs[418]);
    assign outputs[1218] = (layer0_outputs[338]) ^ (layer0_outputs[4558]);
    assign outputs[1219] = (layer0_outputs[2491]) & ~(layer0_outputs[5810]);
    assign outputs[1220] = layer0_outputs[3253];
    assign outputs[1221] = layer0_outputs[2182];
    assign outputs[1222] = ~((layer0_outputs[2968]) | (layer0_outputs[350]));
    assign outputs[1223] = (layer0_outputs[5270]) & (layer0_outputs[2940]);
    assign outputs[1224] = ~(layer0_outputs[3717]);
    assign outputs[1225] = (layer0_outputs[648]) & ~(layer0_outputs[217]);
    assign outputs[1226] = layer0_outputs[4453];
    assign outputs[1227] = ~((layer0_outputs[373]) ^ (layer0_outputs[3007]));
    assign outputs[1228] = (layer0_outputs[7020]) & (layer0_outputs[6468]);
    assign outputs[1229] = (layer0_outputs[664]) ^ (layer0_outputs[6116]);
    assign outputs[1230] = (layer0_outputs[3639]) ^ (layer0_outputs[5621]);
    assign outputs[1231] = ~((layer0_outputs[1539]) ^ (layer0_outputs[3975]));
    assign outputs[1232] = ~(layer0_outputs[5210]);
    assign outputs[1233] = (layer0_outputs[3467]) ^ (layer0_outputs[682]);
    assign outputs[1234] = ~((layer0_outputs[2921]) | (layer0_outputs[3812]));
    assign outputs[1235] = ~((layer0_outputs[4760]) | (layer0_outputs[1552]));
    assign outputs[1236] = layer0_outputs[2492];
    assign outputs[1237] = ~(layer0_outputs[5457]);
    assign outputs[1238] = ~(layer0_outputs[6195]);
    assign outputs[1239] = (layer0_outputs[5226]) & ~(layer0_outputs[4836]);
    assign outputs[1240] = layer0_outputs[6494];
    assign outputs[1241] = layer0_outputs[131];
    assign outputs[1242] = layer0_outputs[5509];
    assign outputs[1243] = 1'b0;
    assign outputs[1244] = (layer0_outputs[5973]) & ~(layer0_outputs[3432]);
    assign outputs[1245] = (layer0_outputs[5811]) & (layer0_outputs[2350]);
    assign outputs[1246] = ~(layer0_outputs[289]);
    assign outputs[1247] = ~(layer0_outputs[3578]);
    assign outputs[1248] = (layer0_outputs[2973]) & ~(layer0_outputs[3686]);
    assign outputs[1249] = (layer0_outputs[626]) & ~(layer0_outputs[5083]);
    assign outputs[1250] = (layer0_outputs[4206]) ^ (layer0_outputs[2280]);
    assign outputs[1251] = (layer0_outputs[4423]) & ~(layer0_outputs[5942]);
    assign outputs[1252] = (layer0_outputs[758]) & ~(layer0_outputs[6199]);
    assign outputs[1253] = (layer0_outputs[4976]) & (layer0_outputs[3928]);
    assign outputs[1254] = layer0_outputs[6388];
    assign outputs[1255] = (layer0_outputs[681]) & (layer0_outputs[1948]);
    assign outputs[1256] = (layer0_outputs[2821]) & ~(layer0_outputs[465]);
    assign outputs[1257] = layer0_outputs[206];
    assign outputs[1258] = (layer0_outputs[4788]) & ~(layer0_outputs[6907]);
    assign outputs[1259] = ~(layer0_outputs[733]);
    assign outputs[1260] = (layer0_outputs[212]) & (layer0_outputs[5452]);
    assign outputs[1261] = layer0_outputs[3971];
    assign outputs[1262] = (layer0_outputs[794]) & (layer0_outputs[2293]);
    assign outputs[1263] = (layer0_outputs[405]) & ~(layer0_outputs[293]);
    assign outputs[1264] = (layer0_outputs[5092]) & ~(layer0_outputs[4376]);
    assign outputs[1265] = ~((layer0_outputs[5487]) | (layer0_outputs[6839]));
    assign outputs[1266] = (layer0_outputs[3130]) & (layer0_outputs[1547]);
    assign outputs[1267] = ~(layer0_outputs[3654]);
    assign outputs[1268] = ~((layer0_outputs[1441]) | (layer0_outputs[3968]));
    assign outputs[1269] = (layer0_outputs[3672]) & (layer0_outputs[454]);
    assign outputs[1270] = (layer0_outputs[1979]) & ~(layer0_outputs[7328]);
    assign outputs[1271] = (layer0_outputs[1964]) & ~(layer0_outputs[3432]);
    assign outputs[1272] = (layer0_outputs[1217]) & ~(layer0_outputs[4813]);
    assign outputs[1273] = ~((layer0_outputs[134]) | (layer0_outputs[4818]));
    assign outputs[1274] = ~(layer0_outputs[1559]);
    assign outputs[1275] = (layer0_outputs[6798]) & ~(layer0_outputs[3318]);
    assign outputs[1276] = layer0_outputs[6236];
    assign outputs[1277] = (layer0_outputs[976]) & ~(layer0_outputs[1507]);
    assign outputs[1278] = (layer0_outputs[1620]) & (layer0_outputs[5914]);
    assign outputs[1279] = layer0_outputs[7657];
    assign outputs[1280] = (layer0_outputs[7429]) ^ (layer0_outputs[4537]);
    assign outputs[1281] = (layer0_outputs[5206]) & ~(layer0_outputs[6275]);
    assign outputs[1282] = (layer0_outputs[1859]) & (layer0_outputs[232]);
    assign outputs[1283] = (layer0_outputs[7515]) & (layer0_outputs[7484]);
    assign outputs[1284] = ~(layer0_outputs[2657]);
    assign outputs[1285] = 1'b0;
    assign outputs[1286] = ~((layer0_outputs[6386]) | (layer0_outputs[7333]));
    assign outputs[1287] = (layer0_outputs[5864]) & ~(layer0_outputs[4639]);
    assign outputs[1288] = layer0_outputs[1724];
    assign outputs[1289] = ~(layer0_outputs[4959]);
    assign outputs[1290] = layer0_outputs[4541];
    assign outputs[1291] = ~(layer0_outputs[6545]);
    assign outputs[1292] = (layer0_outputs[4515]) & ~(layer0_outputs[1106]);
    assign outputs[1293] = (layer0_outputs[4273]) & ~(layer0_outputs[5189]);
    assign outputs[1294] = ~(layer0_outputs[893]);
    assign outputs[1295] = (layer0_outputs[6549]) & ~(layer0_outputs[4738]);
    assign outputs[1296] = (layer0_outputs[6988]) ^ (layer0_outputs[3564]);
    assign outputs[1297] = layer0_outputs[3182];
    assign outputs[1298] = ~((layer0_outputs[4173]) ^ (layer0_outputs[3353]));
    assign outputs[1299] = ~((layer0_outputs[4442]) | (layer0_outputs[5948]));
    assign outputs[1300] = (layer0_outputs[3839]) & ~(layer0_outputs[6626]);
    assign outputs[1301] = layer0_outputs[6025];
    assign outputs[1302] = ~(layer0_outputs[7590]);
    assign outputs[1303] = (layer0_outputs[812]) & (layer0_outputs[1832]);
    assign outputs[1304] = (layer0_outputs[4085]) & ~(layer0_outputs[6597]);
    assign outputs[1305] = (layer0_outputs[6677]) & ~(layer0_outputs[2502]);
    assign outputs[1306] = (layer0_outputs[4004]) & ~(layer0_outputs[2448]);
    assign outputs[1307] = ~(layer0_outputs[2378]);
    assign outputs[1308] = (layer0_outputs[5963]) & ~(layer0_outputs[7075]);
    assign outputs[1309] = 1'b0;
    assign outputs[1310] = (layer0_outputs[6353]) & ~(layer0_outputs[699]);
    assign outputs[1311] = layer0_outputs[6159];
    assign outputs[1312] = (layer0_outputs[3965]) & ~(layer0_outputs[1169]);
    assign outputs[1313] = 1'b0;
    assign outputs[1314] = (layer0_outputs[187]) ^ (layer0_outputs[6468]);
    assign outputs[1315] = 1'b0;
    assign outputs[1316] = layer0_outputs[4912];
    assign outputs[1317] = layer0_outputs[5347];
    assign outputs[1318] = ~((layer0_outputs[6330]) | (layer0_outputs[7537]));
    assign outputs[1319] = (layer0_outputs[173]) & ~(layer0_outputs[5779]);
    assign outputs[1320] = layer0_outputs[1859];
    assign outputs[1321] = (layer0_outputs[2932]) & ~(layer0_outputs[5899]);
    assign outputs[1322] = ~(layer0_outputs[2641]);
    assign outputs[1323] = 1'b0;
    assign outputs[1324] = ~((layer0_outputs[5843]) ^ (layer0_outputs[1110]));
    assign outputs[1325] = ~(layer0_outputs[1333]);
    assign outputs[1326] = (layer0_outputs[1080]) & ~(layer0_outputs[7275]);
    assign outputs[1327] = (layer0_outputs[3963]) & (layer0_outputs[986]);
    assign outputs[1328] = 1'b0;
    assign outputs[1329] = ~(layer0_outputs[3512]);
    assign outputs[1330] = layer0_outputs[1971];
    assign outputs[1331] = ~(layer0_outputs[137]);
    assign outputs[1332] = (layer0_outputs[3971]) & ~(layer0_outputs[7203]);
    assign outputs[1333] = (layer0_outputs[94]) ^ (layer0_outputs[753]);
    assign outputs[1334] = ~(layer0_outputs[2396]);
    assign outputs[1335] = (layer0_outputs[5556]) & ~(layer0_outputs[4740]);
    assign outputs[1336] = ~((layer0_outputs[5367]) ^ (layer0_outputs[6949]));
    assign outputs[1337] = ~((layer0_outputs[5872]) ^ (layer0_outputs[5272]));
    assign outputs[1338] = layer0_outputs[5704];
    assign outputs[1339] = layer0_outputs[2529];
    assign outputs[1340] = (layer0_outputs[6937]) & (layer0_outputs[947]);
    assign outputs[1341] = ~((layer0_outputs[1046]) | (layer0_outputs[6801]));
    assign outputs[1342] = (layer0_outputs[4868]) & (layer0_outputs[4484]);
    assign outputs[1343] = (layer0_outputs[2512]) & ~(layer0_outputs[6328]);
    assign outputs[1344] = ~((layer0_outputs[5630]) | (layer0_outputs[1049]));
    assign outputs[1345] = (layer0_outputs[1415]) & (layer0_outputs[2418]);
    assign outputs[1346] = (layer0_outputs[3540]) & ~(layer0_outputs[3451]);
    assign outputs[1347] = ~((layer0_outputs[2471]) | (layer0_outputs[4806]));
    assign outputs[1348] = (layer0_outputs[3937]) & ~(layer0_outputs[6522]);
    assign outputs[1349] = 1'b0;
    assign outputs[1350] = (layer0_outputs[734]) & ~(layer0_outputs[6135]);
    assign outputs[1351] = (layer0_outputs[6433]) & (layer0_outputs[6762]);
    assign outputs[1352] = (layer0_outputs[2727]) & (layer0_outputs[103]);
    assign outputs[1353] = ~(layer0_outputs[7286]);
    assign outputs[1354] = (layer0_outputs[2095]) & ~(layer0_outputs[4292]);
    assign outputs[1355] = (layer0_outputs[3983]) & (layer0_outputs[4602]);
    assign outputs[1356] = ~((layer0_outputs[809]) | (layer0_outputs[7361]));
    assign outputs[1357] = (layer0_outputs[1572]) ^ (layer0_outputs[2779]);
    assign outputs[1358] = layer0_outputs[670];
    assign outputs[1359] = ~(layer0_outputs[704]);
    assign outputs[1360] = (layer0_outputs[1466]) & ~(layer0_outputs[1432]);
    assign outputs[1361] = layer0_outputs[6667];
    assign outputs[1362] = (layer0_outputs[3723]) & ~(layer0_outputs[2098]);
    assign outputs[1363] = (layer0_outputs[987]) | (layer0_outputs[1271]);
    assign outputs[1364] = 1'b0;
    assign outputs[1365] = ~((layer0_outputs[1225]) | (layer0_outputs[3745]));
    assign outputs[1366] = ~(layer0_outputs[1111]);
    assign outputs[1367] = (layer0_outputs[3041]) ^ (layer0_outputs[5706]);
    assign outputs[1368] = ~(layer0_outputs[1803]);
    assign outputs[1369] = 1'b0;
    assign outputs[1370] = (layer0_outputs[2826]) & (layer0_outputs[2170]);
    assign outputs[1371] = layer0_outputs[4930];
    assign outputs[1372] = layer0_outputs[3079];
    assign outputs[1373] = (layer0_outputs[3985]) & ~(layer0_outputs[1956]);
    assign outputs[1374] = (layer0_outputs[7076]) & ~(layer0_outputs[2745]);
    assign outputs[1375] = ~((layer0_outputs[249]) | (layer0_outputs[3669]));
    assign outputs[1376] = layer0_outputs[2189];
    assign outputs[1377] = layer0_outputs[3555];
    assign outputs[1378] = ~(layer0_outputs[44]);
    assign outputs[1379] = (layer0_outputs[32]) & ~(layer0_outputs[7425]);
    assign outputs[1380] = (layer0_outputs[4954]) & ~(layer0_outputs[4964]);
    assign outputs[1381] = (layer0_outputs[4447]) & ~(layer0_outputs[5162]);
    assign outputs[1382] = (layer0_outputs[5178]) & (layer0_outputs[1711]);
    assign outputs[1383] = layer0_outputs[5837];
    assign outputs[1384] = (layer0_outputs[3562]) & (layer0_outputs[2607]);
    assign outputs[1385] = ~(layer0_outputs[2586]);
    assign outputs[1386] = ~(layer0_outputs[5034]);
    assign outputs[1387] = (layer0_outputs[1083]) & ~(layer0_outputs[5961]);
    assign outputs[1388] = layer0_outputs[2531];
    assign outputs[1389] = ~(layer0_outputs[2702]);
    assign outputs[1390] = ~(layer0_outputs[2637]) | (layer0_outputs[6419]);
    assign outputs[1391] = layer0_outputs[1137];
    assign outputs[1392] = (layer0_outputs[2736]) ^ (layer0_outputs[1407]);
    assign outputs[1393] = ~((layer0_outputs[3724]) ^ (layer0_outputs[4392]));
    assign outputs[1394] = (layer0_outputs[5333]) & ~(layer0_outputs[1534]);
    assign outputs[1395] = (layer0_outputs[1762]) & ~(layer0_outputs[2630]);
    assign outputs[1396] = ~((layer0_outputs[5898]) | (layer0_outputs[2967]));
    assign outputs[1397] = (layer0_outputs[6981]) & (layer0_outputs[904]);
    assign outputs[1398] = (layer0_outputs[3532]) ^ (layer0_outputs[3918]);
    assign outputs[1399] = (layer0_outputs[4441]) & (layer0_outputs[652]);
    assign outputs[1400] = ~(layer0_outputs[56]);
    assign outputs[1401] = layer0_outputs[4903];
    assign outputs[1402] = layer0_outputs[5781];
    assign outputs[1403] = ~(layer0_outputs[140]);
    assign outputs[1404] = ~(layer0_outputs[1266]);
    assign outputs[1405] = (layer0_outputs[5107]) ^ (layer0_outputs[4561]);
    assign outputs[1406] = layer0_outputs[4863];
    assign outputs[1407] = (layer0_outputs[6448]) & ~(layer0_outputs[4503]);
    assign outputs[1408] = (layer0_outputs[7277]) & (layer0_outputs[2825]);
    assign outputs[1409] = (layer0_outputs[478]) ^ (layer0_outputs[3658]);
    assign outputs[1410] = (layer0_outputs[7390]) & ~(layer0_outputs[2987]);
    assign outputs[1411] = ~(layer0_outputs[3675]);
    assign outputs[1412] = ~((layer0_outputs[2173]) | (layer0_outputs[4351]));
    assign outputs[1413] = ~((layer0_outputs[455]) | (layer0_outputs[108]));
    assign outputs[1414] = layer0_outputs[4169];
    assign outputs[1415] = (layer0_outputs[5791]) ^ (layer0_outputs[6092]);
    assign outputs[1416] = (layer0_outputs[5042]) & ~(layer0_outputs[6611]);
    assign outputs[1417] = layer0_outputs[1783];
    assign outputs[1418] = ~((layer0_outputs[5342]) ^ (layer0_outputs[2075]));
    assign outputs[1419] = ~((layer0_outputs[283]) | (layer0_outputs[6083]));
    assign outputs[1420] = ~(layer0_outputs[7018]);
    assign outputs[1421] = (layer0_outputs[579]) & ~(layer0_outputs[4524]);
    assign outputs[1422] = layer0_outputs[3209];
    assign outputs[1423] = (layer0_outputs[6590]) & ~(layer0_outputs[5399]);
    assign outputs[1424] = ~(layer0_outputs[218]);
    assign outputs[1425] = ~((layer0_outputs[1103]) | (layer0_outputs[6840]));
    assign outputs[1426] = ~((layer0_outputs[1848]) ^ (layer0_outputs[1899]));
    assign outputs[1427] = ~(layer0_outputs[4819]);
    assign outputs[1428] = layer0_outputs[3139];
    assign outputs[1429] = layer0_outputs[3883];
    assign outputs[1430] = ~(layer0_outputs[4551]) | (layer0_outputs[1252]);
    assign outputs[1431] = ~((layer0_outputs[6385]) | (layer0_outputs[1381]));
    assign outputs[1432] = (layer0_outputs[2275]) & ~(layer0_outputs[6150]);
    assign outputs[1433] = ~((layer0_outputs[7044]) | (layer0_outputs[6080]));
    assign outputs[1434] = (layer0_outputs[7218]) & ~(layer0_outputs[3427]);
    assign outputs[1435] = (layer0_outputs[5960]) & ~(layer0_outputs[37]);
    assign outputs[1436] = ~((layer0_outputs[7227]) | (layer0_outputs[6654]));
    assign outputs[1437] = layer0_outputs[6754];
    assign outputs[1438] = ~((layer0_outputs[1958]) ^ (layer0_outputs[6835]));
    assign outputs[1439] = layer0_outputs[2677];
    assign outputs[1440] = (layer0_outputs[743]) & ~(layer0_outputs[6046]);
    assign outputs[1441] = ~((layer0_outputs[282]) & (layer0_outputs[4900]));
    assign outputs[1442] = ~(layer0_outputs[2370]) | (layer0_outputs[1301]);
    assign outputs[1443] = (layer0_outputs[5020]) & ~(layer0_outputs[1277]);
    assign outputs[1444] = ~(layer0_outputs[502]);
    assign outputs[1445] = (layer0_outputs[5347]) & ~(layer0_outputs[6385]);
    assign outputs[1446] = (layer0_outputs[604]) & ~(layer0_outputs[927]);
    assign outputs[1447] = ~(layer0_outputs[4653]);
    assign outputs[1448] = (layer0_outputs[4727]) & ~(layer0_outputs[3284]);
    assign outputs[1449] = (layer0_outputs[5828]) ^ (layer0_outputs[1287]);
    assign outputs[1450] = (layer0_outputs[4756]) & (layer0_outputs[1201]);
    assign outputs[1451] = ~(layer0_outputs[6328]);
    assign outputs[1452] = ~(layer0_outputs[7611]);
    assign outputs[1453] = (layer0_outputs[2873]) & (layer0_outputs[7187]);
    assign outputs[1454] = (layer0_outputs[1220]) & ~(layer0_outputs[6836]);
    assign outputs[1455] = (layer0_outputs[3195]) & (layer0_outputs[6345]);
    assign outputs[1456] = layer0_outputs[5574];
    assign outputs[1457] = (layer0_outputs[5685]) & ~(layer0_outputs[3760]);
    assign outputs[1458] = ~(layer0_outputs[2992]);
    assign outputs[1459] = (layer0_outputs[6331]) & ~(layer0_outputs[5971]);
    assign outputs[1460] = (layer0_outputs[3438]) ^ (layer0_outputs[6399]);
    assign outputs[1461] = (layer0_outputs[291]) & ~(layer0_outputs[2965]);
    assign outputs[1462] = layer0_outputs[7655];
    assign outputs[1463] = (layer0_outputs[5577]) ^ (layer0_outputs[5227]);
    assign outputs[1464] = (layer0_outputs[7538]) & ~(layer0_outputs[3350]);
    assign outputs[1465] = (layer0_outputs[1038]) & ~(layer0_outputs[6425]);
    assign outputs[1466] = (layer0_outputs[4314]) & ~(layer0_outputs[5237]);
    assign outputs[1467] = 1'b0;
    assign outputs[1468] = (layer0_outputs[1150]) & (layer0_outputs[4483]);
    assign outputs[1469] = (layer0_outputs[403]) & ~(layer0_outputs[744]);
    assign outputs[1470] = ~(layer0_outputs[122]);
    assign outputs[1471] = (layer0_outputs[3188]) & (layer0_outputs[2426]);
    assign outputs[1472] = (layer0_outputs[3695]) & ~(layer0_outputs[3219]);
    assign outputs[1473] = layer0_outputs[7564];
    assign outputs[1474] = (layer0_outputs[4051]) & ~(layer0_outputs[4078]);
    assign outputs[1475] = (layer0_outputs[1476]) & (layer0_outputs[4067]);
    assign outputs[1476] = layer0_outputs[6148];
    assign outputs[1477] = layer0_outputs[7556];
    assign outputs[1478] = ~((layer0_outputs[631]) ^ (layer0_outputs[4465]));
    assign outputs[1479] = ~(layer0_outputs[2460]) | (layer0_outputs[1234]);
    assign outputs[1480] = 1'b0;
    assign outputs[1481] = (layer0_outputs[6898]) & ~(layer0_outputs[1108]);
    assign outputs[1482] = (layer0_outputs[3550]) & ~(layer0_outputs[327]);
    assign outputs[1483] = (layer0_outputs[49]) ^ (layer0_outputs[4109]);
    assign outputs[1484] = (layer0_outputs[845]) ^ (layer0_outputs[5175]);
    assign outputs[1485] = (layer0_outputs[6214]) & ~(layer0_outputs[7028]);
    assign outputs[1486] = (layer0_outputs[6525]) & (layer0_outputs[6412]);
    assign outputs[1487] = ~(layer0_outputs[5152]);
    assign outputs[1488] = ~((layer0_outputs[1804]) ^ (layer0_outputs[4850]));
    assign outputs[1489] = (layer0_outputs[6407]) ^ (layer0_outputs[1060]);
    assign outputs[1490] = layer0_outputs[1235];
    assign outputs[1491] = (layer0_outputs[5398]) & ~(layer0_outputs[1052]);
    assign outputs[1492] = ~(layer0_outputs[6317]);
    assign outputs[1493] = (layer0_outputs[1187]) & (layer0_outputs[2938]);
    assign outputs[1494] = (layer0_outputs[4130]) & (layer0_outputs[3294]);
    assign outputs[1495] = (layer0_outputs[4557]) ^ (layer0_outputs[2063]);
    assign outputs[1496] = (layer0_outputs[3840]) ^ (layer0_outputs[875]);
    assign outputs[1497] = layer0_outputs[1712];
    assign outputs[1498] = ~((layer0_outputs[6847]) | (layer0_outputs[5021]));
    assign outputs[1499] = (layer0_outputs[842]) & ~(layer0_outputs[5239]);
    assign outputs[1500] = (layer0_outputs[3378]) & (layer0_outputs[1352]);
    assign outputs[1501] = (layer0_outputs[2600]) ^ (layer0_outputs[1465]);
    assign outputs[1502] = (layer0_outputs[1837]) & (layer0_outputs[1660]);
    assign outputs[1503] = (layer0_outputs[1071]) | (layer0_outputs[5510]);
    assign outputs[1504] = layer0_outputs[6185];
    assign outputs[1505] = layer0_outputs[3353];
    assign outputs[1506] = (layer0_outputs[5164]) & (layer0_outputs[4360]);
    assign outputs[1507] = (layer0_outputs[7382]) & ~(layer0_outputs[6075]);
    assign outputs[1508] = (layer0_outputs[436]) & ~(layer0_outputs[321]);
    assign outputs[1509] = ~((layer0_outputs[1893]) ^ (layer0_outputs[6280]));
    assign outputs[1510] = (layer0_outputs[4599]) & ~(layer0_outputs[3400]);
    assign outputs[1511] = ~(layer0_outputs[2039]);
    assign outputs[1512] = (layer0_outputs[2521]) & ~(layer0_outputs[5891]);
    assign outputs[1513] = (layer0_outputs[6060]) & ~(layer0_outputs[732]);
    assign outputs[1514] = layer0_outputs[6616];
    assign outputs[1515] = (layer0_outputs[1921]) ^ (layer0_outputs[6048]);
    assign outputs[1516] = ~((layer0_outputs[2153]) | (layer0_outputs[4202]));
    assign outputs[1517] = layer0_outputs[7396];
    assign outputs[1518] = (layer0_outputs[2393]) & ~(layer0_outputs[3518]);
    assign outputs[1519] = (layer0_outputs[721]) ^ (layer0_outputs[6741]);
    assign outputs[1520] = ~(layer0_outputs[6049]);
    assign outputs[1521] = (layer0_outputs[1729]) & (layer0_outputs[3123]);
    assign outputs[1522] = ~((layer0_outputs[2372]) ^ (layer0_outputs[3036]));
    assign outputs[1523] = 1'b0;
    assign outputs[1524] = (layer0_outputs[5190]) & ~(layer0_outputs[6659]);
    assign outputs[1525] = ~(layer0_outputs[7030]);
    assign outputs[1526] = (layer0_outputs[590]) & ~(layer0_outputs[318]);
    assign outputs[1527] = (layer0_outputs[752]) & ~(layer0_outputs[3569]);
    assign outputs[1528] = ~((layer0_outputs[4608]) & (layer0_outputs[4772]));
    assign outputs[1529] = (layer0_outputs[5500]) & (layer0_outputs[5181]);
    assign outputs[1530] = layer0_outputs[1783];
    assign outputs[1531] = (layer0_outputs[5878]) ^ (layer0_outputs[5112]);
    assign outputs[1532] = (layer0_outputs[2557]) ^ (layer0_outputs[3277]);
    assign outputs[1533] = layer0_outputs[6540];
    assign outputs[1534] = ~(layer0_outputs[1592]);
    assign outputs[1535] = ~((layer0_outputs[3844]) ^ (layer0_outputs[4025]));
    assign outputs[1536] = ~(layer0_outputs[911]) | (layer0_outputs[5601]);
    assign outputs[1537] = ~(layer0_outputs[7309]);
    assign outputs[1538] = ~((layer0_outputs[7065]) ^ (layer0_outputs[276]));
    assign outputs[1539] = layer0_outputs[4497];
    assign outputs[1540] = layer0_outputs[5928];
    assign outputs[1541] = 1'b1;
    assign outputs[1542] = (layer0_outputs[6555]) | (layer0_outputs[3921]);
    assign outputs[1543] = ~(layer0_outputs[445]);
    assign outputs[1544] = ~(layer0_outputs[1097]);
    assign outputs[1545] = layer0_outputs[1874];
    assign outputs[1546] = ~((layer0_outputs[6483]) & (layer0_outputs[6306]));
    assign outputs[1547] = layer0_outputs[2151];
    assign outputs[1548] = (layer0_outputs[2762]) ^ (layer0_outputs[2829]);
    assign outputs[1549] = layer0_outputs[7257];
    assign outputs[1550] = (layer0_outputs[2795]) & ~(layer0_outputs[6442]);
    assign outputs[1551] = ~(layer0_outputs[6052]);
    assign outputs[1552] = (layer0_outputs[1937]) ^ (layer0_outputs[7629]);
    assign outputs[1553] = ~(layer0_outputs[6374]);
    assign outputs[1554] = layer0_outputs[1405];
    assign outputs[1555] = (layer0_outputs[830]) ^ (layer0_outputs[293]);
    assign outputs[1556] = layer0_outputs[1685];
    assign outputs[1557] = ~((layer0_outputs[6853]) & (layer0_outputs[6825]));
    assign outputs[1558] = ~(layer0_outputs[5732]);
    assign outputs[1559] = ~((layer0_outputs[3626]) ^ (layer0_outputs[4028]));
    assign outputs[1560] = ~(layer0_outputs[5224]);
    assign outputs[1561] = (layer0_outputs[2367]) | (layer0_outputs[829]);
    assign outputs[1562] = ~(layer0_outputs[3807]);
    assign outputs[1563] = layer0_outputs[6206];
    assign outputs[1564] = ~((layer0_outputs[100]) | (layer0_outputs[2935]));
    assign outputs[1565] = (layer0_outputs[3366]) & ~(layer0_outputs[5240]);
    assign outputs[1566] = (layer0_outputs[6267]) & ~(layer0_outputs[4641]);
    assign outputs[1567] = (layer0_outputs[3317]) ^ (layer0_outputs[1585]);
    assign outputs[1568] = (layer0_outputs[5757]) | (layer0_outputs[5758]);
    assign outputs[1569] = (layer0_outputs[484]) | (layer0_outputs[6015]);
    assign outputs[1570] = ~(layer0_outputs[2378]) | (layer0_outputs[278]);
    assign outputs[1571] = ~((layer0_outputs[7624]) & (layer0_outputs[5300]));
    assign outputs[1572] = (layer0_outputs[5625]) ^ (layer0_outputs[2353]);
    assign outputs[1573] = ~(layer0_outputs[1876]) | (layer0_outputs[3748]);
    assign outputs[1574] = layer0_outputs[2509];
    assign outputs[1575] = ~(layer0_outputs[2061]) | (layer0_outputs[3669]);
    assign outputs[1576] = ~((layer0_outputs[1693]) ^ (layer0_outputs[3414]));
    assign outputs[1577] = ~(layer0_outputs[2256]);
    assign outputs[1578] = (layer0_outputs[611]) & ~(layer0_outputs[90]);
    assign outputs[1579] = ~(layer0_outputs[4314]) | (layer0_outputs[1200]);
    assign outputs[1580] = ~((layer0_outputs[5587]) ^ (layer0_outputs[7149]));
    assign outputs[1581] = ~(layer0_outputs[5753]) | (layer0_outputs[3744]);
    assign outputs[1582] = ~(layer0_outputs[5467]);
    assign outputs[1583] = (layer0_outputs[1034]) | (layer0_outputs[4145]);
    assign outputs[1584] = layer0_outputs[5513];
    assign outputs[1585] = ~(layer0_outputs[2676]);
    assign outputs[1586] = (layer0_outputs[7674]) & ~(layer0_outputs[1545]);
    assign outputs[1587] = (layer0_outputs[6010]) & (layer0_outputs[3608]);
    assign outputs[1588] = ~((layer0_outputs[118]) & (layer0_outputs[176]));
    assign outputs[1589] = ~((layer0_outputs[5066]) & (layer0_outputs[4352]));
    assign outputs[1590] = ~(layer0_outputs[3071]);
    assign outputs[1591] = ~(layer0_outputs[4557]);
    assign outputs[1592] = ~((layer0_outputs[3283]) ^ (layer0_outputs[1005]));
    assign outputs[1593] = (layer0_outputs[3670]) ^ (layer0_outputs[5628]);
    assign outputs[1594] = ~(layer0_outputs[2203]) | (layer0_outputs[6749]);
    assign outputs[1595] = layer0_outputs[407];
    assign outputs[1596] = (layer0_outputs[2085]) ^ (layer0_outputs[5139]);
    assign outputs[1597] = ~(layer0_outputs[6424]);
    assign outputs[1598] = layer0_outputs[2671];
    assign outputs[1599] = ~(layer0_outputs[4021]) | (layer0_outputs[1167]);
    assign outputs[1600] = (layer0_outputs[7445]) ^ (layer0_outputs[7453]);
    assign outputs[1601] = ~((layer0_outputs[6874]) ^ (layer0_outputs[7407]));
    assign outputs[1602] = layer0_outputs[6227];
    assign outputs[1603] = (layer0_outputs[2506]) & (layer0_outputs[3594]);
    assign outputs[1604] = (layer0_outputs[493]) & ~(layer0_outputs[7014]);
    assign outputs[1605] = ~((layer0_outputs[5435]) | (layer0_outputs[1153]));
    assign outputs[1606] = (layer0_outputs[2711]) ^ (layer0_outputs[7647]);
    assign outputs[1607] = ~(layer0_outputs[4950]) | (layer0_outputs[1690]);
    assign outputs[1608] = ~(layer0_outputs[4752]);
    assign outputs[1609] = ~((layer0_outputs[6188]) ^ (layer0_outputs[4616]));
    assign outputs[1610] = ~(layer0_outputs[1708]);
    assign outputs[1611] = ~(layer0_outputs[3049]);
    assign outputs[1612] = (layer0_outputs[3994]) ^ (layer0_outputs[5329]);
    assign outputs[1613] = (layer0_outputs[3408]) ^ (layer0_outputs[6084]);
    assign outputs[1614] = ~(layer0_outputs[1667]);
    assign outputs[1615] = ~(layer0_outputs[2380]);
    assign outputs[1616] = layer0_outputs[4966];
    assign outputs[1617] = (layer0_outputs[665]) & ~(layer0_outputs[3693]);
    assign outputs[1618] = ~(layer0_outputs[1926]);
    assign outputs[1619] = layer0_outputs[3197];
    assign outputs[1620] = layer0_outputs[6274];
    assign outputs[1621] = ~((layer0_outputs[3842]) ^ (layer0_outputs[6542]));
    assign outputs[1622] = (layer0_outputs[65]) & (layer0_outputs[936]);
    assign outputs[1623] = layer0_outputs[2421];
    assign outputs[1624] = ~(layer0_outputs[7323]) | (layer0_outputs[2467]);
    assign outputs[1625] = ~(layer0_outputs[5675]);
    assign outputs[1626] = ~(layer0_outputs[2059]) | (layer0_outputs[2810]);
    assign outputs[1627] = ~((layer0_outputs[4206]) ^ (layer0_outputs[6417]));
    assign outputs[1628] = ~(layer0_outputs[6562]);
    assign outputs[1629] = ~(layer0_outputs[6844]) | (layer0_outputs[3729]);
    assign outputs[1630] = layer0_outputs[1244];
    assign outputs[1631] = ~(layer0_outputs[5159]) | (layer0_outputs[2554]);
    assign outputs[1632] = layer0_outputs[3384];
    assign outputs[1633] = layer0_outputs[6458];
    assign outputs[1634] = ~(layer0_outputs[362]);
    assign outputs[1635] = (layer0_outputs[3192]) & ~(layer0_outputs[55]);
    assign outputs[1636] = ~((layer0_outputs[3898]) & (layer0_outputs[4802]));
    assign outputs[1637] = ~((layer0_outputs[3736]) & (layer0_outputs[5531]));
    assign outputs[1638] = layer0_outputs[7158];
    assign outputs[1639] = ~(layer0_outputs[1855]);
    assign outputs[1640] = layer0_outputs[717];
    assign outputs[1641] = ~((layer0_outputs[6012]) & (layer0_outputs[3510]));
    assign outputs[1642] = ~(layer0_outputs[1133]) | (layer0_outputs[565]);
    assign outputs[1643] = ~(layer0_outputs[2040]);
    assign outputs[1644] = ~((layer0_outputs[4333]) & (layer0_outputs[6155]));
    assign outputs[1645] = ~((layer0_outputs[7631]) & (layer0_outputs[4848]));
    assign outputs[1646] = ~((layer0_outputs[6789]) ^ (layer0_outputs[3399]));
    assign outputs[1647] = ~(layer0_outputs[550]);
    assign outputs[1648] = (layer0_outputs[1856]) & (layer0_outputs[4393]);
    assign outputs[1649] = layer0_outputs[3121];
    assign outputs[1650] = ~(layer0_outputs[2818]);
    assign outputs[1651] = (layer0_outputs[523]) ^ (layer0_outputs[5772]);
    assign outputs[1652] = ~(layer0_outputs[3480]);
    assign outputs[1653] = (layer0_outputs[6662]) & ~(layer0_outputs[2843]);
    assign outputs[1654] = ~(layer0_outputs[1530]);
    assign outputs[1655] = (layer0_outputs[2944]) ^ (layer0_outputs[1126]);
    assign outputs[1656] = ~(layer0_outputs[7142]) | (layer0_outputs[6967]);
    assign outputs[1657] = layer0_outputs[7437];
    assign outputs[1658] = layer0_outputs[201];
    assign outputs[1659] = ~(layer0_outputs[2210]) | (layer0_outputs[5695]);
    assign outputs[1660] = layer0_outputs[2371];
    assign outputs[1661] = layer0_outputs[4115];
    assign outputs[1662] = (layer0_outputs[4812]) ^ (layer0_outputs[6144]);
    assign outputs[1663] = ~((layer0_outputs[1846]) & (layer0_outputs[3915]));
    assign outputs[1664] = 1'b1;
    assign outputs[1665] = layer0_outputs[5170];
    assign outputs[1666] = (layer0_outputs[2184]) ^ (layer0_outputs[3773]);
    assign outputs[1667] = ~(layer0_outputs[1140]) | (layer0_outputs[3475]);
    assign outputs[1668] = ~(layer0_outputs[6736]);
    assign outputs[1669] = layer0_outputs[6022];
    assign outputs[1670] = ~(layer0_outputs[6552]);
    assign outputs[1671] = ~((layer0_outputs[4413]) ^ (layer0_outputs[4416]));
    assign outputs[1672] = ~(layer0_outputs[7554]);
    assign outputs[1673] = ~(layer0_outputs[2943]);
    assign outputs[1674] = (layer0_outputs[2480]) & ~(layer0_outputs[1316]);
    assign outputs[1675] = layer0_outputs[4959];
    assign outputs[1676] = ~(layer0_outputs[4002]);
    assign outputs[1677] = ~((layer0_outputs[6078]) ^ (layer0_outputs[3016]));
    assign outputs[1678] = ~(layer0_outputs[6689]) | (layer0_outputs[2937]);
    assign outputs[1679] = 1'b1;
    assign outputs[1680] = ~((layer0_outputs[2006]) & (layer0_outputs[5173]));
    assign outputs[1681] = ~((layer0_outputs[1969]) ^ (layer0_outputs[1377]));
    assign outputs[1682] = ~(layer0_outputs[7146]);
    assign outputs[1683] = ~(layer0_outputs[3262]) | (layer0_outputs[3028]);
    assign outputs[1684] = ~((layer0_outputs[3443]) | (layer0_outputs[6463]));
    assign outputs[1685] = ~(layer0_outputs[7296]) | (layer0_outputs[6826]);
    assign outputs[1686] = ~(layer0_outputs[1659]);
    assign outputs[1687] = (layer0_outputs[3613]) | (layer0_outputs[3081]);
    assign outputs[1688] = (layer0_outputs[176]) ^ (layer0_outputs[1081]);
    assign outputs[1689] = ~(layer0_outputs[4254]) | (layer0_outputs[6880]);
    assign outputs[1690] = ~(layer0_outputs[2959]);
    assign outputs[1691] = ~(layer0_outputs[3962]);
    assign outputs[1692] = (layer0_outputs[5738]) ^ (layer0_outputs[379]);
    assign outputs[1693] = layer0_outputs[7518];
    assign outputs[1694] = (layer0_outputs[6491]) & ~(layer0_outputs[4653]);
    assign outputs[1695] = (layer0_outputs[3522]) | (layer0_outputs[5966]);
    assign outputs[1696] = layer0_outputs[4650];
    assign outputs[1697] = ~(layer0_outputs[6246]);
    assign outputs[1698] = ~(layer0_outputs[274]);
    assign outputs[1699] = (layer0_outputs[574]) ^ (layer0_outputs[3365]);
    assign outputs[1700] = ~((layer0_outputs[4124]) & (layer0_outputs[4143]));
    assign outputs[1701] = ~((layer0_outputs[5026]) & (layer0_outputs[3316]));
    assign outputs[1702] = layer0_outputs[2830];
    assign outputs[1703] = ~((layer0_outputs[6947]) & (layer0_outputs[1018]));
    assign outputs[1704] = ~(layer0_outputs[2594]);
    assign outputs[1705] = ~((layer0_outputs[2299]) ^ (layer0_outputs[1715]));
    assign outputs[1706] = layer0_outputs[2893];
    assign outputs[1707] = ~((layer0_outputs[4719]) ^ (layer0_outputs[1680]));
    assign outputs[1708] = layer0_outputs[3147];
    assign outputs[1709] = ~(layer0_outputs[4343]);
    assign outputs[1710] = ~(layer0_outputs[7191]) | (layer0_outputs[3780]);
    assign outputs[1711] = layer0_outputs[7136];
    assign outputs[1712] = layer0_outputs[964];
    assign outputs[1713] = (layer0_outputs[4374]) & (layer0_outputs[5185]);
    assign outputs[1714] = ~(layer0_outputs[6778]) | (layer0_outputs[4474]);
    assign outputs[1715] = ~((layer0_outputs[3811]) ^ (layer0_outputs[1699]));
    assign outputs[1716] = ~(layer0_outputs[6376]) | (layer0_outputs[523]);
    assign outputs[1717] = ~(layer0_outputs[532]);
    assign outputs[1718] = layer0_outputs[4332];
    assign outputs[1719] = layer0_outputs[3841];
    assign outputs[1720] = ~(layer0_outputs[1436]);
    assign outputs[1721] = ~(layer0_outputs[3691]);
    assign outputs[1722] = ~((layer0_outputs[257]) ^ (layer0_outputs[4512]));
    assign outputs[1723] = layer0_outputs[692];
    assign outputs[1724] = ~(layer0_outputs[7053]);
    assign outputs[1725] = layer0_outputs[5679];
    assign outputs[1726] = (layer0_outputs[7567]) & ~(layer0_outputs[3058]);
    assign outputs[1727] = layer0_outputs[6455];
    assign outputs[1728] = ~(layer0_outputs[6857]);
    assign outputs[1729] = layer0_outputs[5050];
    assign outputs[1730] = ~(layer0_outputs[757]);
    assign outputs[1731] = ~(layer0_outputs[5426]);
    assign outputs[1732] = layer0_outputs[6886];
    assign outputs[1733] = ~(layer0_outputs[1083]) | (layer0_outputs[5012]);
    assign outputs[1734] = ~((layer0_outputs[4936]) | (layer0_outputs[6158]));
    assign outputs[1735] = (layer0_outputs[3180]) ^ (layer0_outputs[5989]);
    assign outputs[1736] = (layer0_outputs[5182]) | (layer0_outputs[6376]);
    assign outputs[1737] = ~(layer0_outputs[4213]);
    assign outputs[1738] = ~(layer0_outputs[149]);
    assign outputs[1739] = ~(layer0_outputs[2797]) | (layer0_outputs[4648]);
    assign outputs[1740] = ~((layer0_outputs[3021]) ^ (layer0_outputs[6409]));
    assign outputs[1741] = ~((layer0_outputs[6486]) ^ (layer0_outputs[4176]));
    assign outputs[1742] = ~(layer0_outputs[1363]) | (layer0_outputs[4867]);
    assign outputs[1743] = layer0_outputs[6967];
    assign outputs[1744] = ~((layer0_outputs[5966]) ^ (layer0_outputs[5415]));
    assign outputs[1745] = layer0_outputs[2548];
    assign outputs[1746] = ~((layer0_outputs[1719]) ^ (layer0_outputs[6846]));
    assign outputs[1747] = layer0_outputs[7499];
    assign outputs[1748] = ~(layer0_outputs[3756]);
    assign outputs[1749] = (layer0_outputs[6116]) | (layer0_outputs[5748]);
    assign outputs[1750] = (layer0_outputs[4676]) & (layer0_outputs[964]);
    assign outputs[1751] = ~((layer0_outputs[4890]) & (layer0_outputs[891]));
    assign outputs[1752] = layer0_outputs[2069];
    assign outputs[1753] = ~(layer0_outputs[5405]);
    assign outputs[1754] = layer0_outputs[5265];
    assign outputs[1755] = ~(layer0_outputs[4824]);
    assign outputs[1756] = ~(layer0_outputs[2641]);
    assign outputs[1757] = (layer0_outputs[2137]) & (layer0_outputs[747]);
    assign outputs[1758] = ~(layer0_outputs[5923]);
    assign outputs[1759] = layer0_outputs[220];
    assign outputs[1760] = (layer0_outputs[4285]) & ~(layer0_outputs[7635]);
    assign outputs[1761] = ~(layer0_outputs[5161]);
    assign outputs[1762] = (layer0_outputs[2810]) & ~(layer0_outputs[6299]);
    assign outputs[1763] = 1'b1;
    assign outputs[1764] = ~(layer0_outputs[6752]);
    assign outputs[1765] = ~(layer0_outputs[5581]);
    assign outputs[1766] = ~(layer0_outputs[3249]);
    assign outputs[1767] = (layer0_outputs[3863]) & (layer0_outputs[5802]);
    assign outputs[1768] = ~((layer0_outputs[1557]) | (layer0_outputs[7172]));
    assign outputs[1769] = layer0_outputs[7108];
    assign outputs[1770] = ~(layer0_outputs[5195]) | (layer0_outputs[7019]);
    assign outputs[1771] = ~(layer0_outputs[3018]) | (layer0_outputs[6615]);
    assign outputs[1772] = ~(layer0_outputs[6480]) | (layer0_outputs[2671]);
    assign outputs[1773] = ~(layer0_outputs[1312]);
    assign outputs[1774] = ~((layer0_outputs[4895]) | (layer0_outputs[5668]));
    assign outputs[1775] = ~((layer0_outputs[7488]) ^ (layer0_outputs[5994]));
    assign outputs[1776] = (layer0_outputs[7615]) ^ (layer0_outputs[2369]);
    assign outputs[1777] = layer0_outputs[6458];
    assign outputs[1778] = (layer0_outputs[5448]) ^ (layer0_outputs[7536]);
    assign outputs[1779] = (layer0_outputs[6059]) | (layer0_outputs[6958]);
    assign outputs[1780] = (layer0_outputs[4495]) | (layer0_outputs[6050]);
    assign outputs[1781] = ~((layer0_outputs[376]) & (layer0_outputs[4519]));
    assign outputs[1782] = (layer0_outputs[3175]) & ~(layer0_outputs[1871]);
    assign outputs[1783] = ~(layer0_outputs[534]) | (layer0_outputs[2800]);
    assign outputs[1784] = layer0_outputs[6850];
    assign outputs[1785] = (layer0_outputs[624]) & (layer0_outputs[1563]);
    assign outputs[1786] = (layer0_outputs[864]) ^ (layer0_outputs[1439]);
    assign outputs[1787] = layer0_outputs[6372];
    assign outputs[1788] = layer0_outputs[4722];
    assign outputs[1789] = (layer0_outputs[2543]) ^ (layer0_outputs[7310]);
    assign outputs[1790] = (layer0_outputs[3757]) ^ (layer0_outputs[7494]);
    assign outputs[1791] = ~(layer0_outputs[3920]);
    assign outputs[1792] = layer0_outputs[7504];
    assign outputs[1793] = layer0_outputs[6198];
    assign outputs[1794] = layer0_outputs[5575];
    assign outputs[1795] = ~(layer0_outputs[7135]);
    assign outputs[1796] = (layer0_outputs[27]) | (layer0_outputs[810]);
    assign outputs[1797] = ~(layer0_outputs[683]);
    assign outputs[1798] = ~((layer0_outputs[7550]) ^ (layer0_outputs[3578]));
    assign outputs[1799] = ~(layer0_outputs[5664]);
    assign outputs[1800] = ~(layer0_outputs[4231]);
    assign outputs[1801] = ~((layer0_outputs[6091]) ^ (layer0_outputs[6986]));
    assign outputs[1802] = ~(layer0_outputs[1179]);
    assign outputs[1803] = ~(layer0_outputs[7212]);
    assign outputs[1804] = ~((layer0_outputs[424]) & (layer0_outputs[1665]));
    assign outputs[1805] = (layer0_outputs[6212]) | (layer0_outputs[4689]);
    assign outputs[1806] = ~((layer0_outputs[5232]) ^ (layer0_outputs[437]));
    assign outputs[1807] = layer0_outputs[2356];
    assign outputs[1808] = (layer0_outputs[438]) ^ (layer0_outputs[2200]);
    assign outputs[1809] = ~(layer0_outputs[1493]) | (layer0_outputs[6181]);
    assign outputs[1810] = layer0_outputs[5123];
    assign outputs[1811] = ~(layer0_outputs[6326]) | (layer0_outputs[4983]);
    assign outputs[1812] = ~(layer0_outputs[6631]);
    assign outputs[1813] = ~(layer0_outputs[161]);
    assign outputs[1814] = (layer0_outputs[6817]) ^ (layer0_outputs[2205]);
    assign outputs[1815] = ~((layer0_outputs[4627]) ^ (layer0_outputs[4829]));
    assign outputs[1816] = layer0_outputs[3841];
    assign outputs[1817] = (layer0_outputs[2020]) | (layer0_outputs[1630]);
    assign outputs[1818] = layer0_outputs[4827];
    assign outputs[1819] = layer0_outputs[2352];
    assign outputs[1820] = ~(layer0_outputs[3459]);
    assign outputs[1821] = ~(layer0_outputs[6110]);
    assign outputs[1822] = layer0_outputs[6692];
    assign outputs[1823] = ~(layer0_outputs[3212]) | (layer0_outputs[4749]);
    assign outputs[1824] = ~((layer0_outputs[715]) ^ (layer0_outputs[3390]));
    assign outputs[1825] = ~(layer0_outputs[1428]);
    assign outputs[1826] = layer0_outputs[6329];
    assign outputs[1827] = ~((layer0_outputs[635]) | (layer0_outputs[6709]));
    assign outputs[1828] = layer0_outputs[7583];
    assign outputs[1829] = ~((layer0_outputs[1273]) ^ (layer0_outputs[5100]));
    assign outputs[1830] = (layer0_outputs[1661]) | (layer0_outputs[4775]);
    assign outputs[1831] = ~((layer0_outputs[1223]) ^ (layer0_outputs[486]));
    assign outputs[1832] = (layer0_outputs[6346]) & ~(layer0_outputs[1684]);
    assign outputs[1833] = (layer0_outputs[962]) & ~(layer0_outputs[5698]);
    assign outputs[1834] = (layer0_outputs[3243]) ^ (layer0_outputs[5270]);
    assign outputs[1835] = (layer0_outputs[3728]) ^ (layer0_outputs[6187]);
    assign outputs[1836] = ~(layer0_outputs[3972]);
    assign outputs[1837] = ~((layer0_outputs[7434]) ^ (layer0_outputs[688]));
    assign outputs[1838] = ~((layer0_outputs[2282]) ^ (layer0_outputs[5689]));
    assign outputs[1839] = ~(layer0_outputs[5520]);
    assign outputs[1840] = (layer0_outputs[6965]) ^ (layer0_outputs[5954]);
    assign outputs[1841] = (layer0_outputs[2762]) ^ (layer0_outputs[6224]);
    assign outputs[1842] = ~(layer0_outputs[4049]);
    assign outputs[1843] = ~((layer0_outputs[5551]) ^ (layer0_outputs[7352]));
    assign outputs[1844] = layer0_outputs[4604];
    assign outputs[1845] = ~(layer0_outputs[3888]);
    assign outputs[1846] = (layer0_outputs[1345]) & ~(layer0_outputs[3375]);
    assign outputs[1847] = (layer0_outputs[4755]) ^ (layer0_outputs[1179]);
    assign outputs[1848] = ~(layer0_outputs[6840]);
    assign outputs[1849] = layer0_outputs[1596];
    assign outputs[1850] = (layer0_outputs[2932]) ^ (layer0_outputs[2219]);
    assign outputs[1851] = ~(layer0_outputs[2697]);
    assign outputs[1852] = layer0_outputs[2202];
    assign outputs[1853] = (layer0_outputs[3858]) & ~(layer0_outputs[2934]);
    assign outputs[1854] = ~(layer0_outputs[2504]);
    assign outputs[1855] = ~((layer0_outputs[3398]) ^ (layer0_outputs[6295]));
    assign outputs[1856] = ~(layer0_outputs[6052]) | (layer0_outputs[2464]);
    assign outputs[1857] = ~((layer0_outputs[2725]) ^ (layer0_outputs[3390]));
    assign outputs[1858] = layer0_outputs[7581];
    assign outputs[1859] = (layer0_outputs[7291]) ^ (layer0_outputs[1106]);
    assign outputs[1860] = (layer0_outputs[3110]) ^ (layer0_outputs[3259]);
    assign outputs[1861] = (layer0_outputs[6383]) & ~(layer0_outputs[5208]);
    assign outputs[1862] = (layer0_outputs[5320]) ^ (layer0_outputs[3177]);
    assign outputs[1863] = (layer0_outputs[7209]) ^ (layer0_outputs[6882]);
    assign outputs[1864] = ~(layer0_outputs[1249]) | (layer0_outputs[2685]);
    assign outputs[1865] = ~(layer0_outputs[304]);
    assign outputs[1866] = layer0_outputs[2106];
    assign outputs[1867] = (layer0_outputs[2348]) & (layer0_outputs[328]);
    assign outputs[1868] = (layer0_outputs[6822]) ^ (layer0_outputs[1081]);
    assign outputs[1869] = ~(layer0_outputs[1162]);
    assign outputs[1870] = ~(layer0_outputs[4065]) | (layer0_outputs[7559]);
    assign outputs[1871] = (layer0_outputs[5317]) ^ (layer0_outputs[1011]);
    assign outputs[1872] = (layer0_outputs[5542]) ^ (layer0_outputs[5785]);
    assign outputs[1873] = ~(layer0_outputs[4466]);
    assign outputs[1874] = layer0_outputs[269];
    assign outputs[1875] = layer0_outputs[7134];
    assign outputs[1876] = (layer0_outputs[3062]) & ~(layer0_outputs[5430]);
    assign outputs[1877] = layer0_outputs[4070];
    assign outputs[1878] = (layer0_outputs[2720]) ^ (layer0_outputs[4561]);
    assign outputs[1879] = ~(layer0_outputs[2732]) | (layer0_outputs[85]);
    assign outputs[1880] = (layer0_outputs[5284]) ^ (layer0_outputs[383]);
    assign outputs[1881] = ~(layer0_outputs[7652]);
    assign outputs[1882] = ~(layer0_outputs[6545]);
    assign outputs[1883] = (layer0_outputs[3148]) & ~(layer0_outputs[1210]);
    assign outputs[1884] = layer0_outputs[3260];
    assign outputs[1885] = layer0_outputs[2233];
    assign outputs[1886] = (layer0_outputs[6065]) & (layer0_outputs[2391]);
    assign outputs[1887] = layer0_outputs[3628];
    assign outputs[1888] = layer0_outputs[7090];
    assign outputs[1889] = ~(layer0_outputs[3698]);
    assign outputs[1890] = layer0_outputs[3810];
    assign outputs[1891] = (layer0_outputs[1004]) ^ (layer0_outputs[6191]);
    assign outputs[1892] = ~(layer0_outputs[3534]);
    assign outputs[1893] = ~(layer0_outputs[3733]);
    assign outputs[1894] = ~(layer0_outputs[4892]) | (layer0_outputs[1518]);
    assign outputs[1895] = ~(layer0_outputs[3323]);
    assign outputs[1896] = ~(layer0_outputs[3160]);
    assign outputs[1897] = ~((layer0_outputs[7655]) | (layer0_outputs[6746]));
    assign outputs[1898] = (layer0_outputs[4188]) & ~(layer0_outputs[4282]);
    assign outputs[1899] = ~((layer0_outputs[2033]) ^ (layer0_outputs[5989]));
    assign outputs[1900] = ~((layer0_outputs[1186]) ^ (layer0_outputs[1609]));
    assign outputs[1901] = ~(layer0_outputs[1191]) | (layer0_outputs[1398]);
    assign outputs[1902] = (layer0_outputs[7175]) & (layer0_outputs[1971]);
    assign outputs[1903] = layer0_outputs[5756];
    assign outputs[1904] = ~((layer0_outputs[7248]) & (layer0_outputs[5908]));
    assign outputs[1905] = ~(layer0_outputs[5405]);
    assign outputs[1906] = (layer0_outputs[5059]) ^ (layer0_outputs[5738]);
    assign outputs[1907] = ~(layer0_outputs[25]);
    assign outputs[1908] = ~(layer0_outputs[54]);
    assign outputs[1909] = layer0_outputs[2734];
    assign outputs[1910] = ~(layer0_outputs[6721]);
    assign outputs[1911] = ~(layer0_outputs[716]);
    assign outputs[1912] = ~((layer0_outputs[4160]) | (layer0_outputs[7080]));
    assign outputs[1913] = layer0_outputs[5063];
    assign outputs[1914] = (layer0_outputs[3673]) & ~(layer0_outputs[6703]);
    assign outputs[1915] = ~(layer0_outputs[1689]);
    assign outputs[1916] = (layer0_outputs[5681]) ^ (layer0_outputs[6043]);
    assign outputs[1917] = ~((layer0_outputs[2307]) ^ (layer0_outputs[266]));
    assign outputs[1918] = ~((layer0_outputs[587]) ^ (layer0_outputs[1204]));
    assign outputs[1919] = ~(layer0_outputs[3838]);
    assign outputs[1920] = ~((layer0_outputs[3538]) ^ (layer0_outputs[2701]));
    assign outputs[1921] = (layer0_outputs[2301]) & ~(layer0_outputs[143]);
    assign outputs[1922] = layer0_outputs[2830];
    assign outputs[1923] = (layer0_outputs[2923]) ^ (layer0_outputs[838]);
    assign outputs[1924] = (layer0_outputs[4981]) | (layer0_outputs[5771]);
    assign outputs[1925] = ~((layer0_outputs[1393]) ^ (layer0_outputs[6036]));
    assign outputs[1926] = ~(layer0_outputs[7667]) | (layer0_outputs[5010]);
    assign outputs[1927] = ~(layer0_outputs[7632]) | (layer0_outputs[527]);
    assign outputs[1928] = layer0_outputs[6607];
    assign outputs[1929] = (layer0_outputs[4159]) ^ (layer0_outputs[2855]);
    assign outputs[1930] = ~((layer0_outputs[3853]) ^ (layer0_outputs[2326]));
    assign outputs[1931] = (layer0_outputs[3526]) ^ (layer0_outputs[606]);
    assign outputs[1932] = (layer0_outputs[495]) | (layer0_outputs[3532]);
    assign outputs[1933] = ~(layer0_outputs[170]);
    assign outputs[1934] = ~(layer0_outputs[5390]);
    assign outputs[1935] = (layer0_outputs[4550]) ^ (layer0_outputs[5271]);
    assign outputs[1936] = ~(layer0_outputs[3799]) | (layer0_outputs[7544]);
    assign outputs[1937] = ~(layer0_outputs[2159]);
    assign outputs[1938] = ~(layer0_outputs[1599]);
    assign outputs[1939] = (layer0_outputs[4244]) ^ (layer0_outputs[3575]);
    assign outputs[1940] = ~(layer0_outputs[6121]);
    assign outputs[1941] = ~(layer0_outputs[1344]);
    assign outputs[1942] = (layer0_outputs[3722]) | (layer0_outputs[2456]);
    assign outputs[1943] = ~(layer0_outputs[2343]);
    assign outputs[1944] = layer0_outputs[1039];
    assign outputs[1945] = layer0_outputs[3505];
    assign outputs[1946] = ~(layer0_outputs[4241]);
    assign outputs[1947] = (layer0_outputs[3036]) & ~(layer0_outputs[3160]);
    assign outputs[1948] = ~(layer0_outputs[4066]);
    assign outputs[1949] = layer0_outputs[1439];
    assign outputs[1950] = ~(layer0_outputs[2451]);
    assign outputs[1951] = layer0_outputs[4603];
    assign outputs[1952] = ~((layer0_outputs[4994]) ^ (layer0_outputs[4210]));
    assign outputs[1953] = ~((layer0_outputs[1054]) ^ (layer0_outputs[6622]));
    assign outputs[1954] = layer0_outputs[270];
    assign outputs[1955] = (layer0_outputs[788]) & ~(layer0_outputs[1327]);
    assign outputs[1956] = 1'b1;
    assign outputs[1957] = layer0_outputs[6989];
    assign outputs[1958] = ~((layer0_outputs[4825]) ^ (layer0_outputs[1080]));
    assign outputs[1959] = layer0_outputs[3539];
    assign outputs[1960] = ~(layer0_outputs[2028]);
    assign outputs[1961] = ~(layer0_outputs[3330]);
    assign outputs[1962] = layer0_outputs[1124];
    assign outputs[1963] = ~((layer0_outputs[7288]) | (layer0_outputs[1794]));
    assign outputs[1964] = ~(layer0_outputs[5111]);
    assign outputs[1965] = (layer0_outputs[3310]) | (layer0_outputs[3824]);
    assign outputs[1966] = layer0_outputs[3554];
    assign outputs[1967] = (layer0_outputs[2507]) ^ (layer0_outputs[5887]);
    assign outputs[1968] = layer0_outputs[5541];
    assign outputs[1969] = ~(layer0_outputs[6190]);
    assign outputs[1970] = ~(layer0_outputs[3459]);
    assign outputs[1971] = layer0_outputs[5439];
    assign outputs[1972] = (layer0_outputs[2811]) | (layer0_outputs[5936]);
    assign outputs[1973] = (layer0_outputs[7585]) ^ (layer0_outputs[2665]);
    assign outputs[1974] = layer0_outputs[1897];
    assign outputs[1975] = ~((layer0_outputs[709]) ^ (layer0_outputs[3585]));
    assign outputs[1976] = ~(layer0_outputs[1136]);
    assign outputs[1977] = ~(layer0_outputs[1233]) | (layer0_outputs[114]);
    assign outputs[1978] = ~(layer0_outputs[3151]) | (layer0_outputs[5462]);
    assign outputs[1979] = ~(layer0_outputs[2917]);
    assign outputs[1980] = ~(layer0_outputs[4543]);
    assign outputs[1981] = (layer0_outputs[4691]) ^ (layer0_outputs[309]);
    assign outputs[1982] = layer0_outputs[5977];
    assign outputs[1983] = (layer0_outputs[1482]) & ~(layer0_outputs[5129]);
    assign outputs[1984] = ~(layer0_outputs[3869]);
    assign outputs[1985] = (layer0_outputs[2514]) & ~(layer0_outputs[3910]);
    assign outputs[1986] = ~(layer0_outputs[3343]);
    assign outputs[1987] = layer0_outputs[4044];
    assign outputs[1988] = (layer0_outputs[5476]) & (layer0_outputs[3762]);
    assign outputs[1989] = ~(layer0_outputs[7366]);
    assign outputs[1990] = ~((layer0_outputs[2555]) ^ (layer0_outputs[5540]));
    assign outputs[1991] = ~((layer0_outputs[4263]) | (layer0_outputs[2772]));
    assign outputs[1992] = (layer0_outputs[3247]) ^ (layer0_outputs[7100]);
    assign outputs[1993] = ~(layer0_outputs[7017]);
    assign outputs[1994] = layer0_outputs[6142];
    assign outputs[1995] = layer0_outputs[1525];
    assign outputs[1996] = (layer0_outputs[1261]) | (layer0_outputs[161]);
    assign outputs[1997] = layer0_outputs[5008];
    assign outputs[1998] = ~((layer0_outputs[710]) ^ (layer0_outputs[7469]));
    assign outputs[1999] = ~(layer0_outputs[5627]);
    assign outputs[2000] = ~((layer0_outputs[3718]) ^ (layer0_outputs[6724]));
    assign outputs[2001] = layer0_outputs[6129];
    assign outputs[2002] = ~(layer0_outputs[1773]);
    assign outputs[2003] = (layer0_outputs[597]) ^ (layer0_outputs[151]);
    assign outputs[2004] = layer0_outputs[713];
    assign outputs[2005] = ~(layer0_outputs[1801]);
    assign outputs[2006] = ~(layer0_outputs[5224]);
    assign outputs[2007] = ~((layer0_outputs[806]) ^ (layer0_outputs[1045]));
    assign outputs[2008] = ~(layer0_outputs[3759]);
    assign outputs[2009] = ~((layer0_outputs[3304]) | (layer0_outputs[4664]));
    assign outputs[2010] = layer0_outputs[3038];
    assign outputs[2011] = layer0_outputs[540];
    assign outputs[2012] = (layer0_outputs[3380]) ^ (layer0_outputs[3033]);
    assign outputs[2013] = (layer0_outputs[4671]) & ~(layer0_outputs[7307]);
    assign outputs[2014] = layer0_outputs[3886];
    assign outputs[2015] = ~(layer0_outputs[2334]) | (layer0_outputs[6035]);
    assign outputs[2016] = (layer0_outputs[6873]) & (layer0_outputs[7265]);
    assign outputs[2017] = layer0_outputs[1283];
    assign outputs[2018] = (layer0_outputs[2722]) ^ (layer0_outputs[6361]);
    assign outputs[2019] = ~((layer0_outputs[2178]) & (layer0_outputs[7196]));
    assign outputs[2020] = ~(layer0_outputs[7237]);
    assign outputs[2021] = ~((layer0_outputs[682]) & (layer0_outputs[1634]));
    assign outputs[2022] = ~(layer0_outputs[3466]) | (layer0_outputs[6976]);
    assign outputs[2023] = ~(layer0_outputs[7423]);
    assign outputs[2024] = layer0_outputs[5936];
    assign outputs[2025] = ~((layer0_outputs[1767]) ^ (layer0_outputs[5594]));
    assign outputs[2026] = ~(layer0_outputs[5871]);
    assign outputs[2027] = ~(layer0_outputs[246]) | (layer0_outputs[5909]);
    assign outputs[2028] = layer0_outputs[2966];
    assign outputs[2029] = (layer0_outputs[6167]) ^ (layer0_outputs[4853]);
    assign outputs[2030] = ~((layer0_outputs[7393]) ^ (layer0_outputs[1717]));
    assign outputs[2031] = (layer0_outputs[4828]) | (layer0_outputs[2290]);
    assign outputs[2032] = ~(layer0_outputs[6938]);
    assign outputs[2033] = ~(layer0_outputs[1190]);
    assign outputs[2034] = ~(layer0_outputs[3833]) | (layer0_outputs[6530]);
    assign outputs[2035] = (layer0_outputs[524]) ^ (layer0_outputs[4943]);
    assign outputs[2036] = (layer0_outputs[6054]) & ~(layer0_outputs[6685]);
    assign outputs[2037] = ~(layer0_outputs[7112]);
    assign outputs[2038] = ~((layer0_outputs[1324]) ^ (layer0_outputs[2941]));
    assign outputs[2039] = ~((layer0_outputs[1041]) ^ (layer0_outputs[1636]));
    assign outputs[2040] = layer0_outputs[7466];
    assign outputs[2041] = ~(layer0_outputs[7064]) | (layer0_outputs[3517]);
    assign outputs[2042] = ~((layer0_outputs[7497]) ^ (layer0_outputs[1523]));
    assign outputs[2043] = ~((layer0_outputs[3267]) ^ (layer0_outputs[5845]));
    assign outputs[2044] = ~(layer0_outputs[4159]) | (layer0_outputs[554]);
    assign outputs[2045] = (layer0_outputs[1901]) | (layer0_outputs[88]);
    assign outputs[2046] = layer0_outputs[7136];
    assign outputs[2047] = ~(layer0_outputs[7658]);
    assign outputs[2048] = ~((layer0_outputs[5256]) | (layer0_outputs[5186]));
    assign outputs[2049] = (layer0_outputs[3990]) | (layer0_outputs[7560]);
    assign outputs[2050] = layer0_outputs[7316];
    assign outputs[2051] = (layer0_outputs[2110]) ^ (layer0_outputs[1254]);
    assign outputs[2052] = layer0_outputs[7284];
    assign outputs[2053] = ~(layer0_outputs[1241]);
    assign outputs[2054] = ~((layer0_outputs[2612]) & (layer0_outputs[2070]));
    assign outputs[2055] = layer0_outputs[695];
    assign outputs[2056] = ~(layer0_outputs[3116]);
    assign outputs[2057] = ~((layer0_outputs[5769]) & (layer0_outputs[5612]));
    assign outputs[2058] = ~((layer0_outputs[4225]) ^ (layer0_outputs[3024]));
    assign outputs[2059] = ~(layer0_outputs[1205]);
    assign outputs[2060] = ~((layer0_outputs[7638]) ^ (layer0_outputs[2499]));
    assign outputs[2061] = ~(layer0_outputs[3224]) | (layer0_outputs[2684]);
    assign outputs[2062] = ~(layer0_outputs[6533]);
    assign outputs[2063] = layer0_outputs[1280];
    assign outputs[2064] = ~(layer0_outputs[1828]);
    assign outputs[2065] = ~((layer0_outputs[7165]) ^ (layer0_outputs[361]));
    assign outputs[2066] = ~(layer0_outputs[3736]) | (layer0_outputs[588]);
    assign outputs[2067] = (layer0_outputs[6762]) & ~(layer0_outputs[5301]);
    assign outputs[2068] = (layer0_outputs[3593]) ^ (layer0_outputs[46]);
    assign outputs[2069] = ~((layer0_outputs[199]) ^ (layer0_outputs[7078]));
    assign outputs[2070] = ~(layer0_outputs[3406]);
    assign outputs[2071] = ~((layer0_outputs[1401]) & (layer0_outputs[6027]));
    assign outputs[2072] = layer0_outputs[7465];
    assign outputs[2073] = ~(layer0_outputs[4263]);
    assign outputs[2074] = 1'b1;
    assign outputs[2075] = ~(layer0_outputs[3809]);
    assign outputs[2076] = ~((layer0_outputs[102]) ^ (layer0_outputs[2284]));
    assign outputs[2077] = (layer0_outputs[6255]) ^ (layer0_outputs[4135]);
    assign outputs[2078] = ~((layer0_outputs[3437]) & (layer0_outputs[3270]));
    assign outputs[2079] = ~((layer0_outputs[887]) | (layer0_outputs[6416]));
    assign outputs[2080] = layer0_outputs[6071];
    assign outputs[2081] = ~(layer0_outputs[3446]) | (layer0_outputs[5865]);
    assign outputs[2082] = ~(layer0_outputs[6613]);
    assign outputs[2083] = ~(layer0_outputs[2398]);
    assign outputs[2084] = layer0_outputs[6172];
    assign outputs[2085] = (layer0_outputs[3581]) & ~(layer0_outputs[1282]);
    assign outputs[2086] = ~(layer0_outputs[5355]);
    assign outputs[2087] = layer0_outputs[4794];
    assign outputs[2088] = (layer0_outputs[3620]) & ~(layer0_outputs[7586]);
    assign outputs[2089] = ~(layer0_outputs[4558]);
    assign outputs[2090] = ~((layer0_outputs[2273]) ^ (layer0_outputs[6559]));
    assign outputs[2091] = layer0_outputs[2300];
    assign outputs[2092] = ~(layer0_outputs[7536]);
    assign outputs[2093] = ~(layer0_outputs[5504]) | (layer0_outputs[6242]);
    assign outputs[2094] = ~((layer0_outputs[2577]) ^ (layer0_outputs[1020]));
    assign outputs[2095] = layer0_outputs[7273];
    assign outputs[2096] = layer0_outputs[7391];
    assign outputs[2097] = layer0_outputs[2411];
    assign outputs[2098] = layer0_outputs[3009];
    assign outputs[2099] = ~((layer0_outputs[5955]) | (layer0_outputs[2832]));
    assign outputs[2100] = layer0_outputs[425];
    assign outputs[2101] = ~(layer0_outputs[5584]);
    assign outputs[2102] = ~(layer0_outputs[2288]) | (layer0_outputs[3663]);
    assign outputs[2103] = layer0_outputs[4405];
    assign outputs[2104] = ~(layer0_outputs[512]);
    assign outputs[2105] = ~(layer0_outputs[2138]);
    assign outputs[2106] = layer0_outputs[4011];
    assign outputs[2107] = ~(layer0_outputs[4502]);
    assign outputs[2108] = (layer0_outputs[5986]) ^ (layer0_outputs[6357]);
    assign outputs[2109] = layer0_outputs[1454];
    assign outputs[2110] = layer0_outputs[2683];
    assign outputs[2111] = (layer0_outputs[7675]) ^ (layer0_outputs[983]);
    assign outputs[2112] = ~(layer0_outputs[2845]) | (layer0_outputs[3040]);
    assign outputs[2113] = (layer0_outputs[6189]) ^ (layer0_outputs[5689]);
    assign outputs[2114] = ~((layer0_outputs[6381]) | (layer0_outputs[1468]));
    assign outputs[2115] = (layer0_outputs[6432]) | (layer0_outputs[1077]);
    assign outputs[2116] = ~(layer0_outputs[1838]) | (layer0_outputs[865]);
    assign outputs[2117] = ~(layer0_outputs[6020]) | (layer0_outputs[414]);
    assign outputs[2118] = ~(layer0_outputs[6591]) | (layer0_outputs[6112]);
    assign outputs[2119] = ~(layer0_outputs[7385]);
    assign outputs[2120] = ~(layer0_outputs[4872]);
    assign outputs[2121] = (layer0_outputs[6731]) ^ (layer0_outputs[4649]);
    assign outputs[2122] = ~(layer0_outputs[3641]);
    assign outputs[2123] = ~(layer0_outputs[526]) | (layer0_outputs[6485]);
    assign outputs[2124] = layer0_outputs[5296];
    assign outputs[2125] = (layer0_outputs[2900]) ^ (layer0_outputs[5427]);
    assign outputs[2126] = layer0_outputs[5370];
    assign outputs[2127] = layer0_outputs[2672];
    assign outputs[2128] = layer0_outputs[6546];
    assign outputs[2129] = ~(layer0_outputs[3699]);
    assign outputs[2130] = ~((layer0_outputs[1919]) ^ (layer0_outputs[1954]));
    assign outputs[2131] = layer0_outputs[956];
    assign outputs[2132] = ~(layer0_outputs[6972]);
    assign outputs[2133] = ~(layer0_outputs[4148]);
    assign outputs[2134] = ~(layer0_outputs[5505]) | (layer0_outputs[244]);
    assign outputs[2135] = (layer0_outputs[6]) & ~(layer0_outputs[2091]);
    assign outputs[2136] = (layer0_outputs[5667]) | (layer0_outputs[3984]);
    assign outputs[2137] = ~(layer0_outputs[3361]);
    assign outputs[2138] = ~(layer0_outputs[4926]) | (layer0_outputs[5087]);
    assign outputs[2139] = layer0_outputs[3683];
    assign outputs[2140] = ~(layer0_outputs[6435]);
    assign outputs[2141] = layer0_outputs[3500];
    assign outputs[2142] = ~(layer0_outputs[354]) | (layer0_outputs[4577]);
    assign outputs[2143] = ~(layer0_outputs[5862]);
    assign outputs[2144] = ~((layer0_outputs[562]) ^ (layer0_outputs[771]));
    assign outputs[2145] = ~((layer0_outputs[3305]) & (layer0_outputs[1589]));
    assign outputs[2146] = ~(layer0_outputs[2385]);
    assign outputs[2147] = (layer0_outputs[7217]) ^ (layer0_outputs[1412]);
    assign outputs[2148] = 1'b1;
    assign outputs[2149] = (layer0_outputs[4213]) ^ (layer0_outputs[3331]);
    assign outputs[2150] = (layer0_outputs[1132]) & ~(layer0_outputs[7606]);
    assign outputs[2151] = ~(layer0_outputs[7410]);
    assign outputs[2152] = layer0_outputs[6676];
    assign outputs[2153] = (layer0_outputs[4431]) ^ (layer0_outputs[511]);
    assign outputs[2154] = ~(layer0_outputs[5471]);
    assign outputs[2155] = ~(layer0_outputs[2564]) | (layer0_outputs[3234]);
    assign outputs[2156] = ~((layer0_outputs[5376]) & (layer0_outputs[4403]));
    assign outputs[2157] = ~(layer0_outputs[3662]);
    assign outputs[2158] = (layer0_outputs[6888]) ^ (layer0_outputs[4947]);
    assign outputs[2159] = (layer0_outputs[1749]) & ~(layer0_outputs[3229]);
    assign outputs[2160] = ~((layer0_outputs[4241]) ^ (layer0_outputs[3501]));
    assign outputs[2161] = ~(layer0_outputs[7314]);
    assign outputs[2162] = (layer0_outputs[5588]) ^ (layer0_outputs[2200]);
    assign outputs[2163] = layer0_outputs[4059];
    assign outputs[2164] = layer0_outputs[5038];
    assign outputs[2165] = layer0_outputs[4003];
    assign outputs[2166] = ~(layer0_outputs[3607]) | (layer0_outputs[51]);
    assign outputs[2167] = ~((layer0_outputs[7380]) ^ (layer0_outputs[5292]));
    assign outputs[2168] = (layer0_outputs[2508]) & ~(layer0_outputs[3355]);
    assign outputs[2169] = ~(layer0_outputs[7396]) | (layer0_outputs[5956]);
    assign outputs[2170] = (layer0_outputs[663]) ^ (layer0_outputs[4836]);
    assign outputs[2171] = layer0_outputs[3074];
    assign outputs[2172] = (layer0_outputs[4564]) ^ (layer0_outputs[3496]);
    assign outputs[2173] = ~(layer0_outputs[5711]);
    assign outputs[2174] = (layer0_outputs[288]) & ~(layer0_outputs[2312]);
    assign outputs[2175] = ~((layer0_outputs[6902]) ^ (layer0_outputs[5528]));
    assign outputs[2176] = ~((layer0_outputs[3295]) & (layer0_outputs[2057]));
    assign outputs[2177] = ~(layer0_outputs[1076]) | (layer0_outputs[1950]);
    assign outputs[2178] = ~((layer0_outputs[7097]) & (layer0_outputs[4444]));
    assign outputs[2179] = ~(layer0_outputs[7558]);
    assign outputs[2180] = ~(layer0_outputs[3526]) | (layer0_outputs[7113]);
    assign outputs[2181] = ~(layer0_outputs[7230]);
    assign outputs[2182] = layer0_outputs[2719];
    assign outputs[2183] = layer0_outputs[6216];
    assign outputs[2184] = ~((layer0_outputs[6343]) | (layer0_outputs[2900]));
    assign outputs[2185] = ~((layer0_outputs[3107]) ^ (layer0_outputs[7363]));
    assign outputs[2186] = (layer0_outputs[679]) ^ (layer0_outputs[2310]);
    assign outputs[2187] = ~((layer0_outputs[2233]) ^ (layer0_outputs[2192]));
    assign outputs[2188] = ~(layer0_outputs[5395]);
    assign outputs[2189] = ~((layer0_outputs[4552]) ^ (layer0_outputs[1407]));
    assign outputs[2190] = ~(layer0_outputs[7480]);
    assign outputs[2191] = ~(layer0_outputs[1695]);
    assign outputs[2192] = layer0_outputs[2339];
    assign outputs[2193] = (layer0_outputs[5953]) & ~(layer0_outputs[446]);
    assign outputs[2194] = layer0_outputs[1988];
    assign outputs[2195] = ~(layer0_outputs[4873]) | (layer0_outputs[4459]);
    assign outputs[2196] = layer0_outputs[3418];
    assign outputs[2197] = ~(layer0_outputs[7574]) | (layer0_outputs[4220]);
    assign outputs[2198] = (layer0_outputs[3193]) ^ (layer0_outputs[5279]);
    assign outputs[2199] = ~(layer0_outputs[5326]);
    assign outputs[2200] = ~(layer0_outputs[6923]) | (layer0_outputs[7240]);
    assign outputs[2201] = ~(layer0_outputs[6591]) | (layer0_outputs[4844]);
    assign outputs[2202] = (layer0_outputs[5854]) & (layer0_outputs[2113]);
    assign outputs[2203] = ~((layer0_outputs[5539]) ^ (layer0_outputs[3169]));
    assign outputs[2204] = layer0_outputs[3297];
    assign outputs[2205] = ~(layer0_outputs[741]) | (layer0_outputs[5848]);
    assign outputs[2206] = (layer0_outputs[3388]) ^ (layer0_outputs[48]);
    assign outputs[2207] = layer0_outputs[4413];
    assign outputs[2208] = ~(layer0_outputs[1173]);
    assign outputs[2209] = ~((layer0_outputs[2994]) & (layer0_outputs[5480]));
    assign outputs[2210] = (layer0_outputs[250]) ^ (layer0_outputs[2451]);
    assign outputs[2211] = ~(layer0_outputs[2565]);
    assign outputs[2212] = ~((layer0_outputs[1159]) ^ (layer0_outputs[3325]));
    assign outputs[2213] = layer0_outputs[52];
    assign outputs[2214] = ~(layer0_outputs[1126]);
    assign outputs[2215] = ~(layer0_outputs[81]);
    assign outputs[2216] = layer0_outputs[5400];
    assign outputs[2217] = layer0_outputs[2158];
    assign outputs[2218] = ~((layer0_outputs[569]) | (layer0_outputs[866]));
    assign outputs[2219] = (layer0_outputs[2600]) & ~(layer0_outputs[1976]);
    assign outputs[2220] = (layer0_outputs[993]) ^ (layer0_outputs[7358]);
    assign outputs[2221] = ~(layer0_outputs[2082]) | (layer0_outputs[703]);
    assign outputs[2222] = ~(layer0_outputs[5904]);
    assign outputs[2223] = (layer0_outputs[2155]) ^ (layer0_outputs[2443]);
    assign outputs[2224] = ~(layer0_outputs[7066]) | (layer0_outputs[4270]);
    assign outputs[2225] = layer0_outputs[2116];
    assign outputs[2226] = (layer0_outputs[4259]) & ~(layer0_outputs[4489]);
    assign outputs[2227] = layer0_outputs[397];
    assign outputs[2228] = (layer0_outputs[3944]) & ~(layer0_outputs[194]);
    assign outputs[2229] = (layer0_outputs[5400]) & ~(layer0_outputs[4544]);
    assign outputs[2230] = ~(layer0_outputs[4937]);
    assign outputs[2231] = ~(layer0_outputs[6456]) | (layer0_outputs[6086]);
    assign outputs[2232] = (layer0_outputs[1706]) ^ (layer0_outputs[5599]);
    assign outputs[2233] = (layer0_outputs[2811]) | (layer0_outputs[236]);
    assign outputs[2234] = ~(layer0_outputs[3684]);
    assign outputs[2235] = ~(layer0_outputs[1103]);
    assign outputs[2236] = layer0_outputs[7583];
    assign outputs[2237] = layer0_outputs[4633];
    assign outputs[2238] = ~(layer0_outputs[357]);
    assign outputs[2239] = ~((layer0_outputs[117]) | (layer0_outputs[6391]));
    assign outputs[2240] = (layer0_outputs[201]) & (layer0_outputs[3601]);
    assign outputs[2241] = ~((layer0_outputs[558]) ^ (layer0_outputs[110]));
    assign outputs[2242] = ~((layer0_outputs[5318]) & (layer0_outputs[253]));
    assign outputs[2243] = ~(layer0_outputs[6479]);
    assign outputs[2244] = ~(layer0_outputs[241]);
    assign outputs[2245] = (layer0_outputs[5177]) | (layer0_outputs[4087]);
    assign outputs[2246] = ~(layer0_outputs[2025]);
    assign outputs[2247] = ~((layer0_outputs[4280]) ^ (layer0_outputs[12]));
    assign outputs[2248] = (layer0_outputs[6187]) | (layer0_outputs[5892]);
    assign outputs[2249] = (layer0_outputs[4215]) ^ (layer0_outputs[2786]);
    assign outputs[2250] = layer0_outputs[6495];
    assign outputs[2251] = ~(layer0_outputs[3439]);
    assign outputs[2252] = layer0_outputs[752];
    assign outputs[2253] = ~(layer0_outputs[6895]) | (layer0_outputs[4834]);
    assign outputs[2254] = ~(layer0_outputs[1166]);
    assign outputs[2255] = ~(layer0_outputs[4091]) | (layer0_outputs[2079]);
    assign outputs[2256] = ~(layer0_outputs[1912]);
    assign outputs[2257] = ~((layer0_outputs[1942]) | (layer0_outputs[1731]));
    assign outputs[2258] = ~(layer0_outputs[2021]);
    assign outputs[2259] = (layer0_outputs[6477]) ^ (layer0_outputs[5408]);
    assign outputs[2260] = (layer0_outputs[6284]) | (layer0_outputs[4357]);
    assign outputs[2261] = ~(layer0_outputs[4949]);
    assign outputs[2262] = layer0_outputs[6067];
    assign outputs[2263] = (layer0_outputs[6646]) | (layer0_outputs[3739]);
    assign outputs[2264] = ~((layer0_outputs[502]) | (layer0_outputs[6069]));
    assign outputs[2265] = layer0_outputs[558];
    assign outputs[2266] = ~(layer0_outputs[5596]);
    assign outputs[2267] = (layer0_outputs[5918]) & ~(layer0_outputs[2864]);
    assign outputs[2268] = (layer0_outputs[2108]) & (layer0_outputs[3889]);
    assign outputs[2269] = (layer0_outputs[4146]) ^ (layer0_outputs[7449]);
    assign outputs[2270] = ~(layer0_outputs[3639]);
    assign outputs[2271] = (layer0_outputs[6773]) ^ (layer0_outputs[2930]);
    assign outputs[2272] = ~(layer0_outputs[4563]) | (layer0_outputs[706]);
    assign outputs[2273] = ~(layer0_outputs[4686]);
    assign outputs[2274] = ~((layer0_outputs[75]) | (layer0_outputs[5436]));
    assign outputs[2275] = ~(layer0_outputs[5459]) | (layer0_outputs[655]);
    assign outputs[2276] = ~(layer0_outputs[1195]);
    assign outputs[2277] = ~(layer0_outputs[5306]) | (layer0_outputs[653]);
    assign outputs[2278] = layer0_outputs[6225];
    assign outputs[2279] = ~((layer0_outputs[4907]) & (layer0_outputs[3859]));
    assign outputs[2280] = (layer0_outputs[7604]) ^ (layer0_outputs[3222]);
    assign outputs[2281] = (layer0_outputs[1065]) ^ (layer0_outputs[4183]);
    assign outputs[2282] = (layer0_outputs[813]) & ~(layer0_outputs[3288]);
    assign outputs[2283] = layer0_outputs[971];
    assign outputs[2284] = layer0_outputs[2953];
    assign outputs[2285] = layer0_outputs[1198];
    assign outputs[2286] = ~((layer0_outputs[1400]) ^ (layer0_outputs[7150]));
    assign outputs[2287] = ~((layer0_outputs[6781]) ^ (layer0_outputs[933]));
    assign outputs[2288] = layer0_outputs[7110];
    assign outputs[2289] = ~((layer0_outputs[6772]) ^ (layer0_outputs[5759]));
    assign outputs[2290] = ~(layer0_outputs[1710]);
    assign outputs[2291] = 1'b1;
    assign outputs[2292] = layer0_outputs[7058];
    assign outputs[2293] = layer0_outputs[3147];
    assign outputs[2294] = ~(layer0_outputs[4457]) | (layer0_outputs[4990]);
    assign outputs[2295] = ~((layer0_outputs[5521]) & (layer0_outputs[4704]));
    assign outputs[2296] = layer0_outputs[5495];
    assign outputs[2297] = (layer0_outputs[1523]) ^ (layer0_outputs[6727]);
    assign outputs[2298] = layer0_outputs[6233];
    assign outputs[2299] = ~((layer0_outputs[3595]) | (layer0_outputs[2751]));
    assign outputs[2300] = layer0_outputs[1718];
    assign outputs[2301] = ~(layer0_outputs[512]);
    assign outputs[2302] = layer0_outputs[3022];
    assign outputs[2303] = layer0_outputs[420];
    assign outputs[2304] = layer0_outputs[3801];
    assign outputs[2305] = ~(layer0_outputs[3503]);
    assign outputs[2306] = layer0_outputs[3991];
    assign outputs[2307] = ~(layer0_outputs[6395]) | (layer0_outputs[3307]);
    assign outputs[2308] = (layer0_outputs[375]) & ~(layer0_outputs[6034]);
    assign outputs[2309] = ~(layer0_outputs[6228]) | (layer0_outputs[5953]);
    assign outputs[2310] = ~((layer0_outputs[5835]) | (layer0_outputs[4383]));
    assign outputs[2311] = layer0_outputs[4852];
    assign outputs[2312] = (layer0_outputs[2610]) & ~(layer0_outputs[2587]);
    assign outputs[2313] = (layer0_outputs[7662]) & ~(layer0_outputs[5132]);
    assign outputs[2314] = ~(layer0_outputs[4133]) | (layer0_outputs[7054]);
    assign outputs[2315] = ~(layer0_outputs[3411]) | (layer0_outputs[10]);
    assign outputs[2316] = ~(layer0_outputs[1130]);
    assign outputs[2317] = (layer0_outputs[6109]) & ~(layer0_outputs[239]);
    assign outputs[2318] = ~(layer0_outputs[2907]) | (layer0_outputs[6435]);
    assign outputs[2319] = ~(layer0_outputs[3518]);
    assign outputs[2320] = layer0_outputs[7455];
    assign outputs[2321] = 1'b1;
    assign outputs[2322] = ~((layer0_outputs[5280]) & (layer0_outputs[6314]));
    assign outputs[2323] = ~(layer0_outputs[4681]) | (layer0_outputs[4045]);
    assign outputs[2324] = (layer0_outputs[999]) & ~(layer0_outputs[2687]);
    assign outputs[2325] = (layer0_outputs[2501]) & (layer0_outputs[1239]);
    assign outputs[2326] = layer0_outputs[2328];
    assign outputs[2327] = layer0_outputs[614];
    assign outputs[2328] = (layer0_outputs[4536]) ^ (layer0_outputs[5257]);
    assign outputs[2329] = ~(layer0_outputs[995]) | (layer0_outputs[6641]);
    assign outputs[2330] = layer0_outputs[1365];
    assign outputs[2331] = ~((layer0_outputs[2335]) ^ (layer0_outputs[753]));
    assign outputs[2332] = (layer0_outputs[2476]) | (layer0_outputs[6521]);
    assign outputs[2333] = ~(layer0_outputs[2136]);
    assign outputs[2334] = layer0_outputs[5776];
    assign outputs[2335] = ~(layer0_outputs[4620]) | (layer0_outputs[3648]);
    assign outputs[2336] = (layer0_outputs[7208]) ^ (layer0_outputs[1013]);
    assign outputs[2337] = ~(layer0_outputs[3521]);
    assign outputs[2338] = ~((layer0_outputs[6674]) & (layer0_outputs[4601]));
    assign outputs[2339] = (layer0_outputs[4862]) & ~(layer0_outputs[1097]);
    assign outputs[2340] = layer0_outputs[5498];
    assign outputs[2341] = ~(layer0_outputs[7091]);
    assign outputs[2342] = layer0_outputs[144];
    assign outputs[2343] = ~(layer0_outputs[3374]);
    assign outputs[2344] = (layer0_outputs[2002]) & (layer0_outputs[5975]);
    assign outputs[2345] = ~((layer0_outputs[2464]) ^ (layer0_outputs[4460]));
    assign outputs[2346] = ~((layer0_outputs[7526]) | (layer0_outputs[3458]));
    assign outputs[2347] = (layer0_outputs[3769]) ^ (layer0_outputs[508]);
    assign outputs[2348] = (layer0_outputs[384]) & ~(layer0_outputs[1829]);
    assign outputs[2349] = (layer0_outputs[3595]) ^ (layer0_outputs[5394]);
    assign outputs[2350] = ~(layer0_outputs[6396]);
    assign outputs[2351] = ~((layer0_outputs[3302]) | (layer0_outputs[2123]));
    assign outputs[2352] = ~(layer0_outputs[6370]);
    assign outputs[2353] = ~(layer0_outputs[2816]) | (layer0_outputs[4171]);
    assign outputs[2354] = layer0_outputs[5626];
    assign outputs[2355] = ~(layer0_outputs[4533]);
    assign outputs[2356] = (layer0_outputs[3604]) ^ (layer0_outputs[2890]);
    assign outputs[2357] = ~(layer0_outputs[7027]) | (layer0_outputs[7530]);
    assign outputs[2358] = ~((layer0_outputs[1637]) ^ (layer0_outputs[1383]));
    assign outputs[2359] = ~(layer0_outputs[6239]) | (layer0_outputs[3273]);
    assign outputs[2360] = (layer0_outputs[6386]) ^ (layer0_outputs[6087]);
    assign outputs[2361] = layer0_outputs[4392];
    assign outputs[2362] = layer0_outputs[4039];
    assign outputs[2363] = layer0_outputs[4737];
    assign outputs[2364] = layer0_outputs[97];
    assign outputs[2365] = layer0_outputs[4329];
    assign outputs[2366] = (layer0_outputs[1480]) & ~(layer0_outputs[4131]);
    assign outputs[2367] = ~((layer0_outputs[5093]) ^ (layer0_outputs[7200]));
    assign outputs[2368] = ~(layer0_outputs[1231]);
    assign outputs[2369] = ~(layer0_outputs[5162]);
    assign outputs[2370] = layer0_outputs[7373];
    assign outputs[2371] = ~(layer0_outputs[1717]) | (layer0_outputs[1854]);
    assign outputs[2372] = ~(layer0_outputs[3332]);
    assign outputs[2373] = (layer0_outputs[2812]) | (layer0_outputs[6986]);
    assign outputs[2374] = layer0_outputs[2465];
    assign outputs[2375] = ~(layer0_outputs[2254]);
    assign outputs[2376] = layer0_outputs[4979];
    assign outputs[2377] = (layer0_outputs[4023]) ^ (layer0_outputs[7007]);
    assign outputs[2378] = ~((layer0_outputs[2831]) & (layer0_outputs[3509]));
    assign outputs[2379] = layer0_outputs[4278];
    assign outputs[2380] = ~(layer0_outputs[2482]);
    assign outputs[2381] = ~(layer0_outputs[4501]);
    assign outputs[2382] = ~(layer0_outputs[2308]);
    assign outputs[2383] = (layer0_outputs[5495]) & ~(layer0_outputs[6088]);
    assign outputs[2384] = ~(layer0_outputs[6046]);
    assign outputs[2385] = layer0_outputs[6265];
    assign outputs[2386] = (layer0_outputs[2157]) & (layer0_outputs[6969]);
    assign outputs[2387] = (layer0_outputs[2927]) & ~(layer0_outputs[4660]);
    assign outputs[2388] = ~(layer0_outputs[7255]);
    assign outputs[2389] = layer0_outputs[5640];
    assign outputs[2390] = ~(layer0_outputs[7255]);
    assign outputs[2391] = ~((layer0_outputs[605]) ^ (layer0_outputs[2948]));
    assign outputs[2392] = (layer0_outputs[2401]) ^ (layer0_outputs[4588]);
    assign outputs[2393] = layer0_outputs[3306];
    assign outputs[2394] = ~((layer0_outputs[2476]) ^ (layer0_outputs[6277]));
    assign outputs[2395] = (layer0_outputs[1014]) | (layer0_outputs[2117]);
    assign outputs[2396] = ~(layer0_outputs[3367]);
    assign outputs[2397] = ~((layer0_outputs[7496]) ^ (layer0_outputs[4048]));
    assign outputs[2398] = layer0_outputs[5254];
    assign outputs[2399] = ~(layer0_outputs[453]);
    assign outputs[2400] = ~(layer0_outputs[208]);
    assign outputs[2401] = ~(layer0_outputs[1152]);
    assign outputs[2402] = (layer0_outputs[3716]) & (layer0_outputs[3754]);
    assign outputs[2403] = ~((layer0_outputs[4814]) ^ (layer0_outputs[2358]));
    assign outputs[2404] = ~((layer0_outputs[661]) ^ (layer0_outputs[3959]));
    assign outputs[2405] = (layer0_outputs[157]) | (layer0_outputs[4029]);
    assign outputs[2406] = ~(layer0_outputs[7642]);
    assign outputs[2407] = (layer0_outputs[6844]) ^ (layer0_outputs[7395]);
    assign outputs[2408] = layer0_outputs[3818];
    assign outputs[2409] = ~((layer0_outputs[4800]) ^ (layer0_outputs[5104]));
    assign outputs[2410] = ~((layer0_outputs[5363]) ^ (layer0_outputs[7042]));
    assign outputs[2411] = ~(layer0_outputs[4744]) | (layer0_outputs[4997]);
    assign outputs[2412] = (layer0_outputs[5751]) | (layer0_outputs[5679]);
    assign outputs[2413] = (layer0_outputs[5276]) & ~(layer0_outputs[4789]);
    assign outputs[2414] = (layer0_outputs[4665]) & ~(layer0_outputs[5109]);
    assign outputs[2415] = (layer0_outputs[4680]) ^ (layer0_outputs[5969]);
    assign outputs[2416] = ~(layer0_outputs[6876]);
    assign outputs[2417] = ~((layer0_outputs[5763]) & (layer0_outputs[5804]));
    assign outputs[2418] = (layer0_outputs[6592]) ^ (layer0_outputs[7086]);
    assign outputs[2419] = (layer0_outputs[6895]) | (layer0_outputs[1250]);
    assign outputs[2420] = (layer0_outputs[7507]) & ~(layer0_outputs[1294]);
    assign outputs[2421] = ~((layer0_outputs[1848]) ^ (layer0_outputs[7548]));
    assign outputs[2422] = ~(layer0_outputs[2743]);
    assign outputs[2423] = ~(layer0_outputs[171]);
    assign outputs[2424] = layer0_outputs[961];
    assign outputs[2425] = ~(layer0_outputs[4301]);
    assign outputs[2426] = layer0_outputs[5298];
    assign outputs[2427] = (layer0_outputs[878]) ^ (layer0_outputs[6312]);
    assign outputs[2428] = ~(layer0_outputs[3200]);
    assign outputs[2429] = ~(layer0_outputs[7620]) | (layer0_outputs[6484]);
    assign outputs[2430] = 1'b1;
    assign outputs[2431] = ~(layer0_outputs[2124]) | (layer0_outputs[948]);
    assign outputs[2432] = (layer0_outputs[5649]) & (layer0_outputs[1962]);
    assign outputs[2433] = layer0_outputs[6643];
    assign outputs[2434] = ~(layer0_outputs[3764]) | (layer0_outputs[1]);
    assign outputs[2435] = layer0_outputs[1885];
    assign outputs[2436] = (layer0_outputs[5866]) & ~(layer0_outputs[5533]);
    assign outputs[2437] = ~(layer0_outputs[4307]) | (layer0_outputs[1171]);
    assign outputs[2438] = layer0_outputs[5955];
    assign outputs[2439] = ~((layer0_outputs[3494]) ^ (layer0_outputs[6126]));
    assign outputs[2440] = (layer0_outputs[1731]) ^ (layer0_outputs[3254]);
    assign outputs[2441] = ~(layer0_outputs[886]);
    assign outputs[2442] = (layer0_outputs[3602]) & (layer0_outputs[3535]);
    assign outputs[2443] = (layer0_outputs[5622]) & ~(layer0_outputs[680]);
    assign outputs[2444] = ~(layer0_outputs[1862]);
    assign outputs[2445] = ~(layer0_outputs[4656]);
    assign outputs[2446] = ~(layer0_outputs[3490]);
    assign outputs[2447] = layer0_outputs[6772];
    assign outputs[2448] = 1'b1;
    assign outputs[2449] = (layer0_outputs[2276]) ^ (layer0_outputs[2415]);
    assign outputs[2450] = ~((layer0_outputs[4427]) ^ (layer0_outputs[2669]));
    assign outputs[2451] = ~(layer0_outputs[6288]) | (layer0_outputs[4485]);
    assign outputs[2452] = ~((layer0_outputs[7432]) ^ (layer0_outputs[498]));
    assign outputs[2453] = (layer0_outputs[2966]) ^ (layer0_outputs[3382]);
    assign outputs[2454] = ~(layer0_outputs[5904]);
    assign outputs[2455] = ~((layer0_outputs[7049]) | (layer0_outputs[4226]));
    assign outputs[2456] = layer0_outputs[1394];
    assign outputs[2457] = (layer0_outputs[3158]) ^ (layer0_outputs[1637]);
    assign outputs[2458] = (layer0_outputs[2768]) & ~(layer0_outputs[901]);
    assign outputs[2459] = layer0_outputs[6272];
    assign outputs[2460] = (layer0_outputs[360]) | (layer0_outputs[6788]);
    assign outputs[2461] = (layer0_outputs[4883]) ^ (layer0_outputs[503]);
    assign outputs[2462] = ~(layer0_outputs[868]);
    assign outputs[2463] = ~(layer0_outputs[2824]);
    assign outputs[2464] = ~(layer0_outputs[2945]) | (layer0_outputs[7576]);
    assign outputs[2465] = ~((layer0_outputs[3150]) ^ (layer0_outputs[5872]));
    assign outputs[2466] = ~((layer0_outputs[7381]) ^ (layer0_outputs[737]));
    assign outputs[2467] = ~((layer0_outputs[2333]) ^ (layer0_outputs[7425]));
    assign outputs[2468] = ~((layer0_outputs[49]) & (layer0_outputs[2752]));
    assign outputs[2469] = (layer0_outputs[6606]) ^ (layer0_outputs[5196]);
    assign outputs[2470] = ~((layer0_outputs[785]) ^ (layer0_outputs[2902]));
    assign outputs[2471] = (layer0_outputs[7658]) | (layer0_outputs[5255]);
    assign outputs[2472] = layer0_outputs[2734];
    assign outputs[2473] = layer0_outputs[1442];
    assign outputs[2474] = ~(layer0_outputs[5247]);
    assign outputs[2475] = (layer0_outputs[6302]) ^ (layer0_outputs[6519]);
    assign outputs[2476] = ~(layer0_outputs[6834]) | (layer0_outputs[7605]);
    assign outputs[2477] = ~((layer0_outputs[5661]) ^ (layer0_outputs[3855]));
    assign outputs[2478] = layer0_outputs[6051];
    assign outputs[2479] = ~(layer0_outputs[3344]) | (layer0_outputs[1341]);
    assign outputs[2480] = layer0_outputs[5518];
    assign outputs[2481] = (layer0_outputs[3167]) & ~(layer0_outputs[4239]);
    assign outputs[2482] = layer0_outputs[6241];
    assign outputs[2483] = ~((layer0_outputs[5969]) ^ (layer0_outputs[5928]));
    assign outputs[2484] = ~(layer0_outputs[234]) | (layer0_outputs[1090]);
    assign outputs[2485] = ~(layer0_outputs[3708]) | (layer0_outputs[2974]);
    assign outputs[2486] = ~((layer0_outputs[3530]) ^ (layer0_outputs[3358]));
    assign outputs[2487] = layer0_outputs[2621];
    assign outputs[2488] = 1'b1;
    assign outputs[2489] = ~((layer0_outputs[7435]) & (layer0_outputs[6670]));
    assign outputs[2490] = layer0_outputs[4928];
    assign outputs[2491] = layer0_outputs[5662];
    assign outputs[2492] = ~(layer0_outputs[4326]) | (layer0_outputs[3708]);
    assign outputs[2493] = ~((layer0_outputs[3395]) ^ (layer0_outputs[4255]));
    assign outputs[2494] = (layer0_outputs[7649]) & ~(layer0_outputs[7513]);
    assign outputs[2495] = ~(layer0_outputs[6570]);
    assign outputs[2496] = ~(layer0_outputs[1445]);
    assign outputs[2497] = ~((layer0_outputs[2903]) ^ (layer0_outputs[6342]));
    assign outputs[2498] = (layer0_outputs[4657]) & ~(layer0_outputs[3018]);
    assign outputs[2499] = (layer0_outputs[451]) & (layer0_outputs[1124]);
    assign outputs[2500] = ~(layer0_outputs[1963]);
    assign outputs[2501] = ~((layer0_outputs[846]) ^ (layer0_outputs[668]));
    assign outputs[2502] = (layer0_outputs[7315]) & ~(layer0_outputs[774]);
    assign outputs[2503] = (layer0_outputs[541]) & ~(layer0_outputs[7117]);
    assign outputs[2504] = (layer0_outputs[1563]) & (layer0_outputs[1700]);
    assign outputs[2505] = ~((layer0_outputs[5570]) | (layer0_outputs[3796]));
    assign outputs[2506] = (layer0_outputs[4317]) & ~(layer0_outputs[2942]);
    assign outputs[2507] = (layer0_outputs[5676]) ^ (layer0_outputs[3881]);
    assign outputs[2508] = (layer0_outputs[5438]) & ~(layer0_outputs[3691]);
    assign outputs[2509] = (layer0_outputs[6026]) ^ (layer0_outputs[5207]);
    assign outputs[2510] = (layer0_outputs[2839]) & ~(layer0_outputs[4587]);
    assign outputs[2511] = ~((layer0_outputs[6057]) ^ (layer0_outputs[5134]));
    assign outputs[2512] = ~(layer0_outputs[7424]);
    assign outputs[2513] = ~(layer0_outputs[4297]);
    assign outputs[2514] = ~((layer0_outputs[4295]) | (layer0_outputs[2619]));
    assign outputs[2515] = layer0_outputs[3005];
    assign outputs[2516] = layer0_outputs[1612];
    assign outputs[2517] = layer0_outputs[2797];
    assign outputs[2518] = ~(layer0_outputs[5550]) | (layer0_outputs[6577]);
    assign outputs[2519] = ~(layer0_outputs[4864]);
    assign outputs[2520] = layer0_outputs[3777];
    assign outputs[2521] = ~(layer0_outputs[1351]);
    assign outputs[2522] = layer0_outputs[4973];
    assign outputs[2523] = (layer0_outputs[3610]) & (layer0_outputs[7296]);
    assign outputs[2524] = layer0_outputs[2583];
    assign outputs[2525] = ~(layer0_outputs[1333]) | (layer0_outputs[5323]);
    assign outputs[2526] = ~(layer0_outputs[1161]);
    assign outputs[2527] = ~(layer0_outputs[3730]);
    assign outputs[2528] = ~(layer0_outputs[3909]);
    assign outputs[2529] = ~(layer0_outputs[6157]);
    assign outputs[2530] = ~(layer0_outputs[5356]) | (layer0_outputs[1596]);
    assign outputs[2531] = ~(layer0_outputs[4046]);
    assign outputs[2532] = ~(layer0_outputs[1060]) | (layer0_outputs[1909]);
    assign outputs[2533] = ~(layer0_outputs[1101]) | (layer0_outputs[772]);
    assign outputs[2534] = layer0_outputs[2595];
    assign outputs[2535] = ~(layer0_outputs[1224]);
    assign outputs[2536] = layer0_outputs[2325];
    assign outputs[2537] = (layer0_outputs[2789]) & (layer0_outputs[170]);
    assign outputs[2538] = layer0_outputs[484];
    assign outputs[2539] = ~(layer0_outputs[4581]);
    assign outputs[2540] = ~(layer0_outputs[1213]);
    assign outputs[2541] = (layer0_outputs[2696]) & ~(layer0_outputs[4422]);
    assign outputs[2542] = 1'b1;
    assign outputs[2543] = (layer0_outputs[7041]) | (layer0_outputs[5751]);
    assign outputs[2544] = ~(layer0_outputs[3634]) | (layer0_outputs[3537]);
    assign outputs[2545] = layer0_outputs[1638];
    assign outputs[2546] = (layer0_outputs[3964]) & ~(layer0_outputs[5905]);
    assign outputs[2547] = ~((layer0_outputs[7575]) | (layer0_outputs[1763]));
    assign outputs[2548] = ~(layer0_outputs[4519]) | (layer0_outputs[4285]);
    assign outputs[2549] = layer0_outputs[5246];
    assign outputs[2550] = (layer0_outputs[1965]) ^ (layer0_outputs[4064]);
    assign outputs[2551] = ~(layer0_outputs[4000]);
    assign outputs[2552] = ~(layer0_outputs[582]);
    assign outputs[2553] = (layer0_outputs[6817]) & ~(layer0_outputs[1775]);
    assign outputs[2554] = layer0_outputs[7329];
    assign outputs[2555] = ~((layer0_outputs[4913]) & (layer0_outputs[23]));
    assign outputs[2556] = ~(layer0_outputs[469]);
    assign outputs[2557] = layer0_outputs[676];
    assign outputs[2558] = ~((layer0_outputs[7491]) ^ (layer0_outputs[3342]));
    assign outputs[2559] = ~((layer0_outputs[7125]) & (layer0_outputs[520]));
    assign outputs[2560] = layer0_outputs[2189];
    assign outputs[2561] = ~((layer0_outputs[1517]) ^ (layer0_outputs[5833]));
    assign outputs[2562] = layer0_outputs[6424];
    assign outputs[2563] = (layer0_outputs[3478]) ^ (layer0_outputs[1464]);
    assign outputs[2564] = ~(layer0_outputs[5952]);
    assign outputs[2565] = ~(layer0_outputs[1386]) | (layer0_outputs[4479]);
    assign outputs[2566] = layer0_outputs[4631];
    assign outputs[2567] = ~((layer0_outputs[4652]) & (layer0_outputs[1675]));
    assign outputs[2568] = ~(layer0_outputs[6655]) | (layer0_outputs[6225]);
    assign outputs[2569] = layer0_outputs[1922];
    assign outputs[2570] = ~((layer0_outputs[899]) ^ (layer0_outputs[2979]));
    assign outputs[2571] = layer0_outputs[3251];
    assign outputs[2572] = ~((layer0_outputs[5163]) & (layer0_outputs[1828]));
    assign outputs[2573] = ~((layer0_outputs[6640]) ^ (layer0_outputs[4598]));
    assign outputs[2574] = ~(layer0_outputs[4642]);
    assign outputs[2575] = ~((layer0_outputs[2074]) ^ (layer0_outputs[1750]));
    assign outputs[2576] = ~(layer0_outputs[6864]) | (layer0_outputs[4832]);
    assign outputs[2577] = layer0_outputs[6485];
    assign outputs[2578] = (layer0_outputs[616]) ^ (layer0_outputs[2153]);
    assign outputs[2579] = (layer0_outputs[6301]) ^ (layer0_outputs[2740]);
    assign outputs[2580] = ~((layer0_outputs[5414]) & (layer0_outputs[4984]));
    assign outputs[2581] = ~(layer0_outputs[5364]);
    assign outputs[2582] = ~(layer0_outputs[3238]);
    assign outputs[2583] = layer0_outputs[5129];
    assign outputs[2584] = (layer0_outputs[2207]) | (layer0_outputs[3132]);
    assign outputs[2585] = (layer0_outputs[2881]) | (layer0_outputs[3840]);
    assign outputs[2586] = (layer0_outputs[6917]) | (layer0_outputs[2815]);
    assign outputs[2587] = layer0_outputs[5271];
    assign outputs[2588] = (layer0_outputs[3278]) & ~(layer0_outputs[1491]);
    assign outputs[2589] = layer0_outputs[4945];
    assign outputs[2590] = ~((layer0_outputs[7373]) ^ (layer0_outputs[893]));
    assign outputs[2591] = ~(layer0_outputs[6722]);
    assign outputs[2592] = layer0_outputs[7602];
    assign outputs[2593] = (layer0_outputs[6598]) ^ (layer0_outputs[6169]);
    assign outputs[2594] = layer0_outputs[5496];
    assign outputs[2595] = (layer0_outputs[2285]) ^ (layer0_outputs[4055]);
    assign outputs[2596] = layer0_outputs[6612];
    assign outputs[2597] = ~((layer0_outputs[1538]) ^ (layer0_outputs[3120]));
    assign outputs[2598] = ~((layer0_outputs[7589]) & (layer0_outputs[2269]));
    assign outputs[2599] = ~((layer0_outputs[5164]) ^ (layer0_outputs[513]));
    assign outputs[2600] = ~((layer0_outputs[4217]) ^ (layer0_outputs[6600]));
    assign outputs[2601] = (layer0_outputs[6594]) & ~(layer0_outputs[6136]);
    assign outputs[2602] = layer0_outputs[1120];
    assign outputs[2603] = ~((layer0_outputs[4905]) ^ (layer0_outputs[4248]));
    assign outputs[2604] = (layer0_outputs[1325]) & (layer0_outputs[5395]);
    assign outputs[2605] = ~(layer0_outputs[6679]);
    assign outputs[2606] = ~(layer0_outputs[7297]) | (layer0_outputs[5382]);
    assign outputs[2607] = (layer0_outputs[118]) ^ (layer0_outputs[4946]);
    assign outputs[2608] = layer0_outputs[5237];
    assign outputs[2609] = (layer0_outputs[2234]) & ~(layer0_outputs[7630]);
    assign outputs[2610] = ~((layer0_outputs[4669]) ^ (layer0_outputs[7036]));
    assign outputs[2611] = ~(layer0_outputs[2216]);
    assign outputs[2612] = ~(layer0_outputs[1221]);
    assign outputs[2613] = ~(layer0_outputs[2324]);
    assign outputs[2614] = ~((layer0_outputs[3391]) ^ (layer0_outputs[7105]));
    assign outputs[2615] = ~(layer0_outputs[7298]);
    assign outputs[2616] = (layer0_outputs[1992]) & (layer0_outputs[6556]);
    assign outputs[2617] = (layer0_outputs[4785]) & ~(layer0_outputs[505]);
    assign outputs[2618] = ~(layer0_outputs[1170]);
    assign outputs[2619] = (layer0_outputs[6914]) | (layer0_outputs[7286]);
    assign outputs[2620] = layer0_outputs[866];
    assign outputs[2621] = ~(layer0_outputs[2174]);
    assign outputs[2622] = layer0_outputs[2776];
    assign outputs[2623] = ~(layer0_outputs[476]);
    assign outputs[2624] = (layer0_outputs[6828]) ^ (layer0_outputs[169]);
    assign outputs[2625] = (layer0_outputs[5885]) ^ (layer0_outputs[5870]);
    assign outputs[2626] = ~(layer0_outputs[1174]);
    assign outputs[2627] = ~((layer0_outputs[7334]) ^ (layer0_outputs[7057]));
    assign outputs[2628] = layer0_outputs[7342];
    assign outputs[2629] = (layer0_outputs[920]) ^ (layer0_outputs[4483]);
    assign outputs[2630] = layer0_outputs[5553];
    assign outputs[2631] = ~((layer0_outputs[2893]) ^ (layer0_outputs[360]));
    assign outputs[2632] = (layer0_outputs[438]) & ~(layer0_outputs[6634]);
    assign outputs[2633] = layer0_outputs[1744];
    assign outputs[2634] = (layer0_outputs[1329]) & (layer0_outputs[5932]);
    assign outputs[2635] = ~(layer0_outputs[6144]);
    assign outputs[2636] = ~((layer0_outputs[7093]) | (layer0_outputs[2962]));
    assign outputs[2637] = ~((layer0_outputs[5611]) ^ (layer0_outputs[4724]));
    assign outputs[2638] = layer0_outputs[5755];
    assign outputs[2639] = ~(layer0_outputs[452]);
    assign outputs[2640] = ~(layer0_outputs[2712]);
    assign outputs[2641] = (layer0_outputs[4072]) & ~(layer0_outputs[2578]);
    assign outputs[2642] = ~((layer0_outputs[3740]) ^ (layer0_outputs[6820]));
    assign outputs[2643] = ~(layer0_outputs[6877]);
    assign outputs[2644] = ~(layer0_outputs[2210]) | (layer0_outputs[4045]);
    assign outputs[2645] = ~(layer0_outputs[2862]);
    assign outputs[2646] = (layer0_outputs[3850]) & ~(layer0_outputs[5858]);
    assign outputs[2647] = ~((layer0_outputs[1652]) ^ (layer0_outputs[3685]));
    assign outputs[2648] = ~(layer0_outputs[130]);
    assign outputs[2649] = (layer0_outputs[1652]) & ~(layer0_outputs[6421]);
    assign outputs[2650] = layer0_outputs[2692];
    assign outputs[2651] = ~(layer0_outputs[7048]);
    assign outputs[2652] = ~(layer0_outputs[3029]) | (layer0_outputs[5863]);
    assign outputs[2653] = (layer0_outputs[1456]) ^ (layer0_outputs[7527]);
    assign outputs[2654] = (layer0_outputs[1074]) & ~(layer0_outputs[6618]);
    assign outputs[2655] = layer0_outputs[4636];
    assign outputs[2656] = ~(layer0_outputs[3344]) | (layer0_outputs[7573]);
    assign outputs[2657] = (layer0_outputs[6739]) ^ (layer0_outputs[303]);
    assign outputs[2658] = layer0_outputs[518];
    assign outputs[2659] = ~((layer0_outputs[1509]) ^ (layer0_outputs[1318]));
    assign outputs[2660] = ~((layer0_outputs[93]) | (layer0_outputs[4114]));
    assign outputs[2661] = ~(layer0_outputs[1167]);
    assign outputs[2662] = layer0_outputs[6635];
    assign outputs[2663] = ~((layer0_outputs[4506]) ^ (layer0_outputs[2473]));
    assign outputs[2664] = ~((layer0_outputs[3771]) & (layer0_outputs[6961]));
    assign outputs[2665] = ~((layer0_outputs[5538]) ^ (layer0_outputs[5475]));
    assign outputs[2666] = (layer0_outputs[3056]) & ~(layer0_outputs[6791]);
    assign outputs[2667] = ~((layer0_outputs[2949]) | (layer0_outputs[4736]));
    assign outputs[2668] = (layer0_outputs[2507]) ^ (layer0_outputs[3287]);
    assign outputs[2669] = layer0_outputs[4008];
    assign outputs[2670] = layer0_outputs[2094];
    assign outputs[2671] = ~(layer0_outputs[4504]);
    assign outputs[2672] = layer0_outputs[2406];
    assign outputs[2673] = ~(layer0_outputs[2938]);
    assign outputs[2674] = 1'b1;
    assign outputs[2675] = (layer0_outputs[2704]) ^ (layer0_outputs[3564]);
    assign outputs[2676] = 1'b1;
    assign outputs[2677] = (layer0_outputs[807]) ^ (layer0_outputs[5314]);
    assign outputs[2678] = ~(layer0_outputs[7144]);
    assign outputs[2679] = ~(layer0_outputs[773]);
    assign outputs[2680] = ~((layer0_outputs[3059]) ^ (layer0_outputs[5058]));
    assign outputs[2681] = ~(layer0_outputs[7453]) | (layer0_outputs[6958]);
    assign outputs[2682] = ~((layer0_outputs[5991]) & (layer0_outputs[500]));
    assign outputs[2683] = (layer0_outputs[6572]) ^ (layer0_outputs[6103]);
    assign outputs[2684] = ~(layer0_outputs[1537]);
    assign outputs[2685] = ~((layer0_outputs[3223]) ^ (layer0_outputs[931]));
    assign outputs[2686] = (layer0_outputs[3319]) ^ (layer0_outputs[6991]);
    assign outputs[2687] = ~(layer0_outputs[7181]);
    assign outputs[2688] = ~(layer0_outputs[6113]) | (layer0_outputs[4255]);
    assign outputs[2689] = layer0_outputs[7648];
    assign outputs[2690] = ~(layer0_outputs[6040]);
    assign outputs[2691] = (layer0_outputs[1545]) ^ (layer0_outputs[1072]);
    assign outputs[2692] = (layer0_outputs[5671]) | (layer0_outputs[3247]);
    assign outputs[2693] = ~((layer0_outputs[1386]) | (layer0_outputs[5876]));
    assign outputs[2694] = layer0_outputs[3318];
    assign outputs[2695] = ~(layer0_outputs[5719]);
    assign outputs[2696] = (layer0_outputs[701]) | (layer0_outputs[3090]);
    assign outputs[2697] = ~((layer0_outputs[2363]) ^ (layer0_outputs[1944]));
    assign outputs[2698] = (layer0_outputs[456]) | (layer0_outputs[74]);
    assign outputs[2699] = layer0_outputs[6584];
    assign outputs[2700] = (layer0_outputs[3734]) ^ (layer0_outputs[718]);
    assign outputs[2701] = ~(layer0_outputs[4626]);
    assign outputs[2702] = ~(layer0_outputs[298]) | (layer0_outputs[1573]);
    assign outputs[2703] = (layer0_outputs[6462]) ^ (layer0_outputs[5883]);
    assign outputs[2704] = (layer0_outputs[7194]) ^ (layer0_outputs[2728]);
    assign outputs[2705] = ~(layer0_outputs[7362]);
    assign outputs[2706] = ~(layer0_outputs[693]);
    assign outputs[2707] = layer0_outputs[3163];
    assign outputs[2708] = ~((layer0_outputs[5808]) ^ (layer0_outputs[851]));
    assign outputs[2709] = layer0_outputs[1404];
    assign outputs[2710] = (layer0_outputs[4181]) & ~(layer0_outputs[4295]);
    assign outputs[2711] = ~(layer0_outputs[910]) | (layer0_outputs[371]);
    assign outputs[2712] = (layer0_outputs[1071]) ^ (layer0_outputs[3149]);
    assign outputs[2713] = ~(layer0_outputs[4508]);
    assign outputs[2714] = (layer0_outputs[576]) ^ (layer0_outputs[1540]);
    assign outputs[2715] = ~(layer0_outputs[7309]);
    assign outputs[2716] = ~(layer0_outputs[132]) | (layer0_outputs[5984]);
    assign outputs[2717] = ~((layer0_outputs[414]) ^ (layer0_outputs[1953]));
    assign outputs[2718] = ~((layer0_outputs[5527]) ^ (layer0_outputs[1088]));
    assign outputs[2719] = layer0_outputs[7387];
    assign outputs[2720] = (layer0_outputs[6090]) | (layer0_outputs[638]);
    assign outputs[2721] = ~((layer0_outputs[5613]) & (layer0_outputs[2743]));
    assign outputs[2722] = ~(layer0_outputs[4071]);
    assign outputs[2723] = layer0_outputs[2140];
    assign outputs[2724] = ~(layer0_outputs[5302]) | (layer0_outputs[1304]);
    assign outputs[2725] = ~((layer0_outputs[7321]) | (layer0_outputs[4139]));
    assign outputs[2726] = layer0_outputs[1666];
    assign outputs[2727] = ~((layer0_outputs[2545]) & (layer0_outputs[131]));
    assign outputs[2728] = (layer0_outputs[4668]) & ~(layer0_outputs[2255]);
    assign outputs[2729] = ~(layer0_outputs[6081]) | (layer0_outputs[7103]);
    assign outputs[2730] = ~((layer0_outputs[3236]) ^ (layer0_outputs[615]));
    assign outputs[2731] = (layer0_outputs[4718]) ^ (layer0_outputs[930]);
    assign outputs[2732] = (layer0_outputs[365]) ^ (layer0_outputs[2036]);
    assign outputs[2733] = ~(layer0_outputs[5179]);
    assign outputs[2734] = (layer0_outputs[6196]) ^ (layer0_outputs[4711]);
    assign outputs[2735] = (layer0_outputs[2433]) & ~(layer0_outputs[4151]);
    assign outputs[2736] = ~((layer0_outputs[1614]) ^ (layer0_outputs[2364]));
    assign outputs[2737] = layer0_outputs[7243];
    assign outputs[2738] = ~((layer0_outputs[4428]) ^ (layer0_outputs[2693]));
    assign outputs[2739] = layer0_outputs[2385];
    assign outputs[2740] = (layer0_outputs[2760]) ^ (layer0_outputs[3800]);
    assign outputs[2741] = ~(layer0_outputs[3831]);
    assign outputs[2742] = ~(layer0_outputs[7347]);
    assign outputs[2743] = ~(layer0_outputs[433]) | (layer0_outputs[5242]);
    assign outputs[2744] = (layer0_outputs[3409]) & ~(layer0_outputs[58]);
    assign outputs[2745] = (layer0_outputs[4280]) & ~(layer0_outputs[3883]);
    assign outputs[2746] = ~(layer0_outputs[7051]);
    assign outputs[2747] = layer0_outputs[6087];
    assign outputs[2748] = (layer0_outputs[95]) & ~(layer0_outputs[3166]);
    assign outputs[2749] = layer0_outputs[6691];
    assign outputs[2750] = ~(layer0_outputs[3130]) | (layer0_outputs[2596]);
    assign outputs[2751] = (layer0_outputs[1539]) ^ (layer0_outputs[1799]);
    assign outputs[2752] = ~((layer0_outputs[5699]) | (layer0_outputs[5868]));
    assign outputs[2753] = ~(layer0_outputs[3951]);
    assign outputs[2754] = (layer0_outputs[5716]) & (layer0_outputs[2744]);
    assign outputs[2755] = layer0_outputs[6285];
    assign outputs[2756] = (layer0_outputs[6371]) & ~(layer0_outputs[5655]);
    assign outputs[2757] = layer0_outputs[4907];
    assign outputs[2758] = (layer0_outputs[4655]) ^ (layer0_outputs[5258]);
    assign outputs[2759] = (layer0_outputs[3368]) ^ (layer0_outputs[3413]);
    assign outputs[2760] = ~(layer0_outputs[5703]);
    assign outputs[2761] = ~((layer0_outputs[3619]) ^ (layer0_outputs[5366]));
    assign outputs[2762] = ~((layer0_outputs[1646]) & (layer0_outputs[5145]));
    assign outputs[2763] = ~(layer0_outputs[586]);
    assign outputs[2764] = layer0_outputs[5161];
    assign outputs[2765] = ~(layer0_outputs[2767]);
    assign outputs[2766] = ~(layer0_outputs[6863]);
    assign outputs[2767] = (layer0_outputs[5493]) & ~(layer0_outputs[7199]);
    assign outputs[2768] = layer0_outputs[5005];
    assign outputs[2769] = layer0_outputs[1082];
    assign outputs[2770] = ~(layer0_outputs[5884]);
    assign outputs[2771] = layer0_outputs[4228];
    assign outputs[2772] = (layer0_outputs[230]) | (layer0_outputs[1428]);
    assign outputs[2773] = layer0_outputs[349];
    assign outputs[2774] = ~(layer0_outputs[5463]);
    assign outputs[2775] = ~(layer0_outputs[3987]) | (layer0_outputs[923]);
    assign outputs[2776] = ~(layer0_outputs[2918]);
    assign outputs[2777] = ~((layer0_outputs[550]) ^ (layer0_outputs[1304]));
    assign outputs[2778] = layer0_outputs[2242];
    assign outputs[2779] = (layer0_outputs[1574]) & ~(layer0_outputs[2571]);
    assign outputs[2780] = layer0_outputs[4748];
    assign outputs[2781] = layer0_outputs[1830];
    assign outputs[2782] = layer0_outputs[5444];
    assign outputs[2783] = ~((layer0_outputs[790]) & (layer0_outputs[2758]));
    assign outputs[2784] = (layer0_outputs[4427]) ^ (layer0_outputs[4404]);
    assign outputs[2785] = (layer0_outputs[1852]) & ~(layer0_outputs[2662]);
    assign outputs[2786] = (layer0_outputs[7256]) ^ (layer0_outputs[7]);
    assign outputs[2787] = layer0_outputs[105];
    assign outputs[2788] = ~(layer0_outputs[5789]) | (layer0_outputs[1022]);
    assign outputs[2789] = layer0_outputs[3019];
    assign outputs[2790] = layer0_outputs[7272];
    assign outputs[2791] = layer0_outputs[5762];
    assign outputs[2792] = ~(layer0_outputs[3284]);
    assign outputs[2793] = ~(layer0_outputs[7199]) | (layer0_outputs[345]);
    assign outputs[2794] = ~((layer0_outputs[5444]) ^ (layer0_outputs[5142]));
    assign outputs[2795] = ~(layer0_outputs[7521]) | (layer0_outputs[4807]);
    assign outputs[2796] = (layer0_outputs[4906]) ^ (layer0_outputs[7023]);
    assign outputs[2797] = (layer0_outputs[1604]) & ~(layer0_outputs[7205]);
    assign outputs[2798] = ~(layer0_outputs[4942]);
    assign outputs[2799] = layer0_outputs[5783];
    assign outputs[2800] = ~((layer0_outputs[1785]) ^ (layer0_outputs[7260]));
    assign outputs[2801] = (layer0_outputs[1667]) ^ (layer0_outputs[993]);
    assign outputs[2802] = (layer0_outputs[2824]) ^ (layer0_outputs[1957]);
    assign outputs[2803] = (layer0_outputs[6670]) ^ (layer0_outputs[6355]);
    assign outputs[2804] = (layer0_outputs[6516]) | (layer0_outputs[314]);
    assign outputs[2805] = (layer0_outputs[7420]) ^ (layer0_outputs[786]);
    assign outputs[2806] = ~(layer0_outputs[1670]) | (layer0_outputs[4037]);
    assign outputs[2807] = ~(layer0_outputs[3069]);
    assign outputs[2808] = (layer0_outputs[3227]) & ~(layer0_outputs[4058]);
    assign outputs[2809] = ~(layer0_outputs[4382]) | (layer0_outputs[6710]);
    assign outputs[2810] = ~(layer0_outputs[7043]) | (layer0_outputs[2651]);
    assign outputs[2811] = ~(layer0_outputs[7178]);
    assign outputs[2812] = (layer0_outputs[3895]) & (layer0_outputs[1074]);
    assign outputs[2813] = ~(layer0_outputs[5575]);
    assign outputs[2814] = ~(layer0_outputs[4728]);
    assign outputs[2815] = ~((layer0_outputs[7122]) | (layer0_outputs[1943]));
    assign outputs[2816] = ~((layer0_outputs[4585]) & (layer0_outputs[765]));
    assign outputs[2817] = ~(layer0_outputs[1321]) | (layer0_outputs[756]);
    assign outputs[2818] = (layer0_outputs[5177]) & ~(layer0_outputs[6126]);
    assign outputs[2819] = layer0_outputs[6452];
    assign outputs[2820] = layer0_outputs[6657];
    assign outputs[2821] = ~(layer0_outputs[38]);
    assign outputs[2822] = (layer0_outputs[6711]) ^ (layer0_outputs[2878]);
    assign outputs[2823] = ~(layer0_outputs[2798]);
    assign outputs[2824] = layer0_outputs[2599];
    assign outputs[2825] = (layer0_outputs[4694]) ^ (layer0_outputs[4528]);
    assign outputs[2826] = ~((layer0_outputs[3467]) & (layer0_outputs[1850]));
    assign outputs[2827] = ~((layer0_outputs[1037]) ^ (layer0_outputs[5525]));
    assign outputs[2828] = ~(layer0_outputs[6122]);
    assign outputs[2829] = ~(layer0_outputs[4798]);
    assign outputs[2830] = ~(layer0_outputs[6392]) | (layer0_outputs[7245]);
    assign outputs[2831] = ~(layer0_outputs[5703]);
    assign outputs[2832] = ~(layer0_outputs[1566]) | (layer0_outputs[3969]);
    assign outputs[2833] = ~((layer0_outputs[602]) & (layer0_outputs[1449]));
    assign outputs[2834] = (layer0_outputs[1941]) ^ (layer0_outputs[5054]);
    assign outputs[2835] = layer0_outputs[3453];
    assign outputs[2836] = ~(layer0_outputs[2911]);
    assign outputs[2837] = (layer0_outputs[6788]) & ~(layer0_outputs[469]);
    assign outputs[2838] = (layer0_outputs[3768]) & (layer0_outputs[2270]);
    assign outputs[2839] = layer0_outputs[229];
    assign outputs[2840] = ~(layer0_outputs[1607]);
    assign outputs[2841] = layer0_outputs[2088];
    assign outputs[2842] = layer0_outputs[4767];
    assign outputs[2843] = layer0_outputs[4977];
    assign outputs[2844] = (layer0_outputs[1870]) & ~(layer0_outputs[5843]);
    assign outputs[2845] = (layer0_outputs[1734]) & ~(layer0_outputs[2664]);
    assign outputs[2846] = layer0_outputs[5524];
    assign outputs[2847] = layer0_outputs[7381];
    assign outputs[2848] = layer0_outputs[4574];
    assign outputs[2849] = ~(layer0_outputs[4691]);
    assign outputs[2850] = ~((layer0_outputs[863]) & (layer0_outputs[1209]));
    assign outputs[2851] = ~(layer0_outputs[2995]);
    assign outputs[2852] = ~((layer0_outputs[3506]) ^ (layer0_outputs[2330]));
    assign outputs[2853] = ~(layer0_outputs[6842]);
    assign outputs[2854] = ~(layer0_outputs[5760]);
    assign outputs[2855] = ~((layer0_outputs[1578]) & (layer0_outputs[4527]));
    assign outputs[2856] = ~((layer0_outputs[7337]) ^ (layer0_outputs[6436]));
    assign outputs[2857] = layer0_outputs[3339];
    assign outputs[2858] = ~(layer0_outputs[5413]);
    assign outputs[2859] = layer0_outputs[4209];
    assign outputs[2860] = ~(layer0_outputs[5241]);
    assign outputs[2861] = ~(layer0_outputs[5814]);
    assign outputs[2862] = ~(layer0_outputs[5882]);
    assign outputs[2863] = (layer0_outputs[5412]) ^ (layer0_outputs[1867]);
    assign outputs[2864] = layer0_outputs[7632];
    assign outputs[2865] = (layer0_outputs[826]) & ~(layer0_outputs[7349]);
    assign outputs[2866] = (layer0_outputs[2065]) | (layer0_outputs[754]);
    assign outputs[2867] = ~(layer0_outputs[246]);
    assign outputs[2868] = layer0_outputs[5975];
    assign outputs[2869] = ~((layer0_outputs[3869]) | (layer0_outputs[4306]));
    assign outputs[2870] = ~(layer0_outputs[250]);
    assign outputs[2871] = ~((layer0_outputs[2272]) ^ (layer0_outputs[519]));
    assign outputs[2872] = ~(layer0_outputs[6420]);
    assign outputs[2873] = layer0_outputs[5537];
    assign outputs[2874] = ~((layer0_outputs[7479]) ^ (layer0_outputs[7247]));
    assign outputs[2875] = (layer0_outputs[4148]) & ~(layer0_outputs[7338]);
    assign outputs[2876] = ~((layer0_outputs[1688]) & (layer0_outputs[5699]));
    assign outputs[2877] = ~(layer0_outputs[11]);
    assign outputs[2878] = ~((layer0_outputs[7180]) ^ (layer0_outputs[724]));
    assign outputs[2879] = (layer0_outputs[5362]) & (layer0_outputs[1496]);
    assign outputs[2880] = ~(layer0_outputs[6394]);
    assign outputs[2881] = ~((layer0_outputs[6910]) ^ (layer0_outputs[5785]));
    assign outputs[2882] = ~((layer0_outputs[6663]) | (layer0_outputs[2858]));
    assign outputs[2883] = ~(layer0_outputs[6131]) | (layer0_outputs[7074]);
    assign outputs[2884] = (layer0_outputs[5262]) & ~(layer0_outputs[499]);
    assign outputs[2885] = ~(layer0_outputs[7302]);
    assign outputs[2886] = ~(layer0_outputs[1007]);
    assign outputs[2887] = layer0_outputs[2224];
    assign outputs[2888] = (layer0_outputs[1511]) & ~(layer0_outputs[4778]);
    assign outputs[2889] = ~((layer0_outputs[4573]) ^ (layer0_outputs[7156]));
    assign outputs[2890] = ~((layer0_outputs[2716]) & (layer0_outputs[7337]));
    assign outputs[2891] = ~(layer0_outputs[5328]) | (layer0_outputs[4165]);
    assign outputs[2892] = layer0_outputs[1877];
    assign outputs[2893] = 1'b1;
    assign outputs[2894] = (layer0_outputs[5001]) | (layer0_outputs[1647]);
    assign outputs[2895] = ~(layer0_outputs[978]) | (layer0_outputs[867]);
    assign outputs[2896] = (layer0_outputs[541]) & ~(layer0_outputs[5407]);
    assign outputs[2897] = ~(layer0_outputs[4855]) | (layer0_outputs[1912]);
    assign outputs[2898] = ~((layer0_outputs[759]) ^ (layer0_outputs[138]));
    assign outputs[2899] = ~(layer0_outputs[1688]);
    assign outputs[2900] = layer0_outputs[7533];
    assign outputs[2901] = ~(layer0_outputs[5166]);
    assign outputs[2902] = ~(layer0_outputs[6962]);
    assign outputs[2903] = ~(layer0_outputs[3863]) | (layer0_outputs[1250]);
    assign outputs[2904] = (layer0_outputs[6177]) ^ (layer0_outputs[1730]);
    assign outputs[2905] = ~((layer0_outputs[2372]) ^ (layer0_outputs[6732]));
    assign outputs[2906] = layer0_outputs[3775];
    assign outputs[2907] = ~(layer0_outputs[5888]);
    assign outputs[2908] = layer0_outputs[3484];
    assign outputs[2909] = ~(layer0_outputs[5338]);
    assign outputs[2910] = (layer0_outputs[1153]) & (layer0_outputs[375]);
    assign outputs[2911] = ~(layer0_outputs[6372]);
    assign outputs[2912] = ~((layer0_outputs[2516]) ^ (layer0_outputs[7411]));
    assign outputs[2913] = (layer0_outputs[2357]) & ~(layer0_outputs[6120]);
    assign outputs[2914] = (layer0_outputs[576]) & ~(layer0_outputs[6004]);
    assign outputs[2915] = layer0_outputs[1870];
    assign outputs[2916] = (layer0_outputs[3004]) ^ (layer0_outputs[4238]);
    assign outputs[2917] = (layer0_outputs[222]) & (layer0_outputs[6234]);
    assign outputs[2918] = (layer0_outputs[835]) | (layer0_outputs[2950]);
    assign outputs[2919] = ~((layer0_outputs[1355]) & (layer0_outputs[6404]));
    assign outputs[2920] = ~(layer0_outputs[5054]) | (layer0_outputs[27]);
    assign outputs[2921] = ~(layer0_outputs[7669]);
    assign outputs[2922] = ~(layer0_outputs[4071]);
    assign outputs[2923] = layer0_outputs[4272];
    assign outputs[2924] = (layer0_outputs[1792]) ^ (layer0_outputs[1031]);
    assign outputs[2925] = (layer0_outputs[162]) & (layer0_outputs[1932]);
    assign outputs[2926] = ~((layer0_outputs[6390]) ^ (layer0_outputs[443]));
    assign outputs[2927] = layer0_outputs[7169];
    assign outputs[2928] = ~(layer0_outputs[6149]);
    assign outputs[2929] = (layer0_outputs[1575]) & ~(layer0_outputs[539]);
    assign outputs[2930] = (layer0_outputs[3599]) ^ (layer0_outputs[4910]);
    assign outputs[2931] = layer0_outputs[5775];
    assign outputs[2932] = layer0_outputs[955];
    assign outputs[2933] = (layer0_outputs[6838]) ^ (layer0_outputs[1913]);
    assign outputs[2934] = ~(layer0_outputs[6118]);
    assign outputs[2935] = ~((layer0_outputs[190]) ^ (layer0_outputs[4124]));
    assign outputs[2936] = (layer0_outputs[5847]) ^ (layer0_outputs[3507]);
    assign outputs[2937] = ~((layer0_outputs[1998]) & (layer0_outputs[5197]));
    assign outputs[2938] = layer0_outputs[2178];
    assign outputs[2939] = layer0_outputs[1558];
    assign outputs[2940] = (layer0_outputs[411]) & (layer0_outputs[1217]);
    assign outputs[2941] = layer0_outputs[5009];
    assign outputs[2942] = layer0_outputs[6097];
    assign outputs[2943] = (layer0_outputs[6293]) ^ (layer0_outputs[1805]);
    assign outputs[2944] = layer0_outputs[3272];
    assign outputs[2945] = layer0_outputs[4974];
    assign outputs[2946] = layer0_outputs[5008];
    assign outputs[2947] = (layer0_outputs[1502]) ^ (layer0_outputs[5997]);
    assign outputs[2948] = ~(layer0_outputs[6038]) | (layer0_outputs[4811]);
    assign outputs[2949] = ~(layer0_outputs[4525]);
    assign outputs[2950] = ~((layer0_outputs[5090]) ^ (layer0_outputs[7211]));
    assign outputs[2951] = (layer0_outputs[5416]) & (layer0_outputs[1162]);
    assign outputs[2952] = layer0_outputs[1404];
    assign outputs[2953] = (layer0_outputs[254]) & ~(layer0_outputs[7586]);
    assign outputs[2954] = ~(layer0_outputs[1821]);
    assign outputs[2955] = (layer0_outputs[3357]) ^ (layer0_outputs[3929]);
    assign outputs[2956] = (layer0_outputs[4147]) & ~(layer0_outputs[4055]);
    assign outputs[2957] = ~((layer0_outputs[2315]) ^ (layer0_outputs[2897]));
    assign outputs[2958] = layer0_outputs[3351];
    assign outputs[2959] = ~(layer0_outputs[3861]);
    assign outputs[2960] = (layer0_outputs[335]) & ~(layer0_outputs[2615]);
    assign outputs[2961] = ~(layer0_outputs[1979]);
    assign outputs[2962] = ~(layer0_outputs[7409]) | (layer0_outputs[1883]);
    assign outputs[2963] = ~(layer0_outputs[3383]);
    assign outputs[2964] = ~(layer0_outputs[2204]);
    assign outputs[2965] = ~(layer0_outputs[6171]) | (layer0_outputs[5250]);
    assign outputs[2966] = ~((layer0_outputs[5103]) | (layer0_outputs[3698]));
    assign outputs[2967] = (layer0_outputs[2612]) ^ (layer0_outputs[5917]);
    assign outputs[2968] = layer0_outputs[6642];
    assign outputs[2969] = (layer0_outputs[4061]) & (layer0_outputs[922]);
    assign outputs[2970] = (layer0_outputs[7046]) & ~(layer0_outputs[2742]);
    assign outputs[2971] = ~((layer0_outputs[4616]) ^ (layer0_outputs[1204]));
    assign outputs[2972] = layer0_outputs[5048];
    assign outputs[2973] = layer0_outputs[7328];
    assign outputs[2974] = layer0_outputs[2291];
    assign outputs[2975] = ~((layer0_outputs[2271]) ^ (layer0_outputs[844]));
    assign outputs[2976] = ~(layer0_outputs[3738]);
    assign outputs[2977] = (layer0_outputs[6625]) & ~(layer0_outputs[1381]);
    assign outputs[2978] = ~(layer0_outputs[5525]) | (layer0_outputs[2852]);
    assign outputs[2979] = ~(layer0_outputs[4640]) | (layer0_outputs[5700]);
    assign outputs[2980] = (layer0_outputs[7387]) & ~(layer0_outputs[2783]);
    assign outputs[2981] = layer0_outputs[29];
    assign outputs[2982] = ~(layer0_outputs[6977]);
    assign outputs[2983] = (layer0_outputs[337]) ^ (layer0_outputs[3280]);
    assign outputs[2984] = ~((layer0_outputs[1154]) ^ (layer0_outputs[2503]));
    assign outputs[2985] = ~(layer0_outputs[3919]);
    assign outputs[2986] = ~(layer0_outputs[1681]);
    assign outputs[2987] = layer0_outputs[5617];
    assign outputs[2988] = ~((layer0_outputs[1314]) & (layer0_outputs[2660]));
    assign outputs[2989] = (layer0_outputs[2005]) ^ (layer0_outputs[1564]);
    assign outputs[2990] = ~(layer0_outputs[4953]);
    assign outputs[2991] = layer0_outputs[7164];
    assign outputs[2992] = ~(layer0_outputs[3567]);
    assign outputs[2993] = ~(layer0_outputs[3894]) | (layer0_outputs[3296]);
    assign outputs[2994] = ~((layer0_outputs[7369]) & (layer0_outputs[4665]));
    assign outputs[2995] = layer0_outputs[1342];
    assign outputs[2996] = ~((layer0_outputs[1815]) ^ (layer0_outputs[5818]));
    assign outputs[2997] = ~(layer0_outputs[5665]);
    assign outputs[2998] = ~((layer0_outputs[7512]) ^ (layer0_outputs[827]));
    assign outputs[2999] = ~(layer0_outputs[6662]) | (layer0_outputs[5374]);
    assign outputs[3000] = layer0_outputs[7175];
    assign outputs[3001] = ~(layer0_outputs[3169]);
    assign outputs[3002] = (layer0_outputs[1635]) & ~(layer0_outputs[6394]);
    assign outputs[3003] = (layer0_outputs[5583]) ^ (layer0_outputs[6872]);
    assign outputs[3004] = (layer0_outputs[4077]) & ~(layer0_outputs[7180]);
    assign outputs[3005] = ~(layer0_outputs[5944]);
    assign outputs[3006] = layer0_outputs[3299];
    assign outputs[3007] = ~(layer0_outputs[1795]) | (layer0_outputs[6315]);
    assign outputs[3008] = (layer0_outputs[4428]) | (layer0_outputs[2368]);
    assign outputs[3009] = (layer0_outputs[4048]) ^ (layer0_outputs[2993]);
    assign outputs[3010] = layer0_outputs[4103];
    assign outputs[3011] = layer0_outputs[2535];
    assign outputs[3012] = ~(layer0_outputs[364]);
    assign outputs[3013] = (layer0_outputs[7198]) & ~(layer0_outputs[2890]);
    assign outputs[3014] = layer0_outputs[6235];
    assign outputs[3015] = (layer0_outputs[3419]) & ~(layer0_outputs[4343]);
    assign outputs[3016] = ~(layer0_outputs[2208]);
    assign outputs[3017] = layer0_outputs[4171];
    assign outputs[3018] = ~(layer0_outputs[4446]);
    assign outputs[3019] = layer0_outputs[4726];
    assign outputs[3020] = layer0_outputs[6717];
    assign outputs[3021] = ~(layer0_outputs[3987]);
    assign outputs[3022] = ~((layer0_outputs[5944]) ^ (layer0_outputs[6663]));
    assign outputs[3023] = layer0_outputs[6830];
    assign outputs[3024] = ~((layer0_outputs[3044]) | (layer0_outputs[3060]));
    assign outputs[3025] = (layer0_outputs[1085]) ^ (layer0_outputs[5113]);
    assign outputs[3026] = ~((layer0_outputs[18]) ^ (layer0_outputs[1068]));
    assign outputs[3027] = ~((layer0_outputs[358]) ^ (layer0_outputs[1350]));
    assign outputs[3028] = ~(layer0_outputs[578]);
    assign outputs[3029] = layer0_outputs[6538];
    assign outputs[3030] = layer0_outputs[2478];
    assign outputs[3031] = ~(layer0_outputs[3428]);
    assign outputs[3032] = ~(layer0_outputs[1640]);
    assign outputs[3033] = (layer0_outputs[3401]) ^ (layer0_outputs[2939]);
    assign outputs[3034] = ~(layer0_outputs[2392]) | (layer0_outputs[6604]);
    assign outputs[3035] = ~((layer0_outputs[7038]) ^ (layer0_outputs[2303]));
    assign outputs[3036] = (layer0_outputs[1306]) & ~(layer0_outputs[1034]);
    assign outputs[3037] = ~(layer0_outputs[1152]);
    assign outputs[3038] = (layer0_outputs[2567]) ^ (layer0_outputs[273]);
    assign outputs[3039] = layer0_outputs[723];
    assign outputs[3040] = ~((layer0_outputs[6340]) ^ (layer0_outputs[3167]));
    assign outputs[3041] = (layer0_outputs[1644]) & (layer0_outputs[2593]);
    assign outputs[3042] = ~((layer0_outputs[2337]) ^ (layer0_outputs[1214]));
    assign outputs[3043] = ~(layer0_outputs[886]);
    assign outputs[3044] = ~((layer0_outputs[5421]) ^ (layer0_outputs[4156]));
    assign outputs[3045] = (layer0_outputs[4161]) ^ (layer0_outputs[2237]);
    assign outputs[3046] = ~(layer0_outputs[2628]) | (layer0_outputs[4612]);
    assign outputs[3047] = ~(layer0_outputs[7152]) | (layer0_outputs[6181]);
    assign outputs[3048] = (layer0_outputs[2070]) & (layer0_outputs[686]);
    assign outputs[3049] = (layer0_outputs[890]) ^ (layer0_outputs[1740]);
    assign outputs[3050] = ~((layer0_outputs[6058]) ^ (layer0_outputs[1868]));
    assign outputs[3051] = ~(layer0_outputs[91]);
    assign outputs[3052] = ~(layer0_outputs[1095]) | (layer0_outputs[2533]);
    assign outputs[3053] = layer0_outputs[6236];
    assign outputs[3054] = (layer0_outputs[7139]) & ~(layer0_outputs[410]);
    assign outputs[3055] = (layer0_outputs[4478]) | (layer0_outputs[4841]);
    assign outputs[3056] = ~((layer0_outputs[4446]) ^ (layer0_outputs[314]));
    assign outputs[3057] = ~((layer0_outputs[2592]) & (layer0_outputs[470]));
    assign outputs[3058] = ~(layer0_outputs[6985]);
    assign outputs[3059] = ~((layer0_outputs[374]) ^ (layer0_outputs[5925]));
    assign outputs[3060] = layer0_outputs[5838];
    assign outputs[3061] = ~((layer0_outputs[1256]) ^ (layer0_outputs[811]));
    assign outputs[3062] = ~((layer0_outputs[306]) ^ (layer0_outputs[7052]));
    assign outputs[3063] = ~((layer0_outputs[4883]) ^ (layer0_outputs[1350]));
    assign outputs[3064] = ~(layer0_outputs[302]);
    assign outputs[3065] = ~(layer0_outputs[6460]);
    assign outputs[3066] = (layer0_outputs[6838]) & (layer0_outputs[2909]);
    assign outputs[3067] = (layer0_outputs[5277]) ^ (layer0_outputs[1249]);
    assign outputs[3068] = layer0_outputs[4409];
    assign outputs[3069] = ~((layer0_outputs[4779]) ^ (layer0_outputs[4089]));
    assign outputs[3070] = ~(layer0_outputs[1824]) | (layer0_outputs[795]);
    assign outputs[3071] = (layer0_outputs[2908]) ^ (layer0_outputs[5894]);
    assign outputs[3072] = (layer0_outputs[2995]) & ~(layer0_outputs[2278]);
    assign outputs[3073] = ~((layer0_outputs[3875]) | (layer0_outputs[5056]));
    assign outputs[3074] = (layer0_outputs[2182]) & ~(layer0_outputs[5424]);
    assign outputs[3075] = ~((layer0_outputs[7492]) ^ (layer0_outputs[4369]));
    assign outputs[3076] = ~((layer0_outputs[6641]) | (layer0_outputs[1678]));
    assign outputs[3077] = ~(layer0_outputs[6412]);
    assign outputs[3078] = ~(layer0_outputs[5412]);
    assign outputs[3079] = layer0_outputs[644];
    assign outputs[3080] = layer0_outputs[1161];
    assign outputs[3081] = ~(layer0_outputs[1270]);
    assign outputs[3082] = layer0_outputs[7011];
    assign outputs[3083] = layer0_outputs[4024];
    assign outputs[3084] = ~(layer0_outputs[6764]);
    assign outputs[3085] = layer0_outputs[1623];
    assign outputs[3086] = ~(layer0_outputs[2459]);
    assign outputs[3087] = (layer0_outputs[6147]) ^ (layer0_outputs[7482]);
    assign outputs[3088] = ~(layer0_outputs[2632]);
    assign outputs[3089] = (layer0_outputs[5598]) ^ (layer0_outputs[3992]);
    assign outputs[3090] = (layer0_outputs[5469]) & ~(layer0_outputs[6749]);
    assign outputs[3091] = layer0_outputs[3066];
    assign outputs[3092] = (layer0_outputs[2682]) & ~(layer0_outputs[5317]);
    assign outputs[3093] = ~((layer0_outputs[7466]) | (layer0_outputs[7383]));
    assign outputs[3094] = (layer0_outputs[3535]) & ~(layer0_outputs[7462]);
    assign outputs[3095] = ~(layer0_outputs[6176]);
    assign outputs[3096] = (layer0_outputs[2229]) & ~(layer0_outputs[3522]);
    assign outputs[3097] = ~((layer0_outputs[4766]) ^ (layer0_outputs[3266]));
    assign outputs[3098] = (layer0_outputs[7450]) & (layer0_outputs[7189]);
    assign outputs[3099] = ~((layer0_outputs[3474]) ^ (layer0_outputs[6642]));
    assign outputs[3100] = ~((layer0_outputs[5350]) | (layer0_outputs[4317]));
    assign outputs[3101] = layer0_outputs[5112];
    assign outputs[3102] = ~(layer0_outputs[2835]);
    assign outputs[3103] = layer0_outputs[2839];
    assign outputs[3104] = ~((layer0_outputs[5194]) ^ (layer0_outputs[2800]));
    assign outputs[3105] = ~(layer0_outputs[45]) | (layer0_outputs[1794]);
    assign outputs[3106] = (layer0_outputs[1524]) & ~(layer0_outputs[1880]);
    assign outputs[3107] = ~((layer0_outputs[1650]) | (layer0_outputs[2799]));
    assign outputs[3108] = (layer0_outputs[4952]) | (layer0_outputs[3207]);
    assign outputs[3109] = ~((layer0_outputs[1914]) ^ (layer0_outputs[7415]));
    assign outputs[3110] = layer0_outputs[180];
    assign outputs[3111] = (layer0_outputs[5939]) & ~(layer0_outputs[6550]);
    assign outputs[3112] = ~(layer0_outputs[6496]) | (layer0_outputs[1387]);
    assign outputs[3113] = ~((layer0_outputs[7229]) | (layer0_outputs[2961]));
    assign outputs[3114] = ~((layer0_outputs[4011]) ^ (layer0_outputs[333]));
    assign outputs[3115] = (layer0_outputs[5721]) ^ (layer0_outputs[2282]);
    assign outputs[3116] = ~(layer0_outputs[5725]);
    assign outputs[3117] = (layer0_outputs[7450]) ^ (layer0_outputs[1113]);
    assign outputs[3118] = ~((layer0_outputs[941]) ^ (layer0_outputs[7489]));
    assign outputs[3119] = layer0_outputs[3843];
    assign outputs[3120] = ~((layer0_outputs[5322]) & (layer0_outputs[3667]));
    assign outputs[3121] = (layer0_outputs[5831]) ^ (layer0_outputs[3380]);
    assign outputs[3122] = (layer0_outputs[5806]) & (layer0_outputs[5223]);
    assign outputs[3123] = ~((layer0_outputs[5631]) ^ (layer0_outputs[6504]));
    assign outputs[3124] = ~((layer0_outputs[1323]) | (layer0_outputs[109]));
    assign outputs[3125] = ~((layer0_outputs[6935]) ^ (layer0_outputs[3772]));
    assign outputs[3126] = layer0_outputs[643];
    assign outputs[3127] = ~((layer0_outputs[331]) | (layer0_outputs[2060]));
    assign outputs[3128] = layer0_outputs[5138];
    assign outputs[3129] = ~(layer0_outputs[1464]) | (layer0_outputs[277]);
    assign outputs[3130] = ~((layer0_outputs[1142]) ^ (layer0_outputs[5579]));
    assign outputs[3131] = (layer0_outputs[5464]) | (layer0_outputs[3848]);
    assign outputs[3132] = ~(layer0_outputs[666]);
    assign outputs[3133] = (layer0_outputs[3377]) ^ (layer0_outputs[1928]);
    assign outputs[3134] = ~(layer0_outputs[2361]) | (layer0_outputs[6818]);
    assign outputs[3135] = ~((layer0_outputs[3762]) ^ (layer0_outputs[6154]));
    assign outputs[3136] = ~(layer0_outputs[4167]);
    assign outputs[3137] = ~((layer0_outputs[1788]) ^ (layer0_outputs[4176]));
    assign outputs[3138] = (layer0_outputs[7094]) ^ (layer0_outputs[5585]);
    assign outputs[3139] = ~(layer0_outputs[3285]) | (layer0_outputs[596]);
    assign outputs[3140] = ~(layer0_outputs[159]);
    assign outputs[3141] = ~(layer0_outputs[577]);
    assign outputs[3142] = layer0_outputs[1311];
    assign outputs[3143] = ~((layer0_outputs[4617]) ^ (layer0_outputs[3290]));
    assign outputs[3144] = ~(layer0_outputs[3924]);
    assign outputs[3145] = (layer0_outputs[6238]) & (layer0_outputs[628]);
    assign outputs[3146] = ~((layer0_outputs[1263]) ^ (layer0_outputs[7009]));
    assign outputs[3147] = layer0_outputs[4166];
    assign outputs[3148] = (layer0_outputs[4939]) ^ (layer0_outputs[3755]);
    assign outputs[3149] = ~(layer0_outputs[4996]);
    assign outputs[3150] = (layer0_outputs[6665]) ^ (layer0_outputs[4305]);
    assign outputs[3151] = layer0_outputs[7047];
    assign outputs[3152] = (layer0_outputs[1021]) & ~(layer0_outputs[7501]);
    assign outputs[3153] = layer0_outputs[53];
    assign outputs[3154] = ~((layer0_outputs[4668]) ^ (layer0_outputs[3426]));
    assign outputs[3155] = ~((layer0_outputs[3592]) ^ (layer0_outputs[3290]));
    assign outputs[3156] = ~((layer0_outputs[4741]) | (layer0_outputs[710]));
    assign outputs[3157] = (layer0_outputs[5776]) & ~(layer0_outputs[521]);
    assign outputs[3158] = ~(layer0_outputs[5249]);
    assign outputs[3159] = (layer0_outputs[2913]) | (layer0_outputs[841]);
    assign outputs[3160] = ~(layer0_outputs[7398]) | (layer0_outputs[1617]);
    assign outputs[3161] = layer0_outputs[7537];
    assign outputs[3162] = layer0_outputs[150];
    assign outputs[3163] = (layer0_outputs[918]) & ~(layer0_outputs[2029]);
    assign outputs[3164] = ~(layer0_outputs[6219]) | (layer0_outputs[6702]);
    assign outputs[3165] = layer0_outputs[4140];
    assign outputs[3166] = (layer0_outputs[4043]) & ~(layer0_outputs[4996]);
    assign outputs[3167] = layer0_outputs[2565];
    assign outputs[3168] = (layer0_outputs[5204]) & ~(layer0_outputs[4371]);
    assign outputs[3169] = (layer0_outputs[3092]) & ~(layer0_outputs[1946]);
    assign outputs[3170] = (layer0_outputs[1770]) & ~(layer0_outputs[1764]);
    assign outputs[3171] = layer0_outputs[5857];
    assign outputs[3172] = layer0_outputs[1117];
    assign outputs[3173] = (layer0_outputs[2988]) | (layer0_outputs[2673]);
    assign outputs[3174] = ~((layer0_outputs[7060]) | (layer0_outputs[537]));
    assign outputs[3175] = layer0_outputs[6734];
    assign outputs[3176] = (layer0_outputs[2387]) & (layer0_outputs[2379]);
    assign outputs[3177] = (layer0_outputs[1073]) ^ (layer0_outputs[5243]);
    assign outputs[3178] = (layer0_outputs[247]) & (layer0_outputs[3331]);
    assign outputs[3179] = ~(layer0_outputs[6965]);
    assign outputs[3180] = layer0_outputs[1591];
    assign outputs[3181] = ~((layer0_outputs[142]) ^ (layer0_outputs[2895]));
    assign outputs[3182] = (layer0_outputs[5937]) & ~(layer0_outputs[804]);
    assign outputs[3183] = ~((layer0_outputs[4796]) ^ (layer0_outputs[3943]));
    assign outputs[3184] = layer0_outputs[7096];
    assign outputs[3185] = layer0_outputs[5748];
    assign outputs[3186] = layer0_outputs[7252];
    assign outputs[3187] = (layer0_outputs[1247]) & ~(layer0_outputs[5692]);
    assign outputs[3188] = (layer0_outputs[5469]) ^ (layer0_outputs[1559]);
    assign outputs[3189] = ~(layer0_outputs[4398]);
    assign outputs[3190] = ~((layer0_outputs[3692]) | (layer0_outputs[6878]));
    assign outputs[3191] = layer0_outputs[3857];
    assign outputs[3192] = layer0_outputs[6823];
    assign outputs[3193] = (layer0_outputs[3553]) & (layer0_outputs[6186]);
    assign outputs[3194] = (layer0_outputs[5919]) & ~(layer0_outputs[1784]);
    assign outputs[3195] = (layer0_outputs[1600]) ^ (layer0_outputs[6405]);
    assign outputs[3196] = (layer0_outputs[7268]) & ~(layer0_outputs[3019]);
    assign outputs[3197] = (layer0_outputs[1894]) & ~(layer0_outputs[5996]);
    assign outputs[3198] = ~((layer0_outputs[980]) | (layer0_outputs[4904]));
    assign outputs[3199] = ~(layer0_outputs[5530]);
    assign outputs[3200] = layer0_outputs[6411];
    assign outputs[3201] = (layer0_outputs[7456]) & (layer0_outputs[4494]);
    assign outputs[3202] = ~((layer0_outputs[2176]) ^ (layer0_outputs[1175]));
    assign outputs[3203] = (layer0_outputs[1416]) ^ (layer0_outputs[6268]);
    assign outputs[3204] = ~(layer0_outputs[1723]);
    assign outputs[3205] = ~(layer0_outputs[3412]) | (layer0_outputs[6975]);
    assign outputs[3206] = (layer0_outputs[830]) ^ (layer0_outputs[5958]);
    assign outputs[3207] = ~(layer0_outputs[6198]);
    assign outputs[3208] = ~(layer0_outputs[2634]) | (layer0_outputs[3372]);
    assign outputs[3209] = layer0_outputs[7275];
    assign outputs[3210] = layer0_outputs[4712];
    assign outputs[3211] = layer0_outputs[6455];
    assign outputs[3212] = ~((layer0_outputs[7264]) ^ (layer0_outputs[4922]));
    assign outputs[3213] = (layer0_outputs[3954]) | (layer0_outputs[2390]);
    assign outputs[3214] = ~((layer0_outputs[7278]) ^ (layer0_outputs[2905]));
    assign outputs[3215] = (layer0_outputs[3097]) ^ (layer0_outputs[4036]);
    assign outputs[3216] = ~(layer0_outputs[3491]) | (layer0_outputs[2723]);
    assign outputs[3217] = ~(layer0_outputs[5702]);
    assign outputs[3218] = layer0_outputs[1708];
    assign outputs[3219] = (layer0_outputs[423]) & ~(layer0_outputs[3693]);
    assign outputs[3220] = (layer0_outputs[1347]) ^ (layer0_outputs[5666]);
    assign outputs[3221] = (layer0_outputs[2415]) ^ (layer0_outputs[3967]);
    assign outputs[3222] = (layer0_outputs[831]) ^ (layer0_outputs[7221]);
    assign outputs[3223] = ~((layer0_outputs[2803]) | (layer0_outputs[4661]));
    assign outputs[3224] = (layer0_outputs[6925]) & ~(layer0_outputs[492]);
    assign outputs[3225] = layer0_outputs[958];
    assign outputs[3226] = ~(layer0_outputs[7299]);
    assign outputs[3227] = ~(layer0_outputs[5153]);
    assign outputs[3228] = ~(layer0_outputs[6444]);
    assign outputs[3229] = ~(layer0_outputs[4507]);
    assign outputs[3230] = layer0_outputs[1477];
    assign outputs[3231] = ~(layer0_outputs[3119]);
    assign outputs[3232] = layer0_outputs[4020];
    assign outputs[3233] = (layer0_outputs[384]) & ~(layer0_outputs[5265]);
    assign outputs[3234] = ~((layer0_outputs[2169]) | (layer0_outputs[6993]));
    assign outputs[3235] = (layer0_outputs[5]) ^ (layer0_outputs[4516]);
    assign outputs[3236] = layer0_outputs[4467];
    assign outputs[3237] = ~(layer0_outputs[209]);
    assign outputs[3238] = (layer0_outputs[2519]) ^ (layer0_outputs[6985]);
    assign outputs[3239] = layer0_outputs[3242];
    assign outputs[3240] = layer0_outputs[4027];
    assign outputs[3241] = (layer0_outputs[3172]) ^ (layer0_outputs[7122]);
    assign outputs[3242] = ~(layer0_outputs[1375]);
    assign outputs[3243] = layer0_outputs[2833];
    assign outputs[3244] = layer0_outputs[4795];
    assign outputs[3245] = ~((layer0_outputs[5812]) & (layer0_outputs[6145]));
    assign outputs[3246] = (layer0_outputs[2909]) & (layer0_outputs[6520]);
    assign outputs[3247] = (layer0_outputs[5916]) & ~(layer0_outputs[4818]);
    assign outputs[3248] = layer0_outputs[5912];
    assign outputs[3249] = layer0_outputs[2318];
    assign outputs[3250] = (layer0_outputs[4082]) & ~(layer0_outputs[6216]);
    assign outputs[3251] = ~((layer0_outputs[4377]) ^ (layer0_outputs[7619]));
    assign outputs[3252] = layer0_outputs[1626];
    assign outputs[3253] = ~((layer0_outputs[4670]) | (layer0_outputs[4149]));
    assign outputs[3254] = (layer0_outputs[3150]) ^ (layer0_outputs[5365]);
    assign outputs[3255] = ~((layer0_outputs[6279]) ^ (layer0_outputs[5044]));
    assign outputs[3256] = layer0_outputs[4639];
    assign outputs[3257] = ~(layer0_outputs[4083]);
    assign outputs[3258] = layer0_outputs[6726];
    assign outputs[3259] = (layer0_outputs[3321]) ^ (layer0_outputs[7473]);
    assign outputs[3260] = (layer0_outputs[6734]) & ~(layer0_outputs[2202]);
    assign outputs[3261] = layer0_outputs[388];
    assign outputs[3262] = layer0_outputs[6408];
    assign outputs[3263] = ~((layer0_outputs[1812]) ^ (layer0_outputs[99]));
    assign outputs[3264] = (layer0_outputs[2016]) & ~(layer0_outputs[5834]);
    assign outputs[3265] = ~(layer0_outputs[7250]) | (layer0_outputs[6305]);
    assign outputs[3266] = (layer0_outputs[480]) & ~(layer0_outputs[4114]);
    assign outputs[3267] = (layer0_outputs[7535]) & ~(layer0_outputs[1011]);
    assign outputs[3268] = ~((layer0_outputs[3421]) ^ (layer0_outputs[1342]));
    assign outputs[3269] = ~((layer0_outputs[3896]) ^ (layer0_outputs[226]));
    assign outputs[3270] = (layer0_outputs[6010]) & ~(layer0_outputs[427]);
    assign outputs[3271] = (layer0_outputs[99]) & (layer0_outputs[5483]);
    assign outputs[3272] = (layer0_outputs[1755]) & (layer0_outputs[6213]);
    assign outputs[3273] = (layer0_outputs[919]) ^ (layer0_outputs[2882]);
    assign outputs[3274] = layer0_outputs[7436];
    assign outputs[3275] = (layer0_outputs[4155]) & (layer0_outputs[1005]);
    assign outputs[3276] = ~(layer0_outputs[666]);
    assign outputs[3277] = (layer0_outputs[6295]) ^ (layer0_outputs[193]);
    assign outputs[3278] = (layer0_outputs[1095]) & ~(layer0_outputs[5341]);
    assign outputs[3279] = ~(layer0_outputs[4348]);
    assign outputs[3280] = (layer0_outputs[1037]) ^ (layer0_outputs[2205]);
    assign outputs[3281] = ~((layer0_outputs[3585]) | (layer0_outputs[555]));
    assign outputs[3282] = (layer0_outputs[5498]) & ~(layer0_outputs[6423]);
    assign outputs[3283] = ~((layer0_outputs[6472]) ^ (layer0_outputs[6084]));
    assign outputs[3284] = ~((layer0_outputs[1300]) | (layer0_outputs[6552]));
    assign outputs[3285] = (layer0_outputs[720]) & ~(layer0_outputs[420]);
    assign outputs[3286] = (layer0_outputs[4812]) ^ (layer0_outputs[2790]);
    assign outputs[3287] = ~(layer0_outputs[6257]) | (layer0_outputs[1768]);
    assign outputs[3288] = ~(layer0_outputs[3856]);
    assign outputs[3289] = layer0_outputs[5296];
    assign outputs[3290] = (layer0_outputs[436]) ^ (layer0_outputs[5657]);
    assign outputs[3291] = ~(layer0_outputs[1851]);
    assign outputs[3292] = layer0_outputs[7579];
    assign outputs[3293] = (layer0_outputs[2770]) ^ (layer0_outputs[2347]);
    assign outputs[3294] = (layer0_outputs[6351]) ^ (layer0_outputs[1590]);
    assign outputs[3295] = layer0_outputs[4014];
    assign outputs[3296] = ~((layer0_outputs[5824]) ^ (layer0_outputs[3636]));
    assign outputs[3297] = ~(layer0_outputs[7005]);
    assign outputs[3298] = ~(layer0_outputs[1645]);
    assign outputs[3299] = (layer0_outputs[5345]) & ~(layer0_outputs[2878]);
    assign outputs[3300] = layer0_outputs[7343];
    assign outputs[3301] = (layer0_outputs[7339]) & ~(layer0_outputs[939]);
    assign outputs[3302] = layer0_outputs[2216];
    assign outputs[3303] = ~(layer0_outputs[7492]);
    assign outputs[3304] = ~((layer0_outputs[4134]) & (layer0_outputs[3381]));
    assign outputs[3305] = (layer0_outputs[6821]) ^ (layer0_outputs[1210]);
    assign outputs[3306] = ~(layer0_outputs[4822]);
    assign outputs[3307] = 1'b0;
    assign outputs[3308] = (layer0_outputs[5764]) & (layer0_outputs[4033]);
    assign outputs[3309] = (layer0_outputs[5385]) & (layer0_outputs[1172]);
    assign outputs[3310] = ~((layer0_outputs[4260]) | (layer0_outputs[4785]));
    assign outputs[3311] = layer0_outputs[4168];
    assign outputs[3312] = ~(layer0_outputs[817]);
    assign outputs[3313] = ~(layer0_outputs[7223]);
    assign outputs[3314] = ~(layer0_outputs[2055]);
    assign outputs[3315] = layer0_outputs[5878];
    assign outputs[3316] = 1'b0;
    assign outputs[3317] = ~(layer0_outputs[6115]);
    assign outputs[3318] = layer0_outputs[930];
    assign outputs[3319] = ~(layer0_outputs[1884]);
    assign outputs[3320] = (layer0_outputs[4432]) & ~(layer0_outputs[4026]);
    assign outputs[3321] = ~((layer0_outputs[798]) ^ (layer0_outputs[7118]));
    assign outputs[3322] = ~((layer0_outputs[4136]) | (layer0_outputs[261]));
    assign outputs[3323] = (layer0_outputs[4634]) & ~(layer0_outputs[602]);
    assign outputs[3324] = layer0_outputs[1769];
    assign outputs[3325] = ~((layer0_outputs[3153]) | (layer0_outputs[2837]));
    assign outputs[3326] = (layer0_outputs[2399]) ^ (layer0_outputs[3373]);
    assign outputs[3327] = ~((layer0_outputs[1702]) ^ (layer0_outputs[6498]));
    assign outputs[3328] = 1'b0;
    assign outputs[3329] = ~((layer0_outputs[448]) ^ (layer0_outputs[6742]));
    assign outputs[3330] = ~(layer0_outputs[1568]);
    assign outputs[3331] = ~((layer0_outputs[2806]) & (layer0_outputs[5388]));
    assign outputs[3332] = layer0_outputs[3549];
    assign outputs[3333] = layer0_outputs[2619];
    assign outputs[3334] = layer0_outputs[3133];
    assign outputs[3335] = (layer0_outputs[3405]) & ~(layer0_outputs[1814]);
    assign outputs[3336] = ~(layer0_outputs[4134]);
    assign outputs[3337] = ~((layer0_outputs[5968]) ^ (layer0_outputs[2603]));
    assign outputs[3338] = layer0_outputs[4758];
    assign outputs[3339] = ~(layer0_outputs[3660]) | (layer0_outputs[1058]);
    assign outputs[3340] = ~(layer0_outputs[5990]);
    assign outputs[3341] = (layer0_outputs[2245]) & (layer0_outputs[4043]);
    assign outputs[3342] = layer0_outputs[3444];
    assign outputs[3343] = (layer0_outputs[2289]) & (layer0_outputs[4490]);
    assign outputs[3344] = layer0_outputs[1984];
    assign outputs[3345] = layer0_outputs[6634];
    assign outputs[3346] = (layer0_outputs[1519]) ^ (layer0_outputs[3713]);
    assign outputs[3347] = layer0_outputs[529];
    assign outputs[3348] = ~((layer0_outputs[797]) ^ (layer0_outputs[5667]));
    assign outputs[3349] = ~((layer0_outputs[3876]) | (layer0_outputs[2609]));
    assign outputs[3350] = (layer0_outputs[921]) & ~(layer0_outputs[2291]);
    assign outputs[3351] = layer0_outputs[2391];
    assign outputs[3352] = (layer0_outputs[6011]) & (layer0_outputs[5634]);
    assign outputs[3353] = ~((layer0_outputs[3973]) | (layer0_outputs[1515]));
    assign outputs[3354] = layer0_outputs[4914];
    assign outputs[3355] = ~(layer0_outputs[5082]);
    assign outputs[3356] = (layer0_outputs[2317]) ^ (layer0_outputs[1931]);
    assign outputs[3357] = ~((layer0_outputs[6276]) ^ (layer0_outputs[3618]));
    assign outputs[3358] = layer0_outputs[7679];
    assign outputs[3359] = (layer0_outputs[3973]) ^ (layer0_outputs[6770]);
    assign outputs[3360] = (layer0_outputs[1212]) ^ (layer0_outputs[4542]);
    assign outputs[3361] = (layer0_outputs[3052]) & ~(layer0_outputs[7538]);
    assign outputs[3362] = layer0_outputs[5675];
    assign outputs[3363] = (layer0_outputs[6336]) & (layer0_outputs[335]);
    assign outputs[3364] = ~(layer0_outputs[2975]);
    assign outputs[3365] = (layer0_outputs[4539]) & ~(layer0_outputs[1196]);
    assign outputs[3366] = 1'b1;
    assign outputs[3367] = layer0_outputs[367];
    assign outputs[3368] = (layer0_outputs[1399]) ^ (layer0_outputs[6278]);
    assign outputs[3369] = ~((layer0_outputs[3544]) ^ (layer0_outputs[4031]));
    assign outputs[3370] = ~((layer0_outputs[6349]) | (layer0_outputs[5813]));
    assign outputs[3371] = ~(layer0_outputs[2971]);
    assign outputs[3372] = (layer0_outputs[4651]) & (layer0_outputs[2957]);
    assign outputs[3373] = (layer0_outputs[3146]) ^ (layer0_outputs[1338]);
    assign outputs[3374] = ~((layer0_outputs[3579]) ^ (layer0_outputs[1379]));
    assign outputs[3375] = (layer0_outputs[4723]) & ~(layer0_outputs[6582]);
    assign outputs[3376] = (layer0_outputs[4332]) & ~(layer0_outputs[2298]);
    assign outputs[3377] = (layer0_outputs[3901]) ^ (layer0_outputs[5097]);
    assign outputs[3378] = ~(layer0_outputs[3200]) | (layer0_outputs[2360]);
    assign outputs[3379] = (layer0_outputs[4290]) ^ (layer0_outputs[1585]);
    assign outputs[3380] = ~(layer0_outputs[3229]);
    assign outputs[3381] = (layer0_outputs[1057]) & (layer0_outputs[6919]);
    assign outputs[3382] = ~((layer0_outputs[3128]) & (layer0_outputs[4455]));
    assign outputs[3383] = ~((layer0_outputs[5615]) | (layer0_outputs[6747]));
    assign outputs[3384] = (layer0_outputs[4856]) & ~(layer0_outputs[620]);
    assign outputs[3385] = ~((layer0_outputs[7202]) ^ (layer0_outputs[1297]));
    assign outputs[3386] = layer0_outputs[6574];
    assign outputs[3387] = layer0_outputs[4856];
    assign outputs[3388] = ~(layer0_outputs[6716]);
    assign outputs[3389] = ~(layer0_outputs[7606]);
    assign outputs[3390] = layer0_outputs[567];
    assign outputs[3391] = ~(layer0_outputs[7106]);
    assign outputs[3392] = ~(layer0_outputs[1616]);
    assign outputs[3393] = ~(layer0_outputs[4104]);
    assign outputs[3394] = ~(layer0_outputs[4804]);
    assign outputs[3395] = ~(layer0_outputs[3497]) | (layer0_outputs[1231]);
    assign outputs[3396] = (layer0_outputs[2504]) ^ (layer0_outputs[4305]);
    assign outputs[3397] = (layer0_outputs[7263]) & (layer0_outputs[6680]);
    assign outputs[3398] = (layer0_outputs[3845]) & ~(layer0_outputs[5004]);
    assign outputs[3399] = ~(layer0_outputs[1574]) | (layer0_outputs[6736]);
    assign outputs[3400] = (layer0_outputs[2030]) ^ (layer0_outputs[2330]);
    assign outputs[3401] = (layer0_outputs[5038]) ^ (layer0_outputs[6224]);
    assign outputs[3402] = ~((layer0_outputs[4787]) | (layer0_outputs[6993]));
    assign outputs[3403] = ~(layer0_outputs[5387]) | (layer0_outputs[2076]);
    assign outputs[3404] = layer0_outputs[2695];
    assign outputs[3405] = ~((layer0_outputs[3632]) ^ (layer0_outputs[617]));
    assign outputs[3406] = ~(layer0_outputs[2624]) | (layer0_outputs[3477]);
    assign outputs[3407] = layer0_outputs[6751];
    assign outputs[3408] = (layer0_outputs[7258]) ^ (layer0_outputs[5461]);
    assign outputs[3409] = ~((layer0_outputs[434]) | (layer0_outputs[68]));
    assign outputs[3410] = 1'b0;
    assign outputs[3411] = layer0_outputs[6784];
    assign outputs[3412] = (layer0_outputs[3379]) ^ (layer0_outputs[1362]);
    assign outputs[3413] = (layer0_outputs[1874]) | (layer0_outputs[7524]);
    assign outputs[3414] = (layer0_outputs[2592]) ^ (layer0_outputs[2089]);
    assign outputs[3415] = layer0_outputs[6014];
    assign outputs[3416] = 1'b0;
    assign outputs[3417] = ~((layer0_outputs[6258]) | (layer0_outputs[4541]));
    assign outputs[3418] = (layer0_outputs[344]) & ~(layer0_outputs[5248]);
    assign outputs[3419] = ~(layer0_outputs[5468]) | (layer0_outputs[690]);
    assign outputs[3420] = (layer0_outputs[3464]) & ~(layer0_outputs[6343]);
    assign outputs[3421] = ~((layer0_outputs[1875]) | (layer0_outputs[6650]));
    assign outputs[3422] = ~((layer0_outputs[594]) ^ (layer0_outputs[3012]));
    assign outputs[3423] = ~((layer0_outputs[5046]) | (layer0_outputs[1513]));
    assign outputs[3424] = (layer0_outputs[348]) & ~(layer0_outputs[7311]);
    assign outputs[3425] = ~(layer0_outputs[2294]);
    assign outputs[3426] = layer0_outputs[2972];
    assign outputs[3427] = ~(layer0_outputs[2438]);
    assign outputs[3428] = (layer0_outputs[4197]) ^ (layer0_outputs[2395]);
    assign outputs[3429] = ~(layer0_outputs[106]) | (layer0_outputs[1872]);
    assign outputs[3430] = ~(layer0_outputs[6981]);
    assign outputs[3431] = ~(layer0_outputs[6127]) | (layer0_outputs[5263]);
    assign outputs[3432] = layer0_outputs[7339];
    assign outputs[3433] = ~(layer0_outputs[1891]);
    assign outputs[3434] = ~((layer0_outputs[5454]) ^ (layer0_outputs[5187]));
    assign outputs[3435] = ~((layer0_outputs[3083]) ^ (layer0_outputs[2084]));
    assign outputs[3436] = (layer0_outputs[3558]) ^ (layer0_outputs[7417]);
    assign outputs[3437] = ~(layer0_outputs[2010]);
    assign outputs[3438] = ~(layer0_outputs[5478]);
    assign outputs[3439] = ~((layer0_outputs[1609]) | (layer0_outputs[3081]));
    assign outputs[3440] = (layer0_outputs[5887]) ^ (layer0_outputs[7481]);
    assign outputs[3441] = ~((layer0_outputs[3146]) | (layer0_outputs[4212]));
    assign outputs[3442] = ~((layer0_outputs[6536]) ^ (layer0_outputs[4119]));
    assign outputs[3443] = (layer0_outputs[1709]) ^ (layer0_outputs[3715]);
    assign outputs[3444] = (layer0_outputs[6528]) & ~(layer0_outputs[2879]);
    assign outputs[3445] = ~(layer0_outputs[5434]);
    assign outputs[3446] = layer0_outputs[6593];
    assign outputs[3447] = layer0_outputs[4696];
    assign outputs[3448] = (layer0_outputs[903]) & ~(layer0_outputs[5644]);
    assign outputs[3449] = layer0_outputs[2135];
    assign outputs[3450] = (layer0_outputs[665]) & (layer0_outputs[93]);
    assign outputs[3451] = (layer0_outputs[2004]) & (layer0_outputs[1831]);
    assign outputs[3452] = ~((layer0_outputs[859]) | (layer0_outputs[1664]));
    assign outputs[3453] = (layer0_outputs[6518]) & ~(layer0_outputs[80]);
    assign outputs[3454] = layer0_outputs[6524];
    assign outputs[3455] = layer0_outputs[2629];
    assign outputs[3456] = ~(layer0_outputs[2116]);
    assign outputs[3457] = (layer0_outputs[3524]) & ~(layer0_outputs[5774]);
    assign outputs[3458] = ~(layer0_outputs[4112]);
    assign outputs[3459] = layer0_outputs[1611];
    assign outputs[3460] = ~(layer0_outputs[4748]);
    assign outputs[3461] = (layer0_outputs[3823]) | (layer0_outputs[637]);
    assign outputs[3462] = (layer0_outputs[7206]) ^ (layer0_outputs[6333]);
    assign outputs[3463] = (layer0_outputs[6526]) | (layer0_outputs[1655]);
    assign outputs[3464] = ~(layer0_outputs[4254]);
    assign outputs[3465] = (layer0_outputs[3161]) ^ (layer0_outputs[3376]);
    assign outputs[3466] = (layer0_outputs[1902]) & (layer0_outputs[629]);
    assign outputs[3467] = (layer0_outputs[1251]) ^ (layer0_outputs[2222]);
    assign outputs[3468] = ~((layer0_outputs[6690]) ^ (layer0_outputs[1937]));
    assign outputs[3469] = (layer0_outputs[234]) ^ (layer0_outputs[979]);
    assign outputs[3470] = ~(layer0_outputs[1689]);
    assign outputs[3471] = ~((layer0_outputs[2481]) ^ (layer0_outputs[3571]));
    assign outputs[3472] = layer0_outputs[3400];
    assign outputs[3473] = ~((layer0_outputs[583]) ^ (layer0_outputs[5470]));
    assign outputs[3474] = ~(layer0_outputs[3104]);
    assign outputs[3475] = (layer0_outputs[1155]) & (layer0_outputs[6200]);
    assign outputs[3476] = (layer0_outputs[6906]) ^ (layer0_outputs[525]);
    assign outputs[3477] = ~(layer0_outputs[5589]);
    assign outputs[3478] = (layer0_outputs[647]) ^ (layer0_outputs[6671]);
    assign outputs[3479] = (layer0_outputs[6923]) & ~(layer0_outputs[1712]);
    assign outputs[3480] = ~((layer0_outputs[2060]) | (layer0_outputs[1257]));
    assign outputs[3481] = ~(layer0_outputs[6268]);
    assign outputs[3482] = ~((layer0_outputs[4074]) | (layer0_outputs[2477]));
    assign outputs[3483] = (layer0_outputs[4253]) & ~(layer0_outputs[7302]);
    assign outputs[3484] = ~((layer0_outputs[1164]) ^ (layer0_outputs[6537]));
    assign outputs[3485] = (layer0_outputs[4235]) ^ (layer0_outputs[6081]);
    assign outputs[3486] = (layer0_outputs[7532]) & ~(layer0_outputs[4433]);
    assign outputs[3487] = ~(layer0_outputs[2681]);
    assign outputs[3488] = layer0_outputs[1766];
    assign outputs[3489] = (layer0_outputs[5353]) & (layer0_outputs[4800]);
    assign outputs[3490] = (layer0_outputs[1359]) ^ (layer0_outputs[4080]);
    assign outputs[3491] = ~((layer0_outputs[7083]) | (layer0_outputs[6572]));
    assign outputs[3492] = layer0_outputs[6166];
    assign outputs[3493] = ~((layer0_outputs[7556]) | (layer0_outputs[3770]));
    assign outputs[3494] = ~(layer0_outputs[5074]);
    assign outputs[3495] = layer0_outputs[3201];
    assign outputs[3496] = ~(layer0_outputs[4440]) | (layer0_outputs[2857]);
    assign outputs[3497] = ~((layer0_outputs[4452]) | (layer0_outputs[1967]));
    assign outputs[3498] = ~(layer0_outputs[440]);
    assign outputs[3499] = (layer0_outputs[6483]) & (layer0_outputs[560]);
    assign outputs[3500] = (layer0_outputs[1245]) ^ (layer0_outputs[3732]);
    assign outputs[3501] = (layer0_outputs[5402]) ^ (layer0_outputs[7006]);
    assign outputs[3502] = ~((layer0_outputs[4661]) | (layer0_outputs[2894]));
    assign outputs[3503] = ~(layer0_outputs[807]) | (layer0_outputs[1747]);
    assign outputs[3504] = ~((layer0_outputs[5263]) | (layer0_outputs[1588]));
    assign outputs[3505] = layer0_outputs[2257];
    assign outputs[3506] = ~(layer0_outputs[5023]);
    assign outputs[3507] = ~((layer0_outputs[3571]) ^ (layer0_outputs[444]));
    assign outputs[3508] = layer0_outputs[5761];
    assign outputs[3509] = (layer0_outputs[5865]) & ~(layer0_outputs[1508]);
    assign outputs[3510] = ~(layer0_outputs[5732]);
    assign outputs[3511] = ~(layer0_outputs[83]);
    assign outputs[3512] = ~((layer0_outputs[4609]) ^ (layer0_outputs[2607]));
    assign outputs[3513] = layer0_outputs[304];
    assign outputs[3514] = 1'b0;
    assign outputs[3515] = ~(layer0_outputs[2121]);
    assign outputs[3516] = layer0_outputs[174];
    assign outputs[3517] = ~(layer0_outputs[1809]);
    assign outputs[3518] = layer0_outputs[769];
    assign outputs[3519] = (layer0_outputs[5533]) ^ (layer0_outputs[2081]);
    assign outputs[3520] = layer0_outputs[4719];
    assign outputs[3521] = ~((layer0_outputs[2119]) ^ (layer0_outputs[4461]));
    assign outputs[3522] = ~(layer0_outputs[5597]);
    assign outputs[3523] = (layer0_outputs[2658]) & ~(layer0_outputs[416]);
    assign outputs[3524] = ~(layer0_outputs[4637]);
    assign outputs[3525] = (layer0_outputs[6334]) & ~(layer0_outputs[3103]);
    assign outputs[3526] = ~(layer0_outputs[2030]) | (layer0_outputs[622]);
    assign outputs[3527] = ~(layer0_outputs[2463]);
    assign outputs[3528] = layer0_outputs[1553];
    assign outputs[3529] = ~(layer0_outputs[29]);
    assign outputs[3530] = (layer0_outputs[1240]) & ~(layer0_outputs[7678]);
    assign outputs[3531] = ~(layer0_outputs[5921]);
    assign outputs[3532] = layer0_outputs[4041];
    assign outputs[3533] = (layer0_outputs[2455]) & (layer0_outputs[892]);
    assign outputs[3534] = ~(layer0_outputs[146]);
    assign outputs[3535] = ~(layer0_outputs[2845]) | (layer0_outputs[2136]);
    assign outputs[3536] = (layer0_outputs[2904]) ^ (layer0_outputs[7458]);
    assign outputs[3537] = (layer0_outputs[721]) & ~(layer0_outputs[2090]);
    assign outputs[3538] = ~(layer0_outputs[3611]);
    assign outputs[3539] = ~((layer0_outputs[2847]) ^ (layer0_outputs[6898]));
    assign outputs[3540] = layer0_outputs[4539];
    assign outputs[3541] = ~(layer0_outputs[1701]);
    assign outputs[3542] = ~(layer0_outputs[5187]);
    assign outputs[3543] = layer0_outputs[6905];
    assign outputs[3544] = (layer0_outputs[5389]) & ~(layer0_outputs[6397]);
    assign outputs[3545] = ~((layer0_outputs[5082]) & (layer0_outputs[2281]));
    assign outputs[3546] = ~(layer0_outputs[41]);
    assign outputs[3547] = ~(layer0_outputs[7543]);
    assign outputs[3548] = (layer0_outputs[2969]) ^ (layer0_outputs[1019]);
    assign outputs[3549] = (layer0_outputs[4131]) & ~(layer0_outputs[7430]);
    assign outputs[3550] = layer0_outputs[3037];
    assign outputs[3551] = ~(layer0_outputs[5396]);
    assign outputs[3552] = (layer0_outputs[5620]) & (layer0_outputs[6770]);
    assign outputs[3553] = (layer0_outputs[5165]) | (layer0_outputs[1418]);
    assign outputs[3554] = ~(layer0_outputs[3743]);
    assign outputs[3555] = layer0_outputs[6079];
    assign outputs[3556] = ~(layer0_outputs[5537]);
    assign outputs[3557] = ~((layer0_outputs[4090]) & (layer0_outputs[2292]));
    assign outputs[3558] = ~(layer0_outputs[5288]);
    assign outputs[3559] = ~((layer0_outputs[2420]) ^ (layer0_outputs[2219]));
    assign outputs[3560] = (layer0_outputs[2727]) ^ (layer0_outputs[6456]);
    assign outputs[3561] = ~(layer0_outputs[3829]);
    assign outputs[3562] = ~((layer0_outputs[3580]) ^ (layer0_outputs[1430]));
    assign outputs[3563] = (layer0_outputs[6106]) & ~(layer0_outputs[3761]);
    assign outputs[3564] = (layer0_outputs[4182]) & ~(layer0_outputs[6845]);
    assign outputs[3565] = ~((layer0_outputs[2399]) ^ (layer0_outputs[6608]));
    assign outputs[3566] = ~(layer0_outputs[390]);
    assign outputs[3567] = layer0_outputs[6027];
    assign outputs[3568] = ~((layer0_outputs[7408]) | (layer0_outputs[3269]));
    assign outputs[3569] = (layer0_outputs[6571]) ^ (layer0_outputs[3086]);
    assign outputs[3570] = (layer0_outputs[163]) ^ (layer0_outputs[7427]);
    assign outputs[3571] = (layer0_outputs[3834]) & (layer0_outputs[7589]);
    assign outputs[3572] = ~(layer0_outputs[7269]);
    assign outputs[3573] = layer0_outputs[1356];
    assign outputs[3574] = layer0_outputs[7259];
    assign outputs[3575] = (layer0_outputs[6885]) ^ (layer0_outputs[7426]);
    assign outputs[3576] = ~((layer0_outputs[3354]) | (layer0_outputs[7546]));
    assign outputs[3577] = ~(layer0_outputs[4407]) | (layer0_outputs[7392]);
    assign outputs[3578] = ~(layer0_outputs[197]);
    assign outputs[3579] = (layer0_outputs[5463]) & (layer0_outputs[5801]);
    assign outputs[3580] = (layer0_outputs[5931]) ^ (layer0_outputs[3591]);
    assign outputs[3581] = (layer0_outputs[4713]) & ~(layer0_outputs[7364]);
    assign outputs[3582] = (layer0_outputs[5869]) & ~(layer0_outputs[2036]);
    assign outputs[3583] = ~((layer0_outputs[2181]) | (layer0_outputs[5249]));
    assign outputs[3584] = ~(layer0_outputs[5819]);
    assign outputs[3585] = 1'b0;
    assign outputs[3586] = ~((layer0_outputs[7209]) | (layer0_outputs[5702]));
    assign outputs[3587] = ~(layer0_outputs[2408]);
    assign outputs[3588] = ~(layer0_outputs[2370]) | (layer0_outputs[3885]);
    assign outputs[3589] = (layer0_outputs[3966]) ^ (layer0_outputs[3637]);
    assign outputs[3590] = ~(layer0_outputs[5046]);
    assign outputs[3591] = (layer0_outputs[1770]) & (layer0_outputs[363]);
    assign outputs[3592] = layer0_outputs[2585];
    assign outputs[3593] = ~(layer0_outputs[3741]);
    assign outputs[3594] = ~(layer0_outputs[7595]);
    assign outputs[3595] = (layer0_outputs[4846]) & ~(layer0_outputs[2058]);
    assign outputs[3596] = ~(layer0_outputs[5151]);
    assign outputs[3597] = (layer0_outputs[3492]) | (layer0_outputs[4714]);
    assign outputs[3598] = (layer0_outputs[4593]) & (layer0_outputs[7001]);
    assign outputs[3599] = layer0_outputs[3616];
    assign outputs[3600] = (layer0_outputs[5655]) ^ (layer0_outputs[1003]);
    assign outputs[3601] = ~((layer0_outputs[2572]) ^ (layer0_outputs[3556]));
    assign outputs[3602] = layer0_outputs[1896];
    assign outputs[3603] = ~(layer0_outputs[5578]);
    assign outputs[3604] = ~(layer0_outputs[6270]);
    assign outputs[3605] = (layer0_outputs[16]) & ~(layer0_outputs[316]);
    assign outputs[3606] = ~(layer0_outputs[5736]);
    assign outputs[3607] = (layer0_outputs[5298]) | (layer0_outputs[494]);
    assign outputs[3608] = ~((layer0_outputs[4302]) | (layer0_outputs[7671]));
    assign outputs[3609] = (layer0_outputs[4858]) & ~(layer0_outputs[5110]);
    assign outputs[3610] = ~(layer0_outputs[5676]);
    assign outputs[3611] = (layer0_outputs[4578]) & ~(layer0_outputs[556]);
    assign outputs[3612] = ~((layer0_outputs[7418]) ^ (layer0_outputs[5000]));
    assign outputs[3613] = ~((layer0_outputs[3379]) ^ (layer0_outputs[7164]));
    assign outputs[3614] = ~((layer0_outputs[5691]) ^ (layer0_outputs[5630]));
    assign outputs[3615] = layer0_outputs[1399];
    assign outputs[3616] = ~(layer0_outputs[3214]);
    assign outputs[3617] = layer0_outputs[6841];
    assign outputs[3618] = ~(layer0_outputs[2240]);
    assign outputs[3619] = ~(layer0_outputs[7504]) | (layer0_outputs[3832]);
    assign outputs[3620] = ~((layer0_outputs[3688]) ^ (layer0_outputs[1376]));
    assign outputs[3621] = ~(layer0_outputs[6581]) | (layer0_outputs[3650]);
    assign outputs[3622] = (layer0_outputs[5896]) & (layer0_outputs[1267]);
    assign outputs[3623] = ~(layer0_outputs[5313]);
    assign outputs[3624] = layer0_outputs[4197];
    assign outputs[3625] = (layer0_outputs[3031]) & ~(layer0_outputs[881]);
    assign outputs[3626] = ~(layer0_outputs[5246]);
    assign outputs[3627] = layer0_outputs[5051];
    assign outputs[3628] = (layer0_outputs[914]) | (layer0_outputs[5326]);
    assign outputs[3629] = (layer0_outputs[750]) ^ (layer0_outputs[6942]);
    assign outputs[3630] = layer0_outputs[3033];
    assign outputs[3631] = (layer0_outputs[1736]) & (layer0_outputs[1447]);
    assign outputs[3632] = ~((layer0_outputs[45]) & (layer0_outputs[153]));
    assign outputs[3633] = layer0_outputs[5888];
    assign outputs[3634] = ~(layer0_outputs[1351]);
    assign outputs[3635] = layer0_outputs[2133];
    assign outputs[3636] = ~((layer0_outputs[4628]) ^ (layer0_outputs[1235]));
    assign outputs[3637] = ~(layer0_outputs[219]);
    assign outputs[3638] = (layer0_outputs[6908]) & ~(layer0_outputs[6603]);
    assign outputs[3639] = ~(layer0_outputs[7485]);
    assign outputs[3640] = (layer0_outputs[238]) ^ (layer0_outputs[4685]);
    assign outputs[3641] = ~((layer0_outputs[7213]) ^ (layer0_outputs[514]));
    assign outputs[3642] = ~(layer0_outputs[3438]);
    assign outputs[3643] = ~((layer0_outputs[4753]) ^ (layer0_outputs[4937]));
    assign outputs[3644] = ~(layer0_outputs[185]);
    assign outputs[3645] = (layer0_outputs[741]) & ~(layer0_outputs[352]);
    assign outputs[3646] = ~(layer0_outputs[5492]);
    assign outputs[3647] = (layer0_outputs[4002]) & (layer0_outputs[4632]);
    assign outputs[3648] = ~(layer0_outputs[1616]);
    assign outputs[3649] = (layer0_outputs[1707]) ^ (layer0_outputs[7627]);
    assign outputs[3650] = ~(layer0_outputs[6824]);
    assign outputs[3651] = ~((layer0_outputs[1482]) & (layer0_outputs[4246]));
    assign outputs[3652] = (layer0_outputs[2792]) & ~(layer0_outputs[3465]);
    assign outputs[3653] = ~((layer0_outputs[7511]) ^ (layer0_outputs[5022]));
    assign outputs[3654] = layer0_outputs[5049];
    assign outputs[3655] = ~(layer0_outputs[5646]);
    assign outputs[3656] = (layer0_outputs[377]) & (layer0_outputs[377]);
    assign outputs[3657] = ~((layer0_outputs[72]) ^ (layer0_outputs[7101]));
    assign outputs[3658] = (layer0_outputs[2850]) & ~(layer0_outputs[3046]);
    assign outputs[3659] = ~((layer0_outputs[2866]) ^ (layer0_outputs[5973]));
    assign outputs[3660] = (layer0_outputs[3206]) & ~(layer0_outputs[4154]);
    assign outputs[3661] = ~(layer0_outputs[4872]);
    assign outputs[3662] = (layer0_outputs[1125]) & ~(layer0_outputs[3114]);
    assign outputs[3663] = (layer0_outputs[727]) & (layer0_outputs[5232]);
    assign outputs[3664] = ~((layer0_outputs[2741]) ^ (layer0_outputs[6111]));
    assign outputs[3665] = ~((layer0_outputs[3351]) ^ (layer0_outputs[4537]));
    assign outputs[3666] = ~(layer0_outputs[1222]);
    assign outputs[3667] = layer0_outputs[5714];
    assign outputs[3668] = (layer0_outputs[3202]) ^ (layer0_outputs[7008]);
    assign outputs[3669] = (layer0_outputs[6679]) & ~(layer0_outputs[6113]);
    assign outputs[3670] = (layer0_outputs[693]) & (layer0_outputs[3159]);
    assign outputs[3671] = (layer0_outputs[4651]) & ~(layer0_outputs[1823]);
    assign outputs[3672] = ~((layer0_outputs[222]) ^ (layer0_outputs[4783]));
    assign outputs[3673] = (layer0_outputs[6156]) & ~(layer0_outputs[3137]);
    assign outputs[3674] = layer0_outputs[5754];
    assign outputs[3675] = layer0_outputs[228];
    assign outputs[3676] = ~((layer0_outputs[2605]) ^ (layer0_outputs[2491]));
    assign outputs[3677] = ~(layer0_outputs[4190]);
    assign outputs[3678] = ~(layer0_outputs[6546]);
    assign outputs[3679] = (layer0_outputs[4030]) & ~(layer0_outputs[655]);
    assign outputs[3680] = ~(layer0_outputs[3810]);
    assign outputs[3681] = layer0_outputs[3181];
    assign outputs[3682] = layer0_outputs[3563];
    assign outputs[3683] = ~((layer0_outputs[4732]) ^ (layer0_outputs[888]));
    assign outputs[3684] = layer0_outputs[1620];
    assign outputs[3685] = (layer0_outputs[767]) & ~(layer0_outputs[7004]);
    assign outputs[3686] = layer0_outputs[6089];
    assign outputs[3687] = ~(layer0_outputs[7546]);
    assign outputs[3688] = layer0_outputs[2321];
    assign outputs[3689] = ~(layer0_outputs[1346]);
    assign outputs[3690] = (layer0_outputs[6026]) & ~(layer0_outputs[2836]);
    assign outputs[3691] = ~(layer0_outputs[6561]);
    assign outputs[3692] = ~((layer0_outputs[7402]) ^ (layer0_outputs[1337]));
    assign outputs[3693] = layer0_outputs[5386];
    assign outputs[3694] = (layer0_outputs[87]) & ~(layer0_outputs[5191]);
    assign outputs[3695] = ~((layer0_outputs[3008]) ^ (layer0_outputs[707]));
    assign outputs[3696] = ~((layer0_outputs[1064]) | (layer0_outputs[5705]));
    assign outputs[3697] = layer0_outputs[3367];
    assign outputs[3698] = ~(layer0_outputs[1605]);
    assign outputs[3699] = ~(layer0_outputs[4214]);
    assign outputs[3700] = ~((layer0_outputs[1934]) ^ (layer0_outputs[2470]));
    assign outputs[3701] = ~(layer0_outputs[2981]);
    assign outputs[3702] = ~((layer0_outputs[6341]) ^ (layer0_outputs[3403]));
    assign outputs[3703] = layer0_outputs[5734];
    assign outputs[3704] = (layer0_outputs[4786]) & ~(layer0_outputs[6449]);
    assign outputs[3705] = (layer0_outputs[603]) & ~(layer0_outputs[6421]);
    assign outputs[3706] = (layer0_outputs[5805]) & ~(layer0_outputs[5473]);
    assign outputs[3707] = ~(layer0_outputs[6800]) | (layer0_outputs[6139]);
    assign outputs[3708] = ~(layer0_outputs[1685]);
    assign outputs[3709] = (layer0_outputs[6012]) ^ (layer0_outputs[6650]);
    assign outputs[3710] = layer0_outputs[263];
    assign outputs[3711] = ~(layer0_outputs[5368]);
    assign outputs[3712] = ~((layer0_outputs[5555]) ^ (layer0_outputs[6824]));
    assign outputs[3713] = ~(layer0_outputs[3354]);
    assign outputs[3714] = ~(layer0_outputs[3943]);
    assign outputs[3715] = layer0_outputs[7651];
    assign outputs[3716] = (layer0_outputs[2528]) & ~(layer0_outputs[6693]);
    assign outputs[3717] = layer0_outputs[3993];
    assign outputs[3718] = (layer0_outputs[7552]) & ~(layer0_outputs[901]);
    assign outputs[3719] = layer0_outputs[6917];
    assign outputs[3720] = (layer0_outputs[1700]) ^ (layer0_outputs[3552]);
    assign outputs[3721] = ~((layer0_outputs[4963]) ^ (layer0_outputs[2919]));
    assign outputs[3722] = ~(layer0_outputs[7031]);
    assign outputs[3723] = layer0_outputs[2430];
    assign outputs[3724] = ~((layer0_outputs[1695]) ^ (layer0_outputs[6454]));
    assign outputs[3725] = ~(layer0_outputs[3976]);
    assign outputs[3726] = layer0_outputs[3439];
    assign outputs[3727] = (layer0_outputs[1987]) ^ (layer0_outputs[4707]);
    assign outputs[3728] = (layer0_outputs[988]) ^ (layer0_outputs[1614]);
    assign outputs[3729] = (layer0_outputs[5741]) ^ (layer0_outputs[1930]);
    assign outputs[3730] = layer0_outputs[7265];
    assign outputs[3731] = (layer0_outputs[843]) & (layer0_outputs[2332]);
    assign outputs[3732] = ~(layer0_outputs[398]) | (layer0_outputs[2705]);
    assign outputs[3733] = (layer0_outputs[7146]) & (layer0_outputs[5325]);
    assign outputs[3734] = ~(layer0_outputs[292]);
    assign outputs[3735] = (layer0_outputs[6452]) ^ (layer0_outputs[441]);
    assign outputs[3736] = ~(layer0_outputs[1292]);
    assign outputs[3737] = ~((layer0_outputs[1978]) | (layer0_outputs[5545]));
    assign outputs[3738] = layer0_outputs[2135];
    assign outputs[3739] = ~((layer0_outputs[4172]) ^ (layer0_outputs[4682]));
    assign outputs[3740] = (layer0_outputs[6289]) & ~(layer0_outputs[4509]);
    assign outputs[3741] = layer0_outputs[3259];
    assign outputs[3742] = (layer0_outputs[5840]) ^ (layer0_outputs[6003]);
    assign outputs[3743] = (layer0_outputs[4971]) ^ (layer0_outputs[365]);
    assign outputs[3744] = ~(layer0_outputs[829]);
    assign outputs[3745] = ~(layer0_outputs[4701]) | (layer0_outputs[1811]);
    assign outputs[3746] = layer0_outputs[900];
    assign outputs[3747] = (layer0_outputs[490]) & ~(layer0_outputs[4822]);
    assign outputs[3748] = ~(layer0_outputs[6170]);
    assign outputs[3749] = ~((layer0_outputs[2943]) ^ (layer0_outputs[1777]));
    assign outputs[3750] = (layer0_outputs[6466]) ^ (layer0_outputs[448]);
    assign outputs[3751] = ~((layer0_outputs[1434]) ^ (layer0_outputs[5770]));
    assign outputs[3752] = (layer0_outputs[4960]) & ~(layer0_outputs[3335]);
    assign outputs[3753] = ~(layer0_outputs[7061]) | (layer0_outputs[3998]);
    assign outputs[3754] = ~((layer0_outputs[372]) | (layer0_outputs[7109]));
    assign outputs[3755] = ~(layer0_outputs[1694]);
    assign outputs[3756] = (layer0_outputs[3410]) ^ (layer0_outputs[1042]);
    assign outputs[3757] = layer0_outputs[5043];
    assign outputs[3758] = ~(layer0_outputs[2284]);
    assign outputs[3759] = (layer0_outputs[5859]) ^ (layer0_outputs[7034]);
    assign outputs[3760] = ~(layer0_outputs[1107]);
    assign outputs[3761] = (layer0_outputs[3731]) ^ (layer0_outputs[1901]);
    assign outputs[3762] = (layer0_outputs[7458]) & ~(layer0_outputs[3500]);
    assign outputs[3763] = layer0_outputs[4633];
    assign outputs[3764] = ~((layer0_outputs[6549]) | (layer0_outputs[4417]));
    assign outputs[3765] = layer0_outputs[1862];
    assign outputs[3766] = layer0_outputs[7498];
    assign outputs[3767] = layer0_outputs[5293];
    assign outputs[3768] = ~(layer0_outputs[6611]);
    assign outputs[3769] = layer0_outputs[6948];
    assign outputs[3770] = (layer0_outputs[6684]) ^ (layer0_outputs[1840]);
    assign outputs[3771] = layer0_outputs[3386];
    assign outputs[3772] = ~(layer0_outputs[2630]);
    assign outputs[3773] = (layer0_outputs[6355]) & ~(layer0_outputs[3338]);
    assign outputs[3774] = (layer0_outputs[6587]) ^ (layer0_outputs[5687]);
    assign outputs[3775] = layer0_outputs[4378];
    assign outputs[3776] = ~(layer0_outputs[6938]);
    assign outputs[3777] = (layer0_outputs[452]) | (layer0_outputs[5540]);
    assign outputs[3778] = ~(layer0_outputs[7417]);
    assign outputs[3779] = ~((layer0_outputs[3713]) ^ (layer0_outputs[2137]));
    assign outputs[3780] = ~((layer0_outputs[7565]) & (layer0_outputs[6474]));
    assign outputs[3781] = (layer0_outputs[5107]) & ~(layer0_outputs[7325]);
    assign outputs[3782] = (layer0_outputs[1251]) & (layer0_outputs[3165]);
    assign outputs[3783] = layer0_outputs[3950];
    assign outputs[3784] = ~((layer0_outputs[2828]) ^ (layer0_outputs[5962]));
    assign outputs[3785] = (layer0_outputs[3455]) | (layer0_outputs[4297]);
    assign outputs[3786] = ~(layer0_outputs[5478]);
    assign outputs[3787] = layer0_outputs[2911];
    assign outputs[3788] = layer0_outputs[4497];
    assign outputs[3789] = ~((layer0_outputs[4710]) | (layer0_outputs[3055]));
    assign outputs[3790] = (layer0_outputs[1264]) & ~(layer0_outputs[6854]);
    assign outputs[3791] = layer0_outputs[6124];
    assign outputs[3792] = (layer0_outputs[1658]) & ~(layer0_outputs[1216]);
    assign outputs[3793] = (layer0_outputs[1935]) & ~(layer0_outputs[762]);
    assign outputs[3794] = layer0_outputs[4252];
    assign outputs[3795] = ~((layer0_outputs[284]) | (layer0_outputs[4087]));
    assign outputs[3796] = (layer0_outputs[297]) ^ (layer0_outputs[3952]);
    assign outputs[3797] = layer0_outputs[6047];
    assign outputs[3798] = layer0_outputs[1117];
    assign outputs[3799] = layer0_outputs[4119];
    assign outputs[3800] = ~(layer0_outputs[7578]);
    assign outputs[3801] = (layer0_outputs[92]) ^ (layer0_outputs[2108]);
    assign outputs[3802] = ~(layer0_outputs[5110]);
    assign outputs[3803] = (layer0_outputs[1429]) & ~(layer0_outputs[2011]);
    assign outputs[3804] = ~(layer0_outputs[5547]);
    assign outputs[3805] = (layer0_outputs[2341]) & (layer0_outputs[325]);
    assign outputs[3806] = (layer0_outputs[3573]) & (layer0_outputs[4309]);
    assign outputs[3807] = layer0_outputs[5532];
    assign outputs[3808] = ~((layer0_outputs[407]) | (layer0_outputs[4566]));
    assign outputs[3809] = (layer0_outputs[2176]) & ~(layer0_outputs[1976]);
    assign outputs[3810] = (layer0_outputs[6524]) & (layer0_outputs[5860]);
    assign outputs[3811] = (layer0_outputs[1222]) ^ (layer0_outputs[4695]);
    assign outputs[3812] = (layer0_outputs[889]) & ~(layer0_outputs[7540]);
    assign outputs[3813] = ~((layer0_outputs[3712]) ^ (layer0_outputs[5759]));
    assign outputs[3814] = layer0_outputs[7062];
    assign outputs[3815] = layer0_outputs[475];
    assign outputs[3816] = layer0_outputs[7214];
    assign outputs[3817] = layer0_outputs[4389];
    assign outputs[3818] = ~(layer0_outputs[6700]);
    assign outputs[3819] = (layer0_outputs[4875]) ^ (layer0_outputs[5897]);
    assign outputs[3820] = (layer0_outputs[652]) & (layer0_outputs[787]);
    assign outputs[3821] = ~((layer0_outputs[1945]) ^ (layer0_outputs[2268]));
    assign outputs[3822] = layer0_outputs[4545];
    assign outputs[3823] = layer0_outputs[3395];
    assign outputs[3824] = ~((layer0_outputs[2398]) ^ (layer0_outputs[3739]));
    assign outputs[3825] = layer0_outputs[6950];
    assign outputs[3826] = layer0_outputs[7431];
    assign outputs[3827] = layer0_outputs[7194];
    assign outputs[3828] = layer0_outputs[544];
    assign outputs[3829] = ~((layer0_outputs[2591]) ^ (layer0_outputs[4266]));
    assign outputs[3830] = (layer0_outputs[6255]) & ~(layer0_outputs[6234]);
    assign outputs[3831] = ~(layer0_outputs[3040]);
    assign outputs[3832] = layer0_outputs[3127];
    assign outputs[3833] = layer0_outputs[5301];
    assign outputs[3834] = ~((layer0_outputs[1683]) ^ (layer0_outputs[7259]));
    assign outputs[3835] = (layer0_outputs[4839]) & (layer0_outputs[4359]);
    assign outputs[3836] = ~((layer0_outputs[158]) ^ (layer0_outputs[3808]));
    assign outputs[3837] = ~((layer0_outputs[1444]) ^ (layer0_outputs[6068]));
    assign outputs[3838] = (layer0_outputs[1528]) & (layer0_outputs[328]);
    assign outputs[3839] = (layer0_outputs[945]) & ~(layer0_outputs[4963]);
    assign outputs[3840] = ~(layer0_outputs[107]);
    assign outputs[3841] = (layer0_outputs[368]) | (layer0_outputs[3931]);
    assign outputs[3842] = ~((layer0_outputs[1145]) & (layer0_outputs[3519]));
    assign outputs[3843] = (layer0_outputs[6954]) & ~(layer0_outputs[5762]);
    assign outputs[3844] = ~(layer0_outputs[3615]);
    assign outputs[3845] = ~((layer0_outputs[5428]) & (layer0_outputs[5127]));
    assign outputs[3846] = ~(layer0_outputs[3989]);
    assign outputs[3847] = ~((layer0_outputs[805]) & (layer0_outputs[3871]));
    assign outputs[3848] = (layer0_outputs[1497]) ^ (layer0_outputs[4149]);
    assign outputs[3849] = layer0_outputs[7171];
    assign outputs[3850] = layer0_outputs[3727];
    assign outputs[3851] = ~(layer0_outputs[5879]);
    assign outputs[3852] = ~((layer0_outputs[3456]) ^ (layer0_outputs[5379]));
    assign outputs[3853] = ~((layer0_outputs[7098]) & (layer0_outputs[5084]));
    assign outputs[3854] = ~((layer0_outputs[6054]) | (layer0_outputs[5755]));
    assign outputs[3855] = ~(layer0_outputs[2928]) | (layer0_outputs[2006]);
    assign outputs[3856] = layer0_outputs[2841];
    assign outputs[3857] = ~(layer0_outputs[2034]);
    assign outputs[3858] = ~(layer0_outputs[4457]) | (layer0_outputs[656]);
    assign outputs[3859] = ~((layer0_outputs[4367]) ^ (layer0_outputs[2360]));
    assign outputs[3860] = (layer0_outputs[4341]) ^ (layer0_outputs[2678]);
    assign outputs[3861] = ~((layer0_outputs[5564]) & (layer0_outputs[4270]));
    assign outputs[3862] = layer0_outputs[6246];
    assign outputs[3863] = ~((layer0_outputs[5133]) | (layer0_outputs[5780]));
    assign outputs[3864] = ~((layer0_outputs[4102]) ^ (layer0_outputs[7482]));
    assign outputs[3865] = layer0_outputs[3893];
    assign outputs[3866] = ~(layer0_outputs[4778]);
    assign outputs[3867] = layer0_outputs[1834];
    assign outputs[3868] = (layer0_outputs[5981]) ^ (layer0_outputs[956]);
    assign outputs[3869] = (layer0_outputs[497]) | (layer0_outputs[6930]);
    assign outputs[3870] = ~((layer0_outputs[6080]) ^ (layer0_outputs[6916]));
    assign outputs[3871] = ~(layer0_outputs[882]);
    assign outputs[3872] = ~((layer0_outputs[5605]) ^ (layer0_outputs[3798]));
    assign outputs[3873] = ~((layer0_outputs[2835]) ^ (layer0_outputs[4679]));
    assign outputs[3874] = ~((layer0_outputs[6333]) & (layer0_outputs[6885]));
    assign outputs[3875] = ~(layer0_outputs[3766]);
    assign outputs[3876] = ~(layer0_outputs[1141]) | (layer0_outputs[2774]);
    assign outputs[3877] = ~((layer0_outputs[386]) ^ (layer0_outputs[7198]));
    assign outputs[3878] = (layer0_outputs[2709]) ^ (layer0_outputs[6497]);
    assign outputs[3879] = ~((layer0_outputs[498]) | (layer0_outputs[6075]));
    assign outputs[3880] = ~(layer0_outputs[6921]);
    assign outputs[3881] = ~(layer0_outputs[3396]);
    assign outputs[3882] = (layer0_outputs[3002]) ^ (layer0_outputs[3928]);
    assign outputs[3883] = (layer0_outputs[1562]) | (layer0_outputs[2918]);
    assign outputs[3884] = ~(layer0_outputs[2198]);
    assign outputs[3885] = layer0_outputs[6568];
    assign outputs[3886] = ~((layer0_outputs[4637]) ^ (layer0_outputs[4860]));
    assign outputs[3887] = (layer0_outputs[1889]) & ~(layer0_outputs[6135]);
    assign outputs[3888] = ~((layer0_outputs[571]) ^ (layer0_outputs[3463]));
    assign outputs[3889] = layer0_outputs[7282];
    assign outputs[3890] = (layer0_outputs[4187]) & ~(layer0_outputs[7347]);
    assign outputs[3891] = ~((layer0_outputs[3292]) ^ (layer0_outputs[1904]));
    assign outputs[3892] = (layer0_outputs[5586]) & ~(layer0_outputs[3642]);
    assign outputs[3893] = ~((layer0_outputs[3132]) | (layer0_outputs[4697]));
    assign outputs[3894] = ~((layer0_outputs[3611]) ^ (layer0_outputs[2654]));
    assign outputs[3895] = ~((layer0_outputs[6953]) ^ (layer0_outputs[6960]));
    assign outputs[3896] = ~(layer0_outputs[5654]) | (layer0_outputs[1995]);
    assign outputs[3897] = ~(layer0_outputs[4580]);
    assign outputs[3898] = (layer0_outputs[4701]) & (layer0_outputs[6906]);
    assign outputs[3899] = ~((layer0_outputs[5329]) ^ (layer0_outputs[2396]));
    assign outputs[3900] = layer0_outputs[5470];
    assign outputs[3901] = ~(layer0_outputs[6927]);
    assign outputs[3902] = ~((layer0_outputs[612]) & (layer0_outputs[2611]));
    assign outputs[3903] = ~(layer0_outputs[1990]);
    assign outputs[3904] = ~(layer0_outputs[1994]);
    assign outputs[3905] = ~((layer0_outputs[34]) & (layer0_outputs[668]));
    assign outputs[3906] = ~(layer0_outputs[5906]);
    assign outputs[3907] = ~(layer0_outputs[1579]);
    assign outputs[3908] = ~((layer0_outputs[6912]) ^ (layer0_outputs[5836]));
    assign outputs[3909] = layer0_outputs[6222];
    assign outputs[3910] = ~((layer0_outputs[126]) ^ (layer0_outputs[6564]));
    assign outputs[3911] = ~(layer0_outputs[7559]);
    assign outputs[3912] = ~(layer0_outputs[651]);
    assign outputs[3913] = layer0_outputs[6002];
    assign outputs[3914] = ~(layer0_outputs[2976]);
    assign outputs[3915] = (layer0_outputs[761]) | (layer0_outputs[1605]);
    assign outputs[3916] = ~((layer0_outputs[1919]) ^ (layer0_outputs[406]));
    assign outputs[3917] = (layer0_outputs[7116]) ^ (layer0_outputs[3253]);
    assign outputs[3918] = layer0_outputs[3785];
    assign outputs[3919] = ~(layer0_outputs[2804]);
    assign outputs[3920] = ~(layer0_outputs[4712]);
    assign outputs[3921] = (layer0_outputs[2737]) & (layer0_outputs[2688]);
    assign outputs[3922] = ~(layer0_outputs[1997]);
    assign outputs[3923] = ~(layer0_outputs[5845]);
    assign outputs[3924] = ~((layer0_outputs[6739]) & (layer0_outputs[4370]));
    assign outputs[3925] = layer0_outputs[6567];
    assign outputs[3926] = layer0_outputs[1477];
    assign outputs[3927] = ~(layer0_outputs[1650]);
    assign outputs[3928] = ~(layer0_outputs[3546]);
    assign outputs[3929] = layer0_outputs[4891];
    assign outputs[3930] = (layer0_outputs[4992]) ^ (layer0_outputs[5902]);
    assign outputs[3931] = ~(layer0_outputs[4411]);
    assign outputs[3932] = ~(layer0_outputs[4810]);
    assign outputs[3933] = 1'b1;
    assign outputs[3934] = ~(layer0_outputs[7186]);
    assign outputs[3935] = (layer0_outputs[2052]) & (layer0_outputs[6576]);
    assign outputs[3936] = (layer0_outputs[4224]) & ~(layer0_outputs[2389]);
    assign outputs[3937] = 1'b1;
    assign outputs[3938] = layer0_outputs[2267];
    assign outputs[3939] = ~(layer0_outputs[5381]) | (layer0_outputs[5920]);
    assign outputs[3940] = ~(layer0_outputs[1718]);
    assign outputs[3941] = layer0_outputs[4075];
    assign outputs[3942] = layer0_outputs[4650];
    assign outputs[3943] = ~(layer0_outputs[2344]);
    assign outputs[3944] = (layer0_outputs[7270]) ^ (layer0_outputs[1122]);
    assign outputs[3945] = ~(layer0_outputs[5571]);
    assign outputs[3946] = (layer0_outputs[5311]) ^ (layer0_outputs[1367]);
    assign outputs[3947] = ~(layer0_outputs[2044]);
    assign outputs[3948] = 1'b1;
    assign outputs[3949] = ~(layer0_outputs[833]);
    assign outputs[3950] = ~((layer0_outputs[1766]) ^ (layer0_outputs[5022]));
    assign outputs[3951] = ~(layer0_outputs[1811]);
    assign outputs[3952] = (layer0_outputs[3000]) ^ (layer0_outputs[600]);
    assign outputs[3953] = (layer0_outputs[5600]) & ~(layer0_outputs[5131]);
    assign outputs[3954] = ~(layer0_outputs[4181]);
    assign outputs[3955] = ~((layer0_outputs[4081]) ^ (layer0_outputs[2840]));
    assign outputs[3956] = ~(layer0_outputs[6108]);
    assign outputs[3957] = ~((layer0_outputs[3055]) ^ (layer0_outputs[5844]));
    assign outputs[3958] = ~(layer0_outputs[1929]);
    assign outputs[3959] = (layer0_outputs[1684]) & (layer0_outputs[5713]);
    assign outputs[3960] = (layer0_outputs[3039]) ^ (layer0_outputs[5838]);
    assign outputs[3961] = (layer0_outputs[6569]) & ~(layer0_outputs[460]);
    assign outputs[3962] = ~((layer0_outputs[4575]) ^ (layer0_outputs[5140]));
    assign outputs[3963] = (layer0_outputs[6193]) ^ (layer0_outputs[2848]);
    assign outputs[3964] = ~((layer0_outputs[3728]) ^ (layer0_outputs[4294]));
    assign outputs[3965] = layer0_outputs[4482];
    assign outputs[3966] = (layer0_outputs[4282]) ^ (layer0_outputs[5566]);
    assign outputs[3967] = ~(layer0_outputs[717]);
    assign outputs[3968] = layer0_outputs[1570];
    assign outputs[3969] = ~(layer0_outputs[7125]);
    assign outputs[3970] = (layer0_outputs[354]) & (layer0_outputs[7520]);
    assign outputs[3971] = layer0_outputs[2798];
    assign outputs[3972] = layer0_outputs[1634];
    assign outputs[3973] = (layer0_outputs[1693]) ^ (layer0_outputs[7645]);
    assign outputs[3974] = (layer0_outputs[4764]) ^ (layer0_outputs[957]);
    assign outputs[3975] = ~(layer0_outputs[2577]);
    assign outputs[3976] = layer0_outputs[5453];
    assign outputs[3977] = layer0_outputs[5430];
    assign outputs[3978] = (layer0_outputs[4771]) & ~(layer0_outputs[2805]);
    assign outputs[3979] = layer0_outputs[284];
    assign outputs[3980] = ~((layer0_outputs[938]) & (layer0_outputs[6076]));
    assign outputs[3981] = ~((layer0_outputs[1633]) & (layer0_outputs[673]));
    assign outputs[3982] = ~(layer0_outputs[4672]);
    assign outputs[3983] = ~(layer0_outputs[6809]);
    assign outputs[3984] = ~((layer0_outputs[1946]) | (layer0_outputs[818]));
    assign outputs[3985] = ~((layer0_outputs[3401]) | (layer0_outputs[3891]));
    assign outputs[3986] = layer0_outputs[5530];
    assign outputs[3987] = (layer0_outputs[6561]) ^ (layer0_outputs[920]);
    assign outputs[3988] = ~(layer0_outputs[4780]);
    assign outputs[3989] = ~(layer0_outputs[4618]);
    assign outputs[3990] = ~(layer0_outputs[3576]);
    assign outputs[3991] = layer0_outputs[981];
    assign outputs[3992] = (layer0_outputs[2940]) ^ (layer0_outputs[3527]);
    assign outputs[3993] = layer0_outputs[35];
    assign outputs[3994] = ~(layer0_outputs[4586]);
    assign outputs[3995] = layer0_outputs[434];
    assign outputs[3996] = (layer0_outputs[6887]) | (layer0_outputs[6431]);
    assign outputs[3997] = layer0_outputs[1891];
    assign outputs[3998] = layer0_outputs[1395];
    assign outputs[3999] = ~((layer0_outputs[6636]) ^ (layer0_outputs[4517]));
    assign outputs[4000] = (layer0_outputs[20]) ^ (layer0_outputs[4982]);
    assign outputs[4001] = (layer0_outputs[5991]) ^ (layer0_outputs[7070]);
    assign outputs[4002] = ~((layer0_outputs[4475]) & (layer0_outputs[6]));
    assign outputs[4003] = layer0_outputs[6922];
    assign outputs[4004] = ~(layer0_outputs[6354]);
    assign outputs[4005] = ~(layer0_outputs[3121]);
    assign outputs[4006] = ~((layer0_outputs[6060]) & (layer0_outputs[1338]));
    assign outputs[4007] = (layer0_outputs[3677]) | (layer0_outputs[3237]);
    assign outputs[4008] = (layer0_outputs[6351]) ^ (layer0_outputs[4441]);
    assign outputs[4009] = (layer0_outputs[5724]) ^ (layer0_outputs[7043]);
    assign outputs[4010] = (layer0_outputs[5670]) & (layer0_outputs[932]);
    assign outputs[4011] = ~((layer0_outputs[3449]) & (layer0_outputs[3527]));
    assign outputs[4012] = (layer0_outputs[5985]) ^ (layer0_outputs[3241]);
    assign outputs[4013] = ~(layer0_outputs[4411]);
    assign outputs[4014] = (layer0_outputs[2706]) ^ (layer0_outputs[2193]);
    assign outputs[4015] = ~(layer0_outputs[2300]);
    assign outputs[4016] = ~(layer0_outputs[5934]) | (layer0_outputs[4813]);
    assign outputs[4017] = (layer0_outputs[471]) | (layer0_outputs[3116]);
    assign outputs[4018] = ~(layer0_outputs[5526]);
    assign outputs[4019] = ~(layer0_outputs[1368]);
    assign outputs[4020] = layer0_outputs[5252];
    assign outputs[4021] = ~(layer0_outputs[1865]) | (layer0_outputs[2011]);
    assign outputs[4022] = layer0_outputs[3502];
    assign outputs[4023] = ~(layer0_outputs[2807]);
    assign outputs[4024] = ~(layer0_outputs[5425]);
    assign outputs[4025] = ~((layer0_outputs[6523]) ^ (layer0_outputs[818]));
    assign outputs[4026] = layer0_outputs[3502];
    assign outputs[4027] = ~(layer0_outputs[6300]);
    assign outputs[4028] = layer0_outputs[1493];
    assign outputs[4029] = ~((layer0_outputs[2261]) ^ (layer0_outputs[906]));
    assign outputs[4030] = layer0_outputs[5534];
    assign outputs[4031] = layer0_outputs[4795];
    assign outputs[4032] = layer0_outputs[4555];
    assign outputs[4033] = (layer0_outputs[7138]) ^ (layer0_outputs[6624]);
    assign outputs[4034] = ~(layer0_outputs[4796]) | (layer0_outputs[345]);
    assign outputs[4035] = ~(layer0_outputs[725]);
    assign outputs[4036] = (layer0_outputs[6768]) ^ (layer0_outputs[5946]);
    assign outputs[4037] = layer0_outputs[5075];
    assign outputs[4038] = (layer0_outputs[3226]) ^ (layer0_outputs[3216]);
    assign outputs[4039] = ~(layer0_outputs[209]) | (layer0_outputs[536]);
    assign outputs[4040] = layer0_outputs[3888];
    assign outputs[4041] = (layer0_outputs[749]) ^ (layer0_outputs[1817]);
    assign outputs[4042] = ~((layer0_outputs[1010]) ^ (layer0_outputs[4338]));
    assign outputs[4043] = layer0_outputs[154];
    assign outputs[4044] = (layer0_outputs[1806]) | (layer0_outputs[6951]);
    assign outputs[4045] = ~(layer0_outputs[7403]) | (layer0_outputs[2161]);
    assign outputs[4046] = ~(layer0_outputs[4808]);
    assign outputs[4047] = (layer0_outputs[5568]) & (layer0_outputs[4622]);
    assign outputs[4048] = layer0_outputs[1395];
    assign outputs[4049] = layer0_outputs[3330];
    assign outputs[4050] = ~((layer0_outputs[1730]) ^ (layer0_outputs[4013]));
    assign outputs[4051] = layer0_outputs[5168];
    assign outputs[4052] = layer0_outputs[6629];
    assign outputs[4053] = (layer0_outputs[7184]) & ~(layer0_outputs[1293]);
    assign outputs[4054] = ~(layer0_outputs[6924]);
    assign outputs[4055] = layer0_outputs[5016];
    assign outputs[4056] = ~((layer0_outputs[5096]) ^ (layer0_outputs[6031]));
    assign outputs[4057] = layer0_outputs[1515];
    assign outputs[4058] = (layer0_outputs[323]) ^ (layer0_outputs[4436]);
    assign outputs[4059] = layer0_outputs[984];
    assign outputs[4060] = layer0_outputs[7048];
    assign outputs[4061] = ~(layer0_outputs[6393]);
    assign outputs[4062] = ~(layer0_outputs[7050]);
    assign outputs[4063] = layer0_outputs[370];
    assign outputs[4064] = layer0_outputs[6495];
    assign outputs[4065] = ~((layer0_outputs[2996]) ^ (layer0_outputs[5589]));
    assign outputs[4066] = layer0_outputs[7189];
    assign outputs[4067] = (layer0_outputs[2587]) ^ (layer0_outputs[1422]);
    assign outputs[4068] = ~(layer0_outputs[3833]);
    assign outputs[4069] = (layer0_outputs[2618]) & ~(layer0_outputs[7491]);
    assign outputs[4070] = ~((layer0_outputs[7183]) ^ (layer0_outputs[2002]));
    assign outputs[4071] = layer0_outputs[444];
    assign outputs[4072] = ~((layer0_outputs[5024]) & (layer0_outputs[951]));
    assign outputs[4073] = (layer0_outputs[3825]) ^ (layer0_outputs[2981]);
    assign outputs[4074] = 1'b1;
    assign outputs[4075] = ~((layer0_outputs[974]) & (layer0_outputs[6044]));
    assign outputs[4076] = (layer0_outputs[6754]) ^ (layer0_outputs[52]);
    assign outputs[4077] = ~(layer0_outputs[1506]) | (layer0_outputs[6499]);
    assign outputs[4078] = ~(layer0_outputs[40]);
    assign outputs[4079] = layer0_outputs[2380];
    assign outputs[4080] = (layer0_outputs[3300]) ^ (layer0_outputs[4899]);
    assign outputs[4081] = ~(layer0_outputs[5170]);
    assign outputs[4082] = layer0_outputs[3512];
    assign outputs[4083] = ~((layer0_outputs[255]) ^ (layer0_outputs[1642]));
    assign outputs[4084] = ~((layer0_outputs[158]) ^ (layer0_outputs[4799]));
    assign outputs[4085] = ~((layer0_outputs[1752]) ^ (layer0_outputs[7120]));
    assign outputs[4086] = ~((layer0_outputs[2064]) ^ (layer0_outputs[5594]));
    assign outputs[4087] = (layer0_outputs[1938]) & (layer0_outputs[654]);
    assign outputs[4088] = ~((layer0_outputs[2497]) & (layer0_outputs[4933]));
    assign outputs[4089] = ~(layer0_outputs[700]);
    assign outputs[4090] = (layer0_outputs[3242]) & (layer0_outputs[3481]);
    assign outputs[4091] = ~((layer0_outputs[781]) | (layer0_outputs[4502]));
    assign outputs[4092] = ~(layer0_outputs[5708]);
    assign outputs[4093] = layer0_outputs[3894];
    assign outputs[4094] = ~(layer0_outputs[6946]);
    assign outputs[4095] = layer0_outputs[4443];
    assign outputs[4096] = ~(layer0_outputs[6044]);
    assign outputs[4097] = ~(layer0_outputs[5949]);
    assign outputs[4098] = ~(layer0_outputs[6437]);
    assign outputs[4099] = layer0_outputs[5189];
    assign outputs[4100] = layer0_outputs[2249];
    assign outputs[4101] = ~((layer0_outputs[1166]) ^ (layer0_outputs[2057]));
    assign outputs[4102] = (layer0_outputs[5289]) | (layer0_outputs[4042]);
    assign outputs[4103] = ~((layer0_outputs[7562]) ^ (layer0_outputs[2715]));
    assign outputs[4104] = ~(layer0_outputs[2884]) | (layer0_outputs[5657]);
    assign outputs[4105] = layer0_outputs[172];
    assign outputs[4106] = layer0_outputs[5642];
    assign outputs[4107] = ~((layer0_outputs[3567]) & (layer0_outputs[2898]));
    assign outputs[4108] = layer0_outputs[1986];
    assign outputs[4109] = (layer0_outputs[527]) ^ (layer0_outputs[4459]);
    assign outputs[4110] = layer0_outputs[1711];
    assign outputs[4111] = ~(layer0_outputs[4304]);
    assign outputs[4112] = ~((layer0_outputs[348]) ^ (layer0_outputs[4368]));
    assign outputs[4113] = ~((layer0_outputs[3263]) ^ (layer0_outputs[636]));
    assign outputs[4114] = layer0_outputs[7660];
    assign outputs[4115] = layer0_outputs[296];
    assign outputs[4116] = ~((layer0_outputs[2706]) ^ (layer0_outputs[6362]));
    assign outputs[4117] = (layer0_outputs[308]) ^ (layer0_outputs[5418]);
    assign outputs[4118] = ~(layer0_outputs[1597]);
    assign outputs[4119] = ~(layer0_outputs[3617]);
    assign outputs[4120] = ~(layer0_outputs[7035]);
    assign outputs[4121] = (layer0_outputs[6947]) & ~(layer0_outputs[3817]);
    assign outputs[4122] = ~(layer0_outputs[7506]) | (layer0_outputs[3514]);
    assign outputs[4123] = ~((layer0_outputs[2947]) ^ (layer0_outputs[6182]));
    assign outputs[4124] = (layer0_outputs[4782]) & (layer0_outputs[984]);
    assign outputs[4125] = layer0_outputs[7572];
    assign outputs[4126] = (layer0_outputs[1315]) & ~(layer0_outputs[6033]);
    assign outputs[4127] = layer0_outputs[4760];
    assign outputs[4128] = (layer0_outputs[5487]) ^ (layer0_outputs[679]);
    assign outputs[4129] = ~((layer0_outputs[3234]) | (layer0_outputs[2226]));
    assign outputs[4130] = layer0_outputs[1803];
    assign outputs[4131] = ~(layer0_outputs[1527]);
    assign outputs[4132] = ~((layer0_outputs[7139]) ^ (layer0_outputs[4546]));
    assign outputs[4133] = (layer0_outputs[5062]) ^ (layer0_outputs[2547]);
    assign outputs[4134] = layer0_outputs[3301];
    assign outputs[4135] = ~((layer0_outputs[7098]) & (layer0_outputs[1541]));
    assign outputs[4136] = layer0_outputs[3320];
    assign outputs[4137] = ~((layer0_outputs[6860]) ^ (layer0_outputs[7221]));
    assign outputs[4138] = ~(layer0_outputs[5552]);
    assign outputs[4139] = 1'b1;
    assign outputs[4140] = ~((layer0_outputs[1532]) | (layer0_outputs[213]));
    assign outputs[4141] = ~((layer0_outputs[3409]) ^ (layer0_outputs[2213]));
    assign outputs[4142] = ~(layer0_outputs[1797]);
    assign outputs[4143] = ~(layer0_outputs[4244]);
    assign outputs[4144] = ~((layer0_outputs[5992]) ^ (layer0_outputs[7668]));
    assign outputs[4145] = (layer0_outputs[2479]) ^ (layer0_outputs[6961]);
    assign outputs[4146] = (layer0_outputs[6963]) ^ (layer0_outputs[6000]);
    assign outputs[4147] = layer0_outputs[5853];
    assign outputs[4148] = (layer0_outputs[617]) ^ (layer0_outputs[3511]);
    assign outputs[4149] = layer0_outputs[7660];
    assign outputs[4150] = ~(layer0_outputs[2524]) | (layer0_outputs[5279]);
    assign outputs[4151] = (layer0_outputs[6879]) & ~(layer0_outputs[3722]);
    assign outputs[4152] = (layer0_outputs[3551]) ^ (layer0_outputs[742]);
    assign outputs[4153] = (layer0_outputs[2790]) ^ (layer0_outputs[6717]);
    assign outputs[4154] = ~(layer0_outputs[4262]);
    assign outputs[4155] = ~(layer0_outputs[522]) | (layer0_outputs[3479]);
    assign outputs[4156] = ~((layer0_outputs[5119]) ^ (layer0_outputs[5494]));
    assign outputs[4157] = layer0_outputs[7634];
    assign outputs[4158] = ~(layer0_outputs[2231]) | (layer0_outputs[2541]);
    assign outputs[4159] = ~((layer0_outputs[3032]) ^ (layer0_outputs[2302]));
    assign outputs[4160] = ~(layer0_outputs[4901]);
    assign outputs[4161] = ~(layer0_outputs[5554]) | (layer0_outputs[2935]);
    assign outputs[4162] = ~((layer0_outputs[2611]) ^ (layer0_outputs[561]));
    assign outputs[4163] = layer0_outputs[5135];
    assign outputs[4164] = (layer0_outputs[5633]) & (layer0_outputs[1787]);
    assign outputs[4165] = ~((layer0_outputs[21]) | (layer0_outputs[2674]));
    assign outputs[4166] = ~(layer0_outputs[1839]);
    assign outputs[4167] = ~((layer0_outputs[6729]) ^ (layer0_outputs[237]));
    assign outputs[4168] = ~(layer0_outputs[2405]);
    assign outputs[4169] = ~((layer0_outputs[1297]) ^ (layer0_outputs[6040]));
    assign outputs[4170] = ~((layer0_outputs[4365]) & (layer0_outputs[1485]));
    assign outputs[4171] = ~((layer0_outputs[1610]) & (layer0_outputs[5053]));
    assign outputs[4172] = ~((layer0_outputs[2229]) ^ (layer0_outputs[5199]));
    assign outputs[4173] = (layer0_outputs[2375]) ^ (layer0_outputs[1278]);
    assign outputs[4174] = ~((layer0_outputs[5019]) ^ (layer0_outputs[199]));
    assign outputs[4175] = ~((layer0_outputs[3136]) ^ (layer0_outputs[719]));
    assign outputs[4176] = (layer0_outputs[256]) | (layer0_outputs[7192]);
    assign outputs[4177] = (layer0_outputs[6070]) & (layer0_outputs[7566]);
    assign outputs[4178] = ~(layer0_outputs[1827]);
    assign outputs[4179] = ~((layer0_outputs[7289]) ^ (layer0_outputs[3742]));
    assign outputs[4180] = layer0_outputs[1392];
    assign outputs[4181] = ~((layer0_outputs[6094]) & (layer0_outputs[4039]));
    assign outputs[4182] = ~(layer0_outputs[7222]);
    assign outputs[4183] = layer0_outputs[5504];
    assign outputs[4184] = layer0_outputs[4626];
    assign outputs[4185] = (layer0_outputs[3047]) ^ (layer0_outputs[3173]);
    assign outputs[4186] = ~((layer0_outputs[4885]) | (layer0_outputs[3777]));
    assign outputs[4187] = ~(layer0_outputs[5513]);
    assign outputs[4188] = ~(layer0_outputs[2443]) | (layer0_outputs[521]);
    assign outputs[4189] = ~((layer0_outputs[949]) ^ (layer0_outputs[7115]));
    assign outputs[4190] = ~(layer0_outputs[6310]);
    assign outputs[4191] = layer0_outputs[6758];
    assign outputs[4192] = ~((layer0_outputs[1387]) ^ (layer0_outputs[155]));
    assign outputs[4193] = ~((layer0_outputs[5590]) ^ (layer0_outputs[2429]));
    assign outputs[4194] = layer0_outputs[5048];
    assign outputs[4195] = layer0_outputs[733];
    assign outputs[4196] = ~(layer0_outputs[5294]) | (layer0_outputs[3375]);
    assign outputs[4197] = (layer0_outputs[4615]) & ~(layer0_outputs[1508]);
    assign outputs[4198] = ~((layer0_outputs[1502]) ^ (layer0_outputs[7470]));
    assign outputs[4199] = ~(layer0_outputs[5932]) | (layer0_outputs[1612]);
    assign outputs[4200] = layer0_outputs[869];
    assign outputs[4201] = ~((layer0_outputs[2759]) ^ (layer0_outputs[4832]));
    assign outputs[4202] = ~((layer0_outputs[3884]) & (layer0_outputs[6668]));
    assign outputs[4203] = ~((layer0_outputs[3847]) ^ (layer0_outputs[4574]));
    assign outputs[4204] = ~(layer0_outputs[4571]);
    assign outputs[4205] = ~(layer0_outputs[1704]) | (layer0_outputs[3280]);
    assign outputs[4206] = ~((layer0_outputs[6623]) ^ (layer0_outputs[6118]));
    assign outputs[4207] = ~(layer0_outputs[2787]);
    assign outputs[4208] = (layer0_outputs[7443]) & (layer0_outputs[756]);
    assign outputs[4209] = ~(layer0_outputs[4184]) | (layer0_outputs[6000]);
    assign outputs[4210] = ~(layer0_outputs[4250]);
    assign outputs[4211] = ~((layer0_outputs[7085]) ^ (layer0_outputs[2975]));
    assign outputs[4212] = ~(layer0_outputs[7627]);
    assign outputs[4213] = ~(layer0_outputs[7619]);
    assign outputs[4214] = (layer0_outputs[3974]) & ~(layer0_outputs[646]);
    assign outputs[4215] = layer0_outputs[2179];
    assign outputs[4216] = ~(layer0_outputs[6487]);
    assign outputs[4217] = ~((layer0_outputs[1548]) ^ (layer0_outputs[836]));
    assign outputs[4218] = ~((layer0_outputs[3254]) & (layer0_outputs[5700]));
    assign outputs[4219] = ~(layer0_outputs[1927]);
    assign outputs[4220] = ~(layer0_outputs[2154]);
    assign outputs[4221] = (layer0_outputs[3774]) | (layer0_outputs[4993]);
    assign outputs[4222] = ~(layer0_outputs[3652]);
    assign outputs[4223] = (layer0_outputs[4817]) ^ (layer0_outputs[7643]);
    assign outputs[4224] = layer0_outputs[1096];
    assign outputs[4225] = (layer0_outputs[5198]) & ~(layer0_outputs[7486]);
    assign outputs[4226] = ~(layer0_outputs[6801]);
    assign outputs[4227] = ~((layer0_outputs[4008]) | (layer0_outputs[1160]));
    assign outputs[4228] = ~(layer0_outputs[4787]);
    assign outputs[4229] = (layer0_outputs[6504]) & ~(layer0_outputs[5660]);
    assign outputs[4230] = layer0_outputs[7367];
    assign outputs[4231] = layer0_outputs[2206];
    assign outputs[4232] = layer0_outputs[3406];
    assign outputs[4233] = ~(layer0_outputs[3652]);
    assign outputs[4234] = ~(layer0_outputs[2165]);
    assign outputs[4235] = ~(layer0_outputs[2503]);
    assign outputs[4236] = (layer0_outputs[4019]) & ~(layer0_outputs[3568]);
    assign outputs[4237] = layer0_outputs[6322];
    assign outputs[4238] = ~(layer0_outputs[3349]);
    assign outputs[4239] = ~((layer0_outputs[2880]) ^ (layer0_outputs[2453]));
    assign outputs[4240] = ~((layer0_outputs[1140]) & (layer0_outputs[894]));
    assign outputs[4241] = ~((layer0_outputs[2829]) ^ (layer0_outputs[1053]));
    assign outputs[4242] = layer0_outputs[4535];
    assign outputs[4243] = (layer0_outputs[6720]) ^ (layer0_outputs[4179]);
    assign outputs[4244] = ~(layer0_outputs[506]) | (layer0_outputs[6805]);
    assign outputs[4245] = ~(layer0_outputs[5672]);
    assign outputs[4246] = ~(layer0_outputs[7611]) | (layer0_outputs[5471]);
    assign outputs[4247] = ~(layer0_outputs[1139]);
    assign outputs[4248] = ~(layer0_outputs[2437]);
    assign outputs[4249] = ~(layer0_outputs[3162]);
    assign outputs[4250] = (layer0_outputs[4683]) & (layer0_outputs[2815]);
    assign outputs[4251] = (layer0_outputs[3854]) ^ (layer0_outputs[2942]);
    assign outputs[4252] = ~((layer0_outputs[5353]) ^ (layer0_outputs[571]));
    assign outputs[4253] = ~(layer0_outputs[337]);
    assign outputs[4254] = ~(layer0_outputs[6261]);
    assign outputs[4255] = layer0_outputs[7477];
    assign outputs[4256] = ~((layer0_outputs[5490]) ^ (layer0_outputs[5068]));
    assign outputs[4257] = layer0_outputs[777];
    assign outputs[4258] = layer0_outputs[1922];
    assign outputs[4259] = ~(layer0_outputs[1269]);
    assign outputs[4260] = ~(layer0_outputs[789]);
    assign outputs[4261] = ~((layer0_outputs[1624]) ^ (layer0_outputs[5718]));
    assign outputs[4262] = layer0_outputs[1184];
    assign outputs[4263] = (layer0_outputs[2026]) | (layer0_outputs[32]);
    assign outputs[4264] = (layer0_outputs[3217]) & ~(layer0_outputs[400]);
    assign outputs[4265] = layer0_outputs[5658];
    assign outputs[4266] = ~((layer0_outputs[5041]) & (layer0_outputs[2289]));
    assign outputs[4267] = (layer0_outputs[1385]) & (layer0_outputs[4614]);
    assign outputs[4268] = (layer0_outputs[4487]) | (layer0_outputs[7639]);
    assign outputs[4269] = ~(layer0_outputs[914]);
    assign outputs[4270] = layer0_outputs[3953];
    assign outputs[4271] = layer0_outputs[326];
    assign outputs[4272] = layer0_outputs[6427];
    assign outputs[4273] = ~((layer0_outputs[6154]) ^ (layer0_outputs[1985]));
    assign outputs[4274] = ~((layer0_outputs[4235]) | (layer0_outputs[553]));
    assign outputs[4275] = layer0_outputs[2712];
    assign outputs[4276] = layer0_outputs[2071];
    assign outputs[4277] = ~(layer0_outputs[5561]) | (layer0_outputs[5550]);
    assign outputs[4278] = (layer0_outputs[4501]) | (layer0_outputs[3471]);
    assign outputs[4279] = ~(layer0_outputs[7027]);
    assign outputs[4280] = ~(layer0_outputs[1955]) | (layer0_outputs[782]);
    assign outputs[4281] = ~(layer0_outputs[3845]);
    assign outputs[4282] = (layer0_outputs[4729]) ^ (layer0_outputs[6511]);
    assign outputs[4283] = ~(layer0_outputs[5768]);
    assign outputs[4284] = ~((layer0_outputs[776]) ^ (layer0_outputs[4915]));
    assign outputs[4285] = ~((layer0_outputs[19]) | (layer0_outputs[4121]));
    assign outputs[4286] = ~((layer0_outputs[7219]) & (layer0_outputs[4981]));
    assign outputs[4287] = ~((layer0_outputs[7020]) | (layer0_outputs[6744]));
    assign outputs[4288] = (layer0_outputs[7483]) & (layer0_outputs[2780]);
    assign outputs[4289] = ~(layer0_outputs[2667]);
    assign outputs[4290] = ~(layer0_outputs[263]);
    assign outputs[4291] = layer0_outputs[6398];
    assign outputs[4292] = ~((layer0_outputs[973]) ^ (layer0_outputs[3665]));
    assign outputs[4293] = ~(layer0_outputs[329]);
    assign outputs[4294] = (layer0_outputs[1178]) | (layer0_outputs[5286]);
    assign outputs[4295] = ~((layer0_outputs[6282]) | (layer0_outputs[412]));
    assign outputs[4296] = layer0_outputs[2242];
    assign outputs[4297] = ~(layer0_outputs[4715]) | (layer0_outputs[4140]);
    assign outputs[4298] = layer0_outputs[6401];
    assign outputs[4299] = (layer0_outputs[1359]) ^ (layer0_outputs[6092]);
    assign outputs[4300] = ~(layer0_outputs[95]);
    assign outputs[4301] = ~(layer0_outputs[5772]);
    assign outputs[4302] = ~(layer0_outputs[6104]) | (layer0_outputs[2545]);
    assign outputs[4303] = (layer0_outputs[6001]) | (layer0_outputs[6746]);
    assign outputs[4304] = ~(layer0_outputs[3772]);
    assign outputs[4305] = layer0_outputs[5152];
    assign outputs[4306] = ~((layer0_outputs[2860]) ^ (layer0_outputs[5374]));
    assign outputs[4307] = (layer0_outputs[2885]) & ~(layer0_outputs[1389]);
    assign outputs[4308] = layer0_outputs[1402];
    assign outputs[4309] = layer0_outputs[972];
    assign outputs[4310] = (layer0_outputs[6381]) ^ (layer0_outputs[2274]);
    assign outputs[4311] = ~(layer0_outputs[5221]);
    assign outputs[4312] = (layer0_outputs[6560]) ^ (layer0_outputs[3560]);
    assign outputs[4313] = ~((layer0_outputs[4402]) ^ (layer0_outputs[4328]));
    assign outputs[4314] = (layer0_outputs[1587]) ^ (layer0_outputs[6297]);
    assign outputs[4315] = ~(layer0_outputs[5520]);
    assign outputs[4316] = layer0_outputs[7673];
    assign outputs[4317] = (layer0_outputs[3554]) ^ (layer0_outputs[3388]);
    assign outputs[4318] = ~((layer0_outputs[1212]) | (layer0_outputs[3624]));
    assign outputs[4319] = ~(layer0_outputs[249]);
    assign outputs[4320] = ~(layer0_outputs[1683]) | (layer0_outputs[2956]);
    assign outputs[4321] = ~((layer0_outputs[1471]) ^ (layer0_outputs[3657]));
    assign outputs[4322] = ~(layer0_outputs[3598]);
    assign outputs[4323] = ~((layer0_outputs[4919]) & (layer0_outputs[1565]));
    assign outputs[4324] = ~((layer0_outputs[1816]) ^ (layer0_outputs[3374]));
    assign outputs[4325] = layer0_outputs[211];
    assign outputs[4326] = ~(layer0_outputs[647]) | (layer0_outputs[3748]);
    assign outputs[4327] = ~((layer0_outputs[1424]) & (layer0_outputs[6752]));
    assign outputs[4328] = (layer0_outputs[831]) ^ (layer0_outputs[585]);
    assign outputs[4329] = (layer0_outputs[7479]) | (layer0_outputs[4234]);
    assign outputs[4330] = ~((layer0_outputs[2923]) ^ (layer0_outputs[7602]));
    assign outputs[4331] = ~(layer0_outputs[4467]);
    assign outputs[4332] = layer0_outputs[6298];
    assign outputs[4333] = ~(layer0_outputs[6133]);
    assign outputs[4334] = layer0_outputs[1294];
    assign outputs[4335] = ~((layer0_outputs[4184]) & (layer0_outputs[6016]));
    assign outputs[4336] = ~(layer0_outputs[3864]);
    assign outputs[4337] = (layer0_outputs[607]) & ~(layer0_outputs[2201]);
    assign outputs[4338] = (layer0_outputs[2418]) ^ (layer0_outputs[301]);
    assign outputs[4339] = (layer0_outputs[2568]) ^ (layer0_outputs[6883]);
    assign outputs[4340] = ~((layer0_outputs[6164]) | (layer0_outputs[4931]));
    assign outputs[4341] = ~((layer0_outputs[1045]) & (layer0_outputs[5445]));
    assign outputs[4342] = layer0_outputs[5846];
    assign outputs[4343] = ~(layer0_outputs[5598]);
    assign outputs[4344] = ~(layer0_outputs[549]);
    assign outputs[4345] = (layer0_outputs[2280]) | (layer0_outputs[6441]);
    assign outputs[4346] = ~((layer0_outputs[5413]) & (layer0_outputs[4478]));
    assign outputs[4347] = ~(layer0_outputs[6006]);
    assign outputs[4348] = ~((layer0_outputs[7063]) ^ (layer0_outputs[4358]));
    assign outputs[4349] = (layer0_outputs[1408]) ^ (layer0_outputs[7001]);
    assign outputs[4350] = ~(layer0_outputs[4065]) | (layer0_outputs[6398]);
    assign outputs[4351] = (layer0_outputs[7303]) ^ (layer0_outputs[4768]);
    assign outputs[4352] = (layer0_outputs[7663]) ^ (layer0_outputs[451]);
    assign outputs[4353] = layer0_outputs[6560];
    assign outputs[4354] = layer0_outputs[3077];
    assign outputs[4355] = (layer0_outputs[2409]) & (layer0_outputs[4761]);
    assign outputs[4356] = ~((layer0_outputs[5070]) ^ (layer0_outputs[4851]));
    assign outputs[4357] = ~(layer0_outputs[4554]);
    assign outputs[4358] = (layer0_outputs[370]) & (layer0_outputs[7434]);
    assign outputs[4359] = ~(layer0_outputs[1059]);
    assign outputs[4360] = (layer0_outputs[4716]) & ~(layer0_outputs[1663]);
    assign outputs[4361] = ~((layer0_outputs[6132]) ^ (layer0_outputs[2758]));
    assign outputs[4362] = ~(layer0_outputs[6529]);
    assign outputs[4363] = (layer0_outputs[873]) ^ (layer0_outputs[4908]);
    assign outputs[4364] = ~(layer0_outputs[2931]) | (layer0_outputs[3934]);
    assign outputs[4365] = ~(layer0_outputs[472]);
    assign outputs[4366] = ~(layer0_outputs[196]);
    assign outputs[4367] = ~(layer0_outputs[2844]);
    assign outputs[4368] = (layer0_outputs[1834]) | (layer0_outputs[3622]);
    assign outputs[4369] = ~(layer0_outputs[6490]);
    assign outputs[4370] = ~((layer0_outputs[7361]) | (layer0_outputs[5560]));
    assign outputs[4371] = ~((layer0_outputs[2880]) ^ (layer0_outputs[4600]));
    assign outputs[4372] = (layer0_outputs[4340]) & (layer0_outputs[5330]);
    assign outputs[4373] = (layer0_outputs[1841]) ^ (layer0_outputs[3799]);
    assign outputs[4374] = (layer0_outputs[4692]) ^ (layer0_outputs[5782]);
    assign outputs[4375] = ~((layer0_outputs[7441]) ^ (layer0_outputs[7505]));
    assign outputs[4376] = ~(layer0_outputs[4178]);
    assign outputs[4377] = (layer0_outputs[2029]) & ~(layer0_outputs[7024]);
    assign outputs[4378] = layer0_outputs[2650];
    assign outputs[4379] = layer0_outputs[476];
    assign outputs[4380] = layer0_outputs[4556];
    assign outputs[4381] = layer0_outputs[1735];
    assign outputs[4382] = ~((layer0_outputs[5450]) | (layer0_outputs[4283]));
    assign outputs[4383] = layer0_outputs[3972];
    assign outputs[4384] = ~(layer0_outputs[1007]);
    assign outputs[4385] = ~((layer0_outputs[6627]) ^ (layer0_outputs[2540]));
    assign outputs[4386] = ~((layer0_outputs[644]) & (layer0_outputs[2694]));
    assign outputs[4387] = ~((layer0_outputs[7427]) ^ (layer0_outputs[3577]));
    assign outputs[4388] = ~((layer0_outputs[339]) & (layer0_outputs[7056]));
    assign outputs[4389] = ~(layer0_outputs[645]);
    assign outputs[4390] = ~(layer0_outputs[3189]);
    assign outputs[4391] = ~((layer0_outputs[3250]) ^ (layer0_outputs[3279]));
    assign outputs[4392] = (layer0_outputs[6658]) ^ (layer0_outputs[4654]);
    assign outputs[4393] = (layer0_outputs[6786]) ^ (layer0_outputs[1613]);
    assign outputs[4394] = (layer0_outputs[3262]) & ~(layer0_outputs[1758]);
    assign outputs[4395] = ~(layer0_outputs[6580]) | (layer0_outputs[2172]);
    assign outputs[4396] = layer0_outputs[4245];
    assign outputs[4397] = ~((layer0_outputs[4375]) ^ (layer0_outputs[5410]));
    assign outputs[4398] = (layer0_outputs[1672]) ^ (layer0_outputs[5694]);
    assign outputs[4399] = layer0_outputs[1487];
    assign outputs[4400] = layer0_outputs[2820];
    assign outputs[4401] = (layer0_outputs[1863]) ^ (layer0_outputs[6475]);
    assign outputs[4402] = ~(layer0_outputs[7236]);
    assign outputs[4403] = ~(layer0_outputs[6227]);
    assign outputs[4404] = ~((layer0_outputs[279]) ^ (layer0_outputs[2755]));
    assign outputs[4405] = 1'b1;
    assign outputs[4406] = layer0_outputs[2986];
    assign outputs[4407] = (layer0_outputs[3347]) ^ (layer0_outputs[5908]);
    assign outputs[4408] = ~(layer0_outputs[6059]);
    assign outputs[4409] = (layer0_outputs[7018]) & ~(layer0_outputs[299]);
    assign outputs[4410] = ~(layer0_outputs[2150]);
    assign outputs[4411] = ~(layer0_outputs[4762]);
    assign outputs[4412] = layer0_outputs[869];
    assign outputs[4413] = (layer0_outputs[7332]) & ~(layer0_outputs[5359]);
    assign outputs[4414] = layer0_outputs[3534];
    assign outputs[4415] = ~((layer0_outputs[4105]) | (layer0_outputs[7274]));
    assign outputs[4416] = (layer0_outputs[1112]) | (layer0_outputs[4809]);
    assign outputs[4417] = ~((layer0_outputs[6407]) | (layer0_outputs[1940]));
    assign outputs[4418] = ~(layer0_outputs[59]) | (layer0_outputs[978]);
    assign outputs[4419] = ~(layer0_outputs[6538]);
    assign outputs[4420] = (layer0_outputs[1705]) ^ (layer0_outputs[5859]);
    assign outputs[4421] = (layer0_outputs[4568]) ^ (layer0_outputs[5750]);
    assign outputs[4422] = ~(layer0_outputs[3685]) | (layer0_outputs[4020]);
    assign outputs[4423] = (layer0_outputs[2989]) | (layer0_outputs[1370]);
    assign outputs[4424] = layer0_outputs[3279];
    assign outputs[4425] = (layer0_outputs[760]) ^ (layer0_outputs[6794]);
    assign outputs[4426] = (layer0_outputs[7673]) & ~(layer0_outputs[5976]);
    assign outputs[4427] = (layer0_outputs[3609]) & (layer0_outputs[3757]);
    assign outputs[4428] = ~(layer0_outputs[5796]);
    assign outputs[4429] = ~(layer0_outputs[7437]);
    assign outputs[4430] = ~(layer0_outputs[4521]);
    assign outputs[4431] = ~(layer0_outputs[4754]) | (layer0_outputs[25]);
    assign outputs[4432] = (layer0_outputs[127]) | (layer0_outputs[4746]);
    assign outputs[4433] = layer0_outputs[2495];
    assign outputs[4434] = layer0_outputs[7284];
    assign outputs[4435] = layer0_outputs[2647];
    assign outputs[4436] = (layer0_outputs[1590]) | (layer0_outputs[1860]);
    assign outputs[4437] = ~((layer0_outputs[2636]) & (layer0_outputs[1444]));
    assign outputs[4438] = ~(layer0_outputs[5067]) | (layer0_outputs[3568]);
    assign outputs[4439] = (layer0_outputs[4896]) ^ (layer0_outputs[4549]);
    assign outputs[4440] = ~(layer0_outputs[4549]);
    assign outputs[4441] = (layer0_outputs[6609]) ^ (layer0_outputs[970]);
    assign outputs[4442] = ~((layer0_outputs[5506]) ^ (layer0_outputs[3923]));
    assign outputs[4443] = layer0_outputs[1110];
    assign outputs[4444] = 1'b1;
    assign outputs[4445] = ~((layer0_outputs[7015]) | (layer0_outputs[279]));
    assign outputs[4446] = ~((layer0_outputs[5094]) | (layer0_outputs[1934]));
    assign outputs[4447] = ~(layer0_outputs[5711]);
    assign outputs[4448] = ~(layer0_outputs[1336]) | (layer0_outputs[783]);
    assign outputs[4449] = layer0_outputs[2914];
    assign outputs[4450] = ~(layer0_outputs[1753]);
    assign outputs[4451] = (layer0_outputs[4276]) & ~(layer0_outputs[7493]);
    assign outputs[4452] = ~((layer0_outputs[3006]) ^ (layer0_outputs[4940]));
    assign outputs[4453] = ~(layer0_outputs[6185]);
    assign outputs[4454] = ~((layer0_outputs[1968]) ^ (layer0_outputs[4000]));
    assign outputs[4455] = ~(layer0_outputs[7106]);
    assign outputs[4456] = ~((layer0_outputs[6785]) ^ (layer0_outputs[650]));
    assign outputs[4457] = ~((layer0_outputs[5707]) ^ (layer0_outputs[2648]));
    assign outputs[4458] = ~(layer0_outputs[129]);
    assign outputs[4459] = ~(layer0_outputs[6740]) | (layer0_outputs[7160]);
    assign outputs[4460] = (layer0_outputs[2534]) & ~(layer0_outputs[5529]);
    assign outputs[4461] = ~(layer0_outputs[2554]);
    assign outputs[4462] = ~((layer0_outputs[2267]) ^ (layer0_outputs[4019]));
    assign outputs[4463] = ~(layer0_outputs[7174]);
    assign outputs[4464] = ~(layer0_outputs[7040]);
    assign outputs[4465] = ~(layer0_outputs[1741]);
    assign outputs[4466] = (layer0_outputs[7118]) ^ (layer0_outputs[951]);
    assign outputs[4467] = ~(layer0_outputs[2212]);
    assign outputs[4468] = ~((layer0_outputs[1255]) ^ (layer0_outputs[1038]));
    assign outputs[4469] = ~(layer0_outputs[1403]) | (layer0_outputs[2925]);
    assign outputs[4470] = ~(layer0_outputs[5166]);
    assign outputs[4471] = ~(layer0_outputs[297]);
    assign outputs[4472] = (layer0_outputs[5623]) & ~(layer0_outputs[2969]);
    assign outputs[4473] = ~((layer0_outputs[3415]) ^ (layer0_outputs[4]));
    assign outputs[4474] = layer0_outputs[4933];
    assign outputs[4475] = ~(layer0_outputs[4917]);
    assign outputs[4476] = ~(layer0_outputs[4741]) | (layer0_outputs[3720]);
    assign outputs[4477] = ~(layer0_outputs[639]);
    assign outputs[4478] = ~(layer0_outputs[3505]);
    assign outputs[4479] = (layer0_outputs[2663]) ^ (layer0_outputs[2410]);
    assign outputs[4480] = layer0_outputs[2973];
    assign outputs[4481] = ~(layer0_outputs[6098]);
    assign outputs[4482] = layer0_outputs[2355];
    assign outputs[4483] = layer0_outputs[5609];
    assign outputs[4484] = (layer0_outputs[3776]) ^ (layer0_outputs[597]);
    assign outputs[4485] = ~(layer0_outputs[1098]);
    assign outputs[4486] = (layer0_outputs[3587]) & ~(layer0_outputs[6341]);
    assign outputs[4487] = ~((layer0_outputs[6415]) ^ (layer0_outputs[3945]));
    assign outputs[4488] = ~(layer0_outputs[4310]);
    assign outputs[4489] = ~((layer0_outputs[2364]) ^ (layer0_outputs[5492]));
    assign outputs[4490] = (layer0_outputs[3645]) ^ (layer0_outputs[81]);
    assign outputs[4491] = ~((layer0_outputs[86]) ^ (layer0_outputs[2446]));
    assign outputs[4492] = (layer0_outputs[90]) & ~(layer0_outputs[4619]);
    assign outputs[4493] = layer0_outputs[54];
    assign outputs[4494] = ~(layer0_outputs[7324]);
    assign outputs[4495] = (layer0_outputs[3666]) ^ (layer0_outputs[3731]);
    assign outputs[4496] = layer0_outputs[1453];
    assign outputs[4497] = ~(layer0_outputs[4132]);
    assign outputs[4498] = ~(layer0_outputs[1822]);
    assign outputs[4499] = (layer0_outputs[531]) ^ (layer0_outputs[1586]);
    assign outputs[4500] = (layer0_outputs[5669]) ^ (layer0_outputs[1478]);
    assign outputs[4501] = ~((layer0_outputs[6741]) & (layer0_outputs[2710]));
    assign outputs[4502] = layer0_outputs[3386];
    assign outputs[4503] = ~(layer0_outputs[4375]) | (layer0_outputs[1146]);
    assign outputs[4504] = (layer0_outputs[7572]) & ~(layer0_outputs[101]);
    assign outputs[4505] = ~((layer0_outputs[5968]) ^ (layer0_outputs[5873]));
    assign outputs[4506] = ~((layer0_outputs[6855]) ^ (layer0_outputs[6072]));
    assign outputs[4507] = layer0_outputs[5663];
    assign outputs[4508] = (layer0_outputs[2195]) ^ (layer0_outputs[66]);
    assign outputs[4509] = ~(layer0_outputs[5210]);
    assign outputs[4510] = (layer0_outputs[6167]) ^ (layer0_outputs[4652]);
    assign outputs[4511] = ~(layer0_outputs[5461]) | (layer0_outputs[7235]);
    assign outputs[4512] = ~(layer0_outputs[1763]);
    assign outputs[4513] = (layer0_outputs[3910]) ^ (layer0_outputs[3067]);
    assign outputs[4514] = layer0_outputs[5342];
    assign outputs[4515] = (layer0_outputs[5168]) & ~(layer0_outputs[5827]);
    assign outputs[4516] = ~((layer0_outputs[5916]) ^ (layer0_outputs[1317]));
    assign outputs[4517] = layer0_outputs[2388];
    assign outputs[4518] = layer0_outputs[443];
    assign outputs[4519] = ~((layer0_outputs[2144]) ^ (layer0_outputs[7278]));
    assign outputs[4520] = ~(layer0_outputs[38]);
    assign outputs[4521] = layer0_outputs[2218];
    assign outputs[4522] = (layer0_outputs[503]) & ~(layer0_outputs[3543]);
    assign outputs[4523] = ~(layer0_outputs[2832]);
    assign outputs[4524] = ~((layer0_outputs[415]) ^ (layer0_outputs[5155]));
    assign outputs[4525] = (layer0_outputs[2794]) ^ (layer0_outputs[334]);
    assign outputs[4526] = (layer0_outputs[2868]) | (layer0_outputs[1764]);
    assign outputs[4527] = (layer0_outputs[4373]) ^ (layer0_outputs[4139]);
    assign outputs[4528] = (layer0_outputs[6344]) ^ (layer0_outputs[4820]);
    assign outputs[4529] = ~((layer0_outputs[7376]) ^ (layer0_outputs[3868]));
    assign outputs[4530] = (layer0_outputs[909]) ^ (layer0_outputs[2133]);
    assign outputs[4531] = ~((layer0_outputs[2529]) ^ (layer0_outputs[4136]));
    assign outputs[4532] = ~(layer0_outputs[7631]);
    assign outputs[4533] = layer0_outputs[4348];
    assign outputs[4534] = (layer0_outputs[6204]) ^ (layer0_outputs[6287]);
    assign outputs[4535] = ~(layer0_outputs[6418]);
    assign outputs[4536] = (layer0_outputs[3244]) ^ (layer0_outputs[5114]);
    assign outputs[4537] = layer0_outputs[1755];
    assign outputs[4538] = (layer0_outputs[1308]) | (layer0_outputs[2870]);
    assign outputs[4539] = (layer0_outputs[5950]) ^ (layer0_outputs[7143]);
    assign outputs[4540] = (layer0_outputs[7036]) & ~(layer0_outputs[5794]);
    assign outputs[4541] = (layer0_outputs[7063]) ^ (layer0_outputs[5497]);
    assign outputs[4542] = ~(layer0_outputs[6375]) | (layer0_outputs[2208]);
    assign outputs[4543] = ~((layer0_outputs[7592]) | (layer0_outputs[5025]));
    assign outputs[4544] = ~((layer0_outputs[6660]) & (layer0_outputs[604]));
    assign outputs[4545] = ~((layer0_outputs[1009]) & (layer0_outputs[4211]));
    assign outputs[4546] = ~((layer0_outputs[5656]) ^ (layer0_outputs[2269]));
    assign outputs[4547] = (layer0_outputs[4407]) & (layer0_outputs[5316]);
    assign outputs[4548] = ~((layer0_outputs[6253]) & (layer0_outputs[1170]));
    assign outputs[4549] = ~(layer0_outputs[5690]);
    assign outputs[4550] = layer0_outputs[1290];
    assign outputs[4551] = ~(layer0_outputs[5015]) | (layer0_outputs[7000]);
    assign outputs[4552] = ~(layer0_outputs[6932]);
    assign outputs[4553] = ~(layer0_outputs[7402]);
    assign outputs[4554] = layer0_outputs[2675];
    assign outputs[4555] = layer0_outputs[2236];
    assign outputs[4556] = layer0_outputs[4962];
    assign outputs[4557] = (layer0_outputs[312]) ^ (layer0_outputs[5555]);
    assign outputs[4558] = (layer0_outputs[2050]) ^ (layer0_outputs[4269]);
    assign outputs[4559] = ~((layer0_outputs[3326]) ^ (layer0_outputs[6429]));
    assign outputs[4560] = layer0_outputs[6051];
    assign outputs[4561] = (layer0_outputs[607]) & ~(layer0_outputs[1687]);
    assign outputs[4562] = ~(layer0_outputs[1488]);
    assign outputs[4563] = (layer0_outputs[5379]) ^ (layer0_outputs[531]);
    assign outputs[4564] = ~((layer0_outputs[2483]) & (layer0_outputs[2898]));
    assign outputs[4565] = layer0_outputs[6434];
    assign outputs[4566] = ~((layer0_outputs[4300]) ^ (layer0_outputs[5312]));
    assign outputs[4567] = (layer0_outputs[3750]) ^ (layer0_outputs[5070]);
    assign outputs[4568] = (layer0_outputs[6797]) ^ (layer0_outputs[588]);
    assign outputs[4569] = (layer0_outputs[2954]) & (layer0_outputs[877]);
    assign outputs[4570] = ~((layer0_outputs[2081]) ^ (layer0_outputs[6832]));
    assign outputs[4571] = ~(layer0_outputs[3485]) | (layer0_outputs[4490]);
    assign outputs[4572] = layer0_outputs[3070];
    assign outputs[4573] = (layer0_outputs[2314]) & (layer0_outputs[6513]);
    assign outputs[4574] = (layer0_outputs[1846]) & (layer0_outputs[4437]);
    assign outputs[4575] = ~(layer0_outputs[4141]);
    assign outputs[4576] = (layer0_outputs[5499]) ^ (layer0_outputs[3673]);
    assign outputs[4577] = (layer0_outputs[4563]) & ~(layer0_outputs[2574]);
    assign outputs[4578] = (layer0_outputs[508]) & ~(layer0_outputs[4885]);
    assign outputs[4579] = ~(layer0_outputs[7515]);
    assign outputs[4580] = ~(layer0_outputs[2403]);
    assign outputs[4581] = (layer0_outputs[2817]) | (layer0_outputs[547]);
    assign outputs[4582] = ~((layer0_outputs[4108]) ^ (layer0_outputs[1813]));
    assign outputs[4583] = layer0_outputs[3453];
    assign outputs[4584] = ~((layer0_outputs[5605]) ^ (layer0_outputs[801]));
    assign outputs[4585] = (layer0_outputs[5901]) & (layer0_outputs[3767]);
    assign outputs[4586] = ~(layer0_outputs[6251]);
    assign outputs[4587] = ~(layer0_outputs[784]) | (layer0_outputs[1791]);
    assign outputs[4588] = layer0_outputs[4965];
    assign outputs[4589] = ~((layer0_outputs[691]) ^ (layer0_outputs[5354]));
    assign outputs[4590] = ~((layer0_outputs[1016]) | (layer0_outputs[5791]));
    assign outputs[4591] = ~(layer0_outputs[7008]);
    assign outputs[4592] = ~(layer0_outputs[1648]) | (layer0_outputs[5663]);
    assign outputs[4593] = (layer0_outputs[474]) ^ (layer0_outputs[6608]);
    assign outputs[4594] = layer0_outputs[4138];
    assign outputs[4595] = ~(layer0_outputs[2633]);
    assign outputs[4596] = ~((layer0_outputs[7150]) ^ (layer0_outputs[2386]));
    assign outputs[4597] = ~(layer0_outputs[725]);
    assign outputs[4598] = ~(layer0_outputs[865]) | (layer0_outputs[4052]);
    assign outputs[4599] = ~(layer0_outputs[7357]) | (layer0_outputs[516]);
    assign outputs[4600] = layer0_outputs[3419];
    assign outputs[4601] = (layer0_outputs[7568]) & (layer0_outputs[1926]);
    assign outputs[4602] = (layer0_outputs[5763]) ^ (layer0_outputs[6943]);
    assign outputs[4603] = (layer0_outputs[1076]) & ~(layer0_outputs[1751]);
    assign outputs[4604] = (layer0_outputs[388]) & ~(layer0_outputs[5484]);
    assign outputs[4605] = ~(layer0_outputs[2515]);
    assign outputs[4606] = ~((layer0_outputs[4326]) ^ (layer0_outputs[6759]));
    assign outputs[4607] = layer0_outputs[3917];
    assign outputs[4608] = ~(layer0_outputs[1048]);
    assign outputs[4609] = (layer0_outputs[811]) & (layer0_outputs[2952]);
    assign outputs[4610] = layer0_outputs[4337];
    assign outputs[4611] = ~(layer0_outputs[5669]);
    assign outputs[4612] = ~(layer0_outputs[6036]) | (layer0_outputs[6064]);
    assign outputs[4613] = (layer0_outputs[1233]) | (layer0_outputs[895]);
    assign outputs[4614] = ~((layer0_outputs[7574]) ^ (layer0_outputs[7540]));
    assign outputs[4615] = (layer0_outputs[6834]) & ~(layer0_outputs[4882]);
    assign outputs[4616] = (layer0_outputs[3274]) ^ (layer0_outputs[646]);
    assign outputs[4617] = (layer0_outputs[6019]) ^ (layer0_outputs[1099]);
    assign outputs[4618] = (layer0_outputs[43]) ^ (layer0_outputs[5930]);
    assign outputs[4619] = ~((layer0_outputs[6949]) ^ (layer0_outputs[4967]));
    assign outputs[4620] = (layer0_outputs[4672]) & (layer0_outputs[1577]);
    assign outputs[4621] = ~((layer0_outputs[2325]) & (layer0_outputs[905]));
    assign outputs[4622] = ~(layer0_outputs[6652]) | (layer0_outputs[1737]);
    assign outputs[4623] = layer0_outputs[3328];
    assign outputs[4624] = layer0_outputs[2812];
    assign outputs[4625] = 1'b1;
    assign outputs[4626] = (layer0_outputs[4101]) & ~(layer0_outputs[3186]);
    assign outputs[4627] = ~(layer0_outputs[3654]);
    assign outputs[4628] = layer0_outputs[3064];
    assign outputs[4629] = layer0_outputs[2324];
    assign outputs[4630] = ~(layer0_outputs[7306]);
    assign outputs[4631] = ~(layer0_outputs[2287]);
    assign outputs[4632] = ~(layer0_outputs[2474]);
    assign outputs[4633] = layer0_outputs[4664];
    assign outputs[4634] = ~(layer0_outputs[4396]);
    assign outputs[4635] = ~(layer0_outputs[2145]) | (layer0_outputs[2941]);
    assign outputs[4636] = layer0_outputs[5910];
    assign outputs[4637] = ~(layer0_outputs[2653]);
    assign outputs[4638] = ~((layer0_outputs[1704]) & (layer0_outputs[671]));
    assign outputs[4639] = (layer0_outputs[134]) & ~(layer0_outputs[182]);
    assign outputs[4640] = layer0_outputs[3659];
    assign outputs[4641] = ~(layer0_outputs[6814]);
    assign outputs[4642] = ~(layer0_outputs[3912]);
    assign outputs[4643] = ~(layer0_outputs[2957]);
    assign outputs[4644] = (layer0_outputs[7195]) | (layer0_outputs[3561]);
    assign outputs[4645] = ~(layer0_outputs[2771]);
    assign outputs[4646] = (layer0_outputs[2430]) ^ (layer0_outputs[1746]);
    assign outputs[4647] = ~(layer0_outputs[730]);
    assign outputs[4648] = (layer0_outputs[872]) & (layer0_outputs[5253]);
    assign outputs[4649] = (layer0_outputs[5473]) & ~(layer0_outputs[1054]);
    assign outputs[4650] = ~(layer0_outputs[3706]);
    assign outputs[4651] = ~((layer0_outputs[6630]) | (layer0_outputs[2999]));
    assign outputs[4652] = (layer0_outputs[2639]) ^ (layer0_outputs[2078]);
    assign outputs[4653] = (layer0_outputs[5310]) & ~(layer0_outputs[855]);
    assign outputs[4654] = layer0_outputs[5824];
    assign outputs[4655] = layer0_outputs[6653];
    assign outputs[4656] = ~(layer0_outputs[1093]);
    assign outputs[4657] = ~(layer0_outputs[2143]);
    assign outputs[4658] = layer0_outputs[5851];
    assign outputs[4659] = (layer0_outputs[1522]) & ~(layer0_outputs[174]);
    assign outputs[4660] = ~(layer0_outputs[4281]);
    assign outputs[4661] = layer0_outputs[7375];
    assign outputs[4662] = ~(layer0_outputs[2489]);
    assign outputs[4663] = (layer0_outputs[7613]) ^ (layer0_outputs[766]);
    assign outputs[4664] = (layer0_outputs[1144]) ^ (layer0_outputs[2530]);
    assign outputs[4665] = (layer0_outputs[7299]) & (layer0_outputs[6565]);
    assign outputs[4666] = layer0_outputs[1008];
    assign outputs[4667] = (layer0_outputs[2542]) & ~(layer0_outputs[5757]);
    assign outputs[4668] = ~(layer0_outputs[2561]);
    assign outputs[4669] = layer0_outputs[347];
    assign outputs[4670] = layer0_outputs[7431];
    assign outputs[4671] = ~(layer0_outputs[5866]);
    assign outputs[4672] = ~(layer0_outputs[7244]);
    assign outputs[4673] = ~((layer0_outputs[3601]) ^ (layer0_outputs[7223]));
    assign outputs[4674] = ~(layer0_outputs[504]);
    assign outputs[4675] = (layer0_outputs[5735]) | (layer0_outputs[3068]);
    assign outputs[4676] = ~((layer0_outputs[394]) | (layer0_outputs[1471]));
    assign outputs[4677] = ~(layer0_outputs[4272]);
    assign outputs[4678] = ~((layer0_outputs[5192]) & (layer0_outputs[1397]));
    assign outputs[4679] = ~((layer0_outputs[258]) & (layer0_outputs[2905]));
    assign outputs[4680] = ~((layer0_outputs[1928]) ^ (layer0_outputs[4406]));
    assign outputs[4681] = layer0_outputs[17];
    assign outputs[4682] = (layer0_outputs[1825]) & (layer0_outputs[1594]);
    assign outputs[4683] = (layer0_outputs[6338]) | (layer0_outputs[6281]);
    assign outputs[4684] = (layer0_outputs[2628]) & ~(layer0_outputs[6440]);
    assign outputs[4685] = ~(layer0_outputs[853]);
    assign outputs[4686] = (layer0_outputs[3919]) & ~(layer0_outputs[7392]);
    assign outputs[4687] = layer0_outputs[6558];
    assign outputs[4688] = ~((layer0_outputs[3283]) & (layer0_outputs[1604]));
    assign outputs[4689] = layer0_outputs[1595];
    assign outputs[4690] = (layer0_outputs[4322]) & ~(layer0_outputs[1503]);
    assign outputs[4691] = (layer0_outputs[3141]) & ~(layer0_outputs[4793]);
    assign outputs[4692] = (layer0_outputs[4642]) ^ (layer0_outputs[6750]);
    assign outputs[4693] = (layer0_outputs[4853]) ^ (layer0_outputs[5903]);
    assign outputs[4694] = ~((layer0_outputs[4761]) & (layer0_outputs[6365]));
    assign outputs[4695] = (layer0_outputs[474]) & (layer0_outputs[7282]);
    assign outputs[4696] = (layer0_outputs[700]) | (layer0_outputs[2778]);
    assign outputs[4697] = layer0_outputs[6481];
    assign outputs[4698] = ~((layer0_outputs[6022]) | (layer0_outputs[4780]));
    assign outputs[4699] = ~((layer0_outputs[4850]) & (layer0_outputs[6466]));
    assign outputs[4700] = ~((layer0_outputs[5512]) ^ (layer0_outputs[674]));
    assign outputs[4701] = layer0_outputs[653];
    assign outputs[4702] = ~((layer0_outputs[2047]) | (layer0_outputs[1608]));
    assign outputs[4703] = ~((layer0_outputs[5437]) ^ (layer0_outputs[2181]));
    assign outputs[4704] = layer0_outputs[4409];
    assign outputs[4705] = ~(layer0_outputs[894]);
    assign outputs[4706] = layer0_outputs[5389];
    assign outputs[4707] = layer0_outputs[7155];
    assign outputs[4708] = ~(layer0_outputs[6332]);
    assign outputs[4709] = ~((layer0_outputs[1800]) | (layer0_outputs[5327]));
    assign outputs[4710] = layer0_outputs[239];
    assign outputs[4711] = layer0_outputs[794];
    assign outputs[4712] = layer0_outputs[5910];
    assign outputs[4713] = ~((layer0_outputs[2768]) ^ (layer0_outputs[6656]));
    assign outputs[4714] = (layer0_outputs[4310]) ^ (layer0_outputs[5159]);
    assign outputs[4715] = (layer0_outputs[7628]) & ~(layer0_outputs[5016]);
    assign outputs[4716] = 1'b1;
    assign outputs[4717] = layer0_outputs[1062];
    assign outputs[4718] = ~(layer0_outputs[5278]);
    assign outputs[4719] = ~(layer0_outputs[3681]);
    assign outputs[4720] = (layer0_outputs[593]) & ~(layer0_outputs[7144]);
    assign outputs[4721] = ~(layer0_outputs[1830]);
    assign outputs[4722] = (layer0_outputs[6021]) & ~(layer0_outputs[143]);
    assign outputs[4723] = (layer0_outputs[4150]) & ~(layer0_outputs[1271]);
    assign outputs[4724] = ~(layer0_outputs[6294]) | (layer0_outputs[6619]);
    assign outputs[4725] = (layer0_outputs[2827]) ^ (layer0_outputs[5734]);
    assign outputs[4726] = ~(layer0_outputs[3324]) | (layer0_outputs[568]);
    assign outputs[4727] = ~((layer0_outputs[2203]) ^ (layer0_outputs[1176]));
    assign outputs[4728] = (layer0_outputs[1607]) ^ (layer0_outputs[6924]);
    assign outputs[4729] = (layer0_outputs[1524]) & (layer0_outputs[6571]);
    assign outputs[4730] = layer0_outputs[2539];
    assign outputs[4731] = ~(layer0_outputs[5623]);
    assign outputs[4732] = ~((layer0_outputs[3480]) | (layer0_outputs[7281]));
    assign outputs[4733] = ~((layer0_outputs[7241]) | (layer0_outputs[5188]));
    assign outputs[4734] = ~(layer0_outputs[5394]);
    assign outputs[4735] = ~(layer0_outputs[2550]);
    assign outputs[4736] = ~(layer0_outputs[6136]);
    assign outputs[4737] = (layer0_outputs[1289]) ^ (layer0_outputs[5288]);
    assign outputs[4738] = ~(layer0_outputs[2833]);
    assign outputs[4739] = layer0_outputs[4277];
    assign outputs[4740] = (layer0_outputs[1094]) & ~(layer0_outputs[70]);
    assign outputs[4741] = ~((layer0_outputs[6501]) ^ (layer0_outputs[2639]));
    assign outputs[4742] = layer0_outputs[613];
    assign outputs[4743] = ~(layer0_outputs[6709]);
    assign outputs[4744] = ~(layer0_outputs[552]);
    assign outputs[4745] = layer0_outputs[2180];
    assign outputs[4746] = ~(layer0_outputs[815]);
    assign outputs[4747] = ~(layer0_outputs[2871]) | (layer0_outputs[3939]);
    assign outputs[4748] = ~(layer0_outputs[5225]);
    assign outputs[4749] = ~((layer0_outputs[2273]) ^ (layer0_outputs[6306]));
    assign outputs[4750] = (layer0_outputs[2907]) & ~(layer0_outputs[331]);
    assign outputs[4751] = ~(layer0_outputs[3589]) | (layer0_outputs[1203]);
    assign outputs[4752] = (layer0_outputs[5446]) | (layer0_outputs[4142]);
    assign outputs[4753] = (layer0_outputs[3484]) & (layer0_outputs[7016]);
    assign outputs[4754] = (layer0_outputs[4151]) & ~(layer0_outputs[4770]);
    assign outputs[4755] = layer0_outputs[3961];
    assign outputs[4756] = ~(layer0_outputs[3991]);
    assign outputs[4757] = ~(layer0_outputs[6316]) | (layer0_outputs[5229]);
    assign outputs[4758] = (layer0_outputs[152]) & (layer0_outputs[4526]);
    assign outputs[4759] = ~(layer0_outputs[3540]) | (layer0_outputs[5072]);
    assign outputs[4760] = (layer0_outputs[4915]) ^ (layer0_outputs[2414]);
    assign outputs[4761] = (layer0_outputs[1825]) & ~(layer0_outputs[5833]);
    assign outputs[4762] = (layer0_outputs[5737]) & ~(layer0_outputs[1160]);
    assign outputs[4763] = ~(layer0_outputs[878]);
    assign outputs[4764] = ~((layer0_outputs[351]) | (layer0_outputs[6944]));
    assign outputs[4765] = ~(layer0_outputs[2032]);
    assign outputs[4766] = ~(layer0_outputs[1627]) | (layer0_outputs[6352]);
    assign outputs[4767] = ~((layer0_outputs[6874]) ^ (layer0_outputs[2142]));
    assign outputs[4768] = (layer0_outputs[5282]) ^ (layer0_outputs[1253]);
    assign outputs[4769] = ~(layer0_outputs[2062]);
    assign outputs[4770] = ~((layer0_outputs[3905]) & (layer0_outputs[4786]));
    assign outputs[4771] = ~(layer0_outputs[4403]) | (layer0_outputs[1990]);
    assign outputs[4772] = ~((layer0_outputs[6542]) | (layer0_outputs[6713]));
    assign outputs[4773] = (layer0_outputs[413]) ^ (layer0_outputs[160]);
    assign outputs[4774] = (layer0_outputs[7348]) | (layer0_outputs[2822]);
    assign outputs[4775] = ~(layer0_outputs[3525]);
    assign outputs[4776] = layer0_outputs[3650];
    assign outputs[4777] = (layer0_outputs[1938]) ^ (layer0_outputs[1974]);
    assign outputs[4778] = layer0_outputs[5688];
    assign outputs[4779] = (layer0_outputs[4143]) & ~(layer0_outputs[7292]);
    assign outputs[4780] = (layer0_outputs[5597]) & ~(layer0_outputs[4919]);
    assign outputs[4781] = ~((layer0_outputs[6160]) ^ (layer0_outputs[5510]));
    assign outputs[4782] = ~((layer0_outputs[394]) | (layer0_outputs[6800]));
    assign outputs[4783] = ~(layer0_outputs[2018]);
    assign outputs[4784] = ~((layer0_outputs[5511]) ^ (layer0_outputs[5777]));
    assign outputs[4785] = ~((layer0_outputs[1340]) | (layer0_outputs[4165]));
    assign outputs[4786] = ~(layer0_outputs[3513]);
    assign outputs[4787] = ~((layer0_outputs[4793]) ^ (layer0_outputs[2615]));
    assign outputs[4788] = ~((layer0_outputs[3635]) ^ (layer0_outputs[618]));
    assign outputs[4789] = ~(layer0_outputs[2723]);
    assign outputs[4790] = ~(layer0_outputs[305]);
    assign outputs[4791] = ~(layer0_outputs[5193]);
    assign outputs[4792] = layer0_outputs[281];
    assign outputs[4793] = layer0_outputs[5558];
    assign outputs[4794] = layer0_outputs[7039];
    assign outputs[4795] = ~(layer0_outputs[1292]);
    assign outputs[4796] = ~((layer0_outputs[7326]) | (layer0_outputs[166]));
    assign outputs[4797] = ~(layer0_outputs[3085]);
    assign outputs[4798] = layer0_outputs[5383];
    assign outputs[4799] = ~(layer0_outputs[923]);
    assign outputs[4800] = ~((layer0_outputs[4570]) & (layer0_outputs[4060]));
    assign outputs[4801] = ~(layer0_outputs[7645]) | (layer0_outputs[120]);
    assign outputs[4802] = ~(layer0_outputs[160]);
    assign outputs[4803] = ~(layer0_outputs[3892]);
    assign outputs[4804] = ~((layer0_outputs[1784]) ^ (layer0_outputs[3651]));
    assign outputs[4805] = (layer0_outputs[6777]) & ~(layer0_outputs[4445]);
    assign outputs[4806] = ~(layer0_outputs[6125]);
    assign outputs[4807] = ~(layer0_outputs[247]) | (layer0_outputs[5047]);
    assign outputs[4808] = ~((layer0_outputs[403]) ^ (layer0_outputs[3633]));
    assign outputs[4809] = (layer0_outputs[1577]) & (layer0_outputs[421]);
    assign outputs[4810] = ~(layer0_outputs[1790]);
    assign outputs[4811] = layer0_outputs[1592];
    assign outputs[4812] = layer0_outputs[6459];
    assign outputs[4813] = ~(layer0_outputs[5907]) | (layer0_outputs[6715]);
    assign outputs[4814] = ~(layer0_outputs[6163]);
    assign outputs[4815] = ~(layer0_outputs[3429]);
    assign outputs[4816] = ~(layer0_outputs[4935]) | (layer0_outputs[4406]);
    assign outputs[4817] = layer0_outputs[1300];
    assign outputs[4818] = layer0_outputs[3078];
    assign outputs[4819] = ~((layer0_outputs[6720]) | (layer0_outputs[5747]));
    assign outputs[4820] = layer0_outputs[6029];
    assign outputs[4821] = (layer0_outputs[1895]) & ~(layer0_outputs[7477]);
    assign outputs[4822] = ~(layer0_outputs[7119]);
    assign outputs[4823] = ~(layer0_outputs[2506]) | (layer0_outputs[2933]);
    assign outputs[4824] = layer0_outputs[5304];
    assign outputs[4825] = layer0_outputs[7641];
    assign outputs[4826] = (layer0_outputs[3275]) ^ (layer0_outputs[4372]);
    assign outputs[4827] = ~((layer0_outputs[4418]) ^ (layer0_outputs[1982]));
    assign outputs[4828] = layer0_outputs[7616];
    assign outputs[4829] = ~((layer0_outputs[4881]) ^ (layer0_outputs[5459]));
    assign outputs[4830] = ~((layer0_outputs[6976]) ^ (layer0_outputs[3287]));
    assign outputs[4831] = ~((layer0_outputs[3901]) | (layer0_outputs[3686]));
    assign outputs[4832] = (layer0_outputs[1853]) ^ (layer0_outputs[1163]);
    assign outputs[4833] = ~(layer0_outputs[7516]);
    assign outputs[4834] = ~(layer0_outputs[5717]) | (layer0_outputs[4623]);
    assign outputs[4835] = layer0_outputs[5881];
    assign outputs[4836] = ~(layer0_outputs[3108]);
    assign outputs[4837] = ~((layer0_outputs[1960]) ^ (layer0_outputs[2822]));
    assign outputs[4838] = layer0_outputs[2846];
    assign outputs[4839] = (layer0_outputs[4667]) & ~(layer0_outputs[7524]);
    assign outputs[4840] = ~(layer0_outputs[3938]);
    assign outputs[4841] = ~(layer0_outputs[4716]) | (layer0_outputs[2414]);
    assign outputs[4842] = ~(layer0_outputs[7033]);
    assign outputs[4843] = ~(layer0_outputs[3190]);
    assign outputs[4844] = ~((layer0_outputs[147]) | (layer0_outputs[6897]));
    assign outputs[4845] = ~(layer0_outputs[5643]);
    assign outputs[4846] = layer0_outputs[1580];
    assign outputs[4847] = layer0_outputs[342];
    assign outputs[4848] = ~((layer0_outputs[1032]) | (layer0_outputs[3028]));
    assign outputs[4849] = (layer0_outputs[1285]) & (layer0_outputs[2435]);
    assign outputs[4850] = layer0_outputs[1721];
    assign outputs[4851] = layer0_outputs[2139];
    assign outputs[4852] = ~((layer0_outputs[3813]) & (layer0_outputs[6016]));
    assign outputs[4853] = ~(layer0_outputs[7408]);
    assign outputs[4854] = ~((layer0_outputs[4969]) ^ (layer0_outputs[3232]));
    assign outputs[4855] = layer0_outputs[1832];
    assign outputs[4856] = ~((layer0_outputs[268]) & (layer0_outputs[1988]));
    assign outputs[4857] = (layer0_outputs[4658]) ^ (layer0_outputs[2570]);
    assign outputs[4858] = ~(layer0_outputs[7459]);
    assign outputs[4859] = ~((layer0_outputs[6706]) & (layer0_outputs[4673]));
    assign outputs[4860] = layer0_outputs[4116];
    assign outputs[4861] = (layer0_outputs[684]) | (layer0_outputs[7372]);
    assign outputs[4862] = (layer0_outputs[7609]) & (layer0_outputs[6655]);
    assign outputs[4863] = ~((layer0_outputs[3760]) ^ (layer0_outputs[2985]));
    assign outputs[4864] = (layer0_outputs[4103]) & (layer0_outputs[6877]);
    assign outputs[4865] = ~((layer0_outputs[4898]) ^ (layer0_outputs[3541]));
    assign outputs[4866] = ~((layer0_outputs[998]) | (layer0_outputs[3231]));
    assign outputs[4867] = (layer0_outputs[6674]) & ~(layer0_outputs[2494]);
    assign outputs[4868] = (layer0_outputs[2915]) & ~(layer0_outputs[3334]);
    assign outputs[4869] = layer0_outputs[7162];
    assign outputs[4870] = ~((layer0_outputs[4315]) ^ (layer0_outputs[1118]));
    assign outputs[4871] = layer0_outputs[6681];
    assign outputs[4872] = (layer0_outputs[2623]) | (layer0_outputs[4111]);
    assign outputs[4873] = (layer0_outputs[380]) ^ (layer0_outputs[7568]);
    assign outputs[4874] = (layer0_outputs[6122]) | (layer0_outputs[2086]);
    assign outputs[4875] = ~(layer0_outputs[6431]);
    assign outputs[4876] = ~((layer0_outputs[795]) ^ (layer0_outputs[4864]));
    assign outputs[4877] = ~((layer0_outputs[542]) ^ (layer0_outputs[4621]));
    assign outputs[4878] = layer0_outputs[7338];
    assign outputs[4879] = ~(layer0_outputs[6633]);
    assign outputs[4880] = layer0_outputs[6555];
    assign outputs[4881] = layer0_outputs[79];
    assign outputs[4882] = (layer0_outputs[1654]) & (layer0_outputs[2956]);
    assign outputs[4883] = (layer0_outputs[2122]) & (layer0_outputs[1445]);
    assign outputs[4884] = ~(layer0_outputs[6903]);
    assign outputs[4885] = (layer0_outputs[6776]) | (layer0_outputs[6506]);
    assign outputs[4886] = ~(layer0_outputs[1534]);
    assign outputs[4887] = (layer0_outputs[7433]) ^ (layer0_outputs[5562]);
    assign outputs[4888] = (layer0_outputs[2654]) & ~(layer0_outputs[3709]);
    assign outputs[4889] = ~(layer0_outputs[4312]) | (layer0_outputs[6183]);
    assign outputs[4890] = ~((layer0_outputs[5352]) ^ (layer0_outputs[7555]));
    assign outputs[4891] = layer0_outputs[5695];
    assign outputs[4892] = ~((layer0_outputs[1254]) & (layer0_outputs[123]));
    assign outputs[4893] = ~((layer0_outputs[6250]) ^ (layer0_outputs[5229]));
    assign outputs[4894] = ~((layer0_outputs[2017]) | (layer0_outputs[1664]));
    assign outputs[4895] = ~((layer0_outputs[6647]) ^ (layer0_outputs[5167]));
    assign outputs[4896] = ~(layer0_outputs[2374]);
    assign outputs[4897] = (layer0_outputs[2354]) & (layer0_outputs[53]);
    assign outputs[4898] = ~(layer0_outputs[3850]);
    assign outputs[4899] = layer0_outputs[3065];
    assign outputs[4900] = (layer0_outputs[6992]) ^ (layer0_outputs[1371]);
    assign outputs[4901] = layer0_outputs[3692];
    assign outputs[4902] = layer0_outputs[4022];
    assign outputs[4903] = ~((layer0_outputs[1762]) ^ (layer0_outputs[3410]));
    assign outputs[4904] = ~(layer0_outputs[319]);
    assign outputs[4905] = (layer0_outputs[7399]) | (layer0_outputs[2530]);
    assign outputs[4906] = ~(layer0_outputs[5649]) | (layer0_outputs[872]);
    assign outputs[4907] = (layer0_outputs[6544]) & (layer0_outputs[2581]);
    assign outputs[4908] = ~((layer0_outputs[5041]) ^ (layer0_outputs[6769]));
    assign outputs[4909] = ~(layer0_outputs[5797]) | (layer0_outputs[5547]);
    assign outputs[4910] = ~(layer0_outputs[2160]);
    assign outputs[4911] = layer0_outputs[6249];
    assign outputs[4912] = ~((layer0_outputs[1509]) ^ (layer0_outputs[2266]));
    assign outputs[4913] = (layer0_outputs[1713]) | (layer0_outputs[3466]);
    assign outputs[4914] = (layer0_outputs[6053]) & ~(layer0_outputs[7488]);
    assign outputs[4915] = ~((layer0_outputs[5508]) & (layer0_outputs[4594]));
    assign outputs[4916] = ~(layer0_outputs[3752]) | (layer0_outputs[6656]);
    assign outputs[4917] = ~((layer0_outputs[3590]) ^ (layer0_outputs[3308]));
    assign outputs[4918] = ~(layer0_outputs[2718]);
    assign outputs[4919] = ~(layer0_outputs[3407]) | (layer0_outputs[5803]);
    assign outputs[4920] = layer0_outputs[4154];
    assign outputs[4921] = ~(layer0_outputs[5281]) | (layer0_outputs[619]);
    assign outputs[4922] = ~(layer0_outputs[992]);
    assign outputs[4923] = ~(layer0_outputs[1538]);
    assign outputs[4924] = layer0_outputs[4611];
    assign outputs[4925] = layer0_outputs[412];
    assign outputs[4926] = layer0_outputs[622];
    assign outputs[4927] = layer0_outputs[4238];
    assign outputs[4928] = ~((layer0_outputs[7301]) ^ (layer0_outputs[3383]));
    assign outputs[4929] = (layer0_outputs[5371]) & ~(layer0_outputs[2142]);
    assign outputs[4930] = ~(layer0_outputs[5653]);
    assign outputs[4931] = ~(layer0_outputs[1169]) | (layer0_outputs[1420]);
    assign outputs[4932] = layer0_outputs[6667];
    assign outputs[4933] = ~(layer0_outputs[6548]);
    assign outputs[4934] = layer0_outputs[6437];
    assign outputs[4935] = layer0_outputs[1861];
    assign outputs[4936] = ~((layer0_outputs[2950]) ^ (layer0_outputs[1084]));
    assign outputs[4937] = ~((layer0_outputs[1887]) & (layer0_outputs[7147]));
    assign outputs[4938] = ~((layer0_outputs[4784]) | (layer0_outputs[4102]));
    assign outputs[4939] = (layer0_outputs[6687]) ^ (layer0_outputs[3924]);
    assign outputs[4940] = layer0_outputs[4440];
    assign outputs[4941] = layer0_outputs[7448];
    assign outputs[4942] = layer0_outputs[1789];
    assign outputs[4943] = layer0_outputs[957];
    assign outputs[4944] = (layer0_outputs[4902]) ^ (layer0_outputs[3687]);
    assign outputs[4945] = ~(layer0_outputs[7597]);
    assign outputs[4946] = (layer0_outputs[211]) ^ (layer0_outputs[5421]);
    assign outputs[4947] = layer0_outputs[6062];
    assign outputs[4948] = (layer0_outputs[1995]) ^ (layer0_outputs[4290]);
    assign outputs[4949] = ~(layer0_outputs[6856]);
    assign outputs[4950] = layer0_outputs[7312];
    assign outputs[4951] = layer0_outputs[4113];
    assign outputs[4952] = ~((layer0_outputs[1673]) ^ (layer0_outputs[7075]));
    assign outputs[4953] = (layer0_outputs[336]) | (layer0_outputs[689]);
    assign outputs[4954] = ~((layer0_outputs[518]) & (layer0_outputs[5481]));
    assign outputs[4955] = ~((layer0_outputs[2916]) & (layer0_outputs[5183]));
    assign outputs[4956] = (layer0_outputs[1309]) & ~(layer0_outputs[4781]);
    assign outputs[4957] = ~((layer0_outputs[4040]) ^ (layer0_outputs[1765]));
    assign outputs[4958] = ~((layer0_outputs[672]) ^ (layer0_outputs[96]));
    assign outputs[4959] = ~(layer0_outputs[4683]);
    assign outputs[4960] = (layer0_outputs[7169]) | (layer0_outputs[5954]);
    assign outputs[4961] = (layer0_outputs[2024]) ^ (layer0_outputs[5645]);
    assign outputs[4962] = ~(layer0_outputs[5307]);
    assign outputs[4963] = (layer0_outputs[6089]) & (layer0_outputs[6554]);
    assign outputs[4964] = layer0_outputs[1157];
    assign outputs[4965] = layer0_outputs[7346];
    assign outputs[4966] = ~(layer0_outputs[356]);
    assign outputs[4967] = ~(layer0_outputs[4200]);
    assign outputs[4968] = (layer0_outputs[1460]) & ~(layer0_outputs[6769]);
    assign outputs[4969] = ~((layer0_outputs[2410]) & (layer0_outputs[1230]));
    assign outputs[4970] = (layer0_outputs[3208]) & (layer0_outputs[1896]);
    assign outputs[4971] = layer0_outputs[2031];
    assign outputs[4972] = ~(layer0_outputs[1986]);
    assign outputs[4973] = layer0_outputs[3063];
    assign outputs[4974] = layer0_outputs[4758];
    assign outputs[4975] = (layer0_outputs[4589]) ^ (layer0_outputs[4493]);
    assign outputs[4976] = layer0_outputs[4373];
    assign outputs[4977] = layer0_outputs[2405];
    assign outputs[4978] = ~((layer0_outputs[6460]) ^ (layer0_outputs[3021]));
    assign outputs[4979] = layer0_outputs[7179];
    assign outputs[4980] = (layer0_outputs[3774]) ^ (layer0_outputs[5231]);
    assign outputs[4981] = ~(layer0_outputs[6258]);
    assign outputs[4982] = ~((layer0_outputs[4757]) ^ (layer0_outputs[6996]));
    assign outputs[4983] = ~((layer0_outputs[2039]) | (layer0_outputs[2828]));
    assign outputs[4984] = ~(layer0_outputs[3608]);
    assign outputs[4985] = (layer0_outputs[6271]) ^ (layer0_outputs[1015]);
    assign outputs[4986] = layer0_outputs[3176];
    assign outputs[4987] = ~((layer0_outputs[5417]) | (layer0_outputs[4028]));
    assign outputs[4988] = layer0_outputs[2861];
    assign outputs[4989] = ~(layer0_outputs[3830]);
    assign outputs[4990] = layer0_outputs[213];
    assign outputs[4991] = ~(layer0_outputs[458]);
    assign outputs[4992] = (layer0_outputs[5558]) & ~(layer0_outputs[5299]);
    assign outputs[4993] = layer0_outputs[2038];
    assign outputs[4994] = layer0_outputs[7352];
    assign outputs[4995] = ~((layer0_outputs[6975]) & (layer0_outputs[1866]));
    assign outputs[4996] = ~((layer0_outputs[797]) ^ (layer0_outputs[2193]));
    assign outputs[4997] = ~(layer0_outputs[2001]);
    assign outputs[4998] = layer0_outputs[4278];
    assign outputs[4999] = (layer0_outputs[3647]) ^ (layer0_outputs[3387]);
    assign outputs[5000] = ~(layer0_outputs[971]);
    assign outputs[5001] = ~(layer0_outputs[5616]) | (layer0_outputs[3803]);
    assign outputs[5002] = (layer0_outputs[6841]) & ~(layer0_outputs[465]);
    assign outputs[5003] = layer0_outputs[4613];
    assign outputs[5004] = ~((layer0_outputs[4289]) | (layer0_outputs[1459]));
    assign outputs[5005] = (layer0_outputs[5033]) & ~(layer0_outputs[2736]);
    assign outputs[5006] = (layer0_outputs[2388]) & (layer0_outputs[7225]);
    assign outputs[5007] = ~(layer0_outputs[2550]);
    assign outputs[5008] = (layer0_outputs[7360]) ^ (layer0_outputs[6804]);
    assign outputs[5009] = (layer0_outputs[2877]) ^ (layer0_outputs[796]);
    assign outputs[5010] = ~(layer0_outputs[459]);
    assign outputs[5011] = ~((layer0_outputs[4138]) ^ (layer0_outputs[1115]));
    assign outputs[5012] = layer0_outputs[3824];
    assign outputs[5013] = layer0_outputs[7363];
    assign outputs[5014] = layer0_outputs[6206];
    assign outputs[5015] = ~(layer0_outputs[1403]) | (layer0_outputs[3902]);
    assign outputs[5016] = ~(layer0_outputs[7276]);
    assign outputs[5017] = layer0_outputs[4629];
    assign outputs[5018] = (layer0_outputs[3966]) ^ (layer0_outputs[3338]);
    assign outputs[5019] = ~(layer0_outputs[6096]);
    assign outputs[5020] = ~((layer0_outputs[3385]) | (layer0_outputs[4703]));
    assign outputs[5021] = (layer0_outputs[4974]) ^ (layer0_outputs[1787]);
    assign outputs[5022] = (layer0_outputs[5125]) & (layer0_outputs[2005]);
    assign outputs[5023] = layer0_outputs[5124];
    assign outputs[5024] = layer0_outputs[3849];
    assign outputs[5025] = layer0_outputs[4512];
    assign outputs[5026] = ~(layer0_outputs[3719]);
    assign outputs[5027] = ~(layer0_outputs[4575]);
    assign outputs[5028] = (layer0_outputs[7461]) & ~(layer0_outputs[3257]);
    assign outputs[5029] = ~(layer0_outputs[7590]);
    assign outputs[5030] = ~((layer0_outputs[4694]) | (layer0_outputs[5074]));
    assign outputs[5031] = (layer0_outputs[4359]) & ~(layer0_outputs[916]);
    assign outputs[5032] = ~(layer0_outputs[6900]);
    assign outputs[5033] = layer0_outputs[164];
    assign outputs[5034] = ~(layer0_outputs[2021]);
    assign outputs[5035] = ~(layer0_outputs[6211]);
    assign outputs[5036] = (layer0_outputs[1185]) ^ (layer0_outputs[1127]);
    assign outputs[5037] = ~((layer0_outputs[1127]) ^ (layer0_outputs[3112]));
    assign outputs[5038] = layer0_outputs[1791];
    assign outputs[5039] = layer0_outputs[6920];
    assign outputs[5040] = ~(layer0_outputs[3644]);
    assign outputs[5041] = layer0_outputs[6305];
    assign outputs[5042] = layer0_outputs[5949];
    assign outputs[5043] = ~((layer0_outputs[369]) ^ (layer0_outputs[660]));
    assign outputs[5044] = (layer0_outputs[822]) ^ (layer0_outputs[4623]);
    assign outputs[5045] = ~((layer0_outputs[4092]) | (layer0_outputs[3310]));
    assign outputs[5046] = layer0_outputs[1956];
    assign outputs[5047] = ~((layer0_outputs[7177]) ^ (layer0_outputs[6182]));
    assign outputs[5048] = layer0_outputs[3508];
    assign outputs[5049] = ~((layer0_outputs[5009]) | (layer0_outputs[157]));
    assign outputs[5050] = (layer0_outputs[6968]) & ~(layer0_outputs[2063]);
    assign outputs[5051] = ~(layer0_outputs[3162]);
    assign outputs[5052] = (layer0_outputs[5867]) & (layer0_outputs[817]);
    assign outputs[5053] = (layer0_outputs[5386]) ^ (layer0_outputs[6847]);
    assign outputs[5054] = ~(layer0_outputs[2754]) | (layer0_outputs[5502]);
    assign outputs[5055] = (layer0_outputs[3361]) ^ (layer0_outputs[5259]);
    assign outputs[5056] = ~((layer0_outputs[6004]) | (layer0_outputs[7503]));
    assign outputs[5057] = layer0_outputs[7463];
    assign outputs[5058] = ~(layer0_outputs[2349]);
    assign outputs[5059] = layer0_outputs[5357];
    assign outputs[5060] = ~((layer0_outputs[2061]) ^ (layer0_outputs[2274]));
    assign outputs[5061] = ~(layer0_outputs[5356]);
    assign outputs[5062] = ~(layer0_outputs[3168]);
    assign outputs[5063] = ~((layer0_outputs[6243]) | (layer0_outputs[4128]));
    assign outputs[5064] = ~(layer0_outputs[750]);
    assign outputs[5065] = layer0_outputs[6535];
    assign outputs[5066] = ~(layer0_outputs[1473]);
    assign outputs[5067] = (layer0_outputs[2387]) & ~(layer0_outputs[2887]);
    assign outputs[5068] = layer0_outputs[7074];
    assign outputs[5069] = layer0_outputs[7100];
    assign outputs[5070] = ~(layer0_outputs[2707]) | (layer0_outputs[3098]);
    assign outputs[5071] = (layer0_outputs[5523]) & ~(layer0_outputs[5341]);
    assign outputs[5072] = layer0_outputs[240];
    assign outputs[5073] = layer0_outputs[112];
    assign outputs[5074] = ~(layer0_outputs[3763]);
    assign outputs[5075] = ~(layer0_outputs[6699]);
    assign outputs[5076] = layer0_outputs[7472];
    assign outputs[5077] = (layer0_outputs[6088]) ^ (layer0_outputs[7335]);
    assign outputs[5078] = ~(layer0_outputs[2374]);
    assign outputs[5079] = ~(layer0_outputs[6505]);
    assign outputs[5080] = layer0_outputs[2434];
    assign outputs[5081] = layer0_outputs[6594];
    assign outputs[5082] = ~((layer0_outputs[6303]) | (layer0_outputs[5957]));
    assign outputs[5083] = ~((layer0_outputs[3994]) | (layer0_outputs[7183]));
    assign outputs[5084] = ~(layer0_outputs[3890]);
    assign outputs[5085] = (layer0_outputs[5479]) | (layer0_outputs[1238]);
    assign outputs[5086] = (layer0_outputs[195]) & ~(layer0_outputs[793]);
    assign outputs[5087] = ~((layer0_outputs[4445]) | (layer0_outputs[4262]));
    assign outputs[5088] = (layer0_outputs[2652]) ^ (layer0_outputs[2110]);
    assign outputs[5089] = layer0_outputs[4356];
    assign outputs[5090] = layer0_outputs[592];
    assign outputs[5091] = ~(layer0_outputs[4860]);
    assign outputs[5092] = layer0_outputs[6776];
    assign outputs[5093] = ~(layer0_outputs[5086]);
    assign outputs[5094] = ~((layer0_outputs[6813]) ^ (layer0_outputs[2689]));
    assign outputs[5095] = ~(layer0_outputs[546]);
    assign outputs[5096] = ~(layer0_outputs[3878]);
    assign outputs[5097] = 1'b1;
    assign outputs[5098] = layer0_outputs[47];
    assign outputs[5099] = layer0_outputs[487];
    assign outputs[5100] = (layer0_outputs[6336]) & ~(layer0_outputs[2347]);
    assign outputs[5101] = layer0_outputs[5924];
    assign outputs[5102] = (layer0_outputs[84]) & ~(layer0_outputs[4339]);
    assign outputs[5103] = (layer0_outputs[5835]) ^ (layer0_outputs[188]);
    assign outputs[5104] = (layer0_outputs[7202]) & ~(layer0_outputs[1211]);
    assign outputs[5105] = ~(layer0_outputs[1036]);
    assign outputs[5106] = layer0_outputs[1681];
    assign outputs[5107] = (layer0_outputs[4506]) ^ (layer0_outputs[3196]);
    assign outputs[5108] = layer0_outputs[649];
    assign outputs[5109] = ~((layer0_outputs[6039]) & (layer0_outputs[3261]));
    assign outputs[5110] = (layer0_outputs[2113]) ^ (layer0_outputs[3442]);
    assign outputs[5111] = layer0_outputs[5731];
    assign outputs[5112] = ~(layer0_outputs[7065]);
    assign outputs[5113] = ~(layer0_outputs[260]);
    assign outputs[5114] = ~((layer0_outputs[3612]) & (layer0_outputs[1246]));
    assign outputs[5115] = ~((layer0_outputs[397]) & (layer0_outputs[5013]));
    assign outputs[5116] = (layer0_outputs[2617]) & (layer0_outputs[6581]);
    assign outputs[5117] = ~((layer0_outputs[6177]) ^ (layer0_outputs[5315]));
    assign outputs[5118] = ~(layer0_outputs[6253]) | (layer0_outputs[5727]);
    assign outputs[5119] = ~(layer0_outputs[7464]);
    assign outputs[5120] = ~((layer0_outputs[4690]) | (layer0_outputs[4790]));
    assign outputs[5121] = ~(layer0_outputs[2199]);
    assign outputs[5122] = ~((layer0_outputs[2728]) ^ (layer0_outputs[2931]));
    assign outputs[5123] = ~(layer0_outputs[2805]);
    assign outputs[5124] = ~((layer0_outputs[6862]) | (layer0_outputs[6862]));
    assign outputs[5125] = (layer0_outputs[6353]) & (layer0_outputs[2686]);
    assign outputs[5126] = (layer0_outputs[2759]) ^ (layer0_outputs[31]);
    assign outputs[5127] = ~((layer0_outputs[1431]) ^ (layer0_outputs[5507]));
    assign outputs[5128] = (layer0_outputs[1519]) & ~(layer0_outputs[768]);
    assign outputs[5129] = ~(layer0_outputs[564]);
    assign outputs[5130] = layer0_outputs[2449];
    assign outputs[5131] = ~(layer0_outputs[1593]);
    assign outputs[5132] = layer0_outputs[6892];
    assign outputs[5133] = ~(layer0_outputs[1543]);
    assign outputs[5134] = ~((layer0_outputs[167]) & (layer0_outputs[800]));
    assign outputs[5135] = layer0_outputs[5211];
    assign outputs[5136] = layer0_outputs[1334];
    assign outputs[5137] = ~((layer0_outputs[7206]) ^ (layer0_outputs[5564]));
    assign outputs[5138] = ~((layer0_outputs[6469]) ^ (layer0_outputs[6748]));
    assign outputs[5139] = layer0_outputs[5806];
    assign outputs[5140] = (layer0_outputs[3704]) & (layer0_outputs[1902]);
    assign outputs[5141] = ~(layer0_outputs[1406]) | (layer0_outputs[7603]);
    assign outputs[5142] = (layer0_outputs[5221]) & (layer0_outputs[3332]);
    assign outputs[5143] = layer0_outputs[4725];
    assign outputs[5144] = layer0_outputs[2983];
    assign outputs[5145] = (layer0_outputs[1658]) ^ (layer0_outputs[6696]);
    assign outputs[5146] = ~((layer0_outputs[1533]) | (layer0_outputs[5644]));
    assign outputs[5147] = ~(layer0_outputs[3166]);
    assign outputs[5148] = ~(layer0_outputs[7184]);
    assign outputs[5149] = ~((layer0_outputs[3846]) & (layer0_outputs[1098]));
    assign outputs[5150] = (layer0_outputs[6756]) & ~(layer0_outputs[3404]);
    assign outputs[5151] = (layer0_outputs[6990]) ^ (layer0_outputs[1357]);
    assign outputs[5152] = layer0_outputs[2765];
    assign outputs[5153] = (layer0_outputs[1778]) & ~(layer0_outputs[3194]);
    assign outputs[5154] = (layer0_outputs[958]) | (layer0_outputs[5094]);
    assign outputs[5155] = layer0_outputs[5042];
    assign outputs[5156] = (layer0_outputs[6893]) & (layer0_outputs[1441]);
    assign outputs[5157] = ~(layer0_outputs[5925]) | (layer0_outputs[6024]);
    assign outputs[5158] = ~((layer0_outputs[2381]) ^ (layer0_outputs[6362]));
    assign outputs[5159] = ~((layer0_outputs[373]) ^ (layer0_outputs[1183]));
    assign outputs[5160] = layer0_outputs[4393];
    assign outputs[5161] = layer0_outputs[6310];
    assign outputs[5162] = ~(layer0_outputs[5174]);
    assign outputs[5163] = ~(layer0_outputs[4463]);
    assign outputs[5164] = layer0_outputs[1062];
    assign outputs[5165] = (layer0_outputs[2050]) ^ (layer0_outputs[5332]);
    assign outputs[5166] = (layer0_outputs[6806]) ^ (layer0_outputs[4163]);
    assign outputs[5167] = ~(layer0_outputs[379]);
    assign outputs[5168] = ~(layer0_outputs[6318]);
    assign outputs[5169] = (layer0_outputs[4685]) & ~(layer0_outputs[4936]);
    assign outputs[5170] = ~(layer0_outputs[5146]) | (layer0_outputs[2576]);
    assign outputs[5171] = ~(layer0_outputs[196]);
    assign outputs[5172] = ~((layer0_outputs[2566]) ^ (layer0_outputs[6396]));
    assign outputs[5173] = ~((layer0_outputs[3604]) ^ (layer0_outputs[84]));
    assign outputs[5174] = ~(layer0_outputs[5315]);
    assign outputs[5175] = layer0_outputs[2173];
    assign outputs[5176] = ~((layer0_outputs[4912]) ^ (layer0_outputs[2953]));
    assign outputs[5177] = ~(layer0_outputs[4256]);
    assign outputs[5178] = (layer0_outputs[4275]) & ~(layer0_outputs[2796]);
    assign outputs[5179] = (layer0_outputs[4699]) ^ (layer0_outputs[217]);
    assign outputs[5180] = layer0_outputs[2167];
    assign outputs[5181] = (layer0_outputs[711]) & ~(layer0_outputs[5047]);
    assign outputs[5182] = (layer0_outputs[4029]) ^ (layer0_outputs[3778]);
    assign outputs[5183] = ~(layer0_outputs[55]) | (layer0_outputs[1248]);
    assign outputs[5184] = ~(layer0_outputs[4017]);
    assign outputs[5185] = layer0_outputs[4443];
    assign outputs[5186] = layer0_outputs[4625];
    assign outputs[5187] = (layer0_outputs[3493]) ^ (layer0_outputs[4518]);
    assign outputs[5188] = layer0_outputs[6223];
    assign outputs[5189] = (layer0_outputs[2490]) ^ (layer0_outputs[5201]);
    assign outputs[5190] = ~(layer0_outputs[6462]);
    assign outputs[5191] = layer0_outputs[687];
    assign outputs[5192] = ~(layer0_outputs[1676]);
    assign outputs[5193] = (layer0_outputs[5970]) | (layer0_outputs[3208]);
    assign outputs[5194] = ~(layer0_outputs[5197]);
    assign outputs[5195] = ~((layer0_outputs[5879]) | (layer0_outputs[7313]));
    assign outputs[5196] = layer0_outputs[1260];
    assign outputs[5197] = ~(layer0_outputs[2624]) | (layer0_outputs[5178]);
    assign outputs[5198] = layer0_outputs[2165];
    assign outputs[5199] = (layer0_outputs[3119]) ^ (layer0_outputs[6269]);
    assign outputs[5200] = layer0_outputs[5744];
    assign outputs[5201] = layer0_outputs[2814];
    assign outputs[5202] = ~(layer0_outputs[5079]);
    assign outputs[5203] = (layer0_outputs[4177]) & ~(layer0_outputs[799]);
    assign outputs[5204] = layer0_outputs[6360];
    assign outputs[5205] = ~((layer0_outputs[1088]) | (layer0_outputs[3569]));
    assign outputs[5206] = ~((layer0_outputs[5722]) | (layer0_outputs[2591]));
    assign outputs[5207] = (layer0_outputs[6979]) ^ (layer0_outputs[4928]);
    assign outputs[5208] = (layer0_outputs[1389]) | (layer0_outputs[828]);
    assign outputs[5209] = layer0_outputs[1751];
    assign outputs[5210] = ~(layer0_outputs[5425]) | (layer0_outputs[2363]);
    assign outputs[5211] = ~(layer0_outputs[6713]);
    assign outputs[5212] = ~((layer0_outputs[4961]) ^ (layer0_outputs[3537]));
    assign outputs[5213] = ~(layer0_outputs[5032]);
    assign outputs[5214] = ~(layer0_outputs[5566]) | (layer0_outputs[7438]);
    assign outputs[5215] = (layer0_outputs[3047]) ^ (layer0_outputs[805]);
    assign outputs[5216] = layer0_outputs[5272];
    assign outputs[5217] = (layer0_outputs[6210]) & (layer0_outputs[1857]);
    assign outputs[5218] = (layer0_outputs[1484]) ^ (layer0_outputs[2626]);
    assign outputs[5219] = ~(layer0_outputs[1417]);
    assign outputs[5220] = ~((layer0_outputs[6072]) & (layer0_outputs[7666]));
    assign outputs[5221] = layer0_outputs[7386];
    assign outputs[5222] = layer0_outputs[6291];
    assign outputs[5223] = (layer0_outputs[7517]) & (layer0_outputs[6973]);
    assign outputs[5224] = layer0_outputs[4693];
    assign outputs[5225] = (layer0_outputs[366]) & ~(layer0_outputs[5212]);
    assign outputs[5226] = (layer0_outputs[2747]) & ~(layer0_outputs[5154]);
    assign outputs[5227] = (layer0_outputs[1187]) ^ (layer0_outputs[5752]);
    assign outputs[5228] = ~((layer0_outputs[98]) ^ (layer0_outputs[6478]));
    assign outputs[5229] = ~(layer0_outputs[5175]) | (layer0_outputs[6522]);
    assign outputs[5230] = 1'b1;
    assign outputs[5231] = ~(layer0_outputs[7672]) | (layer0_outputs[3861]);
    assign outputs[5232] = ~(layer0_outputs[5190]);
    assign outputs[5233] = ~(layer0_outputs[3846]);
    assign outputs[5234] = ~(layer0_outputs[755]) | (layer0_outputs[141]);
    assign outputs[5235] = ~((layer0_outputs[4264]) ^ (layer0_outputs[2120]));
    assign outputs[5236] = ~((layer0_outputs[1782]) ^ (layer0_outputs[6085]));
    assign outputs[5237] = layer0_outputs[116];
    assign outputs[5238] = layer0_outputs[6623];
    assign outputs[5239] = ~(layer0_outputs[2191]);
    assign outputs[5240] = (layer0_outputs[3335]) & (layer0_outputs[5568]);
    assign outputs[5241] = layer0_outputs[1413];
    assign outputs[5242] = (layer0_outputs[1560]) & ~(layer0_outputs[4643]);
    assign outputs[5243] = ~((layer0_outputs[5911]) | (layer0_outputs[4781]));
    assign outputs[5244] = layer0_outputs[7588];
    assign outputs[5245] = ~((layer0_outputs[7608]) ^ (layer0_outputs[5142]));
    assign outputs[5246] = layer0_outputs[4921];
    assign outputs[5247] = (layer0_outputs[7340]) ^ (layer0_outputs[1369]);
    assign outputs[5248] = ~(layer0_outputs[7261]);
    assign outputs[5249] = layer0_outputs[5693];
    assign outputs[5250] = (layer0_outputs[1775]) & (layer0_outputs[3122]);
    assign outputs[5251] = (layer0_outputs[7251]) ^ (layer0_outputs[6145]);
    assign outputs[5252] = ~((layer0_outputs[686]) | (layer0_outputs[1746]));
    assign outputs[5253] = layer0_outputs[3921];
    assign outputs[5254] = ~(layer0_outputs[4892]);
    assign outputs[5255] = (layer0_outputs[5693]) & (layer0_outputs[2747]);
    assign outputs[5256] = ~((layer0_outputs[530]) ^ (layer0_outputs[5441]));
    assign outputs[5257] = (layer0_outputs[1067]) & ~(layer0_outputs[7079]);
    assign outputs[5258] = ~((layer0_outputs[106]) ^ (layer0_outputs[2248]));
    assign outputs[5259] = ~(layer0_outputs[1615]);
    assign outputs[5260] = ~(layer0_outputs[3809]) | (layer0_outputs[4730]);
    assign outputs[5261] = (layer0_outputs[5784]) | (layer0_outputs[1425]);
    assign outputs[5262] = (layer0_outputs[3053]) ^ (layer0_outputs[6062]);
    assign outputs[5263] = (layer0_outputs[4837]) & ~(layer0_outputs[3547]);
    assign outputs[5264] = ~((layer0_outputs[6030]) ^ (layer0_outputs[271]));
    assign outputs[5265] = layer0_outputs[2166];
    assign outputs[5266] = ~(layer0_outputs[3716]) | (layer0_outputs[1006]);
    assign outputs[5267] = layer0_outputs[3696];
    assign outputs[5268] = ~(layer0_outputs[4447]);
    assign outputs[5269] = ~((layer0_outputs[516]) | (layer0_outputs[3307]));
    assign outputs[5270] = ~(layer0_outputs[4978]) | (layer0_outputs[58]);
    assign outputs[5271] = ~(layer0_outputs[5225]);
    assign outputs[5272] = (layer0_outputs[1915]) & (layer0_outputs[6277]);
    assign outputs[5273] = ~((layer0_outputs[7028]) & (layer0_outputs[1226]));
    assign outputs[5274] = ~(layer0_outputs[2656]) | (layer0_outputs[1606]);
    assign outputs[5275] = (layer0_outputs[3371]) ^ (layer0_outputs[3087]);
    assign outputs[5276] = ~((layer0_outputs[5621]) ^ (layer0_outputs[3818]));
    assign outputs[5277] = (layer0_outputs[6880]) | (layer0_outputs[190]);
    assign outputs[5278] = ~(layer0_outputs[4985]);
    assign outputs[5279] = ~(layer0_outputs[2749]);
    assign outputs[5280] = ~(layer0_outputs[7523]);
    assign outputs[5281] = layer0_outputs[3];
    assign outputs[5282] = ~((layer0_outputs[481]) | (layer0_outputs[154]));
    assign outputs[5283] = ~((layer0_outputs[4385]) ^ (layer0_outputs[3057]));
    assign outputs[5284] = (layer0_outputs[5455]) | (layer0_outputs[3098]);
    assign outputs[5285] = ~((layer0_outputs[2473]) | (layer0_outputs[2795]));
    assign outputs[5286] = ~(layer0_outputs[1622]);
    assign outputs[5287] = layer0_outputs[910];
    assign outputs[5288] = (layer0_outputs[1521]) & ~(layer0_outputs[1199]);
    assign outputs[5289] = ~(layer0_outputs[7447]);
    assign outputs[5290] = ~(layer0_outputs[5886]);
    assign outputs[5291] = layer0_outputs[3263];
    assign outputs[5292] = ~(layer0_outputs[6043]);
    assign outputs[5293] = ~(layer0_outputs[2696]);
    assign outputs[5294] = (layer0_outputs[5587]) ^ (layer0_outputs[3737]);
    assign outputs[5295] = ~((layer0_outputs[6584]) & (layer0_outputs[5853]));
    assign outputs[5296] = layer0_outputs[4948];
    assign outputs[5297] = ~(layer0_outputs[6714]);
    assign outputs[5298] = layer0_outputs[7240];
    assign outputs[5299] = ~(layer0_outputs[3589]) | (layer0_outputs[1657]);
    assign outputs[5300] = layer0_outputs[5593];
    assign outputs[5301] = (layer0_outputs[2099]) ^ (layer0_outputs[2586]);
    assign outputs[5302] = (layer0_outputs[3896]) ^ (layer0_outputs[6563]);
    assign outputs[5303] = ~(layer0_outputs[7201]);
    assign outputs[5304] = (layer0_outputs[1086]) & ~(layer0_outputs[1802]);
    assign outputs[5305] = (layer0_outputs[6711]) & ~(layer0_outputs[4993]);
    assign outputs[5306] = layer0_outputs[2196];
    assign outputs[5307] = layer0_outputs[6931];
    assign outputs[5308] = layer0_outputs[1035];
    assign outputs[5309] = (layer0_outputs[6233]) ^ (layer0_outputs[13]);
    assign outputs[5310] = ~(layer0_outputs[2823]);
    assign outputs[5311] = (layer0_outputs[3364]) & ~(layer0_outputs[7263]);
    assign outputs[5312] = ~((layer0_outputs[609]) ^ (layer0_outputs[89]));
    assign outputs[5313] = (layer0_outputs[7128]) ^ (layer0_outputs[3433]);
    assign outputs[5314] = layer0_outputs[1997];
    assign outputs[5315] = layer0_outputs[232];
    assign outputs[5316] = ~(layer0_outputs[7467]) | (layer0_outputs[2643]);
    assign outputs[5317] = (layer0_outputs[2840]) ^ (layer0_outputs[2793]);
    assign outputs[5318] = (layer0_outputs[1029]) ^ (layer0_outputs[4292]);
    assign outputs[5319] = ~(layer0_outputs[3264]) | (layer0_outputs[7037]);
    assign outputs[5320] = (layer0_outputs[7634]) & ~(layer0_outputs[3447]);
    assign outputs[5321] = ~(layer0_outputs[7068]) | (layer0_outputs[6148]);
    assign outputs[5322] = layer0_outputs[6982];
    assign outputs[5323] = layer0_outputs[5830];
    assign outputs[5324] = ~((layer0_outputs[4695]) ^ (layer0_outputs[7002]));
    assign outputs[5325] = layer0_outputs[5156];
    assign outputs[5326] = (layer0_outputs[6681]) & ~(layer0_outputs[2186]);
    assign outputs[5327] = ~((layer0_outputs[2937]) ^ (layer0_outputs[834]));
    assign outputs[5328] = layer0_outputs[663];
    assign outputs[5329] = (layer0_outputs[5036]) & ~(layer0_outputs[7676]);
    assign outputs[5330] = ~((layer0_outputs[5987]) ^ (layer0_outputs[382]));
    assign outputs[5331] = (layer0_outputs[104]) ^ (layer0_outputs[7322]);
    assign outputs[5332] = layer0_outputs[5132];
    assign outputs[5333] = ~(layer0_outputs[6439]);
    assign outputs[5334] = ~(layer0_outputs[4469]);
    assign outputs[5335] = layer0_outputs[5619];
    assign outputs[5336] = ~(layer0_outputs[2665]);
    assign outputs[5337] = ~(layer0_outputs[1075]);
    assign outputs[5338] = (layer0_outputs[3448]) & ~(layer0_outputs[4879]);
    assign outputs[5339] = ~(layer0_outputs[5465]);
    assign outputs[5340] = ~(layer0_outputs[3828]);
    assign outputs[5341] = layer0_outputs[4242];
    assign outputs[5342] = layer0_outputs[4189];
    assign outputs[5343] = layer0_outputs[7654];
    assign outputs[5344] = layer0_outputs[1000];
    assign outputs[5345] = layer0_outputs[116];
    assign outputs[5346] = layer0_outputs[3052];
    assign outputs[5347] = (layer0_outputs[1352]) ^ (layer0_outputs[3867]);
    assign outputs[5348] = layer0_outputs[5619];
    assign outputs[5349] = layer0_outputs[4205];
    assign outputs[5350] = ~(layer0_outputs[6447]) | (layer0_outputs[1113]);
    assign outputs[5351] = layer0_outputs[6008];
    assign outputs[5352] = layer0_outputs[4505];
    assign outputs[5353] = layer0_outputs[2670];
    assign outputs[5354] = ~((layer0_outputs[2217]) ^ (layer0_outputs[283]));
    assign outputs[5355] = ~((layer0_outputs[268]) ^ (layer0_outputs[1390]));
    assign outputs[5356] = ~(layer0_outputs[699]);
    assign outputs[5357] = ~(layer0_outputs[6890]);
    assign outputs[5358] = ~(layer0_outputs[4550]);
    assign outputs[5359] = ~(layer0_outputs[5106]);
    assign outputs[5360] = ~(layer0_outputs[6609]);
    assign outputs[5361] = (layer0_outputs[3452]) | (layer0_outputs[7045]);
    assign outputs[5362] = ~((layer0_outputs[4449]) | (layer0_outputs[1856]));
    assign outputs[5363] = ~(layer0_outputs[2]);
    assign outputs[5364] = ~((layer0_outputs[2389]) ^ (layer0_outputs[6064]));
    assign outputs[5365] = ~(layer0_outputs[952]) | (layer0_outputs[1335]);
    assign outputs[5366] = (layer0_outputs[5031]) ^ (layer0_outputs[483]);
    assign outputs[5367] = ~((layer0_outputs[3504]) | (layer0_outputs[2020]));
    assign outputs[5368] = (layer0_outputs[7588]) & ~(layer0_outputs[3925]);
    assign outputs[5369] = (layer0_outputs[7289]) ^ (layer0_outputs[6197]);
    assign outputs[5370] = ~((layer0_outputs[3814]) ^ (layer0_outputs[5052]));
    assign outputs[5371] = ~((layer0_outputs[1679]) ^ (layer0_outputs[7459]));
    assign outputs[5372] = ~(layer0_outputs[4415]);
    assign outputs[5373] = ~(layer0_outputs[1440]) | (layer0_outputs[2664]);
    assign outputs[5374] = layer0_outputs[5680];
    assign outputs[5375] = layer0_outputs[2339];
    assign outputs[5376] = layer0_outputs[4884];
    assign outputs[5377] = layer0_outputs[2493];
    assign outputs[5378] = layer0_outputs[4700];
    assign outputs[5379] = layer0_outputs[1286];
    assign outputs[5380] = layer0_outputs[1819];
    assign outputs[5381] = layer0_outputs[4137];
    assign outputs[5382] = ~(layer0_outputs[3990]);
    assign outputs[5383] = ~(layer0_outputs[1973]) | (layer0_outputs[2897]);
    assign outputs[5384] = (layer0_outputs[6652]) & ~(layer0_outputs[3325]);
    assign outputs[5385] = ~((layer0_outputs[6024]) | (layer0_outputs[6904]));
    assign outputs[5386] = layer0_outputs[7170];
    assign outputs[5387] = ~(layer0_outputs[187]);
    assign outputs[5388] = (layer0_outputs[3583]) & (layer0_outputs[5726]);
    assign outputs[5389] = layer0_outputs[4047];
    assign outputs[5390] = ~(layer0_outputs[1105]);
    assign outputs[5391] = ~(layer0_outputs[2294]);
    assign outputs[5392] = ~((layer0_outputs[5118]) | (layer0_outputs[2156]));
    assign outputs[5393] = layer0_outputs[4276];
    assign outputs[5394] = ~(layer0_outputs[2700]);
    assign outputs[5395] = ~(layer0_outputs[6189]);
    assign outputs[5396] = (layer0_outputs[267]) & (layer0_outputs[2716]);
    assign outputs[5397] = ~(layer0_outputs[4998]);
    assign outputs[5398] = (layer0_outputs[321]) | (layer0_outputs[849]);
    assign outputs[5399] = (layer0_outputs[1608]) ^ (layer0_outputs[2166]);
    assign outputs[5400] = ~(layer0_outputs[1639]);
    assign outputs[5401] = (layer0_outputs[175]) ^ (layer0_outputs[2101]);
    assign outputs[5402] = (layer0_outputs[2717]) & ~(layer0_outputs[425]);
    assign outputs[5403] = (layer0_outputs[5906]) & (layer0_outputs[7672]);
    assign outputs[5404] = ~(layer0_outputs[915]);
    assign outputs[5405] = ~(layer0_outputs[5258]);
    assign outputs[5406] = ~((layer0_outputs[1666]) ^ (layer0_outputs[6529]));
    assign outputs[5407] = (layer0_outputs[6610]) & ~(layer0_outputs[4975]);
    assign outputs[5408] = (layer0_outputs[4951]) & (layer0_outputs[4884]);
    assign outputs[5409] = layer0_outputs[3600];
    assign outputs[5410] = ~(layer0_outputs[387]);
    assign outputs[5411] = ~(layer0_outputs[2122]);
    assign outputs[5412] = ~(layer0_outputs[1238]);
    assign outputs[5413] = ~(layer0_outputs[4402]);
    assign outputs[5414] = ~(layer0_outputs[6037]);
    assign outputs[5415] = layer0_outputs[4016];
    assign outputs[5416] = ~((layer0_outputs[3255]) & (layer0_outputs[7032]));
    assign outputs[5417] = layer0_outputs[3680];
    assign outputs[5418] = layer0_outputs[6521];
    assign outputs[5419] = ~(layer0_outputs[5948]);
    assign outputs[5420] = layer0_outputs[4333];
    assign outputs[5421] = ~((layer0_outputs[5202]) | (layer0_outputs[2731]));
    assign outputs[5422] = ~((layer0_outputs[227]) ^ (layer0_outputs[3735]));
    assign outputs[5423] = ~((layer0_outputs[1019]) ^ (layer0_outputs[4228]));
    assign outputs[5424] = ~(layer0_outputs[3460]);
    assign outputs[5425] = layer0_outputs[2774];
    assign outputs[5426] = 1'b1;
    assign outputs[5427] = (layer0_outputs[4607]) ^ (layer0_outputs[2458]);
    assign outputs[5428] = ~((layer0_outputs[4349]) | (layer0_outputs[3501]));
    assign outputs[5429] = ~(layer0_outputs[245]);
    assign outputs[5430] = (layer0_outputs[1807]) & (layer0_outputs[563]);
    assign outputs[5431] = ~(layer0_outputs[824]);
    assign outputs[5432] = ~(layer0_outputs[5902]);
    assign outputs[5433] = (layer0_outputs[7378]) ^ (layer0_outputs[712]);
    assign outputs[5434] = ~(layer0_outputs[3123]);
    assign outputs[5435] = (layer0_outputs[1649]) & (layer0_outputs[2581]);
    assign outputs[5436] = ~((layer0_outputs[4461]) | (layer0_outputs[1215]));
    assign outputs[5437] = ~(layer0_outputs[6677]);
    assign outputs[5438] = layer0_outputs[7513];
    assign outputs[5439] = layer0_outputs[7034];
    assign outputs[5440] = (layer0_outputs[2707]) & (layer0_outputs[4745]);
    assign outputs[5441] = ~((layer0_outputs[5499]) ^ (layer0_outputs[6492]));
    assign outputs[5442] = ~((layer0_outputs[2764]) | (layer0_outputs[4371]));
    assign outputs[5443] = layer0_outputs[1394];
    assign outputs[5444] = (layer0_outputs[6637]) & (layer0_outputs[5930]);
    assign outputs[5445] = ~(layer0_outputs[7127]) | (layer0_outputs[2961]);
    assign outputs[5446] = ~((layer0_outputs[2448]) ^ (layer0_outputs[1722]));
    assign outputs[5447] = layer0_outputs[2772];
    assign outputs[5448] = layer0_outputs[7633];
    assign outputs[5449] = layer0_outputs[7026];
    assign outputs[5450] = ~(layer0_outputs[5889]);
    assign outputs[5451] = (layer0_outputs[4777]) & ~(layer0_outputs[3819]);
    assign outputs[5452] = ~(layer0_outputs[7129]);
    assign outputs[5453] = (layer0_outputs[3848]) ^ (layer0_outputs[439]);
    assign outputs[5454] = ~((layer0_outputs[1512]) | (layer0_outputs[5901]));
    assign outputs[5455] = ~(layer0_outputs[595]) | (layer0_outputs[1102]);
    assign outputs[5456] = (layer0_outputs[4511]) & ~(layer0_outputs[6657]);
    assign outputs[5457] = (layer0_outputs[6665]) ^ (layer0_outputs[1720]);
    assign outputs[5458] = ~(layer0_outputs[4657]);
    assign outputs[5459] = (layer0_outputs[1483]) ^ (layer0_outputs[4827]);
    assign outputs[5460] = layer0_outputs[6248];
    assign outputs[5461] = ~(layer0_outputs[833]);
    assign outputs[5462] = layer0_outputs[4499];
    assign outputs[5463] = ~(layer0_outputs[4362]);
    assign outputs[5464] = ~(layer0_outputs[745]) | (layer0_outputs[5697]);
    assign outputs[5465] = (layer0_outputs[3128]) ^ (layer0_outputs[1601]);
    assign outputs[5466] = layer0_outputs[1659];
    assign outputs[5467] = ~(layer0_outputs[6445]) | (layer0_outputs[887]);
    assign outputs[5468] = ~((layer0_outputs[6217]) & (layer0_outputs[423]));
    assign outputs[5469] = (layer0_outputs[3192]) ^ (layer0_outputs[296]);
    assign outputs[5470] = ~((layer0_outputs[319]) & (layer0_outputs[3174]));
    assign outputs[5471] = (layer0_outputs[265]) & (layer0_outputs[6797]);
    assign outputs[5472] = ~(layer0_outputs[3448]) | (layer0_outputs[2848]);
    assign outputs[5473] = (layer0_outputs[2515]) & ~(layer0_outputs[2102]);
    assign outputs[5474] = ~(layer0_outputs[5938]);
    assign outputs[5475] = (layer0_outputs[5683]) & ~(layer0_outputs[2152]);
    assign outputs[5476] = (layer0_outputs[3623]) & ~(layer0_outputs[7082]);
    assign outputs[5477] = ~(layer0_outputs[1910]) | (layer0_outputs[552]);
    assign outputs[5478] = ~(layer0_outputs[2642]);
    assign outputs[5479] = (layer0_outputs[5608]) & ~(layer0_outputs[3256]);
    assign outputs[5480] = ~(layer0_outputs[4863]);
    assign outputs[5481] = (layer0_outputs[7087]) & ~(layer0_outputs[2076]);
    assign outputs[5482] = ~(layer0_outputs[2338]) | (layer0_outputs[3010]);
    assign outputs[5483] = ~((layer0_outputs[5209]) ^ (layer0_outputs[6378]));
    assign outputs[5484] = (layer0_outputs[7344]) & (layer0_outputs[4555]);
    assign outputs[5485] = ~(layer0_outputs[1698]);
    assign outputs[5486] = ~((layer0_outputs[7109]) | (layer0_outputs[3860]));
    assign outputs[5487] = layer0_outputs[1963];
    assign outputs[5488] = layer0_outputs[4745];
    assign outputs[5489] = layer0_outputs[852];
    assign outputs[5490] = ~((layer0_outputs[3854]) | (layer0_outputs[148]));
    assign outputs[5491] = ~(layer0_outputs[1384]);
    assign outputs[5492] = (layer0_outputs[4301]) & ~(layer0_outputs[496]);
    assign outputs[5493] = (layer0_outputs[1831]) | (layer0_outputs[7495]);
    assign outputs[5494] = ~(layer0_outputs[5424]);
    assign outputs[5495] = (layer0_outputs[5624]) ^ (layer0_outputs[5223]);
    assign outputs[5496] = (layer0_outputs[6384]) & ~(layer0_outputs[1033]);
    assign outputs[5497] = ~(layer0_outputs[1148]) | (layer0_outputs[5883]);
    assign outputs[5498] = ~((layer0_outputs[1722]) ^ (layer0_outputs[6816]));
    assign outputs[5499] = ~((layer0_outputs[2978]) | (layer0_outputs[1216]));
    assign outputs[5500] = (layer0_outputs[7557]) & (layer0_outputs[4584]);
    assign outputs[5501] = ~((layer0_outputs[4932]) | (layer0_outputs[4111]));
    assign outputs[5502] = layer0_outputs[4187];
    assign outputs[5503] = layer0_outputs[2874];
    assign outputs[5504] = layer0_outputs[2929];
    assign outputs[5505] = layer0_outputs[6215];
    assign outputs[5506] = ~((layer0_outputs[2987]) | (layer0_outputs[7383]));
    assign outputs[5507] = layer0_outputs[6262];
    assign outputs[5508] = layer0_outputs[2008];
    assign outputs[5509] = ~((layer0_outputs[1512]) | (layer0_outputs[2703]));
    assign outputs[5510] = ~(layer0_outputs[5912]);
    assign outputs[5511] = (layer0_outputs[5307]) & (layer0_outputs[1457]);
    assign outputs[5512] = ~((layer0_outputs[112]) ^ (layer0_outputs[6165]));
    assign outputs[5513] = ~(layer0_outputs[4113]);
    assign outputs[5514] = ~((layer0_outputs[4646]) | (layer0_outputs[5803]));
    assign outputs[5515] = layer0_outputs[6532];
    assign outputs[5516] = layer0_outputs[6492];
    assign outputs[5517] = (layer0_outputs[1157]) & ~(layer0_outputs[5364]);
    assign outputs[5518] = layer0_outputs[1361];
    assign outputs[5519] = ~(layer0_outputs[5409]);
    assign outputs[5520] = (layer0_outputs[4894]) & (layer0_outputs[3319]);
    assign outputs[5521] = (layer0_outputs[780]) & ~(layer0_outputs[3083]);
    assign outputs[5522] = (layer0_outputs[2791]) & (layer0_outputs[4246]);
    assign outputs[5523] = ~(layer0_outputs[1525]) | (layer0_outputs[2623]);
    assign outputs[5524] = layer0_outputs[1411];
    assign outputs[5525] = layer0_outputs[7060];
    assign outputs[5526] = layer0_outputs[1641];
    assign outputs[5527] = (layer0_outputs[5674]) & ~(layer0_outputs[4309]);
    assign outputs[5528] = (layer0_outputs[1360]) | (layer0_outputs[4098]);
    assign outputs[5529] = layer0_outputs[3707];
    assign outputs[5530] = ~(layer0_outputs[715]);
    assign outputs[5531] = ~(layer0_outputs[4078]);
    assign outputs[5532] = ~((layer0_outputs[3751]) ^ (layer0_outputs[1330]));
    assign outputs[5533] = layer0_outputs[2658];
    assign outputs[5534] = (layer0_outputs[1553]) | (layer0_outputs[1322]);
    assign outputs[5535] = (layer0_outputs[4059]) ^ (layer0_outputs[4174]);
    assign outputs[5536] = ~((layer0_outputs[709]) | (layer0_outputs[3918]));
    assign outputs[5537] = ~(layer0_outputs[4503]) | (layer0_outputs[864]);
    assign outputs[5538] = ~(layer0_outputs[4013]);
    assign outputs[5539] = ~((layer0_outputs[3305]) | (layer0_outputs[5081]));
    assign outputs[5540] = ~(layer0_outputs[1263]);
    assign outputs[5541] = ~(layer0_outputs[428]);
    assign outputs[5542] = (layer0_outputs[3525]) ^ (layer0_outputs[4464]);
    assign outputs[5543] = ~(layer0_outputs[3582]);
    assign outputs[5544] = (layer0_outputs[6687]) ^ (layer0_outputs[7646]);
    assign outputs[5545] = layer0_outputs[2998];
    assign outputs[5546] = (layer0_outputs[4498]) | (layer0_outputs[4641]);
    assign outputs[5547] = ~((layer0_outputs[156]) ^ (layer0_outputs[2048]));
    assign outputs[5548] = ~(layer0_outputs[2991]);
    assign outputs[5549] = (layer0_outputs[1298]) & ~(layer0_outputs[5502]);
    assign outputs[5550] = layer0_outputs[2141];
    assign outputs[5551] = ~(layer0_outputs[6884]);
    assign outputs[5552] = layer0_outputs[4862];
    assign outputs[5553] = (layer0_outputs[2667]) ^ (layer0_outputs[3171]);
    assign outputs[5554] = layer0_outputs[5729];
    assign outputs[5555] = ~(layer0_outputs[3446]);
    assign outputs[5556] = ~(layer0_outputs[1550]);
    assign outputs[5557] = ~((layer0_outputs[1716]) ^ (layer0_outputs[168]));
    assign outputs[5558] = ~(layer0_outputs[6079]);
    assign outputs[5559] = layer0_outputs[1128];
    assign outputs[5560] = (layer0_outputs[4810]) | (layer0_outputs[1802]);
    assign outputs[5561] = ~(layer0_outputs[2236]) | (layer0_outputs[6598]);
    assign outputs[5562] = layer0_outputs[324];
    assign outputs[5563] = layer0_outputs[6256];
    assign outputs[5564] = layer0_outputs[5918];
    assign outputs[5565] = layer0_outputs[4934];
    assign outputs[5566] = ~(layer0_outputs[4606]);
    assign outputs[5567] = (layer0_outputs[1457]) & ~(layer0_outputs[3422]);
    assign outputs[5568] = ~(layer0_outputs[3333]);
    assign outputs[5569] = (layer0_outputs[6269]) & ~(layer0_outputs[969]);
    assign outputs[5570] = layer0_outputs[3271];
    assign outputs[5571] = (layer0_outputs[1078]) ^ (layer0_outputs[6726]);
    assign outputs[5572] = ~((layer0_outputs[584]) ^ (layer0_outputs[5915]));
    assign outputs[5573] = layer0_outputs[4329];
    assign outputs[5574] = (layer0_outputs[3030]) & (layer0_outputs[3949]);
    assign outputs[5575] = (layer0_outputs[5613]) & (layer0_outputs[6916]);
    assign outputs[5576] = ~((layer0_outputs[3661]) ^ (layer0_outputs[1757]));
    assign outputs[5577] = ~(layer0_outputs[2627]) | (layer0_outputs[3076]);
    assign outputs[5578] = ~(layer0_outputs[2645]);
    assign outputs[5579] = ~((layer0_outputs[3981]) ^ (layer0_outputs[6348]));
    assign outputs[5580] = (layer0_outputs[7059]) & ~(layer0_outputs[2496]);
    assign outputs[5581] = (layer0_outputs[2906]) ^ (layer0_outputs[5443]);
    assign outputs[5582] = layer0_outputs[7067];
    assign outputs[5583] = ~(layer0_outputs[5404]);
    assign outputs[5584] = ~(layer0_outputs[1229]);
    assign outputs[5585] = (layer0_outputs[5136]) & (layer0_outputs[3623]);
    assign outputs[5586] = layer0_outputs[6502];
    assign outputs[5587] = layer0_outputs[3209];
    assign outputs[5588] = (layer0_outputs[5743]) & ~(layer0_outputs[554]);
    assign outputs[5589] = (layer0_outputs[2954]) | (layer0_outputs[7569]);
    assign outputs[5590] = ~((layer0_outputs[4164]) ^ (layer0_outputs[5321]));
    assign outputs[5591] = layer0_outputs[3533];
    assign outputs[5592] = ~(layer0_outputs[1970]) | (layer0_outputs[7285]);
    assign outputs[5593] = ~(layer0_outputs[5593]) | (layer0_outputs[1727]);
    assign outputs[5594] = 1'b0;
    assign outputs[5595] = layer0_outputs[5088];
    assign outputs[5596] = layer0_outputs[7607];
    assign outputs[5597] = (layer0_outputs[2000]) | (layer0_outputs[5638]);
    assign outputs[5598] = layer0_outputs[4784];
    assign outputs[5599] = ~(layer0_outputs[7038]);
    assign outputs[5600] = ~((layer0_outputs[5453]) | (layer0_outputs[3140]));
    assign outputs[5601] = ~(layer0_outputs[5798]);
    assign outputs[5602] = ~((layer0_outputs[80]) | (layer0_outputs[6928]));
    assign outputs[5603] = ~(layer0_outputs[1944]);
    assign outputs[5604] = layer0_outputs[2458];
    assign outputs[5605] = (layer0_outputs[6904]) & ~(layer0_outputs[4511]);
    assign outputs[5606] = (layer0_outputs[6987]) & (layer0_outputs[5283]);
    assign outputs[5607] = ~(layer0_outputs[7077]);
    assign outputs[5608] = ~((layer0_outputs[2453]) ^ (layer0_outputs[2186]));
    assign outputs[5609] = (layer0_outputs[6671]) ^ (layer0_outputs[4347]);
    assign outputs[5610] = (layer0_outputs[7579]) & (layer0_outputs[1001]);
    assign outputs[5611] = ~(layer0_outputs[3853]);
    assign outputs[5612] = layer0_outputs[3574];
    assign outputs[5613] = ~((layer0_outputs[7269]) | (layer0_outputs[3648]));
    assign outputs[5614] = 1'b0;
    assign outputs[5615] = ~((layer0_outputs[1180]) ^ (layer0_outputs[3403]));
    assign outputs[5616] = ~(layer0_outputs[3347]);
    assign outputs[5617] = ~(layer0_outputs[2439]);
    assign outputs[5618] = (layer0_outputs[6393]) ^ (layer0_outputs[1882]);
    assign outputs[5619] = ~((layer0_outputs[4249]) ^ (layer0_outputs[3240]));
    assign outputs[5620] = ~(layer0_outputs[5145]);
    assign outputs[5621] = layer0_outputs[3922];
    assign outputs[5622] = ~(layer0_outputs[775]) | (layer0_outputs[3091]);
    assign outputs[5623] = (layer0_outputs[4848]) & ~(layer0_outputs[4056]);
    assign outputs[5624] = (layer0_outputs[3938]) & ~(layer0_outputs[2979]);
    assign outputs[5625] = (layer0_outputs[7465]) ^ (layer0_outputs[3786]);
    assign outputs[5626] = ~(layer0_outputs[3364]);
    assign outputs[5627] = ~(layer0_outputs[1339]);
    assign outputs[5628] = ~((layer0_outputs[4424]) ^ (layer0_outputs[4474]));
    assign outputs[5629] = layer0_outputs[1975];
    assign outputs[5630] = layer0_outputs[5411];
    assign outputs[5631] = (layer0_outputs[7659]) & ~(layer0_outputs[5577]);
    assign outputs[5632] = ~((layer0_outputs[3321]) ^ (layer0_outputs[2394]));
    assign outputs[5633] = ~(layer0_outputs[667]);
    assign outputs[5634] = ~((layer0_outputs[2434]) | (layer0_outputs[464]));
    assign outputs[5635] = ~(layer0_outputs[2593]);
    assign outputs[5636] = (layer0_outputs[4364]) & ~(layer0_outputs[1374]);
    assign outputs[5637] = layer0_outputs[2089];
    assign outputs[5638] = layer0_outputs[6363];
    assign outputs[5639] = (layer0_outputs[5937]) & ~(layer0_outputs[6138]);
    assign outputs[5640] = ~((layer0_outputs[1638]) ^ (layer0_outputs[2787]));
    assign outputs[5641] = ~(layer0_outputs[7297]);
    assign outputs[5642] = ~(layer0_outputs[4306]);
    assign outputs[5643] = layer0_outputs[4355];
    assign outputs[5644] = ~((layer0_outputs[5464]) | (layer0_outputs[1143]));
    assign outputs[5645] = ~(layer0_outputs[5014]);
    assign outputs[5646] = (layer0_outputs[7400]) & ~(layer0_outputs[148]);
    assign outputs[5647] = ~((layer0_outputs[251]) ^ (layer0_outputs[828]));
    assign outputs[5648] = (layer0_outputs[1018]) ^ (layer0_outputs[442]);
    assign outputs[5649] = layer0_outputs[2744];
    assign outputs[5650] = (layer0_outputs[4142]) & ~(layer0_outputs[7598]);
    assign outputs[5651] = ~((layer0_outputs[3874]) | (layer0_outputs[467]));
    assign outputs[5652] = ~((layer0_outputs[770]) ^ (layer0_outputs[6163]));
    assign outputs[5653] = (layer0_outputs[7484]) & ~(layer0_outputs[7293]);
    assign outputs[5654] = layer0_outputs[5380];
    assign outputs[5655] = ~(layer0_outputs[688]);
    assign outputs[5656] = ~(layer0_outputs[4085]);
    assign outputs[5657] = ~((layer0_outputs[404]) & (layer0_outputs[110]));
    assign outputs[5658] = ~(layer0_outputs[3437]);
    assign outputs[5659] = layer0_outputs[4562];
    assign outputs[5660] = ~((layer0_outputs[5549]) | (layer0_outputs[6617]));
    assign outputs[5661] = ~((layer0_outputs[1945]) ^ (layer0_outputs[0]));
    assign outputs[5662] = ~((layer0_outputs[6633]) & (layer0_outputs[133]));
    assign outputs[5663] = ~(layer0_outputs[3978]);
    assign outputs[5664] = layer0_outputs[2801];
    assign outputs[5665] = ~(layer0_outputs[115]);
    assign outputs[5666] = ~((layer0_outputs[4867]) ^ (layer0_outputs[1303]));
    assign outputs[5667] = (layer0_outputs[1962]) & (layer0_outputs[5476]);
    assign outputs[5668] = ~((layer0_outputs[3064]) | (layer0_outputs[2482]));
    assign outputs[5669] = (layer0_outputs[1139]) & ~(layer0_outputs[398]);
    assign outputs[5670] = layer0_outputs[3832];
    assign outputs[5671] = ~(layer0_outputs[2427]);
    assign outputs[5672] = layer0_outputs[6696];
    assign outputs[5673] = (layer0_outputs[126]) ^ (layer0_outputs[3753]);
    assign outputs[5674] = layer0_outputs[4012];
    assign outputs[5675] = (layer0_outputs[3711]) | (layer0_outputs[3758]);
    assign outputs[5676] = ~(layer0_outputs[1331]);
    assign outputs[5677] = (layer0_outputs[3049]) & ~(layer0_outputs[5418]);
    assign outputs[5678] = ~(layer0_outputs[1305]);
    assign outputs[5679] = (layer0_outputs[1259]) & ~(layer0_outputs[2457]);
    assign outputs[5680] = (layer0_outputs[2775]) & ~(layer0_outputs[3389]);
    assign outputs[5681] = ~(layer0_outputs[4458]) | (layer0_outputs[1494]);
    assign outputs[5682] = ~(layer0_outputs[7460]);
    assign outputs[5683] = (layer0_outputs[87]) & ~(layer0_outputs[82]);
    assign outputs[5684] = ~(layer0_outputs[641]);
    assign outputs[5685] = ~(layer0_outputs[1571]);
    assign outputs[5686] = ~((layer0_outputs[5281]) | (layer0_outputs[1044]));
    assign outputs[5687] = ~((layer0_outputs[6999]) ^ (layer0_outputs[946]));
    assign outputs[5688] = layer0_outputs[4744];
    assign outputs[5689] = layer0_outputs[3653];
    assign outputs[5690] = layer0_outputs[5956];
    assign outputs[5691] = (layer0_outputs[341]) | (layer0_outputs[5018]);
    assign outputs[5692] = (layer0_outputs[7204]) & (layer0_outputs[5029]);
    assign outputs[5693] = (layer0_outputs[1123]) & (layer0_outputs[6041]);
    assign outputs[5694] = layer0_outputs[7230];
    assign outputs[5695] = (layer0_outputs[1964]) ^ (layer0_outputs[2444]);
    assign outputs[5696] = ~(layer0_outputs[4052]);
    assign outputs[5697] = ~(layer0_outputs[2132]) | (layer0_outputs[708]);
    assign outputs[5698] = (layer0_outputs[691]) & (layer0_outputs[1367]);
    assign outputs[5699] = layer0_outputs[4261];
    assign outputs[5700] = (layer0_outputs[819]) ^ (layer0_outputs[2673]);
    assign outputs[5701] = (layer0_outputs[61]) ^ (layer0_outputs[5528]);
    assign outputs[5702] = (layer0_outputs[3529]) & ~(layer0_outputs[3793]);
    assign outputs[5703] = layer0_outputs[2408];
    assign outputs[5704] = (layer0_outputs[4634]) ^ (layer0_outputs[5907]);
    assign outputs[5705] = (layer0_outputs[6980]) & ~(layer0_outputs[5045]);
    assign outputs[5706] = (layer0_outputs[1973]) ^ (layer0_outputs[2589]);
    assign outputs[5707] = ~((layer0_outputs[1749]) ^ (layer0_outputs[3203]));
    assign outputs[5708] = ~(layer0_outputs[6073]);
    assign outputs[5709] = (layer0_outputs[1674]) & (layer0_outputs[140]);
    assign outputs[5710] = ~(layer0_outputs[3945]);
    assign outputs[5711] = layer0_outputs[495];
    assign outputs[5712] = ~((layer0_outputs[2563]) ^ (layer0_outputs[2584]));
    assign outputs[5713] = ~(layer0_outputs[242]);
    assign outputs[5714] = ~(layer0_outputs[6404]) | (layer0_outputs[4182]);
    assign outputs[5715] = ~(layer0_outputs[4523]);
    assign outputs[5716] = ~(layer0_outputs[3014]);
    assign outputs[5717] = ~((layer0_outputs[5403]) ^ (layer0_outputs[4040]));
    assign outputs[5718] = ~(layer0_outputs[395]);
    assign outputs[5719] = (layer0_outputs[3822]) & ~(layer0_outputs[4730]);
    assign outputs[5720] = ~(layer0_outputs[5891]);
    assign outputs[5721] = (layer0_outputs[5864]) ^ (layer0_outputs[6276]);
    assign outputs[5722] = ~((layer0_outputs[7543]) ^ (layer0_outputs[4279]));
    assign outputs[5723] = (layer0_outputs[6201]) & ~(layer0_outputs[799]);
    assign outputs[5724] = layer0_outputs[7102];
    assign outputs[5725] = (layer0_outputs[162]) ^ (layer0_outputs[6850]);
    assign outputs[5726] = layer0_outputs[3276];
    assign outputs[5727] = ~((layer0_outputs[2558]) ^ (layer0_outputs[6653]));
    assign outputs[5728] = (layer0_outputs[6519]) & (layer0_outputs[2159]);
    assign outputs[5729] = (layer0_outputs[5172]) & ~(layer0_outputs[1562]);
    assign outputs[5730] = (layer0_outputs[2441]) & ~(layer0_outputs[695]);
    assign outputs[5731] = ~(layer0_outputs[7451]) | (layer0_outputs[7084]);
    assign outputs[5732] = (layer0_outputs[4456]) & ~(layer0_outputs[4646]);
    assign outputs[5733] = ~(layer0_outputs[221]);
    assign outputs[5734] = ~((layer0_outputs[1099]) ^ (layer0_outputs[6876]));
    assign outputs[5735] = (layer0_outputs[3066]) & (layer0_outputs[4389]);
    assign outputs[5736] = (layer0_outputs[6121]) | (layer0_outputs[850]);
    assign outputs[5737] = ~(layer0_outputs[7272]);
    assign outputs[5738] = (layer0_outputs[7071]) | (layer0_outputs[3470]);
    assign outputs[5739] = ~(layer0_outputs[1769]) | (layer0_outputs[5143]);
    assign outputs[5740] = layer0_outputs[5349];
    assign outputs[5741] = layer0_outputs[4021];
    assign outputs[5742] = ~(layer0_outputs[2885]) | (layer0_outputs[5433]);
    assign outputs[5743] = 1'b0;
    assign outputs[5744] = (layer0_outputs[2864]) & ~(layer0_outputs[155]);
    assign outputs[5745] = (layer0_outputs[7638]) ^ (layer0_outputs[5358]);
    assign outputs[5746] = (layer0_outputs[4999]) ^ (layer0_outputs[2277]);
    assign outputs[5747] = layer0_outputs[5608];
    assign outputs[5748] = ~(layer0_outputs[7449]);
    assign outputs[5749] = (layer0_outputs[105]) & ~(layer0_outputs[5998]);
    assign outputs[5750] = ~(layer0_outputs[2250]);
    assign outputs[5751] = (layer0_outputs[1146]) ^ (layer0_outputs[7023]);
    assign outputs[5752] = ~((layer0_outputs[5911]) | (layer0_outputs[949]));
    assign outputs[5753] = (layer0_outputs[3084]) & ~(layer0_outputs[4192]);
    assign outputs[5754] = layer0_outputs[5850];
    assign outputs[5755] = layer0_outputs[6403];
    assign outputs[5756] = ~(layer0_outputs[5573]);
    assign outputs[5757] = ~(layer0_outputs[5122]);
    assign outputs[5758] = ~((layer0_outputs[4249]) | (layer0_outputs[11]));
    assign outputs[5759] = layer0_outputs[6097];
    assign outputs[5760] = (layer0_outputs[3958]) & ~(layer0_outputs[3035]);
    assign outputs[5761] = layer0_outputs[1469];
    assign outputs[5762] = ~(layer0_outputs[7626]);
    assign outputs[5763] = ~(layer0_outputs[6147]) | (layer0_outputs[3507]);
    assign outputs[5764] = ~((layer0_outputs[4702]) | (layer0_outputs[4349]));
    assign outputs[5765] = layer0_outputs[4995];
    assign outputs[5766] = ~((layer0_outputs[4431]) ^ (layer0_outputs[972]));
    assign outputs[5767] = (layer0_outputs[4521]) & ~(layer0_outputs[4766]);
    assign outputs[5768] = (layer0_outputs[714]) & ~(layer0_outputs[6896]);
    assign outputs[5769] = ~((layer0_outputs[3079]) ^ (layer0_outputs[6843]));
    assign outputs[5770] = ~((layer0_outputs[7147]) ^ (layer0_outputs[4948]));
    assign outputs[5771] = ~(layer0_outputs[6920]);
    assign outputs[5772] = (layer0_outputs[5855]) ^ (layer0_outputs[2485]);
    assign outputs[5773] = ~((layer0_outputs[1727]) ^ (layer0_outputs[5519]));
    assign outputs[5774] = (layer0_outputs[6304]) & ~(layer0_outputs[6360]);
    assign outputs[5775] = (layer0_outputs[979]) ^ (layer0_outputs[4120]);
    assign outputs[5776] = (layer0_outputs[5158]) ^ (layer0_outputs[7377]);
    assign outputs[5777] = (layer0_outputs[2945]) & (layer0_outputs[2249]);
    assign outputs[5778] = (layer0_outputs[724]) & (layer0_outputs[3060]);
    assign outputs[5779] = layer0_outputs[4535];
    assign outputs[5780] = (layer0_outputs[5057]) & ~(layer0_outputs[5959]);
    assign outputs[5781] = ~(layer0_outputs[6625]) | (layer0_outputs[6484]);
    assign outputs[5782] = ~(layer0_outputs[5800]);
    assign outputs[5783] = layer0_outputs[7026];
    assign outputs[5784] = (layer0_outputs[3509]) & (layer0_outputs[4671]);
    assign outputs[5785] = ~((layer0_outputs[1138]) ^ (layer0_outputs[1801]));
    assign outputs[5786] = ~(layer0_outputs[506]) | (layer0_outputs[457]);
    assign outputs[5787] = ~(layer0_outputs[3140]);
    assign outputs[5788] = ~((layer0_outputs[5483]) ^ (layer0_outputs[5375]));
    assign outputs[5789] = ~((layer0_outputs[191]) | (layer0_outputs[4401]));
    assign outputs[5790] = layer0_outputs[2992];
    assign outputs[5791] = layer0_outputs[4026];
    assign outputs[5792] = layer0_outputs[1388];
    assign outputs[5793] = ~(layer0_outputs[4631]);
    assign outputs[5794] = layer0_outputs[73];
    assign outputs[5795] = (layer0_outputs[7127]) & (layer0_outputs[173]);
    assign outputs[5796] = ~((layer0_outputs[6939]) & (layer0_outputs[3726]));
    assign outputs[5797] = ~((layer0_outputs[7664]) ^ (layer0_outputs[2290]));
    assign outputs[5798] = layer0_outputs[515];
    assign outputs[5799] = ~(layer0_outputs[4266]);
    assign outputs[5800] = layer0_outputs[3755];
    assign outputs[5801] = ~(layer0_outputs[4215]);
    assign outputs[5802] = ~((layer0_outputs[6539]) ^ (layer0_outputs[1438]));
    assign outputs[5803] = layer0_outputs[6815];
    assign outputs[5804] = ~((layer0_outputs[1429]) ^ (layer0_outputs[6413]));
    assign outputs[5805] = (layer0_outputs[535]) & ~(layer0_outputs[2357]);
    assign outputs[5806] = layer0_outputs[6157];
    assign outputs[5807] = ~(layer0_outputs[4804]);
    assign outputs[5808] = (layer0_outputs[3871]) ^ (layer0_outputs[3093]);
    assign outputs[5809] = (layer0_outputs[3969]) & ~(layer0_outputs[288]);
    assign outputs[5810] = (layer0_outputs[5672]) | (layer0_outputs[3545]);
    assign outputs[5811] = layer0_outputs[4507];
    assign outputs[5812] = ~(layer0_outputs[5220]);
    assign outputs[5813] = ~(layer0_outputs[2187]) | (layer0_outputs[4893]);
    assign outputs[5814] = (layer0_outputs[1467]) & ~(layer0_outputs[2719]);
    assign outputs[5815] = ~(layer0_outputs[3872]);
    assign outputs[5816] = (layer0_outputs[4336]) & ~(layer0_outputs[6114]);
    assign outputs[5817] = 1'b0;
    assign outputs[5818] = ~((layer0_outputs[4952]) ^ (layer0_outputs[671]));
    assign outputs[5819] = (layer0_outputs[2207]) & ~(layer0_outputs[5040]);
    assign outputs[5820] = (layer0_outputs[6515]) ^ (layer0_outputs[6901]);
    assign outputs[5821] = (layer0_outputs[4488]) ^ (layer0_outputs[2686]);
    assign outputs[5822] = ~((layer0_outputs[3898]) | (layer0_outputs[3311]));
    assign outputs[5823] = layer0_outputs[3849];
    assign outputs[5824] = ~(layer0_outputs[4903]);
    assign outputs[5825] = ~(layer0_outputs[977]);
    assign outputs[5826] = ~(layer0_outputs[1739]);
    assign outputs[5827] = ~((layer0_outputs[3270]) | (layer0_outputs[4580]));
    assign outputs[5828] = (layer0_outputs[3876]) ^ (layer0_outputs[6588]);
    assign outputs[5829] = ~((layer0_outputs[5058]) | (layer0_outputs[4797]));
    assign outputs[5830] = ~((layer0_outputs[4731]) ^ (layer0_outputs[7534]));
    assign outputs[5831] = ~(layer0_outputs[7216]);
    assign outputs[5832] = layer0_outputs[3724];
    assign outputs[5833] = layer0_outputs[2463];
    assign outputs[5834] = ~((layer0_outputs[2912]) | (layer0_outputs[224]));
    assign outputs[5835] = (layer0_outputs[3837]) & ~(layer0_outputs[4861]);
    assign outputs[5836] = ~(layer0_outputs[5514]);
    assign outputs[5837] = ~(layer0_outputs[5153]);
    assign outputs[5838] = ~(layer0_outputs[4335]);
    assign outputs[5839] = layer0_outputs[7321];
    assign outputs[5840] = ~(layer0_outputs[2580]);
    assign outputs[5841] = ~(layer0_outputs[7560]);
    assign outputs[5842] = ~((layer0_outputs[5061]) ^ (layer0_outputs[4231]));
    assign outputs[5843] = ~(layer0_outputs[3298]);
    assign outputs[5844] = ~((layer0_outputs[7514]) ^ (layer0_outputs[4054]));
    assign outputs[5845] = ~(layer0_outputs[3995]);
    assign outputs[5846] = (layer0_outputs[1653]) ^ (layer0_outputs[784]);
    assign outputs[5847] = (layer0_outputs[6959]) & ~(layer0_outputs[4878]);
    assign outputs[5848] = layer0_outputs[3025];
    assign outputs[5849] = layer0_outputs[6887];
    assign outputs[5850] = layer0_outputs[3117];
    assign outputs[5851] = ~(layer0_outputs[4611]);
    assign outputs[5852] = (layer0_outputs[2602]) & ~(layer0_outputs[1364]);
    assign outputs[5853] = ~(layer0_outputs[5861]);
    assign outputs[5854] = (layer0_outputs[6861]) & ~(layer0_outputs[5889]);
    assign outputs[5855] = ~(layer0_outputs[2746]);
    assign outputs[5856] = ~((layer0_outputs[5383]) & (layer0_outputs[7246]));
    assign outputs[5857] = ~(layer0_outputs[524]);
    assign outputs[5858] = ~((layer0_outputs[2939]) ^ (layer0_outputs[7310]));
    assign outputs[5859] = ~((layer0_outputs[5049]) | (layer0_outputs[1738]));
    assign outputs[5860] = ~(layer0_outputs[2846]);
    assign outputs[5861] = (layer0_outputs[3982]) ^ (layer0_outputs[6077]);
    assign outputs[5862] = (layer0_outputs[6765]) & ~(layer0_outputs[5979]);
    assign outputs[5863] = layer0_outputs[2412];
    assign outputs[5864] = ~(layer0_outputs[1269]);
    assign outputs[5865] = (layer0_outputs[6426]) & ~(layer0_outputs[2579]);
    assign outputs[5866] = layer0_outputs[1994];
    assign outputs[5867] = (layer0_outputs[4164]) ^ (layer0_outputs[1194]);
    assign outputs[5868] = ~((layer0_outputs[6807]) ^ (layer0_outputs[2679]));
    assign outputs[5869] = (layer0_outputs[6510]) & (layer0_outputs[1918]);
    assign outputs[5870] = ~(layer0_outputs[5369]) | (layer0_outputs[303]);
    assign outputs[5871] = ~((layer0_outputs[1422]) & (layer0_outputs[4032]));
    assign outputs[5872] = layer0_outputs[3970];
    assign outputs[5873] = ~((layer0_outputs[275]) ^ (layer0_outputs[1481]));
    assign outputs[5874] = (layer0_outputs[4313]) & (layer0_outputs[223]);
    assign outputs[5875] = layer0_outputs[2670];
    assign outputs[5876] = (layer0_outputs[5634]) & (layer0_outputs[2613]);
    assign outputs[5877] = (layer0_outputs[4708]) & ~(layer0_outputs[5584]);
    assign outputs[5878] = layer0_outputs[3882];
    assign outputs[5879] = (layer0_outputs[2514]) & ~(layer0_outputs[960]);
    assign outputs[5880] = ~(layer0_outputs[5553]);
    assign outputs[5881] = (layer0_outputs[2072]) ^ (layer0_outputs[5340]);
    assign outputs[5882] = ~((layer0_outputs[904]) & (layer0_outputs[1087]));
    assign outputs[5883] = ~((layer0_outputs[720]) ^ (layer0_outputs[421]));
    assign outputs[5884] = (layer0_outputs[1799]) ^ (layer0_outputs[4638]);
    assign outputs[5885] = layer0_outputs[4480];
    assign outputs[5886] = layer0_outputs[2737];
    assign outputs[5887] = ~(layer0_outputs[5320]) | (layer0_outputs[1686]);
    assign outputs[5888] = layer0_outputs[2661];
    assign outputs[5889] = (layer0_outputs[2977]) ^ (layer0_outputs[6368]);
    assign outputs[5890] = layer0_outputs[1123];
    assign outputs[5891] = (layer0_outputs[5055]) & ~(layer0_outputs[6984]);
    assign outputs[5892] = ~(layer0_outputs[1067]) | (layer0_outputs[181]);
    assign outputs[5893] = ~((layer0_outputs[3323]) ^ (layer0_outputs[358]));
    assign outputs[5894] = layer0_outputs[7128];
    assign outputs[5895] = (layer0_outputs[363]) & (layer0_outputs[3899]);
    assign outputs[5896] = ~(layer0_outputs[4361]);
    assign outputs[5897] = ~(layer0_outputs[91]);
    assign outputs[5898] = layer0_outputs[7290];
    assign outputs[5899] = layer0_outputs[6836];
    assign outputs[5900] = (layer0_outputs[6544]) & ~(layer0_outputs[1843]);
    assign outputs[5901] = ~((layer0_outputs[24]) ^ (layer0_outputs[658]));
    assign outputs[5902] = layer0_outputs[4199];
    assign outputs[5903] = ~(layer0_outputs[1423]);
    assign outputs[5904] = (layer0_outputs[2915]) & (layer0_outputs[28]);
    assign outputs[5905] = ~(layer0_outputs[2292]);
    assign outputs[5906] = ~((layer0_outputs[3151]) ^ (layer0_outputs[2761]));
    assign outputs[5907] = ~((layer0_outputs[167]) | (layer0_outputs[4538]));
    assign outputs[5908] = layer0_outputs[5434];
    assign outputs[5909] = layer0_outputs[390];
    assign outputs[5910] = (layer0_outputs[1923]) & ~(layer0_outputs[658]);
    assign outputs[5911] = layer0_outputs[1750];
    assign outputs[5912] = layer0_outputs[3679];
    assign outputs[5913] = layer0_outputs[3862];
    assign outputs[5914] = layer0_outputs[1867];
    assign outputs[5915] = ~(layer0_outputs[1584]);
    assign outputs[5916] = ~((layer0_outputs[4068]) | (layer0_outputs[5314]));
    assign outputs[5917] = ~(layer0_outputs[20]);
    assign outputs[5918] = ~((layer0_outputs[3886]) ^ (layer0_outputs[6263]));
    assign outputs[5919] = layer0_outputs[62];
    assign outputs[5920] = (layer0_outputs[7520]) & ~(layer0_outputs[2589]);
    assign outputs[5921] = ~(layer0_outputs[7116]);
    assign outputs[5922] = ~((layer0_outputs[7433]) | (layer0_outputs[7069]));
    assign outputs[5923] = (layer0_outputs[1172]) & (layer0_outputs[1528]);
    assign outputs[5924] = ~(layer0_outputs[6558]);
    assign outputs[5925] = layer0_outputs[1366];
    assign outputs[5926] = layer0_outputs[5730];
    assign outputs[5927] = 1'b0;
    assign outputs[5928] = layer0_outputs[3649];
    assign outputs[5929] = ~((layer0_outputs[816]) ^ (layer0_outputs[5436]));
    assign outputs[5930] = layer0_outputs[1735];
    assign outputs[5931] = ~(layer0_outputs[2860]);
    assign outputs[5932] = ~(layer0_outputs[2913]);
    assign outputs[5933] = ~((layer0_outputs[2351]) & (layer0_outputs[2763]));
    assign outputs[5934] = (layer0_outputs[1191]) & (layer0_outputs[3206]);
    assign outputs[5935] = (layer0_outputs[28]) & (layer0_outputs[2694]);
    assign outputs[5936] = layer0_outputs[5186];
    assign outputs[5937] = (layer0_outputs[6664]) & ~(layer0_outputs[7514]);
    assign outputs[5938] = layer0_outputs[4968];
    assign outputs[5939] = layer0_outputs[2775];
    assign outputs[5940] = layer0_outputs[4195];
    assign outputs[5941] = (layer0_outputs[6842]) & ~(layer0_outputs[5977]);
    assign outputs[5942] = ~(layer0_outputs[4824]);
    assign outputs[5943] = (layer0_outputs[1138]) | (layer0_outputs[3435]);
    assign outputs[5944] = (layer0_outputs[4132]) | (layer0_outputs[4612]);
    assign outputs[5945] = (layer0_outputs[513]) & ~(layer0_outputs[4388]);
    assign outputs[5946] = ~((layer0_outputs[6155]) & (layer0_outputs[2340]));
    assign outputs[5947] = layer0_outputs[6520];
    assign outputs[5948] = (layer0_outputs[6550]) ^ (layer0_outputs[311]);
    assign outputs[5949] = ~(layer0_outputs[179]);
    assign outputs[5950] = ~(layer0_outputs[3857]);
    assign outputs[5951] = ~((layer0_outputs[4647]) ^ (layer0_outputs[4141]));
    assign outputs[5952] = layer0_outputs[2252];
    assign outputs[5953] = (layer0_outputs[1010]) & ~(layer0_outputs[882]);
    assign outputs[5954] = layer0_outputs[4934];
    assign outputs[5955] = ~(layer0_outputs[5640]);
    assign outputs[5956] = (layer0_outputs[2637]) & ~(layer0_outputs[5633]);
    assign outputs[5957] = (layer0_outputs[6719]) & ~(layer0_outputs[7346]);
    assign outputs[5958] = ~(layer0_outputs[4721]);
    assign outputs[5959] = ~(layer0_outputs[896]);
    assign outputs[5960] = layer0_outputs[5586];
    assign outputs[5961] = ~((layer0_outputs[6095]) ^ (layer0_outputs[5336]));
    assign outputs[5962] = ~(layer0_outputs[6832]);
    assign outputs[5963] = ~((layer0_outputs[7153]) | (layer0_outputs[4220]));
    assign outputs[5964] = ~(layer0_outputs[3885]);
    assign outputs[5965] = ~((layer0_outputs[7428]) ^ (layer0_outputs[3606]));
    assign outputs[5966] = (layer0_outputs[2295]) & ~(layer0_outputs[3700]);
    assign outputs[5967] = layer0_outputs[1632];
    assign outputs[5968] = layer0_outputs[3043];
    assign outputs[5969] = ~((layer0_outputs[4331]) | (layer0_outputs[5171]));
    assign outputs[5970] = ~((layer0_outputs[4046]) | (layer0_outputs[3881]));
    assign outputs[5971] = ~(layer0_outputs[2014]);
    assign outputs[5972] = ~(layer0_outputs[6827]);
    assign outputs[5973] = ~((layer0_outputs[6290]) | (layer0_outputs[1458]));
    assign outputs[5974] = (layer0_outputs[4705]) & ~(layer0_outputs[2243]);
    assign outputs[5975] = ~(layer0_outputs[7502]);
    assign outputs[5976] = ~((layer0_outputs[5779]) ^ (layer0_outputs[3044]));
    assign outputs[5977] = (layer0_outputs[6120]) ^ (layer0_outputs[5227]);
    assign outputs[5978] = (layer0_outputs[5810]) & (layer0_outputs[4066]);
    assign outputs[5979] = ~(layer0_outputs[4376]);
    assign outputs[5980] = ~(layer0_outputs[5396]);
    assign outputs[5981] = ~(layer0_outputs[6410]);
    assign outputs[5982] = layer0_outputs[391];
    assign outputs[5983] = (layer0_outputs[6929]) & ~(layer0_outputs[6675]);
    assign outputs[5984] = ~(layer0_outputs[3281]);
    assign outputs[5985] = ~(layer0_outputs[1603]);
    assign outputs[5986] = ~(layer0_outputs[4830]);
    assign outputs[5987] = (layer0_outputs[3575]) ^ (layer0_outputs[2648]);
    assign outputs[5988] = 1'b0;
    assign outputs[5989] = 1'b0;
    assign outputs[5990] = layer0_outputs[2474];
    assign outputs[5991] = layer0_outputs[934];
    assign outputs[5992] = (layer0_outputs[430]) & (layer0_outputs[6300]);
    assign outputs[5993] = layer0_outputs[7414];
    assign outputs[5994] = (layer0_outputs[674]) & ~(layer0_outputs[5602]);
    assign outputs[5995] = ~((layer0_outputs[7267]) ^ (layer0_outputs[1401]));
    assign outputs[5996] = ~(layer0_outputs[3572]) | (layer0_outputs[3362]);
    assign outputs[5997] = (layer0_outputs[3473]) ^ (layer0_outputs[4144]);
    assign outputs[5998] = (layer0_outputs[6539]) & ~(layer0_outputs[7329]);
    assign outputs[5999] = layer0_outputs[4752];
    assign outputs[6000] = (layer0_outputs[6777]) & ~(layer0_outputs[7285]);
    assign outputs[6001] = (layer0_outputs[261]) & (layer0_outputs[4564]);
    assign outputs[6002] = (layer0_outputs[4991]) & ~(layer0_outputs[7662]);
    assign outputs[6003] = ~((layer0_outputs[2035]) | (layer0_outputs[2442]));
    assign outputs[6004] = ~(layer0_outputs[6119]);
    assign outputs[6005] = ~(layer0_outputs[3552]);
    assign outputs[6006] = layer0_outputs[7585];
    assign outputs[6007] = ~((layer0_outputs[7486]) | (layer0_outputs[6093]));
    assign outputs[6008] = (layer0_outputs[6160]) & ~(layer0_outputs[5156]);
    assign outputs[6009] = (layer0_outputs[7059]) ^ (layer0_outputs[1466]);
    assign outputs[6010] = ~(layer0_outputs[6477]) | (layer0_outputs[277]);
    assign outputs[6011] = ~((layer0_outputs[491]) ^ (layer0_outputs[6378]));
    assign outputs[6012] = layer0_outputs[4799];
    assign outputs[6013] = (layer0_outputs[1522]) ^ (layer0_outputs[5765]);
    assign outputs[6014] = (layer0_outputs[2383]) ^ (layer0_outputs[3557]);
    assign outputs[6015] = layer0_outputs[5942];
    assign outputs[6016] = (layer0_outputs[5984]) | (layer0_outputs[2836]);
    assign outputs[6017] = (layer0_outputs[1692]) & ~(layer0_outputs[4340]);
    assign outputs[6018] = ~(layer0_outputs[1065]);
    assign outputs[6019] = (layer0_outputs[1469]) & ~(layer0_outputs[1644]);
    assign outputs[6020] = ~(layer0_outputs[2365]);
    assign outputs[6021] = (layer0_outputs[5796]) & ~(layer0_outputs[2239]);
    assign outputs[6022] = 1'b1;
    assign outputs[6023] = ~(layer0_outputs[689]);
    assign outputs[6024] = (layer0_outputs[1925]) ^ (layer0_outputs[4711]);
    assign outputs[6025] = (layer0_outputs[3887]) & (layer0_outputs[1776]);
    assign outputs[6026] = ~(layer0_outputs[2896]) | (layer0_outputs[519]);
    assign outputs[6027] = (layer0_outputs[2279]) & (layer0_outputs[5002]);
    assign outputs[6028] = layer0_outputs[7633];
    assign outputs[6029] = layer0_outputs[3933];
    assign outputs[6030] = (layer0_outputs[1227]) ^ (layer0_outputs[4887]);
    assign outputs[6031] = (layer0_outputs[3954]) ^ (layer0_outputs[2518]);
    assign outputs[6032] = (layer0_outputs[6208]) & ~(layer0_outputs[7087]);
    assign outputs[6033] = (layer0_outputs[1312]) & ~(layer0_outputs[1228]);
    assign outputs[6034] = ~((layer0_outputs[5335]) | (layer0_outputs[1236]));
    assign outputs[6035] = layer0_outputs[1655];
    assign outputs[6036] = (layer0_outputs[3895]) ^ (layer0_outputs[3826]);
    assign outputs[6037] = layer0_outputs[3688];
    assign outputs[6038] = (layer0_outputs[4987]) ^ (layer0_outputs[625]);
    assign outputs[6039] = ~((layer0_outputs[4054]) ^ (layer0_outputs[3179]));
    assign outputs[6040] = layer0_outputs[4762];
    assign outputs[6041] = (layer0_outputs[430]) & (layer0_outputs[5036]);
    assign outputs[6042] = ~(layer0_outputs[3986]);
    assign outputs[6043] = ~((layer0_outputs[6283]) & (layer0_outputs[3369]));
    assign outputs[6044] = (layer0_outputs[6426]) & ~(layer0_outputs[3258]);
    assign outputs[6045] = ~(layer0_outputs[1725]);
    assign outputs[6046] = ~(layer0_outputs[6247]);
    assign outputs[6047] = (layer0_outputs[1790]) & ~(layer0_outputs[2331]);
    assign outputs[6048] = (layer0_outputs[6262]) ^ (layer0_outputs[6005]);
    assign outputs[6049] = layer0_outputs[3266];
    assign outputs[6050] = ~(layer0_outputs[5766]) | (layer0_outputs[1392]);
    assign outputs[6051] = layer0_outputs[1492];
    assign outputs[6052] = (layer0_outputs[4801]) ^ (layer0_outputs[449]);
    assign outputs[6053] = ~((layer0_outputs[3781]) ^ (layer0_outputs[1623]));
    assign outputs[6054] = ~(layer0_outputs[3134]) | (layer0_outputs[555]);
    assign outputs[6055] = ~((layer0_outputs[3705]) & (layer0_outputs[773]));
    assign outputs[6056] = layer0_outputs[6812];
    assign outputs[6057] = layer0_outputs[6480];
    assign outputs[6058] = layer0_outputs[1171];
    assign outputs[6059] = (layer0_outputs[6365]) & ~(layer0_outputs[4068]);
    assign outputs[6060] = (layer0_outputs[645]) & (layer0_outputs[7351]);
    assign outputs[6061] = ~(layer0_outputs[1645]);
    assign outputs[6062] = ~(layer0_outputs[334]);
    assign outputs[6063] = ~(layer0_outputs[5239]);
    assign outputs[6064] = layer0_outputs[4989];
    assign outputs[6065] = ~(layer0_outputs[7430]);
    assign outputs[6066] = (layer0_outputs[4714]) | (layer0_outputs[1875]);
    assign outputs[6067] = ~((layer0_outputs[2870]) ^ (layer0_outputs[4547]));
    assign outputs[6068] = (layer0_outputs[2687]) ^ (layer0_outputs[792]);
    assign outputs[6069] = layer0_outputs[219];
    assign outputs[6070] = ~(layer0_outputs[2147]);
    assign outputs[6071] = layer0_outputs[1121];
    assign outputs[6072] = (layer0_outputs[533]) & ~(layer0_outputs[2751]);
    assign outputs[6073] = (layer0_outputs[3561]) ^ (layer0_outputs[2859]);
    assign outputs[6074] = ~(layer0_outputs[7521]) | (layer0_outputs[1320]);
    assign outputs[6075] = layer0_outputs[1276];
    assign outputs[6076] = ~((layer0_outputs[2947]) ^ (layer0_outputs[2891]));
    assign outputs[6077] = (layer0_outputs[2015]) ^ (layer0_outputs[4508]);
    assign outputs[6078] = layer0_outputs[7531];
    assign outputs[6079] = (layer0_outputs[3742]) & ~(layer0_outputs[6974]);
    assign outputs[6080] = ~((layer0_outputs[5919]) & (layer0_outputs[125]));
    assign outputs[6081] = ~(layer0_outputs[5556]);
    assign outputs[6082] = ~(layer0_outputs[3175]);
    assign outputs[6083] = layer0_outputs[4070];
    assign outputs[6084] = ~(layer0_outputs[3221]);
    assign outputs[6085] = layer0_outputs[7190];
    assign outputs[6086] = ~((layer0_outputs[1822]) ^ (layer0_outputs[4207]));
    assign outputs[6087] = ~(layer0_outputs[1279]);
    assign outputs[6088] = (layer0_outputs[3313]) & ~(layer0_outputs[6618]);
    assign outputs[6089] = (layer0_outputs[1200]) ^ (layer0_outputs[1109]);
    assign outputs[6090] = layer0_outputs[429];
    assign outputs[6091] = (layer0_outputs[6363]) & ~(layer0_outputs[5034]);
    assign outputs[6092] = ~((layer0_outputs[6151]) | (layer0_outputs[7671]));
    assign outputs[6093] = ~((layer0_outputs[2495]) | (layer0_outputs[6272]));
    assign outputs[6094] = (layer0_outputs[1777]) & ~(layer0_outputs[2177]);
    assign outputs[6095] = (layer0_outputs[5318]) & ~(layer0_outputs[3316]);
    assign outputs[6096] = ~(layer0_outputs[1921]) | (layer0_outputs[7279]);
    assign outputs[6097] = ~(layer0_outputs[195]);
    assign outputs[6098] = ~((layer0_outputs[2851]) ^ (layer0_outputs[4816]));
    assign outputs[6099] = (layer0_outputs[307]) & ~(layer0_outputs[7171]);
    assign outputs[6100] = (layer0_outputs[2228]) ^ (layer0_outputs[6910]);
    assign outputs[6101] = (layer0_outputs[4358]) ^ (layer0_outputs[3566]);
    assign outputs[6102] = layer0_outputs[7584];
    assign outputs[6103] = layer0_outputs[5990];
    assign outputs[6104] = (layer0_outputs[5931]) ^ (layer0_outputs[5368]);
    assign outputs[6105] = ~(layer0_outputs[5830]);
    assign outputs[6106] = ~(layer0_outputs[4234]);
    assign outputs[6107] = ~((layer0_outputs[5482]) | (layer0_outputs[7235]));
    assign outputs[6108] = (layer0_outputs[1244]) ^ (layer0_outputs[7661]);
    assign outputs[6109] = ~(layer0_outputs[2557]);
    assign outputs[6110] = (layer0_outputs[2560]) & ~(layer0_outputs[5429]);
    assign outputs[6111] = ~(layer0_outputs[2322]);
    assign outputs[6112] = layer0_outputs[3491];
    assign outputs[6113] = layer0_outputs[3875];
    assign outputs[6114] = ~(layer0_outputs[2224]);
    assign outputs[6115] = (layer0_outputs[3557]) & (layer0_outputs[1001]);
    assign outputs[6116] = ~((layer0_outputs[3322]) ^ (layer0_outputs[3345]));
    assign outputs[6117] = (layer0_outputs[626]) ^ (layer0_outputs[6427]);
    assign outputs[6118] = (layer0_outputs[3548]) & ~(layer0_outputs[744]);
    assign outputs[6119] = layer0_outputs[5349];
    assign outputs[6120] = ~((layer0_outputs[814]) ^ (layer0_outputs[5309]));
    assign outputs[6121] = ~((layer0_outputs[5641]) ^ (layer0_outputs[2419]));
    assign outputs[6122] = (layer0_outputs[1923]) & ~(layer0_outputs[4911]);
    assign outputs[6123] = (layer0_outputs[6143]) & ~(layer0_outputs[4308]);
    assign outputs[6124] = layer0_outputs[1467];
    assign outputs[6125] = layer0_outputs[2959];
    assign outputs[6126] = layer0_outputs[1993];
    assign outputs[6127] = ~(layer0_outputs[6349]);
    assign outputs[6128] = (layer0_outputs[4805]) & (layer0_outputs[1354]);
    assign outputs[6129] = ~((layer0_outputs[4605]) | (layer0_outputs[1374]));
    assign outputs[6130] = ~(layer0_outputs[3628]);
    assign outputs[6131] = ~(layer0_outputs[2126]);
    assign outputs[6132] = (layer0_outputs[2636]) & ~(layer0_outputs[4722]);
    assign outputs[6133] = (layer0_outputs[514]) ^ (layer0_outputs[3219]);
    assign outputs[6134] = (layer0_outputs[3096]) ^ (layer0_outputs[4627]);
    assign outputs[6135] = layer0_outputs[2552];
    assign outputs[6136] = (layer0_outputs[7669]) & ~(layer0_outputs[1261]);
    assign outputs[6137] = ~(layer0_outputs[220]);
    assign outputs[6138] = layer0_outputs[3043];
    assign outputs[6139] = layer0_outputs[1826];
    assign outputs[6140] = ~((layer0_outputs[4545]) ^ (layer0_outputs[5562]));
    assign outputs[6141] = layer0_outputs[2908];
    assign outputs[6142] = (layer0_outputs[4571]) & ~(layer0_outputs[274]);
    assign outputs[6143] = layer0_outputs[870];
    assign outputs[6144] = (layer0_outputs[83]) ^ (layer0_outputs[6948]);
    assign outputs[6145] = (layer0_outputs[4977]) ^ (layer0_outputs[3915]);
    assign outputs[6146] = layer0_outputs[5856];
    assign outputs[6147] = ~((layer0_outputs[4374]) & (layer0_outputs[282]));
    assign outputs[6148] = (layer0_outputs[6511]) ^ (layer0_outputs[1892]);
    assign outputs[6149] = layer0_outputs[7083];
    assign outputs[6150] = layer0_outputs[2426];
    assign outputs[6151] = (layer0_outputs[501]) & ~(layer0_outputs[450]);
    assign outputs[6152] = layer0_outputs[3953];
    assign outputs[6153] = ~(layer0_outputs[7271]);
    assign outputs[6154] = ~(layer0_outputs[3638]);
    assign outputs[6155] = ~(layer0_outputs[6323]) | (layer0_outputs[4482]);
    assign outputs[6156] = ~(layer0_outputs[1262]) | (layer0_outputs[4708]);
    assign outputs[6157] = layer0_outputs[1500];
    assign outputs[6158] = layer0_outputs[2305];
    assign outputs[6159] = ~((layer0_outputs[6213]) & (layer0_outputs[5855]));
    assign outputs[6160] = (layer0_outputs[5849]) ^ (layer0_outputs[3974]);
    assign outputs[6161] = (layer0_outputs[6042]) | (layer0_outputs[5874]);
    assign outputs[6162] = (layer0_outputs[820]) ^ (layer0_outputs[7058]);
    assign outputs[6163] = (layer0_outputs[6957]) & ~(layer0_outputs[1651]);
    assign outputs[6164] = layer0_outputs[1743];
    assign outputs[6165] = (layer0_outputs[614]) & (layer0_outputs[3620]);
    assign outputs[6166] = ~(layer0_outputs[262]);
    assign outputs[6167] = ~(layer0_outputs[2874]) | (layer0_outputs[5814]);
    assign outputs[6168] = ~((layer0_outputs[5135]) ^ (layer0_outputs[2341]));
    assign outputs[6169] = (layer0_outputs[5546]) & ~(layer0_outputs[4346]);
    assign outputs[6170] = (layer0_outputs[3644]) ^ (layer0_outputs[2520]);
    assign outputs[6171] = ~((layer0_outputs[3348]) ^ (layer0_outputs[3837]));
    assign outputs[6172] = ~(layer0_outputs[5639]) | (layer0_outputs[6645]);
    assign outputs[6173] = ~(layer0_outputs[6900]) | (layer0_outputs[4660]);
    assign outputs[6174] = ~(layer0_outputs[823]);
    assign outputs[6175] = ~((layer0_outputs[3092]) ^ (layer0_outputs[74]));
    assign outputs[6176] = ~(layer0_outputs[5651]);
    assign outputs[6177] = layer0_outputs[4751];
    assign outputs[6178] = layer0_outputs[171];
    assign outputs[6179] = ~(layer0_outputs[1610]);
    assign outputs[6180] = ~(layer0_outputs[2679]);
    assign outputs[6181] = ~(layer0_outputs[988]) | (layer0_outputs[4901]);
    assign outputs[6182] = ~((layer0_outputs[6971]) ^ (layer0_outputs[5766]));
    assign outputs[6183] = ~(layer0_outputs[4844]);
    assign outputs[6184] = ~(layer0_outputs[3045]);
    assign outputs[6185] = ~((layer0_outputs[3249]) ^ (layer0_outputs[4644]));
    assign outputs[6186] = ~(layer0_outputs[6640]) | (layer0_outputs[2601]);
    assign outputs[6187] = (layer0_outputs[3425]) ^ (layer0_outputs[5458]);
    assign outputs[6188] = ~(layer0_outputs[1647]);
    assign outputs[6189] = (layer0_outputs[2194]) & (layer0_outputs[207]);
    assign outputs[6190] = ~(layer0_outputs[2622]) | (layer0_outputs[1892]);
    assign outputs[6191] = ~(layer0_outputs[4749]) | (layer0_outputs[591]);
    assign outputs[6192] = ~(layer0_outputs[1561]);
    assign outputs[6193] = layer0_outputs[7414];
    assign outputs[6194] = ~(layer0_outputs[7341]);
    assign outputs[6195] = (layer0_outputs[5033]) & ~(layer0_outputs[6580]);
    assign outputs[6196] = ~((layer0_outputs[86]) & (layer0_outputs[6816]));
    assign outputs[6197] = layer0_outputs[601];
    assign outputs[6198] = ~(layer0_outputs[5626]);
    assign outputs[6199] = (layer0_outputs[2661]) ^ (layer0_outputs[6174]);
    assign outputs[6200] = ~((layer0_outputs[4567]) ^ (layer0_outputs[943]));
    assign outputs[6201] = ~(layer0_outputs[1093]);
    assign outputs[6202] = (layer0_outputs[1635]) & (layer0_outputs[705]);
    assign outputs[6203] = (layer0_outputs[1992]) | (layer0_outputs[5155]);
    assign outputs[6204] = layer0_outputs[5084];
    assign outputs[6205] = ~((layer0_outputs[2899]) ^ (layer0_outputs[4669]));
    assign outputs[6206] = ~((layer0_outputs[568]) ^ (layer0_outputs[7070]));
    assign outputs[6207] = ~((layer0_outputs[5685]) ^ (layer0_outputs[7628]));
    assign outputs[6208] = ~(layer0_outputs[1888]) | (layer0_outputs[5965]);
    assign outputs[6209] = (layer0_outputs[4286]) ^ (layer0_outputs[1696]);
    assign outputs[6210] = layer0_outputs[3365];
    assign outputs[6211] = layer0_outputs[7333];
    assign outputs[6212] = layer0_outputs[5802];
    assign outputs[6213] = ~(layer0_outputs[5377]);
    assign outputs[6214] = ~(layer0_outputs[3102]);
    assign outputs[6215] = ~((layer0_outputs[1198]) ^ (layer0_outputs[1141]));
    assign outputs[6216] = ~(layer0_outputs[4475]);
    assign outputs[6217] = ~(layer0_outputs[4835]) | (layer0_outputs[4079]);
    assign outputs[6218] = (layer0_outputs[5099]) & ~(layer0_outputs[7550]);
    assign outputs[6219] = ~((layer0_outputs[4970]) ^ (layer0_outputs[7135]));
    assign outputs[6220] = ~(layer0_outputs[5050]);
    assign outputs[6221] = (layer0_outputs[4840]) ^ (layer0_outputs[3682]);
    assign outputs[6222] = (layer0_outputs[4126]) & ~(layer0_outputs[7095]);
    assign outputs[6223] = ~(layer0_outputs[324]);
    assign outputs[6224] = (layer0_outputs[987]) ^ (layer0_outputs[6750]);
    assign outputs[6225] = ~((layer0_outputs[926]) ^ (layer0_outputs[6728]));
    assign outputs[6226] = (layer0_outputs[2631]) & ~(layer0_outputs[3185]);
    assign outputs[6227] = ~(layer0_outputs[7581]) | (layer0_outputs[2132]);
    assign outputs[6228] = (layer0_outputs[4166]) | (layer0_outputs[3541]);
    assign outputs[6229] = ~((layer0_outputs[216]) & (layer0_outputs[6585]));
    assign outputs[6230] = (layer0_outputs[1588]) ^ (layer0_outputs[1996]);
    assign outputs[6231] = (layer0_outputs[3964]) & (layer0_outputs[5754]);
    assign outputs[6232] = ~(layer0_outputs[6318]) | (layer0_outputs[6518]);
    assign outputs[6233] = layer0_outputs[3590];
    assign outputs[6234] = layer0_outputs[6124];
    assign outputs[6235] = layer0_outputs[7218];
    assign outputs[6236] = ~(layer0_outputs[5602]) | (layer0_outputs[4386]);
    assign outputs[6237] = ~(layer0_outputs[2791]) | (layer0_outputs[1772]);
    assign outputs[6238] = ~(layer0_outputs[4086]) | (layer0_outputs[2256]);
    assign outputs[6239] = layer0_outputs[884];
    assign outputs[6240] = (layer0_outputs[1107]) ^ (layer0_outputs[840]);
    assign outputs[6241] = (layer0_outputs[1759]) & ~(layer0_outputs[2309]);
    assign outputs[6242] = ~((layer0_outputs[3026]) | (layer0_outputs[2185]));
    assign outputs[6243] = layer0_outputs[783];
    assign outputs[6244] = (layer0_outputs[1729]) & ~(layer0_outputs[5328]);
    assign outputs[6245] = (layer0_outputs[5825]) & ~(layer0_outputs[1611]);
    assign outputs[6246] = (layer0_outputs[5841]) & (layer0_outputs[5251]);
    assign outputs[6247] = ~((layer0_outputs[6389]) & (layer0_outputs[7280]));
    assign outputs[6248] = layer0_outputs[2536];
    assign outputs[6249] = (layer0_outputs[1176]) ^ (layer0_outputs[6465]);
    assign outputs[6250] = layer0_outputs[6891];
    assign outputs[6251] = ~((layer0_outputs[5204]) ^ (layer0_outputs[4659]));
    assign outputs[6252] = (layer0_outputs[151]) ^ (layer0_outputs[3427]);
    assign outputs[6253] = ~(layer0_outputs[785]);
    assign outputs[6254] = (layer0_outputs[6708]) | (layer0_outputs[5261]);
    assign outputs[6255] = ~(layer0_outputs[6913]);
    assign outputs[6256] = ~(layer0_outputs[6614]);
    assign outputs[6257] = layer0_outputs[1339];
    assign outputs[6258] = layer0_outputs[3468];
    assign outputs[6259] = ~((layer0_outputs[3002]) & (layer0_outputs[3926]));
    assign outputs[6260] = (layer0_outputs[6617]) & ~(layer0_outputs[6266]);
    assign outputs[6261] = (layer0_outputs[6779]) & ~(layer0_outputs[6428]);
    assign outputs[6262] = (layer0_outputs[1298]) & ~(layer0_outputs[5557]);
    assign outputs[6263] = (layer0_outputs[3428]) ^ (layer0_outputs[4458]);
    assign outputs[6264] = ~(layer0_outputs[7610]);
    assign outputs[6265] = (layer0_outputs[3220]) ^ (layer0_outputs[6527]);
    assign outputs[6266] = ~((layer0_outputs[6547]) & (layer0_outputs[1274]));
    assign outputs[6267] = layer0_outputs[3607];
    assign outputs[6268] = (layer0_outputs[1002]) ^ (layer0_outputs[5719]);
    assign outputs[6269] = ~(layer0_outputs[2140]);
    assign outputs[6270] = ~(layer0_outputs[3697]);
    assign outputs[6271] = (layer0_outputs[7664]) & ~(layer0_outputs[5926]);
    assign outputs[6272] = ~(layer0_outputs[4619]);
    assign outputs[6273] = ~(layer0_outputs[3795]) | (layer0_outputs[7604]);
    assign outputs[6274] = ~(layer0_outputs[5682]);
    assign outputs[6275] = ~((layer0_outputs[1680]) | (layer0_outputs[2756]));
    assign outputs[6276] = ~(layer0_outputs[551]);
    assign outputs[6277] = ~(layer0_outputs[6851]) | (layer0_outputs[844]);
    assign outputs[6278] = layer0_outputs[4062];
    assign outputs[6279] = ~(layer0_outputs[40]);
    assign outputs[6280] = layer0_outputs[6748];
    assign outputs[6281] = ~((layer0_outputs[6651]) ^ (layer0_outputs[6228]));
    assign outputs[6282] = ~(layer0_outputs[5139]);
    assign outputs[6283] = ~(layer0_outputs[5235]) | (layer0_outputs[2842]);
    assign outputs[6284] = ~((layer0_outputs[839]) ^ (layer0_outputs[6622]));
    assign outputs[6285] = ~(layer0_outputs[2440]);
    assign outputs[6286] = ~(layer0_outputs[1201]) | (layer0_outputs[1420]);
    assign outputs[6287] = ~(layer0_outputs[2015]);
    assign outputs[6288] = (layer0_outputs[128]) | (layer0_outputs[5277]);
    assign outputs[6289] = ~((layer0_outputs[4596]) | (layer0_outputs[3725]));
    assign outputs[6290] = layer0_outputs[6649];
    assign outputs[6291] = layer0_outputs[7300];
    assign outputs[6292] = (layer0_outputs[5267]) | (layer0_outputs[4303]);
    assign outputs[6293] = ~(layer0_outputs[6972]) | (layer0_outputs[5895]);
    assign outputs[6294] = layer0_outputs[5261];
    assign outputs[6295] = ~(layer0_outputs[6955]) | (layer0_outputs[4]);
    assign outputs[6296] = ~(layer0_outputs[5654]);
    assign outputs[6297] = (layer0_outputs[4438]) ^ (layer0_outputs[5993]);
    assign outputs[6298] = ~(layer0_outputs[7096]);
    assign outputs[6299] = layer0_outputs[6562];
    assign outputs[6300] = ~(layer0_outputs[2668]) | (layer0_outputs[6846]);
    assign outputs[6301] = ~(layer0_outputs[6780]);
    assign outputs[6302] = layer0_outputs[5920];
    assign outputs[6303] = layer0_outputs[1227];
    assign outputs[6304] = ~(layer0_outputs[2490]);
    assign outputs[6305] = (layer0_outputs[2406]) & (layer0_outputs[3523]);
    assign outputs[6306] = (layer0_outputs[7356]) ^ (layer0_outputs[6494]);
    assign outputs[6307] = ~(layer0_outputs[3880]);
    assign outputs[6308] = (layer0_outputs[2657]) & ~(layer0_outputs[4629]);
    assign outputs[6309] = (layer0_outputs[1618]) ^ (layer0_outputs[6796]);
    assign outputs[6310] = ~(layer0_outputs[664]);
    assign outputs[6311] = ~(layer0_outputs[1948]);
    assign outputs[6312] = ~(layer0_outputs[7359]);
    assign outputs[6313] = ~((layer0_outputs[2868]) ^ (layer0_outputs[697]));
    assign outputs[6314] = layer0_outputs[3405];
    assign outputs[6315] = ~((layer0_outputs[1331]) & (layer0_outputs[2820]));
    assign outputs[6316] = (layer0_outputs[6701]) ^ (layer0_outputs[5822]);
    assign outputs[6317] = ~((layer0_outputs[4994]) ^ (layer0_outputs[1303]));
    assign outputs[6318] = (layer0_outputs[3926]) & ~(layer0_outputs[4910]);
    assign outputs[6319] = ~(layer0_outputs[1835]) | (layer0_outputs[4942]);
    assign outputs[6320] = ~((layer0_outputs[5516]) ^ (layer0_outputs[3095]));
    assign outputs[6321] = ~((layer0_outputs[941]) ^ (layer0_outputs[1663]));
    assign outputs[6322] = ~((layer0_outputs[7207]) ^ (layer0_outputs[2185]));
    assign outputs[6323] = (layer0_outputs[7350]) & ~(layer0_outputs[3653]);
    assign outputs[6324] = ~(layer0_outputs[4590]);
    assign outputs[6325] = ~(layer0_outputs[5595]);
    assign outputs[6326] = layer0_outputs[4384];
    assign outputs[6327] = (layer0_outputs[761]) ^ (layer0_outputs[128]);
    assign outputs[6328] = layer0_outputs[1383];
    assign outputs[6329] = ~((layer0_outputs[5497]) ^ (layer0_outputs[1165]));
    assign outputs[6330] = ~(layer0_outputs[3156]) | (layer0_outputs[1372]);
    assign outputs[6331] = ~(layer0_outputs[3545]);
    assign outputs[6332] = ~((layer0_outputs[7015]) | (layer0_outputs[1619]));
    assign outputs[6333] = (layer0_outputs[5287]) ^ (layer0_outputs[599]);
    assign outputs[6334] = (layer0_outputs[3469]) ^ (layer0_outputs[4540]);
    assign outputs[6335] = layer0_outputs[4838];
    assign outputs[6336] = layer0_outputs[3520];
    assign outputs[6337] = ~(layer0_outputs[2222]);
    assign outputs[6338] = ~((layer0_outputs[5397]) ^ (layer0_outputs[7099]));
    assign outputs[6339] = layer0_outputs[7112];
    assign outputs[6340] = (layer0_outputs[5638]) ^ (layer0_outputs[73]);
    assign outputs[6341] = (layer0_outputs[2351]) ^ (layer0_outputs[3154]);
    assign outputs[6342] = (layer0_outputs[4344]) | (layer0_outputs[1234]);
    assign outputs[6343] = ~(layer0_outputs[1682]);
    assign outputs[6344] = ~((layer0_outputs[7334]) | (layer0_outputs[1049]));
    assign outputs[6345] = (layer0_outputs[3462]) | (layer0_outputs[3916]);
    assign outputs[6346] = ~(layer0_outputs[1180]);
    assign outputs[6347] = ~(layer0_outputs[5922]);
    assign outputs[6348] = (layer0_outputs[1556]) & ~(layer0_outputs[4878]);
    assign outputs[6349] = ~((layer0_outputs[1858]) ^ (layer0_outputs[5714]));
    assign outputs[6350] = ~(layer0_outputs[5985]);
    assign outputs[6351] = ~((layer0_outputs[7248]) ^ (layer0_outputs[5789]));
    assign outputs[6352] = (layer0_outputs[6373]) ^ (layer0_outputs[3935]);
    assign outputs[6353] = layer0_outputs[4656];
    assign outputs[6354] = ~((layer0_outputs[4893]) | (layer0_outputs[3434]));
    assign outputs[6355] = ~(layer0_outputs[3889]);
    assign outputs[6356] = ~(layer0_outputs[2141]);
    assign outputs[6357] = (layer0_outputs[1293]) ^ (layer0_outputs[511]);
    assign outputs[6358] = ~(layer0_outputs[7077]);
    assign outputs[6359] = layer0_outputs[4964];
    assign outputs[6360] = ~((layer0_outputs[706]) ^ (layer0_outputs[530]));
    assign outputs[6361] = ~((layer0_outputs[6361]) | (layer0_outputs[3056]));
    assign outputs[6362] = (layer0_outputs[4559]) ^ (layer0_outputs[3584]);
    assign outputs[6363] = ~(layer0_outputs[3138]);
    assign outputs[6364] = ~((layer0_outputs[2568]) ^ (layer0_outputs[7304]));
    assign outputs[6365] = ~(layer0_outputs[862]) | (layer0_outputs[6142]);
    assign outputs[6366] = (layer0_outputs[6600]) ^ (layer0_outputs[3514]);
    assign outputs[6367] = (layer0_outputs[3958]) ^ (layer0_outputs[3157]);
    assign outputs[6368] = (layer0_outputs[5238]) & ~(layer0_outputs[3934]);
    assign outputs[6369] = (layer0_outputs[2976]) & (layer0_outputs[3528]);
    assign outputs[6370] = ~((layer0_outputs[6423]) ^ (layer0_outputs[4649]));
    assign outputs[6371] = layer0_outputs[6940];
    assign outputs[6372] = (layer0_outputs[3102]) ^ (layer0_outputs[2888]);
    assign outputs[6373] = ~(layer0_outputs[6848]);
    assign outputs[6374] = ~(layer0_outputs[5680]);
    assign outputs[6375] = (layer0_outputs[3407]) ^ (layer0_outputs[1911]);
    assign outputs[6376] = ~((layer0_outputs[5362]) ^ (layer0_outputs[854]));
    assign outputs[6377] = ~(layer0_outputs[5108]);
    assign outputs[6378] = ~(layer0_outputs[1029]);
    assign outputs[6379] = ~((layer0_outputs[6592]) & (layer0_outputs[3421]));
    assign outputs[6380] = ~((layer0_outputs[3197]) ^ (layer0_outputs[248]));
    assign outputs[6381] = ~(layer0_outputs[7049]) | (layer0_outputs[5531]);
    assign outputs[6382] = ~(layer0_outputs[7456]);
    assign outputs[6383] = (layer0_outputs[2230]) ^ (layer0_outputs[2007]);
    assign outputs[6384] = (layer0_outputs[396]) & ~(layer0_outputs[1061]);
    assign outputs[6385] = ~((layer0_outputs[3063]) ^ (layer0_outputs[4438]));
    assign outputs[6386] = ~(layer0_outputs[7462]);
    assign outputs[6387] = ~(layer0_outputs[4755]);
    assign outputs[6388] = ~(layer0_outputs[4600]) | (layer0_outputs[5299]);
    assign outputs[6389] = (layer0_outputs[1291]) & (layer0_outputs[3449]);
    assign outputs[6390] = (layer0_outputs[6579]) & ~(layer0_outputs[3198]);
    assign outputs[6391] = ~(layer0_outputs[7005]) | (layer0_outputs[6567]);
    assign outputs[6392] = layer0_outputs[3900];
    assign outputs[6393] = ~((layer0_outputs[594]) ^ (layer0_outputs[1793]));
    assign outputs[6394] = (layer0_outputs[1232]) ^ (layer0_outputs[4606]);
    assign outputs[6395] = (layer0_outputs[5740]) ^ (layer0_outputs[6383]);
    assign outputs[6396] = (layer0_outputs[4772]) | (layer0_outputs[2558]);
    assign outputs[6397] = ~(layer0_outputs[238]);
    assign outputs[6398] = layer0_outputs[2046];
    assign outputs[6399] = ~(layer0_outputs[1674]);
    assign outputs[6400] = ~(layer0_outputs[7522]);
    assign outputs[6401] = (layer0_outputs[4965]) & ~(layer0_outputs[1514]);
    assign outputs[6402] = layer0_outputs[7229];
    assign outputs[6403] = layer0_outputs[3671];
    assign outputs[6404] = (layer0_outputs[2930]) & ~(layer0_outputs[5122]);
    assign outputs[6405] = (layer0_outputs[6288]) | (layer0_outputs[3819]);
    assign outputs[6406] = (layer0_outputs[1400]) & ~(layer0_outputs[5929]);
    assign outputs[6407] = ~(layer0_outputs[6283]);
    assign outputs[6408] = layer0_outputs[4110];
    assign outputs[6409] = ~(layer0_outputs[4161]);
    assign outputs[6410] = (layer0_outputs[3872]) ^ (layer0_outputs[6973]);
    assign outputs[6411] = 1'b1;
    assign outputs[6412] = ~(layer0_outputs[585]);
    assign outputs[6413] = layer0_outputs[6329];
    assign outputs[6414] = (layer0_outputs[5114]) & (layer0_outputs[5840]);
    assign outputs[6415] = layer0_outputs[6061];
    assign outputs[6416] = ~(layer0_outputs[7384]);
    assign outputs[6417] = layer0_outputs[4466];
    assign outputs[6418] = ~(layer0_outputs[3129]);
    assign outputs[6419] = layer0_outputs[7158];
    assign outputs[6420] = ~(layer0_outputs[4367]);
    assign outputs[6421] = layer0_outputs[5668];
    assign outputs[6422] = ~(layer0_outputs[5697]);
    assign outputs[6423] = (layer0_outputs[2435]) ^ (layer0_outputs[3802]);
    assign outputs[6424] = (layer0_outputs[2567]) ^ (layer0_outputs[1323]);
    assign outputs[6425] = layer0_outputs[5039];
    assign outputs[6426] = ~((layer0_outputs[4498]) ^ (layer0_outputs[7439]));
    assign outputs[6427] = (layer0_outputs[3816]) ^ (layer0_outputs[7073]);
    assign outputs[6428] = ~(layer0_outputs[6501]);
    assign outputs[6429] = layer0_outputs[6953];
    assign outputs[6430] = ~(layer0_outputs[3952]);
    assign outputs[6431] = ~((layer0_outputs[6601]) ^ (layer0_outputs[4620]));
    assign outputs[6432] = (layer0_outputs[3965]) & ~(layer0_outputs[1858]);
    assign outputs[6433] = ~((layer0_outputs[3968]) ^ (layer0_outputs[6794]));
    assign outputs[6434] = ~((layer0_outputs[179]) ^ (layer0_outputs[6803]));
    assign outputs[6435] = (layer0_outputs[6260]) ^ (layer0_outputs[6915]);
    assign outputs[6436] = (layer0_outputs[763]) ^ (layer0_outputs[4926]);
    assign outputs[6437] = ~(layer0_outputs[1836]) | (layer0_outputs[916]);
    assign outputs[6438] = ~(layer0_outputs[6614]);
    assign outputs[6439] = layer0_outputs[3520];
    assign outputs[6440] = (layer0_outputs[1550]) & (layer0_outputs[1305]);
    assign outputs[6441] = (layer0_outputs[6070]) ^ (layer0_outputs[5979]);
    assign outputs[6442] = layer0_outputs[1743];
    assign outputs[6443] = ~(layer0_outputs[6015]);
    assign outputs[6444] = (layer0_outputs[7316]) & ~(layer0_outputs[1900]);
    assign outputs[6445] = ~(layer0_outputs[4797]);
    assign outputs[6446] = (layer0_outputs[2763]) & ~(layer0_outputs[72]);
    assign outputs[6447] = layer0_outputs[3709];
    assign outputs[6448] = (layer0_outputs[1597]) ^ (layer0_outputs[2369]);
    assign outputs[6449] = ~(layer0_outputs[5116]) | (layer0_outputs[5451]);
    assign outputs[6450] = (layer0_outputs[1536]) | (layer0_outputs[728]);
    assign outputs[6451] = ~((layer0_outputs[271]) & (layer0_outputs[5432]));
    assign outputs[6452] = ~((layer0_outputs[3402]) & (layer0_outputs[5604]));
    assign outputs[6453] = ~((layer0_outputs[6200]) ^ (layer0_outputs[3936]));
    assign outputs[6454] = ~((layer0_outputs[1087]) ^ (layer0_outputs[5442]));
    assign outputs[6455] = (layer0_outputs[4956]) | (layer0_outputs[6464]);
    assign outputs[6456] = (layer0_outputs[2985]) ^ (layer0_outputs[6406]);
    assign outputs[6457] = ~((layer0_outputs[7287]) ^ (layer0_outputs[1898]));
    assign outputs[6458] = ~((layer0_outputs[3563]) ^ (layer0_outputs[6239]));
    assign outputs[6459] = (layer0_outputs[15]) | (layer0_outputs[5768]);
    assign outputs[6460] = ~(layer0_outputs[633]);
    assign outputs[6461] = ~((layer0_outputs[7166]) ^ (layer0_outputs[4277]));
    assign outputs[6462] = ~(layer0_outputs[7163]) | (layer0_outputs[1899]);
    assign outputs[6463] = ~((layer0_outputs[1213]) | (layer0_outputs[4268]));
    assign outputs[6464] = (layer0_outputs[820]) & (layer0_outputs[3183]);
    assign outputs[6465] = (layer0_outputs[6344]) & (layer0_outputs[6172]);
    assign outputs[6466] = ~(layer0_outputs[2910]);
    assign outputs[6467] = ~(layer0_outputs[3091]) | (layer0_outputs[5588]);
    assign outputs[6468] = (layer0_outputs[2606]) ^ (layer0_outputs[5687]);
    assign outputs[6469] = (layer0_outputs[5005]) & (layer0_outputs[4437]);
    assign outputs[6470] = ~(layer0_outputs[3205]);
    assign outputs[6471] = (layer0_outputs[4614]) & (layer0_outputs[5999]);
    assign outputs[6472] = ~(layer0_outputs[6369]) | (layer0_outputs[7092]);
    assign outputs[6473] = (layer0_outputs[2323]) | (layer0_outputs[4679]);
    assign outputs[6474] = layer0_outputs[4414];
    assign outputs[6475] = ~((layer0_outputs[2416]) ^ (layer0_outputs[2246]));
    assign outputs[6476] = ~((layer0_outputs[5169]) ^ (layer0_outputs[3148]));
    assign outputs[6477] = (layer0_outputs[6443]) ^ (layer0_outputs[2169]);
    assign outputs[6478] = ~(layer0_outputs[2384]) | (layer0_outputs[6137]);
    assign outputs[6479] = layer0_outputs[35];
    assign outputs[6480] = (layer0_outputs[5712]) & ~(layer0_outputs[5401]);
    assign outputs[6481] = (layer0_outputs[1920]) ^ (layer0_outputs[136]);
    assign outputs[6482] = ~(layer0_outputs[3907]);
    assign outputs[6483] = ~((layer0_outputs[2697]) ^ (layer0_outputs[6232]));
    assign outputs[6484] = (layer0_outputs[1668]) | (layer0_outputs[1036]);
    assign outputs[6485] = ~((layer0_outputs[3668]) ^ (layer0_outputs[2691]));
    assign outputs[6486] = ~((layer0_outputs[5947]) & (layer0_outputs[5439]));
    assign outputs[6487] = (layer0_outputs[2328]) ^ (layer0_outputs[5797]);
    assign outputs[6488] = (layer0_outputs[2359]) ^ (layer0_outputs[3458]);
    assign outputs[6489] = ~(layer0_outputs[7636]);
    assign outputs[6490] = (layer0_outputs[940]) & (layer0_outputs[5940]);
    assign outputs[6491] = layer0_outputs[858];
    assign outputs[6492] = ~(layer0_outputs[3001]);
    assign outputs[6493] = ~(layer0_outputs[1189]);
    assign outputs[6494] = (layer0_outputs[3486]) ^ (layer0_outputs[5260]);
    assign outputs[6495] = (layer0_outputs[2823]) & ~(layer0_outputs[7676]);
    assign outputs[6496] = (layer0_outputs[4092]) & (layer0_outputs[7091]);
    assign outputs[6497] = ~((layer0_outputs[1520]) ^ (layer0_outputs[3588]));
    assign outputs[6498] = ~(layer0_outputs[3485]);
    assign outputs[6499] = layer0_outputs[968];
    assign outputs[6500] = ~(layer0_outputs[4621]);
    assign outputs[6501] = ~(layer0_outputs[2338]) | (layer0_outputs[4281]);
    assign outputs[6502] = ~(layer0_outputs[2163]) | (layer0_outputs[7415]);
    assign outputs[6503] = layer0_outputs[4604];
    assign outputs[6504] = ~((layer0_outputs[698]) | (layer0_outputs[895]));
    assign outputs[6505] = layer0_outputs[2982];
    assign outputs[6506] = ~(layer0_outputs[6699]);
    assign outputs[6507] = ~((layer0_outputs[2761]) & (layer0_outputs[6156]));
    assign outputs[6508] = ~(layer0_outputs[889]);
    assign outputs[6509] = (layer0_outputs[5996]) ^ (layer0_outputs[3457]);
    assign outputs[6510] = ~((layer0_outputs[4929]) ^ (layer0_outputs[4670]));
    assign outputs[6511] = (layer0_outputs[7626]) & ~(layer0_outputs[124]);
    assign outputs[6512] = ~((layer0_outputs[7385]) ^ (layer0_outputs[7635]));
    assign outputs[6513] = ~(layer0_outputs[3020]);
    assign outputs[6514] = ~((layer0_outputs[5472]) ^ (layer0_outputs[619]));
    assign outputs[6515] = (layer0_outputs[3196]) | (layer0_outputs[210]);
    assign outputs[6516] = layer0_outputs[1128];
    assign outputs[6517] = ~((layer0_outputs[3289]) & (layer0_outputs[1601]));
    assign outputs[6518] = ~((layer0_outputs[78]) ^ (layer0_outputs[5998]));
    assign outputs[6519] = layer0_outputs[5837];
    assign outputs[6520] = ~(layer0_outputs[2478]);
    assign outputs[6521] = ~(layer0_outputs[5809]) | (layer0_outputs[7281]);
    assign outputs[6522] = ~((layer0_outputs[2003]) ^ (layer0_outputs[2037]));
    assign outputs[6523] = layer0_outputs[3337];
    assign outputs[6524] = (layer0_outputs[5935]) & (layer0_outputs[4925]);
    assign outputs[6525] = layer0_outputs[6557];
    assign outputs[6526] = ~(layer0_outputs[1572]) | (layer0_outputs[4792]);
    assign outputs[6527] = ~(layer0_outputs[600]) | (layer0_outputs[6058]);
    assign outputs[6528] = ~(layer0_outputs[5823]) | (layer0_outputs[711]);
    assign outputs[6529] = (layer0_outputs[1936]) ^ (layer0_outputs[7157]);
    assign outputs[6530] = ~(layer0_outputs[883]);
    assign outputs[6531] = (layer0_outputs[1733]) ^ (layer0_outputs[3656]);
    assign outputs[6532] = ~(layer0_outputs[2297]);
    assign outputs[6533] = ~(layer0_outputs[5313]);
    assign outputs[6534] = (layer0_outputs[5422]) ^ (layer0_outputs[2192]);
    assign outputs[6535] = (layer0_outputs[6517]) & ~(layer0_outputs[4582]);
    assign outputs[6536] = ~(layer0_outputs[5323]);
    assign outputs[6537] = (layer0_outputs[4765]) ^ (layer0_outputs[5628]);
    assign outputs[6538] = ~(layer0_outputs[1903]) | (layer0_outputs[6237]);
    assign outputs[6539] = (layer0_outputs[5786]) ^ (layer0_outputs[6348]);
    assign outputs[6540] = ~(layer0_outputs[4645]);
    assign outputs[6541] = (layer0_outputs[3637]) ^ (layer0_outputs[2465]);
    assign outputs[6542] = ~((layer0_outputs[1546]) | (layer0_outputs[1185]));
    assign outputs[6543] = (layer0_outputs[5946]) | (layer0_outputs[7424]);
    assign outputs[6544] = ~((layer0_outputs[5346]) | (layer0_outputs[1343]));
    assign outputs[6545] = ~((layer0_outputs[6009]) & (layer0_outputs[1781]));
    assign outputs[6546] = layer0_outputs[1668];
    assign outputs[6547] = (layer0_outputs[2098]) ^ (layer0_outputs[1248]);
    assign outputs[6548] = ~((layer0_outputs[897]) & (layer0_outputs[6251]));
    assign outputs[6549] = ~(layer0_outputs[468]);
    assign outputs[6550] = (layer0_outputs[3549]) ^ (layer0_outputs[777]);
    assign outputs[6551] = ~(layer0_outputs[3641]);
    assign outputs[6552] = (layer0_outputs[1646]) | (layer0_outputs[3864]);
    assign outputs[6553] = ~((layer0_outputs[4956]) ^ (layer0_outputs[4077]));
    assign outputs[6554] = (layer0_outputs[6280]) & (layer0_outputs[2753]);
    assign outputs[6555] = ~(layer0_outputs[3914]);
    assign outputs[6556] = ~(layer0_outputs[5665]);
    assign outputs[6557] = (layer0_outputs[1786]) & ~(layer0_outputs[2724]);
    assign outputs[6558] = (layer0_outputs[3744]) ^ (layer0_outputs[3903]);
    assign outputs[6559] = (layer0_outputs[120]) | (layer0_outputs[6020]);
    assign outputs[6560] = ~((layer0_outputs[1345]) ^ (layer0_outputs[3715]));
    assign outputs[6561] = layer0_outputs[1020];
    assign outputs[6562] = ~(layer0_outputs[3127]);
    assign outputs[6563] = (layer0_outputs[3659]) ^ (layer0_outputs[5898]);
    assign outputs[6564] = (layer0_outputs[3646]) | (layer0_outputs[4106]);
    assign outputs[6565] = (layer0_outputs[5344]) & (layer0_outputs[2508]);
    assign outputs[6566] = layer0_outputs[3483];
    assign outputs[6567] = ~(layer0_outputs[5031]);
    assign outputs[6568] = (layer0_outputs[7130]) ^ (layer0_outputs[1197]);
    assign outputs[6569] = ~(layer0_outputs[7500]);
    assign outputs[6570] = ~(layer0_outputs[4416]);
    assign outputs[6571] = ~(layer0_outputs[1100]);
    assign outputs[6572] = (layer0_outputs[7308]) ^ (layer0_outputs[1082]);
    assign outputs[6573] = ~((layer0_outputs[827]) ^ (layer0_outputs[557]));
    assign outputs[6574] = (layer0_outputs[1723]) ^ (layer0_outputs[4097]);
    assign outputs[6575] = (layer0_outputs[2209]) ^ (layer0_outputs[489]);
    assign outputs[6576] = ~(layer0_outputs[3723]) | (layer0_outputs[7167]);
    assign outputs[6577] = (layer0_outputs[4261]) | (layer0_outputs[5420]);
    assign outputs[6578] = ~((layer0_outputs[6008]) ^ (layer0_outputs[6267]));
    assign outputs[6579] = layer0_outputs[1603];
    assign outputs[6580] = 1'b1;
    assign outputs[6581] = ~((layer0_outputs[6763]) ^ (layer0_outputs[5518]));
    assign outputs[6582] = layer0_outputs[991];
    assign outputs[6583] = (layer0_outputs[3378]) & (layer0_outputs[3145]);
    assign outputs[6584] = (layer0_outputs[323]) & (layer0_outputs[4841]);
    assign outputs[6585] = layer0_outputs[896];
    assign outputs[6586] = (layer0_outputs[280]) | (layer0_outputs[2103]);
    assign outputs[6587] = (layer0_outputs[3143]) ^ (layer0_outputs[2582]);
    assign outputs[6588] = layer0_outputs[6296];
    assign outputs[6589] = ~(layer0_outputs[2123]);
    assign outputs[6590] = layer0_outputs[2861];
    assign outputs[6591] = ~(layer0_outputs[2929]);
    assign outputs[6592] = ~((layer0_outputs[4042]) ^ (layer0_outputs[968]));
    assign outputs[6593] = (layer0_outputs[3765]) & (layer0_outputs[353]);
    assign outputs[6594] = layer0_outputs[2365];
    assign outputs[6595] = ~(layer0_outputs[2322]) | (layer0_outputs[302]);
    assign outputs[6596] = ~(layer0_outputs[2804]);
    assign outputs[6597] = ~(layer0_outputs[1908]);
    assign outputs[6598] = ~(layer0_outputs[3336]);
    assign outputs[6599] = (layer0_outputs[1636]) ^ (layer0_outputs[2183]);
    assign outputs[6600] = layer0_outputs[1192];
    assign outputs[6601] = layer0_outputs[4293];
    assign outputs[6602] = layer0_outputs[1639];
    assign outputs[6603] = (layer0_outputs[3984]) ^ (layer0_outputs[3891]);
    assign outputs[6604] = layer0_outputs[5829];
    assign outputs[6605] = ~((layer0_outputs[6482]) ^ (layer0_outputs[4155]));
    assign outputs[6606] = (layer0_outputs[4356]) & (layer0_outputs[1440]);
    assign outputs[6607] = (layer0_outputs[5214]) & (layer0_outputs[422]);
    assign outputs[6608] = ~(layer0_outputs[1320]);
    assign outputs[6609] = ~((layer0_outputs[2090]) | (layer0_outputs[2251]));
    assign outputs[6610] = ~((layer0_outputs[6218]) ^ (layer0_outputs[3855]));
    assign outputs[6611] = ~(layer0_outputs[4007]) | (layer0_outputs[6307]);
    assign outputs[6612] = ~(layer0_outputs[7266]);
    assign outputs[6613] = layer0_outputs[3930];
    assign outputs[6614] = ~(layer0_outputs[4807]);
    assign outputs[6615] = ~((layer0_outputs[6186]) ^ (layer0_outputs[4957]));
    assign outputs[6616] = ~(layer0_outputs[6573]);
    assign outputs[6617] = ~((layer0_outputs[6716]) & (layer0_outputs[3904]));
    assign outputs[6618] = ~(layer0_outputs[6357]) | (layer0_outputs[1929]);
    assign outputs[6619] = ~(layer0_outputs[2245]);
    assign outputs[6620] = layer0_outputs[6998];
    assign outputs[6621] = ~((layer0_outputs[4709]) ^ (layer0_outputs[4152]));
    assign outputs[6622] = layer0_outputs[1814];
    assign outputs[6623] = ~(layer0_outputs[2045]);
    assign outputs[6624] = ~(layer0_outputs[6848]);
    assign outputs[6625] = ~((layer0_outputs[7252]) ^ (layer0_outputs[5275]));
    assign outputs[6626] = ~(layer0_outputs[1111]);
    assign outputs[6627] = (layer0_outputs[781]) ^ (layer0_outputs[601]);
    assign outputs[6628] = ~((layer0_outputs[2042]) | (layer0_outputs[5108]));
    assign outputs[6629] = (layer0_outputs[5578]) ^ (layer0_outputs[7215]);
    assign outputs[6630] = layer0_outputs[1855];
    assign outputs[6631] = ~((layer0_outputs[5635]) | (layer0_outputs[7335]));
    assign outputs[6632] = ~((layer0_outputs[4381]) ^ (layer0_outputs[3184]));
    assign outputs[6633] = (layer0_outputs[4047]) ^ (layer0_outputs[446]);
    assign outputs[6634] = (layer0_outputs[5431]) ^ (layer0_outputs[3643]);
    assign outputs[6635] = ~(layer0_outputs[3826]) | (layer0_outputs[612]);
    assign outputs[6636] = ~((layer0_outputs[2075]) & (layer0_outputs[3072]));
    assign outputs[6637] = (layer0_outputs[6175]) ^ (layer0_outputs[2962]);
    assign outputs[6638] = layer0_outputs[272];
    assign outputs[6639] = (layer0_outputs[3061]) ^ (layer0_outputs[5582]);
    assign outputs[6640] = ~((layer0_outputs[7336]) | (layer0_outputs[6290]));
    assign outputs[6641] = ~(layer0_outputs[769]);
    assign outputs[6642] = layer0_outputs[285];
    assign outputs[6643] = (layer0_outputs[5548]) ^ (layer0_outputs[6111]);
    assign outputs[6644] = ~(layer0_outputs[851]) | (layer0_outputs[2793]);
    assign outputs[6645] = layer0_outputs[6025];
    assign outputs[6646] = (layer0_outputs[6706]) ^ (layer0_outputs[4779]);
    assign outputs[6647] = (layer0_outputs[1486]) ^ (layer0_outputs[6014]);
    assign outputs[6648] = ~((layer0_outputs[4006]) ^ (layer0_outputs[1970]));
    assign outputs[6649] = layer0_outputs[4891];
    assign outputs[6650] = ~(layer0_outputs[1377]) | (layer0_outputs[536]);
    assign outputs[6651] = ~(layer0_outputs[992]);
    assign outputs[6652] = ~((layer0_outputs[7659]) ^ (layer0_outputs[3445]));
    assign outputs[6653] = ~((layer0_outputs[3214]) ^ (layer0_outputs[2920]));
    assign outputs[6654] = (layer0_outputs[6606]) ^ (layer0_outputs[6397]);
    assign outputs[6655] = ~(layer0_outputs[1628]) | (layer0_outputs[4063]);
    assign outputs[6656] = layer0_outputs[2258];
    assign outputs[6657] = (layer0_outputs[3769]) & ~(layer0_outputs[4442]);
    assign outputs[6658] = ~(layer0_outputs[2553]);
    assign outputs[6659] = ~(layer0_outputs[164]);
    assign outputs[6660] = (layer0_outputs[3970]) & ~(layer0_outputs[7133]);
    assign outputs[6661] = layer0_outputs[350];
    assign outputs[6662] = (layer0_outputs[5006]) ^ (layer0_outputs[4826]);
    assign outputs[6663] = (layer0_outputs[6666]) ^ (layer0_outputs[5183]);
    assign outputs[6664] = (layer0_outputs[509]) & ~(layer0_outputs[7648]);
    assign outputs[6665] = ~((layer0_outputs[7366]) ^ (layer0_outputs[7030]));
    assign outputs[6666] = (layer0_outputs[5750]) ^ (layer0_outputs[6405]);
    assign outputs[6667] = (layer0_outputs[6220]) | (layer0_outputs[3671]);
    assign outputs[6668] = layer0_outputs[119];
    assign outputs[6669] = (layer0_outputs[2058]) | (layer0_outputs[5788]);
    assign outputs[6670] = (layer0_outputs[2052]) ^ (layer0_outputs[6724]);
    assign outputs[6671] = (layer0_outputs[2678]) | (layer0_outputs[7114]);
    assign outputs[6672] = ~(layer0_outputs[4086]) | (layer0_outputs[5409]);
    assign outputs[6673] = (layer0_outputs[2735]) ^ (layer0_outputs[5799]);
    assign outputs[6674] = layer0_outputs[6196];
    assign outputs[6675] = ~(layer0_outputs[7487]);
    assign outputs[6676] = (layer0_outputs[114]) ^ (layer0_outputs[2150]);
    assign outputs[6677] = layer0_outputs[6334];
    assign outputs[6678] = (layer0_outputs[4819]) | (layer0_outputs[1058]);
    assign outputs[6679] = ~(layer0_outputs[7601]);
    assign outputs[6680] = 1'b0;
    assign outputs[6681] = ~(layer0_outputs[4313]);
    assign outputs[6682] = ~(layer0_outputs[4576]);
    assign outputs[6683] = ~(layer0_outputs[2513]) | (layer0_outputs[7187]);
    assign outputs[6684] = ~(layer0_outputs[1365]);
    assign outputs[6685] = (layer0_outputs[5184]) ^ (layer0_outputs[6793]);
    assign outputs[6686] = (layer0_outputs[6761]) & (layer0_outputs[2780]);
    assign outputs[6687] = layer0_outputs[7528];
    assign outputs[6688] = ~(layer0_outputs[6256]);
    assign outputs[6689] = ~((layer0_outputs[6753]) ^ (layer0_outputs[2680]));
    assign outputs[6690] = ~(layer0_outputs[4387]) | (layer0_outputs[2901]);
    assign outputs[6691] = (layer0_outputs[669]) | (layer0_outputs[3788]);
    assign outputs[6692] = (layer0_outputs[7525]) & (layer0_outputs[6669]);
    assign outputs[6693] = ~(layer0_outputs[3001]);
    assign outputs[6694] = ~(layer0_outputs[5713]);
    assign outputs[6695] = layer0_outputs[197];
    assign outputs[6696] = (layer0_outputs[2783]) ^ (layer0_outputs[2271]);
    assign outputs[6697] = ~((layer0_outputs[362]) | (layer0_outputs[5404]));
    assign outputs[6698] = (layer0_outputs[859]) ^ (layer0_outputs[3013]);
    assign outputs[6699] = ~((layer0_outputs[4763]) ^ (layer0_outputs[4133]));
    assign outputs[6700] = layer0_outputs[422];
    assign outputs[6701] = ~(layer0_outputs[3315]);
    assign outputs[6702] = ~(layer0_outputs[3989]);
    assign outputs[6703] = layer0_outputs[7548];
    assign outputs[6704] = ~((layer0_outputs[4116]) | (layer0_outputs[2663]));
    assign outputs[6705] = (layer0_outputs[4601]) ^ (layer0_outputs[2056]);
    assign outputs[6706] = ~(layer0_outputs[459]);
    assign outputs[6707] = (layer0_outputs[3285]) & ~(layer0_outputs[3067]);
    assign outputs[6708] = (layer0_outputs[3510]) & (layer0_outputs[7379]);
    assign outputs[6709] = 1'b1;
    assign outputs[6710] = ~((layer0_outputs[2345]) | (layer0_outputs[1871]));
    assign outputs[6711] = (layer0_outputs[3911]) ^ (layer0_outputs[5462]);
    assign outputs[6712] = ~(layer0_outputs[5417]);
    assign outputs[6713] = layer0_outputs[852];
    assign outputs[6714] = (layer0_outputs[2087]) ^ (layer0_outputs[2571]);
    assign outputs[6715] = ~(layer0_outputs[135]) | (layer0_outputs[3743]);
    assign outputs[6716] = layer0_outputs[146];
    assign outputs[6717] = ~(layer0_outputs[1969]) | (layer0_outputs[1040]);
    assign outputs[6718] = layer0_outputs[1889];
    assign outputs[6719] = (layer0_outputs[1382]) & ~(layer0_outputs[63]);
    assign outputs[6720] = 1'b1;
    assign outputs[6721] = layer0_outputs[2948];
    assign outputs[6722] = ~(layer0_outputs[1940]) | (layer0_outputs[3806]);
    assign outputs[6723] = (layer0_outputs[2646]) | (layer0_outputs[1662]);
    assign outputs[6724] = layer0_outputs[6209];
    assign outputs[6725] = ~(layer0_outputs[4842]) | (layer0_outputs[3362]);
    assign outputs[6726] = ~(layer0_outputs[4057]);
    assign outputs[6727] = layer0_outputs[4805];
    assign outputs[6728] = ~(layer0_outputs[6613]);
    assign outputs[6729] = layer0_outputs[3334];
    assign outputs[6730] = ~(layer0_outputs[5595]) | (layer0_outputs[33]);
    assign outputs[6731] = ~(layer0_outputs[7004]);
    assign outputs[6732] = ~(layer0_outputs[6860]) | (layer0_outputs[1079]);
    assign outputs[6733] = ~((layer0_outputs[5620]) ^ (layer0_outputs[6732]));
    assign outputs[6734] = ~((layer0_outputs[251]) & (layer0_outputs[924]));
    assign outputs[6735] = ~(layer0_outputs[5832]) | (layer0_outputs[287]);
    assign outputs[6736] = (layer0_outputs[705]) | (layer0_outputs[4540]);
    assign outputs[6737] = (layer0_outputs[4126]) & (layer0_outputs[7525]);
    assign outputs[6738] = ~(layer0_outputs[1625]);
    assign outputs[6739] = layer0_outputs[2455];
    assign outputs[6740] = ~(layer0_outputs[4531]);
    assign outputs[6741] = ~(layer0_outputs[566]);
    assign outputs[6742] = ~((layer0_outputs[6364]) & (layer0_outputs[4586]));
    assign outputs[6743] = ~((layer0_outputs[7228]) & (layer0_outputs[2894]));
    assign outputs[6744] = layer0_outputs[758];
    assign outputs[6745] = ~(layer0_outputs[3795]);
    assign outputs[6746] = (layer0_outputs[4985]) & ~(layer0_outputs[5460]);
    assign outputs[6747] = (layer0_outputs[2413]) & (layer0_outputs[3603]);
    assign outputs[6748] = ~((layer0_outputs[1193]) ^ (layer0_outputs[7570]));
    assign outputs[6749] = ~((layer0_outputs[3239]) | (layer0_outputs[4590]));
    assign outputs[6750] = layer0_outputs[4035];
    assign outputs[6751] = (layer0_outputs[2433]) & (layer0_outputs[4456]);
    assign outputs[6752] = (layer0_outputs[7495]) ^ (layer0_outputs[2366]);
    assign outputs[6753] = (layer0_outputs[1122]) ^ (layer0_outputs[6066]);
    assign outputs[6754] = ~((layer0_outputs[6937]) ^ (layer0_outputs[1621]));
    assign outputs[6755] = ~((layer0_outputs[5091]) ^ (layer0_outputs[5247]));
    assign outputs[6756] = ~(layer0_outputs[543]);
    assign outputs[6757] = ~(layer0_outputs[3153]);
    assign outputs[6758] = ~((layer0_outputs[8]) ^ (layer0_outputs[4390]));
    assign outputs[6759] = ~(layer0_outputs[150]);
    assign outputs[6760] = ~((layer0_outputs[1949]) ^ (layer0_outputs[1230]));
    assign outputs[6761] = ~((layer0_outputs[986]) & (layer0_outputs[522]));
    assign outputs[6762] = ~((layer0_outputs[4083]) & (layer0_outputs[2281]));
    assign outputs[6763] = ~(layer0_outputs[3998]);
    assign outputs[6764] = ~((layer0_outputs[5254]) & (layer0_outputs[3790]));
    assign outputs[6765] = ~(layer0_outputs[34]);
    assign outputs[6766] = ~(layer0_outputs[3878]) | (layer0_outputs[3783]);
    assign outputs[6767] = ~((layer0_outputs[1947]) ^ (layer0_outputs[6563]));
    assign outputs[6768] = ~(layer0_outputs[2184]);
    assign outputs[6769] = ~((layer0_outputs[1135]) ^ (layer0_outputs[7178]));
    assign outputs[6770] = ~((layer0_outputs[2237]) ^ (layer0_outputs[461]));
    assign outputs[6771] = layer0_outputs[5636];
    assign outputs[6772] = (layer0_outputs[1243]) ^ (layer0_outputs[3528]);
    assign outputs[6773] = layer0_outputs[2883];
    assign outputs[6774] = ~(layer0_outputs[5138]);
    assign outputs[6775] = ~((layer0_outputs[959]) ^ (layer0_outputs[4842]));
    assign outputs[6776] = (layer0_outputs[1836]) ^ (layer0_outputs[6033]);
    assign outputs[6777] = ~(layer0_outputs[7145]);
    assign outputs[6778] = (layer0_outputs[3000]) & (layer0_outputs[5606]);
    assign outputs[6779] = (layer0_outputs[1917]) & ~(layer0_outputs[6356]);
    assign outputs[6780] = (layer0_outputs[1676]) ^ (layer0_outputs[1955]);
    assign outputs[6781] = layer0_outputs[7621];
    assign outputs[6782] = layer0_outputs[6345];
    assign outputs[6783] = ~(layer0_outputs[3574]);
    assign outputs[6784] = ~((layer0_outputs[7468]) ^ (layer0_outputs[4877]));
    assign outputs[6785] = ~((layer0_outputs[5964]) ^ (layer0_outputs[6915]));
    assign outputs[6786] = layer0_outputs[1221];
    assign outputs[6787] = (layer0_outputs[3747]) & ~(layer0_outputs[5661]);
    assign outputs[6788] = ~((layer0_outputs[7416]) ^ (layer0_outputs[5677]));
    assign outputs[6789] = layer0_outputs[7587];
    assign outputs[6790] = ~((layer0_outputs[3210]) ^ (layer0_outputs[5367]));
    assign outputs[6791] = ~((layer0_outputs[3629]) ^ (layer0_outputs[2551]));
    assign outputs[6792] = (layer0_outputs[5710]) ^ (layer0_outputs[5746]);
    assign outputs[6793] = ~((layer0_outputs[2952]) ^ (layer0_outputs[1980]));
    assign outputs[6794] = ~((layer0_outputs[4706]) | (layer0_outputs[6988]));
    assign outputs[6795] = (layer0_outputs[6005]) ^ (layer0_outputs[7599]);
    assign outputs[6796] = ~(layer0_outputs[5203]) | (layer0_outputs[837]);
    assign outputs[6797] = ~(layer0_outputs[346]);
    assign outputs[6798] = layer0_outputs[7161];
    assign outputs[6799] = ~((layer0_outputs[3914]) | (layer0_outputs[1740]));
    assign outputs[6800] = layer0_outputs[3740];
    assign outputs[6801] = ~((layer0_outputs[4918]) | (layer0_outputs[2017]));
    assign outputs[6802] = ~(layer0_outputs[7386]);
    assign outputs[6803] = (layer0_outputs[3581]) ^ (layer0_outputs[5982]);
    assign outputs[6804] = layer0_outputs[1426];
    assign outputs[6805] = layer0_outputs[3942];
    assign outputs[6806] = ~((layer0_outputs[5744]) ^ (layer0_outputs[3746]));
    assign outputs[6807] = ~((layer0_outputs[749]) & (layer0_outputs[7616]));
    assign outputs[6808] = ~((layer0_outputs[1526]) ^ (layer0_outputs[3899]));
    assign outputs[6809] = layer0_outputs[1591];
    assign outputs[6810] = ~((layer0_outputs[6199]) ^ (layer0_outputs[5535]));
    assign outputs[6811] = (layer0_outputs[4946]) ^ (layer0_outputs[294]);
    assign outputs[6812] = (layer0_outputs[5391]) & ~(layer0_outputs[1686]);
    assign outputs[6813] = ~((layer0_outputs[2516]) ^ (layer0_outputs[245]));
    assign outputs[6814] = layer0_outputs[5338];
    assign outputs[6815] = ~(layer0_outputs[2692]);
    assign outputs[6816] = layer0_outputs[4875];
    assign outputs[6817] = layer0_outputs[2794];
    assign outputs[6818] = ~((layer0_outputs[1818]) | (layer0_outputs[2111]));
    assign outputs[6819] = layer0_outputs[4979];
    assign outputs[6820] = (layer0_outputs[3217]) ^ (layer0_outputs[15]);
    assign outputs[6821] = layer0_outputs[294];
    assign outputs[6822] = layer0_outputs[7092];
    assign outputs[6823] = ~((layer0_outputs[4050]) | (layer0_outputs[589]));
    assign outputs[6824] = ~(layer0_outputs[1063]) | (layer0_outputs[3470]);
    assign outputs[6825] = (layer0_outputs[4659]) ^ (layer0_outputs[2808]);
    assign outputs[6826] = layer0_outputs[7273];
    assign outputs[6827] = ~(layer0_outputs[5076]) | (layer0_outputs[1208]);
    assign outputs[6828] = ~(layer0_outputs[4366]) | (layer0_outputs[4980]);
    assign outputs[6829] = layer0_outputs[2239];
    assign outputs[6830] = ~(layer0_outputs[3118]);
    assign outputs[6831] = layer0_outputs[4986];
    assign outputs[6832] = ~(layer0_outputs[6408]);
    assign outputs[6833] = (layer0_outputs[3858]) | (layer0_outputs[7498]);
    assign outputs[6834] = layer0_outputs[6509];
    assign outputs[6835] = ~((layer0_outputs[1003]) ^ (layer0_outputs[6795]));
    assign outputs[6836] = ~((layer0_outputs[4536]) ^ (layer0_outputs[3228]));
    assign outputs[6837] = ~(layer0_outputs[6322]);
    assign outputs[6838] = ~(layer0_outputs[892]);
    assign outputs[6839] = ~(layer0_outputs[7177]);
    assign outputs[6840] = ~((layer0_outputs[4710]) ^ (layer0_outputs[366]));
    assign outputs[6841] = (layer0_outputs[6578]) | (layer0_outputs[1281]);
    assign outputs[6842] = (layer0_outputs[4415]) | (layer0_outputs[2635]);
    assign outputs[6843] = (layer0_outputs[6702]) | (layer0_outputs[4426]);
    assign outputs[6844] = layer0_outputs[7306];
    assign outputs[6845] = ~((layer0_outputs[2539]) ^ (layer0_outputs[6676]));
    assign outputs[6846] = (layer0_outputs[5479]) ^ (layer0_outputs[3756]);
    assign outputs[6847] = ~((layer0_outputs[2644]) | (layer0_outputs[7670]));
    assign outputs[6848] = ~((layer0_outputs[1194]) | (layer0_outputs[2511]));
    assign outputs[6849] = (layer0_outputs[6287]) & (layer0_outputs[7577]);
    assign outputs[6850] = layer0_outputs[6700];
    assign outputs[6851] = layer0_outputs[1348];
    assign outputs[6852] = (layer0_outputs[1618]) ^ (layer0_outputs[3454]);
    assign outputs[6853] = ~(layer0_outputs[5052]) | (layer0_outputs[3632]);
    assign outputs[6854] = ~((layer0_outputs[4991]) ^ (layer0_outputs[1594]));
    assign outputs[6855] = ~(layer0_outputs[5217]) | (layer0_outputs[2074]);
    assign outputs[6856] = ~(layer0_outputs[326]);
    assign outputs[6857] = (layer0_outputs[5707]) & ~(layer0_outputs[7470]);
    assign outputs[6858] = ~((layer0_outputs[6826]) ^ (layer0_outputs[1675]));
    assign outputs[6859] = ~((layer0_outputs[69]) ^ (layer0_outputs[6995]));
    assign outputs[6860] = (layer0_outputs[5021]) ^ (layer0_outputs[6461]);
    assign outputs[6861] = ~(layer0_outputs[1868]);
    assign outputs[6862] = (layer0_outputs[1498]) | (layer0_outputs[1593]);
    assign outputs[6863] = (layer0_outputs[2362]) ^ (layer0_outputs[3822]);
    assign outputs[6864] = (layer0_outputs[7076]) & ~(layer0_outputs[1432]);
    assign outputs[6865] = layer0_outputs[243];
    assign outputs[6866] = ~((layer0_outputs[1427]) ^ (layer0_outputs[1040]));
    assign outputs[6867] = (layer0_outputs[4566]) ^ (layer0_outputs[3343]);
    assign outputs[6868] = layer0_outputs[2901];
    assign outputs[6869] = (layer0_outputs[4492]) ^ (layer0_outputs[7646]);
    assign outputs[6870] = layer0_outputs[7531];
    assign outputs[6871] = ~((layer0_outputs[3683]) | (layer0_outputs[5641]));
    assign outputs[6872] = ~(layer0_outputs[1756]) | (layer0_outputs[236]);
    assign outputs[6873] = ~(layer0_outputs[3369]);
    assign outputs[6874] = ~((layer0_outputs[7291]) | (layer0_outputs[3324]));
    assign outputs[6875] = layer0_outputs[3071];
    assign outputs[6876] = layer0_outputs[3797];
    assign outputs[6877] = ~(layer0_outputs[5673]) | (layer0_outputs[6057]);
    assign outputs[6878] = ~(layer0_outputs[6704]);
    assign outputs[6879] = (layer0_outputs[2546]) ^ (layer0_outputs[4921]);
    assign outputs[6880] = ~(layer0_outputs[1798]);
    assign outputs[6881] = ~(layer0_outputs[6358]) | (layer0_outputs[3058]);
    assign outputs[6882] = ~(layer0_outputs[2302]);
    assign outputs[6883] = ~(layer0_outputs[4053]);
    assign outputs[6884] = ~(layer0_outputs[1810]) | (layer0_outputs[3787]);
    assign outputs[6885] = layer0_outputs[2631];
    assign outputs[6886] = ~(layer0_outputs[5291]) | (layer0_outputs[7446]);
    assign outputs[6887] = layer0_outputs[4269];
    assign outputs[6888] = ~(layer0_outputs[4104]);
    assign outputs[6889] = (layer0_outputs[1941]) ^ (layer0_outputs[1911]);
    assign outputs[6890] = ~((layer0_outputs[6779]) ^ (layer0_outputs[1190]));
    assign outputs[6891] = ~((layer0_outputs[7480]) | (layer0_outputs[6833]));
    assign outputs[6892] = (layer0_outputs[2402]) & (layer0_outputs[4491]);
    assign outputs[6893] = ~(layer0_outputs[4209]);
    assign outputs[6894] = ~((layer0_outputs[6648]) ^ (layer0_outputs[7451]));
    assign outputs[6895] = layer0_outputs[4214];
    assign outputs[6896] = ~((layer0_outputs[3276]) ^ (layer0_outputs[4127]));
    assign outputs[6897] = (layer0_outputs[5913]) ^ (layer0_outputs[2748]);
    assign outputs[6898] = layer0_outputs[4556];
    assign outputs[6899] = ~((layer0_outputs[4514]) & (layer0_outputs[853]));
    assign outputs[6900] = ~(layer0_outputs[3536]);
    assign outputs[6901] = (layer0_outputs[1886]) ^ (layer0_outputs[4735]);
    assign outputs[6902] = layer0_outputs[4450];
    assign outputs[6903] = layer0_outputs[5636];
    assign outputs[6904] = layer0_outputs[1144];
    assign outputs[6905] = (layer0_outputs[4597]) & ~(layer0_outputs[6083]);
    assign outputs[6906] = ~((layer0_outputs[387]) | (layer0_outputs[4932]));
    assign outputs[6907] = (layer0_outputs[3932]) & (layer0_outputs[6569]);
    assign outputs[6908] = layer0_outputs[5158];
    assign outputs[6909] = ~(layer0_outputs[5582]);
    assign outputs[6910] = ~((layer0_outputs[5276]) ^ (layer0_outputs[1879]));
    assign outputs[6911] = layer0_outputs[2535];
    assign outputs[6912] = (layer0_outputs[6913]) & (layer0_outputs[5978]);
    assign outputs[6913] = ~(layer0_outputs[7342]);
    assign outputs[6914] = ~(layer0_outputs[7168]);
    assign outputs[6915] = (layer0_outputs[2739]) ^ (layer0_outputs[4177]);
    assign outputs[6916] = layer0_outputs[1821];
    assign outputs[6917] = (layer0_outputs[5658]) & ~(layer0_outputs[2092]);
    assign outputs[6918] = layer0_outputs[1240];
    assign outputs[6919] = (layer0_outputs[4221]) & ~(layer0_outputs[722]);
    assign outputs[6920] = ~((layer0_outputs[4316]) | (layer0_outputs[6401]));
    assign outputs[6921] = ~((layer0_outputs[378]) ^ (layer0_outputs[6168]));
    assign outputs[6922] = layer0_outputs[2053];
    assign outputs[6923] = ~((layer0_outputs[3312]) & (layer0_outputs[2517]));
    assign outputs[6924] = ~(layer0_outputs[4350]);
    assign outputs[6925] = (layer0_outputs[5881]) & ~(layer0_outputs[5456]);
    assign outputs[6926] = (layer0_outputs[4299]) & ~(layer0_outputs[5538]);
    assign outputs[6927] = (layer0_outputs[138]) ^ (layer0_outputs[1459]);
    assign outputs[6928] = layer0_outputs[5489];
    assign outputs[6929] = ~((layer0_outputs[4153]) ^ (layer0_outputs[7667]));
    assign outputs[6930] = ~(layer0_outputs[2447]);
    assign outputs[6931] = (layer0_outputs[2784]) | (layer0_outputs[6391]);
    assign outputs[6932] = (layer0_outputs[7086]) ^ (layer0_outputs[94]);
    assign outputs[6933] = layer0_outputs[3531];
    assign outputs[6934] = ~((layer0_outputs[4323]) | (layer0_outputs[6465]));
    assign outputs[6935] = (layer0_outputs[2439]) & ~(layer0_outputs[4404]);
    assign outputs[6936] = ~((layer0_outputs[7439]) ^ (layer0_outputs[1211]));
    assign outputs[6937] = ~(layer0_outputs[595]);
    assign outputs[6938] = layer0_outputs[4287];
    assign outputs[6939] = layer0_outputs[4207];
    assign outputs[6940] = ~((layer0_outputs[1265]) ^ (layer0_outputs[2796]));
    assign outputs[6941] = layer0_outputs[4394];
    assign outputs[6942] = ~(layer0_outputs[1302]);
    assign outputs[6943] = (layer0_outputs[4826]) & (layer0_outputs[1754]);
    assign outputs[6944] = (layer0_outputs[4972]) & ~(layer0_outputs[880]);
    assign outputs[6945] = ~(layer0_outputs[257]);
    assign outputs[6946] = (layer0_outputs[4845]) & ~(layer0_outputs[3870]);
    assign outputs[6947] = (layer0_outputs[1273]) & (layer0_outputs[4902]);
    assign outputs[6948] = ~(layer0_outputs[4943]) | (layer0_outputs[2342]);
    assign outputs[6949] = layer0_outputs[7454];
    assign outputs[6950] = ~(layer0_outputs[6673]);
    assign outputs[6951] = ~(layer0_outputs[4425]);
    assign outputs[6952] = ~(layer0_outputs[6535]);
    assign outputs[6953] = ~(layer0_outputs[877]);
    assign outputs[6954] = ~((layer0_outputs[7216]) | (layer0_outputs[1989]));
    assign outputs[6955] = (layer0_outputs[6831]) & ~(layer0_outputs[4233]);
    assign outputs[6956] = (layer0_outputs[6370]) & (layer0_outputs[5029]);
    assign outputs[6957] = ~((layer0_outputs[205]) ^ (layer0_outputs[2134]));
    assign outputs[6958] = layer0_outputs[5686];
    assign outputs[6959] = (layer0_outputs[913]) ^ (layer0_outputs[2054]);
    assign outputs[6960] = (layer0_outputs[5101]) & ~(layer0_outputs[224]);
    assign outputs[6961] = ~(layer0_outputs[7119]);
    assign outputs[6962] = layer0_outputs[5095];
    assign outputs[6963] = ~((layer0_outputs[6242]) ^ (layer0_outputs[6289]));
    assign outputs[6964] = ~(layer0_outputs[6179]);
    assign outputs[6965] = ~(layer0_outputs[7261]) | (layer0_outputs[5123]);
    assign outputs[6966] = ~(layer0_outputs[6119]);
    assign outputs[6967] = (layer0_outputs[1939]) & ~(layer0_outputs[2655]);
    assign outputs[6968] = (layer0_outputs[4505]) ^ (layer0_outputs[2437]);
    assign outputs[6969] = (layer0_outputs[5778]) & (layer0_outputs[4395]);
    assign outputs[6970] = (layer0_outputs[6911]) & ~(layer0_outputs[7448]);
    assign outputs[6971] = ~(layer0_outputs[7376]);
    assign outputs[6972] = layer0_outputs[4581];
    assign outputs[6973] = (layer0_outputs[5957]) & (layer0_outputs[969]);
    assign outputs[6974] = ~((layer0_outputs[7088]) ^ (layer0_outputs[4596]));
    assign outputs[6975] = ~(layer0_outputs[2971]);
    assign outputs[6976] = (layer0_outputs[4410]) ^ (layer0_outputs[1958]);
    assign outputs[6977] = ~(layer0_outputs[5064]);
    assign outputs[6978] = layer0_outputs[2320];
    assign outputs[6979] = ~((layer0_outputs[5236]) | (layer0_outputs[3754]));
    assign outputs[6980] = ~(layer0_outputs[5457]);
    assign outputs[6981] = ~((layer0_outputs[2764]) ^ (layer0_outputs[5228]));
    assign outputs[6982] = (layer0_outputs[7429]) ^ (layer0_outputs[2077]);
    assign outputs[6983] = (layer0_outputs[944]) & (layer0_outputs[7046]);
    assign outputs[6984] = (layer0_outputs[6819]) & (layer0_outputs[3268]);
    assign outputs[6985] = layer0_outputs[3394];
    assign outputs[6986] = ~((layer0_outputs[1454]) ^ (layer0_outputs[4236]));
    assign outputs[6987] = (layer0_outputs[5481]) & ~(layer0_outputs[5826]);
    assign outputs[6988] = (layer0_outputs[6049]) ^ (layer0_outputs[5832]);
    assign outputs[6989] = (layer0_outputs[7244]) & (layer0_outputs[3975]);
    assign outputs[6990] = (layer0_outputs[5115]) & ~(layer0_outputs[6646]);
    assign outputs[6991] = ~((layer0_outputs[2709]) ^ (layer0_outputs[3261]));
    assign outputs[6992] = (layer0_outputs[2597]) & ~(layer0_outputs[4517]);
    assign outputs[6993] = ~((layer0_outputs[6457]) | (layer0_outputs[5003]));
    assign outputs[6994] = ~((layer0_outputs[3665]) | (layer0_outputs[5951]));
    assign outputs[6995] = (layer0_outputs[1474]) | (layer0_outputs[4354]);
    assign outputs[6996] = (layer0_outputs[4589]) ^ (layer0_outputs[2146]);
    assign outputs[6997] = (layer0_outputs[1274]) ^ (layer0_outputs[5934]);
    assign outputs[6998] = ~((layer0_outputs[3884]) ^ (layer0_outputs[7186]));
    assign outputs[6999] = ~((layer0_outputs[4582]) | (layer0_outputs[4454]));
    assign outputs[7000] = ~(layer0_outputs[499]);
    assign outputs[7001] = (layer0_outputs[2852]) & ~(layer0_outputs[4027]);
    assign outputs[7002] = ~(layer0_outputs[6179]);
    assign outputs[7003] = layer0_outputs[1009];
    assign outputs[7004] = ~((layer0_outputs[1961]) | (layer0_outputs[1806]));
    assign outputs[7005] = (layer0_outputs[2299]) & ~(layer0_outputs[912]);
    assign outputs[7006] = ~((layer0_outputs[6994]) & (layer0_outputs[6859]));
    assign outputs[7007] = (layer0_outputs[766]) & ~(layer0_outputs[2621]);
    assign outputs[7008] = (layer0_outputs[6065]) & (layer0_outputs[1156]);
    assign outputs[7009] = ~((layer0_outputs[5018]) | (layer0_outputs[1419]));
    assign outputs[7010] = (layer0_outputs[3859]) & (layer0_outputs[7629]);
    assign outputs[7011] = ~(layer0_outputs[2509]);
    assign outputs[7012] = ~((layer0_outputs[479]) ^ (layer0_outputs[5327]));
    assign outputs[7013] = (layer0_outputs[1920]) ^ (layer0_outputs[6964]);
    assign outputs[7014] = ~((layer0_outputs[4015]) ^ (layer0_outputs[4465]));
    assign outputs[7015] = layer0_outputs[4096];
    assign outputs[7016] = ~(layer0_outputs[4603]);
    assign outputs[7017] = (layer0_outputs[6099]) & ~(layer0_outputs[5351]);
    assign outputs[7018] = ~(layer0_outputs[5093]);
    assign outputs[7019] = (layer0_outputs[1747]) | (layer0_outputs[4773]);
    assign outputs[7020] = (layer0_outputs[4562]) & (layer0_outputs[5303]);
    assign outputs[7021] = layer0_outputs[6742];
    assign outputs[7022] = (layer0_outputs[1633]) ^ (layer0_outputs[1268]);
    assign outputs[7023] = layer0_outputs[713];
    assign outputs[7024] = (layer0_outputs[5285]) ^ (layer0_outputs[5105]);
    assign outputs[7025] = ~(layer0_outputs[6698]);
    assign outputs[7026] = (layer0_outputs[5746]) ^ (layer0_outputs[4379]);
    assign outputs[7027] = ~(layer0_outputs[3700]);
    assign outputs[7028] = (layer0_outputs[5125]) & ~(layer0_outputs[1413]);
    assign outputs[7029] = ~((layer0_outputs[4032]) ^ (layer0_outputs[1707]));
    assign outputs[7030] = ~((layer0_outputs[6366]) & (layer0_outputs[4058]));
    assign outputs[7031] = layer0_outputs[6933];
    assign outputs[7032] = ~((layer0_outputs[4951]) ^ (layer0_outputs[6210]));
    assign outputs[7033] = layer0_outputs[2167];
    assign outputs[7034] = ~((layer0_outputs[2675]) ^ (layer0_outputs[5064]));
    assign outputs[7035] = ~(layer0_outputs[4439]);
    assign outputs[7036] = ~(layer0_outputs[7233]);
    assign outputs[7037] = ~(layer0_outputs[6782]);
    assign outputs[7038] = ~((layer0_outputs[5852]) ^ (layer0_outputs[796]));
    assign outputs[7039] = (layer0_outputs[6304]) ^ (layer0_outputs[4877]);
    assign outputs[7040] = ~((layer0_outputs[7111]) ^ (layer0_outputs[6767]));
    assign outputs[7041] = ~(layer0_outputs[634]);
    assign outputs[7042] = ~(layer0_outputs[5325]) | (layer0_outputs[5335]);
    assign outputs[7043] = layer0_outputs[306];
    assign outputs[7044] = layer0_outputs[5216];
    assign outputs[7045] = ~((layer0_outputs[7228]) | (layer0_outputs[4924]));
    assign outputs[7046] = layer0_outputs[3016];
    assign outputs[7047] = (layer0_outputs[6810]) ^ (layer0_outputs[6810]);
    assign outputs[7048] = ~((layer0_outputs[7650]) ^ (layer0_outputs[4855]));
    assign outputs[7049] = layer0_outputs[5774];
    assign outputs[7050] = (layer0_outputs[1530]) & (layer0_outputs[6793]);
    assign outputs[7051] = (layer0_outputs[5526]) & (layer0_outputs[4318]);
    assign outputs[7052] = (layer0_outputs[5740]) ^ (layer0_outputs[2904]);
    assign outputs[7053] = (layer0_outputs[1972]) ^ (layer0_outputs[4422]);
    assign outputs[7054] = ~((layer0_outputs[3111]) | (layer0_outputs[3302]));
    assign outputs[7055] = layer0_outputs[528];
    assign outputs[7056] = ~((layer0_outputs[662]) ^ (layer0_outputs[2842]));
    assign outputs[7057] = (layer0_outputs[39]) & ~(layer0_outputs[4978]);
    assign outputs[7058] = (layer0_outputs[504]) ^ (layer0_outputs[4481]);
    assign outputs[7059] = ~((layer0_outputs[207]) ^ (layer0_outputs[5599]));
    assign outputs[7060] = layer0_outputs[5172];
    assign outputs[7061] = layer0_outputs[2982];
    assign outputs[7062] = (layer0_outputs[6859]) ^ (layer0_outputs[4935]);
    assign outputs[7063] = layer0_outputs[4595];
    assign outputs[7064] = ~(layer0_outputs[5844]) | (layer0_outputs[2346]);
    assign outputs[7065] = ~(layer0_outputs[376]);
    assign outputs[7066] = ~(layer0_outputs[599]);
    assign outputs[7067] = ~(layer0_outputs[184]);
    assign outputs[7068] = (layer0_outputs[1451]) & ~(layer0_outputs[2821]);
    assign outputs[7069] = (layer0_outputs[2527]) & (layer0_outputs[3852]);
    assign outputs[7070] = (layer0_outputs[7360]) & ~(layer0_outputs[1737]);
    assign outputs[7071] = (layer0_outputs[1908]) & ~(layer0_outputs[248]);
    assign outputs[7072] = (layer0_outputs[1485]) ^ (layer0_outputs[6773]);
    assign outputs[7073] = (layer0_outputs[791]) ^ (layer0_outputs[7021]);
    assign outputs[7074] = layer0_outputs[4448];
    assign outputs[7075] = layer0_outputs[410];
    assign outputs[7076] = layer0_outputs[736];
    assign outputs[7077] = ~(layer0_outputs[4613]);
    assign outputs[7078] = ~(layer0_outputs[6103]);
    assign outputs[7079] = 1'b0;
    assign outputs[7080] = ~(layer0_outputs[7483]);
    assign outputs[7081] = ~(layer0_outputs[4560]);
    assign outputs[7082] = ~(layer0_outputs[3003]);
    assign outputs[7083] = ~((layer0_outputs[774]) ^ (layer0_outputs[3240]));
    assign outputs[7084] = ~(layer0_outputs[6701]);
    assign outputs[7085] = layer0_outputs[1570];
    assign outputs[7086] = ~((layer0_outputs[228]) ^ (layer0_outputs[113]));
    assign outputs[7087] = (layer0_outputs[4227]) ^ (layer0_outputs[6658]);
    assign outputs[7088] = ~((layer0_outputs[2221]) | (layer0_outputs[6068]));
    assign outputs[7089] = (layer0_outputs[5739]) & ~(layer0_outputs[229]);
    assign outputs[7090] = ~(layer0_outputs[378]);
    assign outputs[7091] = layer0_outputs[1479];
    assign outputs[7092] = ~((layer0_outputs[6063]) | (layer0_outputs[2247]));
    assign outputs[7093] = ~(layer0_outputs[4698]) | (layer0_outputs[1380]);
    assign outputs[7094] = layer0_outputs[6309];
    assign outputs[7095] = ~((layer0_outputs[2001]) ^ (layer0_outputs[624]));
    assign outputs[7096] = ~(layer0_outputs[5202]);
    assign outputs[7097] = 1'b0;
    assign outputs[7098] = (layer0_outputs[770]) ^ (layer0_outputs[4350]);
    assign outputs[7099] = layer0_outputs[6620];
    assign outputs[7100] = layer0_outputs[7522];
    assign outputs[7101] = (layer0_outputs[3867]) ^ (layer0_outputs[4434]);
    assign outputs[7102] = layer0_outputs[809];
    assign outputs[7103] = 1'b0;
    assign outputs[7104] = ~(layer0_outputs[1061]);
    assign outputs[7105] = ~((layer0_outputs[1443]) | (layer0_outputs[7156]));
    assign outputs[7106] = layer0_outputs[1069];
    assign outputs[7107] = layer0_outputs[1349];
    assign outputs[7108] = ~(layer0_outputs[4243]);
    assign outputs[7109] = (layer0_outputs[453]) ^ (layer0_outputs[6684]);
    assign outputs[7110] = (layer0_outputs[5992]) ^ (layer0_outputs[3763]);
    assign outputs[7111] = (layer0_outputs[6231]) ^ (layer0_outputs[6612]);
    assign outputs[7112] = ~(layer0_outputs[4100]);
    assign outputs[7113] = ~(layer0_outputs[1851]);
    assign outputs[7114] = (layer0_outputs[6740]) & (layer0_outputs[2922]);
    assign outputs[7115] = layer0_outputs[3687];
    assign outputs[7116] = layer0_outputs[3441];
    assign outputs[7117] = (layer0_outputs[3681]) & ~(layer0_outputs[7082]);
    assign outputs[7118] = ~((layer0_outputs[2264]) | (layer0_outputs[380]));
    assign outputs[7119] = (layer0_outputs[544]) ^ (layer0_outputs[2484]);
    assign outputs[7120] = layer0_outputs[7547];
    assign outputs[7121] = layer0_outputs[4554];
    assign outputs[7122] = ~((layer0_outputs[5964]) | (layer0_outputs[1396]));
    assign outputs[7123] = (layer0_outputs[3729]) ^ (layer0_outputs[1048]);
    assign outputs[7124] = ~(layer0_outputs[6082]);
    assign outputs[7125] = (layer0_outputs[3576]) & (layer0_outputs[3792]);
    assign outputs[7126] = (layer0_outputs[6990]) & ~(layer0_outputs[3440]);
    assign outputs[7127] = layer0_outputs[2109];
    assign outputs[7128] = ~(layer0_outputs[5207]);
    assign outputs[7129] = layer0_outputs[1270];
    assign outputs[7130] = (layer0_outputs[2859]) ^ (layer0_outputs[7554]);
    assign outputs[7131] = ~((layer0_outputs[258]) ^ (layer0_outputs[7149]));
    assign outputs[7132] = ~((layer0_outputs[4274]) ^ (layer0_outputs[3271]));
    assign outputs[7133] = layer0_outputs[3489];
    assign outputs[7134] = layer0_outputs[5698];
    assign outputs[7135] = ~((layer0_outputs[6168]) | (layer0_outputs[1443]));
    assign outputs[7136] = ~(layer0_outputs[3358]);
    assign outputs[7137] = (layer0_outputs[7256]) | (layer0_outputs[3212]);
    assign outputs[7138] = ~(layer0_outputs[7444]);
    assign outputs[7139] = layer0_outputs[2382];
    assign outputs[7140] = layer0_outputs[1446];
    assign outputs[7141] = ~((layer0_outputs[2227]) & (layer0_outputs[735]));
    assign outputs[7142] = ~(layer0_outputs[1372]);
    assign outputs[7143] = ~(layer0_outputs[3697]);
    assign outputs[7144] = layer0_outputs[7639];
    assign outputs[7145] = ~((layer0_outputs[3350]) | (layer0_outputs[1415]));
    assign outputs[7146] = (layer0_outputs[1805]) & (layer0_outputs[3286]);
    assign outputs[7147] = ~(layer0_outputs[2035]);
    assign outputs[7148] = layer0_outputs[6928];
    assign outputs[7149] = (layer0_outputs[1724]) ^ (layer0_outputs[6301]);
    assign outputs[7150] = layer0_outputs[6252];
    assign outputs[7151] = (layer0_outputs[5850]) ^ (layer0_outputs[2536]);
    assign outputs[7152] = layer0_outputs[7412];
    assign outputs[7153] = layer0_outputs[4473];
    assign outputs[7154] = (layer0_outputs[435]) | (layer0_outputs[5868]);
    assign outputs[7155] = (layer0_outputs[7236]) & ~(layer0_outputs[4731]);
    assign outputs[7156] = layer0_outputs[2865];
    assign outputs[7157] = layer0_outputs[5267];
    assign outputs[7158] = layer0_outputs[5218];
    assign outputs[7159] = ~(layer0_outputs[5399]);
    assign outputs[7160] = ~((layer0_outputs[4882]) ^ (layer0_outputs[4037]));
    assign outputs[7161] = (layer0_outputs[2843]) ^ (layer0_outputs[4585]);
    assign outputs[7162] = ~(layer0_outputs[65]);
    assign outputs[7163] = layer0_outputs[847];
    assign outputs[7164] = ~(layer0_outputs[372]);
    assign outputs[7165] = ~(layer0_outputs[701]);
    assign outputs[7166] = ~((layer0_outputs[1125]) | (layer0_outputs[6991]));
    assign outputs[7167] = (layer0_outputs[4809]) & ~(layer0_outputs[2570]);
    assign outputs[7168] = (layer0_outputs[787]) & (layer0_outputs[5622]);
    assign outputs[7169] = (layer0_outputs[3309]) & ~(layer0_outputs[359]);
    assign outputs[7170] = layer0_outputs[4334];
    assign outputs[7171] = (layer0_outputs[2066]) & ~(layer0_outputs[1551]);
    assign outputs[7172] = ~((layer0_outputs[4240]) & (layer0_outputs[4423]));
    assign outputs[7173] = ~(layer0_outputs[4880]);
    assign outputs[7174] = ~(layer0_outputs[4127]);
    assign outputs[7175] = ~((layer0_outputs[6531]) ^ (layer0_outputs[1517]));
    assign outputs[7176] = (layer0_outputs[2717]) & ~(layer0_outputs[6815]);
    assign outputs[7177] = (layer0_outputs[4275]) & (layer0_outputs[3820]);
    assign outputs[7178] = ~((layer0_outputs[1857]) ^ (layer0_outputs[6680]));
    assign outputs[7179] = layer0_outputs[4302];
    assign outputs[7180] = (layer0_outputs[598]) & ~(layer0_outputs[5535]);
    assign outputs[7181] = (layer0_outputs[4522]) & ~(layer0_outputs[343]);
    assign outputs[7182] = (layer0_outputs[1993]) ^ (layer0_outputs[7630]);
    assign outputs[7183] = ~(layer0_outputs[5149]);
    assign outputs[7184] = (layer0_outputs[2000]) & ~(layer0_outputs[2561]);
    assign outputs[7185] = ~((layer0_outputs[2111]) ^ (layer0_outputs[2862]));
    assign outputs[7186] = ~(layer0_outputs[2769]);
    assign outputs[7187] = (layer0_outputs[5705]) ^ (layer0_outputs[2603]);
    assign outputs[7188] = layer0_outputs[286];
    assign outputs[7189] = ~(layer0_outputs[5988]);
    assign outputs[7190] = layer0_outputs[596];
    assign outputs[7191] = (layer0_outputs[7021]) & ~(layer0_outputs[3596]);
    assign outputs[7192] = ~(layer0_outputs[4530]);
    assign outputs[7193] = (layer0_outputs[586]) | (layer0_outputs[1391]);
    assign outputs[7194] = layer0_outputs[5101];
    assign outputs[7195] = (layer0_outputs[3667]) & ~(layer0_outputs[19]);
    assign outputs[7196] = ~(layer0_outputs[4284]);
    assign outputs[7197] = layer0_outputs[6161];
    assign outputs[7198] = layer0_outputs[2710];
    assign outputs[7199] = ~(layer0_outputs[5569]);
    assign outputs[7200] = layer0_outputs[6067];
    assign outputs[7201] = (layer0_outputs[4189]) ^ (layer0_outputs[4130]);
    assign outputs[7202] = layer0_outputs[685];
    assign outputs[7203] = ~(layer0_outputs[1449]) | (layer0_outputs[169]);
    assign outputs[7204] = ~((layer0_outputs[6764]) & (layer0_outputs[4957]));
    assign outputs[7205] = layer0_outputs[7140];
    assign outputs[7206] = layer0_outputs[4185];
    assign outputs[7207] = ~((layer0_outputs[917]) ^ (layer0_outputs[3605]));
    assign outputs[7208] = (layer0_outputs[5182]) ^ (layer0_outputs[5287]);
    assign outputs[7209] = (layer0_outputs[4006]) & (layer0_outputs[2128]);
    assign outputs[7210] = ~(layer0_outputs[5839]);
    assign outputs[7211] = ~((layer0_outputs[696]) | (layer0_outputs[4587]));
    assign outputs[7212] = ~((layer0_outputs[4470]) | (layer0_outputs[1823]));
    assign outputs[7213] = ~((layer0_outputs[2738]) | (layer0_outputs[1641]));
    assign outputs[7214] = ~(layer0_outputs[3293]) | (layer0_outputs[1696]);
    assign outputs[7215] = ~((layer0_outputs[6808]) ^ (layer0_outputs[3412]));
    assign outputs[7216] = 1'b0;
    assign outputs[7217] = ~(layer0_outputs[6766]);
    assign outputs[7218] = (layer0_outputs[7260]) & ~(layer0_outputs[5297]);
    assign outputs[7219] = (layer0_outputs[5727]) ^ (layer0_outputs[3706]);
    assign outputs[7220] = layer0_outputs[3923];
    assign outputs[7221] = layer0_outputs[6139];
    assign outputs[7222] = ~(layer0_outputs[5643]);
    assign outputs[7223] = layer0_outputs[1569];
    assign outputs[7224] = (layer0_outputs[3227]) & (layer0_outputs[1133]);
    assign outputs[7225] = (layer0_outputs[4879]) & ~(layer0_outputs[5542]);
    assign outputs[7226] = ~(layer0_outputs[4576]) | (layer0_outputs[1491]);
    assign outputs[7227] = (layer0_outputs[3012]) & ~(layer0_outputs[416]);
    assign outputs[7228] = layer0_outputs[739];
    assign outputs[7229] = (layer0_outputs[2674]) ^ (layer0_outputs[4172]);
    assign outputs[7230] = layer0_outputs[6442];
    assign outputs[7231] = ~((layer0_outputs[730]) ^ (layer0_outputs[7517]));
    assign outputs[7232] = (layer0_outputs[6007]) ^ (layer0_outputs[2155]);
    assign outputs[7233] = ~(layer0_outputs[3907]);
    assign outputs[7234] = ~((layer0_outputs[2888]) ^ (layer0_outputs[2327]));
    assign outputs[7235] = ~(layer0_outputs[7007]) | (layer0_outputs[4953]);
    assign outputs[7236] = layer0_outputs[4303];
    assign outputs[7237] = (layer0_outputs[6037]) ^ (layer0_outputs[6473]);
    assign outputs[7238] = ~(layer0_outputs[5696]);
    assign outputs[7239] = layer0_outputs[342];
    assign outputs[7240] = (layer0_outputs[7397]) & (layer0_outputs[1833]);
    assign outputs[7241] = ~(layer0_outputs[2368]);
    assign outputs[7242] = layer0_outputs[2027];
    assign outputs[7243] = layer0_outputs[7614];
    assign outputs[7244] = ~(layer0_outputs[2688]);
    assign outputs[7245] = layer0_outputs[3900];
    assign outputs[7246] = ~(layer0_outputs[5607]);
    assign outputs[7247] = (layer0_outputs[6979]) ^ (layer0_outputs[3363]);
    assign outputs[7248] = (layer0_outputs[7571]) ^ (layer0_outputs[2827]);
    assign outputs[7249] = (layer0_outputs[2416]) | (layer0_outputs[1391]);
    assign outputs[7250] = ~((layer0_outputs[7549]) ^ (layer0_outputs[7239]));
    assign outputs[7251] = (layer0_outputs[64]) & ~(layer0_outputs[2086]);
    assign outputs[7252] = ~(layer0_outputs[7501]);
    assign outputs[7253] = ~((layer0_outputs[2626]) ^ (layer0_outputs[2332]));
    assign outputs[7254] = ~((layer0_outputs[4096]) ^ (layer0_outputs[3152]));
    assign outputs[7255] = ~((layer0_outputs[5947]) & (layer0_outputs[605]));
    assign outputs[7256] = ~(layer0_outputs[6013]);
    assign outputs[7257] = (layer0_outputs[2854]) & ~(layer0_outputs[2336]);
    assign outputs[7258] = ~((layer0_outputs[4870]) ^ (layer0_outputs[4552]));
    assign outputs[7259] = ~(layer0_outputs[2813]);
    assign outputs[7260] = (layer0_outputs[5683]) & (layer0_outputs[5235]);
    assign outputs[7261] = ~(layer0_outputs[6509]);
    assign outputs[7262] = ~(layer0_outputs[4774]);
    assign outputs[7263] = (layer0_outputs[3109]) ^ (layer0_outputs[2397]);
    assign outputs[7264] = (layer0_outputs[4009]) ^ (layer0_outputs[447]);
    assign outputs[7265] = layer0_outputs[3193];
    assign outputs[7266] = ~((layer0_outputs[7393]) ^ (layer0_outputs[5808]));
    assign outputs[7267] = (layer0_outputs[789]) & ~(layer0_outputs[7410]);
    assign outputs[7268] = ~(layer0_outputs[31]);
    assign outputs[7269] = ~((layer0_outputs[7509]) | (layer0_outputs[6869]));
    assign outputs[7270] = (layer0_outputs[4751]) ^ (layer0_outputs[1998]);
    assign outputs[7271] = 1'b0;
    assign outputs[7272] = (layer0_outputs[5775]) & (layer0_outputs[5792]);
    assign outputs[7273] = (layer0_outputs[4967]) & ~(layer0_outputs[5200]);
    assign outputs[7274] = (layer0_outputs[5455]) & ~(layer0_outputs[7131]);
    assign outputs[7275] = ~((layer0_outputs[696]) ^ (layer0_outputs[5659]));
    assign outputs[7276] = layer0_outputs[4144];
    assign outputs[7277] = (layer0_outputs[5115]) & (layer0_outputs[3523]);
    assign outputs[7278] = layer0_outputs[313];
    assign outputs[7279] = (layer0_outputs[1567]) & ~(layer0_outputs[5039]);
    assign outputs[7280] = (layer0_outputs[7120]) | (layer0_outputs[1913]);
    assign outputs[7281] = ~(layer0_outputs[6647]);
    assign outputs[7282] = (layer0_outputs[3233]) & ~(layer0_outputs[3785]);
    assign outputs[7283] = (layer0_outputs[1104]) & ~(layer0_outputs[1600]);
    assign outputs[7284] = (layer0_outputs[1625]) & ~(layer0_outputs[7649]);
    assign outputs[7285] = (layer0_outputs[4120]) & (layer0_outputs[2792]);
    assign outputs[7286] = (layer0_outputs[5180]) | (layer0_outputs[486]);
    assign outputs[7287] = layer0_outputs[1561];
    assign outputs[7288] = (layer0_outputs[4153]) & (layer0_outputs[2343]);
    assign outputs[7289] = (layer0_outputs[2537]) ^ (layer0_outputs[623]);
    assign outputs[7290] = ~(layer0_outputs[802]);
    assign outputs[7291] = ~(layer0_outputs[4674]);
    assign outputs[7292] = (layer0_outputs[7226]) ^ (layer0_outputs[7391]);
    assign outputs[7293] = layer0_outputs[6922];
    assign outputs[7294] = ~((layer0_outputs[907]) & (layer0_outputs[13]));
    assign outputs[7295] = layer0_outputs[6379];
    assign outputs[7296] = (layer0_outputs[252]) ^ (layer0_outputs[4704]);
    assign outputs[7297] = ~(layer0_outputs[5860]);
    assign outputs[7298] = (layer0_outputs[3996]) ^ (layer0_outputs[2705]);
    assign outputs[7299] = (layer0_outputs[2766]) ^ (layer0_outputs[3370]);
    assign outputs[7300] = ~((layer0_outputs[2732]) | (layer0_outputs[1433]));
    assign outputs[7301] = (layer0_outputs[3088]) ^ (layer0_outputs[4362]);
    assign outputs[7302] = (layer0_outputs[1643]) & ~(layer0_outputs[3494]);
    assign outputs[7303] = ~(layer0_outputs[125]);
    assign outputs[7304] = ~((layer0_outputs[6100]) ^ (layer0_outputs[5795]));
    assign outputs[7305] = (layer0_outputs[1427]) & (layer0_outputs[4917]);
    assign outputs[7306] = ~((layer0_outputs[418]) ^ (layer0_outputs[677]));
    assign outputs[7307] = ~((layer0_outputs[2588]) | (layer0_outputs[726]));
    assign outputs[7308] = ~(layer0_outputs[975]);
    assign outputs[7309] = ~((layer0_outputs[7509]) | (layer0_outputs[5466]));
    assign outputs[7310] = ~((layer0_outputs[4531]) | (layer0_outputs[6220]));
    assign outputs[7311] = ~(layer0_outputs[1849]);
    assign outputs[7312] = (layer0_outputs[1533]) ^ (layer0_outputs[6249]);
    assign outputs[7313] = (layer0_outputs[419]) & ~(layer0_outputs[1977]);
    assign outputs[7314] = (layer0_outputs[7591]) ^ (layer0_outputs[3787]);
    assign outputs[7315] = (layer0_outputs[4617]) ^ (layer0_outputs[3020]);
    assign outputs[7316] = layer0_outputs[535];
    assign outputs[7317] = (layer0_outputs[215]) & (layer0_outputs[2355]);
    assign outputs[7318] = (layer0_outputs[6176]) ^ (layer0_outputs[2462]);
    assign outputs[7319] = (layer0_outputs[2849]) & (layer0_outputs[2873]);
    assign outputs[7320] = ~(layer0_outputs[6173]) | (layer0_outputs[3425]);
    assign outputs[7321] = ~((layer0_outputs[5384]) | (layer0_outputs[6105]));
    assign outputs[7322] = layer0_outputs[2130];
    assign outputs[7323] = (layer0_outputs[3852]) & (layer0_outputs[858]);
    assign outputs[7324] = (layer0_outputs[3159]) ^ (layer0_outputs[2958]);
    assign outputs[7325] = layer0_outputs[3909];
    assign outputs[7326] = ~(layer0_outputs[3839]);
    assign outputs[7327] = (layer0_outputs[7250]) & ~(layer0_outputs[2475]);
    assign outputs[7328] = ~(layer0_outputs[6411]);
    assign outputs[7329] = ~(layer0_outputs[3154]);
    assign outputs[7330] = ~(layer0_outputs[507]) | (layer0_outputs[4298]);
    assign outputs[7331] = ~(layer0_outputs[3624]);
    assign outputs[7332] = ~(layer0_outputs[3106]);
    assign outputs[7333] = ~(layer0_outputs[3003]);
    assign outputs[7334] = layer0_outputs[1873];
    assign outputs[7335] = (layer0_outputs[5706]) ^ (layer0_outputs[5002]);
    assign outputs[7336] = layer0_outputs[2837];
    assign outputs[7337] = ~((layer0_outputs[3179]) ^ (layer0_outputs[4579]));
    assign outputs[7338] = ~(layer0_outputs[2746]);
    assign outputs[7339] = ~(layer0_outputs[2855]) | (layer0_outputs[3711]);
    assign outputs[7340] = ~((layer0_outputs[731]) | (layer0_outputs[2240]));
    assign outputs[7341] = layer0_outputs[280];
    assign outputs[7342] = ~((layer0_outputs[5827]) | (layer0_outputs[2640]));
    assign outputs[7343] = ~(layer0_outputs[5222]) | (layer0_outputs[2046]);
    assign outputs[7344] = layer0_outputs[6387];
    assign outputs[7345] = (layer0_outputs[6883]) & ~(layer0_outputs[7438]);
    assign outputs[7346] = (layer0_outputs[7516]) & (layer0_outputs[7475]);
    assign outputs[7347] = layer0_outputs[4381];
    assign outputs[7348] = (layer0_outputs[4514]) & ~(layer0_outputs[6006]);
    assign outputs[7349] = ~((layer0_outputs[485]) ^ (layer0_outputs[6737]));
    assign outputs[7350] = (layer0_outputs[299]) & ~(layer0_outputs[5228]);
    assign outputs[7351] = (layer0_outputs[4602]) & ~(layer0_outputs[3090]);
    assign outputs[7352] = layer0_outputs[4298];
    assign outputs[7353] = (layer0_outputs[961]) & (layer0_outputs[2244]);
    assign outputs[7354] = (layer0_outputs[3118]) & ~(layer0_outputs[7113]);
    assign outputs[7355] = ~(layer0_outputs[2432]) | (layer0_outputs[3339]);
    assign outputs[7356] = ~(layer0_outputs[1672]);
    assign outputs[7357] = layer0_outputs[481];
    assign outputs[7358] = ~(layer0_outputs[3422]);
    assign outputs[7359] = ~((layer0_outputs[2668]) ^ (layer0_outputs[3165]));
    assign outputs[7360] = ~((layer0_outputs[1779]) & (layer0_outputs[3631]));
    assign outputs[7361] = ~((layer0_outputs[1725]) ^ (layer0_outputs[2677]));
    assign outputs[7362] = ~((layer0_outputs[309]) & (layer0_outputs[1849]));
    assign outputs[7363] = layer0_outputs[3186];
    assign outputs[7364] = ~(layer0_outputs[4533]);
    assign outputs[7365] = (layer0_outputs[3996]) & ~(layer0_outputs[1405]);
    assign outputs[7366] = ~((layer0_outputs[697]) ^ (layer0_outputs[5297]));
    assign outputs[7367] = (layer0_outputs[927]) & ~(layer0_outputs[7678]);
    assign outputs[7368] = ~(layer0_outputs[5150]);
    assign outputs[7369] = ~((layer0_outputs[5001]) | (layer0_outputs[3392]));
    assign outputs[7370] = (layer0_outputs[3057]) ^ (layer0_outputs[5066]);
    assign outputs[7371] = (layer0_outputs[1039]) ^ (layer0_outputs[1782]);
    assign outputs[7372] = layer0_outputs[6620];
    assign outputs[7373] = (layer0_outputs[3010]) & ~(layer0_outputs[200]);
    assign outputs[7374] = (layer0_outputs[2730]) & (layer0_outputs[947]);
    assign outputs[7375] = layer0_outputs[7130];
    assign outputs[7376] = (layer0_outputs[1072]) | (layer0_outputs[4399]);
    assign outputs[7377] = layer0_outputs[6152];
    assign outputs[7378] = (layer0_outputs[7544]) & ~(layer0_outputs[5006]);
    assign outputs[7379] = ~(layer0_outputs[4645]);
    assign outputs[7380] = (layer0_outputs[3643]) & ~(layer0_outputs[6543]);
    assign outputs[7381] = (layer0_outputs[6833]) ^ (layer0_outputs[826]);
    assign outputs[7382] = layer0_outputs[3181];
    assign outputs[7383] = ~(layer0_outputs[873]);
    assign outputs[7384] = (layer0_outputs[2602]) & ~(layer0_outputs[7287]);
    assign outputs[7385] = layer0_outputs[3005];
    assign outputs[7386] = (layer0_outputs[1853]) & (layer0_outputs[7562]);
    assign outputs[7387] = ~((layer0_outputs[7641]) ^ (layer0_outputs[7173]));
    assign outputs[7388] = ~(layer0_outputs[2721]);
    assign outputs[7389] = (layer0_outputs[5765]) & (layer0_outputs[2718]);
    assign outputs[7390] = (layer0_outputs[6528]) & ~(layer0_outputs[5274]);
    assign outputs[7391] = ~((layer0_outputs[1253]) & (layer0_outputs[3215]));
    assign outputs[7392] = layer0_outputs[832];
    assign outputs[7393] = ~(layer0_outputs[7110]);
    assign outputs[7394] = layer0_outputs[475];
    assign outputs[7395] = (layer0_outputs[4789]) & ~(layer0_outputs[3445]);
    assign outputs[7396] = ~((layer0_outputs[3158]) | (layer0_outputs[751]));
    assign outputs[7397] = ~((layer0_outputs[1981]) | (layer0_outputs[6882]));
    assign outputs[7398] = (layer0_outputs[2460]) & (layer0_outputs[4455]);
    assign outputs[7399] = (layer0_outputs[2066]) & ~(layer0_outputs[2456]);
    assign outputs[7400] = (layer0_outputs[7596]) ^ (layer0_outputs[1551]);
    assign outputs[7401] = ~((layer0_outputs[6153]) ^ (layer0_outputs[6307]));
    assign outputs[7402] = ~(layer0_outputs[2152]);
    assign outputs[7403] = ~(layer0_outputs[768]);
    assign outputs[7404] = layer0_outputs[7196];
    assign outputs[7405] = layer0_outputs[5017];
    assign outputs[7406] = ~((layer0_outputs[6448]) | (layer0_outputs[26]));
    assign outputs[7407] = ~(layer0_outputs[5432]);
    assign outputs[7408] = ~((layer0_outputs[5359]) | (layer0_outputs[1229]));
    assign outputs[7409] = (layer0_outputs[5804]) & ~(layer0_outputs[5909]);
    assign outputs[7410] = (layer0_outputs[22]) & (layer0_outputs[3807]);
    assign outputs[7411] = layer0_outputs[2008];
    assign outputs[7412] = ~(layer0_outputs[4421]);
    assign outputs[7413] = ~((layer0_outputs[4881]) ^ (layer0_outputs[1812]));
    assign outputs[7414] = ~(layer0_outputs[4513]);
    assign outputs[7415] = layer0_outputs[7457];
    assign outputs[7416] = ~(layer0_outputs[7467]);
    assign outputs[7417] = layer0_outputs[7413];
    assign outputs[7418] = ~(layer0_outputs[1654]);
    assign outputs[7419] = ~(layer0_outputs[7553]);
    assign outputs[7420] = ~((layer0_outputs[2080]) | (layer0_outputs[5488]));
    assign outputs[7421] = layer0_outputs[1426];
    assign outputs[7422] = ~((layer0_outputs[1490]) ^ (layer0_outputs[5475]));
    assign outputs[7423] = ~((layer0_outputs[1847]) ^ (layer0_outputs[1939]));
    assign outputs[7424] = (layer0_outputs[399]) & (layer0_outputs[4267]);
    assign outputs[7425] = (layer0_outputs[3349]) | (layer0_outputs[272]);
    assign outputs[7426] = layer0_outputs[7044];
    assign outputs[7427] = ~((layer0_outputs[5068]) ^ (layer0_outputs[2566]));
    assign outputs[7428] = ~(layer0_outputs[4451]) | (layer0_outputs[939]);
    assign outputs[7429] = (layer0_outputs[4984]) ^ (layer0_outputs[6952]);
    assign outputs[7430] = ~(layer0_outputs[6450]);
    assign outputs[7431] = ~(layer0_outputs[4662]);
    assign outputs[7432] = (layer0_outputs[4183]) & ~(layer0_outputs[6811]);
    assign outputs[7433] = ~(layer0_outputs[6223]);
    assign outputs[7434] = (layer0_outputs[3198]) & ~(layer0_outputs[4525]);
    assign outputs[7435] = (layer0_outputs[847]) & ~(layer0_outputs[5971]);
    assign outputs[7436] = ~(layer0_outputs[577]);
    assign outputs[7437] = (layer0_outputs[2104]) ^ (layer0_outputs[2819]);
    assign outputs[7438] = ~(layer0_outputs[6792]);
    assign outputs[7439] = (layer0_outputs[613]) & (layer0_outputs[5500]);
    assign outputs[7440] = (layer0_outputs[6392]) & (layer0_outputs[5742]);
    assign outputs[7441] = ~(layer0_outputs[7582]);
    assign outputs[7442] = ~(layer0_outputs[3551]);
    assign outputs[7443] = layer0_outputs[955];
    assign outputs[7444] = ~((layer0_outputs[5217]) ^ (layer0_outputs[6909]));
    assign outputs[7445] = ~((layer0_outputs[2604]) ^ (layer0_outputs[1004]));
    assign outputs[7446] = layer0_outputs[5758];
    assign outputs[7447] = (layer0_outputs[3794]) ^ (layer0_outputs[4118]);
    assign outputs[7448] = layer0_outputs[5067];
    assign outputs[7449] = ~(layer0_outputs[1734]);
    assign outputs[7450] = (layer0_outputs[7354]) ^ (layer0_outputs[1582]);
    assign outputs[7451] = layer0_outputs[7457];
    assign outputs[7452] = layer0_outputs[1242];
    assign outputs[7453] = (layer0_outputs[850]) ^ (layer0_outputs[726]);
    assign outputs[7454] = ~(layer0_outputs[943]);
    assign outputs[7455] = layer0_outputs[6444];
    assign outputs[7456] = (layer0_outputs[1461]) & ~(layer0_outputs[5065]);
    assign outputs[7457] = (layer0_outputs[5244]) ^ (layer0_outputs[3295]);
    assign outputs[7458] = ~(layer0_outputs[3273]);
    assign outputs[7459] = ~(layer0_outputs[5069]);
    assign outputs[7460] = ~(layer0_outputs[2362]);
    assign outputs[7461] = ~(layer0_outputs[4534]);
    assign outputs[7462] = ~(layer0_outputs[1182]);
    assign outputs[7463] = layer0_outputs[3570];
    assign outputs[7464] = ~((layer0_outputs[5967]) ^ (layer0_outputs[2486]));
    assign outputs[7465] = layer0_outputs[6725];
    assign outputs[7466] = (layer0_outputs[3936]) ^ (layer0_outputs[2377]);
    assign outputs[7467] = ~((layer0_outputs[5717]) | (layer0_outputs[1772]));
    assign outputs[7468] = ~(layer0_outputs[3238]);
    assign outputs[7469] = (layer0_outputs[6925]) & ~(layer0_outputs[10]);
    assign outputs[7470] = ~((layer0_outputs[4308]) ^ (layer0_outputs[2517]));
    assign outputs[7471] = ~((layer0_outputs[5148]) ^ (layer0_outputs[7318]));
    assign outputs[7472] = ~(layer0_outputs[1096]);
    assign outputs[7473] = ~(layer0_outputs[50]);
    assign outputs[7474] = layer0_outputs[7475];
    assign outputs[7475] = ~((layer0_outputs[2488]) | (layer0_outputs[6661]));
    assign outputs[7476] = ~(layer0_outputs[2009]);
    assign outputs[7477] = ~((layer0_outputs[7580]) ^ (layer0_outputs[3112]));
    assign outputs[7478] = layer0_outputs[6508];
    assign outputs[7479] = ~((layer0_outputs[2532]) ^ (layer0_outputs[2262]));
    assign outputs[7480] = ~((layer0_outputs[6873]) | (layer0_outputs[2319]));
    assign outputs[7481] = ~(layer0_outputs[615]);
    assign outputs[7482] = ~((layer0_outputs[3812]) | (layer0_outputs[937]));
    assign outputs[7483] = (layer0_outputs[2735]) & ~(layer0_outputs[4742]);
    assign outputs[7484] = (layer0_outputs[5610]) & (layer0_outputs[2358]);
    assign outputs[7485] = ~(layer0_outputs[6232]);
    assign outputs[7486] = ~((layer0_outputs[473]) | (layer0_outputs[545]));
    assign outputs[7487] = ~(layer0_outputs[5607]);
    assign outputs[7488] = ~((layer0_outputs[1168]) ^ (layer0_outputs[1626]));
    assign outputs[7489] = ~(layer0_outputs[5443]);
    assign outputs[7490] = layer0_outputs[4666];
    assign outputs[7491] = ~(layer0_outputs[3348]);
    assign outputs[7492] = (layer0_outputs[6589]) & (layer0_outputs[7006]);
    assign outputs[7493] = ~(layer0_outputs[3721]);
    assign outputs[7494] = layer0_outputs[3606];
    assign outputs[7495] = ~(layer0_outputs[587]);
    assign outputs[7496] = ~(layer0_outputs[7398]) | (layer0_outputs[1753]);
    assign outputs[7497] = ~(layer0_outputs[4053]);
    assign outputs[7498] = layer0_outputs[1761];
    assign outputs[7499] = ~(layer0_outputs[731]);
    assign outputs[7500] = ~(layer0_outputs[6474]);
    assign outputs[7501] = ~(layer0_outputs[919]) | (layer0_outputs[4488]);
    assign outputs[7502] = ~((layer0_outputs[2293]) & (layer0_outputs[1866]));
    assign outputs[7503] = ~((layer0_outputs[6943]) | (layer0_outputs[4686]));
    assign outputs[7504] = ~(layer0_outputs[4439]);
    assign outputs[7505] = ~((layer0_outputs[4324]) | (layer0_outputs[746]));
    assign outputs[7506] = layer0_outputs[6890];
    assign outputs[7507] = (layer0_outputs[4638]) ^ (layer0_outputs[5264]);
    assign outputs[7508] = ~(layer0_outputs[5060]) | (layer0_outputs[5841]);
    assign outputs[7509] = ~((layer0_outputs[1886]) & (layer0_outputs[6093]));
    assign outputs[7510] = layer0_outputs[1780];
    assign outputs[7511] = (layer0_outputs[2373]) | (layer0_outputs[2726]);
    assign outputs[7512] = ~(layer0_outputs[804]) | (layer0_outputs[2171]);
    assign outputs[7513] = (layer0_outputs[7368]) & ~(layer0_outputs[3256]);
    assign outputs[7514] = layer0_outputs[482];
    assign outputs[7515] = ~((layer0_outputs[4243]) | (layer0_outputs[3111]));
    assign outputs[7516] = (layer0_outputs[156]) ^ (layer0_outputs[5548]);
    assign outputs[7517] = ~((layer0_outputs[3577]) | (layer0_outputs[5403]));
    assign outputs[7518] = (layer0_outputs[7185]) & ~(layer0_outputs[5788]);
    assign outputs[7519] = (layer0_outputs[4718]) & (layer0_outputs[1326]);
    assign outputs[7520] = (layer0_outputs[5893]) ^ (layer0_outputs[4628]);
    assign outputs[7521] = ~((layer0_outputs[545]) ^ (layer0_outputs[1573]));
    assign outputs[7522] = layer0_outputs[4419];
    assign outputs[7523] = layer0_outputs[313];
    assign outputs[7524] = ~(layer0_outputs[867]);
    assign outputs[7525] = layer0_outputs[1173];
    assign outputs[7526] = (layer0_outputs[641]) & (layer0_outputs[6019]);
    assign outputs[7527] = ~((layer0_outputs[5983]) ^ (layer0_outputs[291]));
    assign outputs[7528] = ~((layer0_outputs[6926]) ^ (layer0_outputs[6930]));
    assign outputs[7529] = (layer0_outputs[637]) ^ (layer0_outputs[842]);
    assign outputs[7530] = layer0_outputs[5923];
    assign outputs[7531] = ~((layer0_outputs[4468]) ^ (layer0_outputs[1761]));
    assign outputs[7532] = (layer0_outputs[2865]) & ~(layer0_outputs[5282]);
    assign outputs[7533] = (layer0_outputs[855]) ^ (layer0_outputs[556]);
    assign outputs[7534] = ~(layer0_outputs[7420]);
    assign outputs[7535] = layer0_outputs[2016];
    assign outputs[7536] = layer0_outputs[2323];
    assign outputs[7537] = (layer0_outputs[5111]) ^ (layer0_outputs[3939]);
    assign outputs[7538] = (layer0_outputs[6944]) ^ (layer0_outputs[4098]);
    assign outputs[7539] = ~(layer0_outputs[3978]);
    assign outputs[7540] = ~((layer0_outputs[4110]) ^ (layer0_outputs[3456]));
    assign outputs[7541] = ~(layer0_outputs[5245]);
    assign outputs[7542] = (layer0_outputs[922]) ^ (layer0_outputs[1325]);
    assign outputs[7543] = ~(layer0_outputs[1742]);
    assign outputs[7544] = ~(layer0_outputs[2304]) | (layer0_outputs[4023]);
    assign outputs[7545] = ~((layer0_outputs[2749]) ^ (layer0_outputs[4667]));
    assign outputs[7546] = ~((layer0_outputs[165]) ^ (layer0_outputs[4753]));
    assign outputs[7547] = ~(layer0_outputs[3115]);
    assign outputs[7548] = (layer0_outputs[3416]) & ~(layer0_outputs[2573]);
    assign outputs[7549] = layer0_outputs[4288];
    assign outputs[7550] = (layer0_outputs[4194]) ^ (layer0_outputs[7364]);
    assign outputs[7551] = (layer0_outputs[3524]) & (layer0_outputs[3621]);
    assign outputs[7552] = (layer0_outputs[1598]) & ~(layer0_outputs[7432]);
    assign outputs[7553] = ~(layer0_outputs[2731]);
    assign outputs[7554] = layer0_outputs[3651];
    assign outputs[7555] = ~((layer0_outputs[6356]) | (layer0_outputs[433]));
    assign outputs[7556] = ~((layer0_outputs[4049]) | (layer0_outputs[2440]));
    assign outputs[7557] = layer0_outputs[2105];
    assign outputs[7558] = ~(layer0_outputs[6697]);
    assign outputs[7559] = (layer0_outputs[5965]) & ~(layer0_outputs[3201]);
    assign outputs[7560] = (layer0_outputs[133]) & ~(layer0_outputs[7436]);
    assign outputs[7561] = (layer0_outputs[404]) & (layer0_outputs[2809]);
    assign outputs[7562] = ~(layer0_outputs[2960]);
    assign outputs[7563] = ~(layer0_outputs[6164]);
    assign outputs[7564] = ~((layer0_outputs[3078]) | (layer0_outputs[1335]));
    assign outputs[7565] = (layer0_outputs[4941]) & ~(layer0_outputs[3211]);
    assign outputs[7566] = (layer0_outputs[3927]) & ~(layer0_outputs[2601]);
    assign outputs[7567] = layer0_outputs[2105];
    assign outputs[7568] = (layer0_outputs[5291]) & ~(layer0_outputs[3352]);
    assign outputs[7569] = (layer0_outputs[6765]) & (layer0_outputs[2067]);
    assign outputs[7570] = layer0_outputs[5552];
    assign outputs[7571] = ~(layer0_outputs[2126]);
    assign outputs[7572] = (layer0_outputs[2220]) & ~(layer0_outputs[4095]);
    assign outputs[7573] = layer0_outputs[6358];
    assign outputs[7574] = ~(layer0_outputs[2064]);
    assign outputs[7575] = ~(layer0_outputs[1396]);
    assign outputs[7576] = (layer0_outputs[5283]) ^ (layer0_outputs[4391]);
    assign outputs[7577] = ~((layer0_outputs[3225]) ^ (layer0_outputs[821]));
    assign outputs[7578] = ~((layer0_outputs[2525]) ^ (layer0_outputs[3959]));
    assign outputs[7579] = (layer0_outputs[5987]) ^ (layer0_outputs[3233]);
    assign outputs[7580] = ~((layer0_outputs[5782]) ^ (layer0_outputs[329]));
    assign outputs[7581] = (layer0_outputs[4773]) & (layer0_outputs[4400]);
    assign outputs[7582] = (layer0_outputs[325]) & ~(layer0_outputs[6428]);
    assign outputs[7583] = ~(layer0_outputs[355]);
    assign outputs[7584] = layer0_outputs[5722];
    assign outputs[7585] = (layer0_outputs[2786]) & ~(layer0_outputs[6166]);
    assign outputs[7586] = ~(layer0_outputs[7179]);
    assign outputs[7587] = (layer0_outputs[3865]) & ~(layer0_outputs[3185]);
    assign outputs[7588] = ~((layer0_outputs[2627]) ^ (layer0_outputs[6368]));
    assign outputs[7589] = ~(layer0_outputs[4989]) | (layer0_outputs[6034]);
    assign outputs[7590] = ~((layer0_outputs[764]) ^ (layer0_outputs[3333]));
    assign outputs[7591] = ~(layer0_outputs[4735]);
    assign outputs[7592] = ~((layer0_outputs[6532]) ^ (layer0_outputs[5897]));
    assign outputs[7593] = (layer0_outputs[1064]) & ~(layer0_outputs[4117]);
    assign outputs[7594] = ~(layer0_outputs[4861]);
    assign outputs[7595] = (layer0_outputs[396]) ^ (layer0_outputs[2650]);
    assign outputs[7596] = ~((layer0_outputs[2371]) ^ (layer0_outputs[840]));
    assign outputs[7597] = (layer0_outputs[2532]) & ~(layer0_outputs[5340]);
    assign outputs[7598] = layer0_outputs[1927];
    assign outputs[7599] = ~((layer0_outputs[6308]) | (layer0_outputs[659]));
    assign outputs[7600] = ~((layer0_outputs[1953]) | (layer0_outputs[5370]));
    assign outputs[7601] = (layer0_outputs[4500]) & (layer0_outputs[7620]);
    assign outputs[7602] = ~(layer0_outputs[5798]);
    assign outputs[7603] = (layer0_outputs[5716]) ^ (layer0_outputs[3677]);
    assign outputs[7604] = (layer0_outputs[7012]) & (layer0_outputs[870]);
    assign outputs[7605] = ~(layer0_outputs[5820]);
    assign outputs[7606] = (layer0_outputs[3873]) ^ (layer0_outputs[4211]);
    assign outputs[7607] = layer0_outputs[5321];
    assign outputs[7608] = (layer0_outputs[7245]) & ~(layer0_outputs[1347]);
    assign outputs[7609] = ~(layer0_outputs[2079]);
    assign outputs[7610] = (layer0_outputs[7247]) & (layer0_outputs[2816]);
    assign outputs[7611] = ~((layer0_outputs[548]) ^ (layer0_outputs[3775]));
    assign outputs[7612] = (layer0_outputs[4090]) ^ (layer0_outputs[273]);
    assign outputs[7613] = layer0_outputs[4016];
    assign outputs[7614] = (layer0_outputs[7331]) ^ (layer0_outputs[22]);
    assign outputs[7615] = ~(layer0_outputs[3999]);
    assign outputs[7616] = (layer0_outputs[4888]) ^ (layer0_outputs[5600]);
    assign outputs[7617] = (layer0_outputs[3257]) & ~(layer0_outputs[5012]);
    assign outputs[7618] = ~((layer0_outputs[4747]) | (layer0_outputs[4357]));
    assign outputs[7619] = ~((layer0_outputs[4050]) ^ (layer0_outputs[5077]));
    assign outputs[7620] = layer0_outputs[5777];
    assign outputs[7621] = layer0_outputs[3433];
    assign outputs[7622] = layer0_outputs[7510];
    assign outputs[7623] = layer0_outputs[6143];
    assign outputs[7624] = (layer0_outputs[3908]) ^ (layer0_outputs[2838]);
    assign outputs[7625] = (layer0_outputs[3315]) ^ (layer0_outputs[3917]);
    assign outputs[7626] = (layer0_outputs[260]) & ~(layer0_outputs[6798]);
    assign outputs[7627] = ~((layer0_outputs[3126]) ^ (layer0_outputs[6703]));
    assign outputs[7628] = (layer0_outputs[7214]) & (layer0_outputs[3865]);
    assign outputs[7629] = ~((layer0_outputs[4088]) ^ (layer0_outputs[861]));
    assign outputs[7630] = ~(layer0_outputs[7389]);
    assign outputs[7631] = ~(layer0_outputs[6566]);
    assign outputs[7632] = (layer0_outputs[389]) & ~(layer0_outputs[2340]);
    assign outputs[7633] = (layer0_outputs[3932]) & ~(layer0_outputs[2640]);
    assign outputs[7634] = ~((layer0_outputs[3069]) ^ (layer0_outputs[3605]));
    assign outputs[7635] = ~((layer0_outputs[2590]) & (layer0_outputs[1844]));
    assign outputs[7636] = ~(layer0_outputs[3725]);
    assign outputs[7637] = (layer0_outputs[3645]) ^ (layer0_outputs[6430]);
    assign outputs[7638] = ~((layer0_outputs[4268]) | (layer0_outputs[6692]));
    assign outputs[7639] = ~(layer0_outputs[3099]);
    assign outputs[7640] = ~(layer0_outputs[5815]) | (layer0_outputs[426]);
    assign outputs[7641] = layer0_outputs[2104];
    assign outputs[7642] = layer0_outputs[4342];
    assign outputs[7643] = ~(layer0_outputs[6759]);
    assign outputs[7644] = (layer0_outputs[6275]) | (layer0_outputs[2486]);
    assign outputs[7645] = (layer0_outputs[3109]) ^ (layer0_outputs[6482]);
    assign outputs[7646] = ~(layer0_outputs[5829]);
    assign outputs[7647] = (layer0_outputs[742]) & ~(layer0_outputs[5085]);
    assign outputs[7648] = (layer0_outputs[193]) ^ (layer0_outputs[3288]);
    assign outputs[7649] = (layer0_outputs[1382]) ^ (layer0_outputs[6644]);
    assign outputs[7650] = ~(layer0_outputs[1999]);
    assign outputs[7651] = layer0_outputs[4868];
    assign outputs[7652] = (layer0_outputs[7249]) & ~(layer0_outputs[7401]);
    assign outputs[7653] = ~((layer0_outputs[2172]) ^ (layer0_outputs[1598]));
    assign outputs[7654] = ~((layer0_outputs[0]) | (layer0_outputs[2814]));
    assign outputs[7655] = ~(layer0_outputs[5873]);
    assign outputs[7656] = (layer0_outputs[2946]) ^ (layer0_outputs[339]);
    assign outputs[7657] = ~((layer0_outputs[7117]) ^ (layer0_outputs[6763]));
    assign outputs[7658] = ~(layer0_outputs[6995]);
    assign outputs[7659] = (layer0_outputs[950]) & ~(layer0_outputs[7320]);
    assign outputs[7660] = ~((layer0_outputs[6683]) ^ (layer0_outputs[483]));
    assign outputs[7661] = layer0_outputs[1692];
    assign outputs[7662] = (layer0_outputs[2622]) ^ (layer0_outputs[561]);
    assign outputs[7663] = (layer0_outputs[7294]) & (layer0_outputs[6586]);
    assign outputs[7664] = ~(layer0_outputs[7037]);
    assign outputs[7665] = layer0_outputs[6091];
    assign outputs[7666] = (layer0_outputs[680]) ^ (layer0_outputs[3476]);
    assign outputs[7667] = (layer0_outputs[6170]) ^ (layer0_outputs[1820]);
    assign outputs[7668] = ~(layer0_outputs[4682]) | (layer0_outputs[178]);
    assign outputs[7669] = layer0_outputs[287];
    assign outputs[7670] = (layer0_outputs[265]) & ~(layer0_outputs[5770]);
    assign outputs[7671] = layer0_outputs[1368];
    assign outputs[7672] = ~(layer0_outputs[5974]);
    assign outputs[7673] = ~((layer0_outputs[4080]) & (layer0_outputs[4079]));
    assign outputs[7674] = layer0_outputs[633];
    assign outputs[7675] = ~((layer0_outputs[3741]) ^ (layer0_outputs[3352]));
    assign outputs[7676] = ~(layer0_outputs[1090]);
    assign outputs[7677] = (layer0_outputs[1452]) & (layer0_outputs[745]);
    assign outputs[7678] = ~((layer0_outputs[966]) | (layer0_outputs[4945]));
    assign outputs[7679] = (layer0_outputs[528]) & ~(layer0_outputs[6654]);
endmodule
