library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs: in std_logic_vector(1023 downto 0);
        outputs: out std_logic_vector(9 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs: std_logic_vector(12799 downto 0);

begin
    layer0_outputs(0) <= b and not a;
    layer0_outputs(1) <= not a;
    layer0_outputs(2) <= a xor b;
    layer0_outputs(3) <= a xor b;
    layer0_outputs(4) <= not (a or b);
    layer0_outputs(5) <= a and not b;
    layer0_outputs(6) <= b;
    layer0_outputs(7) <= not (a xor b);
    layer0_outputs(8) <= a and b;
    layer0_outputs(9) <= not (a or b);
    layer0_outputs(10) <= a xor b;
    layer0_outputs(11) <= not a;
    layer0_outputs(12) <= a xor b;
    layer0_outputs(13) <= b and not a;
    layer0_outputs(14) <= b;
    layer0_outputs(15) <= a;
    layer0_outputs(16) <= not (a or b);
    layer0_outputs(17) <= a xor b;
    layer0_outputs(18) <= b;
    layer0_outputs(19) <= not a or b;
    layer0_outputs(20) <= not (a xor b);
    layer0_outputs(21) <= 1'b0;
    layer0_outputs(22) <= not (a xor b);
    layer0_outputs(23) <= b;
    layer0_outputs(24) <= a;
    layer0_outputs(25) <= a xor b;
    layer0_outputs(26) <= not (a or b);
    layer0_outputs(27) <= not b or a;
    layer0_outputs(28) <= b;
    layer0_outputs(29) <= a xor b;
    layer0_outputs(30) <= a or b;
    layer0_outputs(31) <= not (a or b);
    layer0_outputs(32) <= not (a or b);
    layer0_outputs(33) <= not b or a;
    layer0_outputs(34) <= a and not b;
    layer0_outputs(35) <= not (a or b);
    layer0_outputs(36) <= not (a or b);
    layer0_outputs(37) <= b and not a;
    layer0_outputs(38) <= not b;
    layer0_outputs(39) <= not a;
    layer0_outputs(40) <= not b or a;
    layer0_outputs(41) <= a;
    layer0_outputs(42) <= not (a xor b);
    layer0_outputs(43) <= a and b;
    layer0_outputs(44) <= not b or a;
    layer0_outputs(45) <= a;
    layer0_outputs(46) <= not (a and b);
    layer0_outputs(47) <= a xor b;
    layer0_outputs(48) <= a or b;
    layer0_outputs(49) <= not a;
    layer0_outputs(50) <= not b or a;
    layer0_outputs(51) <= not a;
    layer0_outputs(52) <= 1'b0;
    layer0_outputs(53) <= not b or a;
    layer0_outputs(54) <= not b or a;
    layer0_outputs(55) <= a xor b;
    layer0_outputs(56) <= not (a and b);
    layer0_outputs(57) <= not (a or b);
    layer0_outputs(58) <= b and not a;
    layer0_outputs(59) <= not a or b;
    layer0_outputs(60) <= b;
    layer0_outputs(61) <= not (a xor b);
    layer0_outputs(62) <= a xor b;
    layer0_outputs(63) <= a or b;
    layer0_outputs(64) <= not b or a;
    layer0_outputs(65) <= a;
    layer0_outputs(66) <= a or b;
    layer0_outputs(67) <= a xor b;
    layer0_outputs(68) <= 1'b0;
    layer0_outputs(69) <= not b or a;
    layer0_outputs(70) <= a or b;
    layer0_outputs(71) <= not a or b;
    layer0_outputs(72) <= a xor b;
    layer0_outputs(73) <= not (a or b);
    layer0_outputs(74) <= not (a or b);
    layer0_outputs(75) <= not b;
    layer0_outputs(76) <= not (a xor b);
    layer0_outputs(77) <= a and not b;
    layer0_outputs(78) <= a and not b;
    layer0_outputs(79) <= 1'b1;
    layer0_outputs(80) <= not (a xor b);
    layer0_outputs(81) <= a or b;
    layer0_outputs(82) <= not (a or b);
    layer0_outputs(83) <= not (a or b);
    layer0_outputs(84) <= a xor b;
    layer0_outputs(85) <= a or b;
    layer0_outputs(86) <= not b or a;
    layer0_outputs(87) <= b and not a;
    layer0_outputs(88) <= not a;
    layer0_outputs(89) <= b;
    layer0_outputs(90) <= 1'b0;
    layer0_outputs(91) <= b;
    layer0_outputs(92) <= not a;
    layer0_outputs(93) <= a or b;
    layer0_outputs(94) <= not b;
    layer0_outputs(95) <= a xor b;
    layer0_outputs(96) <= b and not a;
    layer0_outputs(97) <= not (a xor b);
    layer0_outputs(98) <= a;
    layer0_outputs(99) <= a xor b;
    layer0_outputs(100) <= b;
    layer0_outputs(101) <= a or b;
    layer0_outputs(102) <= a;
    layer0_outputs(103) <= not a;
    layer0_outputs(104) <= a;
    layer0_outputs(105) <= not b or a;
    layer0_outputs(106) <= a and b;
    layer0_outputs(107) <= not (a xor b);
    layer0_outputs(108) <= not a or b;
    layer0_outputs(109) <= not a or b;
    layer0_outputs(110) <= not (a xor b);
    layer0_outputs(111) <= not (a xor b);
    layer0_outputs(112) <= b;
    layer0_outputs(113) <= a xor b;
    layer0_outputs(114) <= not b;
    layer0_outputs(115) <= not (a xor b);
    layer0_outputs(116) <= a and b;
    layer0_outputs(117) <= not (a xor b);
    layer0_outputs(118) <= not (a and b);
    layer0_outputs(119) <= a xor b;
    layer0_outputs(120) <= not b;
    layer0_outputs(121) <= a;
    layer0_outputs(122) <= a xor b;
    layer0_outputs(123) <= b and not a;
    layer0_outputs(124) <= a;
    layer0_outputs(125) <= a;
    layer0_outputs(126) <= a;
    layer0_outputs(127) <= a;
    layer0_outputs(128) <= not (a xor b);
    layer0_outputs(129) <= not (a or b);
    layer0_outputs(130) <= a xor b;
    layer0_outputs(131) <= a;
    layer0_outputs(132) <= not (a or b);
    layer0_outputs(133) <= not (a xor b);
    layer0_outputs(134) <= b;
    layer0_outputs(135) <= not (a xor b);
    layer0_outputs(136) <= not (a or b);
    layer0_outputs(137) <= a xor b;
    layer0_outputs(138) <= a or b;
    layer0_outputs(139) <= not b;
    layer0_outputs(140) <= b and not a;
    layer0_outputs(141) <= a xor b;
    layer0_outputs(142) <= not b or a;
    layer0_outputs(143) <= not b;
    layer0_outputs(144) <= not (a xor b);
    layer0_outputs(145) <= not a;
    layer0_outputs(146) <= b;
    layer0_outputs(147) <= not (a xor b);
    layer0_outputs(148) <= a or b;
    layer0_outputs(149) <= not (a xor b);
    layer0_outputs(150) <= a and not b;
    layer0_outputs(151) <= a;
    layer0_outputs(152) <= not b;
    layer0_outputs(153) <= not a or b;
    layer0_outputs(154) <= not (a xor b);
    layer0_outputs(155) <= a;
    layer0_outputs(156) <= not (a xor b);
    layer0_outputs(157) <= not (a or b);
    layer0_outputs(158) <= b and not a;
    layer0_outputs(159) <= a and not b;
    layer0_outputs(160) <= a or b;
    layer0_outputs(161) <= a;
    layer0_outputs(162) <= a;
    layer0_outputs(163) <= 1'b0;
    layer0_outputs(164) <= b and not a;
    layer0_outputs(165) <= not (a or b);
    layer0_outputs(166) <= not b or a;
    layer0_outputs(167) <= not (a xor b);
    layer0_outputs(168) <= a or b;
    layer0_outputs(169) <= a;
    layer0_outputs(170) <= not (a or b);
    layer0_outputs(171) <= b and not a;
    layer0_outputs(172) <= not (a xor b);
    layer0_outputs(173) <= b and not a;
    layer0_outputs(174) <= not (a or b);
    layer0_outputs(175) <= not (a and b);
    layer0_outputs(176) <= a;
    layer0_outputs(177) <= b;
    layer0_outputs(178) <= b and not a;
    layer0_outputs(179) <= a and not b;
    layer0_outputs(180) <= a and not b;
    layer0_outputs(181) <= not (a xor b);
    layer0_outputs(182) <= a or b;
    layer0_outputs(183) <= a or b;
    layer0_outputs(184) <= not a or b;
    layer0_outputs(185) <= b;
    layer0_outputs(186) <= b and not a;
    layer0_outputs(187) <= a and not b;
    layer0_outputs(188) <= not b;
    layer0_outputs(189) <= not b;
    layer0_outputs(190) <= a or b;
    layer0_outputs(191) <= not a or b;
    layer0_outputs(192) <= not (a xor b);
    layer0_outputs(193) <= not a or b;
    layer0_outputs(194) <= a xor b;
    layer0_outputs(195) <= a and not b;
    layer0_outputs(196) <= a or b;
    layer0_outputs(197) <= a or b;
    layer0_outputs(198) <= a or b;
    layer0_outputs(199) <= a or b;
    layer0_outputs(200) <= not (a xor b);
    layer0_outputs(201) <= a and not b;
    layer0_outputs(202) <= b and not a;
    layer0_outputs(203) <= not (a xor b);
    layer0_outputs(204) <= 1'b1;
    layer0_outputs(205) <= not a or b;
    layer0_outputs(206) <= a xor b;
    layer0_outputs(207) <= not (a or b);
    layer0_outputs(208) <= b;
    layer0_outputs(209) <= not (a xor b);
    layer0_outputs(210) <= not (a xor b);
    layer0_outputs(211) <= b;
    layer0_outputs(212) <= a or b;
    layer0_outputs(213) <= a and not b;
    layer0_outputs(214) <= a xor b;
    layer0_outputs(215) <= a xor b;
    layer0_outputs(216) <= a and b;
    layer0_outputs(217) <= not a;
    layer0_outputs(218) <= not a or b;
    layer0_outputs(219) <= a;
    layer0_outputs(220) <= not (a or b);
    layer0_outputs(221) <= not b;
    layer0_outputs(222) <= a or b;
    layer0_outputs(223) <= not (a or b);
    layer0_outputs(224) <= not (a xor b);
    layer0_outputs(225) <= not (a or b);
    layer0_outputs(226) <= not b;
    layer0_outputs(227) <= not (a or b);
    layer0_outputs(228) <= a or b;
    layer0_outputs(229) <= not (a or b);
    layer0_outputs(230) <= not b or a;
    layer0_outputs(231) <= not b;
    layer0_outputs(232) <= a or b;
    layer0_outputs(233) <= a;
    layer0_outputs(234) <= 1'b1;
    layer0_outputs(235) <= a xor b;
    layer0_outputs(236) <= not b;
    layer0_outputs(237) <= not (a or b);
    layer0_outputs(238) <= not a or b;
    layer0_outputs(239) <= not (a or b);
    layer0_outputs(240) <= not (a xor b);
    layer0_outputs(241) <= a;
    layer0_outputs(242) <= a or b;
    layer0_outputs(243) <= b and not a;
    layer0_outputs(244) <= not b or a;
    layer0_outputs(245) <= not (a xor b);
    layer0_outputs(246) <= a and not b;
    layer0_outputs(247) <= not a or b;
    layer0_outputs(248) <= not (a or b);
    layer0_outputs(249) <= not b or a;
    layer0_outputs(250) <= a or b;
    layer0_outputs(251) <= not b or a;
    layer0_outputs(252) <= not (a or b);
    layer0_outputs(253) <= a and not b;
    layer0_outputs(254) <= a or b;
    layer0_outputs(255) <= b;
    layer0_outputs(256) <= not (a xor b);
    layer0_outputs(257) <= b;
    layer0_outputs(258) <= not b or a;
    layer0_outputs(259) <= a or b;
    layer0_outputs(260) <= 1'b0;
    layer0_outputs(261) <= not (a or b);
    layer0_outputs(262) <= not (a or b);
    layer0_outputs(263) <= a;
    layer0_outputs(264) <= not (a xor b);
    layer0_outputs(265) <= 1'b1;
    layer0_outputs(266) <= not a;
    layer0_outputs(267) <= b and not a;
    layer0_outputs(268) <= not (a xor b);
    layer0_outputs(269) <= a or b;
    layer0_outputs(270) <= a;
    layer0_outputs(271) <= a and not b;
    layer0_outputs(272) <= a or b;
    layer0_outputs(273) <= not b;
    layer0_outputs(274) <= not a;
    layer0_outputs(275) <= not (a and b);
    layer0_outputs(276) <= b and not a;
    layer0_outputs(277) <= not b or a;
    layer0_outputs(278) <= b;
    layer0_outputs(279) <= not a;
    layer0_outputs(280) <= b and not a;
    layer0_outputs(281) <= not b;
    layer0_outputs(282) <= not a;
    layer0_outputs(283) <= b;
    layer0_outputs(284) <= 1'b0;
    layer0_outputs(285) <= a xor b;
    layer0_outputs(286) <= not (a or b);
    layer0_outputs(287) <= not (a xor b);
    layer0_outputs(288) <= a xor b;
    layer0_outputs(289) <= a xor b;
    layer0_outputs(290) <= a and not b;
    layer0_outputs(291) <= a and not b;
    layer0_outputs(292) <= a and not b;
    layer0_outputs(293) <= a and not b;
    layer0_outputs(294) <= not b or a;
    layer0_outputs(295) <= not (a xor b);
    layer0_outputs(296) <= a;
    layer0_outputs(297) <= not a;
    layer0_outputs(298) <= a xor b;
    layer0_outputs(299) <= a;
    layer0_outputs(300) <= b;
    layer0_outputs(301) <= a and not b;
    layer0_outputs(302) <= a or b;
    layer0_outputs(303) <= b;
    layer0_outputs(304) <= a or b;
    layer0_outputs(305) <= b and not a;
    layer0_outputs(306) <= not a;
    layer0_outputs(307) <= not a or b;
    layer0_outputs(308) <= a and not b;
    layer0_outputs(309) <= not a or b;
    layer0_outputs(310) <= not (a or b);
    layer0_outputs(311) <= a xor b;
    layer0_outputs(312) <= b;
    layer0_outputs(313) <= not a or b;
    layer0_outputs(314) <= a xor b;
    layer0_outputs(315) <= a or b;
    layer0_outputs(316) <= not b or a;
    layer0_outputs(317) <= not (a xor b);
    layer0_outputs(318) <= not a or b;
    layer0_outputs(319) <= not a or b;
    layer0_outputs(320) <= b and not a;
    layer0_outputs(321) <= a or b;
    layer0_outputs(322) <= a;
    layer0_outputs(323) <= b and not a;
    layer0_outputs(324) <= not b or a;
    layer0_outputs(325) <= a xor b;
    layer0_outputs(326) <= not b;
    layer0_outputs(327) <= a or b;
    layer0_outputs(328) <= a;
    layer0_outputs(329) <= not a or b;
    layer0_outputs(330) <= a or b;
    layer0_outputs(331) <= not (a or b);
    layer0_outputs(332) <= 1'b0;
    layer0_outputs(333) <= not b;
    layer0_outputs(334) <= a and not b;
    layer0_outputs(335) <= not b or a;
    layer0_outputs(336) <= not (a xor b);
    layer0_outputs(337) <= a or b;
    layer0_outputs(338) <= not (a and b);
    layer0_outputs(339) <= 1'b0;
    layer0_outputs(340) <= b and not a;
    layer0_outputs(341) <= not a or b;
    layer0_outputs(342) <= a and not b;
    layer0_outputs(343) <= not b;
    layer0_outputs(344) <= a and b;
    layer0_outputs(345) <= not (a xor b);
    layer0_outputs(346) <= b;
    layer0_outputs(347) <= a or b;
    layer0_outputs(348) <= not (a xor b);
    layer0_outputs(349) <= a xor b;
    layer0_outputs(350) <= b;
    layer0_outputs(351) <= not b or a;
    layer0_outputs(352) <= a;
    layer0_outputs(353) <= b and not a;
    layer0_outputs(354) <= not b;
    layer0_outputs(355) <= a;
    layer0_outputs(356) <= a or b;
    layer0_outputs(357) <= a and not b;
    layer0_outputs(358) <= a xor b;
    layer0_outputs(359) <= a;
    layer0_outputs(360) <= b;
    layer0_outputs(361) <= b and not a;
    layer0_outputs(362) <= not b;
    layer0_outputs(363) <= a;
    layer0_outputs(364) <= not a or b;
    layer0_outputs(365) <= b;
    layer0_outputs(366) <= not (a or b);
    layer0_outputs(367) <= b;
    layer0_outputs(368) <= a or b;
    layer0_outputs(369) <= 1'b1;
    layer0_outputs(370) <= not (a xor b);
    layer0_outputs(371) <= b and not a;
    layer0_outputs(372) <= not (a or b);
    layer0_outputs(373) <= not (a or b);
    layer0_outputs(374) <= not a or b;
    layer0_outputs(375) <= not (a or b);
    layer0_outputs(376) <= not (a or b);
    layer0_outputs(377) <= b and not a;
    layer0_outputs(378) <= not (a xor b);
    layer0_outputs(379) <= a or b;
    layer0_outputs(380) <= not (a xor b);
    layer0_outputs(381) <= not (a or b);
    layer0_outputs(382) <= not (a xor b);
    layer0_outputs(383) <= a or b;
    layer0_outputs(384) <= b;
    layer0_outputs(385) <= a and not b;
    layer0_outputs(386) <= b;
    layer0_outputs(387) <= not (a xor b);
    layer0_outputs(388) <= a or b;
    layer0_outputs(389) <= not (a and b);
    layer0_outputs(390) <= a or b;
    layer0_outputs(391) <= a and b;
    layer0_outputs(392) <= a;
    layer0_outputs(393) <= not a;
    layer0_outputs(394) <= not b or a;
    layer0_outputs(395) <= a xor b;
    layer0_outputs(396) <= not b or a;
    layer0_outputs(397) <= a xor b;
    layer0_outputs(398) <= not a;
    layer0_outputs(399) <= not (a xor b);
    layer0_outputs(400) <= a xor b;
    layer0_outputs(401) <= a xor b;
    layer0_outputs(402) <= a;
    layer0_outputs(403) <= 1'b0;
    layer0_outputs(404) <= a or b;
    layer0_outputs(405) <= a or b;
    layer0_outputs(406) <= not a or b;
    layer0_outputs(407) <= a and not b;
    layer0_outputs(408) <= not a or b;
    layer0_outputs(409) <= a xor b;
    layer0_outputs(410) <= a;
    layer0_outputs(411) <= not (a or b);
    layer0_outputs(412) <= not b;
    layer0_outputs(413) <= not b;
    layer0_outputs(414) <= not (a or b);
    layer0_outputs(415) <= not (a xor b);
    layer0_outputs(416) <= not b or a;
    layer0_outputs(417) <= b;
    layer0_outputs(418) <= a;
    layer0_outputs(419) <= a xor b;
    layer0_outputs(420) <= b;
    layer0_outputs(421) <= not a;
    layer0_outputs(422) <= a or b;
    layer0_outputs(423) <= not (a or b);
    layer0_outputs(424) <= a or b;
    layer0_outputs(425) <= a xor b;
    layer0_outputs(426) <= not a or b;
    layer0_outputs(427) <= a and b;
    layer0_outputs(428) <= not b;
    layer0_outputs(429) <= not b;
    layer0_outputs(430) <= a and not b;
    layer0_outputs(431) <= not a;
    layer0_outputs(432) <= not (a or b);
    layer0_outputs(433) <= b and not a;
    layer0_outputs(434) <= not b;
    layer0_outputs(435) <= a or b;
    layer0_outputs(436) <= a and not b;
    layer0_outputs(437) <= a or b;
    layer0_outputs(438) <= not (a xor b);
    layer0_outputs(439) <= not b;
    layer0_outputs(440) <= a;
    layer0_outputs(441) <= not b;
    layer0_outputs(442) <= not a or b;
    layer0_outputs(443) <= not (a xor b);
    layer0_outputs(444) <= not a;
    layer0_outputs(445) <= a or b;
    layer0_outputs(446) <= a xor b;
    layer0_outputs(447) <= not (a or b);
    layer0_outputs(448) <= a or b;
    layer0_outputs(449) <= not (a xor b);
    layer0_outputs(450) <= not b;
    layer0_outputs(451) <= a;
    layer0_outputs(452) <= 1'b0;
    layer0_outputs(453) <= a or b;
    layer0_outputs(454) <= not a or b;
    layer0_outputs(455) <= not a;
    layer0_outputs(456) <= not (a or b);
    layer0_outputs(457) <= a xor b;
    layer0_outputs(458) <= a and b;
    layer0_outputs(459) <= a xor b;
    layer0_outputs(460) <= a xor b;
    layer0_outputs(461) <= not (a or b);
    layer0_outputs(462) <= not b or a;
    layer0_outputs(463) <= not (a xor b);
    layer0_outputs(464) <= a xor b;
    layer0_outputs(465) <= not (a xor b);
    layer0_outputs(466) <= a or b;
    layer0_outputs(467) <= not (a xor b);
    layer0_outputs(468) <= a xor b;
    layer0_outputs(469) <= not a;
    layer0_outputs(470) <= b;
    layer0_outputs(471) <= a xor b;
    layer0_outputs(472) <= a or b;
    layer0_outputs(473) <= not b;
    layer0_outputs(474) <= not a or b;
    layer0_outputs(475) <= a or b;
    layer0_outputs(476) <= a;
    layer0_outputs(477) <= not (a or b);
    layer0_outputs(478) <= a or b;
    layer0_outputs(479) <= a xor b;
    layer0_outputs(480) <= not a;
    layer0_outputs(481) <= a and b;
    layer0_outputs(482) <= not (a xor b);
    layer0_outputs(483) <= not (a xor b);
    layer0_outputs(484) <= not (a xor b);
    layer0_outputs(485) <= a xor b;
    layer0_outputs(486) <= not b or a;
    layer0_outputs(487) <= a;
    layer0_outputs(488) <= not (a or b);
    layer0_outputs(489) <= not b or a;
    layer0_outputs(490) <= not (a or b);
    layer0_outputs(491) <= b;
    layer0_outputs(492) <= a xor b;
    layer0_outputs(493) <= a and not b;
    layer0_outputs(494) <= a xor b;
    layer0_outputs(495) <= 1'b0;
    layer0_outputs(496) <= a or b;
    layer0_outputs(497) <= not (a or b);
    layer0_outputs(498) <= 1'b1;
    layer0_outputs(499) <= b and not a;
    layer0_outputs(500) <= not (a or b);
    layer0_outputs(501) <= not (a or b);
    layer0_outputs(502) <= a xor b;
    layer0_outputs(503) <= a or b;
    layer0_outputs(504) <= a or b;
    layer0_outputs(505) <= a and b;
    layer0_outputs(506) <= a xor b;
    layer0_outputs(507) <= not (a or b);
    layer0_outputs(508) <= a or b;
    layer0_outputs(509) <= a or b;
    layer0_outputs(510) <= b;
    layer0_outputs(511) <= a xor b;
    layer0_outputs(512) <= not (a or b);
    layer0_outputs(513) <= b;
    layer0_outputs(514) <= a or b;
    layer0_outputs(515) <= a and not b;
    layer0_outputs(516) <= b;
    layer0_outputs(517) <= not (a or b);
    layer0_outputs(518) <= not (a or b);
    layer0_outputs(519) <= a xor b;
    layer0_outputs(520) <= b and not a;
    layer0_outputs(521) <= a or b;
    layer0_outputs(522) <= not (a or b);
    layer0_outputs(523) <= not a or b;
    layer0_outputs(524) <= not b or a;
    layer0_outputs(525) <= a or b;
    layer0_outputs(526) <= not b;
    layer0_outputs(527) <= not (a or b);
    layer0_outputs(528) <= a and not b;
    layer0_outputs(529) <= a or b;
    layer0_outputs(530) <= not (a xor b);
    layer0_outputs(531) <= a xor b;
    layer0_outputs(532) <= not (a xor b);
    layer0_outputs(533) <= b and not a;
    layer0_outputs(534) <= a and b;
    layer0_outputs(535) <= b and not a;
    layer0_outputs(536) <= a and not b;
    layer0_outputs(537) <= a and b;
    layer0_outputs(538) <= a or b;
    layer0_outputs(539) <= a or b;
    layer0_outputs(540) <= a or b;
    layer0_outputs(541) <= a xor b;
    layer0_outputs(542) <= not (a xor b);
    layer0_outputs(543) <= not (a xor b);
    layer0_outputs(544) <= not b;
    layer0_outputs(545) <= not (a or b);
    layer0_outputs(546) <= b;
    layer0_outputs(547) <= a xor b;
    layer0_outputs(548) <= not a or b;
    layer0_outputs(549) <= a or b;
    layer0_outputs(550) <= not (a or b);
    layer0_outputs(551) <= b and not a;
    layer0_outputs(552) <= not b or a;
    layer0_outputs(553) <= not b or a;
    layer0_outputs(554) <= not (a or b);
    layer0_outputs(555) <= not (a xor b);
    layer0_outputs(556) <= a and not b;
    layer0_outputs(557) <= a or b;
    layer0_outputs(558) <= not b or a;
    layer0_outputs(559) <= not (a or b);
    layer0_outputs(560) <= not (a xor b);
    layer0_outputs(561) <= not a;
    layer0_outputs(562) <= not b;
    layer0_outputs(563) <= b and not a;
    layer0_outputs(564) <= not (a xor b);
    layer0_outputs(565) <= 1'b0;
    layer0_outputs(566) <= a xor b;
    layer0_outputs(567) <= not (a xor b);
    layer0_outputs(568) <= a or b;
    layer0_outputs(569) <= a;
    layer0_outputs(570) <= a or b;
    layer0_outputs(571) <= a or b;
    layer0_outputs(572) <= a;
    layer0_outputs(573) <= 1'b0;
    layer0_outputs(574) <= a or b;
    layer0_outputs(575) <= not b;
    layer0_outputs(576) <= a or b;
    layer0_outputs(577) <= not b or a;
    layer0_outputs(578) <= not (a or b);
    layer0_outputs(579) <= not b or a;
    layer0_outputs(580) <= a xor b;
    layer0_outputs(581) <= a and not b;
    layer0_outputs(582) <= not b;
    layer0_outputs(583) <= b and not a;
    layer0_outputs(584) <= not (a or b);
    layer0_outputs(585) <= a xor b;
    layer0_outputs(586) <= a or b;
    layer0_outputs(587) <= b and not a;
    layer0_outputs(588) <= 1'b0;
    layer0_outputs(589) <= not b or a;
    layer0_outputs(590) <= a and not b;
    layer0_outputs(591) <= not (a or b);
    layer0_outputs(592) <= not (a xor b);
    layer0_outputs(593) <= a xor b;
    layer0_outputs(594) <= not a;
    layer0_outputs(595) <= b and not a;
    layer0_outputs(596) <= not a or b;
    layer0_outputs(597) <= not (a or b);
    layer0_outputs(598) <= not (a or b);
    layer0_outputs(599) <= b;
    layer0_outputs(600) <= not (a or b);
    layer0_outputs(601) <= a;
    layer0_outputs(602) <= a or b;
    layer0_outputs(603) <= not b;
    layer0_outputs(604) <= b and not a;
    layer0_outputs(605) <= a or b;
    layer0_outputs(606) <= a or b;
    layer0_outputs(607) <= a;
    layer0_outputs(608) <= not (a or b);
    layer0_outputs(609) <= a and not b;
    layer0_outputs(610) <= a or b;
    layer0_outputs(611) <= b;
    layer0_outputs(612) <= 1'b1;
    layer0_outputs(613) <= not a;
    layer0_outputs(614) <= not (a or b);
    layer0_outputs(615) <= a or b;
    layer0_outputs(616) <= b;
    layer0_outputs(617) <= not (a xor b);
    layer0_outputs(618) <= a xor b;
    layer0_outputs(619) <= not (a xor b);
    layer0_outputs(620) <= not b or a;
    layer0_outputs(621) <= a and not b;
    layer0_outputs(622) <= b and not a;
    layer0_outputs(623) <= a or b;
    layer0_outputs(624) <= not (a or b);
    layer0_outputs(625) <= not b or a;
    layer0_outputs(626) <= not (a or b);
    layer0_outputs(627) <= not (a or b);
    layer0_outputs(628) <= not (a xor b);
    layer0_outputs(629) <= not a;
    layer0_outputs(630) <= not (a or b);
    layer0_outputs(631) <= a xor b;
    layer0_outputs(632) <= not b;
    layer0_outputs(633) <= not b or a;
    layer0_outputs(634) <= not a or b;
    layer0_outputs(635) <= not b or a;
    layer0_outputs(636) <= not (a or b);
    layer0_outputs(637) <= not (a xor b);
    layer0_outputs(638) <= not (a xor b);
    layer0_outputs(639) <= 1'b0;
    layer0_outputs(640) <= a xor b;
    layer0_outputs(641) <= not b;
    layer0_outputs(642) <= b;
    layer0_outputs(643) <= not b or a;
    layer0_outputs(644) <= a or b;
    layer0_outputs(645) <= a or b;
    layer0_outputs(646) <= a or b;
    layer0_outputs(647) <= not a;
    layer0_outputs(648) <= a or b;
    layer0_outputs(649) <= not a or b;
    layer0_outputs(650) <= a xor b;
    layer0_outputs(651) <= b and not a;
    layer0_outputs(652) <= not b or a;
    layer0_outputs(653) <= b and not a;
    layer0_outputs(654) <= b;
    layer0_outputs(655) <= not (a xor b);
    layer0_outputs(656) <= not a or b;
    layer0_outputs(657) <= 1'b0;
    layer0_outputs(658) <= 1'b1;
    layer0_outputs(659) <= not (a or b);
    layer0_outputs(660) <= not (a or b);
    layer0_outputs(661) <= a xor b;
    layer0_outputs(662) <= not b;
    layer0_outputs(663) <= not (a or b);
    layer0_outputs(664) <= not (a or b);
    layer0_outputs(665) <= not (a or b);
    layer0_outputs(666) <= not (a xor b);
    layer0_outputs(667) <= not b;
    layer0_outputs(668) <= not a or b;
    layer0_outputs(669) <= 1'b1;
    layer0_outputs(670) <= b;
    layer0_outputs(671) <= not a or b;
    layer0_outputs(672) <= b and not a;
    layer0_outputs(673) <= b and not a;
    layer0_outputs(674) <= a;
    layer0_outputs(675) <= not (a or b);
    layer0_outputs(676) <= 1'b0;
    layer0_outputs(677) <= a or b;
    layer0_outputs(678) <= not a or b;
    layer0_outputs(679) <= b and not a;
    layer0_outputs(680) <= a and not b;
    layer0_outputs(681) <= b;
    layer0_outputs(682) <= not (a or b);
    layer0_outputs(683) <= not a;
    layer0_outputs(684) <= a and not b;
    layer0_outputs(685) <= not (a or b);
    layer0_outputs(686) <= not (a or b);
    layer0_outputs(687) <= not a or b;
    layer0_outputs(688) <= a;
    layer0_outputs(689) <= not a or b;
    layer0_outputs(690) <= not (a xor b);
    layer0_outputs(691) <= not (a or b);
    layer0_outputs(692) <= not a;
    layer0_outputs(693) <= not (a xor b);
    layer0_outputs(694) <= a and not b;
    layer0_outputs(695) <= a or b;
    layer0_outputs(696) <= not a or b;
    layer0_outputs(697) <= not (a xor b);
    layer0_outputs(698) <= b;
    layer0_outputs(699) <= not (a xor b);
    layer0_outputs(700) <= not b;
    layer0_outputs(701) <= b and not a;
    layer0_outputs(702) <= a or b;
    layer0_outputs(703) <= b and not a;
    layer0_outputs(704) <= b;
    layer0_outputs(705) <= a or b;
    layer0_outputs(706) <= not (a xor b);
    layer0_outputs(707) <= b and not a;
    layer0_outputs(708) <= not (a or b);
    layer0_outputs(709) <= b and not a;
    layer0_outputs(710) <= not (a or b);
    layer0_outputs(711) <= a or b;
    layer0_outputs(712) <= not (a or b);
    layer0_outputs(713) <= not a;
    layer0_outputs(714) <= a or b;
    layer0_outputs(715) <= not a;
    layer0_outputs(716) <= b;
    layer0_outputs(717) <= not (a or b);
    layer0_outputs(718) <= a xor b;
    layer0_outputs(719) <= not a;
    layer0_outputs(720) <= b;
    layer0_outputs(721) <= b and not a;
    layer0_outputs(722) <= not b;
    layer0_outputs(723) <= 1'b1;
    layer0_outputs(724) <= not (a xor b);
    layer0_outputs(725) <= not a;
    layer0_outputs(726) <= not b or a;
    layer0_outputs(727) <= a;
    layer0_outputs(728) <= a xor b;
    layer0_outputs(729) <= 1'b1;
    layer0_outputs(730) <= not a;
    layer0_outputs(731) <= not (a and b);
    layer0_outputs(732) <= not a;
    layer0_outputs(733) <= a and b;
    layer0_outputs(734) <= b;
    layer0_outputs(735) <= not (a or b);
    layer0_outputs(736) <= a xor b;
    layer0_outputs(737) <= a xor b;
    layer0_outputs(738) <= not b;
    layer0_outputs(739) <= not b or a;
    layer0_outputs(740) <= a xor b;
    layer0_outputs(741) <= not (a or b);
    layer0_outputs(742) <= a or b;
    layer0_outputs(743) <= not a or b;
    layer0_outputs(744) <= not (a or b);
    layer0_outputs(745) <= not (a xor b);
    layer0_outputs(746) <= a or b;
    layer0_outputs(747) <= b and not a;
    layer0_outputs(748) <= a or b;
    layer0_outputs(749) <= not b or a;
    layer0_outputs(750) <= not (a or b);
    layer0_outputs(751) <= 1'b0;
    layer0_outputs(752) <= not (a or b);
    layer0_outputs(753) <= not (a or b);
    layer0_outputs(754) <= b and not a;
    layer0_outputs(755) <= b;
    layer0_outputs(756) <= b;
    layer0_outputs(757) <= a or b;
    layer0_outputs(758) <= not (a xor b);
    layer0_outputs(759) <= not (a xor b);
    layer0_outputs(760) <= a;
    layer0_outputs(761) <= a;
    layer0_outputs(762) <= a and b;
    layer0_outputs(763) <= a or b;
    layer0_outputs(764) <= a xor b;
    layer0_outputs(765) <= not (a or b);
    layer0_outputs(766) <= not b or a;
    layer0_outputs(767) <= not (a or b);
    layer0_outputs(768) <= 1'b1;
    layer0_outputs(769) <= a and not b;
    layer0_outputs(770) <= b;
    layer0_outputs(771) <= 1'b1;
    layer0_outputs(772) <= not a or b;
    layer0_outputs(773) <= a and not b;
    layer0_outputs(774) <= not a;
    layer0_outputs(775) <= a;
    layer0_outputs(776) <= a xor b;
    layer0_outputs(777) <= not b or a;
    layer0_outputs(778) <= not (a or b);
    layer0_outputs(779) <= a xor b;
    layer0_outputs(780) <= not (a or b);
    layer0_outputs(781) <= a and not b;
    layer0_outputs(782) <= not a;
    layer0_outputs(783) <= not a;
    layer0_outputs(784) <= a;
    layer0_outputs(785) <= not b or a;
    layer0_outputs(786) <= not b;
    layer0_outputs(787) <= not b;
    layer0_outputs(788) <= a xor b;
    layer0_outputs(789) <= 1'b0;
    layer0_outputs(790) <= not a or b;
    layer0_outputs(791) <= not a;
    layer0_outputs(792) <= not (a xor b);
    layer0_outputs(793) <= not (a or b);
    layer0_outputs(794) <= a or b;
    layer0_outputs(795) <= not (a or b);
    layer0_outputs(796) <= not (a xor b);
    layer0_outputs(797) <= a xor b;
    layer0_outputs(798) <= not (a or b);
    layer0_outputs(799) <= not b;
    layer0_outputs(800) <= 1'b1;
    layer0_outputs(801) <= b and not a;
    layer0_outputs(802) <= a and not b;
    layer0_outputs(803) <= not a or b;
    layer0_outputs(804) <= a xor b;
    layer0_outputs(805) <= a or b;
    layer0_outputs(806) <= a;
    layer0_outputs(807) <= a and not b;
    layer0_outputs(808) <= 1'b0;
    layer0_outputs(809) <= a or b;
    layer0_outputs(810) <= 1'b1;
    layer0_outputs(811) <= b;
    layer0_outputs(812) <= a or b;
    layer0_outputs(813) <= 1'b0;
    layer0_outputs(814) <= not b;
    layer0_outputs(815) <= a or b;
    layer0_outputs(816) <= not (a or b);
    layer0_outputs(817) <= a;
    layer0_outputs(818) <= not b;
    layer0_outputs(819) <= a or b;
    layer0_outputs(820) <= not (a xor b);
    layer0_outputs(821) <= a or b;
    layer0_outputs(822) <= 1'b1;
    layer0_outputs(823) <= a or b;
    layer0_outputs(824) <= not a;
    layer0_outputs(825) <= 1'b0;
    layer0_outputs(826) <= a;
    layer0_outputs(827) <= a xor b;
    layer0_outputs(828) <= not (a or b);
    layer0_outputs(829) <= a or b;
    layer0_outputs(830) <= not a;
    layer0_outputs(831) <= not b or a;
    layer0_outputs(832) <= not (a or b);
    layer0_outputs(833) <= not a or b;
    layer0_outputs(834) <= not a or b;
    layer0_outputs(835) <= b;
    layer0_outputs(836) <= not (a xor b);
    layer0_outputs(837) <= a;
    layer0_outputs(838) <= a;
    layer0_outputs(839) <= not a;
    layer0_outputs(840) <= a xor b;
    layer0_outputs(841) <= not b or a;
    layer0_outputs(842) <= not (a or b);
    layer0_outputs(843) <= not b;
    layer0_outputs(844) <= a or b;
    layer0_outputs(845) <= not b or a;
    layer0_outputs(846) <= not b;
    layer0_outputs(847) <= a and not b;
    layer0_outputs(848) <= 1'b0;
    layer0_outputs(849) <= a and b;
    layer0_outputs(850) <= not b;
    layer0_outputs(851) <= not (a xor b);
    layer0_outputs(852) <= not b or a;
    layer0_outputs(853) <= not b;
    layer0_outputs(854) <= not (a or b);
    layer0_outputs(855) <= a;
    layer0_outputs(856) <= not (a xor b);
    layer0_outputs(857) <= not (a xor b);
    layer0_outputs(858) <= a and b;
    layer0_outputs(859) <= 1'b1;
    layer0_outputs(860) <= b and not a;
    layer0_outputs(861) <= b and not a;
    layer0_outputs(862) <= not b;
    layer0_outputs(863) <= not (a or b);
    layer0_outputs(864) <= not (a or b);
    layer0_outputs(865) <= a or b;
    layer0_outputs(866) <= b and not a;
    layer0_outputs(867) <= not b or a;
    layer0_outputs(868) <= b and not a;
    layer0_outputs(869) <= b;
    layer0_outputs(870) <= not (a or b);
    layer0_outputs(871) <= a xor b;
    layer0_outputs(872) <= b;
    layer0_outputs(873) <= a or b;
    layer0_outputs(874) <= not b or a;
    layer0_outputs(875) <= not (a and b);
    layer0_outputs(876) <= not (a or b);
    layer0_outputs(877) <= not b;
    layer0_outputs(878) <= not (a or b);
    layer0_outputs(879) <= a xor b;
    layer0_outputs(880) <= a and not b;
    layer0_outputs(881) <= a and not b;
    layer0_outputs(882) <= a xor b;
    layer0_outputs(883) <= not a or b;
    layer0_outputs(884) <= b and not a;
    layer0_outputs(885) <= a xor b;
    layer0_outputs(886) <= not b;
    layer0_outputs(887) <= a xor b;
    layer0_outputs(888) <= 1'b1;
    layer0_outputs(889) <= a xor b;
    layer0_outputs(890) <= not a;
    layer0_outputs(891) <= a and not b;
    layer0_outputs(892) <= not a or b;
    layer0_outputs(893) <= not a or b;
    layer0_outputs(894) <= a and not b;
    layer0_outputs(895) <= not b;
    layer0_outputs(896) <= a or b;
    layer0_outputs(897) <= not a or b;
    layer0_outputs(898) <= not b;
    layer0_outputs(899) <= a xor b;
    layer0_outputs(900) <= not (a and b);
    layer0_outputs(901) <= a or b;
    layer0_outputs(902) <= not b;
    layer0_outputs(903) <= not (a or b);
    layer0_outputs(904) <= a or b;
    layer0_outputs(905) <= a or b;
    layer0_outputs(906) <= a and not b;
    layer0_outputs(907) <= not a;
    layer0_outputs(908) <= not (a or b);
    layer0_outputs(909) <= not (a xor b);
    layer0_outputs(910) <= b;
    layer0_outputs(911) <= not b;
    layer0_outputs(912) <= not b;
    layer0_outputs(913) <= a or b;
    layer0_outputs(914) <= b;
    layer0_outputs(915) <= not b;
    layer0_outputs(916) <= not b or a;
    layer0_outputs(917) <= not (a or b);
    layer0_outputs(918) <= b;
    layer0_outputs(919) <= a;
    layer0_outputs(920) <= a or b;
    layer0_outputs(921) <= a;
    layer0_outputs(922) <= not a;
    layer0_outputs(923) <= b;
    layer0_outputs(924) <= not b or a;
    layer0_outputs(925) <= a and not b;
    layer0_outputs(926) <= not a;
    layer0_outputs(927) <= a or b;
    layer0_outputs(928) <= not a or b;
    layer0_outputs(929) <= not (a xor b);
    layer0_outputs(930) <= not b;
    layer0_outputs(931) <= a and not b;
    layer0_outputs(932) <= not (a or b);
    layer0_outputs(933) <= a and not b;
    layer0_outputs(934) <= not a or b;
    layer0_outputs(935) <= a or b;
    layer0_outputs(936) <= not (a xor b);
    layer0_outputs(937) <= not b;
    layer0_outputs(938) <= not b or a;
    layer0_outputs(939) <= a or b;
    layer0_outputs(940) <= not a;
    layer0_outputs(941) <= a xor b;
    layer0_outputs(942) <= not (a or b);
    layer0_outputs(943) <= b and not a;
    layer0_outputs(944) <= a and not b;
    layer0_outputs(945) <= not (a xor b);
    layer0_outputs(946) <= not b or a;
    layer0_outputs(947) <= not a or b;
    layer0_outputs(948) <= b and not a;
    layer0_outputs(949) <= a;
    layer0_outputs(950) <= not (a or b);
    layer0_outputs(951) <= not (a and b);
    layer0_outputs(952) <= b and not a;
    layer0_outputs(953) <= not a;
    layer0_outputs(954) <= not a or b;
    layer0_outputs(955) <= a xor b;
    layer0_outputs(956) <= not (a or b);
    layer0_outputs(957) <= a and not b;
    layer0_outputs(958) <= a and not b;
    layer0_outputs(959) <= a;
    layer0_outputs(960) <= not (a and b);
    layer0_outputs(961) <= a and not b;
    layer0_outputs(962) <= not a or b;
    layer0_outputs(963) <= a;
    layer0_outputs(964) <= a or b;
    layer0_outputs(965) <= not a or b;
    layer0_outputs(966) <= b;
    layer0_outputs(967) <= 1'b0;
    layer0_outputs(968) <= not (a xor b);
    layer0_outputs(969) <= not (a or b);
    layer0_outputs(970) <= not (a or b);
    layer0_outputs(971) <= a xor b;
    layer0_outputs(972) <= not b or a;
    layer0_outputs(973) <= a;
    layer0_outputs(974) <= not (a or b);
    layer0_outputs(975) <= not (a and b);
    layer0_outputs(976) <= not (a xor b);
    layer0_outputs(977) <= b;
    layer0_outputs(978) <= b and not a;
    layer0_outputs(979) <= not b or a;
    layer0_outputs(980) <= not b or a;
    layer0_outputs(981) <= not b;
    layer0_outputs(982) <= a and not b;
    layer0_outputs(983) <= not b;
    layer0_outputs(984) <= a or b;
    layer0_outputs(985) <= a or b;
    layer0_outputs(986) <= not b or a;
    layer0_outputs(987) <= a;
    layer0_outputs(988) <= a xor b;
    layer0_outputs(989) <= not a;
    layer0_outputs(990) <= not (a or b);
    layer0_outputs(991) <= not (a or b);
    layer0_outputs(992) <= not (a xor b);
    layer0_outputs(993) <= 1'b1;
    layer0_outputs(994) <= b and not a;
    layer0_outputs(995) <= a or b;
    layer0_outputs(996) <= a or b;
    layer0_outputs(997) <= not (a and b);
    layer0_outputs(998) <= not (a xor b);
    layer0_outputs(999) <= 1'b0;
    layer0_outputs(1000) <= not a or b;
    layer0_outputs(1001) <= b and not a;
    layer0_outputs(1002) <= not a;
    layer0_outputs(1003) <= a or b;
    layer0_outputs(1004) <= a xor b;
    layer0_outputs(1005) <= not a;
    layer0_outputs(1006) <= not a;
    layer0_outputs(1007) <= a;
    layer0_outputs(1008) <= not b or a;
    layer0_outputs(1009) <= a or b;
    layer0_outputs(1010) <= not (a or b);
    layer0_outputs(1011) <= a or b;
    layer0_outputs(1012) <= a xor b;
    layer0_outputs(1013) <= not (a and b);
    layer0_outputs(1014) <= a;
    layer0_outputs(1015) <= b;
    layer0_outputs(1016) <= a xor b;
    layer0_outputs(1017) <= not a;
    layer0_outputs(1018) <= not (a or b);
    layer0_outputs(1019) <= not b or a;
    layer0_outputs(1020) <= a xor b;
    layer0_outputs(1021) <= not a or b;
    layer0_outputs(1022) <= not (a xor b);
    layer0_outputs(1023) <= b and not a;
    layer0_outputs(1024) <= not b;
    layer0_outputs(1025) <= not (a xor b);
    layer0_outputs(1026) <= not b;
    layer0_outputs(1027) <= not b or a;
    layer0_outputs(1028) <= b;
    layer0_outputs(1029) <= b and not a;
    layer0_outputs(1030) <= a xor b;
    layer0_outputs(1031) <= 1'b0;
    layer0_outputs(1032) <= not (a or b);
    layer0_outputs(1033) <= a;
    layer0_outputs(1034) <= not (a and b);
    layer0_outputs(1035) <= a xor b;
    layer0_outputs(1036) <= not b;
    layer0_outputs(1037) <= not (a or b);
    layer0_outputs(1038) <= not (a xor b);
    layer0_outputs(1039) <= 1'b1;
    layer0_outputs(1040) <= not (a and b);
    layer0_outputs(1041) <= b and not a;
    layer0_outputs(1042) <= not (a or b);
    layer0_outputs(1043) <= not b;
    layer0_outputs(1044) <= b;
    layer0_outputs(1045) <= not a or b;
    layer0_outputs(1046) <= a and not b;
    layer0_outputs(1047) <= b and not a;
    layer0_outputs(1048) <= not b;
    layer0_outputs(1049) <= not (a xor b);
    layer0_outputs(1050) <= a xor b;
    layer0_outputs(1051) <= not (a xor b);
    layer0_outputs(1052) <= b;
    layer0_outputs(1053) <= a or b;
    layer0_outputs(1054) <= b and not a;
    layer0_outputs(1055) <= a or b;
    layer0_outputs(1056) <= a and not b;
    layer0_outputs(1057) <= b and not a;
    layer0_outputs(1058) <= not b;
    layer0_outputs(1059) <= a or b;
    layer0_outputs(1060) <= not (a xor b);
    layer0_outputs(1061) <= a;
    layer0_outputs(1062) <= not (a or b);
    layer0_outputs(1063) <= a and not b;
    layer0_outputs(1064) <= b and not a;
    layer0_outputs(1065) <= not b or a;
    layer0_outputs(1066) <= b;
    layer0_outputs(1067) <= a xor b;
    layer0_outputs(1068) <= a xor b;
    layer0_outputs(1069) <= b and not a;
    layer0_outputs(1070) <= not b or a;
    layer0_outputs(1071) <= not (a xor b);
    layer0_outputs(1072) <= a or b;
    layer0_outputs(1073) <= a xor b;
    layer0_outputs(1074) <= a and not b;
    layer0_outputs(1075) <= b and not a;
    layer0_outputs(1076) <= b;
    layer0_outputs(1077) <= not (a or b);
    layer0_outputs(1078) <= not a or b;
    layer0_outputs(1079) <= not (a or b);
    layer0_outputs(1080) <= not b;
    layer0_outputs(1081) <= a or b;
    layer0_outputs(1082) <= a or b;
    layer0_outputs(1083) <= not (a or b);
    layer0_outputs(1084) <= not b or a;
    layer0_outputs(1085) <= 1'b0;
    layer0_outputs(1086) <= a and b;
    layer0_outputs(1087) <= a xor b;
    layer0_outputs(1088) <= b and not a;
    layer0_outputs(1089) <= not (a or b);
    layer0_outputs(1090) <= b;
    layer0_outputs(1091) <= a and not b;
    layer0_outputs(1092) <= a and not b;
    layer0_outputs(1093) <= not (a and b);
    layer0_outputs(1094) <= not a or b;
    layer0_outputs(1095) <= a xor b;
    layer0_outputs(1096) <= a and not b;
    layer0_outputs(1097) <= b;
    layer0_outputs(1098) <= not (a xor b);
    layer0_outputs(1099) <= not a;
    layer0_outputs(1100) <= a or b;
    layer0_outputs(1101) <= a xor b;
    layer0_outputs(1102) <= a and not b;
    layer0_outputs(1103) <= not a;
    layer0_outputs(1104) <= a or b;
    layer0_outputs(1105) <= not (a xor b);
    layer0_outputs(1106) <= not (a or b);
    layer0_outputs(1107) <= not (a or b);
    layer0_outputs(1108) <= not (a xor b);
    layer0_outputs(1109) <= not (a xor b);
    layer0_outputs(1110) <= a or b;
    layer0_outputs(1111) <= a and not b;
    layer0_outputs(1112) <= b and not a;
    layer0_outputs(1113) <= b and not a;
    layer0_outputs(1114) <= a xor b;
    layer0_outputs(1115) <= not b or a;
    layer0_outputs(1116) <= not a;
    layer0_outputs(1117) <= b and not a;
    layer0_outputs(1118) <= b and not a;
    layer0_outputs(1119) <= a xor b;
    layer0_outputs(1120) <= a xor b;
    layer0_outputs(1121) <= not (a or b);
    layer0_outputs(1122) <= a or b;
    layer0_outputs(1123) <= not (a or b);
    layer0_outputs(1124) <= not a;
    layer0_outputs(1125) <= not b or a;
    layer0_outputs(1126) <= 1'b1;
    layer0_outputs(1127) <= a or b;
    layer0_outputs(1128) <= a;
    layer0_outputs(1129) <= not b;
    layer0_outputs(1130) <= not b;
    layer0_outputs(1131) <= not (a and b);
    layer0_outputs(1132) <= a xor b;
    layer0_outputs(1133) <= not b or a;
    layer0_outputs(1134) <= not (a or b);
    layer0_outputs(1135) <= not b;
    layer0_outputs(1136) <= not (a xor b);
    layer0_outputs(1137) <= not (a xor b);
    layer0_outputs(1138) <= a or b;
    layer0_outputs(1139) <= b and not a;
    layer0_outputs(1140) <= a or b;
    layer0_outputs(1141) <= not (a xor b);
    layer0_outputs(1142) <= not a;
    layer0_outputs(1143) <= a;
    layer0_outputs(1144) <= not a;
    layer0_outputs(1145) <= a or b;
    layer0_outputs(1146) <= a or b;
    layer0_outputs(1147) <= not a or b;
    layer0_outputs(1148) <= not b;
    layer0_outputs(1149) <= a or b;
    layer0_outputs(1150) <= a and b;
    layer0_outputs(1151) <= not (a and b);
    layer0_outputs(1152) <= a and not b;
    layer0_outputs(1153) <= not a;
    layer0_outputs(1154) <= a and not b;
    layer0_outputs(1155) <= not b or a;
    layer0_outputs(1156) <= not (a xor b);
    layer0_outputs(1157) <= a or b;
    layer0_outputs(1158) <= b;
    layer0_outputs(1159) <= a and b;
    layer0_outputs(1160) <= b;
    layer0_outputs(1161) <= not a or b;
    layer0_outputs(1162) <= b;
    layer0_outputs(1163) <= not (a xor b);
    layer0_outputs(1164) <= a or b;
    layer0_outputs(1165) <= not a or b;
    layer0_outputs(1166) <= a;
    layer0_outputs(1167) <= not b;
    layer0_outputs(1168) <= not (a or b);
    layer0_outputs(1169) <= not (a or b);
    layer0_outputs(1170) <= 1'b1;
    layer0_outputs(1171) <= b and not a;
    layer0_outputs(1172) <= not (a or b);
    layer0_outputs(1173) <= a or b;
    layer0_outputs(1174) <= not (a or b);
    layer0_outputs(1175) <= not a or b;
    layer0_outputs(1176) <= 1'b0;
    layer0_outputs(1177) <= not b or a;
    layer0_outputs(1178) <= not b;
    layer0_outputs(1179) <= not a;
    layer0_outputs(1180) <= not (a xor b);
    layer0_outputs(1181) <= not a;
    layer0_outputs(1182) <= not b or a;
    layer0_outputs(1183) <= a and not b;
    layer0_outputs(1184) <= not a;
    layer0_outputs(1185) <= not a;
    layer0_outputs(1186) <= a xor b;
    layer0_outputs(1187) <= not (a or b);
    layer0_outputs(1188) <= not b;
    layer0_outputs(1189) <= not b or a;
    layer0_outputs(1190) <= a or b;
    layer0_outputs(1191) <= not a;
    layer0_outputs(1192) <= not (a or b);
    layer0_outputs(1193) <= not (a or b);
    layer0_outputs(1194) <= not a or b;
    layer0_outputs(1195) <= a;
    layer0_outputs(1196) <= a or b;
    layer0_outputs(1197) <= a or b;
    layer0_outputs(1198) <= 1'b1;
    layer0_outputs(1199) <= not (a and b);
    layer0_outputs(1200) <= not a or b;
    layer0_outputs(1201) <= a xor b;
    layer0_outputs(1202) <= not b;
    layer0_outputs(1203) <= a xor b;
    layer0_outputs(1204) <= a xor b;
    layer0_outputs(1205) <= a or b;
    layer0_outputs(1206) <= not a;
    layer0_outputs(1207) <= b;
    layer0_outputs(1208) <= a or b;
    layer0_outputs(1209) <= not b or a;
    layer0_outputs(1210) <= a or b;
    layer0_outputs(1211) <= b;
    layer0_outputs(1212) <= a;
    layer0_outputs(1213) <= 1'b0;
    layer0_outputs(1214) <= not b;
    layer0_outputs(1215) <= not b or a;
    layer0_outputs(1216) <= not (a or b);
    layer0_outputs(1217) <= a and not b;
    layer0_outputs(1218) <= not (a xor b);
    layer0_outputs(1219) <= not a or b;
    layer0_outputs(1220) <= not b;
    layer0_outputs(1221) <= a or b;
    layer0_outputs(1222) <= not (a or b);
    layer0_outputs(1223) <= not a;
    layer0_outputs(1224) <= not a;
    layer0_outputs(1225) <= not (a xor b);
    layer0_outputs(1226) <= a and not b;
    layer0_outputs(1227) <= not b or a;
    layer0_outputs(1228) <= not (a and b);
    layer0_outputs(1229) <= not (a or b);
    layer0_outputs(1230) <= a xor b;
    layer0_outputs(1231) <= 1'b0;
    layer0_outputs(1232) <= not (a xor b);
    layer0_outputs(1233) <= a and b;
    layer0_outputs(1234) <= not b;
    layer0_outputs(1235) <= a;
    layer0_outputs(1236) <= not b;
    layer0_outputs(1237) <= not (a xor b);
    layer0_outputs(1238) <= 1'b1;
    layer0_outputs(1239) <= a or b;
    layer0_outputs(1240) <= a or b;
    layer0_outputs(1241) <= a and b;
    layer0_outputs(1242) <= b;
    layer0_outputs(1243) <= a or b;
    layer0_outputs(1244) <= not b or a;
    layer0_outputs(1245) <= not (a xor b);
    layer0_outputs(1246) <= a;
    layer0_outputs(1247) <= 1'b0;
    layer0_outputs(1248) <= a or b;
    layer0_outputs(1249) <= not b;
    layer0_outputs(1250) <= not (a or b);
    layer0_outputs(1251) <= a xor b;
    layer0_outputs(1252) <= not (a xor b);
    layer0_outputs(1253) <= not b;
    layer0_outputs(1254) <= not b or a;
    layer0_outputs(1255) <= a or b;
    layer0_outputs(1256) <= not a or b;
    layer0_outputs(1257) <= a and not b;
    layer0_outputs(1258) <= a and not b;
    layer0_outputs(1259) <= a or b;
    layer0_outputs(1260) <= not b or a;
    layer0_outputs(1261) <= not b;
    layer0_outputs(1262) <= not (a xor b);
    layer0_outputs(1263) <= a and not b;
    layer0_outputs(1264) <= not b;
    layer0_outputs(1265) <= not (a xor b);
    layer0_outputs(1266) <= a and not b;
    layer0_outputs(1267) <= a xor b;
    layer0_outputs(1268) <= a and not b;
    layer0_outputs(1269) <= not (a xor b);
    layer0_outputs(1270) <= not b;
    layer0_outputs(1271) <= a;
    layer0_outputs(1272) <= not (a xor b);
    layer0_outputs(1273) <= a xor b;
    layer0_outputs(1274) <= a or b;
    layer0_outputs(1275) <= not a;
    layer0_outputs(1276) <= not b or a;
    layer0_outputs(1277) <= a or b;
    layer0_outputs(1278) <= not (a or b);
    layer0_outputs(1279) <= b;
    layer0_outputs(1280) <= a and not b;
    layer0_outputs(1281) <= not (a and b);
    layer0_outputs(1282) <= b and not a;
    layer0_outputs(1283) <= not (a xor b);
    layer0_outputs(1284) <= not (a or b);
    layer0_outputs(1285) <= b;
    layer0_outputs(1286) <= a and not b;
    layer0_outputs(1287) <= b and not a;
    layer0_outputs(1288) <= a;
    layer0_outputs(1289) <= not b or a;
    layer0_outputs(1290) <= not b;
    layer0_outputs(1291) <= not a;
    layer0_outputs(1292) <= b;
    layer0_outputs(1293) <= not b;
    layer0_outputs(1294) <= 1'b0;
    layer0_outputs(1295) <= b and not a;
    layer0_outputs(1296) <= not (a xor b);
    layer0_outputs(1297) <= a;
    layer0_outputs(1298) <= not a;
    layer0_outputs(1299) <= a or b;
    layer0_outputs(1300) <= not b;
    layer0_outputs(1301) <= not (a xor b);
    layer0_outputs(1302) <= a or b;
    layer0_outputs(1303) <= not a or b;
    layer0_outputs(1304) <= a or b;
    layer0_outputs(1305) <= not b;
    layer0_outputs(1306) <= not b or a;
    layer0_outputs(1307) <= not (a xor b);
    layer0_outputs(1308) <= a xor b;
    layer0_outputs(1309) <= not (a or b);
    layer0_outputs(1310) <= not (a or b);
    layer0_outputs(1311) <= not (a or b);
    layer0_outputs(1312) <= not (a or b);
    layer0_outputs(1313) <= a;
    layer0_outputs(1314) <= 1'b0;
    layer0_outputs(1315) <= not (a and b);
    layer0_outputs(1316) <= b and not a;
    layer0_outputs(1317) <= a and not b;
    layer0_outputs(1318) <= a xor b;
    layer0_outputs(1319) <= not (a and b);
    layer0_outputs(1320) <= not (a or b);
    layer0_outputs(1321) <= not a;
    layer0_outputs(1322) <= not (a and b);
    layer0_outputs(1323) <= a or b;
    layer0_outputs(1324) <= a and not b;
    layer0_outputs(1325) <= a or b;
    layer0_outputs(1326) <= a xor b;
    layer0_outputs(1327) <= a;
    layer0_outputs(1328) <= a and not b;
    layer0_outputs(1329) <= not (a or b);
    layer0_outputs(1330) <= not (a xor b);
    layer0_outputs(1331) <= a xor b;
    layer0_outputs(1332) <= not a or b;
    layer0_outputs(1333) <= a and not b;
    layer0_outputs(1334) <= not b;
    layer0_outputs(1335) <= not a or b;
    layer0_outputs(1336) <= not (a xor b);
    layer0_outputs(1337) <= b;
    layer0_outputs(1338) <= not b;
    layer0_outputs(1339) <= not (a or b);
    layer0_outputs(1340) <= a xor b;
    layer0_outputs(1341) <= a or b;
    layer0_outputs(1342) <= a and not b;
    layer0_outputs(1343) <= not (a or b);
    layer0_outputs(1344) <= not (a and b);
    layer0_outputs(1345) <= a xor b;
    layer0_outputs(1346) <= a or b;
    layer0_outputs(1347) <= a;
    layer0_outputs(1348) <= not (a xor b);
    layer0_outputs(1349) <= b;
    layer0_outputs(1350) <= not b;
    layer0_outputs(1351) <= not a;
    layer0_outputs(1352) <= a or b;
    layer0_outputs(1353) <= b;
    layer0_outputs(1354) <= a or b;
    layer0_outputs(1355) <= b;
    layer0_outputs(1356) <= a or b;
    layer0_outputs(1357) <= b;
    layer0_outputs(1358) <= a and not b;
    layer0_outputs(1359) <= a or b;
    layer0_outputs(1360) <= not (a or b);
    layer0_outputs(1361) <= a;
    layer0_outputs(1362) <= not b;
    layer0_outputs(1363) <= not a;
    layer0_outputs(1364) <= not a;
    layer0_outputs(1365) <= not a;
    layer0_outputs(1366) <= b and not a;
    layer0_outputs(1367) <= a xor b;
    layer0_outputs(1368) <= 1'b0;
    layer0_outputs(1369) <= a;
    layer0_outputs(1370) <= b;
    layer0_outputs(1371) <= a or b;
    layer0_outputs(1372) <= a and not b;
    layer0_outputs(1373) <= a and not b;
    layer0_outputs(1374) <= a and not b;
    layer0_outputs(1375) <= not a;
    layer0_outputs(1376) <= b and not a;
    layer0_outputs(1377) <= a or b;
    layer0_outputs(1378) <= not b;
    layer0_outputs(1379) <= b;
    layer0_outputs(1380) <= not a;
    layer0_outputs(1381) <= b and not a;
    layer0_outputs(1382) <= a;
    layer0_outputs(1383) <= a and not b;
    layer0_outputs(1384) <= not a;
    layer0_outputs(1385) <= not a;
    layer0_outputs(1386) <= a or b;
    layer0_outputs(1387) <= not b;
    layer0_outputs(1388) <= a xor b;
    layer0_outputs(1389) <= a xor b;
    layer0_outputs(1390) <= 1'b0;
    layer0_outputs(1391) <= b;
    layer0_outputs(1392) <= a or b;
    layer0_outputs(1393) <= not (a or b);
    layer0_outputs(1394) <= not (a and b);
    layer0_outputs(1395) <= not (a xor b);
    layer0_outputs(1396) <= a or b;
    layer0_outputs(1397) <= not (a xor b);
    layer0_outputs(1398) <= not (a or b);
    layer0_outputs(1399) <= not a;
    layer0_outputs(1400) <= a or b;
    layer0_outputs(1401) <= a and not b;
    layer0_outputs(1402) <= not b;
    layer0_outputs(1403) <= a and not b;
    layer0_outputs(1404) <= not (a and b);
    layer0_outputs(1405) <= not (a or b);
    layer0_outputs(1406) <= not (a or b);
    layer0_outputs(1407) <= b;
    layer0_outputs(1408) <= not (a or b);
    layer0_outputs(1409) <= a or b;
    layer0_outputs(1410) <= not (a or b);
    layer0_outputs(1411) <= not a;
    layer0_outputs(1412) <= a and b;
    layer0_outputs(1413) <= not a;
    layer0_outputs(1414) <= not (a xor b);
    layer0_outputs(1415) <= 1'b1;
    layer0_outputs(1416) <= not b or a;
    layer0_outputs(1417) <= not (a or b);
    layer0_outputs(1418) <= a or b;
    layer0_outputs(1419) <= not (a and b);
    layer0_outputs(1420) <= not b or a;
    layer0_outputs(1421) <= b;
    layer0_outputs(1422) <= not (a or b);
    layer0_outputs(1423) <= not (a or b);
    layer0_outputs(1424) <= a or b;
    layer0_outputs(1425) <= not (a or b);
    layer0_outputs(1426) <= not a or b;
    layer0_outputs(1427) <= not a or b;
    layer0_outputs(1428) <= not b or a;
    layer0_outputs(1429) <= not (a xor b);
    layer0_outputs(1430) <= not b or a;
    layer0_outputs(1431) <= a or b;
    layer0_outputs(1432) <= not (a xor b);
    layer0_outputs(1433) <= a or b;
    layer0_outputs(1434) <= a and not b;
    layer0_outputs(1435) <= 1'b0;
    layer0_outputs(1436) <= not (a or b);
    layer0_outputs(1437) <= not b;
    layer0_outputs(1438) <= not a or b;
    layer0_outputs(1439) <= a and not b;
    layer0_outputs(1440) <= a or b;
    layer0_outputs(1441) <= a xor b;
    layer0_outputs(1442) <= a xor b;
    layer0_outputs(1443) <= not a or b;
    layer0_outputs(1444) <= a xor b;
    layer0_outputs(1445) <= not (a or b);
    layer0_outputs(1446) <= b and not a;
    layer0_outputs(1447) <= a or b;
    layer0_outputs(1448) <= not b;
    layer0_outputs(1449) <= b and not a;
    layer0_outputs(1450) <= not b or a;
    layer0_outputs(1451) <= not (a or b);
    layer0_outputs(1452) <= not a or b;
    layer0_outputs(1453) <= b;
    layer0_outputs(1454) <= a xor b;
    layer0_outputs(1455) <= not (a xor b);
    layer0_outputs(1456) <= not (a xor b);
    layer0_outputs(1457) <= not b or a;
    layer0_outputs(1458) <= a or b;
    layer0_outputs(1459) <= not (a or b);
    layer0_outputs(1460) <= not (a and b);
    layer0_outputs(1461) <= a and not b;
    layer0_outputs(1462) <= not (a xor b);
    layer0_outputs(1463) <= a xor b;
    layer0_outputs(1464) <= not b or a;
    layer0_outputs(1465) <= not (a or b);
    layer0_outputs(1466) <= a;
    layer0_outputs(1467) <= a;
    layer0_outputs(1468) <= a xor b;
    layer0_outputs(1469) <= not a;
    layer0_outputs(1470) <= not (a xor b);
    layer0_outputs(1471) <= a and not b;
    layer0_outputs(1472) <= not (a or b);
    layer0_outputs(1473) <= not b;
    layer0_outputs(1474) <= a and not b;
    layer0_outputs(1475) <= b;
    layer0_outputs(1476) <= not b or a;
    layer0_outputs(1477) <= not (a and b);
    layer0_outputs(1478) <= a and not b;
    layer0_outputs(1479) <= a xor b;
    layer0_outputs(1480) <= not (a or b);
    layer0_outputs(1481) <= not (a xor b);
    layer0_outputs(1482) <= a or b;
    layer0_outputs(1483) <= 1'b1;
    layer0_outputs(1484) <= a or b;
    layer0_outputs(1485) <= a or b;
    layer0_outputs(1486) <= not b or a;
    layer0_outputs(1487) <= b;
    layer0_outputs(1488) <= a or b;
    layer0_outputs(1489) <= not a;
    layer0_outputs(1490) <= not (a xor b);
    layer0_outputs(1491) <= not a or b;
    layer0_outputs(1492) <= a xor b;
    layer0_outputs(1493) <= a or b;
    layer0_outputs(1494) <= not a;
    layer0_outputs(1495) <= not (a or b);
    layer0_outputs(1496) <= not (a xor b);
    layer0_outputs(1497) <= a and not b;
    layer0_outputs(1498) <= not a;
    layer0_outputs(1499) <= a xor b;
    layer0_outputs(1500) <= a and not b;
    layer0_outputs(1501) <= not b;
    layer0_outputs(1502) <= not (a or b);
    layer0_outputs(1503) <= not (a or b);
    layer0_outputs(1504) <= b;
    layer0_outputs(1505) <= not a;
    layer0_outputs(1506) <= a or b;
    layer0_outputs(1507) <= a or b;
    layer0_outputs(1508) <= a or b;
    layer0_outputs(1509) <= not (a and b);
    layer0_outputs(1510) <= not b;
    layer0_outputs(1511) <= not (a xor b);
    layer0_outputs(1512) <= a xor b;
    layer0_outputs(1513) <= not (a and b);
    layer0_outputs(1514) <= not (a or b);
    layer0_outputs(1515) <= a;
    layer0_outputs(1516) <= a xor b;
    layer0_outputs(1517) <= not b or a;
    layer0_outputs(1518) <= 1'b0;
    layer0_outputs(1519) <= not a;
    layer0_outputs(1520) <= not (a xor b);
    layer0_outputs(1521) <= not b;
    layer0_outputs(1522) <= b;
    layer0_outputs(1523) <= a and not b;
    layer0_outputs(1524) <= 1'b0;
    layer0_outputs(1525) <= not a;
    layer0_outputs(1526) <= a and not b;
    layer0_outputs(1527) <= not a;
    layer0_outputs(1528) <= not b or a;
    layer0_outputs(1529) <= a;
    layer0_outputs(1530) <= not b or a;
    layer0_outputs(1531) <= not (a or b);
    layer0_outputs(1532) <= a or b;
    layer0_outputs(1533) <= b and not a;
    layer0_outputs(1534) <= a or b;
    layer0_outputs(1535) <= not b;
    layer0_outputs(1536) <= a xor b;
    layer0_outputs(1537) <= a or b;
    layer0_outputs(1538) <= b and not a;
    layer0_outputs(1539) <= not (a xor b);
    layer0_outputs(1540) <= a xor b;
    layer0_outputs(1541) <= not b;
    layer0_outputs(1542) <= not (a or b);
    layer0_outputs(1543) <= a or b;
    layer0_outputs(1544) <= a or b;
    layer0_outputs(1545) <= a or b;
    layer0_outputs(1546) <= b and not a;
    layer0_outputs(1547) <= a;
    layer0_outputs(1548) <= a and not b;
    layer0_outputs(1549) <= a or b;
    layer0_outputs(1550) <= not (a xor b);
    layer0_outputs(1551) <= b and not a;
    layer0_outputs(1552) <= not b;
    layer0_outputs(1553) <= not (a xor b);
    layer0_outputs(1554) <= b;
    layer0_outputs(1555) <= b;
    layer0_outputs(1556) <= a xor b;
    layer0_outputs(1557) <= a xor b;
    layer0_outputs(1558) <= a and not b;
    layer0_outputs(1559) <= not (a or b);
    layer0_outputs(1560) <= not a or b;
    layer0_outputs(1561) <= not a or b;
    layer0_outputs(1562) <= b;
    layer0_outputs(1563) <= a or b;
    layer0_outputs(1564) <= a and not b;
    layer0_outputs(1565) <= not (a or b);
    layer0_outputs(1566) <= a xor b;
    layer0_outputs(1567) <= not a or b;
    layer0_outputs(1568) <= not b or a;
    layer0_outputs(1569) <= 1'b1;
    layer0_outputs(1570) <= not a;
    layer0_outputs(1571) <= a xor b;
    layer0_outputs(1572) <= not b or a;
    layer0_outputs(1573) <= 1'b0;
    layer0_outputs(1574) <= not (a or b);
    layer0_outputs(1575) <= not (a and b);
    layer0_outputs(1576) <= a and not b;
    layer0_outputs(1577) <= b;
    layer0_outputs(1578) <= not (a or b);
    layer0_outputs(1579) <= not (a or b);
    layer0_outputs(1580) <= not (a xor b);
    layer0_outputs(1581) <= a or b;
    layer0_outputs(1582) <= b and not a;
    layer0_outputs(1583) <= a or b;
    layer0_outputs(1584) <= not (a or b);
    layer0_outputs(1585) <= b;
    layer0_outputs(1586) <= a and b;
    layer0_outputs(1587) <= a and not b;
    layer0_outputs(1588) <= a or b;
    layer0_outputs(1589) <= 1'b0;
    layer0_outputs(1590) <= a or b;
    layer0_outputs(1591) <= a and not b;
    layer0_outputs(1592) <= a or b;
    layer0_outputs(1593) <= a or b;
    layer0_outputs(1594) <= b;
    layer0_outputs(1595) <= a xor b;
    layer0_outputs(1596) <= a xor b;
    layer0_outputs(1597) <= not (a xor b);
    layer0_outputs(1598) <= not a or b;
    layer0_outputs(1599) <= not a;
    layer0_outputs(1600) <= not a or b;
    layer0_outputs(1601) <= not (a xor b);
    layer0_outputs(1602) <= not (a and b);
    layer0_outputs(1603) <= not (a xor b);
    layer0_outputs(1604) <= not b or a;
    layer0_outputs(1605) <= not (a xor b);
    layer0_outputs(1606) <= not (a xor b);
    layer0_outputs(1607) <= not (a or b);
    layer0_outputs(1608) <= not a or b;
    layer0_outputs(1609) <= a xor b;
    layer0_outputs(1610) <= a and not b;
    layer0_outputs(1611) <= not a or b;
    layer0_outputs(1612) <= not b;
    layer0_outputs(1613) <= not (a or b);
    layer0_outputs(1614) <= not b or a;
    layer0_outputs(1615) <= a or b;
    layer0_outputs(1616) <= a;
    layer0_outputs(1617) <= a or b;
    layer0_outputs(1618) <= not a;
    layer0_outputs(1619) <= not b;
    layer0_outputs(1620) <= 1'b0;
    layer0_outputs(1621) <= not (a or b);
    layer0_outputs(1622) <= not a;
    layer0_outputs(1623) <= not b or a;
    layer0_outputs(1624) <= not b;
    layer0_outputs(1625) <= 1'b0;
    layer0_outputs(1626) <= not a or b;
    layer0_outputs(1627) <= not (a or b);
    layer0_outputs(1628) <= not a;
    layer0_outputs(1629) <= b;
    layer0_outputs(1630) <= b;
    layer0_outputs(1631) <= not (a or b);
    layer0_outputs(1632) <= a or b;
    layer0_outputs(1633) <= b;
    layer0_outputs(1634) <= 1'b0;
    layer0_outputs(1635) <= a xor b;
    layer0_outputs(1636) <= b;
    layer0_outputs(1637) <= not a or b;
    layer0_outputs(1638) <= a xor b;
    layer0_outputs(1639) <= a xor b;
    layer0_outputs(1640) <= a or b;
    layer0_outputs(1641) <= not a or b;
    layer0_outputs(1642) <= not b;
    layer0_outputs(1643) <= not (a and b);
    layer0_outputs(1644) <= a and b;
    layer0_outputs(1645) <= not (a or b);
    layer0_outputs(1646) <= not a;
    layer0_outputs(1647) <= not (a xor b);
    layer0_outputs(1648) <= 1'b0;
    layer0_outputs(1649) <= a xor b;
    layer0_outputs(1650) <= a;
    layer0_outputs(1651) <= not (a xor b);
    layer0_outputs(1652) <= not a or b;
    layer0_outputs(1653) <= b;
    layer0_outputs(1654) <= a and not b;
    layer0_outputs(1655) <= not b;
    layer0_outputs(1656) <= a xor b;
    layer0_outputs(1657) <= a xor b;
    layer0_outputs(1658) <= not a;
    layer0_outputs(1659) <= a xor b;
    layer0_outputs(1660) <= a and not b;
    layer0_outputs(1661) <= not b;
    layer0_outputs(1662) <= not b;
    layer0_outputs(1663) <= b;
    layer0_outputs(1664) <= a xor b;
    layer0_outputs(1665) <= a xor b;
    layer0_outputs(1666) <= a;
    layer0_outputs(1667) <= not (a xor b);
    layer0_outputs(1668) <= not b;
    layer0_outputs(1669) <= a xor b;
    layer0_outputs(1670) <= a;
    layer0_outputs(1671) <= a xor b;
    layer0_outputs(1672) <= a xor b;
    layer0_outputs(1673) <= a and not b;
    layer0_outputs(1674) <= not a or b;
    layer0_outputs(1675) <= not (a or b);
    layer0_outputs(1676) <= a or b;
    layer0_outputs(1677) <= b;
    layer0_outputs(1678) <= not (a xor b);
    layer0_outputs(1679) <= b and not a;
    layer0_outputs(1680) <= not b;
    layer0_outputs(1681) <= a xor b;
    layer0_outputs(1682) <= not (a xor b);
    layer0_outputs(1683) <= not (a xor b);
    layer0_outputs(1684) <= a and b;
    layer0_outputs(1685) <= a or b;
    layer0_outputs(1686) <= a;
    layer0_outputs(1687) <= b;
    layer0_outputs(1688) <= b;
    layer0_outputs(1689) <= not (a or b);
    layer0_outputs(1690) <= a and not b;
    layer0_outputs(1691) <= b and not a;
    layer0_outputs(1692) <= not b or a;
    layer0_outputs(1693) <= not a or b;
    layer0_outputs(1694) <= a or b;
    layer0_outputs(1695) <= not a;
    layer0_outputs(1696) <= not b;
    layer0_outputs(1697) <= not (a or b);
    layer0_outputs(1698) <= b;
    layer0_outputs(1699) <= b and not a;
    layer0_outputs(1700) <= not a;
    layer0_outputs(1701) <= not (a xor b);
    layer0_outputs(1702) <= not b or a;
    layer0_outputs(1703) <= not a;
    layer0_outputs(1704) <= a;
    layer0_outputs(1705) <= 1'b0;
    layer0_outputs(1706) <= a xor b;
    layer0_outputs(1707) <= a or b;
    layer0_outputs(1708) <= a or b;
    layer0_outputs(1709) <= not (a xor b);
    layer0_outputs(1710) <= a or b;
    layer0_outputs(1711) <= not (a xor b);
    layer0_outputs(1712) <= a xor b;
    layer0_outputs(1713) <= a or b;
    layer0_outputs(1714) <= not a or b;
    layer0_outputs(1715) <= a and b;
    layer0_outputs(1716) <= a and b;
    layer0_outputs(1717) <= not (a xor b);
    layer0_outputs(1718) <= a;
    layer0_outputs(1719) <= not a or b;
    layer0_outputs(1720) <= not (a and b);
    layer0_outputs(1721) <= not (a xor b);
    layer0_outputs(1722) <= not b or a;
    layer0_outputs(1723) <= not (a xor b);
    layer0_outputs(1724) <= a xor b;
    layer0_outputs(1725) <= a xor b;
    layer0_outputs(1726) <= not (a xor b);
    layer0_outputs(1727) <= a or b;
    layer0_outputs(1728) <= 1'b0;
    layer0_outputs(1729) <= a or b;
    layer0_outputs(1730) <= b;
    layer0_outputs(1731) <= a;
    layer0_outputs(1732) <= not (a or b);
    layer0_outputs(1733) <= not (a or b);
    layer0_outputs(1734) <= not a or b;
    layer0_outputs(1735) <= a and not b;
    layer0_outputs(1736) <= not (a xor b);
    layer0_outputs(1737) <= not (a xor b);
    layer0_outputs(1738) <= not a;
    layer0_outputs(1739) <= not (a xor b);
    layer0_outputs(1740) <= not (a xor b);
    layer0_outputs(1741) <= 1'b0;
    layer0_outputs(1742) <= not (a xor b);
    layer0_outputs(1743) <= a and not b;
    layer0_outputs(1744) <= b;
    layer0_outputs(1745) <= not (a or b);
    layer0_outputs(1746) <= not b;
    layer0_outputs(1747) <= not (a or b);
    layer0_outputs(1748) <= a and not b;
    layer0_outputs(1749) <= b and not a;
    layer0_outputs(1750) <= not a or b;
    layer0_outputs(1751) <= a or b;
    layer0_outputs(1752) <= a and not b;
    layer0_outputs(1753) <= b;
    layer0_outputs(1754) <= a;
    layer0_outputs(1755) <= a and not b;
    layer0_outputs(1756) <= a xor b;
    layer0_outputs(1757) <= a or b;
    layer0_outputs(1758) <= a and b;
    layer0_outputs(1759) <= not (a xor b);
    layer0_outputs(1760) <= not (a or b);
    layer0_outputs(1761) <= not a or b;
    layer0_outputs(1762) <= a;
    layer0_outputs(1763) <= a or b;
    layer0_outputs(1764) <= not (a or b);
    layer0_outputs(1765) <= a or b;
    layer0_outputs(1766) <= a and not b;
    layer0_outputs(1767) <= b;
    layer0_outputs(1768) <= not (a xor b);
    layer0_outputs(1769) <= not b;
    layer0_outputs(1770) <= not (a or b);
    layer0_outputs(1771) <= not (a or b);
    layer0_outputs(1772) <= a;
    layer0_outputs(1773) <= a xor b;
    layer0_outputs(1774) <= a xor b;
    layer0_outputs(1775) <= not b;
    layer0_outputs(1776) <= not b;
    layer0_outputs(1777) <= a xor b;
    layer0_outputs(1778) <= b and not a;
    layer0_outputs(1779) <= a and not b;
    layer0_outputs(1780) <= a or b;
    layer0_outputs(1781) <= not b;
    layer0_outputs(1782) <= not (a xor b);
    layer0_outputs(1783) <= a and b;
    layer0_outputs(1784) <= a and not b;
    layer0_outputs(1785) <= not (a xor b);
    layer0_outputs(1786) <= a or b;
    layer0_outputs(1787) <= not (a or b);
    layer0_outputs(1788) <= not b;
    layer0_outputs(1789) <= a or b;
    layer0_outputs(1790) <= not a;
    layer0_outputs(1791) <= a and not b;
    layer0_outputs(1792) <= a or b;
    layer0_outputs(1793) <= not (a or b);
    layer0_outputs(1794) <= 1'b1;
    layer0_outputs(1795) <= not (a xor b);
    layer0_outputs(1796) <= not (a xor b);
    layer0_outputs(1797) <= not a;
    layer0_outputs(1798) <= not (a xor b);
    layer0_outputs(1799) <= a;
    layer0_outputs(1800) <= not (a or b);
    layer0_outputs(1801) <= a xor b;
    layer0_outputs(1802) <= not (a xor b);
    layer0_outputs(1803) <= not a or b;
    layer0_outputs(1804) <= not (a xor b);
    layer0_outputs(1805) <= a or b;
    layer0_outputs(1806) <= a;
    layer0_outputs(1807) <= not b;
    layer0_outputs(1808) <= b;
    layer0_outputs(1809) <= a and not b;
    layer0_outputs(1810) <= not a;
    layer0_outputs(1811) <= not a;
    layer0_outputs(1812) <= b and not a;
    layer0_outputs(1813) <= b and not a;
    layer0_outputs(1814) <= not (a xor b);
    layer0_outputs(1815) <= a or b;
    layer0_outputs(1816) <= 1'b1;
    layer0_outputs(1817) <= 1'b1;
    layer0_outputs(1818) <= not a or b;
    layer0_outputs(1819) <= a and not b;
    layer0_outputs(1820) <= a or b;
    layer0_outputs(1821) <= a and not b;
    layer0_outputs(1822) <= not (a xor b);
    layer0_outputs(1823) <= not (a or b);
    layer0_outputs(1824) <= b and not a;
    layer0_outputs(1825) <= not b;
    layer0_outputs(1826) <= not (a xor b);
    layer0_outputs(1827) <= not (a or b);
    layer0_outputs(1828) <= not (a or b);
    layer0_outputs(1829) <= not b;
    layer0_outputs(1830) <= not a or b;
    layer0_outputs(1831) <= a and not b;
    layer0_outputs(1832) <= a or b;
    layer0_outputs(1833) <= not a or b;
    layer0_outputs(1834) <= a or b;
    layer0_outputs(1835) <= not (a or b);
    layer0_outputs(1836) <= a;
    layer0_outputs(1837) <= b and not a;
    layer0_outputs(1838) <= not (a or b);
    layer0_outputs(1839) <= b;
    layer0_outputs(1840) <= a;
    layer0_outputs(1841) <= not b;
    layer0_outputs(1842) <= a and not b;
    layer0_outputs(1843) <= not (a and b);
    layer0_outputs(1844) <= 1'b0;
    layer0_outputs(1845) <= not a or b;
    layer0_outputs(1846) <= not b;
    layer0_outputs(1847) <= a or b;
    layer0_outputs(1848) <= not b;
    layer0_outputs(1849) <= not (a or b);
    layer0_outputs(1850) <= a and not b;
    layer0_outputs(1851) <= not a or b;
    layer0_outputs(1852) <= b and not a;
    layer0_outputs(1853) <= not b;
    layer0_outputs(1854) <= a and not b;
    layer0_outputs(1855) <= not (a and b);
    layer0_outputs(1856) <= not a or b;
    layer0_outputs(1857) <= a xor b;
    layer0_outputs(1858) <= not (a xor b);
    layer0_outputs(1859) <= not b;
    layer0_outputs(1860) <= not b;
    layer0_outputs(1861) <= not b;
    layer0_outputs(1862) <= not b or a;
    layer0_outputs(1863) <= not (a or b);
    layer0_outputs(1864) <= not a;
    layer0_outputs(1865) <= a;
    layer0_outputs(1866) <= a xor b;
    layer0_outputs(1867) <= a xor b;
    layer0_outputs(1868) <= a or b;
    layer0_outputs(1869) <= not (a or b);
    layer0_outputs(1870) <= not (a or b);
    layer0_outputs(1871) <= a and not b;
    layer0_outputs(1872) <= not b;
    layer0_outputs(1873) <= not b or a;
    layer0_outputs(1874) <= a and not b;
    layer0_outputs(1875) <= a xor b;
    layer0_outputs(1876) <= b and not a;
    layer0_outputs(1877) <= a and not b;
    layer0_outputs(1878) <= a;
    layer0_outputs(1879) <= not b;
    layer0_outputs(1880) <= not (a or b);
    layer0_outputs(1881) <= not b;
    layer0_outputs(1882) <= 1'b0;
    layer0_outputs(1883) <= a or b;
    layer0_outputs(1884) <= a xor b;
    layer0_outputs(1885) <= a and not b;
    layer0_outputs(1886) <= not b or a;
    layer0_outputs(1887) <= a and not b;
    layer0_outputs(1888) <= not (a or b);
    layer0_outputs(1889) <= not a or b;
    layer0_outputs(1890) <= a and not b;
    layer0_outputs(1891) <= not (a xor b);
    layer0_outputs(1892) <= not a or b;
    layer0_outputs(1893) <= b and not a;
    layer0_outputs(1894) <= not b;
    layer0_outputs(1895) <= a xor b;
    layer0_outputs(1896) <= a and not b;
    layer0_outputs(1897) <= b;
    layer0_outputs(1898) <= not a;
    layer0_outputs(1899) <= a xor b;
    layer0_outputs(1900) <= not a;
    layer0_outputs(1901) <= a and not b;
    layer0_outputs(1902) <= not (a and b);
    layer0_outputs(1903) <= not (a xor b);
    layer0_outputs(1904) <= 1'b1;
    layer0_outputs(1905) <= a;
    layer0_outputs(1906) <= b and not a;
    layer0_outputs(1907) <= a xor b;
    layer0_outputs(1908) <= not b;
    layer0_outputs(1909) <= b and not a;
    layer0_outputs(1910) <= a or b;
    layer0_outputs(1911) <= not (a or b);
    layer0_outputs(1912) <= 1'b1;
    layer0_outputs(1913) <= a and b;
    layer0_outputs(1914) <= not b;
    layer0_outputs(1915) <= not (a or b);
    layer0_outputs(1916) <= not (a or b);
    layer0_outputs(1917) <= not (a or b);
    layer0_outputs(1918) <= not (a or b);
    layer0_outputs(1919) <= not b or a;
    layer0_outputs(1920) <= not a or b;
    layer0_outputs(1921) <= a xor b;
    layer0_outputs(1922) <= a;
    layer0_outputs(1923) <= not a;
    layer0_outputs(1924) <= a or b;
    layer0_outputs(1925) <= a or b;
    layer0_outputs(1926) <= a or b;
    layer0_outputs(1927) <= not (a or b);
    layer0_outputs(1928) <= not b or a;
    layer0_outputs(1929) <= not b;
    layer0_outputs(1930) <= not (a and b);
    layer0_outputs(1931) <= a or b;
    layer0_outputs(1932) <= not a or b;
    layer0_outputs(1933) <= a or b;
    layer0_outputs(1934) <= a or b;
    layer0_outputs(1935) <= a or b;
    layer0_outputs(1936) <= a or b;
    layer0_outputs(1937) <= not (a xor b);
    layer0_outputs(1938) <= a xor b;
    layer0_outputs(1939) <= not a or b;
    layer0_outputs(1940) <= not (a or b);
    layer0_outputs(1941) <= a and b;
    layer0_outputs(1942) <= not (a or b);
    layer0_outputs(1943) <= not a;
    layer0_outputs(1944) <= not a;
    layer0_outputs(1945) <= b;
    layer0_outputs(1946) <= not (a or b);
    layer0_outputs(1947) <= b;
    layer0_outputs(1948) <= not a;
    layer0_outputs(1949) <= a and not b;
    layer0_outputs(1950) <= b and not a;
    layer0_outputs(1951) <= b and not a;
    layer0_outputs(1952) <= not b;
    layer0_outputs(1953) <= not a;
    layer0_outputs(1954) <= a xor b;
    layer0_outputs(1955) <= a and not b;
    layer0_outputs(1956) <= not b or a;
    layer0_outputs(1957) <= not (a xor b);
    layer0_outputs(1958) <= not (a or b);
    layer0_outputs(1959) <= a and not b;
    layer0_outputs(1960) <= a;
    layer0_outputs(1961) <= a and b;
    layer0_outputs(1962) <= b and not a;
    layer0_outputs(1963) <= b;
    layer0_outputs(1964) <= not a or b;
    layer0_outputs(1965) <= not b;
    layer0_outputs(1966) <= a;
    layer0_outputs(1967) <= not (a xor b);
    layer0_outputs(1968) <= a or b;
    layer0_outputs(1969) <= b;
    layer0_outputs(1970) <= a;
    layer0_outputs(1971) <= a and not b;
    layer0_outputs(1972) <= not a;
    layer0_outputs(1973) <= 1'b1;
    layer0_outputs(1974) <= 1'b0;
    layer0_outputs(1975) <= a xor b;
    layer0_outputs(1976) <= b and not a;
    layer0_outputs(1977) <= a or b;
    layer0_outputs(1978) <= not a;
    layer0_outputs(1979) <= b;
    layer0_outputs(1980) <= a and not b;
    layer0_outputs(1981) <= a xor b;
    layer0_outputs(1982) <= b and not a;
    layer0_outputs(1983) <= not a;
    layer0_outputs(1984) <= a and not b;
    layer0_outputs(1985) <= not b or a;
    layer0_outputs(1986) <= not (a or b);
    layer0_outputs(1987) <= not b;
    layer0_outputs(1988) <= a xor b;
    layer0_outputs(1989) <= 1'b0;
    layer0_outputs(1990) <= b and not a;
    layer0_outputs(1991) <= not a or b;
    layer0_outputs(1992) <= not (a or b);
    layer0_outputs(1993) <= not b or a;
    layer0_outputs(1994) <= not a or b;
    layer0_outputs(1995) <= not (a or b);
    layer0_outputs(1996) <= not (a or b);
    layer0_outputs(1997) <= a or b;
    layer0_outputs(1998) <= not b;
    layer0_outputs(1999) <= a or b;
    layer0_outputs(2000) <= b;
    layer0_outputs(2001) <= not a or b;
    layer0_outputs(2002) <= a xor b;
    layer0_outputs(2003) <= not a;
    layer0_outputs(2004) <= a and not b;
    layer0_outputs(2005) <= a;
    layer0_outputs(2006) <= a or b;
    layer0_outputs(2007) <= 1'b1;
    layer0_outputs(2008) <= a xor b;
    layer0_outputs(2009) <= a or b;
    layer0_outputs(2010) <= not a or b;
    layer0_outputs(2011) <= not b;
    layer0_outputs(2012) <= not b or a;
    layer0_outputs(2013) <= not (a or b);
    layer0_outputs(2014) <= a xor b;
    layer0_outputs(2015) <= not b;
    layer0_outputs(2016) <= not (a xor b);
    layer0_outputs(2017) <= not (a xor b);
    layer0_outputs(2018) <= a and b;
    layer0_outputs(2019) <= not a or b;
    layer0_outputs(2020) <= not (a or b);
    layer0_outputs(2021) <= a or b;
    layer0_outputs(2022) <= not a;
    layer0_outputs(2023) <= not a;
    layer0_outputs(2024) <= a or b;
    layer0_outputs(2025) <= 1'b1;
    layer0_outputs(2026) <= not (a or b);
    layer0_outputs(2027) <= a and not b;
    layer0_outputs(2028) <= not a or b;
    layer0_outputs(2029) <= a xor b;
    layer0_outputs(2030) <= not (a xor b);
    layer0_outputs(2031) <= not a;
    layer0_outputs(2032) <= a;
    layer0_outputs(2033) <= a and not b;
    layer0_outputs(2034) <= a xor b;
    layer0_outputs(2035) <= not (a or b);
    layer0_outputs(2036) <= a xor b;
    layer0_outputs(2037) <= a xor b;
    layer0_outputs(2038) <= not b or a;
    layer0_outputs(2039) <= 1'b0;
    layer0_outputs(2040) <= not (a or b);
    layer0_outputs(2041) <= not a;
    layer0_outputs(2042) <= b;
    layer0_outputs(2043) <= a;
    layer0_outputs(2044) <= not (a and b);
    layer0_outputs(2045) <= 1'b1;
    layer0_outputs(2046) <= not (a or b);
    layer0_outputs(2047) <= a and not b;
    layer0_outputs(2048) <= a or b;
    layer0_outputs(2049) <= not a or b;
    layer0_outputs(2050) <= not b;
    layer0_outputs(2051) <= b and not a;
    layer0_outputs(2052) <= not (a or b);
    layer0_outputs(2053) <= b and not a;
    layer0_outputs(2054) <= not (a or b);
    layer0_outputs(2055) <= 1'b0;
    layer0_outputs(2056) <= not b;
    layer0_outputs(2057) <= not b or a;
    layer0_outputs(2058) <= not (a or b);
    layer0_outputs(2059) <= a and not b;
    layer0_outputs(2060) <= not b or a;
    layer0_outputs(2061) <= not (a xor b);
    layer0_outputs(2062) <= a;
    layer0_outputs(2063) <= a or b;
    layer0_outputs(2064) <= a or b;
    layer0_outputs(2065) <= a xor b;
    layer0_outputs(2066) <= not a;
    layer0_outputs(2067) <= a;
    layer0_outputs(2068) <= not (a or b);
    layer0_outputs(2069) <= not (a or b);
    layer0_outputs(2070) <= b and not a;
    layer0_outputs(2071) <= not (a xor b);
    layer0_outputs(2072) <= not a;
    layer0_outputs(2073) <= 1'b1;
    layer0_outputs(2074) <= a or b;
    layer0_outputs(2075) <= not a or b;
    layer0_outputs(2076) <= not b or a;
    layer0_outputs(2077) <= a or b;
    layer0_outputs(2078) <= a xor b;
    layer0_outputs(2079) <= a or b;
    layer0_outputs(2080) <= a;
    layer0_outputs(2081) <= not b;
    layer0_outputs(2082) <= not a or b;
    layer0_outputs(2083) <= a xor b;
    layer0_outputs(2084) <= not a;
    layer0_outputs(2085) <= a xor b;
    layer0_outputs(2086) <= b and not a;
    layer0_outputs(2087) <= b and not a;
    layer0_outputs(2088) <= not a or b;
    layer0_outputs(2089) <= a xor b;
    layer0_outputs(2090) <= a or b;
    layer0_outputs(2091) <= not (a xor b);
    layer0_outputs(2092) <= not (a or b);
    layer0_outputs(2093) <= a xor b;
    layer0_outputs(2094) <= not (a or b);
    layer0_outputs(2095) <= a or b;
    layer0_outputs(2096) <= b and not a;
    layer0_outputs(2097) <= 1'b1;
    layer0_outputs(2098) <= b and not a;
    layer0_outputs(2099) <= not (a and b);
    layer0_outputs(2100) <= 1'b0;
    layer0_outputs(2101) <= not b or a;
    layer0_outputs(2102) <= 1'b0;
    layer0_outputs(2103) <= not (a or b);
    layer0_outputs(2104) <= a xor b;
    layer0_outputs(2105) <= not b;
    layer0_outputs(2106) <= not (a or b);
    layer0_outputs(2107) <= a or b;
    layer0_outputs(2108) <= not b or a;
    layer0_outputs(2109) <= b;
    layer0_outputs(2110) <= b;
    layer0_outputs(2111) <= not a or b;
    layer0_outputs(2112) <= not (a xor b);
    layer0_outputs(2113) <= not b or a;
    layer0_outputs(2114) <= a xor b;
    layer0_outputs(2115) <= a xor b;
    layer0_outputs(2116) <= a xor b;
    layer0_outputs(2117) <= a or b;
    layer0_outputs(2118) <= a xor b;
    layer0_outputs(2119) <= a xor b;
    layer0_outputs(2120) <= a xor b;
    layer0_outputs(2121) <= a or b;
    layer0_outputs(2122) <= not b;
    layer0_outputs(2123) <= not (a xor b);
    layer0_outputs(2124) <= b;
    layer0_outputs(2125) <= not (a xor b);
    layer0_outputs(2126) <= b and not a;
    layer0_outputs(2127) <= not b or a;
    layer0_outputs(2128) <= b;
    layer0_outputs(2129) <= a xor b;
    layer0_outputs(2130) <= a or b;
    layer0_outputs(2131) <= not b;
    layer0_outputs(2132) <= a xor b;
    layer0_outputs(2133) <= a or b;
    layer0_outputs(2134) <= not b;
    layer0_outputs(2135) <= not b or a;
    layer0_outputs(2136) <= a xor b;
    layer0_outputs(2137) <= a and not b;
    layer0_outputs(2138) <= a xor b;
    layer0_outputs(2139) <= not a or b;
    layer0_outputs(2140) <= not a or b;
    layer0_outputs(2141) <= b;
    layer0_outputs(2142) <= not (a or b);
    layer0_outputs(2143) <= not b;
    layer0_outputs(2144) <= not (a xor b);
    layer0_outputs(2145) <= a and b;
    layer0_outputs(2146) <= b and not a;
    layer0_outputs(2147) <= not (a xor b);
    layer0_outputs(2148) <= not (a or b);
    layer0_outputs(2149) <= not b or a;
    layer0_outputs(2150) <= a or b;
    layer0_outputs(2151) <= not (a xor b);
    layer0_outputs(2152) <= not (a xor b);
    layer0_outputs(2153) <= a;
    layer0_outputs(2154) <= not b;
    layer0_outputs(2155) <= a;
    layer0_outputs(2156) <= a or b;
    layer0_outputs(2157) <= a;
    layer0_outputs(2158) <= not b;
    layer0_outputs(2159) <= b and not a;
    layer0_outputs(2160) <= not (a or b);
    layer0_outputs(2161) <= not b;
    layer0_outputs(2162) <= not (a and b);
    layer0_outputs(2163) <= not (a and b);
    layer0_outputs(2164) <= not a;
    layer0_outputs(2165) <= a xor b;
    layer0_outputs(2166) <= a and not b;
    layer0_outputs(2167) <= a xor b;
    layer0_outputs(2168) <= a or b;
    layer0_outputs(2169) <= not (a and b);
    layer0_outputs(2170) <= not (a or b);
    layer0_outputs(2171) <= not a;
    layer0_outputs(2172) <= not (a or b);
    layer0_outputs(2173) <= not a;
    layer0_outputs(2174) <= a or b;
    layer0_outputs(2175) <= not (a and b);
    layer0_outputs(2176) <= not (a or b);
    layer0_outputs(2177) <= 1'b0;
    layer0_outputs(2178) <= not (a xor b);
    layer0_outputs(2179) <= not a;
    layer0_outputs(2180) <= not a;
    layer0_outputs(2181) <= a or b;
    layer0_outputs(2182) <= not a;
    layer0_outputs(2183) <= not (a and b);
    layer0_outputs(2184) <= a;
    layer0_outputs(2185) <= a or b;
    layer0_outputs(2186) <= 1'b0;
    layer0_outputs(2187) <= not (a xor b);
    layer0_outputs(2188) <= not a or b;
    layer0_outputs(2189) <= b;
    layer0_outputs(2190) <= a and not b;
    layer0_outputs(2191) <= b and not a;
    layer0_outputs(2192) <= not (a xor b);
    layer0_outputs(2193) <= a or b;
    layer0_outputs(2194) <= a and not b;
    layer0_outputs(2195) <= not (a or b);
    layer0_outputs(2196) <= not b;
    layer0_outputs(2197) <= not (a or b);
    layer0_outputs(2198) <= not b;
    layer0_outputs(2199) <= a or b;
    layer0_outputs(2200) <= b and not a;
    layer0_outputs(2201) <= not (a or b);
    layer0_outputs(2202) <= b and not a;
    layer0_outputs(2203) <= not (a xor b);
    layer0_outputs(2204) <= a and b;
    layer0_outputs(2205) <= not (a or b);
    layer0_outputs(2206) <= not (a or b);
    layer0_outputs(2207) <= a xor b;
    layer0_outputs(2208) <= not a;
    layer0_outputs(2209) <= b;
    layer0_outputs(2210) <= not (a xor b);
    layer0_outputs(2211) <= not (a or b);
    layer0_outputs(2212) <= a;
    layer0_outputs(2213) <= not (a and b);
    layer0_outputs(2214) <= not a;
    layer0_outputs(2215) <= not b or a;
    layer0_outputs(2216) <= not (a xor b);
    layer0_outputs(2217) <= a and not b;
    layer0_outputs(2218) <= a or b;
    layer0_outputs(2219) <= not (a or b);
    layer0_outputs(2220) <= not (a or b);
    layer0_outputs(2221) <= a;
    layer0_outputs(2222) <= a and not b;
    layer0_outputs(2223) <= a and not b;
    layer0_outputs(2224) <= b;
    layer0_outputs(2225) <= not (a xor b);
    layer0_outputs(2226) <= a or b;
    layer0_outputs(2227) <= b and not a;
    layer0_outputs(2228) <= a;
    layer0_outputs(2229) <= not (a or b);
    layer0_outputs(2230) <= a xor b;
    layer0_outputs(2231) <= a xor b;
    layer0_outputs(2232) <= a or b;
    layer0_outputs(2233) <= not b;
    layer0_outputs(2234) <= a xor b;
    layer0_outputs(2235) <= a and not b;
    layer0_outputs(2236) <= b and not a;
    layer0_outputs(2237) <= not a or b;
    layer0_outputs(2238) <= not (a or b);
    layer0_outputs(2239) <= 1'b0;
    layer0_outputs(2240) <= not (a xor b);
    layer0_outputs(2241) <= not a;
    layer0_outputs(2242) <= b and not a;
    layer0_outputs(2243) <= a xor b;
    layer0_outputs(2244) <= not (a or b);
    layer0_outputs(2245) <= a or b;
    layer0_outputs(2246) <= not b or a;
    layer0_outputs(2247) <= not a;
    layer0_outputs(2248) <= not b or a;
    layer0_outputs(2249) <= not b or a;
    layer0_outputs(2250) <= not (a xor b);
    layer0_outputs(2251) <= a and b;
    layer0_outputs(2252) <= not (a xor b);
    layer0_outputs(2253) <= not (a or b);
    layer0_outputs(2254) <= a xor b;
    layer0_outputs(2255) <= a or b;
    layer0_outputs(2256) <= not a;
    layer0_outputs(2257) <= a xor b;
    layer0_outputs(2258) <= not a or b;
    layer0_outputs(2259) <= b;
    layer0_outputs(2260) <= 1'b0;
    layer0_outputs(2261) <= a xor b;
    layer0_outputs(2262) <= not a or b;
    layer0_outputs(2263) <= a xor b;
    layer0_outputs(2264) <= a and b;
    layer0_outputs(2265) <= not (a and b);
    layer0_outputs(2266) <= 1'b0;
    layer0_outputs(2267) <= not b or a;
    layer0_outputs(2268) <= a or b;
    layer0_outputs(2269) <= a and b;
    layer0_outputs(2270) <= b and not a;
    layer0_outputs(2271) <= 1'b0;
    layer0_outputs(2272) <= not b;
    layer0_outputs(2273) <= a xor b;
    layer0_outputs(2274) <= not (a xor b);
    layer0_outputs(2275) <= a xor b;
    layer0_outputs(2276) <= not (a xor b);
    layer0_outputs(2277) <= a or b;
    layer0_outputs(2278) <= a or b;
    layer0_outputs(2279) <= a or b;
    layer0_outputs(2280) <= b;
    layer0_outputs(2281) <= not a;
    layer0_outputs(2282) <= not (a xor b);
    layer0_outputs(2283) <= b and not a;
    layer0_outputs(2284) <= not a or b;
    layer0_outputs(2285) <= not a or b;
    layer0_outputs(2286) <= not (a or b);
    layer0_outputs(2287) <= not a or b;
    layer0_outputs(2288) <= a and not b;
    layer0_outputs(2289) <= not a or b;
    layer0_outputs(2290) <= b;
    layer0_outputs(2291) <= b;
    layer0_outputs(2292) <= a and not b;
    layer0_outputs(2293) <= not (a or b);
    layer0_outputs(2294) <= not b;
    layer0_outputs(2295) <= not a or b;
    layer0_outputs(2296) <= b and not a;
    layer0_outputs(2297) <= a and not b;
    layer0_outputs(2298) <= a or b;
    layer0_outputs(2299) <= not (a xor b);
    layer0_outputs(2300) <= not (a or b);
    layer0_outputs(2301) <= a;
    layer0_outputs(2302) <= not a or b;
    layer0_outputs(2303) <= a and b;
    layer0_outputs(2304) <= not (a and b);
    layer0_outputs(2305) <= not b or a;
    layer0_outputs(2306) <= not a;
    layer0_outputs(2307) <= b;
    layer0_outputs(2308) <= not a;
    layer0_outputs(2309) <= a and b;
    layer0_outputs(2310) <= not (a or b);
    layer0_outputs(2311) <= a or b;
    layer0_outputs(2312) <= not a or b;
    layer0_outputs(2313) <= a;
    layer0_outputs(2314) <= not (a or b);
    layer0_outputs(2315) <= not b or a;
    layer0_outputs(2316) <= not (a or b);
    layer0_outputs(2317) <= not b or a;
    layer0_outputs(2318) <= not (a or b);
    layer0_outputs(2319) <= 1'b1;
    layer0_outputs(2320) <= not (a xor b);
    layer0_outputs(2321) <= a and b;
    layer0_outputs(2322) <= not b or a;
    layer0_outputs(2323) <= b;
    layer0_outputs(2324) <= not a or b;
    layer0_outputs(2325) <= a or b;
    layer0_outputs(2326) <= a;
    layer0_outputs(2327) <= a;
    layer0_outputs(2328) <= not b;
    layer0_outputs(2329) <= not (a xor b);
    layer0_outputs(2330) <= not a or b;
    layer0_outputs(2331) <= a or b;
    layer0_outputs(2332) <= not (a or b);
    layer0_outputs(2333) <= a and not b;
    layer0_outputs(2334) <= not a or b;
    layer0_outputs(2335) <= not b;
    layer0_outputs(2336) <= not b;
    layer0_outputs(2337) <= not (a or b);
    layer0_outputs(2338) <= not (a or b);
    layer0_outputs(2339) <= not (a or b);
    layer0_outputs(2340) <= a or b;
    layer0_outputs(2341) <= a and not b;
    layer0_outputs(2342) <= not (a xor b);
    layer0_outputs(2343) <= a xor b;
    layer0_outputs(2344) <= a or b;
    layer0_outputs(2345) <= a or b;
    layer0_outputs(2346) <= a xor b;
    layer0_outputs(2347) <= a and not b;
    layer0_outputs(2348) <= a;
    layer0_outputs(2349) <= not (a or b);
    layer0_outputs(2350) <= not a or b;
    layer0_outputs(2351) <= a xor b;
    layer0_outputs(2352) <= not (a and b);
    layer0_outputs(2353) <= a and not b;
    layer0_outputs(2354) <= not a or b;
    layer0_outputs(2355) <= b and not a;
    layer0_outputs(2356) <= not a or b;
    layer0_outputs(2357) <= not a or b;
    layer0_outputs(2358) <= not (a xor b);
    layer0_outputs(2359) <= b and not a;
    layer0_outputs(2360) <= not b;
    layer0_outputs(2361) <= b;
    layer0_outputs(2362) <= not (a or b);
    layer0_outputs(2363) <= not a or b;
    layer0_outputs(2364) <= not b or a;
    layer0_outputs(2365) <= a or b;
    layer0_outputs(2366) <= not (a xor b);
    layer0_outputs(2367) <= b;
    layer0_outputs(2368) <= not (a or b);
    layer0_outputs(2369) <= a xor b;
    layer0_outputs(2370) <= a or b;
    layer0_outputs(2371) <= not b;
    layer0_outputs(2372) <= not b;
    layer0_outputs(2373) <= not b;
    layer0_outputs(2374) <= a xor b;
    layer0_outputs(2375) <= not (a or b);
    layer0_outputs(2376) <= a or b;
    layer0_outputs(2377) <= 1'b0;
    layer0_outputs(2378) <= b;
    layer0_outputs(2379) <= a;
    layer0_outputs(2380) <= b and not a;
    layer0_outputs(2381) <= 1'b0;
    layer0_outputs(2382) <= a or b;
    layer0_outputs(2383) <= not (a xor b);
    layer0_outputs(2384) <= not a or b;
    layer0_outputs(2385) <= a;
    layer0_outputs(2386) <= b and not a;
    layer0_outputs(2387) <= 1'b0;
    layer0_outputs(2388) <= not (a or b);
    layer0_outputs(2389) <= not b or a;
    layer0_outputs(2390) <= not (a xor b);
    layer0_outputs(2391) <= a;
    layer0_outputs(2392) <= a and not b;
    layer0_outputs(2393) <= not a;
    layer0_outputs(2394) <= not (a xor b);
    layer0_outputs(2395) <= a and not b;
    layer0_outputs(2396) <= not a or b;
    layer0_outputs(2397) <= not (a or b);
    layer0_outputs(2398) <= not (a xor b);
    layer0_outputs(2399) <= 1'b1;
    layer0_outputs(2400) <= not b or a;
    layer0_outputs(2401) <= a or b;
    layer0_outputs(2402) <= a and not b;
    layer0_outputs(2403) <= b;
    layer0_outputs(2404) <= b and not a;
    layer0_outputs(2405) <= a xor b;
    layer0_outputs(2406) <= not a;
    layer0_outputs(2407) <= a or b;
    layer0_outputs(2408) <= a and not b;
    layer0_outputs(2409) <= not a or b;
    layer0_outputs(2410) <= not a;
    layer0_outputs(2411) <= b and not a;
    layer0_outputs(2412) <= a;
    layer0_outputs(2413) <= not (a or b);
    layer0_outputs(2414) <= a and not b;
    layer0_outputs(2415) <= a;
    layer0_outputs(2416) <= b and not a;
    layer0_outputs(2417) <= a or b;
    layer0_outputs(2418) <= not (a xor b);
    layer0_outputs(2419) <= not a or b;
    layer0_outputs(2420) <= not a or b;
    layer0_outputs(2421) <= not b or a;
    layer0_outputs(2422) <= not (a xor b);
    layer0_outputs(2423) <= not (a and b);
    layer0_outputs(2424) <= a or b;
    layer0_outputs(2425) <= a;
    layer0_outputs(2426) <= a xor b;
    layer0_outputs(2427) <= not b or a;
    layer0_outputs(2428) <= a or b;
    layer0_outputs(2429) <= a;
    layer0_outputs(2430) <= not (a xor b);
    layer0_outputs(2431) <= a;
    layer0_outputs(2432) <= not (a or b);
    layer0_outputs(2433) <= not (a xor b);
    layer0_outputs(2434) <= b;
    layer0_outputs(2435) <= a xor b;
    layer0_outputs(2436) <= a xor b;
    layer0_outputs(2437) <= a xor b;
    layer0_outputs(2438) <= not (a or b);
    layer0_outputs(2439) <= a or b;
    layer0_outputs(2440) <= a xor b;
    layer0_outputs(2441) <= a xor b;
    layer0_outputs(2442) <= b;
    layer0_outputs(2443) <= a and b;
    layer0_outputs(2444) <= not a or b;
    layer0_outputs(2445) <= a and not b;
    layer0_outputs(2446) <= b;
    layer0_outputs(2447) <= not (a xor b);
    layer0_outputs(2448) <= a or b;
    layer0_outputs(2449) <= a xor b;
    layer0_outputs(2450) <= a;
    layer0_outputs(2451) <= a and not b;
    layer0_outputs(2452) <= a and b;
    layer0_outputs(2453) <= not (a xor b);
    layer0_outputs(2454) <= not (a or b);
    layer0_outputs(2455) <= not a or b;
    layer0_outputs(2456) <= 1'b1;
    layer0_outputs(2457) <= a or b;
    layer0_outputs(2458) <= not a;
    layer0_outputs(2459) <= a or b;
    layer0_outputs(2460) <= a xor b;
    layer0_outputs(2461) <= b and not a;
    layer0_outputs(2462) <= not b or a;
    layer0_outputs(2463) <= a and not b;
    layer0_outputs(2464) <= not (a xor b);
    layer0_outputs(2465) <= not b;
    layer0_outputs(2466) <= a and not b;
    layer0_outputs(2467) <= a xor b;
    layer0_outputs(2468) <= not (a xor b);
    layer0_outputs(2469) <= not (a xor b);
    layer0_outputs(2470) <= b;
    layer0_outputs(2471) <= not (a xor b);
    layer0_outputs(2472) <= not (a or b);
    layer0_outputs(2473) <= not (a xor b);
    layer0_outputs(2474) <= a or b;
    layer0_outputs(2475) <= not (a or b);
    layer0_outputs(2476) <= b and not a;
    layer0_outputs(2477) <= a xor b;
    layer0_outputs(2478) <= a;
    layer0_outputs(2479) <= b and not a;
    layer0_outputs(2480) <= not b;
    layer0_outputs(2481) <= not (a or b);
    layer0_outputs(2482) <= not (a xor b);
    layer0_outputs(2483) <= not b;
    layer0_outputs(2484) <= not a or b;
    layer0_outputs(2485) <= a and not b;
    layer0_outputs(2486) <= a xor b;
    layer0_outputs(2487) <= not b;
    layer0_outputs(2488) <= b and not a;
    layer0_outputs(2489) <= not (a and b);
    layer0_outputs(2490) <= a;
    layer0_outputs(2491) <= a and not b;
    layer0_outputs(2492) <= not b or a;
    layer0_outputs(2493) <= 1'b0;
    layer0_outputs(2494) <= a xor b;
    layer0_outputs(2495) <= b and not a;
    layer0_outputs(2496) <= not b;
    layer0_outputs(2497) <= a xor b;
    layer0_outputs(2498) <= a or b;
    layer0_outputs(2499) <= 1'b1;
    layer0_outputs(2500) <= b;
    layer0_outputs(2501) <= a and not b;
    layer0_outputs(2502) <= a and not b;
    layer0_outputs(2503) <= not a or b;
    layer0_outputs(2504) <= a xor b;
    layer0_outputs(2505) <= b;
    layer0_outputs(2506) <= not b or a;
    layer0_outputs(2507) <= not (a or b);
    layer0_outputs(2508) <= not a;
    layer0_outputs(2509) <= b and not a;
    layer0_outputs(2510) <= not (a or b);
    layer0_outputs(2511) <= not a;
    layer0_outputs(2512) <= a or b;
    layer0_outputs(2513) <= not (a or b);
    layer0_outputs(2514) <= b and not a;
    layer0_outputs(2515) <= not b or a;
    layer0_outputs(2516) <= 1'b0;
    layer0_outputs(2517) <= 1'b0;
    layer0_outputs(2518) <= not b or a;
    layer0_outputs(2519) <= not (a xor b);
    layer0_outputs(2520) <= not (a xor b);
    layer0_outputs(2521) <= a xor b;
    layer0_outputs(2522) <= b and not a;
    layer0_outputs(2523) <= b and not a;
    layer0_outputs(2524) <= a and not b;
    layer0_outputs(2525) <= a and not b;
    layer0_outputs(2526) <= not (a or b);
    layer0_outputs(2527) <= b and not a;
    layer0_outputs(2528) <= b and not a;
    layer0_outputs(2529) <= a or b;
    layer0_outputs(2530) <= a;
    layer0_outputs(2531) <= a xor b;
    layer0_outputs(2532) <= not b or a;
    layer0_outputs(2533) <= not (a xor b);
    layer0_outputs(2534) <= a;
    layer0_outputs(2535) <= not (a xor b);
    layer0_outputs(2536) <= a xor b;
    layer0_outputs(2537) <= a xor b;
    layer0_outputs(2538) <= a or b;
    layer0_outputs(2539) <= not a;
    layer0_outputs(2540) <= not b;
    layer0_outputs(2541) <= a and b;
    layer0_outputs(2542) <= not a;
    layer0_outputs(2543) <= not a;
    layer0_outputs(2544) <= a or b;
    layer0_outputs(2545) <= a xor b;
    layer0_outputs(2546) <= not (a xor b);
    layer0_outputs(2547) <= not b;
    layer0_outputs(2548) <= a and not b;
    layer0_outputs(2549) <= a or b;
    layer0_outputs(2550) <= a and not b;
    layer0_outputs(2551) <= not (a or b);
    layer0_outputs(2552) <= not a or b;
    layer0_outputs(2553) <= not (a xor b);
    layer0_outputs(2554) <= b and not a;
    layer0_outputs(2555) <= a or b;
    layer0_outputs(2556) <= not a or b;
    layer0_outputs(2557) <= a and not b;
    layer0_outputs(2558) <= a and b;
    layer0_outputs(2559) <= not (a or b);
    layer0_outputs(2560) <= b;
    layer0_outputs(2561) <= not (a and b);
    layer0_outputs(2562) <= a or b;
    layer0_outputs(2563) <= a or b;
    layer0_outputs(2564) <= not (a or b);
    layer0_outputs(2565) <= not (a or b);
    layer0_outputs(2566) <= b;
    layer0_outputs(2567) <= not (a xor b);
    layer0_outputs(2568) <= not (a xor b);
    layer0_outputs(2569) <= not (a xor b);
    layer0_outputs(2570) <= a and not b;
    layer0_outputs(2571) <= b and not a;
    layer0_outputs(2572) <= not a;
    layer0_outputs(2573) <= not a;
    layer0_outputs(2574) <= a or b;
    layer0_outputs(2575) <= not (a or b);
    layer0_outputs(2576) <= not b;
    layer0_outputs(2577) <= a xor b;
    layer0_outputs(2578) <= not a;
    layer0_outputs(2579) <= a;
    layer0_outputs(2580) <= not a or b;
    layer0_outputs(2581) <= not b or a;
    layer0_outputs(2582) <= a and not b;
    layer0_outputs(2583) <= not (a or b);
    layer0_outputs(2584) <= not a;
    layer0_outputs(2585) <= not (a xor b);
    layer0_outputs(2586) <= not b or a;
    layer0_outputs(2587) <= a and b;
    layer0_outputs(2588) <= a xor b;
    layer0_outputs(2589) <= not a or b;
    layer0_outputs(2590) <= a or b;
    layer0_outputs(2591) <= a or b;
    layer0_outputs(2592) <= a or b;
    layer0_outputs(2593) <= b;
    layer0_outputs(2594) <= not a;
    layer0_outputs(2595) <= a and not b;
    layer0_outputs(2596) <= a;
    layer0_outputs(2597) <= 1'b1;
    layer0_outputs(2598) <= b and not a;
    layer0_outputs(2599) <= a xor b;
    layer0_outputs(2600) <= b and not a;
    layer0_outputs(2601) <= a xor b;
    layer0_outputs(2602) <= not (a or b);
    layer0_outputs(2603) <= b and not a;
    layer0_outputs(2604) <= b and not a;
    layer0_outputs(2605) <= 1'b1;
    layer0_outputs(2606) <= a xor b;
    layer0_outputs(2607) <= a or b;
    layer0_outputs(2608) <= b and not a;
    layer0_outputs(2609) <= not (a or b);
    layer0_outputs(2610) <= a xor b;
    layer0_outputs(2611) <= a or b;
    layer0_outputs(2612) <= a or b;
    layer0_outputs(2613) <= a or b;
    layer0_outputs(2614) <= not b or a;
    layer0_outputs(2615) <= not (a or b);
    layer0_outputs(2616) <= 1'b1;
    layer0_outputs(2617) <= b and not a;
    layer0_outputs(2618) <= a or b;
    layer0_outputs(2619) <= not a;
    layer0_outputs(2620) <= not a or b;
    layer0_outputs(2621) <= a xor b;
    layer0_outputs(2622) <= not b or a;
    layer0_outputs(2623) <= not b;
    layer0_outputs(2624) <= a or b;
    layer0_outputs(2625) <= not (a or b);
    layer0_outputs(2626) <= a xor b;
    layer0_outputs(2627) <= a and not b;
    layer0_outputs(2628) <= 1'b0;
    layer0_outputs(2629) <= not (a and b);
    layer0_outputs(2630) <= not a;
    layer0_outputs(2631) <= not a or b;
    layer0_outputs(2632) <= b;
    layer0_outputs(2633) <= not (a xor b);
    layer0_outputs(2634) <= a xor b;
    layer0_outputs(2635) <= a and b;
    layer0_outputs(2636) <= b and not a;
    layer0_outputs(2637) <= a or b;
    layer0_outputs(2638) <= a;
    layer0_outputs(2639) <= not (a and b);
    layer0_outputs(2640) <= not (a xor b);
    layer0_outputs(2641) <= not b;
    layer0_outputs(2642) <= not (a or b);
    layer0_outputs(2643) <= not (a xor b);
    layer0_outputs(2644) <= not a or b;
    layer0_outputs(2645) <= not (a or b);
    layer0_outputs(2646) <= not (a xor b);
    layer0_outputs(2647) <= a and not b;
    layer0_outputs(2648) <= b and not a;
    layer0_outputs(2649) <= b;
    layer0_outputs(2650) <= a;
    layer0_outputs(2651) <= a xor b;
    layer0_outputs(2652) <= a or b;
    layer0_outputs(2653) <= not b or a;
    layer0_outputs(2654) <= b and not a;
    layer0_outputs(2655) <= b;
    layer0_outputs(2656) <= not (a and b);
    layer0_outputs(2657) <= not a or b;
    layer0_outputs(2658) <= a and not b;
    layer0_outputs(2659) <= not (a or b);
    layer0_outputs(2660) <= a;
    layer0_outputs(2661) <= a xor b;
    layer0_outputs(2662) <= not (a xor b);
    layer0_outputs(2663) <= not a;
    layer0_outputs(2664) <= not b or a;
    layer0_outputs(2665) <= a xor b;
    layer0_outputs(2666) <= b and not a;
    layer0_outputs(2667) <= not (a or b);
    layer0_outputs(2668) <= a xor b;
    layer0_outputs(2669) <= not b or a;
    layer0_outputs(2670) <= not a or b;
    layer0_outputs(2671) <= not b or a;
    layer0_outputs(2672) <= a xor b;
    layer0_outputs(2673) <= not (a or b);
    layer0_outputs(2674) <= a xor b;
    layer0_outputs(2675) <= not b or a;
    layer0_outputs(2676) <= a and not b;
    layer0_outputs(2677) <= a or b;
    layer0_outputs(2678) <= a or b;
    layer0_outputs(2679) <= not a or b;
    layer0_outputs(2680) <= not (a and b);
    layer0_outputs(2681) <= b;
    layer0_outputs(2682) <= not (a or b);
    layer0_outputs(2683) <= a xor b;
    layer0_outputs(2684) <= not (a and b);
    layer0_outputs(2685) <= a and b;
    layer0_outputs(2686) <= not a;
    layer0_outputs(2687) <= a or b;
    layer0_outputs(2688) <= not (a xor b);
    layer0_outputs(2689) <= not a;
    layer0_outputs(2690) <= a and b;
    layer0_outputs(2691) <= a xor b;
    layer0_outputs(2692) <= not (a xor b);
    layer0_outputs(2693) <= not (a or b);
    layer0_outputs(2694) <= a or b;
    layer0_outputs(2695) <= not (a xor b);
    layer0_outputs(2696) <= a;
    layer0_outputs(2697) <= a;
    layer0_outputs(2698) <= not b;
    layer0_outputs(2699) <= not a;
    layer0_outputs(2700) <= not (a or b);
    layer0_outputs(2701) <= not (a xor b);
    layer0_outputs(2702) <= a and not b;
    layer0_outputs(2703) <= not a or b;
    layer0_outputs(2704) <= b;
    layer0_outputs(2705) <= a and not b;
    layer0_outputs(2706) <= a and b;
    layer0_outputs(2707) <= a and not b;
    layer0_outputs(2708) <= b and not a;
    layer0_outputs(2709) <= not b or a;
    layer0_outputs(2710) <= 1'b0;
    layer0_outputs(2711) <= a or b;
    layer0_outputs(2712) <= a xor b;
    layer0_outputs(2713) <= not (a or b);
    layer0_outputs(2714) <= not (a xor b);
    layer0_outputs(2715) <= b and not a;
    layer0_outputs(2716) <= not b or a;
    layer0_outputs(2717) <= not a;
    layer0_outputs(2718) <= a xor b;
    layer0_outputs(2719) <= not b;
    layer0_outputs(2720) <= b;
    layer0_outputs(2721) <= b;
    layer0_outputs(2722) <= not (a or b);
    layer0_outputs(2723) <= a;
    layer0_outputs(2724) <= a xor b;
    layer0_outputs(2725) <= b;
    layer0_outputs(2726) <= a and not b;
    layer0_outputs(2727) <= a and not b;
    layer0_outputs(2728) <= b;
    layer0_outputs(2729) <= not (a xor b);
    layer0_outputs(2730) <= b and not a;
    layer0_outputs(2731) <= not (a and b);
    layer0_outputs(2732) <= not (a or b);
    layer0_outputs(2733) <= 1'b0;
    layer0_outputs(2734) <= a;
    layer0_outputs(2735) <= a and not b;
    layer0_outputs(2736) <= not a or b;
    layer0_outputs(2737) <= not (a xor b);
    layer0_outputs(2738) <= a xor b;
    layer0_outputs(2739) <= not a;
    layer0_outputs(2740) <= a xor b;
    layer0_outputs(2741) <= not (a or b);
    layer0_outputs(2742) <= not (a or b);
    layer0_outputs(2743) <= not (a xor b);
    layer0_outputs(2744) <= a or b;
    layer0_outputs(2745) <= a and not b;
    layer0_outputs(2746) <= a and b;
    layer0_outputs(2747) <= not (a or b);
    layer0_outputs(2748) <= a xor b;
    layer0_outputs(2749) <= not a or b;
    layer0_outputs(2750) <= a or b;
    layer0_outputs(2751) <= not a;
    layer0_outputs(2752) <= not a;
    layer0_outputs(2753) <= b;
    layer0_outputs(2754) <= a;
    layer0_outputs(2755) <= not (a xor b);
    layer0_outputs(2756) <= not a or b;
    layer0_outputs(2757) <= b;
    layer0_outputs(2758) <= not b or a;
    layer0_outputs(2759) <= not (a xor b);
    layer0_outputs(2760) <= a xor b;
    layer0_outputs(2761) <= a and b;
    layer0_outputs(2762) <= not a;
    layer0_outputs(2763) <= a xor b;
    layer0_outputs(2764) <= 1'b1;
    layer0_outputs(2765) <= b;
    layer0_outputs(2766) <= not (a and b);
    layer0_outputs(2767) <= not (a or b);
    layer0_outputs(2768) <= a or b;
    layer0_outputs(2769) <= not b or a;
    layer0_outputs(2770) <= not a or b;
    layer0_outputs(2771) <= not (a xor b);
    layer0_outputs(2772) <= not b or a;
    layer0_outputs(2773) <= a xor b;
    layer0_outputs(2774) <= a or b;
    layer0_outputs(2775) <= a;
    layer0_outputs(2776) <= not (a xor b);
    layer0_outputs(2777) <= not (a xor b);
    layer0_outputs(2778) <= not b or a;
    layer0_outputs(2779) <= not b;
    layer0_outputs(2780) <= not b or a;
    layer0_outputs(2781) <= not (a xor b);
    layer0_outputs(2782) <= not b or a;
    layer0_outputs(2783) <= a;
    layer0_outputs(2784) <= not b;
    layer0_outputs(2785) <= a and b;
    layer0_outputs(2786) <= a xor b;
    layer0_outputs(2787) <= a or b;
    layer0_outputs(2788) <= not (a and b);
    layer0_outputs(2789) <= not b;
    layer0_outputs(2790) <= not (a or b);
    layer0_outputs(2791) <= not (a xor b);
    layer0_outputs(2792) <= not b or a;
    layer0_outputs(2793) <= a or b;
    layer0_outputs(2794) <= b;
    layer0_outputs(2795) <= not (a or b);
    layer0_outputs(2796) <= not (a xor b);
    layer0_outputs(2797) <= not (a or b);
    layer0_outputs(2798) <= not (a xor b);
    layer0_outputs(2799) <= not a or b;
    layer0_outputs(2800) <= a;
    layer0_outputs(2801) <= b and not a;
    layer0_outputs(2802) <= a or b;
    layer0_outputs(2803) <= not (a and b);
    layer0_outputs(2804) <= not (a xor b);
    layer0_outputs(2805) <= b;
    layer0_outputs(2806) <= not a or b;
    layer0_outputs(2807) <= not (a xor b);
    layer0_outputs(2808) <= not (a xor b);
    layer0_outputs(2809) <= not b;
    layer0_outputs(2810) <= a or b;
    layer0_outputs(2811) <= a or b;
    layer0_outputs(2812) <= not (a or b);
    layer0_outputs(2813) <= not (a xor b);
    layer0_outputs(2814) <= not b or a;
    layer0_outputs(2815) <= not (a xor b);
    layer0_outputs(2816) <= not (a xor b);
    layer0_outputs(2817) <= not (a or b);
    layer0_outputs(2818) <= a or b;
    layer0_outputs(2819) <= a or b;
    layer0_outputs(2820) <= not a or b;
    layer0_outputs(2821) <= not a;
    layer0_outputs(2822) <= 1'b0;
    layer0_outputs(2823) <= a or b;
    layer0_outputs(2824) <= 1'b0;
    layer0_outputs(2825) <= b and not a;
    layer0_outputs(2826) <= b;
    layer0_outputs(2827) <= a;
    layer0_outputs(2828) <= a xor b;
    layer0_outputs(2829) <= a and not b;
    layer0_outputs(2830) <= a or b;
    layer0_outputs(2831) <= 1'b1;
    layer0_outputs(2832) <= not (a xor b);
    layer0_outputs(2833) <= not (a xor b);
    layer0_outputs(2834) <= not (a or b);
    layer0_outputs(2835) <= b and not a;
    layer0_outputs(2836) <= not a or b;
    layer0_outputs(2837) <= a and not b;
    layer0_outputs(2838) <= not a or b;
    layer0_outputs(2839) <= a or b;
    layer0_outputs(2840) <= not a;
    layer0_outputs(2841) <= not (a xor b);
    layer0_outputs(2842) <= a and b;
    layer0_outputs(2843) <= 1'b0;
    layer0_outputs(2844) <= not b or a;
    layer0_outputs(2845) <= a and not b;
    layer0_outputs(2846) <= not a or b;
    layer0_outputs(2847) <= a or b;
    layer0_outputs(2848) <= not a;
    layer0_outputs(2849) <= not a or b;
    layer0_outputs(2850) <= not (a or b);
    layer0_outputs(2851) <= not (a or b);
    layer0_outputs(2852) <= b and not a;
    layer0_outputs(2853) <= not b or a;
    layer0_outputs(2854) <= a or b;
    layer0_outputs(2855) <= a or b;
    layer0_outputs(2856) <= not (a or b);
    layer0_outputs(2857) <= not (a xor b);
    layer0_outputs(2858) <= not b;
    layer0_outputs(2859) <= not (a or b);
    layer0_outputs(2860) <= b and not a;
    layer0_outputs(2861) <= a or b;
    layer0_outputs(2862) <= a or b;
    layer0_outputs(2863) <= a or b;
    layer0_outputs(2864) <= not a or b;
    layer0_outputs(2865) <= a xor b;
    layer0_outputs(2866) <= a and not b;
    layer0_outputs(2867) <= a;
    layer0_outputs(2868) <= a;
    layer0_outputs(2869) <= not (a xor b);
    layer0_outputs(2870) <= not (a or b);
    layer0_outputs(2871) <= a;
    layer0_outputs(2872) <= a and not b;
    layer0_outputs(2873) <= not (a xor b);
    layer0_outputs(2874) <= not a or b;
    layer0_outputs(2875) <= not (a xor b);
    layer0_outputs(2876) <= a xor b;
    layer0_outputs(2877) <= a or b;
    layer0_outputs(2878) <= not (a xor b);
    layer0_outputs(2879) <= not a;
    layer0_outputs(2880) <= not (a or b);
    layer0_outputs(2881) <= not (a or b);
    layer0_outputs(2882) <= 1'b1;
    layer0_outputs(2883) <= a xor b;
    layer0_outputs(2884) <= a;
    layer0_outputs(2885) <= not b or a;
    layer0_outputs(2886) <= a;
    layer0_outputs(2887) <= not (a xor b);
    layer0_outputs(2888) <= b;
    layer0_outputs(2889) <= a and not b;
    layer0_outputs(2890) <= a xor b;
    layer0_outputs(2891) <= not (a or b);
    layer0_outputs(2892) <= a;
    layer0_outputs(2893) <= a xor b;
    layer0_outputs(2894) <= b;
    layer0_outputs(2895) <= a and not b;
    layer0_outputs(2896) <= a;
    layer0_outputs(2897) <= not a or b;
    layer0_outputs(2898) <= not (a or b);
    layer0_outputs(2899) <= a xor b;
    layer0_outputs(2900) <= not (a or b);
    layer0_outputs(2901) <= a xor b;
    layer0_outputs(2902) <= b;
    layer0_outputs(2903) <= 1'b0;
    layer0_outputs(2904) <= not a;
    layer0_outputs(2905) <= a;
    layer0_outputs(2906) <= a xor b;
    layer0_outputs(2907) <= not b or a;
    layer0_outputs(2908) <= a and b;
    layer0_outputs(2909) <= b;
    layer0_outputs(2910) <= a or b;
    layer0_outputs(2911) <= a or b;
    layer0_outputs(2912) <= not a or b;
    layer0_outputs(2913) <= not a;
    layer0_outputs(2914) <= not a or b;
    layer0_outputs(2915) <= not b;
    layer0_outputs(2916) <= a;
    layer0_outputs(2917) <= not a or b;
    layer0_outputs(2918) <= not (a xor b);
    layer0_outputs(2919) <= not (a or b);
    layer0_outputs(2920) <= a and not b;
    layer0_outputs(2921) <= a;
    layer0_outputs(2922) <= not (a xor b);
    layer0_outputs(2923) <= not b;
    layer0_outputs(2924) <= a;
    layer0_outputs(2925) <= not a or b;
    layer0_outputs(2926) <= a or b;
    layer0_outputs(2927) <= not b;
    layer0_outputs(2928) <= not a or b;
    layer0_outputs(2929) <= a or b;
    layer0_outputs(2930) <= not (a or b);
    layer0_outputs(2931) <= not (a or b);
    layer0_outputs(2932) <= not (a xor b);
    layer0_outputs(2933) <= a xor b;
    layer0_outputs(2934) <= not b;
    layer0_outputs(2935) <= a xor b;
    layer0_outputs(2936) <= b and not a;
    layer0_outputs(2937) <= a or b;
    layer0_outputs(2938) <= not (a xor b);
    layer0_outputs(2939) <= not a or b;
    layer0_outputs(2940) <= a;
    layer0_outputs(2941) <= not (a and b);
    layer0_outputs(2942) <= 1'b1;
    layer0_outputs(2943) <= a or b;
    layer0_outputs(2944) <= not (a or b);
    layer0_outputs(2945) <= not (a or b);
    layer0_outputs(2946) <= a and not b;
    layer0_outputs(2947) <= not (a or b);
    layer0_outputs(2948) <= a and not b;
    layer0_outputs(2949) <= a and not b;
    layer0_outputs(2950) <= b and not a;
    layer0_outputs(2951) <= not b or a;
    layer0_outputs(2952) <= 1'b1;
    layer0_outputs(2953) <= not b;
    layer0_outputs(2954) <= not (a xor b);
    layer0_outputs(2955) <= a xor b;
    layer0_outputs(2956) <= a xor b;
    layer0_outputs(2957) <= a xor b;
    layer0_outputs(2958) <= a and b;
    layer0_outputs(2959) <= a and not b;
    layer0_outputs(2960) <= not (a or b);
    layer0_outputs(2961) <= not b or a;
    layer0_outputs(2962) <= a;
    layer0_outputs(2963) <= not a;
    layer0_outputs(2964) <= a xor b;
    layer0_outputs(2965) <= not (a or b);
    layer0_outputs(2966) <= a or b;
    layer0_outputs(2967) <= b;
    layer0_outputs(2968) <= a or b;
    layer0_outputs(2969) <= a xor b;
    layer0_outputs(2970) <= b and not a;
    layer0_outputs(2971) <= not (a and b);
    layer0_outputs(2972) <= a;
    layer0_outputs(2973) <= a;
    layer0_outputs(2974) <= 1'b0;
    layer0_outputs(2975) <= not b;
    layer0_outputs(2976) <= not a;
    layer0_outputs(2977) <= not a or b;
    layer0_outputs(2978) <= not (a or b);
    layer0_outputs(2979) <= b and not a;
    layer0_outputs(2980) <= not b or a;
    layer0_outputs(2981) <= not a;
    layer0_outputs(2982) <= not a;
    layer0_outputs(2983) <= not (a xor b);
    layer0_outputs(2984) <= a xor b;
    layer0_outputs(2985) <= a xor b;
    layer0_outputs(2986) <= not (a xor b);
    layer0_outputs(2987) <= not (a xor b);
    layer0_outputs(2988) <= b;
    layer0_outputs(2989) <= not b or a;
    layer0_outputs(2990) <= a or b;
    layer0_outputs(2991) <= not b or a;
    layer0_outputs(2992) <= a or b;
    layer0_outputs(2993) <= not a or b;
    layer0_outputs(2994) <= not (a xor b);
    layer0_outputs(2995) <= not b or a;
    layer0_outputs(2996) <= a and b;
    layer0_outputs(2997) <= not a;
    layer0_outputs(2998) <= not b or a;
    layer0_outputs(2999) <= not a or b;
    layer0_outputs(3000) <= 1'b1;
    layer0_outputs(3001) <= not b or a;
    layer0_outputs(3002) <= not a;
    layer0_outputs(3003) <= b and not a;
    layer0_outputs(3004) <= not (a or b);
    layer0_outputs(3005) <= not (a xor b);
    layer0_outputs(3006) <= 1'b1;
    layer0_outputs(3007) <= not (a and b);
    layer0_outputs(3008) <= not a;
    layer0_outputs(3009) <= a and not b;
    layer0_outputs(3010) <= b and not a;
    layer0_outputs(3011) <= a and not b;
    layer0_outputs(3012) <= not (a and b);
    layer0_outputs(3013) <= not a;
    layer0_outputs(3014) <= b and not a;
    layer0_outputs(3015) <= a and not b;
    layer0_outputs(3016) <= a;
    layer0_outputs(3017) <= not (a and b);
    layer0_outputs(3018) <= not a;
    layer0_outputs(3019) <= b and not a;
    layer0_outputs(3020) <= 1'b1;
    layer0_outputs(3021) <= b and not a;
    layer0_outputs(3022) <= b;
    layer0_outputs(3023) <= not a or b;
    layer0_outputs(3024) <= a or b;
    layer0_outputs(3025) <= not (a xor b);
    layer0_outputs(3026) <= not (a and b);
    layer0_outputs(3027) <= not b;
    layer0_outputs(3028) <= a or b;
    layer0_outputs(3029) <= not a;
    layer0_outputs(3030) <= not b or a;
    layer0_outputs(3031) <= not b;
    layer0_outputs(3032) <= a and b;
    layer0_outputs(3033) <= a;
    layer0_outputs(3034) <= b;
    layer0_outputs(3035) <= not b;
    layer0_outputs(3036) <= b and not a;
    layer0_outputs(3037) <= not a or b;
    layer0_outputs(3038) <= not b;
    layer0_outputs(3039) <= not a;
    layer0_outputs(3040) <= not (a xor b);
    layer0_outputs(3041) <= a xor b;
    layer0_outputs(3042) <= b and not a;
    layer0_outputs(3043) <= b;
    layer0_outputs(3044) <= a or b;
    layer0_outputs(3045) <= not a;
    layer0_outputs(3046) <= not (a or b);
    layer0_outputs(3047) <= 1'b1;
    layer0_outputs(3048) <= a and b;
    layer0_outputs(3049) <= a and b;
    layer0_outputs(3050) <= a and b;
    layer0_outputs(3051) <= not (a xor b);
    layer0_outputs(3052) <= a xor b;
    layer0_outputs(3053) <= a and not b;
    layer0_outputs(3054) <= not a or b;
    layer0_outputs(3055) <= b;
    layer0_outputs(3056) <= not b;
    layer0_outputs(3057) <= a and b;
    layer0_outputs(3058) <= not b or a;
    layer0_outputs(3059) <= a;
    layer0_outputs(3060) <= a xor b;
    layer0_outputs(3061) <= a or b;
    layer0_outputs(3062) <= not b or a;
    layer0_outputs(3063) <= b;
    layer0_outputs(3064) <= a or b;
    layer0_outputs(3065) <= not a or b;
    layer0_outputs(3066) <= a and b;
    layer0_outputs(3067) <= 1'b1;
    layer0_outputs(3068) <= a xor b;
    layer0_outputs(3069) <= not b or a;
    layer0_outputs(3070) <= a xor b;
    layer0_outputs(3071) <= a or b;
    layer0_outputs(3072) <= b;
    layer0_outputs(3073) <= not b or a;
    layer0_outputs(3074) <= not (a xor b);
    layer0_outputs(3075) <= 1'b1;
    layer0_outputs(3076) <= a;
    layer0_outputs(3077) <= 1'b1;
    layer0_outputs(3078) <= not a;
    layer0_outputs(3079) <= not a;
    layer0_outputs(3080) <= b;
    layer0_outputs(3081) <= not (a xor b);
    layer0_outputs(3082) <= a or b;
    layer0_outputs(3083) <= not b;
    layer0_outputs(3084) <= not a or b;
    layer0_outputs(3085) <= not b;
    layer0_outputs(3086) <= not b;
    layer0_outputs(3087) <= not (a xor b);
    layer0_outputs(3088) <= not (a xor b);
    layer0_outputs(3089) <= a or b;
    layer0_outputs(3090) <= not (a xor b);
    layer0_outputs(3091) <= not (a or b);
    layer0_outputs(3092) <= not (a xor b);
    layer0_outputs(3093) <= not (a or b);
    layer0_outputs(3094) <= not (a xor b);
    layer0_outputs(3095) <= not b;
    layer0_outputs(3096) <= a xor b;
    layer0_outputs(3097) <= b;
    layer0_outputs(3098) <= not b;
    layer0_outputs(3099) <= a;
    layer0_outputs(3100) <= not (a or b);
    layer0_outputs(3101) <= not b;
    layer0_outputs(3102) <= not b or a;
    layer0_outputs(3103) <= not b;
    layer0_outputs(3104) <= not a;
    layer0_outputs(3105) <= a xor b;
    layer0_outputs(3106) <= not (a xor b);
    layer0_outputs(3107) <= a or b;
    layer0_outputs(3108) <= not (a or b);
    layer0_outputs(3109) <= a;
    layer0_outputs(3110) <= not (a or b);
    layer0_outputs(3111) <= a or b;
    layer0_outputs(3112) <= not a;
    layer0_outputs(3113) <= not a or b;
    layer0_outputs(3114) <= not (a or b);
    layer0_outputs(3115) <= a and not b;
    layer0_outputs(3116) <= a or b;
    layer0_outputs(3117) <= not b or a;
    layer0_outputs(3118) <= a xor b;
    layer0_outputs(3119) <= not (a or b);
    layer0_outputs(3120) <= b;
    layer0_outputs(3121) <= a xor b;
    layer0_outputs(3122) <= not (a or b);
    layer0_outputs(3123) <= a xor b;
    layer0_outputs(3124) <= not (a xor b);
    layer0_outputs(3125) <= a xor b;
    layer0_outputs(3126) <= a and b;
    layer0_outputs(3127) <= not (a xor b);
    layer0_outputs(3128) <= b;
    layer0_outputs(3129) <= not a or b;
    layer0_outputs(3130) <= not (a or b);
    layer0_outputs(3131) <= not (a or b);
    layer0_outputs(3132) <= not (a and b);
    layer0_outputs(3133) <= not (a or b);
    layer0_outputs(3134) <= a or b;
    layer0_outputs(3135) <= a and not b;
    layer0_outputs(3136) <= a or b;
    layer0_outputs(3137) <= not (a and b);
    layer0_outputs(3138) <= not a;
    layer0_outputs(3139) <= b;
    layer0_outputs(3140) <= not b;
    layer0_outputs(3141) <= a xor b;
    layer0_outputs(3142) <= a;
    layer0_outputs(3143) <= b;
    layer0_outputs(3144) <= b and not a;
    layer0_outputs(3145) <= b and not a;
    layer0_outputs(3146) <= not b or a;
    layer0_outputs(3147) <= not b or a;
    layer0_outputs(3148) <= a xor b;
    layer0_outputs(3149) <= not (a or b);
    layer0_outputs(3150) <= a or b;
    layer0_outputs(3151) <= a xor b;
    layer0_outputs(3152) <= not (a or b);
    layer0_outputs(3153) <= not b or a;
    layer0_outputs(3154) <= not (a or b);
    layer0_outputs(3155) <= a xor b;
    layer0_outputs(3156) <= not a or b;
    layer0_outputs(3157) <= a;
    layer0_outputs(3158) <= not b;
    layer0_outputs(3159) <= not a or b;
    layer0_outputs(3160) <= not a or b;
    layer0_outputs(3161) <= a and b;
    layer0_outputs(3162) <= not (a xor b);
    layer0_outputs(3163) <= not (a xor b);
    layer0_outputs(3164) <= not (a or b);
    layer0_outputs(3165) <= b and not a;
    layer0_outputs(3166) <= not (a xor b);
    layer0_outputs(3167) <= not (a or b);
    layer0_outputs(3168) <= b and not a;
    layer0_outputs(3169) <= not a;
    layer0_outputs(3170) <= a or b;
    layer0_outputs(3171) <= b and not a;
    layer0_outputs(3172) <= a xor b;
    layer0_outputs(3173) <= a xor b;
    layer0_outputs(3174) <= not a;
    layer0_outputs(3175) <= a and b;
    layer0_outputs(3176) <= b;
    layer0_outputs(3177) <= not b;
    layer0_outputs(3178) <= a xor b;
    layer0_outputs(3179) <= a or b;
    layer0_outputs(3180) <= not (a xor b);
    layer0_outputs(3181) <= not (a or b);
    layer0_outputs(3182) <= a xor b;
    layer0_outputs(3183) <= not b or a;
    layer0_outputs(3184) <= not (a xor b);
    layer0_outputs(3185) <= not (a or b);
    layer0_outputs(3186) <= a xor b;
    layer0_outputs(3187) <= a;
    layer0_outputs(3188) <= a xor b;
    layer0_outputs(3189) <= not b;
    layer0_outputs(3190) <= a;
    layer0_outputs(3191) <= not (a xor b);
    layer0_outputs(3192) <= not (a xor b);
    layer0_outputs(3193) <= a or b;
    layer0_outputs(3194) <= b and not a;
    layer0_outputs(3195) <= a or b;
    layer0_outputs(3196) <= not b or a;
    layer0_outputs(3197) <= not a;
    layer0_outputs(3198) <= a or b;
    layer0_outputs(3199) <= not (a xor b);
    layer0_outputs(3200) <= a or b;
    layer0_outputs(3201) <= a xor b;
    layer0_outputs(3202) <= a and b;
    layer0_outputs(3203) <= not (a or b);
    layer0_outputs(3204) <= b;
    layer0_outputs(3205) <= a;
    layer0_outputs(3206) <= a or b;
    layer0_outputs(3207) <= a;
    layer0_outputs(3208) <= b;
    layer0_outputs(3209) <= a and not b;
    layer0_outputs(3210) <= a or b;
    layer0_outputs(3211) <= a xor b;
    layer0_outputs(3212) <= not (a or b);
    layer0_outputs(3213) <= not b or a;
    layer0_outputs(3214) <= a and not b;
    layer0_outputs(3215) <= not a or b;
    layer0_outputs(3216) <= b;
    layer0_outputs(3217) <= not b;
    layer0_outputs(3218) <= a;
    layer0_outputs(3219) <= not b or a;
    layer0_outputs(3220) <= a and not b;
    layer0_outputs(3221) <= not (a or b);
    layer0_outputs(3222) <= not (a xor b);
    layer0_outputs(3223) <= not (a or b);
    layer0_outputs(3224) <= a;
    layer0_outputs(3225) <= a;
    layer0_outputs(3226) <= not (a xor b);
    layer0_outputs(3227) <= b and not a;
    layer0_outputs(3228) <= not a or b;
    layer0_outputs(3229) <= a xor b;
    layer0_outputs(3230) <= 1'b1;
    layer0_outputs(3231) <= a or b;
    layer0_outputs(3232) <= a or b;
    layer0_outputs(3233) <= 1'b1;
    layer0_outputs(3234) <= not (a or b);
    layer0_outputs(3235) <= b;
    layer0_outputs(3236) <= not (a or b);
    layer0_outputs(3237) <= not b or a;
    layer0_outputs(3238) <= b and not a;
    layer0_outputs(3239) <= not (a or b);
    layer0_outputs(3240) <= a and b;
    layer0_outputs(3241) <= not a or b;
    layer0_outputs(3242) <= not a or b;
    layer0_outputs(3243) <= not (a xor b);
    layer0_outputs(3244) <= not (a xor b);
    layer0_outputs(3245) <= not (a or b);
    layer0_outputs(3246) <= a and b;
    layer0_outputs(3247) <= b;
    layer0_outputs(3248) <= a or b;
    layer0_outputs(3249) <= not (a or b);
    layer0_outputs(3250) <= not (a or b);
    layer0_outputs(3251) <= a xor b;
    layer0_outputs(3252) <= not b;
    layer0_outputs(3253) <= not (a xor b);
    layer0_outputs(3254) <= not a or b;
    layer0_outputs(3255) <= a xor b;
    layer0_outputs(3256) <= a or b;
    layer0_outputs(3257) <= not (a xor b);
    layer0_outputs(3258) <= a or b;
    layer0_outputs(3259) <= b and not a;
    layer0_outputs(3260) <= a and not b;
    layer0_outputs(3261) <= not b or a;
    layer0_outputs(3262) <= not (a or b);
    layer0_outputs(3263) <= not (a xor b);
    layer0_outputs(3264) <= a and not b;
    layer0_outputs(3265) <= a or b;
    layer0_outputs(3266) <= b;
    layer0_outputs(3267) <= a and b;
    layer0_outputs(3268) <= a;
    layer0_outputs(3269) <= not b;
    layer0_outputs(3270) <= not (a xor b);
    layer0_outputs(3271) <= a;
    layer0_outputs(3272) <= not b or a;
    layer0_outputs(3273) <= a and not b;
    layer0_outputs(3274) <= a xor b;
    layer0_outputs(3275) <= not a or b;
    layer0_outputs(3276) <= a or b;
    layer0_outputs(3277) <= not b;
    layer0_outputs(3278) <= a and not b;
    layer0_outputs(3279) <= not a;
    layer0_outputs(3280) <= a;
    layer0_outputs(3281) <= a;
    layer0_outputs(3282) <= not a or b;
    layer0_outputs(3283) <= not (a xor b);
    layer0_outputs(3284) <= not a;
    layer0_outputs(3285) <= not (a xor b);
    layer0_outputs(3286) <= not (a or b);
    layer0_outputs(3287) <= not b;
    layer0_outputs(3288) <= not (a or b);
    layer0_outputs(3289) <= not a or b;
    layer0_outputs(3290) <= a xor b;
    layer0_outputs(3291) <= a;
    layer0_outputs(3292) <= b;
    layer0_outputs(3293) <= a;
    layer0_outputs(3294) <= a or b;
    layer0_outputs(3295) <= not a;
    layer0_outputs(3296) <= a or b;
    layer0_outputs(3297) <= a or b;
    layer0_outputs(3298) <= not (a or b);
    layer0_outputs(3299) <= not (a xor b);
    layer0_outputs(3300) <= a and not b;
    layer0_outputs(3301) <= not b or a;
    layer0_outputs(3302) <= a xor b;
    layer0_outputs(3303) <= not b;
    layer0_outputs(3304) <= not b;
    layer0_outputs(3305) <= b and not a;
    layer0_outputs(3306) <= not b;
    layer0_outputs(3307) <= not (a or b);
    layer0_outputs(3308) <= a xor b;
    layer0_outputs(3309) <= a;
    layer0_outputs(3310) <= b;
    layer0_outputs(3311) <= not (a xor b);
    layer0_outputs(3312) <= not a or b;
    layer0_outputs(3313) <= not (a or b);
    layer0_outputs(3314) <= a xor b;
    layer0_outputs(3315) <= not b or a;
    layer0_outputs(3316) <= a or b;
    layer0_outputs(3317) <= not a or b;
    layer0_outputs(3318) <= b and not a;
    layer0_outputs(3319) <= a xor b;
    layer0_outputs(3320) <= not (a or b);
    layer0_outputs(3321) <= b;
    layer0_outputs(3322) <= a or b;
    layer0_outputs(3323) <= a;
    layer0_outputs(3324) <= a or b;
    layer0_outputs(3325) <= b;
    layer0_outputs(3326) <= not (a xor b);
    layer0_outputs(3327) <= not a or b;
    layer0_outputs(3328) <= not b;
    layer0_outputs(3329) <= not (a xor b);
    layer0_outputs(3330) <= not (a xor b);
    layer0_outputs(3331) <= not (a and b);
    layer0_outputs(3332) <= not a;
    layer0_outputs(3333) <= not (a xor b);
    layer0_outputs(3334) <= not (a or b);
    layer0_outputs(3335) <= a or b;
    layer0_outputs(3336) <= not (a or b);
    layer0_outputs(3337) <= 1'b1;
    layer0_outputs(3338) <= not (a xor b);
    layer0_outputs(3339) <= b and not a;
    layer0_outputs(3340) <= b and not a;
    layer0_outputs(3341) <= not (a xor b);
    layer0_outputs(3342) <= a and not b;
    layer0_outputs(3343) <= b and not a;
    layer0_outputs(3344) <= a or b;
    layer0_outputs(3345) <= not a or b;
    layer0_outputs(3346) <= 1'b0;
    layer0_outputs(3347) <= not b or a;
    layer0_outputs(3348) <= a or b;
    layer0_outputs(3349) <= not (a xor b);
    layer0_outputs(3350) <= b and not a;
    layer0_outputs(3351) <= a xor b;
    layer0_outputs(3352) <= not b;
    layer0_outputs(3353) <= not a;
    layer0_outputs(3354) <= b;
    layer0_outputs(3355) <= not (a xor b);
    layer0_outputs(3356) <= a or b;
    layer0_outputs(3357) <= a or b;
    layer0_outputs(3358) <= not a;
    layer0_outputs(3359) <= not a;
    layer0_outputs(3360) <= not a or b;
    layer0_outputs(3361) <= a or b;
    layer0_outputs(3362) <= not a;
    layer0_outputs(3363) <= not (a xor b);
    layer0_outputs(3364) <= not a or b;
    layer0_outputs(3365) <= a xor b;
    layer0_outputs(3366) <= not a;
    layer0_outputs(3367) <= not (a or b);
    layer0_outputs(3368) <= a or b;
    layer0_outputs(3369) <= not (a or b);
    layer0_outputs(3370) <= not b;
    layer0_outputs(3371) <= not a or b;
    layer0_outputs(3372) <= 1'b0;
    layer0_outputs(3373) <= not (a xor b);
    layer0_outputs(3374) <= not (a or b);
    layer0_outputs(3375) <= not (a or b);
    layer0_outputs(3376) <= not (a or b);
    layer0_outputs(3377) <= a xor b;
    layer0_outputs(3378) <= not (a or b);
    layer0_outputs(3379) <= not b;
    layer0_outputs(3380) <= not a or b;
    layer0_outputs(3381) <= not b or a;
    layer0_outputs(3382) <= not b;
    layer0_outputs(3383) <= not (a xor b);
    layer0_outputs(3384) <= not a or b;
    layer0_outputs(3385) <= 1'b1;
    layer0_outputs(3386) <= a and not b;
    layer0_outputs(3387) <= not a;
    layer0_outputs(3388) <= not (a xor b);
    layer0_outputs(3389) <= not (a xor b);
    layer0_outputs(3390) <= not (a or b);
    layer0_outputs(3391) <= not a or b;
    layer0_outputs(3392) <= not (a or b);
    layer0_outputs(3393) <= a and not b;
    layer0_outputs(3394) <= a or b;
    layer0_outputs(3395) <= a;
    layer0_outputs(3396) <= b and not a;
    layer0_outputs(3397) <= a or b;
    layer0_outputs(3398) <= not (a and b);
    layer0_outputs(3399) <= not a or b;
    layer0_outputs(3400) <= not b;
    layer0_outputs(3401) <= a;
    layer0_outputs(3402) <= not a or b;
    layer0_outputs(3403) <= not b or a;
    layer0_outputs(3404) <= not a or b;
    layer0_outputs(3405) <= not (a or b);
    layer0_outputs(3406) <= not (a xor b);
    layer0_outputs(3407) <= a or b;
    layer0_outputs(3408) <= a and not b;
    layer0_outputs(3409) <= not a;
    layer0_outputs(3410) <= a or b;
    layer0_outputs(3411) <= a;
    layer0_outputs(3412) <= not (a xor b);
    layer0_outputs(3413) <= not b or a;
    layer0_outputs(3414) <= not (a xor b);
    layer0_outputs(3415) <= a or b;
    layer0_outputs(3416) <= a;
    layer0_outputs(3417) <= b;
    layer0_outputs(3418) <= a and not b;
    layer0_outputs(3419) <= not (a or b);
    layer0_outputs(3420) <= a or b;
    layer0_outputs(3421) <= not b or a;
    layer0_outputs(3422) <= not a or b;
    layer0_outputs(3423) <= a or b;
    layer0_outputs(3424) <= a or b;
    layer0_outputs(3425) <= a and not b;
    layer0_outputs(3426) <= a xor b;
    layer0_outputs(3427) <= not (a or b);
    layer0_outputs(3428) <= not b;
    layer0_outputs(3429) <= b;
    layer0_outputs(3430) <= not b;
    layer0_outputs(3431) <= 1'b0;
    layer0_outputs(3432) <= a or b;
    layer0_outputs(3433) <= not b or a;
    layer0_outputs(3434) <= not (a xor b);
    layer0_outputs(3435) <= a and not b;
    layer0_outputs(3436) <= not (a xor b);
    layer0_outputs(3437) <= a or b;
    layer0_outputs(3438) <= a xor b;
    layer0_outputs(3439) <= b and not a;
    layer0_outputs(3440) <= b;
    layer0_outputs(3441) <= a xor b;
    layer0_outputs(3442) <= a and not b;
    layer0_outputs(3443) <= a xor b;
    layer0_outputs(3444) <= not a;
    layer0_outputs(3445) <= not (a or b);
    layer0_outputs(3446) <= not (a or b);
    layer0_outputs(3447) <= not b;
    layer0_outputs(3448) <= a;
    layer0_outputs(3449) <= not (a or b);
    layer0_outputs(3450) <= not (a xor b);
    layer0_outputs(3451) <= not b or a;
    layer0_outputs(3452) <= not (a or b);
    layer0_outputs(3453) <= not b or a;
    layer0_outputs(3454) <= not b;
    layer0_outputs(3455) <= a or b;
    layer0_outputs(3456) <= a xor b;
    layer0_outputs(3457) <= b;
    layer0_outputs(3458) <= not a or b;
    layer0_outputs(3459) <= not a;
    layer0_outputs(3460) <= not b or a;
    layer0_outputs(3461) <= b and not a;
    layer0_outputs(3462) <= b and not a;
    layer0_outputs(3463) <= a and not b;
    layer0_outputs(3464) <= a xor b;
    layer0_outputs(3465) <= a or b;
    layer0_outputs(3466) <= a and not b;
    layer0_outputs(3467) <= not a;
    layer0_outputs(3468) <= not (a xor b);
    layer0_outputs(3469) <= not b or a;
    layer0_outputs(3470) <= not a or b;
    layer0_outputs(3471) <= 1'b0;
    layer0_outputs(3472) <= 1'b1;
    layer0_outputs(3473) <= a and not b;
    layer0_outputs(3474) <= b;
    layer0_outputs(3475) <= b and not a;
    layer0_outputs(3476) <= not (a xor b);
    layer0_outputs(3477) <= not (a or b);
    layer0_outputs(3478) <= a or b;
    layer0_outputs(3479) <= a or b;
    layer0_outputs(3480) <= a xor b;
    layer0_outputs(3481) <= a or b;
    layer0_outputs(3482) <= a;
    layer0_outputs(3483) <= b and not a;
    layer0_outputs(3484) <= not a or b;
    layer0_outputs(3485) <= not (a or b);
    layer0_outputs(3486) <= a;
    layer0_outputs(3487) <= b and not a;
    layer0_outputs(3488) <= not (a or b);
    layer0_outputs(3489) <= not (a xor b);
    layer0_outputs(3490) <= a or b;
    layer0_outputs(3491) <= 1'b1;
    layer0_outputs(3492) <= b;
    layer0_outputs(3493) <= a xor b;
    layer0_outputs(3494) <= not (a or b);
    layer0_outputs(3495) <= not (a and b);
    layer0_outputs(3496) <= not b;
    layer0_outputs(3497) <= a or b;
    layer0_outputs(3498) <= a;
    layer0_outputs(3499) <= a or b;
    layer0_outputs(3500) <= a;
    layer0_outputs(3501) <= not (a xor b);
    layer0_outputs(3502) <= a or b;
    layer0_outputs(3503) <= not a or b;
    layer0_outputs(3504) <= not b;
    layer0_outputs(3505) <= a;
    layer0_outputs(3506) <= b;
    layer0_outputs(3507) <= a and not b;
    layer0_outputs(3508) <= not a or b;
    layer0_outputs(3509) <= a and not b;
    layer0_outputs(3510) <= not (a xor b);
    layer0_outputs(3511) <= a or b;
    layer0_outputs(3512) <= a or b;
    layer0_outputs(3513) <= not a;
    layer0_outputs(3514) <= not (a xor b);
    layer0_outputs(3515) <= a or b;
    layer0_outputs(3516) <= not b or a;
    layer0_outputs(3517) <= a and b;
    layer0_outputs(3518) <= a or b;
    layer0_outputs(3519) <= not a;
    layer0_outputs(3520) <= a or b;
    layer0_outputs(3521) <= a xor b;
    layer0_outputs(3522) <= not (a xor b);
    layer0_outputs(3523) <= not a;
    layer0_outputs(3524) <= a;
    layer0_outputs(3525) <= b;
    layer0_outputs(3526) <= a and not b;
    layer0_outputs(3527) <= b;
    layer0_outputs(3528) <= b;
    layer0_outputs(3529) <= not (a and b);
    layer0_outputs(3530) <= a;
    layer0_outputs(3531) <= not b;
    layer0_outputs(3532) <= b and not a;
    layer0_outputs(3533) <= not (a or b);
    layer0_outputs(3534) <= not (a xor b);
    layer0_outputs(3535) <= not b;
    layer0_outputs(3536) <= a or b;
    layer0_outputs(3537) <= not a or b;
    layer0_outputs(3538) <= not a or b;
    layer0_outputs(3539) <= not (a xor b);
    layer0_outputs(3540) <= not b;
    layer0_outputs(3541) <= not (a xor b);
    layer0_outputs(3542) <= a;
    layer0_outputs(3543) <= a;
    layer0_outputs(3544) <= not b or a;
    layer0_outputs(3545) <= not (a or b);
    layer0_outputs(3546) <= b and not a;
    layer0_outputs(3547) <= a;
    layer0_outputs(3548) <= not (a or b);
    layer0_outputs(3549) <= not (a xor b);
    layer0_outputs(3550) <= not (a xor b);
    layer0_outputs(3551) <= not b;
    layer0_outputs(3552) <= a and not b;
    layer0_outputs(3553) <= a and b;
    layer0_outputs(3554) <= a;
    layer0_outputs(3555) <= a and not b;
    layer0_outputs(3556) <= a xor b;
    layer0_outputs(3557) <= not (a xor b);
    layer0_outputs(3558) <= not (a or b);
    layer0_outputs(3559) <= not b;
    layer0_outputs(3560) <= a xor b;
    layer0_outputs(3561) <= a or b;
    layer0_outputs(3562) <= b and not a;
    layer0_outputs(3563) <= not a or b;
    layer0_outputs(3564) <= not (a xor b);
    layer0_outputs(3565) <= a;
    layer0_outputs(3566) <= a and b;
    layer0_outputs(3567) <= a;
    layer0_outputs(3568) <= not (a or b);
    layer0_outputs(3569) <= not (a xor b);
    layer0_outputs(3570) <= b and not a;
    layer0_outputs(3571) <= not b or a;
    layer0_outputs(3572) <= not a;
    layer0_outputs(3573) <= a;
    layer0_outputs(3574) <= not b;
    layer0_outputs(3575) <= not b or a;
    layer0_outputs(3576) <= b;
    layer0_outputs(3577) <= a;
    layer0_outputs(3578) <= not (a or b);
    layer0_outputs(3579) <= not (a or b);
    layer0_outputs(3580) <= a xor b;
    layer0_outputs(3581) <= not b or a;
    layer0_outputs(3582) <= not b;
    layer0_outputs(3583) <= a xor b;
    layer0_outputs(3584) <= not (a or b);
    layer0_outputs(3585) <= not a or b;
    layer0_outputs(3586) <= not b or a;
    layer0_outputs(3587) <= not (a xor b);
    layer0_outputs(3588) <= a xor b;
    layer0_outputs(3589) <= a and not b;
    layer0_outputs(3590) <= 1'b1;
    layer0_outputs(3591) <= a and b;
    layer0_outputs(3592) <= a xor b;
    layer0_outputs(3593) <= not a;
    layer0_outputs(3594) <= not (a or b);
    layer0_outputs(3595) <= a or b;
    layer0_outputs(3596) <= not a;
    layer0_outputs(3597) <= not b or a;
    layer0_outputs(3598) <= not (a or b);
    layer0_outputs(3599) <= not (a or b);
    layer0_outputs(3600) <= not b or a;
    layer0_outputs(3601) <= a;
    layer0_outputs(3602) <= not b or a;
    layer0_outputs(3603) <= not (a or b);
    layer0_outputs(3604) <= a xor b;
    layer0_outputs(3605) <= b;
    layer0_outputs(3606) <= 1'b0;
    layer0_outputs(3607) <= a or b;
    layer0_outputs(3608) <= not (a or b);
    layer0_outputs(3609) <= not b or a;
    layer0_outputs(3610) <= not (a xor b);
    layer0_outputs(3611) <= a or b;
    layer0_outputs(3612) <= a and b;
    layer0_outputs(3613) <= not b or a;
    layer0_outputs(3614) <= a or b;
    layer0_outputs(3615) <= a or b;
    layer0_outputs(3616) <= a or b;
    layer0_outputs(3617) <= a xor b;
    layer0_outputs(3618) <= not (a and b);
    layer0_outputs(3619) <= a and not b;
    layer0_outputs(3620) <= a and not b;
    layer0_outputs(3621) <= a or b;
    layer0_outputs(3622) <= not (a or b);
    layer0_outputs(3623) <= not (a or b);
    layer0_outputs(3624) <= 1'b1;
    layer0_outputs(3625) <= a;
    layer0_outputs(3626) <= a;
    layer0_outputs(3627) <= not a or b;
    layer0_outputs(3628) <= not (a or b);
    layer0_outputs(3629) <= not a;
    layer0_outputs(3630) <= not (a xor b);
    layer0_outputs(3631) <= not (a or b);
    layer0_outputs(3632) <= not a or b;
    layer0_outputs(3633) <= not a or b;
    layer0_outputs(3634) <= a and not b;
    layer0_outputs(3635) <= 1'b1;
    layer0_outputs(3636) <= a or b;
    layer0_outputs(3637) <= a xor b;
    layer0_outputs(3638) <= b and not a;
    layer0_outputs(3639) <= not a or b;
    layer0_outputs(3640) <= not a;
    layer0_outputs(3641) <= not b;
    layer0_outputs(3642) <= not b;
    layer0_outputs(3643) <= b and not a;
    layer0_outputs(3644) <= not a;
    layer0_outputs(3645) <= b;
    layer0_outputs(3646) <= a;
    layer0_outputs(3647) <= not b;
    layer0_outputs(3648) <= not (a xor b);
    layer0_outputs(3649) <= not (a xor b);
    layer0_outputs(3650) <= a xor b;
    layer0_outputs(3651) <= not a or b;
    layer0_outputs(3652) <= not (a or b);
    layer0_outputs(3653) <= not a or b;
    layer0_outputs(3654) <= a;
    layer0_outputs(3655) <= not (a xor b);
    layer0_outputs(3656) <= a xor b;
    layer0_outputs(3657) <= a;
    layer0_outputs(3658) <= a and b;
    layer0_outputs(3659) <= not (a or b);
    layer0_outputs(3660) <= b and not a;
    layer0_outputs(3661) <= a xor b;
    layer0_outputs(3662) <= 1'b0;
    layer0_outputs(3663) <= not b;
    layer0_outputs(3664) <= 1'b0;
    layer0_outputs(3665) <= a xor b;
    layer0_outputs(3666) <= not a;
    layer0_outputs(3667) <= a xor b;
    layer0_outputs(3668) <= not (a or b);
    layer0_outputs(3669) <= a xor b;
    layer0_outputs(3670) <= not b or a;
    layer0_outputs(3671) <= not (a or b);
    layer0_outputs(3672) <= a and not b;
    layer0_outputs(3673) <= a and not b;
    layer0_outputs(3674) <= not a or b;
    layer0_outputs(3675) <= b;
    layer0_outputs(3676) <= a;
    layer0_outputs(3677) <= a xor b;
    layer0_outputs(3678) <= b and not a;
    layer0_outputs(3679) <= b;
    layer0_outputs(3680) <= not a or b;
    layer0_outputs(3681) <= a;
    layer0_outputs(3682) <= b and not a;
    layer0_outputs(3683) <= a;
    layer0_outputs(3684) <= b and not a;
    layer0_outputs(3685) <= a;
    layer0_outputs(3686) <= not (a or b);
    layer0_outputs(3687) <= not (a or b);
    layer0_outputs(3688) <= not (a or b);
    layer0_outputs(3689) <= a and not b;
    layer0_outputs(3690) <= not (a and b);
    layer0_outputs(3691) <= not a or b;
    layer0_outputs(3692) <= not (a or b);
    layer0_outputs(3693) <= not b or a;
    layer0_outputs(3694) <= not b or a;
    layer0_outputs(3695) <= a xor b;
    layer0_outputs(3696) <= not a or b;
    layer0_outputs(3697) <= a or b;
    layer0_outputs(3698) <= not (a and b);
    layer0_outputs(3699) <= a xor b;
    layer0_outputs(3700) <= b;
    layer0_outputs(3701) <= not (a xor b);
    layer0_outputs(3702) <= a and b;
    layer0_outputs(3703) <= not a or b;
    layer0_outputs(3704) <= not (a or b);
    layer0_outputs(3705) <= a xor b;
    layer0_outputs(3706) <= b and not a;
    layer0_outputs(3707) <= not a or b;
    layer0_outputs(3708) <= not a or b;
    layer0_outputs(3709) <= not (a or b);
    layer0_outputs(3710) <= not a;
    layer0_outputs(3711) <= not b;
    layer0_outputs(3712) <= a and not b;
    layer0_outputs(3713) <= not b or a;
    layer0_outputs(3714) <= not (a or b);
    layer0_outputs(3715) <= not (a or b);
    layer0_outputs(3716) <= b;
    layer0_outputs(3717) <= not a;
    layer0_outputs(3718) <= not b or a;
    layer0_outputs(3719) <= not a;
    layer0_outputs(3720) <= not a;
    layer0_outputs(3721) <= not (a or b);
    layer0_outputs(3722) <= a xor b;
    layer0_outputs(3723) <= not a or b;
    layer0_outputs(3724) <= not b;
    layer0_outputs(3725) <= 1'b0;
    layer0_outputs(3726) <= b and not a;
    layer0_outputs(3727) <= not b;
    layer0_outputs(3728) <= not a or b;
    layer0_outputs(3729) <= not a;
    layer0_outputs(3730) <= not (a or b);
    layer0_outputs(3731) <= not (a xor b);
    layer0_outputs(3732) <= not b;
    layer0_outputs(3733) <= b and not a;
    layer0_outputs(3734) <= not (a xor b);
    layer0_outputs(3735) <= a or b;
    layer0_outputs(3736) <= a and not b;
    layer0_outputs(3737) <= not b or a;
    layer0_outputs(3738) <= not (a or b);
    layer0_outputs(3739) <= a and not b;
    layer0_outputs(3740) <= a;
    layer0_outputs(3741) <= a xor b;
    layer0_outputs(3742) <= not (a or b);
    layer0_outputs(3743) <= a xor b;
    layer0_outputs(3744) <= b and not a;
    layer0_outputs(3745) <= not (a or b);
    layer0_outputs(3746) <= a and not b;
    layer0_outputs(3747) <= a and not b;
    layer0_outputs(3748) <= not (a and b);
    layer0_outputs(3749) <= not (a or b);
    layer0_outputs(3750) <= not a;
    layer0_outputs(3751) <= not (a xor b);
    layer0_outputs(3752) <= not (a xor b);
    layer0_outputs(3753) <= not a or b;
    layer0_outputs(3754) <= a and not b;
    layer0_outputs(3755) <= a or b;
    layer0_outputs(3756) <= not (a xor b);
    layer0_outputs(3757) <= a or b;
    layer0_outputs(3758) <= b;
    layer0_outputs(3759) <= not a;
    layer0_outputs(3760) <= not (a xor b);
    layer0_outputs(3761) <= not a or b;
    layer0_outputs(3762) <= not (a or b);
    layer0_outputs(3763) <= not a or b;
    layer0_outputs(3764) <= not (a or b);
    layer0_outputs(3765) <= not a;
    layer0_outputs(3766) <= not (a or b);
    layer0_outputs(3767) <= not b;
    layer0_outputs(3768) <= not (a and b);
    layer0_outputs(3769) <= not a;
    layer0_outputs(3770) <= not (a or b);
    layer0_outputs(3771) <= a;
    layer0_outputs(3772) <= not (a xor b);
    layer0_outputs(3773) <= a and not b;
    layer0_outputs(3774) <= not (a xor b);
    layer0_outputs(3775) <= not (a or b);
    layer0_outputs(3776) <= a and not b;
    layer0_outputs(3777) <= a;
    layer0_outputs(3778) <= not b or a;
    layer0_outputs(3779) <= a;
    layer0_outputs(3780) <= 1'b1;
    layer0_outputs(3781) <= b and not a;
    layer0_outputs(3782) <= not (a or b);
    layer0_outputs(3783) <= not (a xor b);
    layer0_outputs(3784) <= not (a and b);
    layer0_outputs(3785) <= not a;
    layer0_outputs(3786) <= 1'b0;
    layer0_outputs(3787) <= not a or b;
    layer0_outputs(3788) <= 1'b1;
    layer0_outputs(3789) <= not (a or b);
    layer0_outputs(3790) <= not a;
    layer0_outputs(3791) <= b;
    layer0_outputs(3792) <= a xor b;
    layer0_outputs(3793) <= b;
    layer0_outputs(3794) <= not b or a;
    layer0_outputs(3795) <= b;
    layer0_outputs(3796) <= not (a or b);
    layer0_outputs(3797) <= 1'b0;
    layer0_outputs(3798) <= not (a xor b);
    layer0_outputs(3799) <= b;
    layer0_outputs(3800) <= not a or b;
    layer0_outputs(3801) <= b;
    layer0_outputs(3802) <= not (a or b);
    layer0_outputs(3803) <= b and not a;
    layer0_outputs(3804) <= a or b;
    layer0_outputs(3805) <= a and not b;
    layer0_outputs(3806) <= a and not b;
    layer0_outputs(3807) <= not b;
    layer0_outputs(3808) <= a xor b;
    layer0_outputs(3809) <= a;
    layer0_outputs(3810) <= 1'b1;
    layer0_outputs(3811) <= not b or a;
    layer0_outputs(3812) <= 1'b1;
    layer0_outputs(3813) <= not (a xor b);
    layer0_outputs(3814) <= a xor b;
    layer0_outputs(3815) <= a xor b;
    layer0_outputs(3816) <= not b or a;
    layer0_outputs(3817) <= a and not b;
    layer0_outputs(3818) <= not b;
    layer0_outputs(3819) <= not b;
    layer0_outputs(3820) <= not (a or b);
    layer0_outputs(3821) <= a;
    layer0_outputs(3822) <= b;
    layer0_outputs(3823) <= not b or a;
    layer0_outputs(3824) <= a and not b;
    layer0_outputs(3825) <= not (a or b);
    layer0_outputs(3826) <= a or b;
    layer0_outputs(3827) <= not (a or b);
    layer0_outputs(3828) <= 1'b1;
    layer0_outputs(3829) <= a xor b;
    layer0_outputs(3830) <= a or b;
    layer0_outputs(3831) <= a xor b;
    layer0_outputs(3832) <= a xor b;
    layer0_outputs(3833) <= 1'b0;
    layer0_outputs(3834) <= b;
    layer0_outputs(3835) <= not a or b;
    layer0_outputs(3836) <= a or b;
    layer0_outputs(3837) <= not (a or b);
    layer0_outputs(3838) <= b;
    layer0_outputs(3839) <= b;
    layer0_outputs(3840) <= a or b;
    layer0_outputs(3841) <= not (a or b);
    layer0_outputs(3842) <= a and not b;
    layer0_outputs(3843) <= not b;
    layer0_outputs(3844) <= b and not a;
    layer0_outputs(3845) <= not (a or b);
    layer0_outputs(3846) <= not (a or b);
    layer0_outputs(3847) <= not (a or b);
    layer0_outputs(3848) <= a and not b;
    layer0_outputs(3849) <= 1'b1;
    layer0_outputs(3850) <= not b;
    layer0_outputs(3851) <= not b;
    layer0_outputs(3852) <= not a;
    layer0_outputs(3853) <= a xor b;
    layer0_outputs(3854) <= not b;
    layer0_outputs(3855) <= b;
    layer0_outputs(3856) <= a;
    layer0_outputs(3857) <= a;
    layer0_outputs(3858) <= not (a or b);
    layer0_outputs(3859) <= not (a xor b);
    layer0_outputs(3860) <= not b;
    layer0_outputs(3861) <= a or b;
    layer0_outputs(3862) <= not b;
    layer0_outputs(3863) <= not (a xor b);
    layer0_outputs(3864) <= a;
    layer0_outputs(3865) <= not (a xor b);
    layer0_outputs(3866) <= a xor b;
    layer0_outputs(3867) <= not (a xor b);
    layer0_outputs(3868) <= not b;
    layer0_outputs(3869) <= not (a and b);
    layer0_outputs(3870) <= a and b;
    layer0_outputs(3871) <= not b;
    layer0_outputs(3872) <= a or b;
    layer0_outputs(3873) <= not (a or b);
    layer0_outputs(3874) <= not b;
    layer0_outputs(3875) <= 1'b1;
    layer0_outputs(3876) <= b and not a;
    layer0_outputs(3877) <= not (a or b);
    layer0_outputs(3878) <= not (a or b);
    layer0_outputs(3879) <= a and not b;
    layer0_outputs(3880) <= not b or a;
    layer0_outputs(3881) <= not a or b;
    layer0_outputs(3882) <= not (a xor b);
    layer0_outputs(3883) <= a and not b;
    layer0_outputs(3884) <= a or b;
    layer0_outputs(3885) <= not b;
    layer0_outputs(3886) <= not a or b;
    layer0_outputs(3887) <= a xor b;
    layer0_outputs(3888) <= not (a or b);
    layer0_outputs(3889) <= a or b;
    layer0_outputs(3890) <= not (a or b);
    layer0_outputs(3891) <= not (a or b);
    layer0_outputs(3892) <= not (a xor b);
    layer0_outputs(3893) <= not (a or b);
    layer0_outputs(3894) <= a xor b;
    layer0_outputs(3895) <= not a;
    layer0_outputs(3896) <= not b or a;
    layer0_outputs(3897) <= b and not a;
    layer0_outputs(3898) <= b and not a;
    layer0_outputs(3899) <= b;
    layer0_outputs(3900) <= not (a and b);
    layer0_outputs(3901) <= not a or b;
    layer0_outputs(3902) <= a and not b;
    layer0_outputs(3903) <= a;
    layer0_outputs(3904) <= not (a or b);
    layer0_outputs(3905) <= a and not b;
    layer0_outputs(3906) <= b;
    layer0_outputs(3907) <= not (a xor b);
    layer0_outputs(3908) <= not (a or b);
    layer0_outputs(3909) <= a and not b;
    layer0_outputs(3910) <= not (a or b);
    layer0_outputs(3911) <= a xor b;
    layer0_outputs(3912) <= not (a or b);
    layer0_outputs(3913) <= not (a xor b);
    layer0_outputs(3914) <= not a;
    layer0_outputs(3915) <= not (a or b);
    layer0_outputs(3916) <= b;
    layer0_outputs(3917) <= a and not b;
    layer0_outputs(3918) <= 1'b1;
    layer0_outputs(3919) <= b and not a;
    layer0_outputs(3920) <= not (a or b);
    layer0_outputs(3921) <= not a or b;
    layer0_outputs(3922) <= not (a xor b);
    layer0_outputs(3923) <= not (a or b);
    layer0_outputs(3924) <= not b or a;
    layer0_outputs(3925) <= b;
    layer0_outputs(3926) <= b and not a;
    layer0_outputs(3927) <= b and not a;
    layer0_outputs(3928) <= not (a or b);
    layer0_outputs(3929) <= not (a xor b);
    layer0_outputs(3930) <= not b or a;
    layer0_outputs(3931) <= not a;
    layer0_outputs(3932) <= not (a or b);
    layer0_outputs(3933) <= a and b;
    layer0_outputs(3934) <= not b or a;
    layer0_outputs(3935) <= a xor b;
    layer0_outputs(3936) <= a xor b;
    layer0_outputs(3937) <= not a or b;
    layer0_outputs(3938) <= a or b;
    layer0_outputs(3939) <= b and not a;
    layer0_outputs(3940) <= b;
    layer0_outputs(3941) <= a and not b;
    layer0_outputs(3942) <= a and b;
    layer0_outputs(3943) <= a or b;
    layer0_outputs(3944) <= a and not b;
    layer0_outputs(3945) <= not (a xor b);
    layer0_outputs(3946) <= b;
    layer0_outputs(3947) <= a or b;
    layer0_outputs(3948) <= not b;
    layer0_outputs(3949) <= a and not b;
    layer0_outputs(3950) <= a and not b;
    layer0_outputs(3951) <= a xor b;
    layer0_outputs(3952) <= a;
    layer0_outputs(3953) <= a xor b;
    layer0_outputs(3954) <= a xor b;
    layer0_outputs(3955) <= not (a xor b);
    layer0_outputs(3956) <= not b or a;
    layer0_outputs(3957) <= not a;
    layer0_outputs(3958) <= b;
    layer0_outputs(3959) <= b;
    layer0_outputs(3960) <= not a;
    layer0_outputs(3961) <= not b;
    layer0_outputs(3962) <= not (a or b);
    layer0_outputs(3963) <= not a;
    layer0_outputs(3964) <= not (a or b);
    layer0_outputs(3965) <= a xor b;
    layer0_outputs(3966) <= a and not b;
    layer0_outputs(3967) <= not a or b;
    layer0_outputs(3968) <= not a;
    layer0_outputs(3969) <= a xor b;
    layer0_outputs(3970) <= a or b;
    layer0_outputs(3971) <= a xor b;
    layer0_outputs(3972) <= a or b;
    layer0_outputs(3973) <= not a;
    layer0_outputs(3974) <= a and not b;
    layer0_outputs(3975) <= a and not b;
    layer0_outputs(3976) <= a or b;
    layer0_outputs(3977) <= not (a xor b);
    layer0_outputs(3978) <= not a;
    layer0_outputs(3979) <= b and not a;
    layer0_outputs(3980) <= not b;
    layer0_outputs(3981) <= not (a xor b);
    layer0_outputs(3982) <= a or b;
    layer0_outputs(3983) <= a and b;
    layer0_outputs(3984) <= not b;
    layer0_outputs(3985) <= not a or b;
    layer0_outputs(3986) <= a xor b;
    layer0_outputs(3987) <= not (a xor b);
    layer0_outputs(3988) <= not (a or b);
    layer0_outputs(3989) <= not b;
    layer0_outputs(3990) <= not (a or b);
    layer0_outputs(3991) <= not (a or b);
    layer0_outputs(3992) <= a;
    layer0_outputs(3993) <= not (a or b);
    layer0_outputs(3994) <= a and not b;
    layer0_outputs(3995) <= not a;
    layer0_outputs(3996) <= a;
    layer0_outputs(3997) <= not (a or b);
    layer0_outputs(3998) <= not (a or b);
    layer0_outputs(3999) <= not a;
    layer0_outputs(4000) <= b;
    layer0_outputs(4001) <= not (a xor b);
    layer0_outputs(4002) <= not (a xor b);
    layer0_outputs(4003) <= not b;
    layer0_outputs(4004) <= not (a or b);
    layer0_outputs(4005) <= a or b;
    layer0_outputs(4006) <= a xor b;
    layer0_outputs(4007) <= not a;
    layer0_outputs(4008) <= not (a and b);
    layer0_outputs(4009) <= not (a and b);
    layer0_outputs(4010) <= a xor b;
    layer0_outputs(4011) <= a and not b;
    layer0_outputs(4012) <= a xor b;
    layer0_outputs(4013) <= b and not a;
    layer0_outputs(4014) <= not b;
    layer0_outputs(4015) <= a xor b;
    layer0_outputs(4016) <= a or b;
    layer0_outputs(4017) <= a and b;
    layer0_outputs(4018) <= not a or b;
    layer0_outputs(4019) <= 1'b0;
    layer0_outputs(4020) <= not (a or b);
    layer0_outputs(4021) <= not (a or b);
    layer0_outputs(4022) <= not (a or b);
    layer0_outputs(4023) <= not a;
    layer0_outputs(4024) <= not (a or b);
    layer0_outputs(4025) <= a;
    layer0_outputs(4026) <= a and b;
    layer0_outputs(4027) <= b;
    layer0_outputs(4028) <= a or b;
    layer0_outputs(4029) <= a and not b;
    layer0_outputs(4030) <= not (a xor b);
    layer0_outputs(4031) <= not (a xor b);
    layer0_outputs(4032) <= a;
    layer0_outputs(4033) <= not (a xor b);
    layer0_outputs(4034) <= a and b;
    layer0_outputs(4035) <= not (a or b);
    layer0_outputs(4036) <= not (a or b);
    layer0_outputs(4037) <= a;
    layer0_outputs(4038) <= not a or b;
    layer0_outputs(4039) <= a;
    layer0_outputs(4040) <= not a;
    layer0_outputs(4041) <= not (a or b);
    layer0_outputs(4042) <= a or b;
    layer0_outputs(4043) <= not a;
    layer0_outputs(4044) <= not a;
    layer0_outputs(4045) <= a xor b;
    layer0_outputs(4046) <= 1'b0;
    layer0_outputs(4047) <= not (a or b);
    layer0_outputs(4048) <= not (a or b);
    layer0_outputs(4049) <= a and b;
    layer0_outputs(4050) <= not (a xor b);
    layer0_outputs(4051) <= not (a xor b);
    layer0_outputs(4052) <= a xor b;
    layer0_outputs(4053) <= not a or b;
    layer0_outputs(4054) <= not (a or b);
    layer0_outputs(4055) <= a or b;
    layer0_outputs(4056) <= not (a xor b);
    layer0_outputs(4057) <= not (a or b);
    layer0_outputs(4058) <= not b or a;
    layer0_outputs(4059) <= 1'b0;
    layer0_outputs(4060) <= not (a or b);
    layer0_outputs(4061) <= a;
    layer0_outputs(4062) <= 1'b1;
    layer0_outputs(4063) <= not a;
    layer0_outputs(4064) <= 1'b0;
    layer0_outputs(4065) <= b;
    layer0_outputs(4066) <= not a;
    layer0_outputs(4067) <= a or b;
    layer0_outputs(4068) <= a;
    layer0_outputs(4069) <= not b or a;
    layer0_outputs(4070) <= not (a xor b);
    layer0_outputs(4071) <= not b or a;
    layer0_outputs(4072) <= not a;
    layer0_outputs(4073) <= not (a xor b);
    layer0_outputs(4074) <= a or b;
    layer0_outputs(4075) <= b and not a;
    layer0_outputs(4076) <= a and not b;
    layer0_outputs(4077) <= a xor b;
    layer0_outputs(4078) <= b;
    layer0_outputs(4079) <= a xor b;
    layer0_outputs(4080) <= not b;
    layer0_outputs(4081) <= a or b;
    layer0_outputs(4082) <= not b;
    layer0_outputs(4083) <= not a;
    layer0_outputs(4084) <= not a or b;
    layer0_outputs(4085) <= not (a xor b);
    layer0_outputs(4086) <= a;
    layer0_outputs(4087) <= not a;
    layer0_outputs(4088) <= not (a or b);
    layer0_outputs(4089) <= a or b;
    layer0_outputs(4090) <= not b;
    layer0_outputs(4091) <= a or b;
    layer0_outputs(4092) <= a and not b;
    layer0_outputs(4093) <= not (a xor b);
    layer0_outputs(4094) <= a or b;
    layer0_outputs(4095) <= 1'b0;
    layer0_outputs(4096) <= not a;
    layer0_outputs(4097) <= a xor b;
    layer0_outputs(4098) <= a and b;
    layer0_outputs(4099) <= not a or b;
    layer0_outputs(4100) <= not a or b;
    layer0_outputs(4101) <= not b or a;
    layer0_outputs(4102) <= not (a or b);
    layer0_outputs(4103) <= a or b;
    layer0_outputs(4104) <= not b or a;
    layer0_outputs(4105) <= a and not b;
    layer0_outputs(4106) <= not (a or b);
    layer0_outputs(4107) <= a and not b;
    layer0_outputs(4108) <= not (a xor b);
    layer0_outputs(4109) <= 1'b1;
    layer0_outputs(4110) <= not (a xor b);
    layer0_outputs(4111) <= not (a or b);
    layer0_outputs(4112) <= a or b;
    layer0_outputs(4113) <= not b;
    layer0_outputs(4114) <= a and b;
    layer0_outputs(4115) <= not (a or b);
    layer0_outputs(4116) <= not a or b;
    layer0_outputs(4117) <= a and not b;
    layer0_outputs(4118) <= not (a xor b);
    layer0_outputs(4119) <= not b or a;
    layer0_outputs(4120) <= not a;
    layer0_outputs(4121) <= b;
    layer0_outputs(4122) <= not a;
    layer0_outputs(4123) <= not (a xor b);
    layer0_outputs(4124) <= not a or b;
    layer0_outputs(4125) <= 1'b1;
    layer0_outputs(4126) <= b;
    layer0_outputs(4127) <= b and not a;
    layer0_outputs(4128) <= not (a or b);
    layer0_outputs(4129) <= a;
    layer0_outputs(4130) <= b and not a;
    layer0_outputs(4131) <= a or b;
    layer0_outputs(4132) <= b and not a;
    layer0_outputs(4133) <= not (a xor b);
    layer0_outputs(4134) <= not a;
    layer0_outputs(4135) <= a and not b;
    layer0_outputs(4136) <= not a or b;
    layer0_outputs(4137) <= not a or b;
    layer0_outputs(4138) <= a or b;
    layer0_outputs(4139) <= not a or b;
    layer0_outputs(4140) <= not (a xor b);
    layer0_outputs(4141) <= not b;
    layer0_outputs(4142) <= a or b;
    layer0_outputs(4143) <= a and b;
    layer0_outputs(4144) <= not (a or b);
    layer0_outputs(4145) <= not (a or b);
    layer0_outputs(4146) <= 1'b0;
    layer0_outputs(4147) <= a or b;
    layer0_outputs(4148) <= b;
    layer0_outputs(4149) <= not (a xor b);
    layer0_outputs(4150) <= not a or b;
    layer0_outputs(4151) <= a or b;
    layer0_outputs(4152) <= not (a and b);
    layer0_outputs(4153) <= b and not a;
    layer0_outputs(4154) <= not (a xor b);
    layer0_outputs(4155) <= not b;
    layer0_outputs(4156) <= b and not a;
    layer0_outputs(4157) <= not a or b;
    layer0_outputs(4158) <= not (a or b);
    layer0_outputs(4159) <= b and not a;
    layer0_outputs(4160) <= not b;
    layer0_outputs(4161) <= a xor b;
    layer0_outputs(4162) <= not b;
    layer0_outputs(4163) <= 1'b1;
    layer0_outputs(4164) <= 1'b0;
    layer0_outputs(4165) <= not b;
    layer0_outputs(4166) <= a or b;
    layer0_outputs(4167) <= b;
    layer0_outputs(4168) <= not a or b;
    layer0_outputs(4169) <= not b or a;
    layer0_outputs(4170) <= a or b;
    layer0_outputs(4171) <= a xor b;
    layer0_outputs(4172) <= 1'b0;
    layer0_outputs(4173) <= a or b;
    layer0_outputs(4174) <= not b or a;
    layer0_outputs(4175) <= not b or a;
    layer0_outputs(4176) <= a;
    layer0_outputs(4177) <= a or b;
    layer0_outputs(4178) <= a or b;
    layer0_outputs(4179) <= a and not b;
    layer0_outputs(4180) <= a or b;
    layer0_outputs(4181) <= a xor b;
    layer0_outputs(4182) <= not b or a;
    layer0_outputs(4183) <= a and not b;
    layer0_outputs(4184) <= 1'b0;
    layer0_outputs(4185) <= a or b;
    layer0_outputs(4186) <= not a or b;
    layer0_outputs(4187) <= not b;
    layer0_outputs(4188) <= not a;
    layer0_outputs(4189) <= not b;
    layer0_outputs(4190) <= not a;
    layer0_outputs(4191) <= b and not a;
    layer0_outputs(4192) <= b and not a;
    layer0_outputs(4193) <= 1'b0;
    layer0_outputs(4194) <= a and not b;
    layer0_outputs(4195) <= not a;
    layer0_outputs(4196) <= not (a or b);
    layer0_outputs(4197) <= not (a and b);
    layer0_outputs(4198) <= not a or b;
    layer0_outputs(4199) <= not (a or b);
    layer0_outputs(4200) <= not (a and b);
    layer0_outputs(4201) <= not a or b;
    layer0_outputs(4202) <= a;
    layer0_outputs(4203) <= b;
    layer0_outputs(4204) <= a xor b;
    layer0_outputs(4205) <= a and b;
    layer0_outputs(4206) <= not a or b;
    layer0_outputs(4207) <= not (a or b);
    layer0_outputs(4208) <= b and not a;
    layer0_outputs(4209) <= not b;
    layer0_outputs(4210) <= 1'b0;
    layer0_outputs(4211) <= not b or a;
    layer0_outputs(4212) <= not a or b;
    layer0_outputs(4213) <= not a;
    layer0_outputs(4214) <= a;
    layer0_outputs(4215) <= not a;
    layer0_outputs(4216) <= a or b;
    layer0_outputs(4217) <= a or b;
    layer0_outputs(4218) <= not (a xor b);
    layer0_outputs(4219) <= not a;
    layer0_outputs(4220) <= not (a or b);
    layer0_outputs(4221) <= a and b;
    layer0_outputs(4222) <= a and not b;
    layer0_outputs(4223) <= not b;
    layer0_outputs(4224) <= not (a or b);
    layer0_outputs(4225) <= not (a xor b);
    layer0_outputs(4226) <= 1'b1;
    layer0_outputs(4227) <= b;
    layer0_outputs(4228) <= a or b;
    layer0_outputs(4229) <= not (a or b);
    layer0_outputs(4230) <= a xor b;
    layer0_outputs(4231) <= b and not a;
    layer0_outputs(4232) <= not (a or b);
    layer0_outputs(4233) <= a;
    layer0_outputs(4234) <= a or b;
    layer0_outputs(4235) <= not (a or b);
    layer0_outputs(4236) <= not (a or b);
    layer0_outputs(4237) <= a;
    layer0_outputs(4238) <= a and b;
    layer0_outputs(4239) <= b;
    layer0_outputs(4240) <= b;
    layer0_outputs(4241) <= b and not a;
    layer0_outputs(4242) <= not b;
    layer0_outputs(4243) <= not (a xor b);
    layer0_outputs(4244) <= not b;
    layer0_outputs(4245) <= not (a or b);
    layer0_outputs(4246) <= not a or b;
    layer0_outputs(4247) <= a;
    layer0_outputs(4248) <= a or b;
    layer0_outputs(4249) <= b;
    layer0_outputs(4250) <= not b;
    layer0_outputs(4251) <= a and not b;
    layer0_outputs(4252) <= a or b;
    layer0_outputs(4253) <= not a;
    layer0_outputs(4254) <= not a;
    layer0_outputs(4255) <= not a;
    layer0_outputs(4256) <= not (a xor b);
    layer0_outputs(4257) <= a or b;
    layer0_outputs(4258) <= b and not a;
    layer0_outputs(4259) <= a xor b;
    layer0_outputs(4260) <= not a;
    layer0_outputs(4261) <= a or b;
    layer0_outputs(4262) <= a and not b;
    layer0_outputs(4263) <= a and b;
    layer0_outputs(4264) <= not a;
    layer0_outputs(4265) <= not a;
    layer0_outputs(4266) <= not a or b;
    layer0_outputs(4267) <= not a;
    layer0_outputs(4268) <= a and b;
    layer0_outputs(4269) <= not b or a;
    layer0_outputs(4270) <= a;
    layer0_outputs(4271) <= a or b;
    layer0_outputs(4272) <= not a or b;
    layer0_outputs(4273) <= a xor b;
    layer0_outputs(4274) <= a or b;
    layer0_outputs(4275) <= not a or b;
    layer0_outputs(4276) <= not b or a;
    layer0_outputs(4277) <= not (a or b);
    layer0_outputs(4278) <= 1'b1;
    layer0_outputs(4279) <= a xor b;
    layer0_outputs(4280) <= 1'b0;
    layer0_outputs(4281) <= a or b;
    layer0_outputs(4282) <= not b or a;
    layer0_outputs(4283) <= not b;
    layer0_outputs(4284) <= b;
    layer0_outputs(4285) <= not (a xor b);
    layer0_outputs(4286) <= b and not a;
    layer0_outputs(4287) <= not a;
    layer0_outputs(4288) <= not (a xor b);
    layer0_outputs(4289) <= b and not a;
    layer0_outputs(4290) <= not (a xor b);
    layer0_outputs(4291) <= not a or b;
    layer0_outputs(4292) <= not a;
    layer0_outputs(4293) <= not a or b;
    layer0_outputs(4294) <= not (a xor b);
    layer0_outputs(4295) <= a xor b;
    layer0_outputs(4296) <= a and not b;
    layer0_outputs(4297) <= b and not a;
    layer0_outputs(4298) <= a and not b;
    layer0_outputs(4299) <= a xor b;
    layer0_outputs(4300) <= not b or a;
    layer0_outputs(4301) <= a or b;
    layer0_outputs(4302) <= not (a or b);
    layer0_outputs(4303) <= b and not a;
    layer0_outputs(4304) <= not a or b;
    layer0_outputs(4305) <= not a;
    layer0_outputs(4306) <= not (a xor b);
    layer0_outputs(4307) <= a and b;
    layer0_outputs(4308) <= not a;
    layer0_outputs(4309) <= 1'b1;
    layer0_outputs(4310) <= not (a or b);
    layer0_outputs(4311) <= a;
    layer0_outputs(4312) <= b and not a;
    layer0_outputs(4313) <= b and not a;
    layer0_outputs(4314) <= a;
    layer0_outputs(4315) <= not (a or b);
    layer0_outputs(4316) <= a xor b;
    layer0_outputs(4317) <= not b;
    layer0_outputs(4318) <= a or b;
    layer0_outputs(4319) <= b;
    layer0_outputs(4320) <= not (a or b);
    layer0_outputs(4321) <= not a;
    layer0_outputs(4322) <= a or b;
    layer0_outputs(4323) <= b;
    layer0_outputs(4324) <= a xor b;
    layer0_outputs(4325) <= not (a or b);
    layer0_outputs(4326) <= a and not b;
    layer0_outputs(4327) <= a xor b;
    layer0_outputs(4328) <= a xor b;
    layer0_outputs(4329) <= a;
    layer0_outputs(4330) <= not (a or b);
    layer0_outputs(4331) <= not (a or b);
    layer0_outputs(4332) <= a xor b;
    layer0_outputs(4333) <= not a or b;
    layer0_outputs(4334) <= 1'b1;
    layer0_outputs(4335) <= a or b;
    layer0_outputs(4336) <= not (a or b);
    layer0_outputs(4337) <= not (a and b);
    layer0_outputs(4338) <= not (a or b);
    layer0_outputs(4339) <= not (a xor b);
    layer0_outputs(4340) <= not (a and b);
    layer0_outputs(4341) <= not (a xor b);
    layer0_outputs(4342) <= not (a and b);
    layer0_outputs(4343) <= not b;
    layer0_outputs(4344) <= not b or a;
    layer0_outputs(4345) <= not b or a;
    layer0_outputs(4346) <= not (a xor b);
    layer0_outputs(4347) <= not b;
    layer0_outputs(4348) <= a xor b;
    layer0_outputs(4349) <= 1'b0;
    layer0_outputs(4350) <= not a;
    layer0_outputs(4351) <= a and b;
    layer0_outputs(4352) <= not a or b;
    layer0_outputs(4353) <= not (a xor b);
    layer0_outputs(4354) <= a and b;
    layer0_outputs(4355) <= a xor b;
    layer0_outputs(4356) <= not a;
    layer0_outputs(4357) <= a xor b;
    layer0_outputs(4358) <= not a;
    layer0_outputs(4359) <= b and not a;
    layer0_outputs(4360) <= b;
    layer0_outputs(4361) <= not (a xor b);
    layer0_outputs(4362) <= a and b;
    layer0_outputs(4363) <= b;
    layer0_outputs(4364) <= not (a xor b);
    layer0_outputs(4365) <= not a or b;
    layer0_outputs(4366) <= not (a or b);
    layer0_outputs(4367) <= a and not b;
    layer0_outputs(4368) <= b and not a;
    layer0_outputs(4369) <= not a or b;
    layer0_outputs(4370) <= 1'b0;
    layer0_outputs(4371) <= b and not a;
    layer0_outputs(4372) <= not (a or b);
    layer0_outputs(4373) <= a xor b;
    layer0_outputs(4374) <= a or b;
    layer0_outputs(4375) <= not a;
    layer0_outputs(4376) <= not (a or b);
    layer0_outputs(4377) <= a or b;
    layer0_outputs(4378) <= not (a xor b);
    layer0_outputs(4379) <= b and not a;
    layer0_outputs(4380) <= 1'b0;
    layer0_outputs(4381) <= a or b;
    layer0_outputs(4382) <= b and not a;
    layer0_outputs(4383) <= a and not b;
    layer0_outputs(4384) <= a xor b;
    layer0_outputs(4385) <= not b or a;
    layer0_outputs(4386) <= a xor b;
    layer0_outputs(4387) <= a and not b;
    layer0_outputs(4388) <= a and not b;
    layer0_outputs(4389) <= not a or b;
    layer0_outputs(4390) <= not (a xor b);
    layer0_outputs(4391) <= not (a xor b);
    layer0_outputs(4392) <= a xor b;
    layer0_outputs(4393) <= not b or a;
    layer0_outputs(4394) <= a or b;
    layer0_outputs(4395) <= b;
    layer0_outputs(4396) <= not a;
    layer0_outputs(4397) <= a;
    layer0_outputs(4398) <= not b;
    layer0_outputs(4399) <= not (a or b);
    layer0_outputs(4400) <= a;
    layer0_outputs(4401) <= not b;
    layer0_outputs(4402) <= not a;
    layer0_outputs(4403) <= a or b;
    layer0_outputs(4404) <= not b or a;
    layer0_outputs(4405) <= not a;
    layer0_outputs(4406) <= a and b;
    layer0_outputs(4407) <= b and not a;
    layer0_outputs(4408) <= not (a xor b);
    layer0_outputs(4409) <= not a;
    layer0_outputs(4410) <= 1'b0;
    layer0_outputs(4411) <= b;
    layer0_outputs(4412) <= a or b;
    layer0_outputs(4413) <= a xor b;
    layer0_outputs(4414) <= not (a xor b);
    layer0_outputs(4415) <= a;
    layer0_outputs(4416) <= a and not b;
    layer0_outputs(4417) <= not a;
    layer0_outputs(4418) <= a;
    layer0_outputs(4419) <= a or b;
    layer0_outputs(4420) <= not (a or b);
    layer0_outputs(4421) <= a xor b;
    layer0_outputs(4422) <= not (a xor b);
    layer0_outputs(4423) <= a xor b;
    layer0_outputs(4424) <= a;
    layer0_outputs(4425) <= b and not a;
    layer0_outputs(4426) <= not (a or b);
    layer0_outputs(4427) <= not (a or b);
    layer0_outputs(4428) <= b and not a;
    layer0_outputs(4429) <= b and not a;
    layer0_outputs(4430) <= not (a xor b);
    layer0_outputs(4431) <= 1'b1;
    layer0_outputs(4432) <= a;
    layer0_outputs(4433) <= not a or b;
    layer0_outputs(4434) <= not b;
    layer0_outputs(4435) <= b and not a;
    layer0_outputs(4436) <= a or b;
    layer0_outputs(4437) <= not (a or b);
    layer0_outputs(4438) <= not (a or b);
    layer0_outputs(4439) <= not (a xor b);
    layer0_outputs(4440) <= b;
    layer0_outputs(4441) <= not b or a;
    layer0_outputs(4442) <= a or b;
    layer0_outputs(4443) <= not a;
    layer0_outputs(4444) <= a;
    layer0_outputs(4445) <= a or b;
    layer0_outputs(4446) <= a xor b;
    layer0_outputs(4447) <= a or b;
    layer0_outputs(4448) <= a;
    layer0_outputs(4449) <= b;
    layer0_outputs(4450) <= a xor b;
    layer0_outputs(4451) <= not (a or b);
    layer0_outputs(4452) <= b and not a;
    layer0_outputs(4453) <= a xor b;
    layer0_outputs(4454) <= a or b;
    layer0_outputs(4455) <= a xor b;
    layer0_outputs(4456) <= a xor b;
    layer0_outputs(4457) <= not (a xor b);
    layer0_outputs(4458) <= a and not b;
    layer0_outputs(4459) <= b;
    layer0_outputs(4460) <= a and not b;
    layer0_outputs(4461) <= a or b;
    layer0_outputs(4462) <= a and b;
    layer0_outputs(4463) <= b and not a;
    layer0_outputs(4464) <= not (a or b);
    layer0_outputs(4465) <= b;
    layer0_outputs(4466) <= not a;
    layer0_outputs(4467) <= not (a xor b);
    layer0_outputs(4468) <= not a or b;
    layer0_outputs(4469) <= a and not b;
    layer0_outputs(4470) <= a;
    layer0_outputs(4471) <= 1'b1;
    layer0_outputs(4472) <= a xor b;
    layer0_outputs(4473) <= not (a or b);
    layer0_outputs(4474) <= a;
    layer0_outputs(4475) <= not (a xor b);
    layer0_outputs(4476) <= a or b;
    layer0_outputs(4477) <= a;
    layer0_outputs(4478) <= a and not b;
    layer0_outputs(4479) <= not b or a;
    layer0_outputs(4480) <= a xor b;
    layer0_outputs(4481) <= b and not a;
    layer0_outputs(4482) <= not b;
    layer0_outputs(4483) <= not (a or b);
    layer0_outputs(4484) <= not a or b;
    layer0_outputs(4485) <= not (a or b);
    layer0_outputs(4486) <= a xor b;
    layer0_outputs(4487) <= a and not b;
    layer0_outputs(4488) <= a and not b;
    layer0_outputs(4489) <= b;
    layer0_outputs(4490) <= a and not b;
    layer0_outputs(4491) <= a or b;
    layer0_outputs(4492) <= b and not a;
    layer0_outputs(4493) <= not (a or b);
    layer0_outputs(4494) <= not b;
    layer0_outputs(4495) <= not (a or b);
    layer0_outputs(4496) <= not (a or b);
    layer0_outputs(4497) <= b;
    layer0_outputs(4498) <= a xor b;
    layer0_outputs(4499) <= a;
    layer0_outputs(4500) <= a;
    layer0_outputs(4501) <= not (a xor b);
    layer0_outputs(4502) <= not b;
    layer0_outputs(4503) <= not b or a;
    layer0_outputs(4504) <= a or b;
    layer0_outputs(4505) <= a;
    layer0_outputs(4506) <= b and not a;
    layer0_outputs(4507) <= not b;
    layer0_outputs(4508) <= not (a xor b);
    layer0_outputs(4509) <= not (a xor b);
    layer0_outputs(4510) <= not a;
    layer0_outputs(4511) <= not (a xor b);
    layer0_outputs(4512) <= not (a xor b);
    layer0_outputs(4513) <= not (a xor b);
    layer0_outputs(4514) <= not b or a;
    layer0_outputs(4515) <= not a;
    layer0_outputs(4516) <= 1'b0;
    layer0_outputs(4517) <= not (a and b);
    layer0_outputs(4518) <= not (a or b);
    layer0_outputs(4519) <= not (a or b);
    layer0_outputs(4520) <= not a;
    layer0_outputs(4521) <= b;
    layer0_outputs(4522) <= b and not a;
    layer0_outputs(4523) <= a and not b;
    layer0_outputs(4524) <= b;
    layer0_outputs(4525) <= a xor b;
    layer0_outputs(4526) <= a or b;
    layer0_outputs(4527) <= a and b;
    layer0_outputs(4528) <= a and not b;
    layer0_outputs(4529) <= a xor b;
    layer0_outputs(4530) <= a or b;
    layer0_outputs(4531) <= a or b;
    layer0_outputs(4532) <= b;
    layer0_outputs(4533) <= not (a or b);
    layer0_outputs(4534) <= b;
    layer0_outputs(4535) <= a xor b;
    layer0_outputs(4536) <= not a or b;
    layer0_outputs(4537) <= not (a or b);
    layer0_outputs(4538) <= not (a or b);
    layer0_outputs(4539) <= not b or a;
    layer0_outputs(4540) <= not (a or b);
    layer0_outputs(4541) <= not (a or b);
    layer0_outputs(4542) <= b;
    layer0_outputs(4543) <= not b;
    layer0_outputs(4544) <= not (a xor b);
    layer0_outputs(4545) <= b and not a;
    layer0_outputs(4546) <= not b;
    layer0_outputs(4547) <= a xor b;
    layer0_outputs(4548) <= a or b;
    layer0_outputs(4549) <= not b or a;
    layer0_outputs(4550) <= not b;
    layer0_outputs(4551) <= not b;
    layer0_outputs(4552) <= a;
    layer0_outputs(4553) <= not b;
    layer0_outputs(4554) <= not (a or b);
    layer0_outputs(4555) <= a and not b;
    layer0_outputs(4556) <= a;
    layer0_outputs(4557) <= not a;
    layer0_outputs(4558) <= a and not b;
    layer0_outputs(4559) <= not b or a;
    layer0_outputs(4560) <= a or b;
    layer0_outputs(4561) <= a and not b;
    layer0_outputs(4562) <= a or b;
    layer0_outputs(4563) <= not (a xor b);
    layer0_outputs(4564) <= 1'b1;
    layer0_outputs(4565) <= not (a or b);
    layer0_outputs(4566) <= b;
    layer0_outputs(4567) <= a or b;
    layer0_outputs(4568) <= not a or b;
    layer0_outputs(4569) <= a or b;
    layer0_outputs(4570) <= not b or a;
    layer0_outputs(4571) <= a or b;
    layer0_outputs(4572) <= a;
    layer0_outputs(4573) <= not (a xor b);
    layer0_outputs(4574) <= not (a or b);
    layer0_outputs(4575) <= a;
    layer0_outputs(4576) <= b and not a;
    layer0_outputs(4577) <= not b or a;
    layer0_outputs(4578) <= not a or b;
    layer0_outputs(4579) <= not b or a;
    layer0_outputs(4580) <= b and not a;
    layer0_outputs(4581) <= b and not a;
    layer0_outputs(4582) <= not b;
    layer0_outputs(4583) <= a xor b;
    layer0_outputs(4584) <= not a;
    layer0_outputs(4585) <= a;
    layer0_outputs(4586) <= a and not b;
    layer0_outputs(4587) <= not b;
    layer0_outputs(4588) <= a;
    layer0_outputs(4589) <= not (a xor b);
    layer0_outputs(4590) <= a and not b;
    layer0_outputs(4591) <= a xor b;
    layer0_outputs(4592) <= not a or b;
    layer0_outputs(4593) <= not a;
    layer0_outputs(4594) <= a;
    layer0_outputs(4595) <= 1'b1;
    layer0_outputs(4596) <= not b or a;
    layer0_outputs(4597) <= not b;
    layer0_outputs(4598) <= 1'b1;
    layer0_outputs(4599) <= not a;
    layer0_outputs(4600) <= not b;
    layer0_outputs(4601) <= a xor b;
    layer0_outputs(4602) <= b and not a;
    layer0_outputs(4603) <= not a or b;
    layer0_outputs(4604) <= a;
    layer0_outputs(4605) <= not (a xor b);
    layer0_outputs(4606) <= b;
    layer0_outputs(4607) <= b;
    layer0_outputs(4608) <= not (a or b);
    layer0_outputs(4609) <= not (a xor b);
    layer0_outputs(4610) <= not a;
    layer0_outputs(4611) <= a or b;
    layer0_outputs(4612) <= b and not a;
    layer0_outputs(4613) <= b;
    layer0_outputs(4614) <= a xor b;
    layer0_outputs(4615) <= a xor b;
    layer0_outputs(4616) <= a and not b;
    layer0_outputs(4617) <= 1'b1;
    layer0_outputs(4618) <= not (a xor b);
    layer0_outputs(4619) <= a or b;
    layer0_outputs(4620) <= not a or b;
    layer0_outputs(4621) <= b;
    layer0_outputs(4622) <= b;
    layer0_outputs(4623) <= not (a xor b);
    layer0_outputs(4624) <= b;
    layer0_outputs(4625) <= not (a or b);
    layer0_outputs(4626) <= a xor b;
    layer0_outputs(4627) <= a or b;
    layer0_outputs(4628) <= not (a xor b);
    layer0_outputs(4629) <= a;
    layer0_outputs(4630) <= not b or a;
    layer0_outputs(4631) <= not (a and b);
    layer0_outputs(4632) <= a or b;
    layer0_outputs(4633) <= not (a or b);
    layer0_outputs(4634) <= not (a xor b);
    layer0_outputs(4635) <= not (a or b);
    layer0_outputs(4636) <= a or b;
    layer0_outputs(4637) <= b and not a;
    layer0_outputs(4638) <= not (a xor b);
    layer0_outputs(4639) <= not (a xor b);
    layer0_outputs(4640) <= not (a xor b);
    layer0_outputs(4641) <= a xor b;
    layer0_outputs(4642) <= a or b;
    layer0_outputs(4643) <= not (a xor b);
    layer0_outputs(4644) <= not a or b;
    layer0_outputs(4645) <= a;
    layer0_outputs(4646) <= a;
    layer0_outputs(4647) <= a;
    layer0_outputs(4648) <= a or b;
    layer0_outputs(4649) <= not (a xor b);
    layer0_outputs(4650) <= a xor b;
    layer0_outputs(4651) <= not a or b;
    layer0_outputs(4652) <= not b;
    layer0_outputs(4653) <= not a or b;
    layer0_outputs(4654) <= not a or b;
    layer0_outputs(4655) <= not (a or b);
    layer0_outputs(4656) <= 1'b1;
    layer0_outputs(4657) <= a or b;
    layer0_outputs(4658) <= a or b;
    layer0_outputs(4659) <= not b or a;
    layer0_outputs(4660) <= not a;
    layer0_outputs(4661) <= not (a xor b);
    layer0_outputs(4662) <= not a or b;
    layer0_outputs(4663) <= a or b;
    layer0_outputs(4664) <= not b;
    layer0_outputs(4665) <= a xor b;
    layer0_outputs(4666) <= b;
    layer0_outputs(4667) <= not (a xor b);
    layer0_outputs(4668) <= not (a or b);
    layer0_outputs(4669) <= not a or b;
    layer0_outputs(4670) <= not b or a;
    layer0_outputs(4671) <= b and not a;
    layer0_outputs(4672) <= not b or a;
    layer0_outputs(4673) <= not a;
    layer0_outputs(4674) <= not (a xor b);
    layer0_outputs(4675) <= 1'b0;
    layer0_outputs(4676) <= not b;
    layer0_outputs(4677) <= 1'b0;
    layer0_outputs(4678) <= not (a xor b);
    layer0_outputs(4679) <= not a;
    layer0_outputs(4680) <= not (a xor b);
    layer0_outputs(4681) <= a;
    layer0_outputs(4682) <= a and b;
    layer0_outputs(4683) <= not b or a;
    layer0_outputs(4684) <= not (a xor b);
    layer0_outputs(4685) <= not b;
    layer0_outputs(4686) <= not (a xor b);
    layer0_outputs(4687) <= a and not b;
    layer0_outputs(4688) <= a;
    layer0_outputs(4689) <= a or b;
    layer0_outputs(4690) <= not (a or b);
    layer0_outputs(4691) <= not a;
    layer0_outputs(4692) <= b and not a;
    layer0_outputs(4693) <= a;
    layer0_outputs(4694) <= a and not b;
    layer0_outputs(4695) <= not b or a;
    layer0_outputs(4696) <= not (a and b);
    layer0_outputs(4697) <= b and not a;
    layer0_outputs(4698) <= not b or a;
    layer0_outputs(4699) <= a xor b;
    layer0_outputs(4700) <= not b or a;
    layer0_outputs(4701) <= b;
    layer0_outputs(4702) <= a or b;
    layer0_outputs(4703) <= 1'b0;
    layer0_outputs(4704) <= a or b;
    layer0_outputs(4705) <= not a or b;
    layer0_outputs(4706) <= not b;
    layer0_outputs(4707) <= not (a or b);
    layer0_outputs(4708) <= not a or b;
    layer0_outputs(4709) <= not (a or b);
    layer0_outputs(4710) <= a or b;
    layer0_outputs(4711) <= not a or b;
    layer0_outputs(4712) <= not (a xor b);
    layer0_outputs(4713) <= a xor b;
    layer0_outputs(4714) <= not (a xor b);
    layer0_outputs(4715) <= not a;
    layer0_outputs(4716) <= a xor b;
    layer0_outputs(4717) <= not (a xor b);
    layer0_outputs(4718) <= not (a or b);
    layer0_outputs(4719) <= not (a or b);
    layer0_outputs(4720) <= not b;
    layer0_outputs(4721) <= a and not b;
    layer0_outputs(4722) <= a or b;
    layer0_outputs(4723) <= not b;
    layer0_outputs(4724) <= a;
    layer0_outputs(4725) <= b and not a;
    layer0_outputs(4726) <= a or b;
    layer0_outputs(4727) <= b and not a;
    layer0_outputs(4728) <= not a;
    layer0_outputs(4729) <= a or b;
    layer0_outputs(4730) <= b;
    layer0_outputs(4731) <= 1'b0;
    layer0_outputs(4732) <= not (a xor b);
    layer0_outputs(4733) <= a or b;
    layer0_outputs(4734) <= not (a or b);
    layer0_outputs(4735) <= a xor b;
    layer0_outputs(4736) <= a;
    layer0_outputs(4737) <= a xor b;
    layer0_outputs(4738) <= not b or a;
    layer0_outputs(4739) <= a xor b;
    layer0_outputs(4740) <= a;
    layer0_outputs(4741) <= b and not a;
    layer0_outputs(4742) <= not a;
    layer0_outputs(4743) <= a;
    layer0_outputs(4744) <= not a or b;
    layer0_outputs(4745) <= a xor b;
    layer0_outputs(4746) <= not (a xor b);
    layer0_outputs(4747) <= not b;
    layer0_outputs(4748) <= not a;
    layer0_outputs(4749) <= b;
    layer0_outputs(4750) <= not a;
    layer0_outputs(4751) <= not b;
    layer0_outputs(4752) <= not a;
    layer0_outputs(4753) <= a or b;
    layer0_outputs(4754) <= b;
    layer0_outputs(4755) <= not (a or b);
    layer0_outputs(4756) <= not b;
    layer0_outputs(4757) <= not a;
    layer0_outputs(4758) <= not (a or b);
    layer0_outputs(4759) <= a xor b;
    layer0_outputs(4760) <= a or b;
    layer0_outputs(4761) <= not b;
    layer0_outputs(4762) <= a and not b;
    layer0_outputs(4763) <= not (a or b);
    layer0_outputs(4764) <= not (a xor b);
    layer0_outputs(4765) <= not a;
    layer0_outputs(4766) <= a;
    layer0_outputs(4767) <= not (a or b);
    layer0_outputs(4768) <= not (a xor b);
    layer0_outputs(4769) <= not a or b;
    layer0_outputs(4770) <= a or b;
    layer0_outputs(4771) <= not (a and b);
    layer0_outputs(4772) <= 1'b0;
    layer0_outputs(4773) <= not (a xor b);
    layer0_outputs(4774) <= a and not b;
    layer0_outputs(4775) <= b and not a;
    layer0_outputs(4776) <= b;
    layer0_outputs(4777) <= not (a or b);
    layer0_outputs(4778) <= a xor b;
    layer0_outputs(4779) <= not b;
    layer0_outputs(4780) <= a or b;
    layer0_outputs(4781) <= b;
    layer0_outputs(4782) <= not (a or b);
    layer0_outputs(4783) <= not (a xor b);
    layer0_outputs(4784) <= b;
    layer0_outputs(4785) <= a xor b;
    layer0_outputs(4786) <= not b or a;
    layer0_outputs(4787) <= not b or a;
    layer0_outputs(4788) <= not b or a;
    layer0_outputs(4789) <= a or b;
    layer0_outputs(4790) <= not (a xor b);
    layer0_outputs(4791) <= not (a or b);
    layer0_outputs(4792) <= a xor b;
    layer0_outputs(4793) <= b;
    layer0_outputs(4794) <= not (a xor b);
    layer0_outputs(4795) <= b;
    layer0_outputs(4796) <= a or b;
    layer0_outputs(4797) <= a xor b;
    layer0_outputs(4798) <= not (a xor b);
    layer0_outputs(4799) <= not b;
    layer0_outputs(4800) <= not a;
    layer0_outputs(4801) <= not (a or b);
    layer0_outputs(4802) <= not b or a;
    layer0_outputs(4803) <= 1'b0;
    layer0_outputs(4804) <= not (a or b);
    layer0_outputs(4805) <= a xor b;
    layer0_outputs(4806) <= a or b;
    layer0_outputs(4807) <= not b or a;
    layer0_outputs(4808) <= a;
    layer0_outputs(4809) <= a or b;
    layer0_outputs(4810) <= b;
    layer0_outputs(4811) <= a;
    layer0_outputs(4812) <= not b or a;
    layer0_outputs(4813) <= a or b;
    layer0_outputs(4814) <= b and not a;
    layer0_outputs(4815) <= not b;
    layer0_outputs(4816) <= not (a xor b);
    layer0_outputs(4817) <= a or b;
    layer0_outputs(4818) <= a and not b;
    layer0_outputs(4819) <= not (a xor b);
    layer0_outputs(4820) <= a;
    layer0_outputs(4821) <= not a;
    layer0_outputs(4822) <= not a;
    layer0_outputs(4823) <= not a;
    layer0_outputs(4824) <= a;
    layer0_outputs(4825) <= a and not b;
    layer0_outputs(4826) <= not (a or b);
    layer0_outputs(4827) <= a or b;
    layer0_outputs(4828) <= b and not a;
    layer0_outputs(4829) <= b;
    layer0_outputs(4830) <= not b;
    layer0_outputs(4831) <= a xor b;
    layer0_outputs(4832) <= 1'b1;
    layer0_outputs(4833) <= not (a or b);
    layer0_outputs(4834) <= a;
    layer0_outputs(4835) <= a;
    layer0_outputs(4836) <= a xor b;
    layer0_outputs(4837) <= not a;
    layer0_outputs(4838) <= b;
    layer0_outputs(4839) <= 1'b1;
    layer0_outputs(4840) <= a or b;
    layer0_outputs(4841) <= a and not b;
    layer0_outputs(4842) <= a and not b;
    layer0_outputs(4843) <= a xor b;
    layer0_outputs(4844) <= not (a or b);
    layer0_outputs(4845) <= not (a or b);
    layer0_outputs(4846) <= a xor b;
    layer0_outputs(4847) <= a;
    layer0_outputs(4848) <= a or b;
    layer0_outputs(4849) <= a or b;
    layer0_outputs(4850) <= not (a or b);
    layer0_outputs(4851) <= not (a xor b);
    layer0_outputs(4852) <= a and not b;
    layer0_outputs(4853) <= a or b;
    layer0_outputs(4854) <= not a or b;
    layer0_outputs(4855) <= not (a xor b);
    layer0_outputs(4856) <= b;
    layer0_outputs(4857) <= not b or a;
    layer0_outputs(4858) <= a or b;
    layer0_outputs(4859) <= a or b;
    layer0_outputs(4860) <= not (a xor b);
    layer0_outputs(4861) <= not b;
    layer0_outputs(4862) <= not (a or b);
    layer0_outputs(4863) <= not (a or b);
    layer0_outputs(4864) <= not b;
    layer0_outputs(4865) <= not a or b;
    layer0_outputs(4866) <= 1'b0;
    layer0_outputs(4867) <= not b or a;
    layer0_outputs(4868) <= not b;
    layer0_outputs(4869) <= a;
    layer0_outputs(4870) <= not (a xor b);
    layer0_outputs(4871) <= a or b;
    layer0_outputs(4872) <= not (a xor b);
    layer0_outputs(4873) <= a or b;
    layer0_outputs(4874) <= a xor b;
    layer0_outputs(4875) <= a or b;
    layer0_outputs(4876) <= b;
    layer0_outputs(4877) <= not (a or b);
    layer0_outputs(4878) <= not a;
    layer0_outputs(4879) <= not b;
    layer0_outputs(4880) <= a and not b;
    layer0_outputs(4881) <= a xor b;
    layer0_outputs(4882) <= a or b;
    layer0_outputs(4883) <= a or b;
    layer0_outputs(4884) <= b;
    layer0_outputs(4885) <= a;
    layer0_outputs(4886) <= not (a and b);
    layer0_outputs(4887) <= not (a xor b);
    layer0_outputs(4888) <= 1'b0;
    layer0_outputs(4889) <= a or b;
    layer0_outputs(4890) <= b;
    layer0_outputs(4891) <= not a;
    layer0_outputs(4892) <= a and not b;
    layer0_outputs(4893) <= not a or b;
    layer0_outputs(4894) <= not (a or b);
    layer0_outputs(4895) <= not (a or b);
    layer0_outputs(4896) <= a and not b;
    layer0_outputs(4897) <= not (a xor b);
    layer0_outputs(4898) <= a or b;
    layer0_outputs(4899) <= not (a xor b);
    layer0_outputs(4900) <= b;
    layer0_outputs(4901) <= b and not a;
    layer0_outputs(4902) <= a xor b;
    layer0_outputs(4903) <= a xor b;
    layer0_outputs(4904) <= not b;
    layer0_outputs(4905) <= b;
    layer0_outputs(4906) <= not a or b;
    layer0_outputs(4907) <= not (a or b);
    layer0_outputs(4908) <= not (a xor b);
    layer0_outputs(4909) <= a;
    layer0_outputs(4910) <= not (a or b);
    layer0_outputs(4911) <= a;
    layer0_outputs(4912) <= a or b;
    layer0_outputs(4913) <= not (a and b);
    layer0_outputs(4914) <= b;
    layer0_outputs(4915) <= a and not b;
    layer0_outputs(4916) <= a and b;
    layer0_outputs(4917) <= a xor b;
    layer0_outputs(4918) <= a xor b;
    layer0_outputs(4919) <= not (a xor b);
    layer0_outputs(4920) <= a or b;
    layer0_outputs(4921) <= not a or b;
    layer0_outputs(4922) <= a or b;
    layer0_outputs(4923) <= a xor b;
    layer0_outputs(4924) <= not b;
    layer0_outputs(4925) <= a;
    layer0_outputs(4926) <= 1'b0;
    layer0_outputs(4927) <= a or b;
    layer0_outputs(4928) <= a or b;
    layer0_outputs(4929) <= not a or b;
    layer0_outputs(4930) <= b;
    layer0_outputs(4931) <= a;
    layer0_outputs(4932) <= not b;
    layer0_outputs(4933) <= a xor b;
    layer0_outputs(4934) <= a;
    layer0_outputs(4935) <= not b;
    layer0_outputs(4936) <= a xor b;
    layer0_outputs(4937) <= not b or a;
    layer0_outputs(4938) <= a or b;
    layer0_outputs(4939) <= a and b;
    layer0_outputs(4940) <= a or b;
    layer0_outputs(4941) <= a;
    layer0_outputs(4942) <= not a or b;
    layer0_outputs(4943) <= a;
    layer0_outputs(4944) <= not (a or b);
    layer0_outputs(4945) <= a;
    layer0_outputs(4946) <= a or b;
    layer0_outputs(4947) <= a xor b;
    layer0_outputs(4948) <= a and b;
    layer0_outputs(4949) <= a xor b;
    layer0_outputs(4950) <= b and not a;
    layer0_outputs(4951) <= a or b;
    layer0_outputs(4952) <= not b or a;
    layer0_outputs(4953) <= a;
    layer0_outputs(4954) <= not (a xor b);
    layer0_outputs(4955) <= not b or a;
    layer0_outputs(4956) <= not a;
    layer0_outputs(4957) <= a or b;
    layer0_outputs(4958) <= a xor b;
    layer0_outputs(4959) <= a and not b;
    layer0_outputs(4960) <= not a;
    layer0_outputs(4961) <= not a or b;
    layer0_outputs(4962) <= a xor b;
    layer0_outputs(4963) <= not (a or b);
    layer0_outputs(4964) <= b;
    layer0_outputs(4965) <= not b or a;
    layer0_outputs(4966) <= a and b;
    layer0_outputs(4967) <= not b;
    layer0_outputs(4968) <= b;
    layer0_outputs(4969) <= a and b;
    layer0_outputs(4970) <= not b or a;
    layer0_outputs(4971) <= not b or a;
    layer0_outputs(4972) <= not (a xor b);
    layer0_outputs(4973) <= not (a and b);
    layer0_outputs(4974) <= a;
    layer0_outputs(4975) <= not (a or b);
    layer0_outputs(4976) <= a and not b;
    layer0_outputs(4977) <= not b or a;
    layer0_outputs(4978) <= a xor b;
    layer0_outputs(4979) <= b;
    layer0_outputs(4980) <= not (a and b);
    layer0_outputs(4981) <= not b;
    layer0_outputs(4982) <= b;
    layer0_outputs(4983) <= a;
    layer0_outputs(4984) <= a and not b;
    layer0_outputs(4985) <= not b;
    layer0_outputs(4986) <= a xor b;
    layer0_outputs(4987) <= b;
    layer0_outputs(4988) <= b;
    layer0_outputs(4989) <= a or b;
    layer0_outputs(4990) <= not (a and b);
    layer0_outputs(4991) <= not (a or b);
    layer0_outputs(4992) <= a;
    layer0_outputs(4993) <= not a or b;
    layer0_outputs(4994) <= b and not a;
    layer0_outputs(4995) <= not b;
    layer0_outputs(4996) <= a;
    layer0_outputs(4997) <= 1'b1;
    layer0_outputs(4998) <= a xor b;
    layer0_outputs(4999) <= not a;
    layer0_outputs(5000) <= not a or b;
    layer0_outputs(5001) <= not (a or b);
    layer0_outputs(5002) <= not (a or b);
    layer0_outputs(5003) <= not b or a;
    layer0_outputs(5004) <= b and not a;
    layer0_outputs(5005) <= b;
    layer0_outputs(5006) <= a;
    layer0_outputs(5007) <= b;
    layer0_outputs(5008) <= not (a xor b);
    layer0_outputs(5009) <= a or b;
    layer0_outputs(5010) <= a and not b;
    layer0_outputs(5011) <= not (a or b);
    layer0_outputs(5012) <= not (a xor b);
    layer0_outputs(5013) <= not a or b;
    layer0_outputs(5014) <= b and not a;
    layer0_outputs(5015) <= not (a and b);
    layer0_outputs(5016) <= a and not b;
    layer0_outputs(5017) <= not b or a;
    layer0_outputs(5018) <= a xor b;
    layer0_outputs(5019) <= not (a and b);
    layer0_outputs(5020) <= not (a xor b);
    layer0_outputs(5021) <= a and not b;
    layer0_outputs(5022) <= b;
    layer0_outputs(5023) <= b;
    layer0_outputs(5024) <= 1'b0;
    layer0_outputs(5025) <= not a;
    layer0_outputs(5026) <= a xor b;
    layer0_outputs(5027) <= not a;
    layer0_outputs(5028) <= not (a or b);
    layer0_outputs(5029) <= a and not b;
    layer0_outputs(5030) <= not b;
    layer0_outputs(5031) <= b and not a;
    layer0_outputs(5032) <= not (a xor b);
    layer0_outputs(5033) <= not (a or b);
    layer0_outputs(5034) <= not (a xor b);
    layer0_outputs(5035) <= not (a and b);
    layer0_outputs(5036) <= not b or a;
    layer0_outputs(5037) <= a and not b;
    layer0_outputs(5038) <= not a or b;
    layer0_outputs(5039) <= a or b;
    layer0_outputs(5040) <= not b;
    layer0_outputs(5041) <= not b or a;
    layer0_outputs(5042) <= a and b;
    layer0_outputs(5043) <= a and not b;
    layer0_outputs(5044) <= not (a xor b);
    layer0_outputs(5045) <= not (a xor b);
    layer0_outputs(5046) <= a or b;
    layer0_outputs(5047) <= b and not a;
    layer0_outputs(5048) <= b;
    layer0_outputs(5049) <= a xor b;
    layer0_outputs(5050) <= a or b;
    layer0_outputs(5051) <= not (a xor b);
    layer0_outputs(5052) <= not a;
    layer0_outputs(5053) <= not (a xor b);
    layer0_outputs(5054) <= b and not a;
    layer0_outputs(5055) <= b;
    layer0_outputs(5056) <= 1'b0;
    layer0_outputs(5057) <= not (a or b);
    layer0_outputs(5058) <= b;
    layer0_outputs(5059) <= b and not a;
    layer0_outputs(5060) <= a;
    layer0_outputs(5061) <= 1'b0;
    layer0_outputs(5062) <= a and not b;
    layer0_outputs(5063) <= not a;
    layer0_outputs(5064) <= not a or b;
    layer0_outputs(5065) <= not a or b;
    layer0_outputs(5066) <= not a;
    layer0_outputs(5067) <= a;
    layer0_outputs(5068) <= not a;
    layer0_outputs(5069) <= not (a xor b);
    layer0_outputs(5070) <= a or b;
    layer0_outputs(5071) <= a xor b;
    layer0_outputs(5072) <= not a or b;
    layer0_outputs(5073) <= not b or a;
    layer0_outputs(5074) <= a;
    layer0_outputs(5075) <= a or b;
    layer0_outputs(5076) <= not b or a;
    layer0_outputs(5077) <= not a;
    layer0_outputs(5078) <= not b or a;
    layer0_outputs(5079) <= b and not a;
    layer0_outputs(5080) <= a;
    layer0_outputs(5081) <= not (a or b);
    layer0_outputs(5082) <= not (a xor b);
    layer0_outputs(5083) <= not (a xor b);
    layer0_outputs(5084) <= b and not a;
    layer0_outputs(5085) <= a xor b;
    layer0_outputs(5086) <= not b or a;
    layer0_outputs(5087) <= not (a or b);
    layer0_outputs(5088) <= not (a or b);
    layer0_outputs(5089) <= a xor b;
    layer0_outputs(5090) <= not (a xor b);
    layer0_outputs(5091) <= a xor b;
    layer0_outputs(5092) <= not a;
    layer0_outputs(5093) <= a or b;
    layer0_outputs(5094) <= a xor b;
    layer0_outputs(5095) <= a or b;
    layer0_outputs(5096) <= 1'b0;
    layer0_outputs(5097) <= not (a xor b);
    layer0_outputs(5098) <= a or b;
    layer0_outputs(5099) <= a or b;
    layer0_outputs(5100) <= not b;
    layer0_outputs(5101) <= not b or a;
    layer0_outputs(5102) <= a or b;
    layer0_outputs(5103) <= a or b;
    layer0_outputs(5104) <= a and b;
    layer0_outputs(5105) <= a xor b;
    layer0_outputs(5106) <= a;
    layer0_outputs(5107) <= not (a or b);
    layer0_outputs(5108) <= a or b;
    layer0_outputs(5109) <= not a or b;
    layer0_outputs(5110) <= b;
    layer0_outputs(5111) <= a xor b;
    layer0_outputs(5112) <= b and not a;
    layer0_outputs(5113) <= a or b;
    layer0_outputs(5114) <= a or b;
    layer0_outputs(5115) <= not (a or b);
    layer0_outputs(5116) <= not a or b;
    layer0_outputs(5117) <= not (a or b);
    layer0_outputs(5118) <= not b;
    layer0_outputs(5119) <= not (a xor b);
    layer0_outputs(5120) <= a or b;
    layer0_outputs(5121) <= not (a or b);
    layer0_outputs(5122) <= not (a xor b);
    layer0_outputs(5123) <= 1'b1;
    layer0_outputs(5124) <= not (a xor b);
    layer0_outputs(5125) <= 1'b1;
    layer0_outputs(5126) <= a or b;
    layer0_outputs(5127) <= a xor b;
    layer0_outputs(5128) <= not a;
    layer0_outputs(5129) <= not (a or b);
    layer0_outputs(5130) <= not (a or b);
    layer0_outputs(5131) <= not (a or b);
    layer0_outputs(5132) <= a or b;
    layer0_outputs(5133) <= b and not a;
    layer0_outputs(5134) <= not (a or b);
    layer0_outputs(5135) <= a and not b;
    layer0_outputs(5136) <= not b;
    layer0_outputs(5137) <= a;
    layer0_outputs(5138) <= 1'b0;
    layer0_outputs(5139) <= a or b;
    layer0_outputs(5140) <= not b or a;
    layer0_outputs(5141) <= not b;
    layer0_outputs(5142) <= b;
    layer0_outputs(5143) <= a and not b;
    layer0_outputs(5144) <= not b or a;
    layer0_outputs(5145) <= not a or b;
    layer0_outputs(5146) <= not b or a;
    layer0_outputs(5147) <= a xor b;
    layer0_outputs(5148) <= a xor b;
    layer0_outputs(5149) <= not b or a;
    layer0_outputs(5150) <= a or b;
    layer0_outputs(5151) <= a;
    layer0_outputs(5152) <= not b;
    layer0_outputs(5153) <= b and not a;
    layer0_outputs(5154) <= a and b;
    layer0_outputs(5155) <= a;
    layer0_outputs(5156) <= a;
    layer0_outputs(5157) <= a and not b;
    layer0_outputs(5158) <= a xor b;
    layer0_outputs(5159) <= not b or a;
    layer0_outputs(5160) <= not a or b;
    layer0_outputs(5161) <= not b or a;
    layer0_outputs(5162) <= 1'b0;
    layer0_outputs(5163) <= not (a xor b);
    layer0_outputs(5164) <= a or b;
    layer0_outputs(5165) <= 1'b0;
    layer0_outputs(5166) <= not (a and b);
    layer0_outputs(5167) <= 1'b1;
    layer0_outputs(5168) <= a and b;
    layer0_outputs(5169) <= not (a xor b);
    layer0_outputs(5170) <= not (a and b);
    layer0_outputs(5171) <= a or b;
    layer0_outputs(5172) <= not (a or b);
    layer0_outputs(5173) <= a and not b;
    layer0_outputs(5174) <= not (a xor b);
    layer0_outputs(5175) <= b and not a;
    layer0_outputs(5176) <= a or b;
    layer0_outputs(5177) <= b;
    layer0_outputs(5178) <= not (a or b);
    layer0_outputs(5179) <= not a;
    layer0_outputs(5180) <= not a;
    layer0_outputs(5181) <= a or b;
    layer0_outputs(5182) <= a and b;
    layer0_outputs(5183) <= not (a xor b);
    layer0_outputs(5184) <= a xor b;
    layer0_outputs(5185) <= not (a or b);
    layer0_outputs(5186) <= a or b;
    layer0_outputs(5187) <= not (a or b);
    layer0_outputs(5188) <= not b or a;
    layer0_outputs(5189) <= not (a or b);
    layer0_outputs(5190) <= b and not a;
    layer0_outputs(5191) <= not (a or b);
    layer0_outputs(5192) <= not (a or b);
    layer0_outputs(5193) <= a or b;
    layer0_outputs(5194) <= not (a xor b);
    layer0_outputs(5195) <= not b or a;
    layer0_outputs(5196) <= not (a or b);
    layer0_outputs(5197) <= 1'b0;
    layer0_outputs(5198) <= a and not b;
    layer0_outputs(5199) <= not (a xor b);
    layer0_outputs(5200) <= a xor b;
    layer0_outputs(5201) <= b and not a;
    layer0_outputs(5202) <= a and not b;
    layer0_outputs(5203) <= not b or a;
    layer0_outputs(5204) <= a or b;
    layer0_outputs(5205) <= a and not b;
    layer0_outputs(5206) <= a or b;
    layer0_outputs(5207) <= not a or b;
    layer0_outputs(5208) <= not (a xor b);
    layer0_outputs(5209) <= not a;
    layer0_outputs(5210) <= not a or b;
    layer0_outputs(5211) <= not (a or b);
    layer0_outputs(5212) <= not (a xor b);
    layer0_outputs(5213) <= a xor b;
    layer0_outputs(5214) <= a or b;
    layer0_outputs(5215) <= not (a or b);
    layer0_outputs(5216) <= a or b;
    layer0_outputs(5217) <= not (a or b);
    layer0_outputs(5218) <= a;
    layer0_outputs(5219) <= not b or a;
    layer0_outputs(5220) <= a;
    layer0_outputs(5221) <= not (a or b);
    layer0_outputs(5222) <= not a;
    layer0_outputs(5223) <= a or b;
    layer0_outputs(5224) <= b;
    layer0_outputs(5225) <= 1'b1;
    layer0_outputs(5226) <= not (a or b);
    layer0_outputs(5227) <= not (a xor b);
    layer0_outputs(5228) <= not b;
    layer0_outputs(5229) <= not b;
    layer0_outputs(5230) <= a;
    layer0_outputs(5231) <= not a;
    layer0_outputs(5232) <= a;
    layer0_outputs(5233) <= b and not a;
    layer0_outputs(5234) <= not b;
    layer0_outputs(5235) <= a or b;
    layer0_outputs(5236) <= a and not b;
    layer0_outputs(5237) <= not (a or b);
    layer0_outputs(5238) <= a xor b;
    layer0_outputs(5239) <= not b;
    layer0_outputs(5240) <= a and not b;
    layer0_outputs(5241) <= not b;
    layer0_outputs(5242) <= not b;
    layer0_outputs(5243) <= not b or a;
    layer0_outputs(5244) <= not (a xor b);
    layer0_outputs(5245) <= a or b;
    layer0_outputs(5246) <= a;
    layer0_outputs(5247) <= a and not b;
    layer0_outputs(5248) <= not (a or b);
    layer0_outputs(5249) <= b and not a;
    layer0_outputs(5250) <= not (a or b);
    layer0_outputs(5251) <= b;
    layer0_outputs(5252) <= a xor b;
    layer0_outputs(5253) <= not b or a;
    layer0_outputs(5254) <= a xor b;
    layer0_outputs(5255) <= a or b;
    layer0_outputs(5256) <= a;
    layer0_outputs(5257) <= a and not b;
    layer0_outputs(5258) <= a or b;
    layer0_outputs(5259) <= a xor b;
    layer0_outputs(5260) <= not b or a;
    layer0_outputs(5261) <= b and not a;
    layer0_outputs(5262) <= a and not b;
    layer0_outputs(5263) <= a and not b;
    layer0_outputs(5264) <= not a or b;
    layer0_outputs(5265) <= not (a or b);
    layer0_outputs(5266) <= not a or b;
    layer0_outputs(5267) <= b;
    layer0_outputs(5268) <= b and not a;
    layer0_outputs(5269) <= not (a or b);
    layer0_outputs(5270) <= b and not a;
    layer0_outputs(5271) <= not (a xor b);
    layer0_outputs(5272) <= a xor b;
    layer0_outputs(5273) <= not b;
    layer0_outputs(5274) <= a;
    layer0_outputs(5275) <= not b;
    layer0_outputs(5276) <= not b or a;
    layer0_outputs(5277) <= not (a and b);
    layer0_outputs(5278) <= not (a xor b);
    layer0_outputs(5279) <= a xor b;
    layer0_outputs(5280) <= not (a or b);
    layer0_outputs(5281) <= not (a xor b);
    layer0_outputs(5282) <= not (a or b);
    layer0_outputs(5283) <= a and b;
    layer0_outputs(5284) <= not a;
    layer0_outputs(5285) <= 1'b0;
    layer0_outputs(5286) <= a;
    layer0_outputs(5287) <= a xor b;
    layer0_outputs(5288) <= a;
    layer0_outputs(5289) <= a or b;
    layer0_outputs(5290) <= not b;
    layer0_outputs(5291) <= b and not a;
    layer0_outputs(5292) <= not (a xor b);
    layer0_outputs(5293) <= not (a xor b);
    layer0_outputs(5294) <= b;
    layer0_outputs(5295) <= a or b;
    layer0_outputs(5296) <= a and not b;
    layer0_outputs(5297) <= a xor b;
    layer0_outputs(5298) <= not (a xor b);
    layer0_outputs(5299) <= a or b;
    layer0_outputs(5300) <= not a or b;
    layer0_outputs(5301) <= a;
    layer0_outputs(5302) <= not a;
    layer0_outputs(5303) <= not (a xor b);
    layer0_outputs(5304) <= b;
    layer0_outputs(5305) <= a or b;
    layer0_outputs(5306) <= not a or b;
    layer0_outputs(5307) <= a and not b;
    layer0_outputs(5308) <= not (a and b);
    layer0_outputs(5309) <= not (a or b);
    layer0_outputs(5310) <= not a;
    layer0_outputs(5311) <= a;
    layer0_outputs(5312) <= not (a and b);
    layer0_outputs(5313) <= a;
    layer0_outputs(5314) <= not (a xor b);
    layer0_outputs(5315) <= a or b;
    layer0_outputs(5316) <= a;
    layer0_outputs(5317) <= a and not b;
    layer0_outputs(5318) <= a xor b;
    layer0_outputs(5319) <= 1'b0;
    layer0_outputs(5320) <= a and not b;
    layer0_outputs(5321) <= a or b;
    layer0_outputs(5322) <= not a;
    layer0_outputs(5323) <= b and not a;
    layer0_outputs(5324) <= not a or b;
    layer0_outputs(5325) <= not b or a;
    layer0_outputs(5326) <= a or b;
    layer0_outputs(5327) <= b and not a;
    layer0_outputs(5328) <= not b;
    layer0_outputs(5329) <= a or b;
    layer0_outputs(5330) <= not (a or b);
    layer0_outputs(5331) <= a or b;
    layer0_outputs(5332) <= not (a or b);
    layer0_outputs(5333) <= not (a or b);
    layer0_outputs(5334) <= not a;
    layer0_outputs(5335) <= a xor b;
    layer0_outputs(5336) <= b;
    layer0_outputs(5337) <= a and not b;
    layer0_outputs(5338) <= b and not a;
    layer0_outputs(5339) <= b and not a;
    layer0_outputs(5340) <= a or b;
    layer0_outputs(5341) <= a;
    layer0_outputs(5342) <= not a;
    layer0_outputs(5343) <= b and not a;
    layer0_outputs(5344) <= not (a xor b);
    layer0_outputs(5345) <= a or b;
    layer0_outputs(5346) <= not (a or b);
    layer0_outputs(5347) <= not a;
    layer0_outputs(5348) <= a and not b;
    layer0_outputs(5349) <= not (a and b);
    layer0_outputs(5350) <= a xor b;
    layer0_outputs(5351) <= b and not a;
    layer0_outputs(5352) <= a and not b;
    layer0_outputs(5353) <= a and not b;
    layer0_outputs(5354) <= b;
    layer0_outputs(5355) <= 1'b1;
    layer0_outputs(5356) <= not (a or b);
    layer0_outputs(5357) <= b and not a;
    layer0_outputs(5358) <= not b or a;
    layer0_outputs(5359) <= not a;
    layer0_outputs(5360) <= a;
    layer0_outputs(5361) <= b;
    layer0_outputs(5362) <= a xor b;
    layer0_outputs(5363) <= b;
    layer0_outputs(5364) <= not (a xor b);
    layer0_outputs(5365) <= a xor b;
    layer0_outputs(5366) <= b and not a;
    layer0_outputs(5367) <= a or b;
    layer0_outputs(5368) <= not (a xor b);
    layer0_outputs(5369) <= b;
    layer0_outputs(5370) <= not (a or b);
    layer0_outputs(5371) <= not (a or b);
    layer0_outputs(5372) <= a or b;
    layer0_outputs(5373) <= not b or a;
    layer0_outputs(5374) <= not a or b;
    layer0_outputs(5375) <= not (a or b);
    layer0_outputs(5376) <= b;
    layer0_outputs(5377) <= not (a xor b);
    layer0_outputs(5378) <= a xor b;
    layer0_outputs(5379) <= a xor b;
    layer0_outputs(5380) <= a and not b;
    layer0_outputs(5381) <= b;
    layer0_outputs(5382) <= a and b;
    layer0_outputs(5383) <= a or b;
    layer0_outputs(5384) <= not b;
    layer0_outputs(5385) <= not a;
    layer0_outputs(5386) <= a xor b;
    layer0_outputs(5387) <= not (a xor b);
    layer0_outputs(5388) <= not (a or b);
    layer0_outputs(5389) <= a or b;
    layer0_outputs(5390) <= a or b;
    layer0_outputs(5391) <= not b or a;
    layer0_outputs(5392) <= a or b;
    layer0_outputs(5393) <= not b;
    layer0_outputs(5394) <= a or b;
    layer0_outputs(5395) <= a xor b;
    layer0_outputs(5396) <= b;
    layer0_outputs(5397) <= not b;
    layer0_outputs(5398) <= not (a or b);
    layer0_outputs(5399) <= a xor b;
    layer0_outputs(5400) <= not b or a;
    layer0_outputs(5401) <= not a;
    layer0_outputs(5402) <= not (a or b);
    layer0_outputs(5403) <= a;
    layer0_outputs(5404) <= a xor b;
    layer0_outputs(5405) <= a;
    layer0_outputs(5406) <= a or b;
    layer0_outputs(5407) <= a and not b;
    layer0_outputs(5408) <= not (a or b);
    layer0_outputs(5409) <= not b;
    layer0_outputs(5410) <= a and b;
    layer0_outputs(5411) <= a xor b;
    layer0_outputs(5412) <= 1'b1;
    layer0_outputs(5413) <= not (a xor b);
    layer0_outputs(5414) <= a xor b;
    layer0_outputs(5415) <= b;
    layer0_outputs(5416) <= not (a xor b);
    layer0_outputs(5417) <= not (a or b);
    layer0_outputs(5418) <= a;
    layer0_outputs(5419) <= not b or a;
    layer0_outputs(5420) <= 1'b0;
    layer0_outputs(5421) <= not (a and b);
    layer0_outputs(5422) <= not b or a;
    layer0_outputs(5423) <= not (a or b);
    layer0_outputs(5424) <= not a;
    layer0_outputs(5425) <= a and b;
    layer0_outputs(5426) <= b;
    layer0_outputs(5427) <= a;
    layer0_outputs(5428) <= not (a or b);
    layer0_outputs(5429) <= a;
    layer0_outputs(5430) <= a or b;
    layer0_outputs(5431) <= 1'b1;
    layer0_outputs(5432) <= not a;
    layer0_outputs(5433) <= not (a and b);
    layer0_outputs(5434) <= not a;
    layer0_outputs(5435) <= b;
    layer0_outputs(5436) <= b;
    layer0_outputs(5437) <= b;
    layer0_outputs(5438) <= not (a or b);
    layer0_outputs(5439) <= 1'b0;
    layer0_outputs(5440) <= b;
    layer0_outputs(5441) <= a xor b;
    layer0_outputs(5442) <= a and not b;
    layer0_outputs(5443) <= not (a or b);
    layer0_outputs(5444) <= 1'b1;
    layer0_outputs(5445) <= b and not a;
    layer0_outputs(5446) <= a or b;
    layer0_outputs(5447) <= a or b;
    layer0_outputs(5448) <= a xor b;
    layer0_outputs(5449) <= b;
    layer0_outputs(5450) <= a;
    layer0_outputs(5451) <= b and not a;
    layer0_outputs(5452) <= a and not b;
    layer0_outputs(5453) <= not (a or b);
    layer0_outputs(5454) <= a xor b;
    layer0_outputs(5455) <= a xor b;
    layer0_outputs(5456) <= not a or b;
    layer0_outputs(5457) <= not b or a;
    layer0_outputs(5458) <= a xor b;
    layer0_outputs(5459) <= a or b;
    layer0_outputs(5460) <= a or b;
    layer0_outputs(5461) <= not b;
    layer0_outputs(5462) <= not a;
    layer0_outputs(5463) <= 1'b1;
    layer0_outputs(5464) <= not b;
    layer0_outputs(5465) <= not (a or b);
    layer0_outputs(5466) <= a or b;
    layer0_outputs(5467) <= a xor b;
    layer0_outputs(5468) <= a or b;
    layer0_outputs(5469) <= not (a xor b);
    layer0_outputs(5470) <= not (a or b);
    layer0_outputs(5471) <= a or b;
    layer0_outputs(5472) <= not b;
    layer0_outputs(5473) <= a and not b;
    layer0_outputs(5474) <= a or b;
    layer0_outputs(5475) <= not a;
    layer0_outputs(5476) <= a or b;
    layer0_outputs(5477) <= a and not b;
    layer0_outputs(5478) <= b and not a;
    layer0_outputs(5479) <= not a or b;
    layer0_outputs(5480) <= a;
    layer0_outputs(5481) <= a and not b;
    layer0_outputs(5482) <= a and b;
    layer0_outputs(5483) <= b and not a;
    layer0_outputs(5484) <= a xor b;
    layer0_outputs(5485) <= a and b;
    layer0_outputs(5486) <= a xor b;
    layer0_outputs(5487) <= not (a xor b);
    layer0_outputs(5488) <= not (a or b);
    layer0_outputs(5489) <= a and not b;
    layer0_outputs(5490) <= a xor b;
    layer0_outputs(5491) <= a xor b;
    layer0_outputs(5492) <= not a or b;
    layer0_outputs(5493) <= not a or b;
    layer0_outputs(5494) <= a xor b;
    layer0_outputs(5495) <= a and b;
    layer0_outputs(5496) <= not (a xor b);
    layer0_outputs(5497) <= a and not b;
    layer0_outputs(5498) <= not (a xor b);
    layer0_outputs(5499) <= a or b;
    layer0_outputs(5500) <= not (a xor b);
    layer0_outputs(5501) <= a xor b;
    layer0_outputs(5502) <= a and not b;
    layer0_outputs(5503) <= not (a or b);
    layer0_outputs(5504) <= a or b;
    layer0_outputs(5505) <= not b;
    layer0_outputs(5506) <= b and not a;
    layer0_outputs(5507) <= not b;
    layer0_outputs(5508) <= not b or a;
    layer0_outputs(5509) <= not (a xor b);
    layer0_outputs(5510) <= not b or a;
    layer0_outputs(5511) <= not (a or b);
    layer0_outputs(5512) <= not b or a;
    layer0_outputs(5513) <= 1'b0;
    layer0_outputs(5514) <= not a;
    layer0_outputs(5515) <= a xor b;
    layer0_outputs(5516) <= not b or a;
    layer0_outputs(5517) <= not b or a;
    layer0_outputs(5518) <= a;
    layer0_outputs(5519) <= b and not a;
    layer0_outputs(5520) <= a or b;
    layer0_outputs(5521) <= a;
    layer0_outputs(5522) <= a or b;
    layer0_outputs(5523) <= not b or a;
    layer0_outputs(5524) <= b and not a;
    layer0_outputs(5525) <= not b;
    layer0_outputs(5526) <= b;
    layer0_outputs(5527) <= not (a or b);
    layer0_outputs(5528) <= b and not a;
    layer0_outputs(5529) <= 1'b1;
    layer0_outputs(5530) <= a or b;
    layer0_outputs(5531) <= a and not b;
    layer0_outputs(5532) <= not (a xor b);
    layer0_outputs(5533) <= a;
    layer0_outputs(5534) <= not a or b;
    layer0_outputs(5535) <= a and not b;
    layer0_outputs(5536) <= not a;
    layer0_outputs(5537) <= a;
    layer0_outputs(5538) <= not a or b;
    layer0_outputs(5539) <= not (a xor b);
    layer0_outputs(5540) <= not (a or b);
    layer0_outputs(5541) <= not b or a;
    layer0_outputs(5542) <= not a;
    layer0_outputs(5543) <= a and b;
    layer0_outputs(5544) <= not (a or b);
    layer0_outputs(5545) <= not (a xor b);
    layer0_outputs(5546) <= a;
    layer0_outputs(5547) <= a and not b;
    layer0_outputs(5548) <= not b or a;
    layer0_outputs(5549) <= b;
    layer0_outputs(5550) <= not a;
    layer0_outputs(5551) <= a and not b;
    layer0_outputs(5552) <= a and not b;
    layer0_outputs(5553) <= not a;
    layer0_outputs(5554) <= 1'b1;
    layer0_outputs(5555) <= b;
    layer0_outputs(5556) <= not b;
    layer0_outputs(5557) <= not (a xor b);
    layer0_outputs(5558) <= not (a or b);
    layer0_outputs(5559) <= b and not a;
    layer0_outputs(5560) <= not b or a;
    layer0_outputs(5561) <= not (a or b);
    layer0_outputs(5562) <= a or b;
    layer0_outputs(5563) <= 1'b0;
    layer0_outputs(5564) <= a and b;
    layer0_outputs(5565) <= not a or b;
    layer0_outputs(5566) <= not a;
    layer0_outputs(5567) <= a;
    layer0_outputs(5568) <= a xor b;
    layer0_outputs(5569) <= not (a and b);
    layer0_outputs(5570) <= a or b;
    layer0_outputs(5571) <= a xor b;
    layer0_outputs(5572) <= not (a xor b);
    layer0_outputs(5573) <= not a;
    layer0_outputs(5574) <= a and b;
    layer0_outputs(5575) <= a and not b;
    layer0_outputs(5576) <= a and not b;
    layer0_outputs(5577) <= not b;
    layer0_outputs(5578) <= not a or b;
    layer0_outputs(5579) <= not (a xor b);
    layer0_outputs(5580) <= not (a or b);
    layer0_outputs(5581) <= not b or a;
    layer0_outputs(5582) <= a xor b;
    layer0_outputs(5583) <= a and b;
    layer0_outputs(5584) <= a xor b;
    layer0_outputs(5585) <= not (a or b);
    layer0_outputs(5586) <= a or b;
    layer0_outputs(5587) <= not (a or b);
    layer0_outputs(5588) <= not (a or b);
    layer0_outputs(5589) <= a or b;
    layer0_outputs(5590) <= not a;
    layer0_outputs(5591) <= not a or b;
    layer0_outputs(5592) <= b and not a;
    layer0_outputs(5593) <= not b or a;
    layer0_outputs(5594) <= a xor b;
    layer0_outputs(5595) <= not b;
    layer0_outputs(5596) <= a or b;
    layer0_outputs(5597) <= a xor b;
    layer0_outputs(5598) <= a or b;
    layer0_outputs(5599) <= b;
    layer0_outputs(5600) <= b and not a;
    layer0_outputs(5601) <= not (a xor b);
    layer0_outputs(5602) <= b;
    layer0_outputs(5603) <= not (a xor b);
    layer0_outputs(5604) <= not a or b;
    layer0_outputs(5605) <= a;
    layer0_outputs(5606) <= not b;
    layer0_outputs(5607) <= not b or a;
    layer0_outputs(5608) <= not b;
    layer0_outputs(5609) <= b;
    layer0_outputs(5610) <= a or b;
    layer0_outputs(5611) <= not b or a;
    layer0_outputs(5612) <= a and b;
    layer0_outputs(5613) <= not b or a;
    layer0_outputs(5614) <= a xor b;
    layer0_outputs(5615) <= not (a or b);
    layer0_outputs(5616) <= not (a or b);
    layer0_outputs(5617) <= not a or b;
    layer0_outputs(5618) <= not a or b;
    layer0_outputs(5619) <= a and not b;
    layer0_outputs(5620) <= b;
    layer0_outputs(5621) <= b and not a;
    layer0_outputs(5622) <= not a;
    layer0_outputs(5623) <= b;
    layer0_outputs(5624) <= not a;
    layer0_outputs(5625) <= not a;
    layer0_outputs(5626) <= not b or a;
    layer0_outputs(5627) <= b;
    layer0_outputs(5628) <= not (a xor b);
    layer0_outputs(5629) <= 1'b1;
    layer0_outputs(5630) <= a or b;
    layer0_outputs(5631) <= 1'b0;
    layer0_outputs(5632) <= not b or a;
    layer0_outputs(5633) <= not (a or b);
    layer0_outputs(5634) <= not b or a;
    layer0_outputs(5635) <= b and not a;
    layer0_outputs(5636) <= b and not a;
    layer0_outputs(5637) <= a;
    layer0_outputs(5638) <= not (a or b);
    layer0_outputs(5639) <= not (a or b);
    layer0_outputs(5640) <= 1'b0;
    layer0_outputs(5641) <= not b;
    layer0_outputs(5642) <= a or b;
    layer0_outputs(5643) <= not b;
    layer0_outputs(5644) <= not (a or b);
    layer0_outputs(5645) <= a xor b;
    layer0_outputs(5646) <= a or b;
    layer0_outputs(5647) <= not b or a;
    layer0_outputs(5648) <= a or b;
    layer0_outputs(5649) <= not (a or b);
    layer0_outputs(5650) <= a;
    layer0_outputs(5651) <= a or b;
    layer0_outputs(5652) <= not (a xor b);
    layer0_outputs(5653) <= not (a xor b);
    layer0_outputs(5654) <= a;
    layer0_outputs(5655) <= a or b;
    layer0_outputs(5656) <= not b;
    layer0_outputs(5657) <= b and not a;
    layer0_outputs(5658) <= not b;
    layer0_outputs(5659) <= not b;
    layer0_outputs(5660) <= not (a and b);
    layer0_outputs(5661) <= not (a or b);
    layer0_outputs(5662) <= not a;
    layer0_outputs(5663) <= not b or a;
    layer0_outputs(5664) <= a xor b;
    layer0_outputs(5665) <= not b or a;
    layer0_outputs(5666) <= a or b;
    layer0_outputs(5667) <= not a;
    layer0_outputs(5668) <= a or b;
    layer0_outputs(5669) <= not b or a;
    layer0_outputs(5670) <= not a or b;
    layer0_outputs(5671) <= a and not b;
    layer0_outputs(5672) <= a or b;
    layer0_outputs(5673) <= not (a or b);
    layer0_outputs(5674) <= not a;
    layer0_outputs(5675) <= a xor b;
    layer0_outputs(5676) <= b and not a;
    layer0_outputs(5677) <= a xor b;
    layer0_outputs(5678) <= not a;
    layer0_outputs(5679) <= a;
    layer0_outputs(5680) <= a or b;
    layer0_outputs(5681) <= not b;
    layer0_outputs(5682) <= b;
    layer0_outputs(5683) <= a and b;
    layer0_outputs(5684) <= not (a or b);
    layer0_outputs(5685) <= a xor b;
    layer0_outputs(5686) <= b;
    layer0_outputs(5687) <= not (a or b);
    layer0_outputs(5688) <= a or b;
    layer0_outputs(5689) <= not (a xor b);
    layer0_outputs(5690) <= not (a or b);
    layer0_outputs(5691) <= a xor b;
    layer0_outputs(5692) <= not a or b;
    layer0_outputs(5693) <= not b or a;
    layer0_outputs(5694) <= a;
    layer0_outputs(5695) <= b and not a;
    layer0_outputs(5696) <= a or b;
    layer0_outputs(5697) <= 1'b1;
    layer0_outputs(5698) <= not b or a;
    layer0_outputs(5699) <= not (a and b);
    layer0_outputs(5700) <= a or b;
    layer0_outputs(5701) <= a or b;
    layer0_outputs(5702) <= not (a or b);
    layer0_outputs(5703) <= not a;
    layer0_outputs(5704) <= a or b;
    layer0_outputs(5705) <= not b;
    layer0_outputs(5706) <= not a;
    layer0_outputs(5707) <= a xor b;
    layer0_outputs(5708) <= not (a and b);
    layer0_outputs(5709) <= not (a or b);
    layer0_outputs(5710) <= not (a xor b);
    layer0_outputs(5711) <= b and not a;
    layer0_outputs(5712) <= not (a or b);
    layer0_outputs(5713) <= a and not b;
    layer0_outputs(5714) <= a xor b;
    layer0_outputs(5715) <= a or b;
    layer0_outputs(5716) <= a;
    layer0_outputs(5717) <= a and not b;
    layer0_outputs(5718) <= not (a or b);
    layer0_outputs(5719) <= a or b;
    layer0_outputs(5720) <= not b or a;
    layer0_outputs(5721) <= not (a or b);
    layer0_outputs(5722) <= not (a xor b);
    layer0_outputs(5723) <= not (a xor b);
    layer0_outputs(5724) <= not b;
    layer0_outputs(5725) <= not a or b;
    layer0_outputs(5726) <= not b;
    layer0_outputs(5727) <= a or b;
    layer0_outputs(5728) <= a or b;
    layer0_outputs(5729) <= not (a or b);
    layer0_outputs(5730) <= b and not a;
    layer0_outputs(5731) <= not b;
    layer0_outputs(5732) <= not b;
    layer0_outputs(5733) <= a or b;
    layer0_outputs(5734) <= not (a xor b);
    layer0_outputs(5735) <= not (a or b);
    layer0_outputs(5736) <= not (a xor b);
    layer0_outputs(5737) <= not (a or b);
    layer0_outputs(5738) <= not a or b;
    layer0_outputs(5739) <= not (a or b);
    layer0_outputs(5740) <= a;
    layer0_outputs(5741) <= a;
    layer0_outputs(5742) <= a and not b;
    layer0_outputs(5743) <= not (a or b);
    layer0_outputs(5744) <= a and b;
    layer0_outputs(5745) <= a;
    layer0_outputs(5746) <= a;
    layer0_outputs(5747) <= a;
    layer0_outputs(5748) <= b;
    layer0_outputs(5749) <= not (a xor b);
    layer0_outputs(5750) <= not a or b;
    layer0_outputs(5751) <= not (a or b);
    layer0_outputs(5752) <= not (a or b);
    layer0_outputs(5753) <= not a or b;
    layer0_outputs(5754) <= b;
    layer0_outputs(5755) <= a and not b;
    layer0_outputs(5756) <= a and not b;
    layer0_outputs(5757) <= 1'b1;
    layer0_outputs(5758) <= b and not a;
    layer0_outputs(5759) <= not (a and b);
    layer0_outputs(5760) <= a and not b;
    layer0_outputs(5761) <= a;
    layer0_outputs(5762) <= a xor b;
    layer0_outputs(5763) <= not (a and b);
    layer0_outputs(5764) <= a or b;
    layer0_outputs(5765) <= not (a or b);
    layer0_outputs(5766) <= not (a xor b);
    layer0_outputs(5767) <= b;
    layer0_outputs(5768) <= not a or b;
    layer0_outputs(5769) <= not a;
    layer0_outputs(5770) <= b and not a;
    layer0_outputs(5771) <= a and b;
    layer0_outputs(5772) <= a;
    layer0_outputs(5773) <= a and not b;
    layer0_outputs(5774) <= a xor b;
    layer0_outputs(5775) <= not b;
    layer0_outputs(5776) <= b;
    layer0_outputs(5777) <= a;
    layer0_outputs(5778) <= not a or b;
    layer0_outputs(5779) <= not (a or b);
    layer0_outputs(5780) <= not a;
    layer0_outputs(5781) <= not b;
    layer0_outputs(5782) <= a;
    layer0_outputs(5783) <= not a;
    layer0_outputs(5784) <= not b or a;
    layer0_outputs(5785) <= not (a xor b);
    layer0_outputs(5786) <= not (a or b);
    layer0_outputs(5787) <= not a;
    layer0_outputs(5788) <= a;
    layer0_outputs(5789) <= not b;
    layer0_outputs(5790) <= not b;
    layer0_outputs(5791) <= not a;
    layer0_outputs(5792) <= a xor b;
    layer0_outputs(5793) <= not (a xor b);
    layer0_outputs(5794) <= a xor b;
    layer0_outputs(5795) <= a and not b;
    layer0_outputs(5796) <= not (a or b);
    layer0_outputs(5797) <= not (a or b);
    layer0_outputs(5798) <= a;
    layer0_outputs(5799) <= a and not b;
    layer0_outputs(5800) <= a and not b;
    layer0_outputs(5801) <= not b;
    layer0_outputs(5802) <= not (a or b);
    layer0_outputs(5803) <= b;
    layer0_outputs(5804) <= a or b;
    layer0_outputs(5805) <= not (a or b);
    layer0_outputs(5806) <= not (a xor b);
    layer0_outputs(5807) <= not a or b;
    layer0_outputs(5808) <= a;
    layer0_outputs(5809) <= not a;
    layer0_outputs(5810) <= not (a xor b);
    layer0_outputs(5811) <= not a;
    layer0_outputs(5812) <= not a or b;
    layer0_outputs(5813) <= not b or a;
    layer0_outputs(5814) <= not b or a;
    layer0_outputs(5815) <= not (a xor b);
    layer0_outputs(5816) <= a xor b;
    layer0_outputs(5817) <= not b or a;
    layer0_outputs(5818) <= not a or b;
    layer0_outputs(5819) <= a xor b;
    layer0_outputs(5820) <= not (a xor b);
    layer0_outputs(5821) <= a and not b;
    layer0_outputs(5822) <= not b or a;
    layer0_outputs(5823) <= not b;
    layer0_outputs(5824) <= not (a or b);
    layer0_outputs(5825) <= a xor b;
    layer0_outputs(5826) <= not a;
    layer0_outputs(5827) <= not a or b;
    layer0_outputs(5828) <= a;
    layer0_outputs(5829) <= not a;
    layer0_outputs(5830) <= not b or a;
    layer0_outputs(5831) <= b and not a;
    layer0_outputs(5832) <= b and not a;
    layer0_outputs(5833) <= a;
    layer0_outputs(5834) <= not (a or b);
    layer0_outputs(5835) <= b;
    layer0_outputs(5836) <= not (a xor b);
    layer0_outputs(5837) <= not b or a;
    layer0_outputs(5838) <= not a or b;
    layer0_outputs(5839) <= not (a and b);
    layer0_outputs(5840) <= a xor b;
    layer0_outputs(5841) <= a or b;
    layer0_outputs(5842) <= b;
    layer0_outputs(5843) <= not (a or b);
    layer0_outputs(5844) <= not (a xor b);
    layer0_outputs(5845) <= not a or b;
    layer0_outputs(5846) <= a xor b;
    layer0_outputs(5847) <= not a;
    layer0_outputs(5848) <= b;
    layer0_outputs(5849) <= not (a or b);
    layer0_outputs(5850) <= a xor b;
    layer0_outputs(5851) <= not b;
    layer0_outputs(5852) <= not b;
    layer0_outputs(5853) <= not (a xor b);
    layer0_outputs(5854) <= not (a or b);
    layer0_outputs(5855) <= not (a or b);
    layer0_outputs(5856) <= a xor b;
    layer0_outputs(5857) <= b;
    layer0_outputs(5858) <= not a or b;
    layer0_outputs(5859) <= not (a or b);
    layer0_outputs(5860) <= a xor b;
    layer0_outputs(5861) <= b;
    layer0_outputs(5862) <= b;
    layer0_outputs(5863) <= not (a xor b);
    layer0_outputs(5864) <= not a;
    layer0_outputs(5865) <= not (a xor b);
    layer0_outputs(5866) <= a or b;
    layer0_outputs(5867) <= a xor b;
    layer0_outputs(5868) <= not (a or b);
    layer0_outputs(5869) <= not (a or b);
    layer0_outputs(5870) <= a;
    layer0_outputs(5871) <= not b or a;
    layer0_outputs(5872) <= b;
    layer0_outputs(5873) <= a xor b;
    layer0_outputs(5874) <= a or b;
    layer0_outputs(5875) <= not b;
    layer0_outputs(5876) <= a or b;
    layer0_outputs(5877) <= not a or b;
    layer0_outputs(5878) <= not (a or b);
    layer0_outputs(5879) <= not (a or b);
    layer0_outputs(5880) <= a xor b;
    layer0_outputs(5881) <= a and not b;
    layer0_outputs(5882) <= not a or b;
    layer0_outputs(5883) <= a xor b;
    layer0_outputs(5884) <= a or b;
    layer0_outputs(5885) <= b;
    layer0_outputs(5886) <= not b or a;
    layer0_outputs(5887) <= not b or a;
    layer0_outputs(5888) <= a xor b;
    layer0_outputs(5889) <= a;
    layer0_outputs(5890) <= not (a or b);
    layer0_outputs(5891) <= b and not a;
    layer0_outputs(5892) <= a and not b;
    layer0_outputs(5893) <= a and not b;
    layer0_outputs(5894) <= not a or b;
    layer0_outputs(5895) <= not b or a;
    layer0_outputs(5896) <= not (a xor b);
    layer0_outputs(5897) <= not b or a;
    layer0_outputs(5898) <= not b or a;
    layer0_outputs(5899) <= not (a or b);
    layer0_outputs(5900) <= not b or a;
    layer0_outputs(5901) <= b and not a;
    layer0_outputs(5902) <= not a;
    layer0_outputs(5903) <= a or b;
    layer0_outputs(5904) <= not b;
    layer0_outputs(5905) <= a xor b;
    layer0_outputs(5906) <= a and not b;
    layer0_outputs(5907) <= not b;
    layer0_outputs(5908) <= a and not b;
    layer0_outputs(5909) <= not (a xor b);
    layer0_outputs(5910) <= not a or b;
    layer0_outputs(5911) <= b;
    layer0_outputs(5912) <= not (a xor b);
    layer0_outputs(5913) <= a;
    layer0_outputs(5914) <= not (a or b);
    layer0_outputs(5915) <= not b or a;
    layer0_outputs(5916) <= not a;
    layer0_outputs(5917) <= b and not a;
    layer0_outputs(5918) <= not b or a;
    layer0_outputs(5919) <= a xor b;
    layer0_outputs(5920) <= b;
    layer0_outputs(5921) <= 1'b0;
    layer0_outputs(5922) <= not (a xor b);
    layer0_outputs(5923) <= a and b;
    layer0_outputs(5924) <= b and not a;
    layer0_outputs(5925) <= not (a xor b);
    layer0_outputs(5926) <= not a or b;
    layer0_outputs(5927) <= a and b;
    layer0_outputs(5928) <= not (a or b);
    layer0_outputs(5929) <= a xor b;
    layer0_outputs(5930) <= a;
    layer0_outputs(5931) <= not b or a;
    layer0_outputs(5932) <= a or b;
    layer0_outputs(5933) <= a and not b;
    layer0_outputs(5934) <= not (a xor b);
    layer0_outputs(5935) <= not (a or b);
    layer0_outputs(5936) <= not (a or b);
    layer0_outputs(5937) <= not b or a;
    layer0_outputs(5938) <= not (a or b);
    layer0_outputs(5939) <= a;
    layer0_outputs(5940) <= b and not a;
    layer0_outputs(5941) <= not a;
    layer0_outputs(5942) <= not (a or b);
    layer0_outputs(5943) <= a xor b;
    layer0_outputs(5944) <= not b or a;
    layer0_outputs(5945) <= not b or a;
    layer0_outputs(5946) <= not b;
    layer0_outputs(5947) <= a and b;
    layer0_outputs(5948) <= not (a or b);
    layer0_outputs(5949) <= not (a or b);
    layer0_outputs(5950) <= not b;
    layer0_outputs(5951) <= not a or b;
    layer0_outputs(5952) <= not b or a;
    layer0_outputs(5953) <= not (a or b);
    layer0_outputs(5954) <= b;
    layer0_outputs(5955) <= a and not b;
    layer0_outputs(5956) <= b and not a;
    layer0_outputs(5957) <= not a;
    layer0_outputs(5958) <= a;
    layer0_outputs(5959) <= 1'b0;
    layer0_outputs(5960) <= a or b;
    layer0_outputs(5961) <= b;
    layer0_outputs(5962) <= not (a or b);
    layer0_outputs(5963) <= a and not b;
    layer0_outputs(5964) <= a and not b;
    layer0_outputs(5965) <= not a;
    layer0_outputs(5966) <= not b;
    layer0_outputs(5967) <= a or b;
    layer0_outputs(5968) <= not a;
    layer0_outputs(5969) <= not b;
    layer0_outputs(5970) <= not b or a;
    layer0_outputs(5971) <= not b;
    layer0_outputs(5972) <= not a;
    layer0_outputs(5973) <= not b;
    layer0_outputs(5974) <= not (a and b);
    layer0_outputs(5975) <= a xor b;
    layer0_outputs(5976) <= not b;
    layer0_outputs(5977) <= a;
    layer0_outputs(5978) <= a or b;
    layer0_outputs(5979) <= a and not b;
    layer0_outputs(5980) <= a xor b;
    layer0_outputs(5981) <= not (a xor b);
    layer0_outputs(5982) <= a and not b;
    layer0_outputs(5983) <= a or b;
    layer0_outputs(5984) <= b and not a;
    layer0_outputs(5985) <= a or b;
    layer0_outputs(5986) <= not (a xor b);
    layer0_outputs(5987) <= not (a xor b);
    layer0_outputs(5988) <= a xor b;
    layer0_outputs(5989) <= a or b;
    layer0_outputs(5990) <= b;
    layer0_outputs(5991) <= not (a or b);
    layer0_outputs(5992) <= not (a or b);
    layer0_outputs(5993) <= a xor b;
    layer0_outputs(5994) <= a;
    layer0_outputs(5995) <= not (a xor b);
    layer0_outputs(5996) <= not a or b;
    layer0_outputs(5997) <= not (a or b);
    layer0_outputs(5998) <= a xor b;
    layer0_outputs(5999) <= a xor b;
    layer0_outputs(6000) <= b and not a;
    layer0_outputs(6001) <= 1'b1;
    layer0_outputs(6002) <= b;
    layer0_outputs(6003) <= not b or a;
    layer0_outputs(6004) <= not b;
    layer0_outputs(6005) <= not a or b;
    layer0_outputs(6006) <= a and b;
    layer0_outputs(6007) <= a or b;
    layer0_outputs(6008) <= a;
    layer0_outputs(6009) <= not b;
    layer0_outputs(6010) <= a and not b;
    layer0_outputs(6011) <= not (a and b);
    layer0_outputs(6012) <= a xor b;
    layer0_outputs(6013) <= not (a xor b);
    layer0_outputs(6014) <= not (a xor b);
    layer0_outputs(6015) <= not b;
    layer0_outputs(6016) <= a;
    layer0_outputs(6017) <= not a or b;
    layer0_outputs(6018) <= not (a or b);
    layer0_outputs(6019) <= not (a or b);
    layer0_outputs(6020) <= a or b;
    layer0_outputs(6021) <= not a or b;
    layer0_outputs(6022) <= a xor b;
    layer0_outputs(6023) <= not b;
    layer0_outputs(6024) <= 1'b1;
    layer0_outputs(6025) <= a xor b;
    layer0_outputs(6026) <= b and not a;
    layer0_outputs(6027) <= not b;
    layer0_outputs(6028) <= not (a xor b);
    layer0_outputs(6029) <= not (a or b);
    layer0_outputs(6030) <= not a;
    layer0_outputs(6031) <= not (a and b);
    layer0_outputs(6032) <= a and b;
    layer0_outputs(6033) <= a or b;
    layer0_outputs(6034) <= b;
    layer0_outputs(6035) <= not (a xor b);
    layer0_outputs(6036) <= not (a xor b);
    layer0_outputs(6037) <= 1'b1;
    layer0_outputs(6038) <= a or b;
    layer0_outputs(6039) <= not a or b;
    layer0_outputs(6040) <= a or b;
    layer0_outputs(6041) <= not b;
    layer0_outputs(6042) <= b;
    layer0_outputs(6043) <= not (a or b);
    layer0_outputs(6044) <= b and not a;
    layer0_outputs(6045) <= not a or b;
    layer0_outputs(6046) <= not b;
    layer0_outputs(6047) <= not a;
    layer0_outputs(6048) <= not (a or b);
    layer0_outputs(6049) <= b;
    layer0_outputs(6050) <= a;
    layer0_outputs(6051) <= b and not a;
    layer0_outputs(6052) <= not (a xor b);
    layer0_outputs(6053) <= not (a or b);
    layer0_outputs(6054) <= a or b;
    layer0_outputs(6055) <= a;
    layer0_outputs(6056) <= 1'b1;
    layer0_outputs(6057) <= not (a xor b);
    layer0_outputs(6058) <= a xor b;
    layer0_outputs(6059) <= not a or b;
    layer0_outputs(6060) <= a or b;
    layer0_outputs(6061) <= not (a or b);
    layer0_outputs(6062) <= not (a xor b);
    layer0_outputs(6063) <= not (a xor b);
    layer0_outputs(6064) <= not a or b;
    layer0_outputs(6065) <= not (a or b);
    layer0_outputs(6066) <= not (a or b);
    layer0_outputs(6067) <= not b;
    layer0_outputs(6068) <= not (a xor b);
    layer0_outputs(6069) <= a and not b;
    layer0_outputs(6070) <= not b;
    layer0_outputs(6071) <= a xor b;
    layer0_outputs(6072) <= not b;
    layer0_outputs(6073) <= b and not a;
    layer0_outputs(6074) <= a xor b;
    layer0_outputs(6075) <= a and not b;
    layer0_outputs(6076) <= not (a xor b);
    layer0_outputs(6077) <= not b or a;
    layer0_outputs(6078) <= not b or a;
    layer0_outputs(6079) <= not (a or b);
    layer0_outputs(6080) <= not b or a;
    layer0_outputs(6081) <= not a or b;
    layer0_outputs(6082) <= not a;
    layer0_outputs(6083) <= not a;
    layer0_outputs(6084) <= 1'b0;
    layer0_outputs(6085) <= a and b;
    layer0_outputs(6086) <= not (a or b);
    layer0_outputs(6087) <= a;
    layer0_outputs(6088) <= not b;
    layer0_outputs(6089) <= a and not b;
    layer0_outputs(6090) <= not a or b;
    layer0_outputs(6091) <= not a;
    layer0_outputs(6092) <= a or b;
    layer0_outputs(6093) <= b;
    layer0_outputs(6094) <= a or b;
    layer0_outputs(6095) <= not (a or b);
    layer0_outputs(6096) <= a xor b;
    layer0_outputs(6097) <= not (a or b);
    layer0_outputs(6098) <= not b;
    layer0_outputs(6099) <= not (a xor b);
    layer0_outputs(6100) <= not a or b;
    layer0_outputs(6101) <= a or b;
    layer0_outputs(6102) <= 1'b0;
    layer0_outputs(6103) <= a xor b;
    layer0_outputs(6104) <= not (a xor b);
    layer0_outputs(6105) <= not (a or b);
    layer0_outputs(6106) <= b and not a;
    layer0_outputs(6107) <= a or b;
    layer0_outputs(6108) <= a and not b;
    layer0_outputs(6109) <= not b or a;
    layer0_outputs(6110) <= b and not a;
    layer0_outputs(6111) <= b and not a;
    layer0_outputs(6112) <= not a;
    layer0_outputs(6113) <= a xor b;
    layer0_outputs(6114) <= a;
    layer0_outputs(6115) <= not b or a;
    layer0_outputs(6116) <= a;
    layer0_outputs(6117) <= not a or b;
    layer0_outputs(6118) <= b;
    layer0_outputs(6119) <= not a or b;
    layer0_outputs(6120) <= not (a or b);
    layer0_outputs(6121) <= b and not a;
    layer0_outputs(6122) <= b;
    layer0_outputs(6123) <= a or b;
    layer0_outputs(6124) <= not (a xor b);
    layer0_outputs(6125) <= a;
    layer0_outputs(6126) <= b;
    layer0_outputs(6127) <= not (a xor b);
    layer0_outputs(6128) <= not (a xor b);
    layer0_outputs(6129) <= a or b;
    layer0_outputs(6130) <= a xor b;
    layer0_outputs(6131) <= not (a or b);
    layer0_outputs(6132) <= a;
    layer0_outputs(6133) <= a;
    layer0_outputs(6134) <= not a;
    layer0_outputs(6135) <= not (a xor b);
    layer0_outputs(6136) <= not b;
    layer0_outputs(6137) <= 1'b1;
    layer0_outputs(6138) <= a and not b;
    layer0_outputs(6139) <= not (a and b);
    layer0_outputs(6140) <= a;
    layer0_outputs(6141) <= not b;
    layer0_outputs(6142) <= not (a or b);
    layer0_outputs(6143) <= not (a or b);
    layer0_outputs(6144) <= a or b;
    layer0_outputs(6145) <= not (a or b);
    layer0_outputs(6146) <= a xor b;
    layer0_outputs(6147) <= b and not a;
    layer0_outputs(6148) <= not b or a;
    layer0_outputs(6149) <= not (a xor b);
    layer0_outputs(6150) <= not b;
    layer0_outputs(6151) <= a or b;
    layer0_outputs(6152) <= a or b;
    layer0_outputs(6153) <= 1'b0;
    layer0_outputs(6154) <= not a;
    layer0_outputs(6155) <= not (a xor b);
    layer0_outputs(6156) <= b;
    layer0_outputs(6157) <= a and not b;
    layer0_outputs(6158) <= a or b;
    layer0_outputs(6159) <= not (a or b);
    layer0_outputs(6160) <= b and not a;
    layer0_outputs(6161) <= not a;
    layer0_outputs(6162) <= not a;
    layer0_outputs(6163) <= not (a or b);
    layer0_outputs(6164) <= not b or a;
    layer0_outputs(6165) <= a;
    layer0_outputs(6166) <= not (a or b);
    layer0_outputs(6167) <= a;
    layer0_outputs(6168) <= b and not a;
    layer0_outputs(6169) <= not (a xor b);
    layer0_outputs(6170) <= a and not b;
    layer0_outputs(6171) <= 1'b0;
    layer0_outputs(6172) <= 1'b0;
    layer0_outputs(6173) <= not (a xor b);
    layer0_outputs(6174) <= b and not a;
    layer0_outputs(6175) <= a xor b;
    layer0_outputs(6176) <= not (a or b);
    layer0_outputs(6177) <= not (a xor b);
    layer0_outputs(6178) <= a;
    layer0_outputs(6179) <= b and not a;
    layer0_outputs(6180) <= not (a and b);
    layer0_outputs(6181) <= 1'b1;
    layer0_outputs(6182) <= not (a and b);
    layer0_outputs(6183) <= not b or a;
    layer0_outputs(6184) <= 1'b1;
    layer0_outputs(6185) <= b and not a;
    layer0_outputs(6186) <= a and not b;
    layer0_outputs(6187) <= a or b;
    layer0_outputs(6188) <= not (a xor b);
    layer0_outputs(6189) <= 1'b0;
    layer0_outputs(6190) <= a and not b;
    layer0_outputs(6191) <= b and not a;
    layer0_outputs(6192) <= not b;
    layer0_outputs(6193) <= b and not a;
    layer0_outputs(6194) <= a or b;
    layer0_outputs(6195) <= not b or a;
    layer0_outputs(6196) <= a xor b;
    layer0_outputs(6197) <= a;
    layer0_outputs(6198) <= not a or b;
    layer0_outputs(6199) <= not b or a;
    layer0_outputs(6200) <= not (a xor b);
    layer0_outputs(6201) <= not (a or b);
    layer0_outputs(6202) <= not a;
    layer0_outputs(6203) <= not (a or b);
    layer0_outputs(6204) <= b and not a;
    layer0_outputs(6205) <= not b;
    layer0_outputs(6206) <= a or b;
    layer0_outputs(6207) <= a xor b;
    layer0_outputs(6208) <= b;
    layer0_outputs(6209) <= not a;
    layer0_outputs(6210) <= a or b;
    layer0_outputs(6211) <= b and not a;
    layer0_outputs(6212) <= b;
    layer0_outputs(6213) <= 1'b1;
    layer0_outputs(6214) <= a or b;
    layer0_outputs(6215) <= not b;
    layer0_outputs(6216) <= not b or a;
    layer0_outputs(6217) <= a xor b;
    layer0_outputs(6218) <= a or b;
    layer0_outputs(6219) <= a xor b;
    layer0_outputs(6220) <= not (a xor b);
    layer0_outputs(6221) <= not a;
    layer0_outputs(6222) <= not (a xor b);
    layer0_outputs(6223) <= not (a xor b);
    layer0_outputs(6224) <= a and not b;
    layer0_outputs(6225) <= a;
    layer0_outputs(6226) <= not (a xor b);
    layer0_outputs(6227) <= b and not a;
    layer0_outputs(6228) <= not (a xor b);
    layer0_outputs(6229) <= not b;
    layer0_outputs(6230) <= a xor b;
    layer0_outputs(6231) <= not a;
    layer0_outputs(6232) <= not a;
    layer0_outputs(6233) <= b;
    layer0_outputs(6234) <= not (a or b);
    layer0_outputs(6235) <= b and not a;
    layer0_outputs(6236) <= not (a xor b);
    layer0_outputs(6237) <= a xor b;
    layer0_outputs(6238) <= a xor b;
    layer0_outputs(6239) <= not (a xor b);
    layer0_outputs(6240) <= not b or a;
    layer0_outputs(6241) <= not (a or b);
    layer0_outputs(6242) <= not (a or b);
    layer0_outputs(6243) <= a and not b;
    layer0_outputs(6244) <= a and b;
    layer0_outputs(6245) <= not b;
    layer0_outputs(6246) <= not (a or b);
    layer0_outputs(6247) <= not b;
    layer0_outputs(6248) <= a;
    layer0_outputs(6249) <= not a;
    layer0_outputs(6250) <= not a or b;
    layer0_outputs(6251) <= not (a xor b);
    layer0_outputs(6252) <= not a or b;
    layer0_outputs(6253) <= b and not a;
    layer0_outputs(6254) <= not a or b;
    layer0_outputs(6255) <= 1'b0;
    layer0_outputs(6256) <= not a;
    layer0_outputs(6257) <= b;
    layer0_outputs(6258) <= a or b;
    layer0_outputs(6259) <= b;
    layer0_outputs(6260) <= not a or b;
    layer0_outputs(6261) <= not (a or b);
    layer0_outputs(6262) <= not (a xor b);
    layer0_outputs(6263) <= not a;
    layer0_outputs(6264) <= a and not b;
    layer0_outputs(6265) <= 1'b0;
    layer0_outputs(6266) <= a and not b;
    layer0_outputs(6267) <= a or b;
    layer0_outputs(6268) <= b and not a;
    layer0_outputs(6269) <= not b or a;
    layer0_outputs(6270) <= not a or b;
    layer0_outputs(6271) <= a xor b;
    layer0_outputs(6272) <= a xor b;
    layer0_outputs(6273) <= not a or b;
    layer0_outputs(6274) <= not a;
    layer0_outputs(6275) <= b and not a;
    layer0_outputs(6276) <= a;
    layer0_outputs(6277) <= 1'b1;
    layer0_outputs(6278) <= a;
    layer0_outputs(6279) <= not a;
    layer0_outputs(6280) <= not (a or b);
    layer0_outputs(6281) <= not a or b;
    layer0_outputs(6282) <= not b or a;
    layer0_outputs(6283) <= b;
    layer0_outputs(6284) <= a;
    layer0_outputs(6285) <= not a;
    layer0_outputs(6286) <= not a;
    layer0_outputs(6287) <= not b or a;
    layer0_outputs(6288) <= not (a xor b);
    layer0_outputs(6289) <= not a or b;
    layer0_outputs(6290) <= a and b;
    layer0_outputs(6291) <= a and not b;
    layer0_outputs(6292) <= 1'b0;
    layer0_outputs(6293) <= not a;
    layer0_outputs(6294) <= not (a or b);
    layer0_outputs(6295) <= not (a xor b);
    layer0_outputs(6296) <= a or b;
    layer0_outputs(6297) <= a xor b;
    layer0_outputs(6298) <= not b;
    layer0_outputs(6299) <= not a;
    layer0_outputs(6300) <= not (a or b);
    layer0_outputs(6301) <= a xor b;
    layer0_outputs(6302) <= not b;
    layer0_outputs(6303) <= not (a xor b);
    layer0_outputs(6304) <= not a or b;
    layer0_outputs(6305) <= a and not b;
    layer0_outputs(6306) <= a xor b;
    layer0_outputs(6307) <= not b;
    layer0_outputs(6308) <= a and not b;
    layer0_outputs(6309) <= 1'b0;
    layer0_outputs(6310) <= not a;
    layer0_outputs(6311) <= not a;
    layer0_outputs(6312) <= not (a xor b);
    layer0_outputs(6313) <= a xor b;
    layer0_outputs(6314) <= not a or b;
    layer0_outputs(6315) <= not (a or b);
    layer0_outputs(6316) <= not b or a;
    layer0_outputs(6317) <= a or b;
    layer0_outputs(6318) <= not (a or b);
    layer0_outputs(6319) <= a or b;
    layer0_outputs(6320) <= not (a xor b);
    layer0_outputs(6321) <= a or b;
    layer0_outputs(6322) <= a xor b;
    layer0_outputs(6323) <= a;
    layer0_outputs(6324) <= a xor b;
    layer0_outputs(6325) <= a or b;
    layer0_outputs(6326) <= a or b;
    layer0_outputs(6327) <= not b or a;
    layer0_outputs(6328) <= b;
    layer0_outputs(6329) <= not (a and b);
    layer0_outputs(6330) <= not a;
    layer0_outputs(6331) <= not a or b;
    layer0_outputs(6332) <= a and not b;
    layer0_outputs(6333) <= a and not b;
    layer0_outputs(6334) <= a;
    layer0_outputs(6335) <= b and not a;
    layer0_outputs(6336) <= not (a and b);
    layer0_outputs(6337) <= a;
    layer0_outputs(6338) <= not b or a;
    layer0_outputs(6339) <= not (a xor b);
    layer0_outputs(6340) <= 1'b1;
    layer0_outputs(6341) <= a or b;
    layer0_outputs(6342) <= not (a xor b);
    layer0_outputs(6343) <= not (a xor b);
    layer0_outputs(6344) <= not b;
    layer0_outputs(6345) <= not a or b;
    layer0_outputs(6346) <= a or b;
    layer0_outputs(6347) <= not (a or b);
    layer0_outputs(6348) <= b;
    layer0_outputs(6349) <= a or b;
    layer0_outputs(6350) <= b;
    layer0_outputs(6351) <= not b or a;
    layer0_outputs(6352) <= not b;
    layer0_outputs(6353) <= not b or a;
    layer0_outputs(6354) <= b;
    layer0_outputs(6355) <= a or b;
    layer0_outputs(6356) <= not (a xor b);
    layer0_outputs(6357) <= not (a xor b);
    layer0_outputs(6358) <= b;
    layer0_outputs(6359) <= a;
    layer0_outputs(6360) <= not (a xor b);
    layer0_outputs(6361) <= a or b;
    layer0_outputs(6362) <= not (a or b);
    layer0_outputs(6363) <= b;
    layer0_outputs(6364) <= not b or a;
    layer0_outputs(6365) <= a or b;
    layer0_outputs(6366) <= b;
    layer0_outputs(6367) <= a or b;
    layer0_outputs(6368) <= not a;
    layer0_outputs(6369) <= not b or a;
    layer0_outputs(6370) <= 1'b0;
    layer0_outputs(6371) <= not b or a;
    layer0_outputs(6372) <= a and not b;
    layer0_outputs(6373) <= a or b;
    layer0_outputs(6374) <= not (a xor b);
    layer0_outputs(6375) <= not a;
    layer0_outputs(6376) <= not (a xor b);
    layer0_outputs(6377) <= not b or a;
    layer0_outputs(6378) <= a;
    layer0_outputs(6379) <= 1'b1;
    layer0_outputs(6380) <= a and b;
    layer0_outputs(6381) <= not (a xor b);
    layer0_outputs(6382) <= not b;
    layer0_outputs(6383) <= a or b;
    layer0_outputs(6384) <= a;
    layer0_outputs(6385) <= b and not a;
    layer0_outputs(6386) <= a and b;
    layer0_outputs(6387) <= a and not b;
    layer0_outputs(6388) <= a or b;
    layer0_outputs(6389) <= not b or a;
    layer0_outputs(6390) <= a xor b;
    layer0_outputs(6391) <= a;
    layer0_outputs(6392) <= not (a or b);
    layer0_outputs(6393) <= b and not a;
    layer0_outputs(6394) <= not (a xor b);
    layer0_outputs(6395) <= a xor b;
    layer0_outputs(6396) <= b and not a;
    layer0_outputs(6397) <= not (a xor b);
    layer0_outputs(6398) <= not (a or b);
    layer0_outputs(6399) <= not (a and b);
    layer0_outputs(6400) <= not b;
    layer0_outputs(6401) <= a or b;
    layer0_outputs(6402) <= not b;
    layer0_outputs(6403) <= b;
    layer0_outputs(6404) <= 1'b0;
    layer0_outputs(6405) <= a xor b;
    layer0_outputs(6406) <= b and not a;
    layer0_outputs(6407) <= not (a xor b);
    layer0_outputs(6408) <= a;
    layer0_outputs(6409) <= not a or b;
    layer0_outputs(6410) <= b;
    layer0_outputs(6411) <= b;
    layer0_outputs(6412) <= a or b;
    layer0_outputs(6413) <= not (a xor b);
    layer0_outputs(6414) <= not b or a;
    layer0_outputs(6415) <= a;
    layer0_outputs(6416) <= a;
    layer0_outputs(6417) <= a or b;
    layer0_outputs(6418) <= not (a or b);
    layer0_outputs(6419) <= not b or a;
    layer0_outputs(6420) <= not (a xor b);
    layer0_outputs(6421) <= a or b;
    layer0_outputs(6422) <= a xor b;
    layer0_outputs(6423) <= a or b;
    layer0_outputs(6424) <= b and not a;
    layer0_outputs(6425) <= not (a or b);
    layer0_outputs(6426) <= not (a and b);
    layer0_outputs(6427) <= a and b;
    layer0_outputs(6428) <= a xor b;
    layer0_outputs(6429) <= not (a or b);
    layer0_outputs(6430) <= b;
    layer0_outputs(6431) <= not b;
    layer0_outputs(6432) <= a or b;
    layer0_outputs(6433) <= a xor b;
    layer0_outputs(6434) <= a xor b;
    layer0_outputs(6435) <= a and not b;
    layer0_outputs(6436) <= not (a or b);
    layer0_outputs(6437) <= b and not a;
    layer0_outputs(6438) <= not b or a;
    layer0_outputs(6439) <= a or b;
    layer0_outputs(6440) <= a and b;
    layer0_outputs(6441) <= not a or b;
    layer0_outputs(6442) <= b;
    layer0_outputs(6443) <= a or b;
    layer0_outputs(6444) <= a;
    layer0_outputs(6445) <= not a;
    layer0_outputs(6446) <= b and not a;
    layer0_outputs(6447) <= not (a xor b);
    layer0_outputs(6448) <= a and not b;
    layer0_outputs(6449) <= not a or b;
    layer0_outputs(6450) <= not b;
    layer0_outputs(6451) <= b and not a;
    layer0_outputs(6452) <= b;
    layer0_outputs(6453) <= not (a or b);
    layer0_outputs(6454) <= b;
    layer0_outputs(6455) <= b;
    layer0_outputs(6456) <= a xor b;
    layer0_outputs(6457) <= 1'b1;
    layer0_outputs(6458) <= not a or b;
    layer0_outputs(6459) <= b and not a;
    layer0_outputs(6460) <= not (a and b);
    layer0_outputs(6461) <= b and not a;
    layer0_outputs(6462) <= a and not b;
    layer0_outputs(6463) <= a;
    layer0_outputs(6464) <= not (a and b);
    layer0_outputs(6465) <= not (a or b);
    layer0_outputs(6466) <= not b;
    layer0_outputs(6467) <= not (a or b);
    layer0_outputs(6468) <= a or b;
    layer0_outputs(6469) <= a and not b;
    layer0_outputs(6470) <= not a;
    layer0_outputs(6471) <= a xor b;
    layer0_outputs(6472) <= not a or b;
    layer0_outputs(6473) <= a or b;
    layer0_outputs(6474) <= not (a or b);
    layer0_outputs(6475) <= not (a xor b);
    layer0_outputs(6476) <= b;
    layer0_outputs(6477) <= b and not a;
    layer0_outputs(6478) <= 1'b1;
    layer0_outputs(6479) <= b and not a;
    layer0_outputs(6480) <= a and not b;
    layer0_outputs(6481) <= b and not a;
    layer0_outputs(6482) <= a or b;
    layer0_outputs(6483) <= not a or b;
    layer0_outputs(6484) <= not (a and b);
    layer0_outputs(6485) <= b and not a;
    layer0_outputs(6486) <= not (a or b);
    layer0_outputs(6487) <= not (a xor b);
    layer0_outputs(6488) <= not (a or b);
    layer0_outputs(6489) <= not a;
    layer0_outputs(6490) <= a xor b;
    layer0_outputs(6491) <= 1'b0;
    layer0_outputs(6492) <= not (a xor b);
    layer0_outputs(6493) <= not b or a;
    layer0_outputs(6494) <= a and b;
    layer0_outputs(6495) <= not b;
    layer0_outputs(6496) <= b;
    layer0_outputs(6497) <= a xor b;
    layer0_outputs(6498) <= not (a xor b);
    layer0_outputs(6499) <= not b;
    layer0_outputs(6500) <= not a;
    layer0_outputs(6501) <= not (a xor b);
    layer0_outputs(6502) <= not b or a;
    layer0_outputs(6503) <= not (a or b);
    layer0_outputs(6504) <= not b or a;
    layer0_outputs(6505) <= a or b;
    layer0_outputs(6506) <= not (a or b);
    layer0_outputs(6507) <= not b;
    layer0_outputs(6508) <= not (a or b);
    layer0_outputs(6509) <= a and not b;
    layer0_outputs(6510) <= not a or b;
    layer0_outputs(6511) <= not b;
    layer0_outputs(6512) <= not b;
    layer0_outputs(6513) <= a and not b;
    layer0_outputs(6514) <= not (a and b);
    layer0_outputs(6515) <= not (a or b);
    layer0_outputs(6516) <= not b or a;
    layer0_outputs(6517) <= a xor b;
    layer0_outputs(6518) <= b and not a;
    layer0_outputs(6519) <= a or b;
    layer0_outputs(6520) <= not (a or b);
    layer0_outputs(6521) <= b and not a;
    layer0_outputs(6522) <= not a or b;
    layer0_outputs(6523) <= not (a and b);
    layer0_outputs(6524) <= a or b;
    layer0_outputs(6525) <= not a;
    layer0_outputs(6526) <= a xor b;
    layer0_outputs(6527) <= a or b;
    layer0_outputs(6528) <= 1'b0;
    layer0_outputs(6529) <= not (a xor b);
    layer0_outputs(6530) <= a or b;
    layer0_outputs(6531) <= a xor b;
    layer0_outputs(6532) <= not (a xor b);
    layer0_outputs(6533) <= not a;
    layer0_outputs(6534) <= not a or b;
    layer0_outputs(6535) <= a xor b;
    layer0_outputs(6536) <= a;
    layer0_outputs(6537) <= a and not b;
    layer0_outputs(6538) <= 1'b0;
    layer0_outputs(6539) <= not b;
    layer0_outputs(6540) <= a;
    layer0_outputs(6541) <= a xor b;
    layer0_outputs(6542) <= not a or b;
    layer0_outputs(6543) <= a xor b;
    layer0_outputs(6544) <= not a or b;
    layer0_outputs(6545) <= not (a or b);
    layer0_outputs(6546) <= not (a xor b);
    layer0_outputs(6547) <= a or b;
    layer0_outputs(6548) <= not (a or b);
    layer0_outputs(6549) <= not (a xor b);
    layer0_outputs(6550) <= b and not a;
    layer0_outputs(6551) <= not (a xor b);
    layer0_outputs(6552) <= not (a or b);
    layer0_outputs(6553) <= a or b;
    layer0_outputs(6554) <= a and not b;
    layer0_outputs(6555) <= not a or b;
    layer0_outputs(6556) <= b;
    layer0_outputs(6557) <= not a or b;
    layer0_outputs(6558) <= not (a xor b);
    layer0_outputs(6559) <= 1'b1;
    layer0_outputs(6560) <= not a;
    layer0_outputs(6561) <= not (a and b);
    layer0_outputs(6562) <= a xor b;
    layer0_outputs(6563) <= not (a xor b);
    layer0_outputs(6564) <= 1'b0;
    layer0_outputs(6565) <= a xor b;
    layer0_outputs(6566) <= b;
    layer0_outputs(6567) <= 1'b1;
    layer0_outputs(6568) <= not (a or b);
    layer0_outputs(6569) <= 1'b0;
    layer0_outputs(6570) <= b and not a;
    layer0_outputs(6571) <= a xor b;
    layer0_outputs(6572) <= a and not b;
    layer0_outputs(6573) <= a or b;
    layer0_outputs(6574) <= a;
    layer0_outputs(6575) <= not a;
    layer0_outputs(6576) <= a;
    layer0_outputs(6577) <= not (a or b);
    layer0_outputs(6578) <= not a or b;
    layer0_outputs(6579) <= not b;
    layer0_outputs(6580) <= a and not b;
    layer0_outputs(6581) <= b;
    layer0_outputs(6582) <= not (a xor b);
    layer0_outputs(6583) <= a and b;
    layer0_outputs(6584) <= not a;
    layer0_outputs(6585) <= a;
    layer0_outputs(6586) <= not (a xor b);
    layer0_outputs(6587) <= a and not b;
    layer0_outputs(6588) <= not b;
    layer0_outputs(6589) <= a or b;
    layer0_outputs(6590) <= a and not b;
    layer0_outputs(6591) <= not a or b;
    layer0_outputs(6592) <= not (a and b);
    layer0_outputs(6593) <= not (a xor b);
    layer0_outputs(6594) <= not b;
    layer0_outputs(6595) <= b;
    layer0_outputs(6596) <= not a or b;
    layer0_outputs(6597) <= a or b;
    layer0_outputs(6598) <= a or b;
    layer0_outputs(6599) <= a or b;
    layer0_outputs(6600) <= not (a xor b);
    layer0_outputs(6601) <= not a;
    layer0_outputs(6602) <= a xor b;
    layer0_outputs(6603) <= a and not b;
    layer0_outputs(6604) <= b;
    layer0_outputs(6605) <= 1'b0;
    layer0_outputs(6606) <= not a or b;
    layer0_outputs(6607) <= a or b;
    layer0_outputs(6608) <= a xor b;
    layer0_outputs(6609) <= not b or a;
    layer0_outputs(6610) <= not a;
    layer0_outputs(6611) <= not b or a;
    layer0_outputs(6612) <= not b or a;
    layer0_outputs(6613) <= not b;
    layer0_outputs(6614) <= not b or a;
    layer0_outputs(6615) <= not b;
    layer0_outputs(6616) <= not (a xor b);
    layer0_outputs(6617) <= a xor b;
    layer0_outputs(6618) <= b and not a;
    layer0_outputs(6619) <= not (a or b);
    layer0_outputs(6620) <= a and not b;
    layer0_outputs(6621) <= a xor b;
    layer0_outputs(6622) <= not (a xor b);
    layer0_outputs(6623) <= not (a and b);
    layer0_outputs(6624) <= not b or a;
    layer0_outputs(6625) <= a xor b;
    layer0_outputs(6626) <= not (a or b);
    layer0_outputs(6627) <= not (a or b);
    layer0_outputs(6628) <= not b or a;
    layer0_outputs(6629) <= b;
    layer0_outputs(6630) <= a and not b;
    layer0_outputs(6631) <= not b;
    layer0_outputs(6632) <= a or b;
    layer0_outputs(6633) <= 1'b0;
    layer0_outputs(6634) <= not (a xor b);
    layer0_outputs(6635) <= a and b;
    layer0_outputs(6636) <= not (a or b);
    layer0_outputs(6637) <= 1'b0;
    layer0_outputs(6638) <= 1'b0;
    layer0_outputs(6639) <= a and not b;
    layer0_outputs(6640) <= a or b;
    layer0_outputs(6641) <= b;
    layer0_outputs(6642) <= not b or a;
    layer0_outputs(6643) <= b;
    layer0_outputs(6644) <= not (a and b);
    layer0_outputs(6645) <= not a;
    layer0_outputs(6646) <= a and not b;
    layer0_outputs(6647) <= not (a xor b);
    layer0_outputs(6648) <= b and not a;
    layer0_outputs(6649) <= a or b;
    layer0_outputs(6650) <= b and not a;
    layer0_outputs(6651) <= a or b;
    layer0_outputs(6652) <= a xor b;
    layer0_outputs(6653) <= a xor b;
    layer0_outputs(6654) <= not b;
    layer0_outputs(6655) <= a;
    layer0_outputs(6656) <= not (a xor b);
    layer0_outputs(6657) <= a;
    layer0_outputs(6658) <= a or b;
    layer0_outputs(6659) <= not (a or b);
    layer0_outputs(6660) <= a xor b;
    layer0_outputs(6661) <= not a;
    layer0_outputs(6662) <= a;
    layer0_outputs(6663) <= a xor b;
    layer0_outputs(6664) <= b and not a;
    layer0_outputs(6665) <= b and not a;
    layer0_outputs(6666) <= a and b;
    layer0_outputs(6667) <= not b;
    layer0_outputs(6668) <= not (a or b);
    layer0_outputs(6669) <= not a or b;
    layer0_outputs(6670) <= not (a xor b);
    layer0_outputs(6671) <= not b or a;
    layer0_outputs(6672) <= a xor b;
    layer0_outputs(6673) <= a xor b;
    layer0_outputs(6674) <= not b or a;
    layer0_outputs(6675) <= a or b;
    layer0_outputs(6676) <= a or b;
    layer0_outputs(6677) <= not a;
    layer0_outputs(6678) <= a and b;
    layer0_outputs(6679) <= a or b;
    layer0_outputs(6680) <= 1'b0;
    layer0_outputs(6681) <= a xor b;
    layer0_outputs(6682) <= a;
    layer0_outputs(6683) <= not a or b;
    layer0_outputs(6684) <= not (a or b);
    layer0_outputs(6685) <= b;
    layer0_outputs(6686) <= a and not b;
    layer0_outputs(6687) <= b and not a;
    layer0_outputs(6688) <= a and b;
    layer0_outputs(6689) <= not (a or b);
    layer0_outputs(6690) <= not a;
    layer0_outputs(6691) <= b and not a;
    layer0_outputs(6692) <= not (a xor b);
    layer0_outputs(6693) <= b;
    layer0_outputs(6694) <= not b;
    layer0_outputs(6695) <= b and not a;
    layer0_outputs(6696) <= a and b;
    layer0_outputs(6697) <= not (a or b);
    layer0_outputs(6698) <= not (a xor b);
    layer0_outputs(6699) <= not (a xor b);
    layer0_outputs(6700) <= a or b;
    layer0_outputs(6701) <= b;
    layer0_outputs(6702) <= not (a or b);
    layer0_outputs(6703) <= b;
    layer0_outputs(6704) <= not (a or b);
    layer0_outputs(6705) <= not (a xor b);
    layer0_outputs(6706) <= a and not b;
    layer0_outputs(6707) <= not (a xor b);
    layer0_outputs(6708) <= not (a or b);
    layer0_outputs(6709) <= not a or b;
    layer0_outputs(6710) <= a and not b;
    layer0_outputs(6711) <= not a;
    layer0_outputs(6712) <= a or b;
    layer0_outputs(6713) <= not (a or b);
    layer0_outputs(6714) <= not (a xor b);
    layer0_outputs(6715) <= not b or a;
    layer0_outputs(6716) <= not b;
    layer0_outputs(6717) <= not (a xor b);
    layer0_outputs(6718) <= not b or a;
    layer0_outputs(6719) <= a and b;
    layer0_outputs(6720) <= not (a or b);
    layer0_outputs(6721) <= a or b;
    layer0_outputs(6722) <= a or b;
    layer0_outputs(6723) <= 1'b1;
    layer0_outputs(6724) <= a;
    layer0_outputs(6725) <= not (a xor b);
    layer0_outputs(6726) <= a;
    layer0_outputs(6727) <= not a;
    layer0_outputs(6728) <= not b;
    layer0_outputs(6729) <= not (a xor b);
    layer0_outputs(6730) <= b;
    layer0_outputs(6731) <= not a;
    layer0_outputs(6732) <= a xor b;
    layer0_outputs(6733) <= a and b;
    layer0_outputs(6734) <= b;
    layer0_outputs(6735) <= not a;
    layer0_outputs(6736) <= not (a or b);
    layer0_outputs(6737) <= 1'b1;
    layer0_outputs(6738) <= b;
    layer0_outputs(6739) <= not (a or b);
    layer0_outputs(6740) <= not b;
    layer0_outputs(6741) <= not (a and b);
    layer0_outputs(6742) <= not b or a;
    layer0_outputs(6743) <= 1'b1;
    layer0_outputs(6744) <= a xor b;
    layer0_outputs(6745) <= b;
    layer0_outputs(6746) <= b and not a;
    layer0_outputs(6747) <= not b or a;
    layer0_outputs(6748) <= a and not b;
    layer0_outputs(6749) <= b and not a;
    layer0_outputs(6750) <= not a;
    layer0_outputs(6751) <= not (a or b);
    layer0_outputs(6752) <= 1'b0;
    layer0_outputs(6753) <= not a or b;
    layer0_outputs(6754) <= not (a xor b);
    layer0_outputs(6755) <= not (a xor b);
    layer0_outputs(6756) <= not (a xor b);
    layer0_outputs(6757) <= not b;
    layer0_outputs(6758) <= a or b;
    layer0_outputs(6759) <= not b or a;
    layer0_outputs(6760) <= 1'b0;
    layer0_outputs(6761) <= not b or a;
    layer0_outputs(6762) <= not b;
    layer0_outputs(6763) <= not a;
    layer0_outputs(6764) <= not a or b;
    layer0_outputs(6765) <= b and not a;
    layer0_outputs(6766) <= b and not a;
    layer0_outputs(6767) <= a xor b;
    layer0_outputs(6768) <= not b;
    layer0_outputs(6769) <= not (a xor b);
    layer0_outputs(6770) <= not b;
    layer0_outputs(6771) <= not (a or b);
    layer0_outputs(6772) <= not (a xor b);
    layer0_outputs(6773) <= a xor b;
    layer0_outputs(6774) <= not (a or b);
    layer0_outputs(6775) <= not b or a;
    layer0_outputs(6776) <= a and b;
    layer0_outputs(6777) <= a and b;
    layer0_outputs(6778) <= b and not a;
    layer0_outputs(6779) <= a;
    layer0_outputs(6780) <= a;
    layer0_outputs(6781) <= not a;
    layer0_outputs(6782) <= not (a xor b);
    layer0_outputs(6783) <= b and not a;
    layer0_outputs(6784) <= not b or a;
    layer0_outputs(6785) <= a or b;
    layer0_outputs(6786) <= not b;
    layer0_outputs(6787) <= not (a or b);
    layer0_outputs(6788) <= not b or a;
    layer0_outputs(6789) <= a and b;
    layer0_outputs(6790) <= not (a or b);
    layer0_outputs(6791) <= not a;
    layer0_outputs(6792) <= not (a or b);
    layer0_outputs(6793) <= not (a or b);
    layer0_outputs(6794) <= not (a and b);
    layer0_outputs(6795) <= b;
    layer0_outputs(6796) <= a and b;
    layer0_outputs(6797) <= not (a or b);
    layer0_outputs(6798) <= a xor b;
    layer0_outputs(6799) <= not (a xor b);
    layer0_outputs(6800) <= a or b;
    layer0_outputs(6801) <= 1'b0;
    layer0_outputs(6802) <= a;
    layer0_outputs(6803) <= not b or a;
    layer0_outputs(6804) <= a and b;
    layer0_outputs(6805) <= b and not a;
    layer0_outputs(6806) <= 1'b0;
    layer0_outputs(6807) <= a xor b;
    layer0_outputs(6808) <= not b;
    layer0_outputs(6809) <= not (a xor b);
    layer0_outputs(6810) <= a or b;
    layer0_outputs(6811) <= not (a xor b);
    layer0_outputs(6812) <= not (a or b);
    layer0_outputs(6813) <= not (a or b);
    layer0_outputs(6814) <= b and not a;
    layer0_outputs(6815) <= not (a xor b);
    layer0_outputs(6816) <= not a;
    layer0_outputs(6817) <= a xor b;
    layer0_outputs(6818) <= b;
    layer0_outputs(6819) <= not (a or b);
    layer0_outputs(6820) <= a or b;
    layer0_outputs(6821) <= b;
    layer0_outputs(6822) <= not a;
    layer0_outputs(6823) <= not (a xor b);
    layer0_outputs(6824) <= 1'b0;
    layer0_outputs(6825) <= not b or a;
    layer0_outputs(6826) <= not b;
    layer0_outputs(6827) <= b and not a;
    layer0_outputs(6828) <= not a or b;
    layer0_outputs(6829) <= not (a xor b);
    layer0_outputs(6830) <= a xor b;
    layer0_outputs(6831) <= a xor b;
    layer0_outputs(6832) <= not (a or b);
    layer0_outputs(6833) <= a and not b;
    layer0_outputs(6834) <= not (a or b);
    layer0_outputs(6835) <= a xor b;
    layer0_outputs(6836) <= a or b;
    layer0_outputs(6837) <= not (a or b);
    layer0_outputs(6838) <= a or b;
    layer0_outputs(6839) <= not (a or b);
    layer0_outputs(6840) <= not a or b;
    layer0_outputs(6841) <= a or b;
    layer0_outputs(6842) <= a and not b;
    layer0_outputs(6843) <= not (a xor b);
    layer0_outputs(6844) <= a xor b;
    layer0_outputs(6845) <= not (a xor b);
    layer0_outputs(6846) <= b and not a;
    layer0_outputs(6847) <= a;
    layer0_outputs(6848) <= a xor b;
    layer0_outputs(6849) <= not a or b;
    layer0_outputs(6850) <= not b;
    layer0_outputs(6851) <= b and not a;
    layer0_outputs(6852) <= a xor b;
    layer0_outputs(6853) <= not (a or b);
    layer0_outputs(6854) <= not b;
    layer0_outputs(6855) <= a and not b;
    layer0_outputs(6856) <= not a or b;
    layer0_outputs(6857) <= b;
    layer0_outputs(6858) <= 1'b0;
    layer0_outputs(6859) <= a or b;
    layer0_outputs(6860) <= not b;
    layer0_outputs(6861) <= not a or b;
    layer0_outputs(6862) <= not b;
    layer0_outputs(6863) <= not a or b;
    layer0_outputs(6864) <= a xor b;
    layer0_outputs(6865) <= a or b;
    layer0_outputs(6866) <= 1'b0;
    layer0_outputs(6867) <= not (a xor b);
    layer0_outputs(6868) <= a or b;
    layer0_outputs(6869) <= not (a or b);
    layer0_outputs(6870) <= a xor b;
    layer0_outputs(6871) <= a and not b;
    layer0_outputs(6872) <= not (a or b);
    layer0_outputs(6873) <= not b or a;
    layer0_outputs(6874) <= not (a xor b);
    layer0_outputs(6875) <= b and not a;
    layer0_outputs(6876) <= b;
    layer0_outputs(6877) <= not (a and b);
    layer0_outputs(6878) <= not a or b;
    layer0_outputs(6879) <= a or b;
    layer0_outputs(6880) <= not (a xor b);
    layer0_outputs(6881) <= a xor b;
    layer0_outputs(6882) <= not (a and b);
    layer0_outputs(6883) <= not b or a;
    layer0_outputs(6884) <= a or b;
    layer0_outputs(6885) <= 1'b1;
    layer0_outputs(6886) <= not (a and b);
    layer0_outputs(6887) <= a;
    layer0_outputs(6888) <= a xor b;
    layer0_outputs(6889) <= not b;
    layer0_outputs(6890) <= a or b;
    layer0_outputs(6891) <= not a or b;
    layer0_outputs(6892) <= a xor b;
    layer0_outputs(6893) <= b and not a;
    layer0_outputs(6894) <= not b;
    layer0_outputs(6895) <= not a or b;
    layer0_outputs(6896) <= a or b;
    layer0_outputs(6897) <= a and not b;
    layer0_outputs(6898) <= 1'b1;
    layer0_outputs(6899) <= a and not b;
    layer0_outputs(6900) <= not a;
    layer0_outputs(6901) <= a or b;
    layer0_outputs(6902) <= not a;
    layer0_outputs(6903) <= not (a or b);
    layer0_outputs(6904) <= not b or a;
    layer0_outputs(6905) <= not (a or b);
    layer0_outputs(6906) <= b;
    layer0_outputs(6907) <= not b or a;
    layer0_outputs(6908) <= not b;
    layer0_outputs(6909) <= not (a xor b);
    layer0_outputs(6910) <= not (a or b);
    layer0_outputs(6911) <= not (a xor b);
    layer0_outputs(6912) <= a or b;
    layer0_outputs(6913) <= not (a xor b);
    layer0_outputs(6914) <= a and not b;
    layer0_outputs(6915) <= 1'b0;
    layer0_outputs(6916) <= a or b;
    layer0_outputs(6917) <= a xor b;
    layer0_outputs(6918) <= b and not a;
    layer0_outputs(6919) <= not (a or b);
    layer0_outputs(6920) <= a or b;
    layer0_outputs(6921) <= not a;
    layer0_outputs(6922) <= a or b;
    layer0_outputs(6923) <= a or b;
    layer0_outputs(6924) <= not (a or b);
    layer0_outputs(6925) <= not (a or b);
    layer0_outputs(6926) <= not b or a;
    layer0_outputs(6927) <= a or b;
    layer0_outputs(6928) <= not b;
    layer0_outputs(6929) <= a xor b;
    layer0_outputs(6930) <= a or b;
    layer0_outputs(6931) <= a and not b;
    layer0_outputs(6932) <= not (a xor b);
    layer0_outputs(6933) <= a;
    layer0_outputs(6934) <= not (a xor b);
    layer0_outputs(6935) <= not (a xor b);
    layer0_outputs(6936) <= not (a xor b);
    layer0_outputs(6937) <= not (a or b);
    layer0_outputs(6938) <= a xor b;
    layer0_outputs(6939) <= not a or b;
    layer0_outputs(6940) <= not a or b;
    layer0_outputs(6941) <= not (a and b);
    layer0_outputs(6942) <= not b or a;
    layer0_outputs(6943) <= b and not a;
    layer0_outputs(6944) <= a and b;
    layer0_outputs(6945) <= not (a or b);
    layer0_outputs(6946) <= b and not a;
    layer0_outputs(6947) <= not b or a;
    layer0_outputs(6948) <= not b;
    layer0_outputs(6949) <= not (a and b);
    layer0_outputs(6950) <= a;
    layer0_outputs(6951) <= b;
    layer0_outputs(6952) <= not b;
    layer0_outputs(6953) <= not (a or b);
    layer0_outputs(6954) <= b and not a;
    layer0_outputs(6955) <= not b or a;
    layer0_outputs(6956) <= not a;
    layer0_outputs(6957) <= not a;
    layer0_outputs(6958) <= not a;
    layer0_outputs(6959) <= not a;
    layer0_outputs(6960) <= a and not b;
    layer0_outputs(6961) <= a or b;
    layer0_outputs(6962) <= a or b;
    layer0_outputs(6963) <= not (a xor b);
    layer0_outputs(6964) <= not (a or b);
    layer0_outputs(6965) <= not a;
    layer0_outputs(6966) <= not b;
    layer0_outputs(6967) <= not b;
    layer0_outputs(6968) <= not b;
    layer0_outputs(6969) <= a or b;
    layer0_outputs(6970) <= a or b;
    layer0_outputs(6971) <= a or b;
    layer0_outputs(6972) <= a or b;
    layer0_outputs(6973) <= not (a or b);
    layer0_outputs(6974) <= not (a xor b);
    layer0_outputs(6975) <= b and not a;
    layer0_outputs(6976) <= b;
    layer0_outputs(6977) <= b and not a;
    layer0_outputs(6978) <= a xor b;
    layer0_outputs(6979) <= not (a xor b);
    layer0_outputs(6980) <= a xor b;
    layer0_outputs(6981) <= a xor b;
    layer0_outputs(6982) <= a;
    layer0_outputs(6983) <= not b or a;
    layer0_outputs(6984) <= a and b;
    layer0_outputs(6985) <= not (a xor b);
    layer0_outputs(6986) <= a xor b;
    layer0_outputs(6987) <= a or b;
    layer0_outputs(6988) <= a xor b;
    layer0_outputs(6989) <= a or b;
    layer0_outputs(6990) <= not a;
    layer0_outputs(6991) <= not a or b;
    layer0_outputs(6992) <= a;
    layer0_outputs(6993) <= b;
    layer0_outputs(6994) <= a;
    layer0_outputs(6995) <= not (a or b);
    layer0_outputs(6996) <= b and not a;
    layer0_outputs(6997) <= not (a or b);
    layer0_outputs(6998) <= a xor b;
    layer0_outputs(6999) <= a or b;
    layer0_outputs(7000) <= not a;
    layer0_outputs(7001) <= 1'b1;
    layer0_outputs(7002) <= a xor b;
    layer0_outputs(7003) <= not b or a;
    layer0_outputs(7004) <= a xor b;
    layer0_outputs(7005) <= not a or b;
    layer0_outputs(7006) <= a xor b;
    layer0_outputs(7007) <= not (a or b);
    layer0_outputs(7008) <= not b or a;
    layer0_outputs(7009) <= a or b;
    layer0_outputs(7010) <= not (a xor b);
    layer0_outputs(7011) <= a;
    layer0_outputs(7012) <= not (a xor b);
    layer0_outputs(7013) <= b;
    layer0_outputs(7014) <= not (a or b);
    layer0_outputs(7015) <= a and b;
    layer0_outputs(7016) <= not b;
    layer0_outputs(7017) <= not a;
    layer0_outputs(7018) <= a or b;
    layer0_outputs(7019) <= 1'b0;
    layer0_outputs(7020) <= a or b;
    layer0_outputs(7021) <= not (a and b);
    layer0_outputs(7022) <= b;
    layer0_outputs(7023) <= b and not a;
    layer0_outputs(7024) <= not a or b;
    layer0_outputs(7025) <= not (a xor b);
    layer0_outputs(7026) <= not (a xor b);
    layer0_outputs(7027) <= not a;
    layer0_outputs(7028) <= b and not a;
    layer0_outputs(7029) <= a or b;
    layer0_outputs(7030) <= a and b;
    layer0_outputs(7031) <= not (a xor b);
    layer0_outputs(7032) <= a or b;
    layer0_outputs(7033) <= not a;
    layer0_outputs(7034) <= not (a xor b);
    layer0_outputs(7035) <= not (a xor b);
    layer0_outputs(7036) <= not a or b;
    layer0_outputs(7037) <= not (a xor b);
    layer0_outputs(7038) <= not a;
    layer0_outputs(7039) <= a and b;
    layer0_outputs(7040) <= a xor b;
    layer0_outputs(7041) <= b;
    layer0_outputs(7042) <= a or b;
    layer0_outputs(7043) <= a;
    layer0_outputs(7044) <= not (a xor b);
    layer0_outputs(7045) <= not b;
    layer0_outputs(7046) <= not (a xor b);
    layer0_outputs(7047) <= a xor b;
    layer0_outputs(7048) <= not a;
    layer0_outputs(7049) <= a xor b;
    layer0_outputs(7050) <= b and not a;
    layer0_outputs(7051) <= not a or b;
    layer0_outputs(7052) <= b;
    layer0_outputs(7053) <= a and not b;
    layer0_outputs(7054) <= a or b;
    layer0_outputs(7055) <= a;
    layer0_outputs(7056) <= b and not a;
    layer0_outputs(7057) <= a xor b;
    layer0_outputs(7058) <= b;
    layer0_outputs(7059) <= not b;
    layer0_outputs(7060) <= not (a xor b);
    layer0_outputs(7061) <= a;
    layer0_outputs(7062) <= a xor b;
    layer0_outputs(7063) <= a and not b;
    layer0_outputs(7064) <= not (a or b);
    layer0_outputs(7065) <= b and not a;
    layer0_outputs(7066) <= not a or b;
    layer0_outputs(7067) <= b;
    layer0_outputs(7068) <= a or b;
    layer0_outputs(7069) <= not a;
    layer0_outputs(7070) <= not a;
    layer0_outputs(7071) <= a or b;
    layer0_outputs(7072) <= not b;
    layer0_outputs(7073) <= not b;
    layer0_outputs(7074) <= b and not a;
    layer0_outputs(7075) <= a or b;
    layer0_outputs(7076) <= not a;
    layer0_outputs(7077) <= a xor b;
    layer0_outputs(7078) <= not b or a;
    layer0_outputs(7079) <= not b;
    layer0_outputs(7080) <= a and not b;
    layer0_outputs(7081) <= not b;
    layer0_outputs(7082) <= a and not b;
    layer0_outputs(7083) <= b;
    layer0_outputs(7084) <= not (a and b);
    layer0_outputs(7085) <= not (a or b);
    layer0_outputs(7086) <= not a;
    layer0_outputs(7087) <= a and b;
    layer0_outputs(7088) <= not (a or b);
    layer0_outputs(7089) <= not a;
    layer0_outputs(7090) <= not (a xor b);
    layer0_outputs(7091) <= b and not a;
    layer0_outputs(7092) <= not (a or b);
    layer0_outputs(7093) <= not (a or b);
    layer0_outputs(7094) <= a xor b;
    layer0_outputs(7095) <= 1'b0;
    layer0_outputs(7096) <= a;
    layer0_outputs(7097) <= not (a or b);
    layer0_outputs(7098) <= not a;
    layer0_outputs(7099) <= not b or a;
    layer0_outputs(7100) <= b;
    layer0_outputs(7101) <= not (a or b);
    layer0_outputs(7102) <= a;
    layer0_outputs(7103) <= not b;
    layer0_outputs(7104) <= a or b;
    layer0_outputs(7105) <= b and not a;
    layer0_outputs(7106) <= b;
    layer0_outputs(7107) <= not (a and b);
    layer0_outputs(7108) <= b and not a;
    layer0_outputs(7109) <= 1'b1;
    layer0_outputs(7110) <= a and not b;
    layer0_outputs(7111) <= a;
    layer0_outputs(7112) <= b and not a;
    layer0_outputs(7113) <= not b;
    layer0_outputs(7114) <= a xor b;
    layer0_outputs(7115) <= not (a or b);
    layer0_outputs(7116) <= a or b;
    layer0_outputs(7117) <= not b;
    layer0_outputs(7118) <= a xor b;
    layer0_outputs(7119) <= a or b;
    layer0_outputs(7120) <= a or b;
    layer0_outputs(7121) <= a xor b;
    layer0_outputs(7122) <= b;
    layer0_outputs(7123) <= a xor b;
    layer0_outputs(7124) <= a and not b;
    layer0_outputs(7125) <= not b;
    layer0_outputs(7126) <= not b;
    layer0_outputs(7127) <= not a;
    layer0_outputs(7128) <= not (a xor b);
    layer0_outputs(7129) <= not a;
    layer0_outputs(7130) <= not b;
    layer0_outputs(7131) <= not b;
    layer0_outputs(7132) <= not (a or b);
    layer0_outputs(7133) <= not (a xor b);
    layer0_outputs(7134) <= b and not a;
    layer0_outputs(7135) <= not b;
    layer0_outputs(7136) <= not a or b;
    layer0_outputs(7137) <= not b or a;
    layer0_outputs(7138) <= b;
    layer0_outputs(7139) <= not a;
    layer0_outputs(7140) <= a xor b;
    layer0_outputs(7141) <= not b;
    layer0_outputs(7142) <= a or b;
    layer0_outputs(7143) <= not (a xor b);
    layer0_outputs(7144) <= not a or b;
    layer0_outputs(7145) <= 1'b0;
    layer0_outputs(7146) <= not (a or b);
    layer0_outputs(7147) <= a;
    layer0_outputs(7148) <= not b;
    layer0_outputs(7149) <= not (a or b);
    layer0_outputs(7150) <= not (a and b);
    layer0_outputs(7151) <= not (a xor b);
    layer0_outputs(7152) <= not (a xor b);
    layer0_outputs(7153) <= a or b;
    layer0_outputs(7154) <= not a;
    layer0_outputs(7155) <= not (a or b);
    layer0_outputs(7156) <= not (a xor b);
    layer0_outputs(7157) <= not (a xor b);
    layer0_outputs(7158) <= not (a xor b);
    layer0_outputs(7159) <= not (a and b);
    layer0_outputs(7160) <= a xor b;
    layer0_outputs(7161) <= a or b;
    layer0_outputs(7162) <= not (a xor b);
    layer0_outputs(7163) <= not (a xor b);
    layer0_outputs(7164) <= a;
    layer0_outputs(7165) <= a xor b;
    layer0_outputs(7166) <= not a or b;
    layer0_outputs(7167) <= a xor b;
    layer0_outputs(7168) <= a;
    layer0_outputs(7169) <= not a;
    layer0_outputs(7170) <= b and not a;
    layer0_outputs(7171) <= not (a or b);
    layer0_outputs(7172) <= a and not b;
    layer0_outputs(7173) <= a xor b;
    layer0_outputs(7174) <= a or b;
    layer0_outputs(7175) <= 1'b0;
    layer0_outputs(7176) <= b and not a;
    layer0_outputs(7177) <= a and not b;
    layer0_outputs(7178) <= not a or b;
    layer0_outputs(7179) <= not (a xor b);
    layer0_outputs(7180) <= not b;
    layer0_outputs(7181) <= b;
    layer0_outputs(7182) <= not a or b;
    layer0_outputs(7183) <= a and not b;
    layer0_outputs(7184) <= not a;
    layer0_outputs(7185) <= b;
    layer0_outputs(7186) <= a and not b;
    layer0_outputs(7187) <= not (a or b);
    layer0_outputs(7188) <= a or b;
    layer0_outputs(7189) <= a and not b;
    layer0_outputs(7190) <= not (a or b);
    layer0_outputs(7191) <= a or b;
    layer0_outputs(7192) <= 1'b0;
    layer0_outputs(7193) <= not a or b;
    layer0_outputs(7194) <= not (a xor b);
    layer0_outputs(7195) <= not a;
    layer0_outputs(7196) <= a and not b;
    layer0_outputs(7197) <= a or b;
    layer0_outputs(7198) <= a or b;
    layer0_outputs(7199) <= not b;
    layer0_outputs(7200) <= not (a or b);
    layer0_outputs(7201) <= not (a xor b);
    layer0_outputs(7202) <= not (a or b);
    layer0_outputs(7203) <= a or b;
    layer0_outputs(7204) <= not b or a;
    layer0_outputs(7205) <= not (a and b);
    layer0_outputs(7206) <= b and not a;
    layer0_outputs(7207) <= not a;
    layer0_outputs(7208) <= not (a or b);
    layer0_outputs(7209) <= 1'b0;
    layer0_outputs(7210) <= not (a or b);
    layer0_outputs(7211) <= not (a xor b);
    layer0_outputs(7212) <= not (a xor b);
    layer0_outputs(7213) <= not (a and b);
    layer0_outputs(7214) <= not b;
    layer0_outputs(7215) <= b and not a;
    layer0_outputs(7216) <= a xor b;
    layer0_outputs(7217) <= b;
    layer0_outputs(7218) <= a or b;
    layer0_outputs(7219) <= a xor b;
    layer0_outputs(7220) <= not (a xor b);
    layer0_outputs(7221) <= a and not b;
    layer0_outputs(7222) <= a xor b;
    layer0_outputs(7223) <= not a;
    layer0_outputs(7224) <= not a;
    layer0_outputs(7225) <= not b;
    layer0_outputs(7226) <= not a;
    layer0_outputs(7227) <= not (a or b);
    layer0_outputs(7228) <= b;
    layer0_outputs(7229) <= b;
    layer0_outputs(7230) <= not a;
    layer0_outputs(7231) <= a;
    layer0_outputs(7232) <= not b or a;
    layer0_outputs(7233) <= not (a or b);
    layer0_outputs(7234) <= not (a or b);
    layer0_outputs(7235) <= b and not a;
    layer0_outputs(7236) <= b;
    layer0_outputs(7237) <= a or b;
    layer0_outputs(7238) <= a and not b;
    layer0_outputs(7239) <= a;
    layer0_outputs(7240) <= not (a xor b);
    layer0_outputs(7241) <= not (a xor b);
    layer0_outputs(7242) <= not a;
    layer0_outputs(7243) <= not b or a;
    layer0_outputs(7244) <= b and not a;
    layer0_outputs(7245) <= a and not b;
    layer0_outputs(7246) <= not a or b;
    layer0_outputs(7247) <= not a;
    layer0_outputs(7248) <= not a or b;
    layer0_outputs(7249) <= not a or b;
    layer0_outputs(7250) <= not (a xor b);
    layer0_outputs(7251) <= not (a or b);
    layer0_outputs(7252) <= not (a or b);
    layer0_outputs(7253) <= a xor b;
    layer0_outputs(7254) <= not (a xor b);
    layer0_outputs(7255) <= not (a or b);
    layer0_outputs(7256) <= not (a xor b);
    layer0_outputs(7257) <= a or b;
    layer0_outputs(7258) <= a xor b;
    layer0_outputs(7259) <= b and not a;
    layer0_outputs(7260) <= not (a or b);
    layer0_outputs(7261) <= 1'b1;
    layer0_outputs(7262) <= not b or a;
    layer0_outputs(7263) <= not (a xor b);
    layer0_outputs(7264) <= not (a xor b);
    layer0_outputs(7265) <= b;
    layer0_outputs(7266) <= not (a xor b);
    layer0_outputs(7267) <= a or b;
    layer0_outputs(7268) <= not (a xor b);
    layer0_outputs(7269) <= not (a or b);
    layer0_outputs(7270) <= not (a or b);
    layer0_outputs(7271) <= not (a and b);
    layer0_outputs(7272) <= a and not b;
    layer0_outputs(7273) <= not (a xor b);
    layer0_outputs(7274) <= not (a xor b);
    layer0_outputs(7275) <= a or b;
    layer0_outputs(7276) <= not a or b;
    layer0_outputs(7277) <= a or b;
    layer0_outputs(7278) <= not (a or b);
    layer0_outputs(7279) <= a or b;
    layer0_outputs(7280) <= not b or a;
    layer0_outputs(7281) <= a or b;
    layer0_outputs(7282) <= a xor b;
    layer0_outputs(7283) <= a and not b;
    layer0_outputs(7284) <= a or b;
    layer0_outputs(7285) <= a or b;
    layer0_outputs(7286) <= not b;
    layer0_outputs(7287) <= not b;
    layer0_outputs(7288) <= not a or b;
    layer0_outputs(7289) <= not a or b;
    layer0_outputs(7290) <= not (a xor b);
    layer0_outputs(7291) <= not b;
    layer0_outputs(7292) <= b;
    layer0_outputs(7293) <= not (a xor b);
    layer0_outputs(7294) <= a;
    layer0_outputs(7295) <= a xor b;
    layer0_outputs(7296) <= 1'b1;
    layer0_outputs(7297) <= not a;
    layer0_outputs(7298) <= not a or b;
    layer0_outputs(7299) <= not b or a;
    layer0_outputs(7300) <= a xor b;
    layer0_outputs(7301) <= not (a or b);
    layer0_outputs(7302) <= b and not a;
    layer0_outputs(7303) <= not (a or b);
    layer0_outputs(7304) <= a or b;
    layer0_outputs(7305) <= a xor b;
    layer0_outputs(7306) <= a or b;
    layer0_outputs(7307) <= a and not b;
    layer0_outputs(7308) <= a or b;
    layer0_outputs(7309) <= not b or a;
    layer0_outputs(7310) <= not (a or b);
    layer0_outputs(7311) <= not a or b;
    layer0_outputs(7312) <= not a;
    layer0_outputs(7313) <= not (a and b);
    layer0_outputs(7314) <= not b;
    layer0_outputs(7315) <= not (a or b);
    layer0_outputs(7316) <= a xor b;
    layer0_outputs(7317) <= 1'b0;
    layer0_outputs(7318) <= a xor b;
    layer0_outputs(7319) <= a and not b;
    layer0_outputs(7320) <= a;
    layer0_outputs(7321) <= not b or a;
    layer0_outputs(7322) <= not a or b;
    layer0_outputs(7323) <= a or b;
    layer0_outputs(7324) <= a;
    layer0_outputs(7325) <= a xor b;
    layer0_outputs(7326) <= not a;
    layer0_outputs(7327) <= 1'b1;
    layer0_outputs(7328) <= not (a xor b);
    layer0_outputs(7329) <= not b or a;
    layer0_outputs(7330) <= b and not a;
    layer0_outputs(7331) <= a or b;
    layer0_outputs(7332) <= not b or a;
    layer0_outputs(7333) <= not a or b;
    layer0_outputs(7334) <= a xor b;
    layer0_outputs(7335) <= not b or a;
    layer0_outputs(7336) <= not a;
    layer0_outputs(7337) <= not (a or b);
    layer0_outputs(7338) <= a;
    layer0_outputs(7339) <= not (a xor b);
    layer0_outputs(7340) <= not (a xor b);
    layer0_outputs(7341) <= a or b;
    layer0_outputs(7342) <= b and not a;
    layer0_outputs(7343) <= not b or a;
    layer0_outputs(7344) <= a;
    layer0_outputs(7345) <= not (a or b);
    layer0_outputs(7346) <= 1'b0;
    layer0_outputs(7347) <= a and not b;
    layer0_outputs(7348) <= b and not a;
    layer0_outputs(7349) <= not b;
    layer0_outputs(7350) <= not (a or b);
    layer0_outputs(7351) <= a and b;
    layer0_outputs(7352) <= b;
    layer0_outputs(7353) <= b;
    layer0_outputs(7354) <= not a or b;
    layer0_outputs(7355) <= a xor b;
    layer0_outputs(7356) <= not b;
    layer0_outputs(7357) <= a xor b;
    layer0_outputs(7358) <= b;
    layer0_outputs(7359) <= not a or b;
    layer0_outputs(7360) <= not (a or b);
    layer0_outputs(7361) <= not a;
    layer0_outputs(7362) <= not b or a;
    layer0_outputs(7363) <= not a;
    layer0_outputs(7364) <= not (a xor b);
    layer0_outputs(7365) <= a xor b;
    layer0_outputs(7366) <= not b or a;
    layer0_outputs(7367) <= b and not a;
    layer0_outputs(7368) <= b;
    layer0_outputs(7369) <= b and not a;
    layer0_outputs(7370) <= a;
    layer0_outputs(7371) <= not a;
    layer0_outputs(7372) <= a and not b;
    layer0_outputs(7373) <= not a or b;
    layer0_outputs(7374) <= b and not a;
    layer0_outputs(7375) <= not (a or b);
    layer0_outputs(7376) <= not (a or b);
    layer0_outputs(7377) <= not a;
    layer0_outputs(7378) <= not a or b;
    layer0_outputs(7379) <= not b or a;
    layer0_outputs(7380) <= a and not b;
    layer0_outputs(7381) <= a;
    layer0_outputs(7382) <= not b or a;
    layer0_outputs(7383) <= a xor b;
    layer0_outputs(7384) <= a and not b;
    layer0_outputs(7385) <= a;
    layer0_outputs(7386) <= b;
    layer0_outputs(7387) <= not (a xor b);
    layer0_outputs(7388) <= a or b;
    layer0_outputs(7389) <= not a or b;
    layer0_outputs(7390) <= not a;
    layer0_outputs(7391) <= not (a xor b);
    layer0_outputs(7392) <= b;
    layer0_outputs(7393) <= a;
    layer0_outputs(7394) <= not b;
    layer0_outputs(7395) <= not (a or b);
    layer0_outputs(7396) <= b and not a;
    layer0_outputs(7397) <= b and not a;
    layer0_outputs(7398) <= a or b;
    layer0_outputs(7399) <= not a;
    layer0_outputs(7400) <= b;
    layer0_outputs(7401) <= not (a or b);
    layer0_outputs(7402) <= not a or b;
    layer0_outputs(7403) <= 1'b0;
    layer0_outputs(7404) <= not (a xor b);
    layer0_outputs(7405) <= not a;
    layer0_outputs(7406) <= b;
    layer0_outputs(7407) <= b and not a;
    layer0_outputs(7408) <= not (a or b);
    layer0_outputs(7409) <= not b or a;
    layer0_outputs(7410) <= a and b;
    layer0_outputs(7411) <= not (a xor b);
    layer0_outputs(7412) <= b;
    layer0_outputs(7413) <= not b or a;
    layer0_outputs(7414) <= not (a xor b);
    layer0_outputs(7415) <= a and not b;
    layer0_outputs(7416) <= a or b;
    layer0_outputs(7417) <= not b;
    layer0_outputs(7418) <= a and b;
    layer0_outputs(7419) <= a;
    layer0_outputs(7420) <= a;
    layer0_outputs(7421) <= b and not a;
    layer0_outputs(7422) <= not (a xor b);
    layer0_outputs(7423) <= a or b;
    layer0_outputs(7424) <= not (a xor b);
    layer0_outputs(7425) <= not a;
    layer0_outputs(7426) <= not (a xor b);
    layer0_outputs(7427) <= b and not a;
    layer0_outputs(7428) <= a xor b;
    layer0_outputs(7429) <= b and not a;
    layer0_outputs(7430) <= not (a xor b);
    layer0_outputs(7431) <= a xor b;
    layer0_outputs(7432) <= a or b;
    layer0_outputs(7433) <= not a or b;
    layer0_outputs(7434) <= not (a xor b);
    layer0_outputs(7435) <= a or b;
    layer0_outputs(7436) <= not a;
    layer0_outputs(7437) <= a xor b;
    layer0_outputs(7438) <= a and b;
    layer0_outputs(7439) <= not a;
    layer0_outputs(7440) <= not (a or b);
    layer0_outputs(7441) <= not a;
    layer0_outputs(7442) <= a;
    layer0_outputs(7443) <= not (a or b);
    layer0_outputs(7444) <= not b or a;
    layer0_outputs(7445) <= not b or a;
    layer0_outputs(7446) <= b;
    layer0_outputs(7447) <= a and not b;
    layer0_outputs(7448) <= not (a or b);
    layer0_outputs(7449) <= b;
    layer0_outputs(7450) <= not b;
    layer0_outputs(7451) <= not (a xor b);
    layer0_outputs(7452) <= not (a or b);
    layer0_outputs(7453) <= a and b;
    layer0_outputs(7454) <= a xor b;
    layer0_outputs(7455) <= 1'b1;
    layer0_outputs(7456) <= a or b;
    layer0_outputs(7457) <= a;
    layer0_outputs(7458) <= a and not b;
    layer0_outputs(7459) <= not a;
    layer0_outputs(7460) <= a and not b;
    layer0_outputs(7461) <= not a;
    layer0_outputs(7462) <= a and not b;
    layer0_outputs(7463) <= not (a or b);
    layer0_outputs(7464) <= not (a or b);
    layer0_outputs(7465) <= a or b;
    layer0_outputs(7466) <= not b;
    layer0_outputs(7467) <= a and not b;
    layer0_outputs(7468) <= a or b;
    layer0_outputs(7469) <= a or b;
    layer0_outputs(7470) <= a or b;
    layer0_outputs(7471) <= a and not b;
    layer0_outputs(7472) <= b and not a;
    layer0_outputs(7473) <= not b or a;
    layer0_outputs(7474) <= a or b;
    layer0_outputs(7475) <= a or b;
    layer0_outputs(7476) <= a or b;
    layer0_outputs(7477) <= not a or b;
    layer0_outputs(7478) <= a and not b;
    layer0_outputs(7479) <= a xor b;
    layer0_outputs(7480) <= a or b;
    layer0_outputs(7481) <= b and not a;
    layer0_outputs(7482) <= not (a or b);
    layer0_outputs(7483) <= a xor b;
    layer0_outputs(7484) <= a and b;
    layer0_outputs(7485) <= not a;
    layer0_outputs(7486) <= a and not b;
    layer0_outputs(7487) <= 1'b0;
    layer0_outputs(7488) <= not a or b;
    layer0_outputs(7489) <= b;
    layer0_outputs(7490) <= not b or a;
    layer0_outputs(7491) <= a xor b;
    layer0_outputs(7492) <= not a or b;
    layer0_outputs(7493) <= a xor b;
    layer0_outputs(7494) <= not b or a;
    layer0_outputs(7495) <= a xor b;
    layer0_outputs(7496) <= not (a and b);
    layer0_outputs(7497) <= not b or a;
    layer0_outputs(7498) <= not (a or b);
    layer0_outputs(7499) <= not a;
    layer0_outputs(7500) <= b;
    layer0_outputs(7501) <= not a or b;
    layer0_outputs(7502) <= a xor b;
    layer0_outputs(7503) <= a;
    layer0_outputs(7504) <= not a;
    layer0_outputs(7505) <= not (a xor b);
    layer0_outputs(7506) <= b and not a;
    layer0_outputs(7507) <= 1'b0;
    layer0_outputs(7508) <= not a;
    layer0_outputs(7509) <= not b;
    layer0_outputs(7510) <= not a;
    layer0_outputs(7511) <= b and not a;
    layer0_outputs(7512) <= not (a or b);
    layer0_outputs(7513) <= a xor b;
    layer0_outputs(7514) <= a xor b;
    layer0_outputs(7515) <= a or b;
    layer0_outputs(7516) <= a;
    layer0_outputs(7517) <= not (a or b);
    layer0_outputs(7518) <= not b;
    layer0_outputs(7519) <= not b;
    layer0_outputs(7520) <= not b;
    layer0_outputs(7521) <= a and not b;
    layer0_outputs(7522) <= a or b;
    layer0_outputs(7523) <= a and b;
    layer0_outputs(7524) <= a xor b;
    layer0_outputs(7525) <= b and not a;
    layer0_outputs(7526) <= 1'b1;
    layer0_outputs(7527) <= not a;
    layer0_outputs(7528) <= 1'b0;
    layer0_outputs(7529) <= not b;
    layer0_outputs(7530) <= 1'b0;
    layer0_outputs(7531) <= not a;
    layer0_outputs(7532) <= not a;
    layer0_outputs(7533) <= a or b;
    layer0_outputs(7534) <= not (a xor b);
    layer0_outputs(7535) <= not a;
    layer0_outputs(7536) <= not a;
    layer0_outputs(7537) <= a or b;
    layer0_outputs(7538) <= a xor b;
    layer0_outputs(7539) <= b;
    layer0_outputs(7540) <= b and not a;
    layer0_outputs(7541) <= a and b;
    layer0_outputs(7542) <= not b;
    layer0_outputs(7543) <= a or b;
    layer0_outputs(7544) <= not b;
    layer0_outputs(7545) <= not (a xor b);
    layer0_outputs(7546) <= not b;
    layer0_outputs(7547) <= a or b;
    layer0_outputs(7548) <= a or b;
    layer0_outputs(7549) <= not (a or b);
    layer0_outputs(7550) <= not a;
    layer0_outputs(7551) <= a or b;
    layer0_outputs(7552) <= a and not b;
    layer0_outputs(7553) <= not a or b;
    layer0_outputs(7554) <= b;
    layer0_outputs(7555) <= b and not a;
    layer0_outputs(7556) <= not b or a;
    layer0_outputs(7557) <= 1'b1;
    layer0_outputs(7558) <= 1'b0;
    layer0_outputs(7559) <= not a or b;
    layer0_outputs(7560) <= not (a or b);
    layer0_outputs(7561) <= not (a or b);
    layer0_outputs(7562) <= a xor b;
    layer0_outputs(7563) <= not b;
    layer0_outputs(7564) <= a xor b;
    layer0_outputs(7565) <= not a or b;
    layer0_outputs(7566) <= not b;
    layer0_outputs(7567) <= a;
    layer0_outputs(7568) <= a and not b;
    layer0_outputs(7569) <= not b or a;
    layer0_outputs(7570) <= not (a or b);
    layer0_outputs(7571) <= not b;
    layer0_outputs(7572) <= b and not a;
    layer0_outputs(7573) <= a and not b;
    layer0_outputs(7574) <= not (a or b);
    layer0_outputs(7575) <= not a;
    layer0_outputs(7576) <= a xor b;
    layer0_outputs(7577) <= b;
    layer0_outputs(7578) <= a xor b;
    layer0_outputs(7579) <= 1'b0;
    layer0_outputs(7580) <= b and not a;
    layer0_outputs(7581) <= not b;
    layer0_outputs(7582) <= a or b;
    layer0_outputs(7583) <= a;
    layer0_outputs(7584) <= not b or a;
    layer0_outputs(7585) <= a and not b;
    layer0_outputs(7586) <= 1'b1;
    layer0_outputs(7587) <= not (a xor b);
    layer0_outputs(7588) <= not b;
    layer0_outputs(7589) <= not a or b;
    layer0_outputs(7590) <= not a or b;
    layer0_outputs(7591) <= a xor b;
    layer0_outputs(7592) <= a;
    layer0_outputs(7593) <= b and not a;
    layer0_outputs(7594) <= a or b;
    layer0_outputs(7595) <= not a;
    layer0_outputs(7596) <= not (a or b);
    layer0_outputs(7597) <= not (a or b);
    layer0_outputs(7598) <= not (a or b);
    layer0_outputs(7599) <= b;
    layer0_outputs(7600) <= not (a or b);
    layer0_outputs(7601) <= not (a or b);
    layer0_outputs(7602) <= a and b;
    layer0_outputs(7603) <= a;
    layer0_outputs(7604) <= b;
    layer0_outputs(7605) <= not a or b;
    layer0_outputs(7606) <= not a;
    layer0_outputs(7607) <= a and not b;
    layer0_outputs(7608) <= b;
    layer0_outputs(7609) <= not b or a;
    layer0_outputs(7610) <= a or b;
    layer0_outputs(7611) <= not (a and b);
    layer0_outputs(7612) <= 1'b0;
    layer0_outputs(7613) <= a xor b;
    layer0_outputs(7614) <= not (a or b);
    layer0_outputs(7615) <= a and not b;
    layer0_outputs(7616) <= a or b;
    layer0_outputs(7617) <= not b or a;
    layer0_outputs(7618) <= not b;
    layer0_outputs(7619) <= not (a or b);
    layer0_outputs(7620) <= not a;
    layer0_outputs(7621) <= not (a or b);
    layer0_outputs(7622) <= a;
    layer0_outputs(7623) <= not (a or b);
    layer0_outputs(7624) <= b;
    layer0_outputs(7625) <= b and not a;
    layer0_outputs(7626) <= a or b;
    layer0_outputs(7627) <= not (a xor b);
    layer0_outputs(7628) <= not b or a;
    layer0_outputs(7629) <= b;
    layer0_outputs(7630) <= a and not b;
    layer0_outputs(7631) <= a or b;
    layer0_outputs(7632) <= not b;
    layer0_outputs(7633) <= a or b;
    layer0_outputs(7634) <= a or b;
    layer0_outputs(7635) <= not (a or b);
    layer0_outputs(7636) <= a or b;
    layer0_outputs(7637) <= not (a and b);
    layer0_outputs(7638) <= 1'b1;
    layer0_outputs(7639) <= a or b;
    layer0_outputs(7640) <= a;
    layer0_outputs(7641) <= a;
    layer0_outputs(7642) <= not a;
    layer0_outputs(7643) <= a or b;
    layer0_outputs(7644) <= b and not a;
    layer0_outputs(7645) <= b and not a;
    layer0_outputs(7646) <= a and not b;
    layer0_outputs(7647) <= a xor b;
    layer0_outputs(7648) <= a or b;
    layer0_outputs(7649) <= not (a or b);
    layer0_outputs(7650) <= not (a xor b);
    layer0_outputs(7651) <= a and not b;
    layer0_outputs(7652) <= b and not a;
    layer0_outputs(7653) <= not (a or b);
    layer0_outputs(7654) <= b;
    layer0_outputs(7655) <= b and not a;
    layer0_outputs(7656) <= not a;
    layer0_outputs(7657) <= a or b;
    layer0_outputs(7658) <= a xor b;
    layer0_outputs(7659) <= b and not a;
    layer0_outputs(7660) <= a xor b;
    layer0_outputs(7661) <= a or b;
    layer0_outputs(7662) <= a and not b;
    layer0_outputs(7663) <= b;
    layer0_outputs(7664) <= b and not a;
    layer0_outputs(7665) <= a and not b;
    layer0_outputs(7666) <= 1'b1;
    layer0_outputs(7667) <= a and not b;
    layer0_outputs(7668) <= not b;
    layer0_outputs(7669) <= not b or a;
    layer0_outputs(7670) <= a xor b;
    layer0_outputs(7671) <= a;
    layer0_outputs(7672) <= a;
    layer0_outputs(7673) <= b;
    layer0_outputs(7674) <= a;
    layer0_outputs(7675) <= a or b;
    layer0_outputs(7676) <= a and b;
    layer0_outputs(7677) <= b and not a;
    layer0_outputs(7678) <= a xor b;
    layer0_outputs(7679) <= not (a xor b);
    layer0_outputs(7680) <= b and not a;
    layer0_outputs(7681) <= b;
    layer0_outputs(7682) <= not a or b;
    layer0_outputs(7683) <= not (a and b);
    layer0_outputs(7684) <= not b or a;
    layer0_outputs(7685) <= not (a xor b);
    layer0_outputs(7686) <= 1'b0;
    layer0_outputs(7687) <= not b;
    layer0_outputs(7688) <= not b or a;
    layer0_outputs(7689) <= not (a or b);
    layer0_outputs(7690) <= not a or b;
    layer0_outputs(7691) <= a;
    layer0_outputs(7692) <= not (a or b);
    layer0_outputs(7693) <= not (a and b);
    layer0_outputs(7694) <= a and not b;
    layer0_outputs(7695) <= a and b;
    layer0_outputs(7696) <= not (a xor b);
    layer0_outputs(7697) <= a;
    layer0_outputs(7698) <= not b;
    layer0_outputs(7699) <= a or b;
    layer0_outputs(7700) <= not a;
    layer0_outputs(7701) <= not (a xor b);
    layer0_outputs(7702) <= a;
    layer0_outputs(7703) <= a or b;
    layer0_outputs(7704) <= not b;
    layer0_outputs(7705) <= a and not b;
    layer0_outputs(7706) <= b and not a;
    layer0_outputs(7707) <= b;
    layer0_outputs(7708) <= a xor b;
    layer0_outputs(7709) <= b;
    layer0_outputs(7710) <= a or b;
    layer0_outputs(7711) <= a xor b;
    layer0_outputs(7712) <= not (a or b);
    layer0_outputs(7713) <= a xor b;
    layer0_outputs(7714) <= a xor b;
    layer0_outputs(7715) <= not (a or b);
    layer0_outputs(7716) <= not (a or b);
    layer0_outputs(7717) <= not a;
    layer0_outputs(7718) <= not a;
    layer0_outputs(7719) <= not (a xor b);
    layer0_outputs(7720) <= a or b;
    layer0_outputs(7721) <= a or b;
    layer0_outputs(7722) <= a and not b;
    layer0_outputs(7723) <= a;
    layer0_outputs(7724) <= not (a xor b);
    layer0_outputs(7725) <= not b;
    layer0_outputs(7726) <= not b;
    layer0_outputs(7727) <= a xor b;
    layer0_outputs(7728) <= not a;
    layer0_outputs(7729) <= b and not a;
    layer0_outputs(7730) <= a or b;
    layer0_outputs(7731) <= a;
    layer0_outputs(7732) <= a and not b;
    layer0_outputs(7733) <= b;
    layer0_outputs(7734) <= not b;
    layer0_outputs(7735) <= not b;
    layer0_outputs(7736) <= not (a or b);
    layer0_outputs(7737) <= not b or a;
    layer0_outputs(7738) <= a or b;
    layer0_outputs(7739) <= not (a and b);
    layer0_outputs(7740) <= not (a xor b);
    layer0_outputs(7741) <= not (a or b);
    layer0_outputs(7742) <= not (a xor b);
    layer0_outputs(7743) <= b;
    layer0_outputs(7744) <= a or b;
    layer0_outputs(7745) <= not b;
    layer0_outputs(7746) <= a and not b;
    layer0_outputs(7747) <= a or b;
    layer0_outputs(7748) <= 1'b0;
    layer0_outputs(7749) <= 1'b0;
    layer0_outputs(7750) <= not b;
    layer0_outputs(7751) <= not (a or b);
    layer0_outputs(7752) <= not b;
    layer0_outputs(7753) <= a and not b;
    layer0_outputs(7754) <= a or b;
    layer0_outputs(7755) <= not (a or b);
    layer0_outputs(7756) <= not (a or b);
    layer0_outputs(7757) <= not (a xor b);
    layer0_outputs(7758) <= a or b;
    layer0_outputs(7759) <= a xor b;
    layer0_outputs(7760) <= not (a or b);
    layer0_outputs(7761) <= 1'b0;
    layer0_outputs(7762) <= a or b;
    layer0_outputs(7763) <= b;
    layer0_outputs(7764) <= not a;
    layer0_outputs(7765) <= not (a or b);
    layer0_outputs(7766) <= not a;
    layer0_outputs(7767) <= a xor b;
    layer0_outputs(7768) <= not (a or b);
    layer0_outputs(7769) <= a or b;
    layer0_outputs(7770) <= b;
    layer0_outputs(7771) <= b and not a;
    layer0_outputs(7772) <= a xor b;
    layer0_outputs(7773) <= not b or a;
    layer0_outputs(7774) <= a and not b;
    layer0_outputs(7775) <= not b;
    layer0_outputs(7776) <= a;
    layer0_outputs(7777) <= not (a or b);
    layer0_outputs(7778) <= a xor b;
    layer0_outputs(7779) <= 1'b0;
    layer0_outputs(7780) <= not (a xor b);
    layer0_outputs(7781) <= a xor b;
    layer0_outputs(7782) <= not b or a;
    layer0_outputs(7783) <= not b or a;
    layer0_outputs(7784) <= a or b;
    layer0_outputs(7785) <= b;
    layer0_outputs(7786) <= a or b;
    layer0_outputs(7787) <= a or b;
    layer0_outputs(7788) <= a xor b;
    layer0_outputs(7789) <= b and not a;
    layer0_outputs(7790) <= not (a xor b);
    layer0_outputs(7791) <= not (a xor b);
    layer0_outputs(7792) <= b and not a;
    layer0_outputs(7793) <= not b or a;
    layer0_outputs(7794) <= not b;
    layer0_outputs(7795) <= b;
    layer0_outputs(7796) <= a or b;
    layer0_outputs(7797) <= not a;
    layer0_outputs(7798) <= not a;
    layer0_outputs(7799) <= a and b;
    layer0_outputs(7800) <= not (a and b);
    layer0_outputs(7801) <= not a or b;
    layer0_outputs(7802) <= not (a xor b);
    layer0_outputs(7803) <= not (a xor b);
    layer0_outputs(7804) <= not a;
    layer0_outputs(7805) <= b;
    layer0_outputs(7806) <= a and not b;
    layer0_outputs(7807) <= a xor b;
    layer0_outputs(7808) <= not (a or b);
    layer0_outputs(7809) <= b;
    layer0_outputs(7810) <= a and not b;
    layer0_outputs(7811) <= not a or b;
    layer0_outputs(7812) <= not a or b;
    layer0_outputs(7813) <= not (a xor b);
    layer0_outputs(7814) <= a or b;
    layer0_outputs(7815) <= a and not b;
    layer0_outputs(7816) <= a or b;
    layer0_outputs(7817) <= a or b;
    layer0_outputs(7818) <= not b;
    layer0_outputs(7819) <= b and not a;
    layer0_outputs(7820) <= not (a xor b);
    layer0_outputs(7821) <= not b;
    layer0_outputs(7822) <= not (a xor b);
    layer0_outputs(7823) <= b;
    layer0_outputs(7824) <= not b or a;
    layer0_outputs(7825) <= 1'b1;
    layer0_outputs(7826) <= not (a xor b);
    layer0_outputs(7827) <= not b;
    layer0_outputs(7828) <= not b or a;
    layer0_outputs(7829) <= 1'b0;
    layer0_outputs(7830) <= not b or a;
    layer0_outputs(7831) <= a xor b;
    layer0_outputs(7832) <= b and not a;
    layer0_outputs(7833) <= not a;
    layer0_outputs(7834) <= a or b;
    layer0_outputs(7835) <= 1'b1;
    layer0_outputs(7836) <= not b;
    layer0_outputs(7837) <= not b;
    layer0_outputs(7838) <= not (a or b);
    layer0_outputs(7839) <= not a or b;
    layer0_outputs(7840) <= 1'b1;
    layer0_outputs(7841) <= a;
    layer0_outputs(7842) <= a or b;
    layer0_outputs(7843) <= not (a or b);
    layer0_outputs(7844) <= a and not b;
    layer0_outputs(7845) <= not (a xor b);
    layer0_outputs(7846) <= a or b;
    layer0_outputs(7847) <= not b;
    layer0_outputs(7848) <= not b or a;
    layer0_outputs(7849) <= not (a or b);
    layer0_outputs(7850) <= not (a or b);
    layer0_outputs(7851) <= not a or b;
    layer0_outputs(7852) <= not (a xor b);
    layer0_outputs(7853) <= 1'b0;
    layer0_outputs(7854) <= a;
    layer0_outputs(7855) <= not a or b;
    layer0_outputs(7856) <= b and not a;
    layer0_outputs(7857) <= 1'b0;
    layer0_outputs(7858) <= not a or b;
    layer0_outputs(7859) <= not a;
    layer0_outputs(7860) <= not (a and b);
    layer0_outputs(7861) <= not (a or b);
    layer0_outputs(7862) <= not a or b;
    layer0_outputs(7863) <= not a;
    layer0_outputs(7864) <= not b or a;
    layer0_outputs(7865) <= a or b;
    layer0_outputs(7866) <= b and not a;
    layer0_outputs(7867) <= not (a or b);
    layer0_outputs(7868) <= a or b;
    layer0_outputs(7869) <= b and not a;
    layer0_outputs(7870) <= 1'b0;
    layer0_outputs(7871) <= not b;
    layer0_outputs(7872) <= not b;
    layer0_outputs(7873) <= a;
    layer0_outputs(7874) <= a xor b;
    layer0_outputs(7875) <= a xor b;
    layer0_outputs(7876) <= a xor b;
    layer0_outputs(7877) <= a xor b;
    layer0_outputs(7878) <= not (a xor b);
    layer0_outputs(7879) <= a xor b;
    layer0_outputs(7880) <= a and not b;
    layer0_outputs(7881) <= a;
    layer0_outputs(7882) <= 1'b1;
    layer0_outputs(7883) <= b;
    layer0_outputs(7884) <= a;
    layer0_outputs(7885) <= a and not b;
    layer0_outputs(7886) <= b;
    layer0_outputs(7887) <= a or b;
    layer0_outputs(7888) <= not a;
    layer0_outputs(7889) <= not (a or b);
    layer0_outputs(7890) <= a xor b;
    layer0_outputs(7891) <= a or b;
    layer0_outputs(7892) <= not a;
    layer0_outputs(7893) <= not (a xor b);
    layer0_outputs(7894) <= not (a or b);
    layer0_outputs(7895) <= a and not b;
    layer0_outputs(7896) <= a or b;
    layer0_outputs(7897) <= not (a or b);
    layer0_outputs(7898) <= not (a or b);
    layer0_outputs(7899) <= not b or a;
    layer0_outputs(7900) <= not (a xor b);
    layer0_outputs(7901) <= a;
    layer0_outputs(7902) <= a or b;
    layer0_outputs(7903) <= not (a or b);
    layer0_outputs(7904) <= a or b;
    layer0_outputs(7905) <= not (a or b);
    layer0_outputs(7906) <= b and not a;
    layer0_outputs(7907) <= a or b;
    layer0_outputs(7908) <= b;
    layer0_outputs(7909) <= not (a and b);
    layer0_outputs(7910) <= a xor b;
    layer0_outputs(7911) <= not a or b;
    layer0_outputs(7912) <= a xor b;
    layer0_outputs(7913) <= a or b;
    layer0_outputs(7914) <= a or b;
    layer0_outputs(7915) <= a;
    layer0_outputs(7916) <= not (a xor b);
    layer0_outputs(7917) <= a and not b;
    layer0_outputs(7918) <= not b;
    layer0_outputs(7919) <= not a or b;
    layer0_outputs(7920) <= a or b;
    layer0_outputs(7921) <= a xor b;
    layer0_outputs(7922) <= not b or a;
    layer0_outputs(7923) <= not b or a;
    layer0_outputs(7924) <= a and not b;
    layer0_outputs(7925) <= a or b;
    layer0_outputs(7926) <= a or b;
    layer0_outputs(7927) <= a;
    layer0_outputs(7928) <= a xor b;
    layer0_outputs(7929) <= a or b;
    layer0_outputs(7930) <= not (a or b);
    layer0_outputs(7931) <= not (a or b);
    layer0_outputs(7932) <= not (a or b);
    layer0_outputs(7933) <= a xor b;
    layer0_outputs(7934) <= not a or b;
    layer0_outputs(7935) <= a xor b;
    layer0_outputs(7936) <= b and not a;
    layer0_outputs(7937) <= a and not b;
    layer0_outputs(7938) <= a xor b;
    layer0_outputs(7939) <= not (a xor b);
    layer0_outputs(7940) <= b;
    layer0_outputs(7941) <= not (a or b);
    layer0_outputs(7942) <= b;
    layer0_outputs(7943) <= not (a or b);
    layer0_outputs(7944) <= a and not b;
    layer0_outputs(7945) <= not (a or b);
    layer0_outputs(7946) <= not b;
    layer0_outputs(7947) <= not (a xor b);
    layer0_outputs(7948) <= not (a or b);
    layer0_outputs(7949) <= a xor b;
    layer0_outputs(7950) <= a or b;
    layer0_outputs(7951) <= b and not a;
    layer0_outputs(7952) <= not (a or b);
    layer0_outputs(7953) <= not (a or b);
    layer0_outputs(7954) <= b;
    layer0_outputs(7955) <= a xor b;
    layer0_outputs(7956) <= a xor b;
    layer0_outputs(7957) <= not (a xor b);
    layer0_outputs(7958) <= not (a xor b);
    layer0_outputs(7959) <= not a;
    layer0_outputs(7960) <= not b;
    layer0_outputs(7961) <= not a;
    layer0_outputs(7962) <= not (a xor b);
    layer0_outputs(7963) <= 1'b0;
    layer0_outputs(7964) <= a or b;
    layer0_outputs(7965) <= b and not a;
    layer0_outputs(7966) <= b and not a;
    layer0_outputs(7967) <= 1'b0;
    layer0_outputs(7968) <= a and not b;
    layer0_outputs(7969) <= not (a xor b);
    layer0_outputs(7970) <= b and not a;
    layer0_outputs(7971) <= a or b;
    layer0_outputs(7972) <= not b or a;
    layer0_outputs(7973) <= a;
    layer0_outputs(7974) <= 1'b1;
    layer0_outputs(7975) <= a xor b;
    layer0_outputs(7976) <= not (a or b);
    layer0_outputs(7977) <= 1'b1;
    layer0_outputs(7978) <= b;
    layer0_outputs(7979) <= a;
    layer0_outputs(7980) <= b;
    layer0_outputs(7981) <= not (a xor b);
    layer0_outputs(7982) <= not (a or b);
    layer0_outputs(7983) <= not a or b;
    layer0_outputs(7984) <= not (a or b);
    layer0_outputs(7985) <= a or b;
    layer0_outputs(7986) <= a xor b;
    layer0_outputs(7987) <= a or b;
    layer0_outputs(7988) <= not (a or b);
    layer0_outputs(7989) <= not (a xor b);
    layer0_outputs(7990) <= b and not a;
    layer0_outputs(7991) <= not b;
    layer0_outputs(7992) <= a or b;
    layer0_outputs(7993) <= not (a xor b);
    layer0_outputs(7994) <= a xor b;
    layer0_outputs(7995) <= not b;
    layer0_outputs(7996) <= a and not b;
    layer0_outputs(7997) <= a or b;
    layer0_outputs(7998) <= a and not b;
    layer0_outputs(7999) <= a xor b;
    layer0_outputs(8000) <= not a or b;
    layer0_outputs(8001) <= not (a and b);
    layer0_outputs(8002) <= not a or b;
    layer0_outputs(8003) <= b and not a;
    layer0_outputs(8004) <= not (a xor b);
    layer0_outputs(8005) <= a;
    layer0_outputs(8006) <= not (a or b);
    layer0_outputs(8007) <= a and not b;
    layer0_outputs(8008) <= not a;
    layer0_outputs(8009) <= not (a xor b);
    layer0_outputs(8010) <= a;
    layer0_outputs(8011) <= not a or b;
    layer0_outputs(8012) <= a or b;
    layer0_outputs(8013) <= 1'b1;
    layer0_outputs(8014) <= not b or a;
    layer0_outputs(8015) <= not (a or b);
    layer0_outputs(8016) <= not (a or b);
    layer0_outputs(8017) <= not (a xor b);
    layer0_outputs(8018) <= b;
    layer0_outputs(8019) <= not b or a;
    layer0_outputs(8020) <= a;
    layer0_outputs(8021) <= not (a xor b);
    layer0_outputs(8022) <= not b;
    layer0_outputs(8023) <= a and not b;
    layer0_outputs(8024) <= b;
    layer0_outputs(8025) <= a and b;
    layer0_outputs(8026) <= b and not a;
    layer0_outputs(8027) <= b and not a;
    layer0_outputs(8028) <= a or b;
    layer0_outputs(8029) <= b and not a;
    layer0_outputs(8030) <= not (a or b);
    layer0_outputs(8031) <= a xor b;
    layer0_outputs(8032) <= 1'b0;
    layer0_outputs(8033) <= a;
    layer0_outputs(8034) <= not (a xor b);
    layer0_outputs(8035) <= not b or a;
    layer0_outputs(8036) <= b and not a;
    layer0_outputs(8037) <= a and not b;
    layer0_outputs(8038) <= a;
    layer0_outputs(8039) <= a and b;
    layer0_outputs(8040) <= 1'b0;
    layer0_outputs(8041) <= b;
    layer0_outputs(8042) <= not (a or b);
    layer0_outputs(8043) <= not (a or b);
    layer0_outputs(8044) <= not a or b;
    layer0_outputs(8045) <= a xor b;
    layer0_outputs(8046) <= a or b;
    layer0_outputs(8047) <= not b;
    layer0_outputs(8048) <= not b or a;
    layer0_outputs(8049) <= b and not a;
    layer0_outputs(8050) <= a and not b;
    layer0_outputs(8051) <= b and not a;
    layer0_outputs(8052) <= not a;
    layer0_outputs(8053) <= a and b;
    layer0_outputs(8054) <= not a;
    layer0_outputs(8055) <= not (a or b);
    layer0_outputs(8056) <= a and not b;
    layer0_outputs(8057) <= b and not a;
    layer0_outputs(8058) <= not (a or b);
    layer0_outputs(8059) <= a and not b;
    layer0_outputs(8060) <= not (a or b);
    layer0_outputs(8061) <= a or b;
    layer0_outputs(8062) <= not a;
    layer0_outputs(8063) <= a or b;
    layer0_outputs(8064) <= not (a or b);
    layer0_outputs(8065) <= a xor b;
    layer0_outputs(8066) <= a xor b;
    layer0_outputs(8067) <= not (a xor b);
    layer0_outputs(8068) <= not (a or b);
    layer0_outputs(8069) <= a and not b;
    layer0_outputs(8070) <= not a;
    layer0_outputs(8071) <= a or b;
    layer0_outputs(8072) <= not (a or b);
    layer0_outputs(8073) <= not a or b;
    layer0_outputs(8074) <= not (a and b);
    layer0_outputs(8075) <= not b or a;
    layer0_outputs(8076) <= b and not a;
    layer0_outputs(8077) <= not b;
    layer0_outputs(8078) <= not b;
    layer0_outputs(8079) <= not (a or b);
    layer0_outputs(8080) <= a and not b;
    layer0_outputs(8081) <= a;
    layer0_outputs(8082) <= a xor b;
    layer0_outputs(8083) <= 1'b1;
    layer0_outputs(8084) <= a or b;
    layer0_outputs(8085) <= a;
    layer0_outputs(8086) <= not b or a;
    layer0_outputs(8087) <= not (a xor b);
    layer0_outputs(8088) <= a xor b;
    layer0_outputs(8089) <= a;
    layer0_outputs(8090) <= 1'b0;
    layer0_outputs(8091) <= b and not a;
    layer0_outputs(8092) <= not (a or b);
    layer0_outputs(8093) <= a xor b;
    layer0_outputs(8094) <= a xor b;
    layer0_outputs(8095) <= a and not b;
    layer0_outputs(8096) <= not (a xor b);
    layer0_outputs(8097) <= not (a or b);
    layer0_outputs(8098) <= not b;
    layer0_outputs(8099) <= not b;
    layer0_outputs(8100) <= not a or b;
    layer0_outputs(8101) <= a or b;
    layer0_outputs(8102) <= a xor b;
    layer0_outputs(8103) <= b and not a;
    layer0_outputs(8104) <= not (a or b);
    layer0_outputs(8105) <= b;
    layer0_outputs(8106) <= a or b;
    layer0_outputs(8107) <= not (a xor b);
    layer0_outputs(8108) <= a xor b;
    layer0_outputs(8109) <= not a;
    layer0_outputs(8110) <= a xor b;
    layer0_outputs(8111) <= 1'b0;
    layer0_outputs(8112) <= not (a or b);
    layer0_outputs(8113) <= not (a or b);
    layer0_outputs(8114) <= not (a and b);
    layer0_outputs(8115) <= a;
    layer0_outputs(8116) <= b;
    layer0_outputs(8117) <= not (a xor b);
    layer0_outputs(8118) <= not b or a;
    layer0_outputs(8119) <= a and b;
    layer0_outputs(8120) <= a;
    layer0_outputs(8121) <= not b or a;
    layer0_outputs(8122) <= not b or a;
    layer0_outputs(8123) <= not b;
    layer0_outputs(8124) <= a xor b;
    layer0_outputs(8125) <= a or b;
    layer0_outputs(8126) <= not b or a;
    layer0_outputs(8127) <= not (a or b);
    layer0_outputs(8128) <= not (a xor b);
    layer0_outputs(8129) <= a xor b;
    layer0_outputs(8130) <= not (a xor b);
    layer0_outputs(8131) <= b and not a;
    layer0_outputs(8132) <= not (a and b);
    layer0_outputs(8133) <= not (a xor b);
    layer0_outputs(8134) <= a or b;
    layer0_outputs(8135) <= not b or a;
    layer0_outputs(8136) <= not (a xor b);
    layer0_outputs(8137) <= not (a xor b);
    layer0_outputs(8138) <= a or b;
    layer0_outputs(8139) <= 1'b0;
    layer0_outputs(8140) <= b;
    layer0_outputs(8141) <= a;
    layer0_outputs(8142) <= a xor b;
    layer0_outputs(8143) <= not b or a;
    layer0_outputs(8144) <= a;
    layer0_outputs(8145) <= not a or b;
    layer0_outputs(8146) <= not b;
    layer0_outputs(8147) <= b;
    layer0_outputs(8148) <= not (a and b);
    layer0_outputs(8149) <= not a;
    layer0_outputs(8150) <= a or b;
    layer0_outputs(8151) <= not (a or b);
    layer0_outputs(8152) <= a or b;
    layer0_outputs(8153) <= not (a or b);
    layer0_outputs(8154) <= not b or a;
    layer0_outputs(8155) <= a xor b;
    layer0_outputs(8156) <= a xor b;
    layer0_outputs(8157) <= a and b;
    layer0_outputs(8158) <= not (a xor b);
    layer0_outputs(8159) <= a;
    layer0_outputs(8160) <= not (a xor b);
    layer0_outputs(8161) <= not (a xor b);
    layer0_outputs(8162) <= not (a or b);
    layer0_outputs(8163) <= a xor b;
    layer0_outputs(8164) <= a or b;
    layer0_outputs(8165) <= not (a or b);
    layer0_outputs(8166) <= a or b;
    layer0_outputs(8167) <= not a or b;
    layer0_outputs(8168) <= a or b;
    layer0_outputs(8169) <= not (a and b);
    layer0_outputs(8170) <= b;
    layer0_outputs(8171) <= a and not b;
    layer0_outputs(8172) <= a or b;
    layer0_outputs(8173) <= b and not a;
    layer0_outputs(8174) <= not a or b;
    layer0_outputs(8175) <= not b or a;
    layer0_outputs(8176) <= not a;
    layer0_outputs(8177) <= not a;
    layer0_outputs(8178) <= 1'b0;
    layer0_outputs(8179) <= a xor b;
    layer0_outputs(8180) <= not a;
    layer0_outputs(8181) <= b and not a;
    layer0_outputs(8182) <= 1'b0;
    layer0_outputs(8183) <= a and not b;
    layer0_outputs(8184) <= not b;
    layer0_outputs(8185) <= a xor b;
    layer0_outputs(8186) <= not (a or b);
    layer0_outputs(8187) <= not b or a;
    layer0_outputs(8188) <= not a or b;
    layer0_outputs(8189) <= not b;
    layer0_outputs(8190) <= a and not b;
    layer0_outputs(8191) <= a or b;
    layer0_outputs(8192) <= a xor b;
    layer0_outputs(8193) <= a or b;
    layer0_outputs(8194) <= not (a or b);
    layer0_outputs(8195) <= a xor b;
    layer0_outputs(8196) <= a or b;
    layer0_outputs(8197) <= not (a or b);
    layer0_outputs(8198) <= a xor b;
    layer0_outputs(8199) <= a and not b;
    layer0_outputs(8200) <= not (a or b);
    layer0_outputs(8201) <= b and not a;
    layer0_outputs(8202) <= 1'b0;
    layer0_outputs(8203) <= a and not b;
    layer0_outputs(8204) <= a or b;
    layer0_outputs(8205) <= a and not b;
    layer0_outputs(8206) <= not (a and b);
    layer0_outputs(8207) <= not b or a;
    layer0_outputs(8208) <= b and not a;
    layer0_outputs(8209) <= a or b;
    layer0_outputs(8210) <= a and not b;
    layer0_outputs(8211) <= a or b;
    layer0_outputs(8212) <= not (a or b);
    layer0_outputs(8213) <= not a;
    layer0_outputs(8214) <= not b;
    layer0_outputs(8215) <= not a or b;
    layer0_outputs(8216) <= not (a xor b);
    layer0_outputs(8217) <= not a;
    layer0_outputs(8218) <= b and not a;
    layer0_outputs(8219) <= not (a or b);
    layer0_outputs(8220) <= b;
    layer0_outputs(8221) <= 1'b0;
    layer0_outputs(8222) <= not (a xor b);
    layer0_outputs(8223) <= a or b;
    layer0_outputs(8224) <= not b or a;
    layer0_outputs(8225) <= not a;
    layer0_outputs(8226) <= a xor b;
    layer0_outputs(8227) <= not (a xor b);
    layer0_outputs(8228) <= a xor b;
    layer0_outputs(8229) <= not a;
    layer0_outputs(8230) <= a;
    layer0_outputs(8231) <= not b;
    layer0_outputs(8232) <= a xor b;
    layer0_outputs(8233) <= not (a or b);
    layer0_outputs(8234) <= not (a or b);
    layer0_outputs(8235) <= not (a or b);
    layer0_outputs(8236) <= a;
    layer0_outputs(8237) <= not b;
    layer0_outputs(8238) <= a or b;
    layer0_outputs(8239) <= not a or b;
    layer0_outputs(8240) <= b and not a;
    layer0_outputs(8241) <= not (a xor b);
    layer0_outputs(8242) <= 1'b1;
    layer0_outputs(8243) <= not a;
    layer0_outputs(8244) <= not (a xor b);
    layer0_outputs(8245) <= not (a xor b);
    layer0_outputs(8246) <= a or b;
    layer0_outputs(8247) <= a and b;
    layer0_outputs(8248) <= a;
    layer0_outputs(8249) <= b and not a;
    layer0_outputs(8250) <= b;
    layer0_outputs(8251) <= a and not b;
    layer0_outputs(8252) <= 1'b1;
    layer0_outputs(8253) <= not b or a;
    layer0_outputs(8254) <= a xor b;
    layer0_outputs(8255) <= not (a or b);
    layer0_outputs(8256) <= not (a xor b);
    layer0_outputs(8257) <= a and not b;
    layer0_outputs(8258) <= a and b;
    layer0_outputs(8259) <= a xor b;
    layer0_outputs(8260) <= a and not b;
    layer0_outputs(8261) <= not a;
    layer0_outputs(8262) <= a;
    layer0_outputs(8263) <= not b;
    layer0_outputs(8264) <= b and not a;
    layer0_outputs(8265) <= a xor b;
    layer0_outputs(8266) <= a;
    layer0_outputs(8267) <= not (a and b);
    layer0_outputs(8268) <= a and b;
    layer0_outputs(8269) <= not (a or b);
    layer0_outputs(8270) <= a;
    layer0_outputs(8271) <= not a or b;
    layer0_outputs(8272) <= not b;
    layer0_outputs(8273) <= a xor b;
    layer0_outputs(8274) <= a or b;
    layer0_outputs(8275) <= not (a or b);
    layer0_outputs(8276) <= a xor b;
    layer0_outputs(8277) <= a or b;
    layer0_outputs(8278) <= 1'b0;
    layer0_outputs(8279) <= a or b;
    layer0_outputs(8280) <= a xor b;
    layer0_outputs(8281) <= not (a xor b);
    layer0_outputs(8282) <= a and not b;
    layer0_outputs(8283) <= not b or a;
    layer0_outputs(8284) <= a or b;
    layer0_outputs(8285) <= b;
    layer0_outputs(8286) <= a;
    layer0_outputs(8287) <= not (a or b);
    layer0_outputs(8288) <= b;
    layer0_outputs(8289) <= not (a or b);
    layer0_outputs(8290) <= a and not b;
    layer0_outputs(8291) <= a and not b;
    layer0_outputs(8292) <= a and not b;
    layer0_outputs(8293) <= not (a xor b);
    layer0_outputs(8294) <= a;
    layer0_outputs(8295) <= a xor b;
    layer0_outputs(8296) <= not (a xor b);
    layer0_outputs(8297) <= a or b;
    layer0_outputs(8298) <= a xor b;
    layer0_outputs(8299) <= not b;
    layer0_outputs(8300) <= not (a or b);
    layer0_outputs(8301) <= not b or a;
    layer0_outputs(8302) <= a xor b;
    layer0_outputs(8303) <= not b;
    layer0_outputs(8304) <= not b or a;
    layer0_outputs(8305) <= a;
    layer0_outputs(8306) <= a xor b;
    layer0_outputs(8307) <= not (a or b);
    layer0_outputs(8308) <= a xor b;
    layer0_outputs(8309) <= not (a or b);
    layer0_outputs(8310) <= a xor b;
    layer0_outputs(8311) <= not b or a;
    layer0_outputs(8312) <= not (a xor b);
    layer0_outputs(8313) <= not b;
    layer0_outputs(8314) <= a or b;
    layer0_outputs(8315) <= 1'b0;
    layer0_outputs(8316) <= a and b;
    layer0_outputs(8317) <= b;
    layer0_outputs(8318) <= a or b;
    layer0_outputs(8319) <= not (a and b);
    layer0_outputs(8320) <= not (a xor b);
    layer0_outputs(8321) <= b;
    layer0_outputs(8322) <= b;
    layer0_outputs(8323) <= not (a or b);
    layer0_outputs(8324) <= a or b;
    layer0_outputs(8325) <= a;
    layer0_outputs(8326) <= a or b;
    layer0_outputs(8327) <= a and not b;
    layer0_outputs(8328) <= not (a or b);
    layer0_outputs(8329) <= a and not b;
    layer0_outputs(8330) <= not b;
    layer0_outputs(8331) <= 1'b0;
    layer0_outputs(8332) <= not b;
    layer0_outputs(8333) <= not (a or b);
    layer0_outputs(8334) <= b and not a;
    layer0_outputs(8335) <= a or b;
    layer0_outputs(8336) <= a xor b;
    layer0_outputs(8337) <= a and not b;
    layer0_outputs(8338) <= a or b;
    layer0_outputs(8339) <= not (a xor b);
    layer0_outputs(8340) <= b and not a;
    layer0_outputs(8341) <= not b;
    layer0_outputs(8342) <= not a or b;
    layer0_outputs(8343) <= a or b;
    layer0_outputs(8344) <= not a;
    layer0_outputs(8345) <= a;
    layer0_outputs(8346) <= a and not b;
    layer0_outputs(8347) <= not b or a;
    layer0_outputs(8348) <= a or b;
    layer0_outputs(8349) <= not (a or b);
    layer0_outputs(8350) <= not (a or b);
    layer0_outputs(8351) <= a or b;
    layer0_outputs(8352) <= a or b;
    layer0_outputs(8353) <= not (a or b);
    layer0_outputs(8354) <= not (a or b);
    layer0_outputs(8355) <= not b or a;
    layer0_outputs(8356) <= not (a or b);
    layer0_outputs(8357) <= a and b;
    layer0_outputs(8358) <= a xor b;
    layer0_outputs(8359) <= b and not a;
    layer0_outputs(8360) <= a or b;
    layer0_outputs(8361) <= not b or a;
    layer0_outputs(8362) <= a and not b;
    layer0_outputs(8363) <= not (a or b);
    layer0_outputs(8364) <= 1'b0;
    layer0_outputs(8365) <= b and not a;
    layer0_outputs(8366) <= not (a xor b);
    layer0_outputs(8367) <= not b;
    layer0_outputs(8368) <= not b;
    layer0_outputs(8369) <= a or b;
    layer0_outputs(8370) <= 1'b1;
    layer0_outputs(8371) <= not (a or b);
    layer0_outputs(8372) <= not b;
    layer0_outputs(8373) <= not a or b;
    layer0_outputs(8374) <= not (a and b);
    layer0_outputs(8375) <= not (a xor b);
    layer0_outputs(8376) <= not b;
    layer0_outputs(8377) <= not a or b;
    layer0_outputs(8378) <= a or b;
    layer0_outputs(8379) <= not (a xor b);
    layer0_outputs(8380) <= a and not b;
    layer0_outputs(8381) <= a;
    layer0_outputs(8382) <= a or b;
    layer0_outputs(8383) <= not (a or b);
    layer0_outputs(8384) <= not (a and b);
    layer0_outputs(8385) <= not a or b;
    layer0_outputs(8386) <= not a or b;
    layer0_outputs(8387) <= not b;
    layer0_outputs(8388) <= not b or a;
    layer0_outputs(8389) <= not a;
    layer0_outputs(8390) <= a or b;
    layer0_outputs(8391) <= not (a xor b);
    layer0_outputs(8392) <= a or b;
    layer0_outputs(8393) <= a and not b;
    layer0_outputs(8394) <= a or b;
    layer0_outputs(8395) <= not b;
    layer0_outputs(8396) <= not a or b;
    layer0_outputs(8397) <= b and not a;
    layer0_outputs(8398) <= not a;
    layer0_outputs(8399) <= b and not a;
    layer0_outputs(8400) <= not b or a;
    layer0_outputs(8401) <= not (a or b);
    layer0_outputs(8402) <= not b or a;
    layer0_outputs(8403) <= b and not a;
    layer0_outputs(8404) <= not (a xor b);
    layer0_outputs(8405) <= a or b;
    layer0_outputs(8406) <= not (a or b);
    layer0_outputs(8407) <= not (a and b);
    layer0_outputs(8408) <= not a;
    layer0_outputs(8409) <= not b or a;
    layer0_outputs(8410) <= not (a xor b);
    layer0_outputs(8411) <= not (a xor b);
    layer0_outputs(8412) <= b;
    layer0_outputs(8413) <= a;
    layer0_outputs(8414) <= b and not a;
    layer0_outputs(8415) <= not (a or b);
    layer0_outputs(8416) <= a or b;
    layer0_outputs(8417) <= a;
    layer0_outputs(8418) <= not b;
    layer0_outputs(8419) <= b and not a;
    layer0_outputs(8420) <= a xor b;
    layer0_outputs(8421) <= b and not a;
    layer0_outputs(8422) <= a xor b;
    layer0_outputs(8423) <= not (a or b);
    layer0_outputs(8424) <= not a or b;
    layer0_outputs(8425) <= a and not b;
    layer0_outputs(8426) <= not a;
    layer0_outputs(8427) <= not (a xor b);
    layer0_outputs(8428) <= 1'b1;
    layer0_outputs(8429) <= a and not b;
    layer0_outputs(8430) <= not b;
    layer0_outputs(8431) <= a xor b;
    layer0_outputs(8432) <= not b or a;
    layer0_outputs(8433) <= a;
    layer0_outputs(8434) <= not (a xor b);
    layer0_outputs(8435) <= a or b;
    layer0_outputs(8436) <= not b;
    layer0_outputs(8437) <= a;
    layer0_outputs(8438) <= not a or b;
    layer0_outputs(8439) <= a or b;
    layer0_outputs(8440) <= b and not a;
    layer0_outputs(8441) <= a and not b;
    layer0_outputs(8442) <= not b or a;
    layer0_outputs(8443) <= not (a or b);
    layer0_outputs(8444) <= a xor b;
    layer0_outputs(8445) <= a xor b;
    layer0_outputs(8446) <= 1'b1;
    layer0_outputs(8447) <= not a;
    layer0_outputs(8448) <= not a;
    layer0_outputs(8449) <= a or b;
    layer0_outputs(8450) <= not a or b;
    layer0_outputs(8451) <= not (a xor b);
    layer0_outputs(8452) <= not (a xor b);
    layer0_outputs(8453) <= a and not b;
    layer0_outputs(8454) <= a xor b;
    layer0_outputs(8455) <= not (a xor b);
    layer0_outputs(8456) <= not (a and b);
    layer0_outputs(8457) <= not (a or b);
    layer0_outputs(8458) <= not a;
    layer0_outputs(8459) <= a and not b;
    layer0_outputs(8460) <= a and not b;
    layer0_outputs(8461) <= 1'b0;
    layer0_outputs(8462) <= not a;
    layer0_outputs(8463) <= not (a xor b);
    layer0_outputs(8464) <= a or b;
    layer0_outputs(8465) <= b;
    layer0_outputs(8466) <= not b;
    layer0_outputs(8467) <= a and not b;
    layer0_outputs(8468) <= not (a xor b);
    layer0_outputs(8469) <= not (a or b);
    layer0_outputs(8470) <= 1'b1;
    layer0_outputs(8471) <= not a;
    layer0_outputs(8472) <= not (a or b);
    layer0_outputs(8473) <= not (a xor b);
    layer0_outputs(8474) <= a;
    layer0_outputs(8475) <= not (a xor b);
    layer0_outputs(8476) <= a and b;
    layer0_outputs(8477) <= a xor b;
    layer0_outputs(8478) <= not (a or b);
    layer0_outputs(8479) <= a or b;
    layer0_outputs(8480) <= a or b;
    layer0_outputs(8481) <= a and not b;
    layer0_outputs(8482) <= not (a or b);
    layer0_outputs(8483) <= not (a and b);
    layer0_outputs(8484) <= not a or b;
    layer0_outputs(8485) <= a;
    layer0_outputs(8486) <= not b or a;
    layer0_outputs(8487) <= a and not b;
    layer0_outputs(8488) <= a and b;
    layer0_outputs(8489) <= a and not b;
    layer0_outputs(8490) <= not (a or b);
    layer0_outputs(8491) <= a or b;
    layer0_outputs(8492) <= not (a or b);
    layer0_outputs(8493) <= a or b;
    layer0_outputs(8494) <= a and not b;
    layer0_outputs(8495) <= a xor b;
    layer0_outputs(8496) <= a xor b;
    layer0_outputs(8497) <= not b or a;
    layer0_outputs(8498) <= a;
    layer0_outputs(8499) <= not (a or b);
    layer0_outputs(8500) <= not (a or b);
    layer0_outputs(8501) <= not (a xor b);
    layer0_outputs(8502) <= b;
    layer0_outputs(8503) <= a xor b;
    layer0_outputs(8504) <= b;
    layer0_outputs(8505) <= a and not b;
    layer0_outputs(8506) <= not (a or b);
    layer0_outputs(8507) <= a or b;
    layer0_outputs(8508) <= not (a or b);
    layer0_outputs(8509) <= a or b;
    layer0_outputs(8510) <= not a or b;
    layer0_outputs(8511) <= not (a or b);
    layer0_outputs(8512) <= not (a or b);
    layer0_outputs(8513) <= a;
    layer0_outputs(8514) <= a and not b;
    layer0_outputs(8515) <= 1'b1;
    layer0_outputs(8516) <= a or b;
    layer0_outputs(8517) <= a or b;
    layer0_outputs(8518) <= a and not b;
    layer0_outputs(8519) <= a xor b;
    layer0_outputs(8520) <= a xor b;
    layer0_outputs(8521) <= a or b;
    layer0_outputs(8522) <= b and not a;
    layer0_outputs(8523) <= not (a or b);
    layer0_outputs(8524) <= a and b;
    layer0_outputs(8525) <= not (a or b);
    layer0_outputs(8526) <= not b;
    layer0_outputs(8527) <= a or b;
    layer0_outputs(8528) <= not b or a;
    layer0_outputs(8529) <= not b;
    layer0_outputs(8530) <= b;
    layer0_outputs(8531) <= not (a or b);
    layer0_outputs(8532) <= not (a xor b);
    layer0_outputs(8533) <= a and b;
    layer0_outputs(8534) <= a or b;
    layer0_outputs(8535) <= a;
    layer0_outputs(8536) <= a xor b;
    layer0_outputs(8537) <= not b;
    layer0_outputs(8538) <= not (a and b);
    layer0_outputs(8539) <= a and not b;
    layer0_outputs(8540) <= not b or a;
    layer0_outputs(8541) <= not (a or b);
    layer0_outputs(8542) <= not (a xor b);
    layer0_outputs(8543) <= a or b;
    layer0_outputs(8544) <= not (a xor b);
    layer0_outputs(8545) <= a or b;
    layer0_outputs(8546) <= a and not b;
    layer0_outputs(8547) <= not (a or b);
    layer0_outputs(8548) <= b;
    layer0_outputs(8549) <= not a;
    layer0_outputs(8550) <= b and not a;
    layer0_outputs(8551) <= not b or a;
    layer0_outputs(8552) <= not b;
    layer0_outputs(8553) <= not (a xor b);
    layer0_outputs(8554) <= not (a or b);
    layer0_outputs(8555) <= not (a xor b);
    layer0_outputs(8556) <= not (a and b);
    layer0_outputs(8557) <= a and not b;
    layer0_outputs(8558) <= a xor b;
    layer0_outputs(8559) <= a xor b;
    layer0_outputs(8560) <= not b;
    layer0_outputs(8561) <= not a;
    layer0_outputs(8562) <= a xor b;
    layer0_outputs(8563) <= b and not a;
    layer0_outputs(8564) <= a or b;
    layer0_outputs(8565) <= not a;
    layer0_outputs(8566) <= a xor b;
    layer0_outputs(8567) <= 1'b0;
    layer0_outputs(8568) <= not a;
    layer0_outputs(8569) <= not a;
    layer0_outputs(8570) <= a or b;
    layer0_outputs(8571) <= not a or b;
    layer0_outputs(8572) <= not (a and b);
    layer0_outputs(8573) <= b and not a;
    layer0_outputs(8574) <= not (a or b);
    layer0_outputs(8575) <= b and not a;
    layer0_outputs(8576) <= not (a or b);
    layer0_outputs(8577) <= not (a or b);
    layer0_outputs(8578) <= not a or b;
    layer0_outputs(8579) <= not b;
    layer0_outputs(8580) <= b and not a;
    layer0_outputs(8581) <= a xor b;
    layer0_outputs(8582) <= b and not a;
    layer0_outputs(8583) <= 1'b1;
    layer0_outputs(8584) <= not (a or b);
    layer0_outputs(8585) <= not (a xor b);
    layer0_outputs(8586) <= not (a xor b);
    layer0_outputs(8587) <= not b;
    layer0_outputs(8588) <= b;
    layer0_outputs(8589) <= not (a or b);
    layer0_outputs(8590) <= b and not a;
    layer0_outputs(8591) <= 1'b0;
    layer0_outputs(8592) <= a and not b;
    layer0_outputs(8593) <= not b or a;
    layer0_outputs(8594) <= b;
    layer0_outputs(8595) <= not a;
    layer0_outputs(8596) <= a or b;
    layer0_outputs(8597) <= a and not b;
    layer0_outputs(8598) <= b;
    layer0_outputs(8599) <= a;
    layer0_outputs(8600) <= a xor b;
    layer0_outputs(8601) <= not b;
    layer0_outputs(8602) <= b and not a;
    layer0_outputs(8603) <= not (a or b);
    layer0_outputs(8604) <= not a or b;
    layer0_outputs(8605) <= a and not b;
    layer0_outputs(8606) <= not a;
    layer0_outputs(8607) <= not b;
    layer0_outputs(8608) <= not b or a;
    layer0_outputs(8609) <= a xor b;
    layer0_outputs(8610) <= a and not b;
    layer0_outputs(8611) <= not a;
    layer0_outputs(8612) <= not (a xor b);
    layer0_outputs(8613) <= a or b;
    layer0_outputs(8614) <= not a;
    layer0_outputs(8615) <= not b;
    layer0_outputs(8616) <= a or b;
    layer0_outputs(8617) <= not b;
    layer0_outputs(8618) <= not a;
    layer0_outputs(8619) <= not (a xor b);
    layer0_outputs(8620) <= not (a xor b);
    layer0_outputs(8621) <= not (a xor b);
    layer0_outputs(8622) <= b;
    layer0_outputs(8623) <= a or b;
    layer0_outputs(8624) <= not (a or b);
    layer0_outputs(8625) <= not (a xor b);
    layer0_outputs(8626) <= a and not b;
    layer0_outputs(8627) <= not (a or b);
    layer0_outputs(8628) <= a;
    layer0_outputs(8629) <= not a;
    layer0_outputs(8630) <= a;
    layer0_outputs(8631) <= a xor b;
    layer0_outputs(8632) <= not (a or b);
    layer0_outputs(8633) <= 1'b1;
    layer0_outputs(8634) <= not (a or b);
    layer0_outputs(8635) <= not b;
    layer0_outputs(8636) <= a or b;
    layer0_outputs(8637) <= a;
    layer0_outputs(8638) <= not (a and b);
    layer0_outputs(8639) <= a xor b;
    layer0_outputs(8640) <= not a or b;
    layer0_outputs(8641) <= b and not a;
    layer0_outputs(8642) <= not (a or b);
    layer0_outputs(8643) <= not b;
    layer0_outputs(8644) <= b;
    layer0_outputs(8645) <= b and not a;
    layer0_outputs(8646) <= not a;
    layer0_outputs(8647) <= a xor b;
    layer0_outputs(8648) <= not a or b;
    layer0_outputs(8649) <= a or b;
    layer0_outputs(8650) <= a or b;
    layer0_outputs(8651) <= a or b;
    layer0_outputs(8652) <= a xor b;
    layer0_outputs(8653) <= a xor b;
    layer0_outputs(8654) <= a or b;
    layer0_outputs(8655) <= not (a or b);
    layer0_outputs(8656) <= not (a or b);
    layer0_outputs(8657) <= not (a or b);
    layer0_outputs(8658) <= b and not a;
    layer0_outputs(8659) <= not a;
    layer0_outputs(8660) <= not (a xor b);
    layer0_outputs(8661) <= a or b;
    layer0_outputs(8662) <= a and not b;
    layer0_outputs(8663) <= 1'b1;
    layer0_outputs(8664) <= b and not a;
    layer0_outputs(8665) <= b;
    layer0_outputs(8666) <= not b;
    layer0_outputs(8667) <= not b or a;
    layer0_outputs(8668) <= b and not a;
    layer0_outputs(8669) <= b and not a;
    layer0_outputs(8670) <= not a or b;
    layer0_outputs(8671) <= not (a xor b);
    layer0_outputs(8672) <= not (a or b);
    layer0_outputs(8673) <= not (a or b);
    layer0_outputs(8674) <= a or b;
    layer0_outputs(8675) <= not (a xor b);
    layer0_outputs(8676) <= 1'b1;
    layer0_outputs(8677) <= a;
    layer0_outputs(8678) <= a xor b;
    layer0_outputs(8679) <= b and not a;
    layer0_outputs(8680) <= a;
    layer0_outputs(8681) <= a or b;
    layer0_outputs(8682) <= not (a or b);
    layer0_outputs(8683) <= a or b;
    layer0_outputs(8684) <= b;
    layer0_outputs(8685) <= a;
    layer0_outputs(8686) <= not a;
    layer0_outputs(8687) <= a and not b;
    layer0_outputs(8688) <= not a;
    layer0_outputs(8689) <= not a;
    layer0_outputs(8690) <= b;
    layer0_outputs(8691) <= not (a or b);
    layer0_outputs(8692) <= not a;
    layer0_outputs(8693) <= not b;
    layer0_outputs(8694) <= a xor b;
    layer0_outputs(8695) <= a or b;
    layer0_outputs(8696) <= not b or a;
    layer0_outputs(8697) <= a xor b;
    layer0_outputs(8698) <= not b or a;
    layer0_outputs(8699) <= a;
    layer0_outputs(8700) <= a xor b;
    layer0_outputs(8701) <= not b;
    layer0_outputs(8702) <= not a or b;
    layer0_outputs(8703) <= a or b;
    layer0_outputs(8704) <= not b;
    layer0_outputs(8705) <= a xor b;
    layer0_outputs(8706) <= b;
    layer0_outputs(8707) <= not (a or b);
    layer0_outputs(8708) <= a xor b;
    layer0_outputs(8709) <= not b or a;
    layer0_outputs(8710) <= not (a or b);
    layer0_outputs(8711) <= not a;
    layer0_outputs(8712) <= not b or a;
    layer0_outputs(8713) <= not (a or b);
    layer0_outputs(8714) <= a and b;
    layer0_outputs(8715) <= not (a or b);
    layer0_outputs(8716) <= a or b;
    layer0_outputs(8717) <= not (a or b);
    layer0_outputs(8718) <= b and not a;
    layer0_outputs(8719) <= a xor b;
    layer0_outputs(8720) <= not a;
    layer0_outputs(8721) <= a and not b;
    layer0_outputs(8722) <= not (a xor b);
    layer0_outputs(8723) <= a;
    layer0_outputs(8724) <= not (a xor b);
    layer0_outputs(8725) <= not (a xor b);
    layer0_outputs(8726) <= a xor b;
    layer0_outputs(8727) <= a xor b;
    layer0_outputs(8728) <= a or b;
    layer0_outputs(8729) <= a or b;
    layer0_outputs(8730) <= a or b;
    layer0_outputs(8731) <= 1'b1;
    layer0_outputs(8732) <= a or b;
    layer0_outputs(8733) <= not a;
    layer0_outputs(8734) <= not (a xor b);
    layer0_outputs(8735) <= a or b;
    layer0_outputs(8736) <= not a or b;
    layer0_outputs(8737) <= not a or b;
    layer0_outputs(8738) <= a or b;
    layer0_outputs(8739) <= not b;
    layer0_outputs(8740) <= not (a or b);
    layer0_outputs(8741) <= not (a and b);
    layer0_outputs(8742) <= not (a xor b);
    layer0_outputs(8743) <= a and not b;
    layer0_outputs(8744) <= not b or a;
    layer0_outputs(8745) <= not (a xor b);
    layer0_outputs(8746) <= not a;
    layer0_outputs(8747) <= a or b;
    layer0_outputs(8748) <= b and not a;
    layer0_outputs(8749) <= a xor b;
    layer0_outputs(8750) <= not (a xor b);
    layer0_outputs(8751) <= not (a or b);
    layer0_outputs(8752) <= not b;
    layer0_outputs(8753) <= 1'b1;
    layer0_outputs(8754) <= a and b;
    layer0_outputs(8755) <= not b;
    layer0_outputs(8756) <= a;
    layer0_outputs(8757) <= a;
    layer0_outputs(8758) <= a or b;
    layer0_outputs(8759) <= 1'b1;
    layer0_outputs(8760) <= not a or b;
    layer0_outputs(8761) <= a or b;
    layer0_outputs(8762) <= b and not a;
    layer0_outputs(8763) <= a or b;
    layer0_outputs(8764) <= a and b;
    layer0_outputs(8765) <= not (a xor b);
    layer0_outputs(8766) <= a xor b;
    layer0_outputs(8767) <= not b;
    layer0_outputs(8768) <= a;
    layer0_outputs(8769) <= a;
    layer0_outputs(8770) <= a;
    layer0_outputs(8771) <= a or b;
    layer0_outputs(8772) <= not b or a;
    layer0_outputs(8773) <= not a or b;
    layer0_outputs(8774) <= a or b;
    layer0_outputs(8775) <= b;
    layer0_outputs(8776) <= b and not a;
    layer0_outputs(8777) <= not (a xor b);
    layer0_outputs(8778) <= b;
    layer0_outputs(8779) <= a xor b;
    layer0_outputs(8780) <= not (a xor b);
    layer0_outputs(8781) <= a;
    layer0_outputs(8782) <= a xor b;
    layer0_outputs(8783) <= b;
    layer0_outputs(8784) <= 1'b1;
    layer0_outputs(8785) <= b and not a;
    layer0_outputs(8786) <= b and not a;
    layer0_outputs(8787) <= not (a or b);
    layer0_outputs(8788) <= not a or b;
    layer0_outputs(8789) <= not b or a;
    layer0_outputs(8790) <= b and not a;
    layer0_outputs(8791) <= not (a xor b);
    layer0_outputs(8792) <= 1'b0;
    layer0_outputs(8793) <= a xor b;
    layer0_outputs(8794) <= a and not b;
    layer0_outputs(8795) <= not (a xor b);
    layer0_outputs(8796) <= not b or a;
    layer0_outputs(8797) <= a and not b;
    layer0_outputs(8798) <= a xor b;
    layer0_outputs(8799) <= not (a xor b);
    layer0_outputs(8800) <= not b;
    layer0_outputs(8801) <= not a or b;
    layer0_outputs(8802) <= a and b;
    layer0_outputs(8803) <= not (a xor b);
    layer0_outputs(8804) <= a and b;
    layer0_outputs(8805) <= not (a or b);
    layer0_outputs(8806) <= not (a or b);
    layer0_outputs(8807) <= not b;
    layer0_outputs(8808) <= not (a xor b);
    layer0_outputs(8809) <= a and b;
    layer0_outputs(8810) <= not a;
    layer0_outputs(8811) <= not b or a;
    layer0_outputs(8812) <= a;
    layer0_outputs(8813) <= not a or b;
    layer0_outputs(8814) <= not a;
    layer0_outputs(8815) <= a and not b;
    layer0_outputs(8816) <= not a;
    layer0_outputs(8817) <= a or b;
    layer0_outputs(8818) <= not (a or b);
    layer0_outputs(8819) <= a;
    layer0_outputs(8820) <= not a;
    layer0_outputs(8821) <= not (a xor b);
    layer0_outputs(8822) <= 1'b0;
    layer0_outputs(8823) <= a or b;
    layer0_outputs(8824) <= 1'b1;
    layer0_outputs(8825) <= b and not a;
    layer0_outputs(8826) <= not (a or b);
    layer0_outputs(8827) <= 1'b0;
    layer0_outputs(8828) <= b;
    layer0_outputs(8829) <= not a or b;
    layer0_outputs(8830) <= a and not b;
    layer0_outputs(8831) <= not a or b;
    layer0_outputs(8832) <= not (a xor b);
    layer0_outputs(8833) <= a or b;
    layer0_outputs(8834) <= not b or a;
    layer0_outputs(8835) <= not b or a;
    layer0_outputs(8836) <= b;
    layer0_outputs(8837) <= not (a xor b);
    layer0_outputs(8838) <= a or b;
    layer0_outputs(8839) <= a xor b;
    layer0_outputs(8840) <= not (a and b);
    layer0_outputs(8841) <= not (a or b);
    layer0_outputs(8842) <= a xor b;
    layer0_outputs(8843) <= a and not b;
    layer0_outputs(8844) <= a or b;
    layer0_outputs(8845) <= not (a or b);
    layer0_outputs(8846) <= a or b;
    layer0_outputs(8847) <= not b;
    layer0_outputs(8848) <= not (a or b);
    layer0_outputs(8849) <= a or b;
    layer0_outputs(8850) <= a or b;
    layer0_outputs(8851) <= not a or b;
    layer0_outputs(8852) <= b;
    layer0_outputs(8853) <= not (a or b);
    layer0_outputs(8854) <= 1'b1;
    layer0_outputs(8855) <= not a;
    layer0_outputs(8856) <= not b;
    layer0_outputs(8857) <= not a or b;
    layer0_outputs(8858) <= not (a and b);
    layer0_outputs(8859) <= not (a or b);
    layer0_outputs(8860) <= not (a or b);
    layer0_outputs(8861) <= not b or a;
    layer0_outputs(8862) <= a or b;
    layer0_outputs(8863) <= b;
    layer0_outputs(8864) <= a xor b;
    layer0_outputs(8865) <= a and not b;
    layer0_outputs(8866) <= b;
    layer0_outputs(8867) <= not (a or b);
    layer0_outputs(8868) <= a xor b;
    layer0_outputs(8869) <= b and not a;
    layer0_outputs(8870) <= b and not a;
    layer0_outputs(8871) <= not a;
    layer0_outputs(8872) <= not (a or b);
    layer0_outputs(8873) <= not (a xor b);
    layer0_outputs(8874) <= not b;
    layer0_outputs(8875) <= not b;
    layer0_outputs(8876) <= a xor b;
    layer0_outputs(8877) <= not b or a;
    layer0_outputs(8878) <= a or b;
    layer0_outputs(8879) <= a;
    layer0_outputs(8880) <= a or b;
    layer0_outputs(8881) <= b;
    layer0_outputs(8882) <= not (a or b);
    layer0_outputs(8883) <= a xor b;
    layer0_outputs(8884) <= a and not b;
    layer0_outputs(8885) <= b and not a;
    layer0_outputs(8886) <= a;
    layer0_outputs(8887) <= b and not a;
    layer0_outputs(8888) <= a and not b;
    layer0_outputs(8889) <= not (a or b);
    layer0_outputs(8890) <= not a or b;
    layer0_outputs(8891) <= not a;
    layer0_outputs(8892) <= not b;
    layer0_outputs(8893) <= not (a or b);
    layer0_outputs(8894) <= not (a xor b);
    layer0_outputs(8895) <= b;
    layer0_outputs(8896) <= a xor b;
    layer0_outputs(8897) <= not b;
    layer0_outputs(8898) <= a or b;
    layer0_outputs(8899) <= a and not b;
    layer0_outputs(8900) <= not a;
    layer0_outputs(8901) <= a xor b;
    layer0_outputs(8902) <= not a or b;
    layer0_outputs(8903) <= b;
    layer0_outputs(8904) <= a or b;
    layer0_outputs(8905) <= a xor b;
    layer0_outputs(8906) <= not b;
    layer0_outputs(8907) <= a;
    layer0_outputs(8908) <= 1'b0;
    layer0_outputs(8909) <= a and not b;
    layer0_outputs(8910) <= b and not a;
    layer0_outputs(8911) <= not (a xor b);
    layer0_outputs(8912) <= b and not a;
    layer0_outputs(8913) <= a xor b;
    layer0_outputs(8914) <= b;
    layer0_outputs(8915) <= a;
    layer0_outputs(8916) <= a xor b;
    layer0_outputs(8917) <= not (a xor b);
    layer0_outputs(8918) <= a xor b;
    layer0_outputs(8919) <= a;
    layer0_outputs(8920) <= not (a or b);
    layer0_outputs(8921) <= a xor b;
    layer0_outputs(8922) <= b;
    layer0_outputs(8923) <= a xor b;
    layer0_outputs(8924) <= a or b;
    layer0_outputs(8925) <= 1'b1;
    layer0_outputs(8926) <= b and not a;
    layer0_outputs(8927) <= not a;
    layer0_outputs(8928) <= not (a and b);
    layer0_outputs(8929) <= not (a and b);
    layer0_outputs(8930) <= a xor b;
    layer0_outputs(8931) <= b and not a;
    layer0_outputs(8932) <= not b or a;
    layer0_outputs(8933) <= 1'b0;
    layer0_outputs(8934) <= a or b;
    layer0_outputs(8935) <= a and b;
    layer0_outputs(8936) <= not (a xor b);
    layer0_outputs(8937) <= a;
    layer0_outputs(8938) <= a xor b;
    layer0_outputs(8939) <= a and not b;
    layer0_outputs(8940) <= b;
    layer0_outputs(8941) <= not a;
    layer0_outputs(8942) <= not (a or b);
    layer0_outputs(8943) <= not a;
    layer0_outputs(8944) <= not a or b;
    layer0_outputs(8945) <= not b;
    layer0_outputs(8946) <= a;
    layer0_outputs(8947) <= b and not a;
    layer0_outputs(8948) <= a and b;
    layer0_outputs(8949) <= not b;
    layer0_outputs(8950) <= not b;
    layer0_outputs(8951) <= not (a xor b);
    layer0_outputs(8952) <= 1'b0;
    layer0_outputs(8953) <= not (a or b);
    layer0_outputs(8954) <= not (a or b);
    layer0_outputs(8955) <= a xor b;
    layer0_outputs(8956) <= a and b;
    layer0_outputs(8957) <= a and not b;
    layer0_outputs(8958) <= not (a xor b);
    layer0_outputs(8959) <= a and b;
    layer0_outputs(8960) <= not a or b;
    layer0_outputs(8961) <= a;
    layer0_outputs(8962) <= b;
    layer0_outputs(8963) <= not (a or b);
    layer0_outputs(8964) <= a;
    layer0_outputs(8965) <= b and not a;
    layer0_outputs(8966) <= not (a and b);
    layer0_outputs(8967) <= a or b;
    layer0_outputs(8968) <= not a;
    layer0_outputs(8969) <= a or b;
    layer0_outputs(8970) <= a xor b;
    layer0_outputs(8971) <= a xor b;
    layer0_outputs(8972) <= not (a and b);
    layer0_outputs(8973) <= a or b;
    layer0_outputs(8974) <= not b or a;
    layer0_outputs(8975) <= not (a or b);
    layer0_outputs(8976) <= a or b;
    layer0_outputs(8977) <= not b or a;
    layer0_outputs(8978) <= b;
    layer0_outputs(8979) <= not b or a;
    layer0_outputs(8980) <= b and not a;
    layer0_outputs(8981) <= not b or a;
    layer0_outputs(8982) <= a and b;
    layer0_outputs(8983) <= b;
    layer0_outputs(8984) <= not b;
    layer0_outputs(8985) <= a and not b;
    layer0_outputs(8986) <= 1'b0;
    layer0_outputs(8987) <= b;
    layer0_outputs(8988) <= a and not b;
    layer0_outputs(8989) <= a or b;
    layer0_outputs(8990) <= b;
    layer0_outputs(8991) <= not b or a;
    layer0_outputs(8992) <= 1'b0;
    layer0_outputs(8993) <= b and not a;
    layer0_outputs(8994) <= b;
    layer0_outputs(8995) <= a;
    layer0_outputs(8996) <= not a or b;
    layer0_outputs(8997) <= not b;
    layer0_outputs(8998) <= not (a or b);
    layer0_outputs(8999) <= a and not b;
    layer0_outputs(9000) <= a xor b;
    layer0_outputs(9001) <= not b or a;
    layer0_outputs(9002) <= b;
    layer0_outputs(9003) <= b and not a;
    layer0_outputs(9004) <= not (a xor b);
    layer0_outputs(9005) <= 1'b1;
    layer0_outputs(9006) <= not a or b;
    layer0_outputs(9007) <= b;
    layer0_outputs(9008) <= not a or b;
    layer0_outputs(9009) <= not b;
    layer0_outputs(9010) <= a or b;
    layer0_outputs(9011) <= not (a xor b);
    layer0_outputs(9012) <= a and b;
    layer0_outputs(9013) <= a or b;
    layer0_outputs(9014) <= b and not a;
    layer0_outputs(9015) <= not b or a;
    layer0_outputs(9016) <= 1'b0;
    layer0_outputs(9017) <= a or b;
    layer0_outputs(9018) <= b;
    layer0_outputs(9019) <= not (a or b);
    layer0_outputs(9020) <= a or b;
    layer0_outputs(9021) <= not (a and b);
    layer0_outputs(9022) <= not a or b;
    layer0_outputs(9023) <= not b;
    layer0_outputs(9024) <= not (a xor b);
    layer0_outputs(9025) <= not a or b;
    layer0_outputs(9026) <= not b or a;
    layer0_outputs(9027) <= not b;
    layer0_outputs(9028) <= not a;
    layer0_outputs(9029) <= b and not a;
    layer0_outputs(9030) <= not (a or b);
    layer0_outputs(9031) <= not (a xor b);
    layer0_outputs(9032) <= b;
    layer0_outputs(9033) <= not a or b;
    layer0_outputs(9034) <= not b or a;
    layer0_outputs(9035) <= b;
    layer0_outputs(9036) <= not b or a;
    layer0_outputs(9037) <= not b;
    layer0_outputs(9038) <= a;
    layer0_outputs(9039) <= b and not a;
    layer0_outputs(9040) <= a and not b;
    layer0_outputs(9041) <= b and not a;
    layer0_outputs(9042) <= not b or a;
    layer0_outputs(9043) <= b and not a;
    layer0_outputs(9044) <= not b;
    layer0_outputs(9045) <= b;
    layer0_outputs(9046) <= a or b;
    layer0_outputs(9047) <= not b or a;
    layer0_outputs(9048) <= a and not b;
    layer0_outputs(9049) <= b;
    layer0_outputs(9050) <= b and not a;
    layer0_outputs(9051) <= a;
    layer0_outputs(9052) <= a;
    layer0_outputs(9053) <= not (a xor b);
    layer0_outputs(9054) <= a;
    layer0_outputs(9055) <= a or b;
    layer0_outputs(9056) <= b and not a;
    layer0_outputs(9057) <= a;
    layer0_outputs(9058) <= not (a xor b);
    layer0_outputs(9059) <= not b or a;
    layer0_outputs(9060) <= not b or a;
    layer0_outputs(9061) <= a xor b;
    layer0_outputs(9062) <= not b or a;
    layer0_outputs(9063) <= b;
    layer0_outputs(9064) <= a and not b;
    layer0_outputs(9065) <= a xor b;
    layer0_outputs(9066) <= not a or b;
    layer0_outputs(9067) <= not a or b;
    layer0_outputs(9068) <= not b or a;
    layer0_outputs(9069) <= a xor b;
    layer0_outputs(9070) <= b;
    layer0_outputs(9071) <= not a;
    layer0_outputs(9072) <= not (a xor b);
    layer0_outputs(9073) <= a;
    layer0_outputs(9074) <= 1'b0;
    layer0_outputs(9075) <= not a or b;
    layer0_outputs(9076) <= a xor b;
    layer0_outputs(9077) <= b and not a;
    layer0_outputs(9078) <= not b;
    layer0_outputs(9079) <= b;
    layer0_outputs(9080) <= a or b;
    layer0_outputs(9081) <= not b;
    layer0_outputs(9082) <= not (a or b);
    layer0_outputs(9083) <= not (a xor b);
    layer0_outputs(9084) <= a or b;
    layer0_outputs(9085) <= not (a xor b);
    layer0_outputs(9086) <= a;
    layer0_outputs(9087) <= not (a or b);
    layer0_outputs(9088) <= a xor b;
    layer0_outputs(9089) <= 1'b0;
    layer0_outputs(9090) <= not (a xor b);
    layer0_outputs(9091) <= not b or a;
    layer0_outputs(9092) <= not (a xor b);
    layer0_outputs(9093) <= a;
    layer0_outputs(9094) <= not b;
    layer0_outputs(9095) <= not (a xor b);
    layer0_outputs(9096) <= not (a xor b);
    layer0_outputs(9097) <= a xor b;
    layer0_outputs(9098) <= a xor b;
    layer0_outputs(9099) <= a or b;
    layer0_outputs(9100) <= a and not b;
    layer0_outputs(9101) <= b;
    layer0_outputs(9102) <= a xor b;
    layer0_outputs(9103) <= a or b;
    layer0_outputs(9104) <= not a;
    layer0_outputs(9105) <= a or b;
    layer0_outputs(9106) <= not (a or b);
    layer0_outputs(9107) <= not (a or b);
    layer0_outputs(9108) <= not a;
    layer0_outputs(9109) <= a;
    layer0_outputs(9110) <= not a or b;
    layer0_outputs(9111) <= a or b;
    layer0_outputs(9112) <= a and b;
    layer0_outputs(9113) <= not a or b;
    layer0_outputs(9114) <= not b;
    layer0_outputs(9115) <= not a or b;
    layer0_outputs(9116) <= a or b;
    layer0_outputs(9117) <= a or b;
    layer0_outputs(9118) <= not (a or b);
    layer0_outputs(9119) <= not (a or b);
    layer0_outputs(9120) <= not b or a;
    layer0_outputs(9121) <= a and not b;
    layer0_outputs(9122) <= a xor b;
    layer0_outputs(9123) <= not a or b;
    layer0_outputs(9124) <= not a;
    layer0_outputs(9125) <= a;
    layer0_outputs(9126) <= not a or b;
    layer0_outputs(9127) <= not (a xor b);
    layer0_outputs(9128) <= b and not a;
    layer0_outputs(9129) <= not b;
    layer0_outputs(9130) <= not b or a;
    layer0_outputs(9131) <= not b;
    layer0_outputs(9132) <= not (a or b);
    layer0_outputs(9133) <= a xor b;
    layer0_outputs(9134) <= a xor b;
    layer0_outputs(9135) <= not (a xor b);
    layer0_outputs(9136) <= not a;
    layer0_outputs(9137) <= not (a or b);
    layer0_outputs(9138) <= a or b;
    layer0_outputs(9139) <= not (a xor b);
    layer0_outputs(9140) <= a or b;
    layer0_outputs(9141) <= a or b;
    layer0_outputs(9142) <= a xor b;
    layer0_outputs(9143) <= b;
    layer0_outputs(9144) <= a xor b;
    layer0_outputs(9145) <= not a or b;
    layer0_outputs(9146) <= a xor b;
    layer0_outputs(9147) <= 1'b1;
    layer0_outputs(9148) <= a xor b;
    layer0_outputs(9149) <= a xor b;
    layer0_outputs(9150) <= not (a xor b);
    layer0_outputs(9151) <= not (a or b);
    layer0_outputs(9152) <= not a or b;
    layer0_outputs(9153) <= not (a or b);
    layer0_outputs(9154) <= a xor b;
    layer0_outputs(9155) <= a xor b;
    layer0_outputs(9156) <= b;
    layer0_outputs(9157) <= not b or a;
    layer0_outputs(9158) <= a xor b;
    layer0_outputs(9159) <= not b;
    layer0_outputs(9160) <= b;
    layer0_outputs(9161) <= a or b;
    layer0_outputs(9162) <= not (a xor b);
    layer0_outputs(9163) <= not b or a;
    layer0_outputs(9164) <= a or b;
    layer0_outputs(9165) <= 1'b1;
    layer0_outputs(9166) <= a or b;
    layer0_outputs(9167) <= not a or b;
    layer0_outputs(9168) <= not b;
    layer0_outputs(9169) <= b and not a;
    layer0_outputs(9170) <= b and not a;
    layer0_outputs(9171) <= not b;
    layer0_outputs(9172) <= b;
    layer0_outputs(9173) <= not a;
    layer0_outputs(9174) <= a or b;
    layer0_outputs(9175) <= a or b;
    layer0_outputs(9176) <= 1'b0;
    layer0_outputs(9177) <= b and not a;
    layer0_outputs(9178) <= not b or a;
    layer0_outputs(9179) <= not (a or b);
    layer0_outputs(9180) <= a and not b;
    layer0_outputs(9181) <= a or b;
    layer0_outputs(9182) <= a;
    layer0_outputs(9183) <= a and b;
    layer0_outputs(9184) <= 1'b0;
    layer0_outputs(9185) <= not (a or b);
    layer0_outputs(9186) <= not (a or b);
    layer0_outputs(9187) <= a or b;
    layer0_outputs(9188) <= not a;
    layer0_outputs(9189) <= not (a or b);
    layer0_outputs(9190) <= not (a xor b);
    layer0_outputs(9191) <= not a or b;
    layer0_outputs(9192) <= a or b;
    layer0_outputs(9193) <= a or b;
    layer0_outputs(9194) <= a and not b;
    layer0_outputs(9195) <= b and not a;
    layer0_outputs(9196) <= a or b;
    layer0_outputs(9197) <= b and not a;
    layer0_outputs(9198) <= a xor b;
    layer0_outputs(9199) <= not (a xor b);
    layer0_outputs(9200) <= a;
    layer0_outputs(9201) <= a or b;
    layer0_outputs(9202) <= not b or a;
    layer0_outputs(9203) <= not a;
    layer0_outputs(9204) <= not b or a;
    layer0_outputs(9205) <= b and not a;
    layer0_outputs(9206) <= not b or a;
    layer0_outputs(9207) <= not (a or b);
    layer0_outputs(9208) <= not a;
    layer0_outputs(9209) <= b and not a;
    layer0_outputs(9210) <= a;
    layer0_outputs(9211) <= b;
    layer0_outputs(9212) <= not (a xor b);
    layer0_outputs(9213) <= not (a or b);
    layer0_outputs(9214) <= a;
    layer0_outputs(9215) <= not (a or b);
    layer0_outputs(9216) <= not b;
    layer0_outputs(9217) <= a or b;
    layer0_outputs(9218) <= not (a xor b);
    layer0_outputs(9219) <= not a or b;
    layer0_outputs(9220) <= not b;
    layer0_outputs(9221) <= not (a xor b);
    layer0_outputs(9222) <= a;
    layer0_outputs(9223) <= not (a and b);
    layer0_outputs(9224) <= not (a or b);
    layer0_outputs(9225) <= not b or a;
    layer0_outputs(9226) <= a xor b;
    layer0_outputs(9227) <= a or b;
    layer0_outputs(9228) <= a and not b;
    layer0_outputs(9229) <= a or b;
    layer0_outputs(9230) <= a xor b;
    layer0_outputs(9231) <= b and not a;
    layer0_outputs(9232) <= a;
    layer0_outputs(9233) <= not a;
    layer0_outputs(9234) <= not (a xor b);
    layer0_outputs(9235) <= a or b;
    layer0_outputs(9236) <= 1'b0;
    layer0_outputs(9237) <= a xor b;
    layer0_outputs(9238) <= a or b;
    layer0_outputs(9239) <= not (a or b);
    layer0_outputs(9240) <= not (a or b);
    layer0_outputs(9241) <= not b or a;
    layer0_outputs(9242) <= b and not a;
    layer0_outputs(9243) <= not (a or b);
    layer0_outputs(9244) <= a and not b;
    layer0_outputs(9245) <= b and not a;
    layer0_outputs(9246) <= b;
    layer0_outputs(9247) <= a or b;
    layer0_outputs(9248) <= a;
    layer0_outputs(9249) <= b and not a;
    layer0_outputs(9250) <= not b;
    layer0_outputs(9251) <= a or b;
    layer0_outputs(9252) <= not (a xor b);
    layer0_outputs(9253) <= not a or b;
    layer0_outputs(9254) <= not (a xor b);
    layer0_outputs(9255) <= not a;
    layer0_outputs(9256) <= a xor b;
    layer0_outputs(9257) <= a xor b;
    layer0_outputs(9258) <= a and not b;
    layer0_outputs(9259) <= not b;
    layer0_outputs(9260) <= a and not b;
    layer0_outputs(9261) <= not a or b;
    layer0_outputs(9262) <= a or b;
    layer0_outputs(9263) <= a and not b;
    layer0_outputs(9264) <= not (a or b);
    layer0_outputs(9265) <= a or b;
    layer0_outputs(9266) <= b;
    layer0_outputs(9267) <= not (a and b);
    layer0_outputs(9268) <= a;
    layer0_outputs(9269) <= a or b;
    layer0_outputs(9270) <= a or b;
    layer0_outputs(9271) <= 1'b0;
    layer0_outputs(9272) <= not b or a;
    layer0_outputs(9273) <= not (a or b);
    layer0_outputs(9274) <= not (a or b);
    layer0_outputs(9275) <= not b or a;
    layer0_outputs(9276) <= not (a and b);
    layer0_outputs(9277) <= not (a xor b);
    layer0_outputs(9278) <= a or b;
    layer0_outputs(9279) <= not (a or b);
    layer0_outputs(9280) <= a or b;
    layer0_outputs(9281) <= a or b;
    layer0_outputs(9282) <= a or b;
    layer0_outputs(9283) <= not a or b;
    layer0_outputs(9284) <= not b;
    layer0_outputs(9285) <= a and not b;
    layer0_outputs(9286) <= a and not b;
    layer0_outputs(9287) <= not (a xor b);
    layer0_outputs(9288) <= a and not b;
    layer0_outputs(9289) <= a xor b;
    layer0_outputs(9290) <= a and not b;
    layer0_outputs(9291) <= not (a xor b);
    layer0_outputs(9292) <= not (a xor b);
    layer0_outputs(9293) <= not b or a;
    layer0_outputs(9294) <= a xor b;
    layer0_outputs(9295) <= a and not b;
    layer0_outputs(9296) <= not (a or b);
    layer0_outputs(9297) <= not (a or b);
    layer0_outputs(9298) <= a and not b;
    layer0_outputs(9299) <= a and not b;
    layer0_outputs(9300) <= a xor b;
    layer0_outputs(9301) <= a or b;
    layer0_outputs(9302) <= a xor b;
    layer0_outputs(9303) <= a xor b;
    layer0_outputs(9304) <= a or b;
    layer0_outputs(9305) <= not (a xor b);
    layer0_outputs(9306) <= not (a and b);
    layer0_outputs(9307) <= a or b;
    layer0_outputs(9308) <= not a or b;
    layer0_outputs(9309) <= a;
    layer0_outputs(9310) <= a or b;
    layer0_outputs(9311) <= a xor b;
    layer0_outputs(9312) <= not (a or b);
    layer0_outputs(9313) <= not a;
    layer0_outputs(9314) <= a xor b;
    layer0_outputs(9315) <= a;
    layer0_outputs(9316) <= not (a xor b);
    layer0_outputs(9317) <= b;
    layer0_outputs(9318) <= not b;
    layer0_outputs(9319) <= 1'b0;
    layer0_outputs(9320) <= not (a xor b);
    layer0_outputs(9321) <= not b or a;
    layer0_outputs(9322) <= not (a or b);
    layer0_outputs(9323) <= not a;
    layer0_outputs(9324) <= not (a or b);
    layer0_outputs(9325) <= not (a xor b);
    layer0_outputs(9326) <= a or b;
    layer0_outputs(9327) <= a;
    layer0_outputs(9328) <= a or b;
    layer0_outputs(9329) <= a and b;
    layer0_outputs(9330) <= not (a xor b);
    layer0_outputs(9331) <= not a or b;
    layer0_outputs(9332) <= not b;
    layer0_outputs(9333) <= a or b;
    layer0_outputs(9334) <= b;
    layer0_outputs(9335) <= a and b;
    layer0_outputs(9336) <= a;
    layer0_outputs(9337) <= not (a xor b);
    layer0_outputs(9338) <= not (a or b);
    layer0_outputs(9339) <= a;
    layer0_outputs(9340) <= not (a or b);
    layer0_outputs(9341) <= a or b;
    layer0_outputs(9342) <= not a;
    layer0_outputs(9343) <= not b or a;
    layer0_outputs(9344) <= not (a or b);
    layer0_outputs(9345) <= not (a xor b);
    layer0_outputs(9346) <= not (a xor b);
    layer0_outputs(9347) <= b;
    layer0_outputs(9348) <= a or b;
    layer0_outputs(9349) <= not (a and b);
    layer0_outputs(9350) <= b and not a;
    layer0_outputs(9351) <= b;
    layer0_outputs(9352) <= not a;
    layer0_outputs(9353) <= a xor b;
    layer0_outputs(9354) <= not b;
    layer0_outputs(9355) <= a and not b;
    layer0_outputs(9356) <= not (a xor b);
    layer0_outputs(9357) <= a xor b;
    layer0_outputs(9358) <= b and not a;
    layer0_outputs(9359) <= a or b;
    layer0_outputs(9360) <= not (a xor b);
    layer0_outputs(9361) <= 1'b0;
    layer0_outputs(9362) <= a or b;
    layer0_outputs(9363) <= a or b;
    layer0_outputs(9364) <= a;
    layer0_outputs(9365) <= b;
    layer0_outputs(9366) <= b;
    layer0_outputs(9367) <= not (a or b);
    layer0_outputs(9368) <= not (a or b);
    layer0_outputs(9369) <= a xor b;
    layer0_outputs(9370) <= not (a or b);
    layer0_outputs(9371) <= not (a or b);
    layer0_outputs(9372) <= a or b;
    layer0_outputs(9373) <= not (a xor b);
    layer0_outputs(9374) <= not b or a;
    layer0_outputs(9375) <= not (a xor b);
    layer0_outputs(9376) <= a or b;
    layer0_outputs(9377) <= not a;
    layer0_outputs(9378) <= not (a xor b);
    layer0_outputs(9379) <= not b;
    layer0_outputs(9380) <= not (a or b);
    layer0_outputs(9381) <= not (a or b);
    layer0_outputs(9382) <= b and not a;
    layer0_outputs(9383) <= not b;
    layer0_outputs(9384) <= a xor b;
    layer0_outputs(9385) <= not (a or b);
    layer0_outputs(9386) <= not b or a;
    layer0_outputs(9387) <= b and not a;
    layer0_outputs(9388) <= a;
    layer0_outputs(9389) <= not b;
    layer0_outputs(9390) <= not b or a;
    layer0_outputs(9391) <= not (a xor b);
    layer0_outputs(9392) <= a or b;
    layer0_outputs(9393) <= not a or b;
    layer0_outputs(9394) <= a or b;
    layer0_outputs(9395) <= not a;
    layer0_outputs(9396) <= a and not b;
    layer0_outputs(9397) <= not a or b;
    layer0_outputs(9398) <= a and b;
    layer0_outputs(9399) <= b and not a;
    layer0_outputs(9400) <= 1'b1;
    layer0_outputs(9401) <= a or b;
    layer0_outputs(9402) <= not a;
    layer0_outputs(9403) <= a xor b;
    layer0_outputs(9404) <= a or b;
    layer0_outputs(9405) <= not a;
    layer0_outputs(9406) <= b and not a;
    layer0_outputs(9407) <= not a or b;
    layer0_outputs(9408) <= not (a or b);
    layer0_outputs(9409) <= not (a xor b);
    layer0_outputs(9410) <= not b;
    layer0_outputs(9411) <= not (a and b);
    layer0_outputs(9412) <= a or b;
    layer0_outputs(9413) <= a and b;
    layer0_outputs(9414) <= b;
    layer0_outputs(9415) <= a and not b;
    layer0_outputs(9416) <= 1'b0;
    layer0_outputs(9417) <= not (a and b);
    layer0_outputs(9418) <= not b or a;
    layer0_outputs(9419) <= not a or b;
    layer0_outputs(9420) <= a and b;
    layer0_outputs(9421) <= not (a xor b);
    layer0_outputs(9422) <= a or b;
    layer0_outputs(9423) <= not (a or b);
    layer0_outputs(9424) <= not (a xor b);
    layer0_outputs(9425) <= b;
    layer0_outputs(9426) <= a or b;
    layer0_outputs(9427) <= not (a or b);
    layer0_outputs(9428) <= not (a or b);
    layer0_outputs(9429) <= a xor b;
    layer0_outputs(9430) <= b and not a;
    layer0_outputs(9431) <= not (a xor b);
    layer0_outputs(9432) <= not (a or b);
    layer0_outputs(9433) <= not a;
    layer0_outputs(9434) <= a or b;
    layer0_outputs(9435) <= not b or a;
    layer0_outputs(9436) <= not (a xor b);
    layer0_outputs(9437) <= not b;
    layer0_outputs(9438) <= not (a xor b);
    layer0_outputs(9439) <= not b or a;
    layer0_outputs(9440) <= not b;
    layer0_outputs(9441) <= not a;
    layer0_outputs(9442) <= not b or a;
    layer0_outputs(9443) <= not (a xor b);
    layer0_outputs(9444) <= b;
    layer0_outputs(9445) <= not (a or b);
    layer0_outputs(9446) <= not (a or b);
    layer0_outputs(9447) <= b and not a;
    layer0_outputs(9448) <= a or b;
    layer0_outputs(9449) <= a xor b;
    layer0_outputs(9450) <= not (a and b);
    layer0_outputs(9451) <= not (a xor b);
    layer0_outputs(9452) <= a;
    layer0_outputs(9453) <= a and not b;
    layer0_outputs(9454) <= a or b;
    layer0_outputs(9455) <= a or b;
    layer0_outputs(9456) <= not (a or b);
    layer0_outputs(9457) <= not a or b;
    layer0_outputs(9458) <= not a;
    layer0_outputs(9459) <= not (a xor b);
    layer0_outputs(9460) <= a or b;
    layer0_outputs(9461) <= a or b;
    layer0_outputs(9462) <= b;
    layer0_outputs(9463) <= not (a xor b);
    layer0_outputs(9464) <= not (a xor b);
    layer0_outputs(9465) <= not (a or b);
    layer0_outputs(9466) <= not (a and b);
    layer0_outputs(9467) <= 1'b0;
    layer0_outputs(9468) <= 1'b0;
    layer0_outputs(9469) <= a or b;
    layer0_outputs(9470) <= not (a or b);
    layer0_outputs(9471) <= not b or a;
    layer0_outputs(9472) <= a or b;
    layer0_outputs(9473) <= b;
    layer0_outputs(9474) <= not (a or b);
    layer0_outputs(9475) <= 1'b0;
    layer0_outputs(9476) <= a;
    layer0_outputs(9477) <= b;
    layer0_outputs(9478) <= not a;
    layer0_outputs(9479) <= not (a or b);
    layer0_outputs(9480) <= b and not a;
    layer0_outputs(9481) <= a;
    layer0_outputs(9482) <= not (a or b);
    layer0_outputs(9483) <= b;
    layer0_outputs(9484) <= a and not b;
    layer0_outputs(9485) <= a and not b;
    layer0_outputs(9486) <= a or b;
    layer0_outputs(9487) <= not (a or b);
    layer0_outputs(9488) <= a;
    layer0_outputs(9489) <= a xor b;
    layer0_outputs(9490) <= not b or a;
    layer0_outputs(9491) <= not (a or b);
    layer0_outputs(9492) <= a and b;
    layer0_outputs(9493) <= b;
    layer0_outputs(9494) <= a xor b;
    layer0_outputs(9495) <= not (a or b);
    layer0_outputs(9496) <= not b;
    layer0_outputs(9497) <= not (a xor b);
    layer0_outputs(9498) <= a;
    layer0_outputs(9499) <= a and b;
    layer0_outputs(9500) <= a and not b;
    layer0_outputs(9501) <= not (a or b);
    layer0_outputs(9502) <= not (a xor b);
    layer0_outputs(9503) <= b;
    layer0_outputs(9504) <= 1'b0;
    layer0_outputs(9505) <= 1'b0;
    layer0_outputs(9506) <= not (a xor b);
    layer0_outputs(9507) <= not a or b;
    layer0_outputs(9508) <= 1'b0;
    layer0_outputs(9509) <= not (a or b);
    layer0_outputs(9510) <= not (a or b);
    layer0_outputs(9511) <= a and not b;
    layer0_outputs(9512) <= a and b;
    layer0_outputs(9513) <= a or b;
    layer0_outputs(9514) <= 1'b0;
    layer0_outputs(9515) <= not b;
    layer0_outputs(9516) <= not (a or b);
    layer0_outputs(9517) <= b;
    layer0_outputs(9518) <= a xor b;
    layer0_outputs(9519) <= not a;
    layer0_outputs(9520) <= not (a xor b);
    layer0_outputs(9521) <= a;
    layer0_outputs(9522) <= not (a xor b);
    layer0_outputs(9523) <= not b;
    layer0_outputs(9524) <= b;
    layer0_outputs(9525) <= not (a or b);
    layer0_outputs(9526) <= b;
    layer0_outputs(9527) <= not (a or b);
    layer0_outputs(9528) <= not (a xor b);
    layer0_outputs(9529) <= not a;
    layer0_outputs(9530) <= b;
    layer0_outputs(9531) <= a and b;
    layer0_outputs(9532) <= a or b;
    layer0_outputs(9533) <= not b or a;
    layer0_outputs(9534) <= not b or a;
    layer0_outputs(9535) <= a;
    layer0_outputs(9536) <= not (a xor b);
    layer0_outputs(9537) <= b and not a;
    layer0_outputs(9538) <= a or b;
    layer0_outputs(9539) <= a and not b;
    layer0_outputs(9540) <= not a;
    layer0_outputs(9541) <= not b;
    layer0_outputs(9542) <= not a or b;
    layer0_outputs(9543) <= a xor b;
    layer0_outputs(9544) <= not (a xor b);
    layer0_outputs(9545) <= 1'b0;
    layer0_outputs(9546) <= a or b;
    layer0_outputs(9547) <= b;
    layer0_outputs(9548) <= b and not a;
    layer0_outputs(9549) <= b;
    layer0_outputs(9550) <= not a or b;
    layer0_outputs(9551) <= not (a xor b);
    layer0_outputs(9552) <= a xor b;
    layer0_outputs(9553) <= b;
    layer0_outputs(9554) <= not b or a;
    layer0_outputs(9555) <= not (a or b);
    layer0_outputs(9556) <= a or b;
    layer0_outputs(9557) <= a xor b;
    layer0_outputs(9558) <= not (a or b);
    layer0_outputs(9559) <= a and not b;
    layer0_outputs(9560) <= not (a or b);
    layer0_outputs(9561) <= b;
    layer0_outputs(9562) <= not (a or b);
    layer0_outputs(9563) <= 1'b1;
    layer0_outputs(9564) <= not a;
    layer0_outputs(9565) <= 1'b0;
    layer0_outputs(9566) <= a or b;
    layer0_outputs(9567) <= not (a xor b);
    layer0_outputs(9568) <= not (a xor b);
    layer0_outputs(9569) <= a xor b;
    layer0_outputs(9570) <= a xor b;
    layer0_outputs(9571) <= a and b;
    layer0_outputs(9572) <= a xor b;
    layer0_outputs(9573) <= not a;
    layer0_outputs(9574) <= a or b;
    layer0_outputs(9575) <= a xor b;
    layer0_outputs(9576) <= b and not a;
    layer0_outputs(9577) <= a and b;
    layer0_outputs(9578) <= 1'b1;
    layer0_outputs(9579) <= not a or b;
    layer0_outputs(9580) <= b;
    layer0_outputs(9581) <= a or b;
    layer0_outputs(9582) <= b;
    layer0_outputs(9583) <= not (a xor b);
    layer0_outputs(9584) <= a and not b;
    layer0_outputs(9585) <= not a;
    layer0_outputs(9586) <= not a or b;
    layer0_outputs(9587) <= not (a xor b);
    layer0_outputs(9588) <= not (a xor b);
    layer0_outputs(9589) <= a xor b;
    layer0_outputs(9590) <= not (a xor b);
    layer0_outputs(9591) <= a or b;
    layer0_outputs(9592) <= b;
    layer0_outputs(9593) <= b and not a;
    layer0_outputs(9594) <= b;
    layer0_outputs(9595) <= b and not a;
    layer0_outputs(9596) <= b and not a;
    layer0_outputs(9597) <= b;
    layer0_outputs(9598) <= a;
    layer0_outputs(9599) <= b and not a;
    layer0_outputs(9600) <= not b;
    layer0_outputs(9601) <= a or b;
    layer0_outputs(9602) <= 1'b0;
    layer0_outputs(9603) <= 1'b1;
    layer0_outputs(9604) <= not b;
    layer0_outputs(9605) <= not a;
    layer0_outputs(9606) <= a or b;
    layer0_outputs(9607) <= a;
    layer0_outputs(9608) <= not (a xor b);
    layer0_outputs(9609) <= not (a or b);
    layer0_outputs(9610) <= b and not a;
    layer0_outputs(9611) <= a xor b;
    layer0_outputs(9612) <= 1'b0;
    layer0_outputs(9613) <= b;
    layer0_outputs(9614) <= b and not a;
    layer0_outputs(9615) <= b;
    layer0_outputs(9616) <= not b;
    layer0_outputs(9617) <= not (a xor b);
    layer0_outputs(9618) <= not a;
    layer0_outputs(9619) <= not (a xor b);
    layer0_outputs(9620) <= a or b;
    layer0_outputs(9621) <= not a;
    layer0_outputs(9622) <= not (a or b);
    layer0_outputs(9623) <= not (a xor b);
    layer0_outputs(9624) <= not (a or b);
    layer0_outputs(9625) <= b;
    layer0_outputs(9626) <= not a;
    layer0_outputs(9627) <= a or b;
    layer0_outputs(9628) <= a xor b;
    layer0_outputs(9629) <= not (a or b);
    layer0_outputs(9630) <= 1'b1;
    layer0_outputs(9631) <= a xor b;
    layer0_outputs(9632) <= a xor b;
    layer0_outputs(9633) <= not (a or b);
    layer0_outputs(9634) <= a or b;
    layer0_outputs(9635) <= a or b;
    layer0_outputs(9636) <= not (a xor b);
    layer0_outputs(9637) <= a or b;
    layer0_outputs(9638) <= a or b;
    layer0_outputs(9639) <= b and not a;
    layer0_outputs(9640) <= 1'b1;
    layer0_outputs(9641) <= not (a xor b);
    layer0_outputs(9642) <= not b;
    layer0_outputs(9643) <= a or b;
    layer0_outputs(9644) <= not (a or b);
    layer0_outputs(9645) <= b;
    layer0_outputs(9646) <= not (a xor b);
    layer0_outputs(9647) <= not (a or b);
    layer0_outputs(9648) <= b and not a;
    layer0_outputs(9649) <= not a or b;
    layer0_outputs(9650) <= not (a xor b);
    layer0_outputs(9651) <= a;
    layer0_outputs(9652) <= b and not a;
    layer0_outputs(9653) <= a xor b;
    layer0_outputs(9654) <= a and not b;
    layer0_outputs(9655) <= a xor b;
    layer0_outputs(9656) <= a and not b;
    layer0_outputs(9657) <= not (a xor b);
    layer0_outputs(9658) <= not b;
    layer0_outputs(9659) <= not b or a;
    layer0_outputs(9660) <= not a;
    layer0_outputs(9661) <= not (a or b);
    layer0_outputs(9662) <= not (a or b);
    layer0_outputs(9663) <= a and b;
    layer0_outputs(9664) <= b and not a;
    layer0_outputs(9665) <= not (a xor b);
    layer0_outputs(9666) <= a or b;
    layer0_outputs(9667) <= a or b;
    layer0_outputs(9668) <= a or b;
    layer0_outputs(9669) <= a or b;
    layer0_outputs(9670) <= not b or a;
    layer0_outputs(9671) <= a or b;
    layer0_outputs(9672) <= not (a and b);
    layer0_outputs(9673) <= not (a and b);
    layer0_outputs(9674) <= not b or a;
    layer0_outputs(9675) <= a xor b;
    layer0_outputs(9676) <= not a or b;
    layer0_outputs(9677) <= not a;
    layer0_outputs(9678) <= not a or b;
    layer0_outputs(9679) <= not (a or b);
    layer0_outputs(9680) <= not (a or b);
    layer0_outputs(9681) <= a or b;
    layer0_outputs(9682) <= b and not a;
    layer0_outputs(9683) <= not a or b;
    layer0_outputs(9684) <= a xor b;
    layer0_outputs(9685) <= not (a or b);
    layer0_outputs(9686) <= a or b;
    layer0_outputs(9687) <= a;
    layer0_outputs(9688) <= b;
    layer0_outputs(9689) <= a or b;
    layer0_outputs(9690) <= a or b;
    layer0_outputs(9691) <= not b;
    layer0_outputs(9692) <= a or b;
    layer0_outputs(9693) <= a xor b;
    layer0_outputs(9694) <= a and not b;
    layer0_outputs(9695) <= a or b;
    layer0_outputs(9696) <= a xor b;
    layer0_outputs(9697) <= not b;
    layer0_outputs(9698) <= not a;
    layer0_outputs(9699) <= b;
    layer0_outputs(9700) <= not a;
    layer0_outputs(9701) <= not b or a;
    layer0_outputs(9702) <= not (a or b);
    layer0_outputs(9703) <= b;
    layer0_outputs(9704) <= not (a or b);
    layer0_outputs(9705) <= a xor b;
    layer0_outputs(9706) <= not b or a;
    layer0_outputs(9707) <= a or b;
    layer0_outputs(9708) <= 1'b0;
    layer0_outputs(9709) <= not (a or b);
    layer0_outputs(9710) <= not (a or b);
    layer0_outputs(9711) <= a xor b;
    layer0_outputs(9712) <= a xor b;
    layer0_outputs(9713) <= a or b;
    layer0_outputs(9714) <= a or b;
    layer0_outputs(9715) <= not (a or b);
    layer0_outputs(9716) <= not b or a;
    layer0_outputs(9717) <= not b;
    layer0_outputs(9718) <= not a or b;
    layer0_outputs(9719) <= 1'b1;
    layer0_outputs(9720) <= a and not b;
    layer0_outputs(9721) <= not (a xor b);
    layer0_outputs(9722) <= not (a xor b);
    layer0_outputs(9723) <= not b or a;
    layer0_outputs(9724) <= a or b;
    layer0_outputs(9725) <= not b or a;
    layer0_outputs(9726) <= not b or a;
    layer0_outputs(9727) <= a and not b;
    layer0_outputs(9728) <= a and not b;
    layer0_outputs(9729) <= b;
    layer0_outputs(9730) <= b;
    layer0_outputs(9731) <= not (a or b);
    layer0_outputs(9732) <= a or b;
    layer0_outputs(9733) <= a;
    layer0_outputs(9734) <= not a or b;
    layer0_outputs(9735) <= a and not b;
    layer0_outputs(9736) <= not a or b;
    layer0_outputs(9737) <= a and b;
    layer0_outputs(9738) <= a xor b;
    layer0_outputs(9739) <= not (a or b);
    layer0_outputs(9740) <= not (a xor b);
    layer0_outputs(9741) <= not a;
    layer0_outputs(9742) <= not (a or b);
    layer0_outputs(9743) <= a;
    layer0_outputs(9744) <= a or b;
    layer0_outputs(9745) <= not b or a;
    layer0_outputs(9746) <= a or b;
    layer0_outputs(9747) <= not (a or b);
    layer0_outputs(9748) <= 1'b0;
    layer0_outputs(9749) <= not (a xor b);
    layer0_outputs(9750) <= not a;
    layer0_outputs(9751) <= not (a xor b);
    layer0_outputs(9752) <= b and not a;
    layer0_outputs(9753) <= not (a or b);
    layer0_outputs(9754) <= not (a xor b);
    layer0_outputs(9755) <= not (a or b);
    layer0_outputs(9756) <= a or b;
    layer0_outputs(9757) <= a or b;
    layer0_outputs(9758) <= 1'b1;
    layer0_outputs(9759) <= a;
    layer0_outputs(9760) <= a xor b;
    layer0_outputs(9761) <= a or b;
    layer0_outputs(9762) <= not (a xor b);
    layer0_outputs(9763) <= not (a or b);
    layer0_outputs(9764) <= not b;
    layer0_outputs(9765) <= not a or b;
    layer0_outputs(9766) <= a xor b;
    layer0_outputs(9767) <= not (a or b);
    layer0_outputs(9768) <= not (a or b);
    layer0_outputs(9769) <= not (a or b);
    layer0_outputs(9770) <= not (a or b);
    layer0_outputs(9771) <= not (a xor b);
    layer0_outputs(9772) <= b;
    layer0_outputs(9773) <= b;
    layer0_outputs(9774) <= not (a xor b);
    layer0_outputs(9775) <= b and not a;
    layer0_outputs(9776) <= not a or b;
    layer0_outputs(9777) <= a and not b;
    layer0_outputs(9778) <= a and not b;
    layer0_outputs(9779) <= a or b;
    layer0_outputs(9780) <= a and b;
    layer0_outputs(9781) <= b and not a;
    layer0_outputs(9782) <= a or b;
    layer0_outputs(9783) <= not b or a;
    layer0_outputs(9784) <= a and not b;
    layer0_outputs(9785) <= a xor b;
    layer0_outputs(9786) <= not a or b;
    layer0_outputs(9787) <= not b;
    layer0_outputs(9788) <= a or b;
    layer0_outputs(9789) <= not (a or b);
    layer0_outputs(9790) <= not a or b;
    layer0_outputs(9791) <= not (a xor b);
    layer0_outputs(9792) <= 1'b0;
    layer0_outputs(9793) <= not b;
    layer0_outputs(9794) <= b and not a;
    layer0_outputs(9795) <= a and not b;
    layer0_outputs(9796) <= a or b;
    layer0_outputs(9797) <= not b or a;
    layer0_outputs(9798) <= a xor b;
    layer0_outputs(9799) <= not (a xor b);
    layer0_outputs(9800) <= a or b;
    layer0_outputs(9801) <= not b;
    layer0_outputs(9802) <= b and not a;
    layer0_outputs(9803) <= b;
    layer0_outputs(9804) <= not b;
    layer0_outputs(9805) <= a or b;
    layer0_outputs(9806) <= not (a xor b);
    layer0_outputs(9807) <= b and not a;
    layer0_outputs(9808) <= a xor b;
    layer0_outputs(9809) <= not a;
    layer0_outputs(9810) <= not (a or b);
    layer0_outputs(9811) <= a;
    layer0_outputs(9812) <= b;
    layer0_outputs(9813) <= not b;
    layer0_outputs(9814) <= not a;
    layer0_outputs(9815) <= not b;
    layer0_outputs(9816) <= a or b;
    layer0_outputs(9817) <= not (a or b);
    layer0_outputs(9818) <= a;
    layer0_outputs(9819) <= not a;
    layer0_outputs(9820) <= a and not b;
    layer0_outputs(9821) <= a xor b;
    layer0_outputs(9822) <= a and not b;
    layer0_outputs(9823) <= a or b;
    layer0_outputs(9824) <= not (a xor b);
    layer0_outputs(9825) <= not (a or b);
    layer0_outputs(9826) <= a or b;
    layer0_outputs(9827) <= not (a xor b);
    layer0_outputs(9828) <= a or b;
    layer0_outputs(9829) <= 1'b0;
    layer0_outputs(9830) <= b;
    layer0_outputs(9831) <= a;
    layer0_outputs(9832) <= not b or a;
    layer0_outputs(9833) <= not a;
    layer0_outputs(9834) <= not a;
    layer0_outputs(9835) <= a xor b;
    layer0_outputs(9836) <= a;
    layer0_outputs(9837) <= a xor b;
    layer0_outputs(9838) <= not b;
    layer0_outputs(9839) <= a or b;
    layer0_outputs(9840) <= a;
    layer0_outputs(9841) <= b and not a;
    layer0_outputs(9842) <= a;
    layer0_outputs(9843) <= not (a or b);
    layer0_outputs(9844) <= not b;
    layer0_outputs(9845) <= b and not a;
    layer0_outputs(9846) <= a and b;
    layer0_outputs(9847) <= not (a and b);
    layer0_outputs(9848) <= not (a xor b);
    layer0_outputs(9849) <= not b;
    layer0_outputs(9850) <= b;
    layer0_outputs(9851) <= not (a xor b);
    layer0_outputs(9852) <= a;
    layer0_outputs(9853) <= not (a xor b);
    layer0_outputs(9854) <= a and b;
    layer0_outputs(9855) <= not a;
    layer0_outputs(9856) <= a xor b;
    layer0_outputs(9857) <= a or b;
    layer0_outputs(9858) <= not (a or b);
    layer0_outputs(9859) <= not a or b;
    layer0_outputs(9860) <= not b or a;
    layer0_outputs(9861) <= 1'b0;
    layer0_outputs(9862) <= 1'b0;
    layer0_outputs(9863) <= b;
    layer0_outputs(9864) <= 1'b0;
    layer0_outputs(9865) <= not (a or b);
    layer0_outputs(9866) <= a xor b;
    layer0_outputs(9867) <= not (a xor b);
    layer0_outputs(9868) <= b and not a;
    layer0_outputs(9869) <= a or b;
    layer0_outputs(9870) <= not a;
    layer0_outputs(9871) <= not (a xor b);
    layer0_outputs(9872) <= a or b;
    layer0_outputs(9873) <= b;
    layer0_outputs(9874) <= not (a or b);
    layer0_outputs(9875) <= a;
    layer0_outputs(9876) <= not (a xor b);
    layer0_outputs(9877) <= not b;
    layer0_outputs(9878) <= a xor b;
    layer0_outputs(9879) <= not (a or b);
    layer0_outputs(9880) <= a xor b;
    layer0_outputs(9881) <= a;
    layer0_outputs(9882) <= not (a or b);
    layer0_outputs(9883) <= b;
    layer0_outputs(9884) <= a or b;
    layer0_outputs(9885) <= not b;
    layer0_outputs(9886) <= not a or b;
    layer0_outputs(9887) <= 1'b1;
    layer0_outputs(9888) <= not (a xor b);
    layer0_outputs(9889) <= 1'b1;
    layer0_outputs(9890) <= a or b;
    layer0_outputs(9891) <= b;
    layer0_outputs(9892) <= not a;
    layer0_outputs(9893) <= a xor b;
    layer0_outputs(9894) <= a or b;
    layer0_outputs(9895) <= not b;
    layer0_outputs(9896) <= not (a or b);
    layer0_outputs(9897) <= b and not a;
    layer0_outputs(9898) <= not b;
    layer0_outputs(9899) <= not a or b;
    layer0_outputs(9900) <= a and b;
    layer0_outputs(9901) <= not b;
    layer0_outputs(9902) <= 1'b1;
    layer0_outputs(9903) <= a;
    layer0_outputs(9904) <= b and not a;
    layer0_outputs(9905) <= a or b;
    layer0_outputs(9906) <= a;
    layer0_outputs(9907) <= not a or b;
    layer0_outputs(9908) <= not b or a;
    layer0_outputs(9909) <= a;
    layer0_outputs(9910) <= a or b;
    layer0_outputs(9911) <= not (a or b);
    layer0_outputs(9912) <= not b or a;
    layer0_outputs(9913) <= not b or a;
    layer0_outputs(9914) <= not a;
    layer0_outputs(9915) <= a xor b;
    layer0_outputs(9916) <= not b or a;
    layer0_outputs(9917) <= 1'b1;
    layer0_outputs(9918) <= not (a or b);
    layer0_outputs(9919) <= a and b;
    layer0_outputs(9920) <= a or b;
    layer0_outputs(9921) <= not a;
    layer0_outputs(9922) <= a xor b;
    layer0_outputs(9923) <= a and b;
    layer0_outputs(9924) <= not a or b;
    layer0_outputs(9925) <= a and not b;
    layer0_outputs(9926) <= a xor b;
    layer0_outputs(9927) <= a or b;
    layer0_outputs(9928) <= a xor b;
    layer0_outputs(9929) <= not (a xor b);
    layer0_outputs(9930) <= a or b;
    layer0_outputs(9931) <= a and b;
    layer0_outputs(9932) <= not (a and b);
    layer0_outputs(9933) <= a and not b;
    layer0_outputs(9934) <= not (a xor b);
    layer0_outputs(9935) <= not b or a;
    layer0_outputs(9936) <= a xor b;
    layer0_outputs(9937) <= not a or b;
    layer0_outputs(9938) <= a xor b;
    layer0_outputs(9939) <= a xor b;
    layer0_outputs(9940) <= not (a or b);
    layer0_outputs(9941) <= not (a xor b);
    layer0_outputs(9942) <= not (a xor b);
    layer0_outputs(9943) <= a or b;
    layer0_outputs(9944) <= a xor b;
    layer0_outputs(9945) <= a and not b;
    layer0_outputs(9946) <= a xor b;
    layer0_outputs(9947) <= not a;
    layer0_outputs(9948) <= not (a or b);
    layer0_outputs(9949) <= a or b;
    layer0_outputs(9950) <= a or b;
    layer0_outputs(9951) <= a;
    layer0_outputs(9952) <= a;
    layer0_outputs(9953) <= a and not b;
    layer0_outputs(9954) <= not b;
    layer0_outputs(9955) <= not (a or b);
    layer0_outputs(9956) <= a or b;
    layer0_outputs(9957) <= a and b;
    layer0_outputs(9958) <= not a;
    layer0_outputs(9959) <= not b;
    layer0_outputs(9960) <= a and not b;
    layer0_outputs(9961) <= b and not a;
    layer0_outputs(9962) <= not a;
    layer0_outputs(9963) <= not (a or b);
    layer0_outputs(9964) <= not (a xor b);
    layer0_outputs(9965) <= not a;
    layer0_outputs(9966) <= a or b;
    layer0_outputs(9967) <= a and not b;
    layer0_outputs(9968) <= a and not b;
    layer0_outputs(9969) <= b;
    layer0_outputs(9970) <= b and not a;
    layer0_outputs(9971) <= not (a xor b);
    layer0_outputs(9972) <= not (a xor b);
    layer0_outputs(9973) <= not a;
    layer0_outputs(9974) <= not (a or b);
    layer0_outputs(9975) <= not b;
    layer0_outputs(9976) <= a and not b;
    layer0_outputs(9977) <= b and not a;
    layer0_outputs(9978) <= a and not b;
    layer0_outputs(9979) <= not b or a;
    layer0_outputs(9980) <= not b;
    layer0_outputs(9981) <= not a;
    layer0_outputs(9982) <= a or b;
    layer0_outputs(9983) <= not (a and b);
    layer0_outputs(9984) <= b and not a;
    layer0_outputs(9985) <= a and not b;
    layer0_outputs(9986) <= b;
    layer0_outputs(9987) <= not (a or b);
    layer0_outputs(9988) <= a or b;
    layer0_outputs(9989) <= a xor b;
    layer0_outputs(9990) <= not a;
    layer0_outputs(9991) <= not (a or b);
    layer0_outputs(9992) <= a xor b;
    layer0_outputs(9993) <= not a;
    layer0_outputs(9994) <= not (a or b);
    layer0_outputs(9995) <= not (a xor b);
    layer0_outputs(9996) <= not (a xor b);
    layer0_outputs(9997) <= b;
    layer0_outputs(9998) <= not b;
    layer0_outputs(9999) <= b and not a;
    layer0_outputs(10000) <= not (a or b);
    layer0_outputs(10001) <= a and not b;
    layer0_outputs(10002) <= a xor b;
    layer0_outputs(10003) <= b;
    layer0_outputs(10004) <= a and not b;
    layer0_outputs(10005) <= a;
    layer0_outputs(10006) <= not (a or b);
    layer0_outputs(10007) <= b;
    layer0_outputs(10008) <= not (a or b);
    layer0_outputs(10009) <= a or b;
    layer0_outputs(10010) <= not b;
    layer0_outputs(10011) <= not b;
    layer0_outputs(10012) <= not a or b;
    layer0_outputs(10013) <= b and not a;
    layer0_outputs(10014) <= not (a xor b);
    layer0_outputs(10015) <= not (a xor b);
    layer0_outputs(10016) <= a or b;
    layer0_outputs(10017) <= a xor b;
    layer0_outputs(10018) <= a;
    layer0_outputs(10019) <= not (a or b);
    layer0_outputs(10020) <= a or b;
    layer0_outputs(10021) <= not a or b;
    layer0_outputs(10022) <= a and not b;
    layer0_outputs(10023) <= not (a or b);
    layer0_outputs(10024) <= not (a xor b);
    layer0_outputs(10025) <= a or b;
    layer0_outputs(10026) <= not (a or b);
    layer0_outputs(10027) <= not a or b;
    layer0_outputs(10028) <= a xor b;
    layer0_outputs(10029) <= not a;
    layer0_outputs(10030) <= a xor b;
    layer0_outputs(10031) <= b and not a;
    layer0_outputs(10032) <= b and not a;
    layer0_outputs(10033) <= not (a or b);
    layer0_outputs(10034) <= not (a xor b);
    layer0_outputs(10035) <= not (a or b);
    layer0_outputs(10036) <= a;
    layer0_outputs(10037) <= not b or a;
    layer0_outputs(10038) <= not a or b;
    layer0_outputs(10039) <= not (a or b);
    layer0_outputs(10040) <= not a or b;
    layer0_outputs(10041) <= a xor b;
    layer0_outputs(10042) <= not b;
    layer0_outputs(10043) <= a or b;
    layer0_outputs(10044) <= a or b;
    layer0_outputs(10045) <= not (a or b);
    layer0_outputs(10046) <= b;
    layer0_outputs(10047) <= not b or a;
    layer0_outputs(10048) <= a or b;
    layer0_outputs(10049) <= not (a or b);
    layer0_outputs(10050) <= 1'b1;
    layer0_outputs(10051) <= not a;
    layer0_outputs(10052) <= a xor b;
    layer0_outputs(10053) <= not b or a;
    layer0_outputs(10054) <= not a or b;
    layer0_outputs(10055) <= not a;
    layer0_outputs(10056) <= not a or b;
    layer0_outputs(10057) <= a and not b;
    layer0_outputs(10058) <= not (a or b);
    layer0_outputs(10059) <= a or b;
    layer0_outputs(10060) <= not (a or b);
    layer0_outputs(10061) <= not a or b;
    layer0_outputs(10062) <= b;
    layer0_outputs(10063) <= a or b;
    layer0_outputs(10064) <= not a or b;
    layer0_outputs(10065) <= a;
    layer0_outputs(10066) <= b;
    layer0_outputs(10067) <= not (a or b);
    layer0_outputs(10068) <= a and not b;
    layer0_outputs(10069) <= a xor b;
    layer0_outputs(10070) <= not b;
    layer0_outputs(10071) <= not b;
    layer0_outputs(10072) <= not (a or b);
    layer0_outputs(10073) <= a xor b;
    layer0_outputs(10074) <= not (a xor b);
    layer0_outputs(10075) <= a and not b;
    layer0_outputs(10076) <= 1'b1;
    layer0_outputs(10077) <= not (a or b);
    layer0_outputs(10078) <= not a or b;
    layer0_outputs(10079) <= a and b;
    layer0_outputs(10080) <= not (a or b);
    layer0_outputs(10081) <= b and not a;
    layer0_outputs(10082) <= a xor b;
    layer0_outputs(10083) <= a or b;
    layer0_outputs(10084) <= a and b;
    layer0_outputs(10085) <= a and not b;
    layer0_outputs(10086) <= a;
    layer0_outputs(10087) <= not (a xor b);
    layer0_outputs(10088) <= not b or a;
    layer0_outputs(10089) <= a xor b;
    layer0_outputs(10090) <= a or b;
    layer0_outputs(10091) <= b and not a;
    layer0_outputs(10092) <= a;
    layer0_outputs(10093) <= a or b;
    layer0_outputs(10094) <= not b;
    layer0_outputs(10095) <= not a or b;
    layer0_outputs(10096) <= not (a and b);
    layer0_outputs(10097) <= not a or b;
    layer0_outputs(10098) <= not a;
    layer0_outputs(10099) <= not a or b;
    layer0_outputs(10100) <= 1'b0;
    layer0_outputs(10101) <= a xor b;
    layer0_outputs(10102) <= a;
    layer0_outputs(10103) <= not (a xor b);
    layer0_outputs(10104) <= a and not b;
    layer0_outputs(10105) <= not (a or b);
    layer0_outputs(10106) <= b and not a;
    layer0_outputs(10107) <= a;
    layer0_outputs(10108) <= not b;
    layer0_outputs(10109) <= not (a xor b);
    layer0_outputs(10110) <= a xor b;
    layer0_outputs(10111) <= b and not a;
    layer0_outputs(10112) <= not (a or b);
    layer0_outputs(10113) <= not a;
    layer0_outputs(10114) <= not b;
    layer0_outputs(10115) <= not (a and b);
    layer0_outputs(10116) <= not a;
    layer0_outputs(10117) <= b;
    layer0_outputs(10118) <= not (a or b);
    layer0_outputs(10119) <= not (a or b);
    layer0_outputs(10120) <= not a;
    layer0_outputs(10121) <= a;
    layer0_outputs(10122) <= a xor b;
    layer0_outputs(10123) <= 1'b0;
    layer0_outputs(10124) <= not b;
    layer0_outputs(10125) <= not a or b;
    layer0_outputs(10126) <= not (a xor b);
    layer0_outputs(10127) <= a xor b;
    layer0_outputs(10128) <= not (a xor b);
    layer0_outputs(10129) <= not (a or b);
    layer0_outputs(10130) <= a or b;
    layer0_outputs(10131) <= not (a or b);
    layer0_outputs(10132) <= a and b;
    layer0_outputs(10133) <= a or b;
    layer0_outputs(10134) <= a xor b;
    layer0_outputs(10135) <= 1'b0;
    layer0_outputs(10136) <= not (a xor b);
    layer0_outputs(10137) <= not b;
    layer0_outputs(10138) <= not b or a;
    layer0_outputs(10139) <= a;
    layer0_outputs(10140) <= not (a or b);
    layer0_outputs(10141) <= not b or a;
    layer0_outputs(10142) <= a;
    layer0_outputs(10143) <= not b;
    layer0_outputs(10144) <= 1'b1;
    layer0_outputs(10145) <= not b;
    layer0_outputs(10146) <= a xor b;
    layer0_outputs(10147) <= a xor b;
    layer0_outputs(10148) <= not (a or b);
    layer0_outputs(10149) <= a;
    layer0_outputs(10150) <= not (a or b);
    layer0_outputs(10151) <= not a;
    layer0_outputs(10152) <= not b or a;
    layer0_outputs(10153) <= not (a xor b);
    layer0_outputs(10154) <= not (a or b);
    layer0_outputs(10155) <= a or b;
    layer0_outputs(10156) <= a or b;
    layer0_outputs(10157) <= not (a xor b);
    layer0_outputs(10158) <= a or b;
    layer0_outputs(10159) <= a xor b;
    layer0_outputs(10160) <= not b or a;
    layer0_outputs(10161) <= b;
    layer0_outputs(10162) <= not (a and b);
    layer0_outputs(10163) <= not a or b;
    layer0_outputs(10164) <= a xor b;
    layer0_outputs(10165) <= not (a or b);
    layer0_outputs(10166) <= not (a xor b);
    layer0_outputs(10167) <= a and not b;
    layer0_outputs(10168) <= not (a xor b);
    layer0_outputs(10169) <= not (a or b);
    layer0_outputs(10170) <= a or b;
    layer0_outputs(10171) <= not (a xor b);
    layer0_outputs(10172) <= a xor b;
    layer0_outputs(10173) <= not (a xor b);
    layer0_outputs(10174) <= a or b;
    layer0_outputs(10175) <= not (a or b);
    layer0_outputs(10176) <= not (a or b);
    layer0_outputs(10177) <= b and not a;
    layer0_outputs(10178) <= not (a or b);
    layer0_outputs(10179) <= not (a and b);
    layer0_outputs(10180) <= not (a or b);
    layer0_outputs(10181) <= 1'b0;
    layer0_outputs(10182) <= not b;
    layer0_outputs(10183) <= a;
    layer0_outputs(10184) <= b and not a;
    layer0_outputs(10185) <= not (a xor b);
    layer0_outputs(10186) <= not a or b;
    layer0_outputs(10187) <= b;
    layer0_outputs(10188) <= a and not b;
    layer0_outputs(10189) <= a and b;
    layer0_outputs(10190) <= not a or b;
    layer0_outputs(10191) <= not a;
    layer0_outputs(10192) <= not a;
    layer0_outputs(10193) <= a xor b;
    layer0_outputs(10194) <= a xor b;
    layer0_outputs(10195) <= not b or a;
    layer0_outputs(10196) <= a and b;
    layer0_outputs(10197) <= not a or b;
    layer0_outputs(10198) <= not a;
    layer0_outputs(10199) <= not b;
    layer0_outputs(10200) <= not (a and b);
    layer0_outputs(10201) <= a or b;
    layer0_outputs(10202) <= b;
    layer0_outputs(10203) <= a;
    layer0_outputs(10204) <= not (a or b);
    layer0_outputs(10205) <= b;
    layer0_outputs(10206) <= not (a or b);
    layer0_outputs(10207) <= not (a or b);
    layer0_outputs(10208) <= b;
    layer0_outputs(10209) <= not a;
    layer0_outputs(10210) <= not (a or b);
    layer0_outputs(10211) <= not a;
    layer0_outputs(10212) <= a or b;
    layer0_outputs(10213) <= not b or a;
    layer0_outputs(10214) <= not a;
    layer0_outputs(10215) <= b and not a;
    layer0_outputs(10216) <= a;
    layer0_outputs(10217) <= not b;
    layer0_outputs(10218) <= b and not a;
    layer0_outputs(10219) <= a or b;
    layer0_outputs(10220) <= a or b;
    layer0_outputs(10221) <= not (a and b);
    layer0_outputs(10222) <= a or b;
    layer0_outputs(10223) <= not (a xor b);
    layer0_outputs(10224) <= b;
    layer0_outputs(10225) <= a and not b;
    layer0_outputs(10226) <= a xor b;
    layer0_outputs(10227) <= not (a or b);
    layer0_outputs(10228) <= not a or b;
    layer0_outputs(10229) <= not (a and b);
    layer0_outputs(10230) <= not (a xor b);
    layer0_outputs(10231) <= a xor b;
    layer0_outputs(10232) <= a;
    layer0_outputs(10233) <= a xor b;
    layer0_outputs(10234) <= a xor b;
    layer0_outputs(10235) <= a or b;
    layer0_outputs(10236) <= b and not a;
    layer0_outputs(10237) <= not a;
    layer0_outputs(10238) <= b;
    layer0_outputs(10239) <= a;
    layer0_outputs(10240) <= a xor b;
    layer0_outputs(10241) <= not (a or b);
    layer0_outputs(10242) <= 1'b0;
    layer0_outputs(10243) <= a xor b;
    layer0_outputs(10244) <= not (a or b);
    layer0_outputs(10245) <= not (a xor b);
    layer0_outputs(10246) <= not (a or b);
    layer0_outputs(10247) <= b and not a;
    layer0_outputs(10248) <= not (a or b);
    layer0_outputs(10249) <= not a or b;
    layer0_outputs(10250) <= a xor b;
    layer0_outputs(10251) <= not (a xor b);
    layer0_outputs(10252) <= not (a or b);
    layer0_outputs(10253) <= not b;
    layer0_outputs(10254) <= a;
    layer0_outputs(10255) <= not (a xor b);
    layer0_outputs(10256) <= not (a or b);
    layer0_outputs(10257) <= not b or a;
    layer0_outputs(10258) <= not (a or b);
    layer0_outputs(10259) <= a;
    layer0_outputs(10260) <= a;
    layer0_outputs(10261) <= not (a xor b);
    layer0_outputs(10262) <= a or b;
    layer0_outputs(10263) <= not a or b;
    layer0_outputs(10264) <= a and not b;
    layer0_outputs(10265) <= not (a xor b);
    layer0_outputs(10266) <= 1'b0;
    layer0_outputs(10267) <= not (a or b);
    layer0_outputs(10268) <= a and not b;
    layer0_outputs(10269) <= not (a or b);
    layer0_outputs(10270) <= a or b;
    layer0_outputs(10271) <= not (a or b);
    layer0_outputs(10272) <= a and not b;
    layer0_outputs(10273) <= b and not a;
    layer0_outputs(10274) <= b and not a;
    layer0_outputs(10275) <= a and not b;
    layer0_outputs(10276) <= not (a and b);
    layer0_outputs(10277) <= not b or a;
    layer0_outputs(10278) <= not a or b;
    layer0_outputs(10279) <= a xor b;
    layer0_outputs(10280) <= b;
    layer0_outputs(10281) <= b;
    layer0_outputs(10282) <= a;
    layer0_outputs(10283) <= b;
    layer0_outputs(10284) <= a xor b;
    layer0_outputs(10285) <= not (a xor b);
    layer0_outputs(10286) <= a;
    layer0_outputs(10287) <= a xor b;
    layer0_outputs(10288) <= not (a or b);
    layer0_outputs(10289) <= not (a and b);
    layer0_outputs(10290) <= a and not b;
    layer0_outputs(10291) <= a xor b;
    layer0_outputs(10292) <= 1'b1;
    layer0_outputs(10293) <= not a;
    layer0_outputs(10294) <= not a or b;
    layer0_outputs(10295) <= a or b;
    layer0_outputs(10296) <= not b;
    layer0_outputs(10297) <= a and not b;
    layer0_outputs(10298) <= not (a xor b);
    layer0_outputs(10299) <= a;
    layer0_outputs(10300) <= a;
    layer0_outputs(10301) <= not a;
    layer0_outputs(10302) <= not b or a;
    layer0_outputs(10303) <= not (a or b);
    layer0_outputs(10304) <= not (a or b);
    layer0_outputs(10305) <= not (a and b);
    layer0_outputs(10306) <= not b;
    layer0_outputs(10307) <= a;
    layer0_outputs(10308) <= a;
    layer0_outputs(10309) <= a or b;
    layer0_outputs(10310) <= not (a and b);
    layer0_outputs(10311) <= 1'b1;
    layer0_outputs(10312) <= not (a xor b);
    layer0_outputs(10313) <= a or b;
    layer0_outputs(10314) <= a xor b;
    layer0_outputs(10315) <= a;
    layer0_outputs(10316) <= a or b;
    layer0_outputs(10317) <= not a;
    layer0_outputs(10318) <= not (a or b);
    layer0_outputs(10319) <= not (a or b);
    layer0_outputs(10320) <= a;
    layer0_outputs(10321) <= 1'b1;
    layer0_outputs(10322) <= a or b;
    layer0_outputs(10323) <= not a;
    layer0_outputs(10324) <= not a;
    layer0_outputs(10325) <= a or b;
    layer0_outputs(10326) <= not (a xor b);
    layer0_outputs(10327) <= not a or b;
    layer0_outputs(10328) <= not b or a;
    layer0_outputs(10329) <= not a or b;
    layer0_outputs(10330) <= a or b;
    layer0_outputs(10331) <= a;
    layer0_outputs(10332) <= 1'b0;
    layer0_outputs(10333) <= a;
    layer0_outputs(10334) <= not b;
    layer0_outputs(10335) <= not (a and b);
    layer0_outputs(10336) <= b and not a;
    layer0_outputs(10337) <= not (a xor b);
    layer0_outputs(10338) <= b;
    layer0_outputs(10339) <= a xor b;
    layer0_outputs(10340) <= a or b;
    layer0_outputs(10341) <= a and not b;
    layer0_outputs(10342) <= a;
    layer0_outputs(10343) <= a and not b;
    layer0_outputs(10344) <= not (a or b);
    layer0_outputs(10345) <= 1'b0;
    layer0_outputs(10346) <= a;
    layer0_outputs(10347) <= a or b;
    layer0_outputs(10348) <= not a;
    layer0_outputs(10349) <= a;
    layer0_outputs(10350) <= not a;
    layer0_outputs(10351) <= not (a or b);
    layer0_outputs(10352) <= not a or b;
    layer0_outputs(10353) <= a or b;
    layer0_outputs(10354) <= not b;
    layer0_outputs(10355) <= not (a xor b);
    layer0_outputs(10356) <= a xor b;
    layer0_outputs(10357) <= a or b;
    layer0_outputs(10358) <= not b;
    layer0_outputs(10359) <= not (a or b);
    layer0_outputs(10360) <= not (a xor b);
    layer0_outputs(10361) <= not a;
    layer0_outputs(10362) <= not (a xor b);
    layer0_outputs(10363) <= not (a xor b);
    layer0_outputs(10364) <= b;
    layer0_outputs(10365) <= not b or a;
    layer0_outputs(10366) <= not (a or b);
    layer0_outputs(10367) <= a xor b;
    layer0_outputs(10368) <= not a or b;
    layer0_outputs(10369) <= a or b;
    layer0_outputs(10370) <= a or b;
    layer0_outputs(10371) <= a or b;
    layer0_outputs(10372) <= not b;
    layer0_outputs(10373) <= not (a or b);
    layer0_outputs(10374) <= not (a or b);
    layer0_outputs(10375) <= not a or b;
    layer0_outputs(10376) <= a;
    layer0_outputs(10377) <= not (a xor b);
    layer0_outputs(10378) <= not (a xor b);
    layer0_outputs(10379) <= a or b;
    layer0_outputs(10380) <= a or b;
    layer0_outputs(10381) <= b and not a;
    layer0_outputs(10382) <= not (a xor b);
    layer0_outputs(10383) <= b and not a;
    layer0_outputs(10384) <= not b;
    layer0_outputs(10385) <= not b or a;
    layer0_outputs(10386) <= not a;
    layer0_outputs(10387) <= a or b;
    layer0_outputs(10388) <= not b or a;
    layer0_outputs(10389) <= a xor b;
    layer0_outputs(10390) <= a or b;
    layer0_outputs(10391) <= not b or a;
    layer0_outputs(10392) <= 1'b0;
    layer0_outputs(10393) <= a or b;
    layer0_outputs(10394) <= a or b;
    layer0_outputs(10395) <= a xor b;
    layer0_outputs(10396) <= a xor b;
    layer0_outputs(10397) <= not b or a;
    layer0_outputs(10398) <= not (a or b);
    layer0_outputs(10399) <= a and not b;
    layer0_outputs(10400) <= 1'b0;
    layer0_outputs(10401) <= not (a xor b);
    layer0_outputs(10402) <= b and not a;
    layer0_outputs(10403) <= b and not a;
    layer0_outputs(10404) <= not a or b;
    layer0_outputs(10405) <= a xor b;
    layer0_outputs(10406) <= a and not b;
    layer0_outputs(10407) <= b;
    layer0_outputs(10408) <= not (a and b);
    layer0_outputs(10409) <= a;
    layer0_outputs(10410) <= a;
    layer0_outputs(10411) <= a or b;
    layer0_outputs(10412) <= not b;
    layer0_outputs(10413) <= a or b;
    layer0_outputs(10414) <= not (a or b);
    layer0_outputs(10415) <= a and not b;
    layer0_outputs(10416) <= not b;
    layer0_outputs(10417) <= a and b;
    layer0_outputs(10418) <= not b;
    layer0_outputs(10419) <= b;
    layer0_outputs(10420) <= a and b;
    layer0_outputs(10421) <= a or b;
    layer0_outputs(10422) <= not (a or b);
    layer0_outputs(10423) <= a and b;
    layer0_outputs(10424) <= not (a xor b);
    layer0_outputs(10425) <= not (a xor b);
    layer0_outputs(10426) <= 1'b1;
    layer0_outputs(10427) <= a or b;
    layer0_outputs(10428) <= a;
    layer0_outputs(10429) <= not (a or b);
    layer0_outputs(10430) <= a and b;
    layer0_outputs(10431) <= not a or b;
    layer0_outputs(10432) <= not a;
    layer0_outputs(10433) <= a xor b;
    layer0_outputs(10434) <= not a or b;
    layer0_outputs(10435) <= a or b;
    layer0_outputs(10436) <= b;
    layer0_outputs(10437) <= not b;
    layer0_outputs(10438) <= b and not a;
    layer0_outputs(10439) <= not a or b;
    layer0_outputs(10440) <= b and not a;
    layer0_outputs(10441) <= not a;
    layer0_outputs(10442) <= not b;
    layer0_outputs(10443) <= a xor b;
    layer0_outputs(10444) <= not (a xor b);
    layer0_outputs(10445) <= not (a xor b);
    layer0_outputs(10446) <= a xor b;
    layer0_outputs(10447) <= b;
    layer0_outputs(10448) <= b;
    layer0_outputs(10449) <= not a or b;
    layer0_outputs(10450) <= a or b;
    layer0_outputs(10451) <= not b or a;
    layer0_outputs(10452) <= a or b;
    layer0_outputs(10453) <= b;
    layer0_outputs(10454) <= not a or b;
    layer0_outputs(10455) <= not b or a;
    layer0_outputs(10456) <= not (a or b);
    layer0_outputs(10457) <= a and not b;
    layer0_outputs(10458) <= a or b;
    layer0_outputs(10459) <= a and not b;
    layer0_outputs(10460) <= b;
    layer0_outputs(10461) <= a or b;
    layer0_outputs(10462) <= b;
    layer0_outputs(10463) <= not a or b;
    layer0_outputs(10464) <= 1'b0;
    layer0_outputs(10465) <= not a or b;
    layer0_outputs(10466) <= not a;
    layer0_outputs(10467) <= a xor b;
    layer0_outputs(10468) <= a or b;
    layer0_outputs(10469) <= not (a or b);
    layer0_outputs(10470) <= 1'b1;
    layer0_outputs(10471) <= b and not a;
    layer0_outputs(10472) <= not b or a;
    layer0_outputs(10473) <= a and b;
    layer0_outputs(10474) <= not (a or b);
    layer0_outputs(10475) <= a;
    layer0_outputs(10476) <= not a or b;
    layer0_outputs(10477) <= not b;
    layer0_outputs(10478) <= not (a xor b);
    layer0_outputs(10479) <= not (a or b);
    layer0_outputs(10480) <= not a;
    layer0_outputs(10481) <= 1'b0;
    layer0_outputs(10482) <= a or b;
    layer0_outputs(10483) <= not a;
    layer0_outputs(10484) <= not a;
    layer0_outputs(10485) <= not (a xor b);
    layer0_outputs(10486) <= 1'b0;
    layer0_outputs(10487) <= a or b;
    layer0_outputs(10488) <= not b or a;
    layer0_outputs(10489) <= not b;
    layer0_outputs(10490) <= a xor b;
    layer0_outputs(10491) <= b;
    layer0_outputs(10492) <= a or b;
    layer0_outputs(10493) <= a xor b;
    layer0_outputs(10494) <= b;
    layer0_outputs(10495) <= a or b;
    layer0_outputs(10496) <= a or b;
    layer0_outputs(10497) <= not (a or b);
    layer0_outputs(10498) <= a;
    layer0_outputs(10499) <= b;
    layer0_outputs(10500) <= 1'b0;
    layer0_outputs(10501) <= not b or a;
    layer0_outputs(10502) <= not b or a;
    layer0_outputs(10503) <= not (a xor b);
    layer0_outputs(10504) <= not (a xor b);
    layer0_outputs(10505) <= b and not a;
    layer0_outputs(10506) <= b;
    layer0_outputs(10507) <= not a or b;
    layer0_outputs(10508) <= b;
    layer0_outputs(10509) <= not (a xor b);
    layer0_outputs(10510) <= not (a xor b);
    layer0_outputs(10511) <= not b;
    layer0_outputs(10512) <= not (a or b);
    layer0_outputs(10513) <= a or b;
    layer0_outputs(10514) <= a xor b;
    layer0_outputs(10515) <= a or b;
    layer0_outputs(10516) <= not b or a;
    layer0_outputs(10517) <= a xor b;
    layer0_outputs(10518) <= a or b;
    layer0_outputs(10519) <= b;
    layer0_outputs(10520) <= b;
    layer0_outputs(10521) <= not (a xor b);
    layer0_outputs(10522) <= 1'b1;
    layer0_outputs(10523) <= not a;
    layer0_outputs(10524) <= b and not a;
    layer0_outputs(10525) <= a or b;
    layer0_outputs(10526) <= not (a or b);
    layer0_outputs(10527) <= not a;
    layer0_outputs(10528) <= not (a xor b);
    layer0_outputs(10529) <= a and not b;
    layer0_outputs(10530) <= not a or b;
    layer0_outputs(10531) <= b;
    layer0_outputs(10532) <= a xor b;
    layer0_outputs(10533) <= not (a or b);
    layer0_outputs(10534) <= b;
    layer0_outputs(10535) <= b;
    layer0_outputs(10536) <= not (a xor b);
    layer0_outputs(10537) <= a;
    layer0_outputs(10538) <= 1'b1;
    layer0_outputs(10539) <= not (a or b);
    layer0_outputs(10540) <= a and b;
    layer0_outputs(10541) <= not (a xor b);
    layer0_outputs(10542) <= not b;
    layer0_outputs(10543) <= not (a xor b);
    layer0_outputs(10544) <= not b;
    layer0_outputs(10545) <= not (a or b);
    layer0_outputs(10546) <= 1'b0;
    layer0_outputs(10547) <= not b or a;
    layer0_outputs(10548) <= not (a and b);
    layer0_outputs(10549) <= a or b;
    layer0_outputs(10550) <= not b or a;
    layer0_outputs(10551) <= a or b;
    layer0_outputs(10552) <= a and b;
    layer0_outputs(10553) <= a or b;
    layer0_outputs(10554) <= not (a xor b);
    layer0_outputs(10555) <= a xor b;
    layer0_outputs(10556) <= a xor b;
    layer0_outputs(10557) <= b;
    layer0_outputs(10558) <= b and not a;
    layer0_outputs(10559) <= not a or b;
    layer0_outputs(10560) <= a and b;
    layer0_outputs(10561) <= not b or a;
    layer0_outputs(10562) <= b and not a;
    layer0_outputs(10563) <= a;
    layer0_outputs(10564) <= not b;
    layer0_outputs(10565) <= b and not a;
    layer0_outputs(10566) <= not a or b;
    layer0_outputs(10567) <= a xor b;
    layer0_outputs(10568) <= not b;
    layer0_outputs(10569) <= b;
    layer0_outputs(10570) <= b and not a;
    layer0_outputs(10571) <= not a or b;
    layer0_outputs(10572) <= not (a xor b);
    layer0_outputs(10573) <= not b or a;
    layer0_outputs(10574) <= not b or a;
    layer0_outputs(10575) <= not b or a;
    layer0_outputs(10576) <= b;
    layer0_outputs(10577) <= 1'b1;
    layer0_outputs(10578) <= not (a and b);
    layer0_outputs(10579) <= a or b;
    layer0_outputs(10580) <= a;
    layer0_outputs(10581) <= a xor b;
    layer0_outputs(10582) <= not (a or b);
    layer0_outputs(10583) <= not a or b;
    layer0_outputs(10584) <= not (a or b);
    layer0_outputs(10585) <= not b;
    layer0_outputs(10586) <= not (a xor b);
    layer0_outputs(10587) <= not a or b;
    layer0_outputs(10588) <= not (a or b);
    layer0_outputs(10589) <= a or b;
    layer0_outputs(10590) <= not (a xor b);
    layer0_outputs(10591) <= not b;
    layer0_outputs(10592) <= a and not b;
    layer0_outputs(10593) <= a and b;
    layer0_outputs(10594) <= not (a or b);
    layer0_outputs(10595) <= a;
    layer0_outputs(10596) <= not (a or b);
    layer0_outputs(10597) <= not (a xor b);
    layer0_outputs(10598) <= not b or a;
    layer0_outputs(10599) <= not (a or b);
    layer0_outputs(10600) <= 1'b0;
    layer0_outputs(10601) <= a or b;
    layer0_outputs(10602) <= not (a or b);
    layer0_outputs(10603) <= b;
    layer0_outputs(10604) <= a xor b;
    layer0_outputs(10605) <= not (a and b);
    layer0_outputs(10606) <= a;
    layer0_outputs(10607) <= not (a and b);
    layer0_outputs(10608) <= not b;
    layer0_outputs(10609) <= b and not a;
    layer0_outputs(10610) <= 1'b0;
    layer0_outputs(10611) <= a;
    layer0_outputs(10612) <= not (a xor b);
    layer0_outputs(10613) <= b;
    layer0_outputs(10614) <= not b;
    layer0_outputs(10615) <= not (a or b);
    layer0_outputs(10616) <= a xor b;
    layer0_outputs(10617) <= not b;
    layer0_outputs(10618) <= a and not b;
    layer0_outputs(10619) <= a or b;
    layer0_outputs(10620) <= not a or b;
    layer0_outputs(10621) <= b;
    layer0_outputs(10622) <= 1'b0;
    layer0_outputs(10623) <= not b;
    layer0_outputs(10624) <= a xor b;
    layer0_outputs(10625) <= a;
    layer0_outputs(10626) <= not (a and b);
    layer0_outputs(10627) <= not b or a;
    layer0_outputs(10628) <= a xor b;
    layer0_outputs(10629) <= a;
    layer0_outputs(10630) <= b;
    layer0_outputs(10631) <= not (a or b);
    layer0_outputs(10632) <= a or b;
    layer0_outputs(10633) <= not a or b;
    layer0_outputs(10634) <= not b or a;
    layer0_outputs(10635) <= not a or b;
    layer0_outputs(10636) <= not (a or b);
    layer0_outputs(10637) <= not (a or b);
    layer0_outputs(10638) <= b;
    layer0_outputs(10639) <= not a;
    layer0_outputs(10640) <= a and b;
    layer0_outputs(10641) <= not (a xor b);
    layer0_outputs(10642) <= 1'b1;
    layer0_outputs(10643) <= not b or a;
    layer0_outputs(10644) <= b and not a;
    layer0_outputs(10645) <= not a;
    layer0_outputs(10646) <= not a or b;
    layer0_outputs(10647) <= a xor b;
    layer0_outputs(10648) <= b;
    layer0_outputs(10649) <= not (a xor b);
    layer0_outputs(10650) <= a xor b;
    layer0_outputs(10651) <= not b or a;
    layer0_outputs(10652) <= a and not b;
    layer0_outputs(10653) <= not (a and b);
    layer0_outputs(10654) <= not (a or b);
    layer0_outputs(10655) <= not (a or b);
    layer0_outputs(10656) <= not b;
    layer0_outputs(10657) <= not a or b;
    layer0_outputs(10658) <= b;
    layer0_outputs(10659) <= b and not a;
    layer0_outputs(10660) <= a and not b;
    layer0_outputs(10661) <= 1'b1;
    layer0_outputs(10662) <= not (a or b);
    layer0_outputs(10663) <= not b;
    layer0_outputs(10664) <= not b;
    layer0_outputs(10665) <= b;
    layer0_outputs(10666) <= 1'b0;
    layer0_outputs(10667) <= not (a or b);
    layer0_outputs(10668) <= not a;
    layer0_outputs(10669) <= not (a xor b);
    layer0_outputs(10670) <= not (a and b);
    layer0_outputs(10671) <= a and b;
    layer0_outputs(10672) <= b;
    layer0_outputs(10673) <= a or b;
    layer0_outputs(10674) <= not a;
    layer0_outputs(10675) <= not b;
    layer0_outputs(10676) <= not a;
    layer0_outputs(10677) <= not b or a;
    layer0_outputs(10678) <= a;
    layer0_outputs(10679) <= not (a xor b);
    layer0_outputs(10680) <= not (a xor b);
    layer0_outputs(10681) <= not (a or b);
    layer0_outputs(10682) <= not (a xor b);
    layer0_outputs(10683) <= a;
    layer0_outputs(10684) <= b;
    layer0_outputs(10685) <= a;
    layer0_outputs(10686) <= a or b;
    layer0_outputs(10687) <= not b;
    layer0_outputs(10688) <= a and not b;
    layer0_outputs(10689) <= not b;
    layer0_outputs(10690) <= a or b;
    layer0_outputs(10691) <= a and not b;
    layer0_outputs(10692) <= a or b;
    layer0_outputs(10693) <= a and not b;
    layer0_outputs(10694) <= a or b;
    layer0_outputs(10695) <= a xor b;
    layer0_outputs(10696) <= not a;
    layer0_outputs(10697) <= not b;
    layer0_outputs(10698) <= not (a or b);
    layer0_outputs(10699) <= b and not a;
    layer0_outputs(10700) <= a xor b;
    layer0_outputs(10701) <= not b or a;
    layer0_outputs(10702) <= not (a xor b);
    layer0_outputs(10703) <= not a or b;
    layer0_outputs(10704) <= not b;
    layer0_outputs(10705) <= 1'b1;
    layer0_outputs(10706) <= not (a or b);
    layer0_outputs(10707) <= not (a or b);
    layer0_outputs(10708) <= b;
    layer0_outputs(10709) <= a xor b;
    layer0_outputs(10710) <= not (a or b);
    layer0_outputs(10711) <= not (a xor b);
    layer0_outputs(10712) <= 1'b0;
    layer0_outputs(10713) <= a;
    layer0_outputs(10714) <= not a or b;
    layer0_outputs(10715) <= not (a xor b);
    layer0_outputs(10716) <= a or b;
    layer0_outputs(10717) <= not (a and b);
    layer0_outputs(10718) <= a or b;
    layer0_outputs(10719) <= not b or a;
    layer0_outputs(10720) <= not b;
    layer0_outputs(10721) <= a xor b;
    layer0_outputs(10722) <= a;
    layer0_outputs(10723) <= a xor b;
    layer0_outputs(10724) <= not (a and b);
    layer0_outputs(10725) <= b and not a;
    layer0_outputs(10726) <= not b;
    layer0_outputs(10727) <= not b;
    layer0_outputs(10728) <= not (a or b);
    layer0_outputs(10729) <= not (a or b);
    layer0_outputs(10730) <= b;
    layer0_outputs(10731) <= not (a xor b);
    layer0_outputs(10732) <= not (a or b);
    layer0_outputs(10733) <= a;
    layer0_outputs(10734) <= not b or a;
    layer0_outputs(10735) <= a or b;
    layer0_outputs(10736) <= not (a or b);
    layer0_outputs(10737) <= not (a xor b);
    layer0_outputs(10738) <= not a or b;
    layer0_outputs(10739) <= not a or b;
    layer0_outputs(10740) <= not (a or b);
    layer0_outputs(10741) <= not a or b;
    layer0_outputs(10742) <= not (a xor b);
    layer0_outputs(10743) <= a and not b;
    layer0_outputs(10744) <= not b;
    layer0_outputs(10745) <= not (a xor b);
    layer0_outputs(10746) <= b;
    layer0_outputs(10747) <= b and not a;
    layer0_outputs(10748) <= not (a xor b);
    layer0_outputs(10749) <= a or b;
    layer0_outputs(10750) <= 1'b1;
    layer0_outputs(10751) <= not (a or b);
    layer0_outputs(10752) <= not b;
    layer0_outputs(10753) <= 1'b0;
    layer0_outputs(10754) <= a;
    layer0_outputs(10755) <= a xor b;
    layer0_outputs(10756) <= not (a and b);
    layer0_outputs(10757) <= a and not b;
    layer0_outputs(10758) <= a;
    layer0_outputs(10759) <= not (a xor b);
    layer0_outputs(10760) <= a and not b;
    layer0_outputs(10761) <= b;
    layer0_outputs(10762) <= not b or a;
    layer0_outputs(10763) <= not b or a;
    layer0_outputs(10764) <= not b;
    layer0_outputs(10765) <= not b;
    layer0_outputs(10766) <= a or b;
    layer0_outputs(10767) <= not (a or b);
    layer0_outputs(10768) <= b;
    layer0_outputs(10769) <= not b;
    layer0_outputs(10770) <= not b;
    layer0_outputs(10771) <= b and not a;
    layer0_outputs(10772) <= a;
    layer0_outputs(10773) <= not (a or b);
    layer0_outputs(10774) <= a;
    layer0_outputs(10775) <= not b;
    layer0_outputs(10776) <= a or b;
    layer0_outputs(10777) <= not a;
    layer0_outputs(10778) <= a xor b;
    layer0_outputs(10779) <= a xor b;
    layer0_outputs(10780) <= not a or b;
    layer0_outputs(10781) <= a or b;
    layer0_outputs(10782) <= b;
    layer0_outputs(10783) <= not b or a;
    layer0_outputs(10784) <= a and not b;
    layer0_outputs(10785) <= b;
    layer0_outputs(10786) <= b and not a;
    layer0_outputs(10787) <= a or b;
    layer0_outputs(10788) <= b and not a;
    layer0_outputs(10789) <= b and not a;
    layer0_outputs(10790) <= a xor b;
    layer0_outputs(10791) <= not b or a;
    layer0_outputs(10792) <= not (a or b);
    layer0_outputs(10793) <= a and b;
    layer0_outputs(10794) <= not b;
    layer0_outputs(10795) <= not b;
    layer0_outputs(10796) <= a;
    layer0_outputs(10797) <= a or b;
    layer0_outputs(10798) <= not a;
    layer0_outputs(10799) <= not b;
    layer0_outputs(10800) <= not (a and b);
    layer0_outputs(10801) <= b and not a;
    layer0_outputs(10802) <= not (a and b);
    layer0_outputs(10803) <= a or b;
    layer0_outputs(10804) <= a and not b;
    layer0_outputs(10805) <= not (a xor b);
    layer0_outputs(10806) <= not a;
    layer0_outputs(10807) <= 1'b1;
    layer0_outputs(10808) <= not (a xor b);
    layer0_outputs(10809) <= not a or b;
    layer0_outputs(10810) <= not b;
    layer0_outputs(10811) <= not b or a;
    layer0_outputs(10812) <= not b or a;
    layer0_outputs(10813) <= not b;
    layer0_outputs(10814) <= a;
    layer0_outputs(10815) <= not (a xor b);
    layer0_outputs(10816) <= a or b;
    layer0_outputs(10817) <= a and b;
    layer0_outputs(10818) <= a or b;
    layer0_outputs(10819) <= not a or b;
    layer0_outputs(10820) <= 1'b1;
    layer0_outputs(10821) <= a;
    layer0_outputs(10822) <= not a;
    layer0_outputs(10823) <= not (a or b);
    layer0_outputs(10824) <= a or b;
    layer0_outputs(10825) <= not a or b;
    layer0_outputs(10826) <= a or b;
    layer0_outputs(10827) <= not b;
    layer0_outputs(10828) <= b and not a;
    layer0_outputs(10829) <= not b;
    layer0_outputs(10830) <= a xor b;
    layer0_outputs(10831) <= a;
    layer0_outputs(10832) <= not (a xor b);
    layer0_outputs(10833) <= not b;
    layer0_outputs(10834) <= a or b;
    layer0_outputs(10835) <= a and not b;
    layer0_outputs(10836) <= a or b;
    layer0_outputs(10837) <= not b;
    layer0_outputs(10838) <= a or b;
    layer0_outputs(10839) <= a and not b;
    layer0_outputs(10840) <= not (a or b);
    layer0_outputs(10841) <= a or b;
    layer0_outputs(10842) <= a and b;
    layer0_outputs(10843) <= b;
    layer0_outputs(10844) <= not (a or b);
    layer0_outputs(10845) <= not (a xor b);
    layer0_outputs(10846) <= a xor b;
    layer0_outputs(10847) <= a or b;
    layer0_outputs(10848) <= not (a or b);
    layer0_outputs(10849) <= a and not b;
    layer0_outputs(10850) <= a xor b;
    layer0_outputs(10851) <= a;
    layer0_outputs(10852) <= not b or a;
    layer0_outputs(10853) <= a or b;
    layer0_outputs(10854) <= not b;
    layer0_outputs(10855) <= not b or a;
    layer0_outputs(10856) <= a xor b;
    layer0_outputs(10857) <= a and not b;
    layer0_outputs(10858) <= not b or a;
    layer0_outputs(10859) <= b and not a;
    layer0_outputs(10860) <= b;
    layer0_outputs(10861) <= a and not b;
    layer0_outputs(10862) <= not (a xor b);
    layer0_outputs(10863) <= a xor b;
    layer0_outputs(10864) <= not a or b;
    layer0_outputs(10865) <= not b;
    layer0_outputs(10866) <= not (a or b);
    layer0_outputs(10867) <= a or b;
    layer0_outputs(10868) <= not b or a;
    layer0_outputs(10869) <= not (a xor b);
    layer0_outputs(10870) <= not b or a;
    layer0_outputs(10871) <= not (a or b);
    layer0_outputs(10872) <= not (a xor b);
    layer0_outputs(10873) <= not (a or b);
    layer0_outputs(10874) <= not b;
    layer0_outputs(10875) <= not b or a;
    layer0_outputs(10876) <= a;
    layer0_outputs(10877) <= not (a or b);
    layer0_outputs(10878) <= not b;
    layer0_outputs(10879) <= a and b;
    layer0_outputs(10880) <= a;
    layer0_outputs(10881) <= a or b;
    layer0_outputs(10882) <= not (a and b);
    layer0_outputs(10883) <= not (a xor b);
    layer0_outputs(10884) <= 1'b1;
    layer0_outputs(10885) <= 1'b1;
    layer0_outputs(10886) <= not (a or b);
    layer0_outputs(10887) <= a xor b;
    layer0_outputs(10888) <= not b or a;
    layer0_outputs(10889) <= a or b;
    layer0_outputs(10890) <= a or b;
    layer0_outputs(10891) <= not (a or b);
    layer0_outputs(10892) <= not (a xor b);
    layer0_outputs(10893) <= not a or b;
    layer0_outputs(10894) <= not a;
    layer0_outputs(10895) <= a and not b;
    layer0_outputs(10896) <= 1'b0;
    layer0_outputs(10897) <= not (a or b);
    layer0_outputs(10898) <= a or b;
    layer0_outputs(10899) <= a or b;
    layer0_outputs(10900) <= b;
    layer0_outputs(10901) <= not b;
    layer0_outputs(10902) <= not (a xor b);
    layer0_outputs(10903) <= not a or b;
    layer0_outputs(10904) <= not b;
    layer0_outputs(10905) <= a xor b;
    layer0_outputs(10906) <= not a or b;
    layer0_outputs(10907) <= not b or a;
    layer0_outputs(10908) <= not a;
    layer0_outputs(10909) <= a or b;
    layer0_outputs(10910) <= not a or b;
    layer0_outputs(10911) <= not a or b;
    layer0_outputs(10912) <= a or b;
    layer0_outputs(10913) <= not (a xor b);
    layer0_outputs(10914) <= not a;
    layer0_outputs(10915) <= b;
    layer0_outputs(10916) <= a or b;
    layer0_outputs(10917) <= a or b;
    layer0_outputs(10918) <= a and b;
    layer0_outputs(10919) <= not b or a;
    layer0_outputs(10920) <= not (a and b);
    layer0_outputs(10921) <= a or b;
    layer0_outputs(10922) <= not a;
    layer0_outputs(10923) <= a and not b;
    layer0_outputs(10924) <= not a;
    layer0_outputs(10925) <= b and not a;
    layer0_outputs(10926) <= a or b;
    layer0_outputs(10927) <= not b or a;
    layer0_outputs(10928) <= a xor b;
    layer0_outputs(10929) <= a and b;
    layer0_outputs(10930) <= a or b;
    layer0_outputs(10931) <= a or b;
    layer0_outputs(10932) <= not (a xor b);
    layer0_outputs(10933) <= not a;
    layer0_outputs(10934) <= a and not b;
    layer0_outputs(10935) <= not (a or b);
    layer0_outputs(10936) <= not (a or b);
    layer0_outputs(10937) <= not (a or b);
    layer0_outputs(10938) <= not a or b;
    layer0_outputs(10939) <= b and not a;
    layer0_outputs(10940) <= 1'b0;
    layer0_outputs(10941) <= not a or b;
    layer0_outputs(10942) <= not b or a;
    layer0_outputs(10943) <= not b or a;
    layer0_outputs(10944) <= a and b;
    layer0_outputs(10945) <= not (a xor b);
    layer0_outputs(10946) <= not (a and b);
    layer0_outputs(10947) <= not b or a;
    layer0_outputs(10948) <= a or b;
    layer0_outputs(10949) <= not a or b;
    layer0_outputs(10950) <= b and not a;
    layer0_outputs(10951) <= not b;
    layer0_outputs(10952) <= a and b;
    layer0_outputs(10953) <= a or b;
    layer0_outputs(10954) <= a;
    layer0_outputs(10955) <= not b or a;
    layer0_outputs(10956) <= b;
    layer0_outputs(10957) <= a xor b;
    layer0_outputs(10958) <= not a;
    layer0_outputs(10959) <= a and not b;
    layer0_outputs(10960) <= a or b;
    layer0_outputs(10961) <= a or b;
    layer0_outputs(10962) <= b and not a;
    layer0_outputs(10963) <= a;
    layer0_outputs(10964) <= not b or a;
    layer0_outputs(10965) <= a xor b;
    layer0_outputs(10966) <= not a;
    layer0_outputs(10967) <= a or b;
    layer0_outputs(10968) <= not (a xor b);
    layer0_outputs(10969) <= a or b;
    layer0_outputs(10970) <= not (a xor b);
    layer0_outputs(10971) <= not (a or b);
    layer0_outputs(10972) <= not b or a;
    layer0_outputs(10973) <= not (a xor b);
    layer0_outputs(10974) <= not b;
    layer0_outputs(10975) <= not (a or b);
    layer0_outputs(10976) <= b;
    layer0_outputs(10977) <= a or b;
    layer0_outputs(10978) <= a and not b;
    layer0_outputs(10979) <= not (a or b);
    layer0_outputs(10980) <= b;
    layer0_outputs(10981) <= not a or b;
    layer0_outputs(10982) <= not (a xor b);
    layer0_outputs(10983) <= not (a or b);
    layer0_outputs(10984) <= b;
    layer0_outputs(10985) <= a and b;
    layer0_outputs(10986) <= b and not a;
    layer0_outputs(10987) <= b and not a;
    layer0_outputs(10988) <= a or b;
    layer0_outputs(10989) <= a and b;
    layer0_outputs(10990) <= a and not b;
    layer0_outputs(10991) <= not b or a;
    layer0_outputs(10992) <= a or b;
    layer0_outputs(10993) <= not (a xor b);
    layer0_outputs(10994) <= not b;
    layer0_outputs(10995) <= b and not a;
    layer0_outputs(10996) <= not (a xor b);
    layer0_outputs(10997) <= b and not a;
    layer0_outputs(10998) <= not b or a;
    layer0_outputs(10999) <= a or b;
    layer0_outputs(11000) <= b and not a;
    layer0_outputs(11001) <= not a or b;
    layer0_outputs(11002) <= a and not b;
    layer0_outputs(11003) <= not a;
    layer0_outputs(11004) <= not (a xor b);
    layer0_outputs(11005) <= a;
    layer0_outputs(11006) <= b;
    layer0_outputs(11007) <= a;
    layer0_outputs(11008) <= not b or a;
    layer0_outputs(11009) <= a or b;
    layer0_outputs(11010) <= a;
    layer0_outputs(11011) <= a and not b;
    layer0_outputs(11012) <= not (a or b);
    layer0_outputs(11013) <= a xor b;
    layer0_outputs(11014) <= b and not a;
    layer0_outputs(11015) <= 1'b0;
    layer0_outputs(11016) <= not b or a;
    layer0_outputs(11017) <= a;
    layer0_outputs(11018) <= a xor b;
    layer0_outputs(11019) <= b and not a;
    layer0_outputs(11020) <= not b or a;
    layer0_outputs(11021) <= not b;
    layer0_outputs(11022) <= not b;
    layer0_outputs(11023) <= not a;
    layer0_outputs(11024) <= a xor b;
    layer0_outputs(11025) <= a xor b;
    layer0_outputs(11026) <= not (a xor b);
    layer0_outputs(11027) <= not (a xor b);
    layer0_outputs(11028) <= not a or b;
    layer0_outputs(11029) <= not (a or b);
    layer0_outputs(11030) <= b and not a;
    layer0_outputs(11031) <= 1'b1;
    layer0_outputs(11032) <= not a or b;
    layer0_outputs(11033) <= not a or b;
    layer0_outputs(11034) <= not a or b;
    layer0_outputs(11035) <= not b;
    layer0_outputs(11036) <= b;
    layer0_outputs(11037) <= not b;
    layer0_outputs(11038) <= not (a xor b);
    layer0_outputs(11039) <= a and not b;
    layer0_outputs(11040) <= not (a or b);
    layer0_outputs(11041) <= a or b;
    layer0_outputs(11042) <= a and not b;
    layer0_outputs(11043) <= a and not b;
    layer0_outputs(11044) <= not a;
    layer0_outputs(11045) <= not (a xor b);
    layer0_outputs(11046) <= not b or a;
    layer0_outputs(11047) <= not (a xor b);
    layer0_outputs(11048) <= a xor b;
    layer0_outputs(11049) <= a xor b;
    layer0_outputs(11050) <= a or b;
    layer0_outputs(11051) <= not b;
    layer0_outputs(11052) <= not (a or b);
    layer0_outputs(11053) <= a xor b;
    layer0_outputs(11054) <= not (a xor b);
    layer0_outputs(11055) <= not b or a;
    layer0_outputs(11056) <= b;
    layer0_outputs(11057) <= a or b;
    layer0_outputs(11058) <= a xor b;
    layer0_outputs(11059) <= not (a or b);
    layer0_outputs(11060) <= a;
    layer0_outputs(11061) <= a or b;
    layer0_outputs(11062) <= b and not a;
    layer0_outputs(11063) <= a xor b;
    layer0_outputs(11064) <= a xor b;
    layer0_outputs(11065) <= not (a xor b);
    layer0_outputs(11066) <= not (a xor b);
    layer0_outputs(11067) <= b and not a;
    layer0_outputs(11068) <= a xor b;
    layer0_outputs(11069) <= not (a xor b);
    layer0_outputs(11070) <= a or b;
    layer0_outputs(11071) <= a or b;
    layer0_outputs(11072) <= not (a or b);
    layer0_outputs(11073) <= not (a or b);
    layer0_outputs(11074) <= not (a or b);
    layer0_outputs(11075) <= a and not b;
    layer0_outputs(11076) <= not b or a;
    layer0_outputs(11077) <= a and not b;
    layer0_outputs(11078) <= not (a xor b);
    layer0_outputs(11079) <= not (a xor b);
    layer0_outputs(11080) <= b and not a;
    layer0_outputs(11081) <= a or b;
    layer0_outputs(11082) <= a xor b;
    layer0_outputs(11083) <= not a or b;
    layer0_outputs(11084) <= not (a or b);
    layer0_outputs(11085) <= a and not b;
    layer0_outputs(11086) <= b and not a;
    layer0_outputs(11087) <= a;
    layer0_outputs(11088) <= b;
    layer0_outputs(11089) <= b and not a;
    layer0_outputs(11090) <= a xor b;
    layer0_outputs(11091) <= not (a or b);
    layer0_outputs(11092) <= a xor b;
    layer0_outputs(11093) <= a xor b;
    layer0_outputs(11094) <= a and not b;
    layer0_outputs(11095) <= a xor b;
    layer0_outputs(11096) <= a xor b;
    layer0_outputs(11097) <= a xor b;
    layer0_outputs(11098) <= not a;
    layer0_outputs(11099) <= not a or b;
    layer0_outputs(11100) <= not (a or b);
    layer0_outputs(11101) <= a xor b;
    layer0_outputs(11102) <= not a;
    layer0_outputs(11103) <= not (a xor b);
    layer0_outputs(11104) <= a;
    layer0_outputs(11105) <= a xor b;
    layer0_outputs(11106) <= not a or b;
    layer0_outputs(11107) <= a xor b;
    layer0_outputs(11108) <= b and not a;
    layer0_outputs(11109) <= b and not a;
    layer0_outputs(11110) <= a or b;
    layer0_outputs(11111) <= not (a xor b);
    layer0_outputs(11112) <= not b or a;
    layer0_outputs(11113) <= not (a or b);
    layer0_outputs(11114) <= not (a or b);
    layer0_outputs(11115) <= b;
    layer0_outputs(11116) <= not b or a;
    layer0_outputs(11117) <= not b;
    layer0_outputs(11118) <= a;
    layer0_outputs(11119) <= not a or b;
    layer0_outputs(11120) <= not b or a;
    layer0_outputs(11121) <= a or b;
    layer0_outputs(11122) <= a;
    layer0_outputs(11123) <= not a;
    layer0_outputs(11124) <= not b or a;
    layer0_outputs(11125) <= 1'b1;
    layer0_outputs(11126) <= b and not a;
    layer0_outputs(11127) <= not a;
    layer0_outputs(11128) <= not b or a;
    layer0_outputs(11129) <= not a or b;
    layer0_outputs(11130) <= not (a xor b);
    layer0_outputs(11131) <= not (a xor b);
    layer0_outputs(11132) <= not a;
    layer0_outputs(11133) <= a and not b;
    layer0_outputs(11134) <= not (a xor b);
    layer0_outputs(11135) <= b;
    layer0_outputs(11136) <= a and not b;
    layer0_outputs(11137) <= not (a and b);
    layer0_outputs(11138) <= a xor b;
    layer0_outputs(11139) <= a or b;
    layer0_outputs(11140) <= not (a or b);
    layer0_outputs(11141) <= b and not a;
    layer0_outputs(11142) <= a or b;
    layer0_outputs(11143) <= not (a or b);
    layer0_outputs(11144) <= not b or a;
    layer0_outputs(11145) <= not a;
    layer0_outputs(11146) <= not a or b;
    layer0_outputs(11147) <= a or b;
    layer0_outputs(11148) <= not a or b;
    layer0_outputs(11149) <= 1'b0;
    layer0_outputs(11150) <= not (a xor b);
    layer0_outputs(11151) <= b and not a;
    layer0_outputs(11152) <= not (a xor b);
    layer0_outputs(11153) <= not b or a;
    layer0_outputs(11154) <= not b;
    layer0_outputs(11155) <= not a or b;
    layer0_outputs(11156) <= not b or a;
    layer0_outputs(11157) <= a or b;
    layer0_outputs(11158) <= 1'b0;
    layer0_outputs(11159) <= a and b;
    layer0_outputs(11160) <= not (a or b);
    layer0_outputs(11161) <= not (a xor b);
    layer0_outputs(11162) <= not (a xor b);
    layer0_outputs(11163) <= a and not b;
    layer0_outputs(11164) <= not (a xor b);
    layer0_outputs(11165) <= a;
    layer0_outputs(11166) <= not b;
    layer0_outputs(11167) <= a xor b;
    layer0_outputs(11168) <= not (a xor b);
    layer0_outputs(11169) <= b and not a;
    layer0_outputs(11170) <= a or b;
    layer0_outputs(11171) <= a xor b;
    layer0_outputs(11172) <= a xor b;
    layer0_outputs(11173) <= not b;
    layer0_outputs(11174) <= b;
    layer0_outputs(11175) <= not a;
    layer0_outputs(11176) <= not b or a;
    layer0_outputs(11177) <= not b or a;
    layer0_outputs(11178) <= not (a or b);
    layer0_outputs(11179) <= not (a xor b);
    layer0_outputs(11180) <= not a or b;
    layer0_outputs(11181) <= a;
    layer0_outputs(11182) <= not (a xor b);
    layer0_outputs(11183) <= not b;
    layer0_outputs(11184) <= a and not b;
    layer0_outputs(11185) <= a or b;
    layer0_outputs(11186) <= a and b;
    layer0_outputs(11187) <= a xor b;
    layer0_outputs(11188) <= a and not b;
    layer0_outputs(11189) <= a or b;
    layer0_outputs(11190) <= not (a or b);
    layer0_outputs(11191) <= a xor b;
    layer0_outputs(11192) <= a xor b;
    layer0_outputs(11193) <= not (a or b);
    layer0_outputs(11194) <= b;
    layer0_outputs(11195) <= not a;
    layer0_outputs(11196) <= a;
    layer0_outputs(11197) <= not b;
    layer0_outputs(11198) <= a and not b;
    layer0_outputs(11199) <= not (a xor b);
    layer0_outputs(11200) <= not (a or b);
    layer0_outputs(11201) <= not (a xor b);
    layer0_outputs(11202) <= 1'b0;
    layer0_outputs(11203) <= b and not a;
    layer0_outputs(11204) <= a and not b;
    layer0_outputs(11205) <= b and not a;
    layer0_outputs(11206) <= a or b;
    layer0_outputs(11207) <= a or b;
    layer0_outputs(11208) <= not (a or b);
    layer0_outputs(11209) <= a;
    layer0_outputs(11210) <= a xor b;
    layer0_outputs(11211) <= not (a or b);
    layer0_outputs(11212) <= not (a xor b);
    layer0_outputs(11213) <= not a or b;
    layer0_outputs(11214) <= not b or a;
    layer0_outputs(11215) <= not b;
    layer0_outputs(11216) <= b and not a;
    layer0_outputs(11217) <= not b;
    layer0_outputs(11218) <= not (a xor b);
    layer0_outputs(11219) <= a and b;
    layer0_outputs(11220) <= b and not a;
    layer0_outputs(11221) <= not b or a;
    layer0_outputs(11222) <= a xor b;
    layer0_outputs(11223) <= a and not b;
    layer0_outputs(11224) <= a;
    layer0_outputs(11225) <= a;
    layer0_outputs(11226) <= b and not a;
    layer0_outputs(11227) <= not (a or b);
    layer0_outputs(11228) <= a or b;
    layer0_outputs(11229) <= a and not b;
    layer0_outputs(11230) <= 1'b0;
    layer0_outputs(11231) <= not b or a;
    layer0_outputs(11232) <= a xor b;
    layer0_outputs(11233) <= a and b;
    layer0_outputs(11234) <= a xor b;
    layer0_outputs(11235) <= a and not b;
    layer0_outputs(11236) <= not (a xor b);
    layer0_outputs(11237) <= b and not a;
    layer0_outputs(11238) <= not (a xor b);
    layer0_outputs(11239) <= a and not b;
    layer0_outputs(11240) <= a;
    layer0_outputs(11241) <= not b or a;
    layer0_outputs(11242) <= not b or a;
    layer0_outputs(11243) <= not b or a;
    layer0_outputs(11244) <= a or b;
    layer0_outputs(11245) <= a xor b;
    layer0_outputs(11246) <= a and not b;
    layer0_outputs(11247) <= not (a or b);
    layer0_outputs(11248) <= not a;
    layer0_outputs(11249) <= not (a or b);
    layer0_outputs(11250) <= a or b;
    layer0_outputs(11251) <= not a or b;
    layer0_outputs(11252) <= b and not a;
    layer0_outputs(11253) <= 1'b1;
    layer0_outputs(11254) <= a xor b;
    layer0_outputs(11255) <= a;
    layer0_outputs(11256) <= not b or a;
    layer0_outputs(11257) <= not (a or b);
    layer0_outputs(11258) <= b;
    layer0_outputs(11259) <= not (a xor b);
    layer0_outputs(11260) <= not a;
    layer0_outputs(11261) <= not a or b;
    layer0_outputs(11262) <= not (a xor b);
    layer0_outputs(11263) <= a and b;
    layer0_outputs(11264) <= not a or b;
    layer0_outputs(11265) <= a or b;
    layer0_outputs(11266) <= 1'b0;
    layer0_outputs(11267) <= not (a xor b);
    layer0_outputs(11268) <= a and not b;
    layer0_outputs(11269) <= not b;
    layer0_outputs(11270) <= a and b;
    layer0_outputs(11271) <= a;
    layer0_outputs(11272) <= not (a or b);
    layer0_outputs(11273) <= not (a or b);
    layer0_outputs(11274) <= not b;
    layer0_outputs(11275) <= a or b;
    layer0_outputs(11276) <= a and b;
    layer0_outputs(11277) <= not (a xor b);
    layer0_outputs(11278) <= not a;
    layer0_outputs(11279) <= a xor b;
    layer0_outputs(11280) <= not a;
    layer0_outputs(11281) <= a and not b;
    layer0_outputs(11282) <= not a;
    layer0_outputs(11283) <= not (a or b);
    layer0_outputs(11284) <= not a;
    layer0_outputs(11285) <= b;
    layer0_outputs(11286) <= a or b;
    layer0_outputs(11287) <= not a;
    layer0_outputs(11288) <= not a;
    layer0_outputs(11289) <= b and not a;
    layer0_outputs(11290) <= not a or b;
    layer0_outputs(11291) <= not (a xor b);
    layer0_outputs(11292) <= a and not b;
    layer0_outputs(11293) <= a or b;
    layer0_outputs(11294) <= not b or a;
    layer0_outputs(11295) <= not a;
    layer0_outputs(11296) <= not a;
    layer0_outputs(11297) <= b;
    layer0_outputs(11298) <= not (a xor b);
    layer0_outputs(11299) <= not a;
    layer0_outputs(11300) <= a and b;
    layer0_outputs(11301) <= a and not b;
    layer0_outputs(11302) <= not (a and b);
    layer0_outputs(11303) <= a or b;
    layer0_outputs(11304) <= not b;
    layer0_outputs(11305) <= a xor b;
    layer0_outputs(11306) <= a xor b;
    layer0_outputs(11307) <= not (a xor b);
    layer0_outputs(11308) <= not b;
    layer0_outputs(11309) <= not (a or b);
    layer0_outputs(11310) <= not a or b;
    layer0_outputs(11311) <= a and b;
    layer0_outputs(11312) <= not a;
    layer0_outputs(11313) <= not (a or b);
    layer0_outputs(11314) <= a or b;
    layer0_outputs(11315) <= not (a xor b);
    layer0_outputs(11316) <= a;
    layer0_outputs(11317) <= a and b;
    layer0_outputs(11318) <= b and not a;
    layer0_outputs(11319) <= b and not a;
    layer0_outputs(11320) <= b;
    layer0_outputs(11321) <= not (a or b);
    layer0_outputs(11322) <= not (a or b);
    layer0_outputs(11323) <= not (a xor b);
    layer0_outputs(11324) <= not b or a;
    layer0_outputs(11325) <= a or b;
    layer0_outputs(11326) <= not b;
    layer0_outputs(11327) <= not b or a;
    layer0_outputs(11328) <= a or b;
    layer0_outputs(11329) <= not a or b;
    layer0_outputs(11330) <= not (a or b);
    layer0_outputs(11331) <= a or b;
    layer0_outputs(11332) <= 1'b0;
    layer0_outputs(11333) <= not b;
    layer0_outputs(11334) <= 1'b1;
    layer0_outputs(11335) <= not a;
    layer0_outputs(11336) <= not a;
    layer0_outputs(11337) <= not b;
    layer0_outputs(11338) <= not (a or b);
    layer0_outputs(11339) <= a and b;
    layer0_outputs(11340) <= not (a or b);
    layer0_outputs(11341) <= not b or a;
    layer0_outputs(11342) <= b and not a;
    layer0_outputs(11343) <= not b;
    layer0_outputs(11344) <= a or b;
    layer0_outputs(11345) <= a xor b;
    layer0_outputs(11346) <= not (a or b);
    layer0_outputs(11347) <= a or b;
    layer0_outputs(11348) <= not (a xor b);
    layer0_outputs(11349) <= not (a xor b);
    layer0_outputs(11350) <= not (a or b);
    layer0_outputs(11351) <= not a or b;
    layer0_outputs(11352) <= not a;
    layer0_outputs(11353) <= a or b;
    layer0_outputs(11354) <= a and not b;
    layer0_outputs(11355) <= a;
    layer0_outputs(11356) <= not b or a;
    layer0_outputs(11357) <= not (a or b);
    layer0_outputs(11358) <= a;
    layer0_outputs(11359) <= a or b;
    layer0_outputs(11360) <= a or b;
    layer0_outputs(11361) <= a or b;
    layer0_outputs(11362) <= not (a xor b);
    layer0_outputs(11363) <= not b;
    layer0_outputs(11364) <= 1'b1;
    layer0_outputs(11365) <= b and not a;
    layer0_outputs(11366) <= a or b;
    layer0_outputs(11367) <= not (a xor b);
    layer0_outputs(11368) <= a or b;
    layer0_outputs(11369) <= 1'b1;
    layer0_outputs(11370) <= not (a or b);
    layer0_outputs(11371) <= b;
    layer0_outputs(11372) <= not b or a;
    layer0_outputs(11373) <= 1'b0;
    layer0_outputs(11374) <= a or b;
    layer0_outputs(11375) <= b;
    layer0_outputs(11376) <= a and not b;
    layer0_outputs(11377) <= b and not a;
    layer0_outputs(11378) <= a;
    layer0_outputs(11379) <= b and not a;
    layer0_outputs(11380) <= not (a or b);
    layer0_outputs(11381) <= not (a and b);
    layer0_outputs(11382) <= b;
    layer0_outputs(11383) <= a xor b;
    layer0_outputs(11384) <= not (a xor b);
    layer0_outputs(11385) <= a xor b;
    layer0_outputs(11386) <= not a;
    layer0_outputs(11387) <= not (a or b);
    layer0_outputs(11388) <= not a;
    layer0_outputs(11389) <= b;
    layer0_outputs(11390) <= not b;
    layer0_outputs(11391) <= a and b;
    layer0_outputs(11392) <= not (a or b);
    layer0_outputs(11393) <= a and not b;
    layer0_outputs(11394) <= not b or a;
    layer0_outputs(11395) <= a or b;
    layer0_outputs(11396) <= b;
    layer0_outputs(11397) <= a xor b;
    layer0_outputs(11398) <= not b or a;
    layer0_outputs(11399) <= not (a or b);
    layer0_outputs(11400) <= a or b;
    layer0_outputs(11401) <= not (a or b);
    layer0_outputs(11402) <= not b or a;
    layer0_outputs(11403) <= 1'b0;
    layer0_outputs(11404) <= a xor b;
    layer0_outputs(11405) <= not b;
    layer0_outputs(11406) <= not (a xor b);
    layer0_outputs(11407) <= not b;
    layer0_outputs(11408) <= not (a or b);
    layer0_outputs(11409) <= a and not b;
    layer0_outputs(11410) <= not (a or b);
    layer0_outputs(11411) <= a or b;
    layer0_outputs(11412) <= not a or b;
    layer0_outputs(11413) <= not a;
    layer0_outputs(11414) <= b;
    layer0_outputs(11415) <= a or b;
    layer0_outputs(11416) <= not a;
    layer0_outputs(11417) <= b;
    layer0_outputs(11418) <= b;
    layer0_outputs(11419) <= not (a xor b);
    layer0_outputs(11420) <= a and not b;
    layer0_outputs(11421) <= b and not a;
    layer0_outputs(11422) <= a xor b;
    layer0_outputs(11423) <= not a;
    layer0_outputs(11424) <= a or b;
    layer0_outputs(11425) <= not a;
    layer0_outputs(11426) <= a or b;
    layer0_outputs(11427) <= not a or b;
    layer0_outputs(11428) <= a or b;
    layer0_outputs(11429) <= not a or b;
    layer0_outputs(11430) <= not (a or b);
    layer0_outputs(11431) <= not b or a;
    layer0_outputs(11432) <= b;
    layer0_outputs(11433) <= a and b;
    layer0_outputs(11434) <= not (a or b);
    layer0_outputs(11435) <= a xor b;
    layer0_outputs(11436) <= 1'b0;
    layer0_outputs(11437) <= a and not b;
    layer0_outputs(11438) <= not (a xor b);
    layer0_outputs(11439) <= not a;
    layer0_outputs(11440) <= b and not a;
    layer0_outputs(11441) <= b;
    layer0_outputs(11442) <= a and b;
    layer0_outputs(11443) <= a xor b;
    layer0_outputs(11444) <= not a or b;
    layer0_outputs(11445) <= 1'b1;
    layer0_outputs(11446) <= a;
    layer0_outputs(11447) <= not b or a;
    layer0_outputs(11448) <= not (a xor b);
    layer0_outputs(11449) <= b;
    layer0_outputs(11450) <= b and not a;
    layer0_outputs(11451) <= not b or a;
    layer0_outputs(11452) <= a or b;
    layer0_outputs(11453) <= not a;
    layer0_outputs(11454) <= not a or b;
    layer0_outputs(11455) <= a xor b;
    layer0_outputs(11456) <= a or b;
    layer0_outputs(11457) <= not b;
    layer0_outputs(11458) <= b and not a;
    layer0_outputs(11459) <= not b or a;
    layer0_outputs(11460) <= not b;
    layer0_outputs(11461) <= b and not a;
    layer0_outputs(11462) <= not b or a;
    layer0_outputs(11463) <= a or b;
    layer0_outputs(11464) <= a xor b;
    layer0_outputs(11465) <= a or b;
    layer0_outputs(11466) <= a;
    layer0_outputs(11467) <= not b or a;
    layer0_outputs(11468) <= not b;
    layer0_outputs(11469) <= a xor b;
    layer0_outputs(11470) <= a and b;
    layer0_outputs(11471) <= not (a xor b);
    layer0_outputs(11472) <= b;
    layer0_outputs(11473) <= not a or b;
    layer0_outputs(11474) <= not (a xor b);
    layer0_outputs(11475) <= b;
    layer0_outputs(11476) <= not (a or b);
    layer0_outputs(11477) <= a;
    layer0_outputs(11478) <= b and not a;
    layer0_outputs(11479) <= a or b;
    layer0_outputs(11480) <= not b or a;
    layer0_outputs(11481) <= a or b;
    layer0_outputs(11482) <= not (a or b);
    layer0_outputs(11483) <= not a;
    layer0_outputs(11484) <= not b;
    layer0_outputs(11485) <= not (a and b);
    layer0_outputs(11486) <= a xor b;
    layer0_outputs(11487) <= 1'b0;
    layer0_outputs(11488) <= a xor b;
    layer0_outputs(11489) <= a or b;
    layer0_outputs(11490) <= not b or a;
    layer0_outputs(11491) <= not a;
    layer0_outputs(11492) <= b;
    layer0_outputs(11493) <= not b or a;
    layer0_outputs(11494) <= not b or a;
    layer0_outputs(11495) <= a and not b;
    layer0_outputs(11496) <= a or b;
    layer0_outputs(11497) <= 1'b0;
    layer0_outputs(11498) <= a xor b;
    layer0_outputs(11499) <= 1'b1;
    layer0_outputs(11500) <= not a or b;
    layer0_outputs(11501) <= not (a xor b);
    layer0_outputs(11502) <= a or b;
    layer0_outputs(11503) <= not (a or b);
    layer0_outputs(11504) <= not (a or b);
    layer0_outputs(11505) <= a and not b;
    layer0_outputs(11506) <= a or b;
    layer0_outputs(11507) <= a or b;
    layer0_outputs(11508) <= not (a or b);
    layer0_outputs(11509) <= a xor b;
    layer0_outputs(11510) <= b;
    layer0_outputs(11511) <= a or b;
    layer0_outputs(11512) <= a and not b;
    layer0_outputs(11513) <= not b or a;
    layer0_outputs(11514) <= not a;
    layer0_outputs(11515) <= not a or b;
    layer0_outputs(11516) <= a or b;
    layer0_outputs(11517) <= b;
    layer0_outputs(11518) <= not (a or b);
    layer0_outputs(11519) <= not (a xor b);
    layer0_outputs(11520) <= not a;
    layer0_outputs(11521) <= a xor b;
    layer0_outputs(11522) <= not (a or b);
    layer0_outputs(11523) <= 1'b1;
    layer0_outputs(11524) <= not b or a;
    layer0_outputs(11525) <= a or b;
    layer0_outputs(11526) <= not (a or b);
    layer0_outputs(11527) <= a or b;
    layer0_outputs(11528) <= a and b;
    layer0_outputs(11529) <= a and b;
    layer0_outputs(11530) <= b;
    layer0_outputs(11531) <= not (a or b);
    layer0_outputs(11532) <= not (a and b);
    layer0_outputs(11533) <= b and not a;
    layer0_outputs(11534) <= not (a or b);
    layer0_outputs(11535) <= b;
    layer0_outputs(11536) <= a or b;
    layer0_outputs(11537) <= not (a or b);
    layer0_outputs(11538) <= a;
    layer0_outputs(11539) <= a and not b;
    layer0_outputs(11540) <= a or b;
    layer0_outputs(11541) <= b and not a;
    layer0_outputs(11542) <= b;
    layer0_outputs(11543) <= a and not b;
    layer0_outputs(11544) <= not (a xor b);
    layer0_outputs(11545) <= not (a xor b);
    layer0_outputs(11546) <= a and not b;
    layer0_outputs(11547) <= a xor b;
    layer0_outputs(11548) <= a;
    layer0_outputs(11549) <= a or b;
    layer0_outputs(11550) <= a or b;
    layer0_outputs(11551) <= not (a or b);
    layer0_outputs(11552) <= not b or a;
    layer0_outputs(11553) <= a;
    layer0_outputs(11554) <= a xor b;
    layer0_outputs(11555) <= not (a or b);
    layer0_outputs(11556) <= not b;
    layer0_outputs(11557) <= not b or a;
    layer0_outputs(11558) <= a or b;
    layer0_outputs(11559) <= not (a and b);
    layer0_outputs(11560) <= not a;
    layer0_outputs(11561) <= not (a or b);
    layer0_outputs(11562) <= not (a or b);
    layer0_outputs(11563) <= a xor b;
    layer0_outputs(11564) <= a xor b;
    layer0_outputs(11565) <= 1'b1;
    layer0_outputs(11566) <= not (a or b);
    layer0_outputs(11567) <= not (a xor b);
    layer0_outputs(11568) <= a and not b;
    layer0_outputs(11569) <= a or b;
    layer0_outputs(11570) <= b and not a;
    layer0_outputs(11571) <= a and not b;
    layer0_outputs(11572) <= a xor b;
    layer0_outputs(11573) <= a or b;
    layer0_outputs(11574) <= not (a xor b);
    layer0_outputs(11575) <= b;
    layer0_outputs(11576) <= a or b;
    layer0_outputs(11577) <= not (a or b);
    layer0_outputs(11578) <= not a or b;
    layer0_outputs(11579) <= a;
    layer0_outputs(11580) <= a xor b;
    layer0_outputs(11581) <= not b;
    layer0_outputs(11582) <= not a;
    layer0_outputs(11583) <= not a;
    layer0_outputs(11584) <= not b or a;
    layer0_outputs(11585) <= not a;
    layer0_outputs(11586) <= not b;
    layer0_outputs(11587) <= not a;
    layer0_outputs(11588) <= not b;
    layer0_outputs(11589) <= not (a or b);
    layer0_outputs(11590) <= b and not a;
    layer0_outputs(11591) <= b and not a;
    layer0_outputs(11592) <= not b;
    layer0_outputs(11593) <= not (a or b);
    layer0_outputs(11594) <= a or b;
    layer0_outputs(11595) <= not (a xor b);
    layer0_outputs(11596) <= a;
    layer0_outputs(11597) <= b;
    layer0_outputs(11598) <= not b or a;
    layer0_outputs(11599) <= not (a xor b);
    layer0_outputs(11600) <= not (a xor b);
    layer0_outputs(11601) <= a or b;
    layer0_outputs(11602) <= a or b;
    layer0_outputs(11603) <= not (a xor b);
    layer0_outputs(11604) <= a;
    layer0_outputs(11605) <= not (a xor b);
    layer0_outputs(11606) <= a or b;
    layer0_outputs(11607) <= not b or a;
    layer0_outputs(11608) <= not (a or b);
    layer0_outputs(11609) <= not (a or b);
    layer0_outputs(11610) <= a xor b;
    layer0_outputs(11611) <= b and not a;
    layer0_outputs(11612) <= b and not a;
    layer0_outputs(11613) <= not a or b;
    layer0_outputs(11614) <= not (a xor b);
    layer0_outputs(11615) <= not a or b;
    layer0_outputs(11616) <= not (a or b);
    layer0_outputs(11617) <= a and not b;
    layer0_outputs(11618) <= a or b;
    layer0_outputs(11619) <= not b;
    layer0_outputs(11620) <= a or b;
    layer0_outputs(11621) <= a;
    layer0_outputs(11622) <= not b;
    layer0_outputs(11623) <= not b or a;
    layer0_outputs(11624) <= a xor b;
    layer0_outputs(11625) <= not a or b;
    layer0_outputs(11626) <= a;
    layer0_outputs(11627) <= a and not b;
    layer0_outputs(11628) <= a;
    layer0_outputs(11629) <= a xor b;
    layer0_outputs(11630) <= not (a or b);
    layer0_outputs(11631) <= not (a or b);
    layer0_outputs(11632) <= a;
    layer0_outputs(11633) <= not b;
    layer0_outputs(11634) <= not b or a;
    layer0_outputs(11635) <= a xor b;
    layer0_outputs(11636) <= b;
    layer0_outputs(11637) <= not (a or b);
    layer0_outputs(11638) <= a xor b;
    layer0_outputs(11639) <= 1'b1;
    layer0_outputs(11640) <= not (a or b);
    layer0_outputs(11641) <= not a or b;
    layer0_outputs(11642) <= b;
    layer0_outputs(11643) <= a;
    layer0_outputs(11644) <= not b or a;
    layer0_outputs(11645) <= not (a or b);
    layer0_outputs(11646) <= a;
    layer0_outputs(11647) <= a xor b;
    layer0_outputs(11648) <= not b;
    layer0_outputs(11649) <= a;
    layer0_outputs(11650) <= not b or a;
    layer0_outputs(11651) <= a or b;
    layer0_outputs(11652) <= 1'b0;
    layer0_outputs(11653) <= not a;
    layer0_outputs(11654) <= a and not b;
    layer0_outputs(11655) <= not (a xor b);
    layer0_outputs(11656) <= b and not a;
    layer0_outputs(11657) <= not (a and b);
    layer0_outputs(11658) <= b and not a;
    layer0_outputs(11659) <= not (a or b);
    layer0_outputs(11660) <= a xor b;
    layer0_outputs(11661) <= 1'b0;
    layer0_outputs(11662) <= not (a or b);
    layer0_outputs(11663) <= a or b;
    layer0_outputs(11664) <= not a;
    layer0_outputs(11665) <= a;
    layer0_outputs(11666) <= b and not a;
    layer0_outputs(11667) <= a and not b;
    layer0_outputs(11668) <= b;
    layer0_outputs(11669) <= not (a or b);
    layer0_outputs(11670) <= a;
    layer0_outputs(11671) <= not (a or b);
    layer0_outputs(11672) <= not b or a;
    layer0_outputs(11673) <= 1'b1;
    layer0_outputs(11674) <= a;
    layer0_outputs(11675) <= 1'b1;
    layer0_outputs(11676) <= not a or b;
    layer0_outputs(11677) <= a xor b;
    layer0_outputs(11678) <= not b or a;
    layer0_outputs(11679) <= not (a xor b);
    layer0_outputs(11680) <= b;
    layer0_outputs(11681) <= not b;
    layer0_outputs(11682) <= not (a xor b);
    layer0_outputs(11683) <= not (a xor b);
    layer0_outputs(11684) <= not (a or b);
    layer0_outputs(11685) <= not (a or b);
    layer0_outputs(11686) <= not (a or b);
    layer0_outputs(11687) <= not (a xor b);
    layer0_outputs(11688) <= not (a or b);
    layer0_outputs(11689) <= not (a or b);
    layer0_outputs(11690) <= not a;
    layer0_outputs(11691) <= a or b;
    layer0_outputs(11692) <= a and b;
    layer0_outputs(11693) <= b and not a;
    layer0_outputs(11694) <= not (a or b);
    layer0_outputs(11695) <= a or b;
    layer0_outputs(11696) <= not a;
    layer0_outputs(11697) <= 1'b1;
    layer0_outputs(11698) <= a;
    layer0_outputs(11699) <= b;
    layer0_outputs(11700) <= not (a or b);
    layer0_outputs(11701) <= 1'b0;
    layer0_outputs(11702) <= not (a or b);
    layer0_outputs(11703) <= not (a xor b);
    layer0_outputs(11704) <= b and not a;
    layer0_outputs(11705) <= b and not a;
    layer0_outputs(11706) <= a xor b;
    layer0_outputs(11707) <= not (a xor b);
    layer0_outputs(11708) <= b and not a;
    layer0_outputs(11709) <= not b or a;
    layer0_outputs(11710) <= a;
    layer0_outputs(11711) <= a;
    layer0_outputs(11712) <= b and not a;
    layer0_outputs(11713) <= b;
    layer0_outputs(11714) <= not (a or b);
    layer0_outputs(11715) <= not (a or b);
    layer0_outputs(11716) <= not (a or b);
    layer0_outputs(11717) <= 1'b0;
    layer0_outputs(11718) <= not (a or b);
    layer0_outputs(11719) <= not b;
    layer0_outputs(11720) <= not a;
    layer0_outputs(11721) <= b and not a;
    layer0_outputs(11722) <= 1'b0;
    layer0_outputs(11723) <= a xor b;
    layer0_outputs(11724) <= a and not b;
    layer0_outputs(11725) <= a or b;
    layer0_outputs(11726) <= a or b;
    layer0_outputs(11727) <= a and b;
    layer0_outputs(11728) <= a;
    layer0_outputs(11729) <= 1'b1;
    layer0_outputs(11730) <= a xor b;
    layer0_outputs(11731) <= a xor b;
    layer0_outputs(11732) <= not (a xor b);
    layer0_outputs(11733) <= not (a or b);
    layer0_outputs(11734) <= a xor b;
    layer0_outputs(11735) <= b and not a;
    layer0_outputs(11736) <= not b;
    layer0_outputs(11737) <= not a or b;
    layer0_outputs(11738) <= not b or a;
    layer0_outputs(11739) <= not (a or b);
    layer0_outputs(11740) <= not (a xor b);
    layer0_outputs(11741) <= not (a xor b);
    layer0_outputs(11742) <= not (a xor b);
    layer0_outputs(11743) <= b;
    layer0_outputs(11744) <= a xor b;
    layer0_outputs(11745) <= not (a or b);
    layer0_outputs(11746) <= b and not a;
    layer0_outputs(11747) <= a and not b;
    layer0_outputs(11748) <= not a or b;
    layer0_outputs(11749) <= b and not a;
    layer0_outputs(11750) <= not (a or b);
    layer0_outputs(11751) <= a or b;
    layer0_outputs(11752) <= a and not b;
    layer0_outputs(11753) <= a;
    layer0_outputs(11754) <= a xor b;
    layer0_outputs(11755) <= b;
    layer0_outputs(11756) <= not (a or b);
    layer0_outputs(11757) <= not (a xor b);
    layer0_outputs(11758) <= not (a or b);
    layer0_outputs(11759) <= b;
    layer0_outputs(11760) <= a or b;
    layer0_outputs(11761) <= not (a or b);
    layer0_outputs(11762) <= a or b;
    layer0_outputs(11763) <= a or b;
    layer0_outputs(11764) <= a and not b;
    layer0_outputs(11765) <= a or b;
    layer0_outputs(11766) <= b;
    layer0_outputs(11767) <= not a;
    layer0_outputs(11768) <= a xor b;
    layer0_outputs(11769) <= a xor b;
    layer0_outputs(11770) <= 1'b1;
    layer0_outputs(11771) <= not (a xor b);
    layer0_outputs(11772) <= not (a or b);
    layer0_outputs(11773) <= a;
    layer0_outputs(11774) <= b;
    layer0_outputs(11775) <= not (a or b);
    layer0_outputs(11776) <= not b or a;
    layer0_outputs(11777) <= a xor b;
    layer0_outputs(11778) <= not (a xor b);
    layer0_outputs(11779) <= not (a or b);
    layer0_outputs(11780) <= not (a xor b);
    layer0_outputs(11781) <= a xor b;
    layer0_outputs(11782) <= a or b;
    layer0_outputs(11783) <= a and b;
    layer0_outputs(11784) <= not (a or b);
    layer0_outputs(11785) <= not a or b;
    layer0_outputs(11786) <= a or b;
    layer0_outputs(11787) <= a and not b;
    layer0_outputs(11788) <= not a;
    layer0_outputs(11789) <= a or b;
    layer0_outputs(11790) <= a xor b;
    layer0_outputs(11791) <= a xor b;
    layer0_outputs(11792) <= not a or b;
    layer0_outputs(11793) <= a or b;
    layer0_outputs(11794) <= a or b;
    layer0_outputs(11795) <= a or b;
    layer0_outputs(11796) <= not (a or b);
    layer0_outputs(11797) <= not (a or b);
    layer0_outputs(11798) <= not b or a;
    layer0_outputs(11799) <= a;
    layer0_outputs(11800) <= not (a xor b);
    layer0_outputs(11801) <= a and not b;
    layer0_outputs(11802) <= not a or b;
    layer0_outputs(11803) <= not (a xor b);
    layer0_outputs(11804) <= a or b;
    layer0_outputs(11805) <= not (a or b);
    layer0_outputs(11806) <= a xor b;
    layer0_outputs(11807) <= not (a or b);
    layer0_outputs(11808) <= not a;
    layer0_outputs(11809) <= not b;
    layer0_outputs(11810) <= not a or b;
    layer0_outputs(11811) <= a;
    layer0_outputs(11812) <= a and not b;
    layer0_outputs(11813) <= not (a xor b);
    layer0_outputs(11814) <= a xor b;
    layer0_outputs(11815) <= a;
    layer0_outputs(11816) <= a xor b;
    layer0_outputs(11817) <= not (a xor b);
    layer0_outputs(11818) <= b and not a;
    layer0_outputs(11819) <= not a;
    layer0_outputs(11820) <= not (a or b);
    layer0_outputs(11821) <= a;
    layer0_outputs(11822) <= not b or a;
    layer0_outputs(11823) <= not b;
    layer0_outputs(11824) <= b;
    layer0_outputs(11825) <= a or b;
    layer0_outputs(11826) <= not (a or b);
    layer0_outputs(11827) <= b;
    layer0_outputs(11828) <= not (a or b);
    layer0_outputs(11829) <= a;
    layer0_outputs(11830) <= a and not b;
    layer0_outputs(11831) <= not (a xor b);
    layer0_outputs(11832) <= b;
    layer0_outputs(11833) <= a xor b;
    layer0_outputs(11834) <= not b or a;
    layer0_outputs(11835) <= not a;
    layer0_outputs(11836) <= not (a or b);
    layer0_outputs(11837) <= a xor b;
    layer0_outputs(11838) <= not (a or b);
    layer0_outputs(11839) <= not a;
    layer0_outputs(11840) <= a;
    layer0_outputs(11841) <= b and not a;
    layer0_outputs(11842) <= not a or b;
    layer0_outputs(11843) <= a and b;
    layer0_outputs(11844) <= b and not a;
    layer0_outputs(11845) <= not (a xor b);
    layer0_outputs(11846) <= b;
    layer0_outputs(11847) <= 1'b1;
    layer0_outputs(11848) <= not (a xor b);
    layer0_outputs(11849) <= a;
    layer0_outputs(11850) <= not (a xor b);
    layer0_outputs(11851) <= not (a xor b);
    layer0_outputs(11852) <= a or b;
    layer0_outputs(11853) <= not (a or b);
    layer0_outputs(11854) <= not (a or b);
    layer0_outputs(11855) <= a xor b;
    layer0_outputs(11856) <= a and not b;
    layer0_outputs(11857) <= not b;
    layer0_outputs(11858) <= a and not b;
    layer0_outputs(11859) <= not b;
    layer0_outputs(11860) <= not (a or b);
    layer0_outputs(11861) <= 1'b0;
    layer0_outputs(11862) <= a;
    layer0_outputs(11863) <= a or b;
    layer0_outputs(11864) <= not b;
    layer0_outputs(11865) <= not a or b;
    layer0_outputs(11866) <= b;
    layer0_outputs(11867) <= a xor b;
    layer0_outputs(11868) <= a and not b;
    layer0_outputs(11869) <= a xor b;
    layer0_outputs(11870) <= b;
    layer0_outputs(11871) <= a or b;
    layer0_outputs(11872) <= not (a xor b);
    layer0_outputs(11873) <= not a;
    layer0_outputs(11874) <= not (a xor b);
    layer0_outputs(11875) <= b and not a;
    layer0_outputs(11876) <= b and not a;
    layer0_outputs(11877) <= not (a xor b);
    layer0_outputs(11878) <= a and not b;
    layer0_outputs(11879) <= not (a or b);
    layer0_outputs(11880) <= not a;
    layer0_outputs(11881) <= a or b;
    layer0_outputs(11882) <= not (a and b);
    layer0_outputs(11883) <= a xor b;
    layer0_outputs(11884) <= b and not a;
    layer0_outputs(11885) <= a xor b;
    layer0_outputs(11886) <= a;
    layer0_outputs(11887) <= not a;
    layer0_outputs(11888) <= not (a or b);
    layer0_outputs(11889) <= b and not a;
    layer0_outputs(11890) <= a xor b;
    layer0_outputs(11891) <= a or b;
    layer0_outputs(11892) <= a xor b;
    layer0_outputs(11893) <= b;
    layer0_outputs(11894) <= a and b;
    layer0_outputs(11895) <= b and not a;
    layer0_outputs(11896) <= not (a or b);
    layer0_outputs(11897) <= a;
    layer0_outputs(11898) <= not (a xor b);
    layer0_outputs(11899) <= not b;
    layer0_outputs(11900) <= not (a xor b);
    layer0_outputs(11901) <= not (a xor b);
    layer0_outputs(11902) <= not (a and b);
    layer0_outputs(11903) <= a and b;
    layer0_outputs(11904) <= b;
    layer0_outputs(11905) <= a xor b;
    layer0_outputs(11906) <= a and b;
    layer0_outputs(11907) <= b;
    layer0_outputs(11908) <= a or b;
    layer0_outputs(11909) <= a or b;
    layer0_outputs(11910) <= a xor b;
    layer0_outputs(11911) <= a or b;
    layer0_outputs(11912) <= not (a xor b);
    layer0_outputs(11913) <= not (a xor b);
    layer0_outputs(11914) <= not (a and b);
    layer0_outputs(11915) <= a and not b;
    layer0_outputs(11916) <= a and not b;
    layer0_outputs(11917) <= a xor b;
    layer0_outputs(11918) <= not (a or b);
    layer0_outputs(11919) <= a and not b;
    layer0_outputs(11920) <= a or b;
    layer0_outputs(11921) <= not a;
    layer0_outputs(11922) <= b and not a;
    layer0_outputs(11923) <= a or b;
    layer0_outputs(11924) <= a xor b;
    layer0_outputs(11925) <= a and b;
    layer0_outputs(11926) <= not (a or b);
    layer0_outputs(11927) <= not (a xor b);
    layer0_outputs(11928) <= b;
    layer0_outputs(11929) <= a;
    layer0_outputs(11930) <= b;
    layer0_outputs(11931) <= a or b;
    layer0_outputs(11932) <= b and not a;
    layer0_outputs(11933) <= b;
    layer0_outputs(11934) <= a and b;
    layer0_outputs(11935) <= b and not a;
    layer0_outputs(11936) <= not b;
    layer0_outputs(11937) <= not a;
    layer0_outputs(11938) <= b;
    layer0_outputs(11939) <= not a;
    layer0_outputs(11940) <= not (a and b);
    layer0_outputs(11941) <= not b;
    layer0_outputs(11942) <= not (a xor b);
    layer0_outputs(11943) <= a or b;
    layer0_outputs(11944) <= not a;
    layer0_outputs(11945) <= not (a or b);
    layer0_outputs(11946) <= 1'b1;
    layer0_outputs(11947) <= a and b;
    layer0_outputs(11948) <= not b;
    layer0_outputs(11949) <= not (a xor b);
    layer0_outputs(11950) <= not (a xor b);
    layer0_outputs(11951) <= a or b;
    layer0_outputs(11952) <= a and not b;
    layer0_outputs(11953) <= a xor b;
    layer0_outputs(11954) <= a;
    layer0_outputs(11955) <= b and not a;
    layer0_outputs(11956) <= not (a xor b);
    layer0_outputs(11957) <= not (a or b);
    layer0_outputs(11958) <= not (a or b);
    layer0_outputs(11959) <= not (a xor b);
    layer0_outputs(11960) <= b and not a;
    layer0_outputs(11961) <= 1'b1;
    layer0_outputs(11962) <= a xor b;
    layer0_outputs(11963) <= a and not b;
    layer0_outputs(11964) <= not a;
    layer0_outputs(11965) <= b and not a;
    layer0_outputs(11966) <= a and not b;
    layer0_outputs(11967) <= a and b;
    layer0_outputs(11968) <= not (a or b);
    layer0_outputs(11969) <= not b;
    layer0_outputs(11970) <= 1'b1;
    layer0_outputs(11971) <= not a;
    layer0_outputs(11972) <= not (a or b);
    layer0_outputs(11973) <= not b;
    layer0_outputs(11974) <= a or b;
    layer0_outputs(11975) <= a and not b;
    layer0_outputs(11976) <= not a;
    layer0_outputs(11977) <= not b;
    layer0_outputs(11978) <= not (a or b);
    layer0_outputs(11979) <= not (a or b);
    layer0_outputs(11980) <= 1'b0;
    layer0_outputs(11981) <= 1'b0;
    layer0_outputs(11982) <= not (a xor b);
    layer0_outputs(11983) <= not b;
    layer0_outputs(11984) <= not a;
    layer0_outputs(11985) <= not (a xor b);
    layer0_outputs(11986) <= a xor b;
    layer0_outputs(11987) <= a or b;
    layer0_outputs(11988) <= not b or a;
    layer0_outputs(11989) <= not a;
    layer0_outputs(11990) <= a or b;
    layer0_outputs(11991) <= b and not a;
    layer0_outputs(11992) <= not (a xor b);
    layer0_outputs(11993) <= not (a xor b);
    layer0_outputs(11994) <= not b;
    layer0_outputs(11995) <= a and not b;
    layer0_outputs(11996) <= not (a or b);
    layer0_outputs(11997) <= a and not b;
    layer0_outputs(11998) <= a xor b;
    layer0_outputs(11999) <= not a or b;
    layer0_outputs(12000) <= not a or b;
    layer0_outputs(12001) <= not a;
    layer0_outputs(12002) <= not (a or b);
    layer0_outputs(12003) <= not a or b;
    layer0_outputs(12004) <= not a;
    layer0_outputs(12005) <= not b;
    layer0_outputs(12006) <= not (a or b);
    layer0_outputs(12007) <= b and not a;
    layer0_outputs(12008) <= a or b;
    layer0_outputs(12009) <= a or b;
    layer0_outputs(12010) <= not (a xor b);
    layer0_outputs(12011) <= not (a xor b);
    layer0_outputs(12012) <= a and not b;
    layer0_outputs(12013) <= a or b;
    layer0_outputs(12014) <= not (a xor b);
    layer0_outputs(12015) <= a or b;
    layer0_outputs(12016) <= a xor b;
    layer0_outputs(12017) <= not (a or b);
    layer0_outputs(12018) <= b and not a;
    layer0_outputs(12019) <= a xor b;
    layer0_outputs(12020) <= b;
    layer0_outputs(12021) <= not (a xor b);
    layer0_outputs(12022) <= not a;
    layer0_outputs(12023) <= not a or b;
    layer0_outputs(12024) <= not (a and b);
    layer0_outputs(12025) <= 1'b0;
    layer0_outputs(12026) <= not a;
    layer0_outputs(12027) <= not a or b;
    layer0_outputs(12028) <= 1'b0;
    layer0_outputs(12029) <= b;
    layer0_outputs(12030) <= b and not a;
    layer0_outputs(12031) <= a or b;
    layer0_outputs(12032) <= not (a or b);
    layer0_outputs(12033) <= not a;
    layer0_outputs(12034) <= not a or b;
    layer0_outputs(12035) <= a xor b;
    layer0_outputs(12036) <= not (a xor b);
    layer0_outputs(12037) <= not (a xor b);
    layer0_outputs(12038) <= a xor b;
    layer0_outputs(12039) <= not b;
    layer0_outputs(12040) <= a xor b;
    layer0_outputs(12041) <= a;
    layer0_outputs(12042) <= a xor b;
    layer0_outputs(12043) <= a and b;
    layer0_outputs(12044) <= a or b;
    layer0_outputs(12045) <= not b;
    layer0_outputs(12046) <= not b or a;
    layer0_outputs(12047) <= not a;
    layer0_outputs(12048) <= a and not b;
    layer0_outputs(12049) <= a or b;
    layer0_outputs(12050) <= b and not a;
    layer0_outputs(12051) <= not a or b;
    layer0_outputs(12052) <= not a;
    layer0_outputs(12053) <= a or b;
    layer0_outputs(12054) <= not (a or b);
    layer0_outputs(12055) <= not b;
    layer0_outputs(12056) <= not a or b;
    layer0_outputs(12057) <= a xor b;
    layer0_outputs(12058) <= b;
    layer0_outputs(12059) <= a xor b;
    layer0_outputs(12060) <= b and not a;
    layer0_outputs(12061) <= not (a or b);
    layer0_outputs(12062) <= not b;
    layer0_outputs(12063) <= not (a or b);
    layer0_outputs(12064) <= not a or b;
    layer0_outputs(12065) <= b;
    layer0_outputs(12066) <= not a or b;
    layer0_outputs(12067) <= a xor b;
    layer0_outputs(12068) <= not b or a;
    layer0_outputs(12069) <= not (a or b);
    layer0_outputs(12070) <= not b or a;
    layer0_outputs(12071) <= 1'b0;
    layer0_outputs(12072) <= b;
    layer0_outputs(12073) <= 1'b0;
    layer0_outputs(12074) <= a or b;
    layer0_outputs(12075) <= not (a and b);
    layer0_outputs(12076) <= not (a xor b);
    layer0_outputs(12077) <= a or b;
    layer0_outputs(12078) <= not a or b;
    layer0_outputs(12079) <= not b or a;
    layer0_outputs(12080) <= not b or a;
    layer0_outputs(12081) <= not (a xor b);
    layer0_outputs(12082) <= a or b;
    layer0_outputs(12083) <= not b or a;
    layer0_outputs(12084) <= a;
    layer0_outputs(12085) <= not b or a;
    layer0_outputs(12086) <= not a or b;
    layer0_outputs(12087) <= b and not a;
    layer0_outputs(12088) <= a or b;
    layer0_outputs(12089) <= not (a or b);
    layer0_outputs(12090) <= not a;
    layer0_outputs(12091) <= a;
    layer0_outputs(12092) <= not (a and b);
    layer0_outputs(12093) <= a xor b;
    layer0_outputs(12094) <= a;
    layer0_outputs(12095) <= not a or b;
    layer0_outputs(12096) <= b and not a;
    layer0_outputs(12097) <= b and not a;
    layer0_outputs(12098) <= not a;
    layer0_outputs(12099) <= not (a and b);
    layer0_outputs(12100) <= b and not a;
    layer0_outputs(12101) <= a or b;
    layer0_outputs(12102) <= not a;
    layer0_outputs(12103) <= not (a xor b);
    layer0_outputs(12104) <= not a;
    layer0_outputs(12105) <= b and not a;
    layer0_outputs(12106) <= a or b;
    layer0_outputs(12107) <= not a or b;
    layer0_outputs(12108) <= not b or a;
    layer0_outputs(12109) <= b;
    layer0_outputs(12110) <= not (a or b);
    layer0_outputs(12111) <= a;
    layer0_outputs(12112) <= a xor b;
    layer0_outputs(12113) <= 1'b0;
    layer0_outputs(12114) <= not a;
    layer0_outputs(12115) <= not a or b;
    layer0_outputs(12116) <= not a;
    layer0_outputs(12117) <= not b;
    layer0_outputs(12118) <= a or b;
    layer0_outputs(12119) <= b;
    layer0_outputs(12120) <= a xor b;
    layer0_outputs(12121) <= not (a xor b);
    layer0_outputs(12122) <= not (a or b);
    layer0_outputs(12123) <= a or b;
    layer0_outputs(12124) <= a or b;
    layer0_outputs(12125) <= a xor b;
    layer0_outputs(12126) <= a or b;
    layer0_outputs(12127) <= a or b;
    layer0_outputs(12128) <= a or b;
    layer0_outputs(12129) <= not (a xor b);
    layer0_outputs(12130) <= a xor b;
    layer0_outputs(12131) <= not (a or b);
    layer0_outputs(12132) <= a xor b;
    layer0_outputs(12133) <= a or b;
    layer0_outputs(12134) <= a;
    layer0_outputs(12135) <= a;
    layer0_outputs(12136) <= not b or a;
    layer0_outputs(12137) <= b and not a;
    layer0_outputs(12138) <= a;
    layer0_outputs(12139) <= a and not b;
    layer0_outputs(12140) <= not (a xor b);
    layer0_outputs(12141) <= b;
    layer0_outputs(12142) <= b and not a;
    layer0_outputs(12143) <= 1'b1;
    layer0_outputs(12144) <= a and not b;
    layer0_outputs(12145) <= b and not a;
    layer0_outputs(12146) <= not a or b;
    layer0_outputs(12147) <= a or b;
    layer0_outputs(12148) <= not (a xor b);
    layer0_outputs(12149) <= a xor b;
    layer0_outputs(12150) <= not (a or b);
    layer0_outputs(12151) <= a xor b;
    layer0_outputs(12152) <= b and not a;
    layer0_outputs(12153) <= not (a and b);
    layer0_outputs(12154) <= not (a or b);
    layer0_outputs(12155) <= a xor b;
    layer0_outputs(12156) <= a and not b;
    layer0_outputs(12157) <= not (a xor b);
    layer0_outputs(12158) <= not a or b;
    layer0_outputs(12159) <= not a or b;
    layer0_outputs(12160) <= not a;
    layer0_outputs(12161) <= b and not a;
    layer0_outputs(12162) <= not (a xor b);
    layer0_outputs(12163) <= b;
    layer0_outputs(12164) <= a xor b;
    layer0_outputs(12165) <= a;
    layer0_outputs(12166) <= not (a or b);
    layer0_outputs(12167) <= a or b;
    layer0_outputs(12168) <= not (a or b);
    layer0_outputs(12169) <= a or b;
    layer0_outputs(12170) <= 1'b1;
    layer0_outputs(12171) <= not a or b;
    layer0_outputs(12172) <= a;
    layer0_outputs(12173) <= not (a or b);
    layer0_outputs(12174) <= not (a or b);
    layer0_outputs(12175) <= a or b;
    layer0_outputs(12176) <= not (a and b);
    layer0_outputs(12177) <= b;
    layer0_outputs(12178) <= a or b;
    layer0_outputs(12179) <= not (a or b);
    layer0_outputs(12180) <= a and not b;
    layer0_outputs(12181) <= a or b;
    layer0_outputs(12182) <= a and not b;
    layer0_outputs(12183) <= not (a or b);
    layer0_outputs(12184) <= a or b;
    layer0_outputs(12185) <= not (a or b);
    layer0_outputs(12186) <= not (a xor b);
    layer0_outputs(12187) <= a xor b;
    layer0_outputs(12188) <= a xor b;
    layer0_outputs(12189) <= a or b;
    layer0_outputs(12190) <= a or b;
    layer0_outputs(12191) <= a xor b;
    layer0_outputs(12192) <= not a or b;
    layer0_outputs(12193) <= not b or a;
    layer0_outputs(12194) <= not (a or b);
    layer0_outputs(12195) <= not a;
    layer0_outputs(12196) <= a and not b;
    layer0_outputs(12197) <= a and not b;
    layer0_outputs(12198) <= not a;
    layer0_outputs(12199) <= not (a xor b);
    layer0_outputs(12200) <= b and not a;
    layer0_outputs(12201) <= not (a or b);
    layer0_outputs(12202) <= a and not b;
    layer0_outputs(12203) <= not (a or b);
    layer0_outputs(12204) <= a;
    layer0_outputs(12205) <= a xor b;
    layer0_outputs(12206) <= not (a or b);
    layer0_outputs(12207) <= not (a and b);
    layer0_outputs(12208) <= b and not a;
    layer0_outputs(12209) <= not (a and b);
    layer0_outputs(12210) <= not a;
    layer0_outputs(12211) <= a and not b;
    layer0_outputs(12212) <= not (a or b);
    layer0_outputs(12213) <= 1'b0;
    layer0_outputs(12214) <= a or b;
    layer0_outputs(12215) <= a xor b;
    layer0_outputs(12216) <= not (a or b);
    layer0_outputs(12217) <= a or b;
    layer0_outputs(12218) <= not (a or b);
    layer0_outputs(12219) <= b and not a;
    layer0_outputs(12220) <= not a;
    layer0_outputs(12221) <= not b;
    layer0_outputs(12222) <= not a;
    layer0_outputs(12223) <= a or b;
    layer0_outputs(12224) <= a and not b;
    layer0_outputs(12225) <= a and b;
    layer0_outputs(12226) <= a and not b;
    layer0_outputs(12227) <= a or b;
    layer0_outputs(12228) <= a xor b;
    layer0_outputs(12229) <= 1'b1;
    layer0_outputs(12230) <= not a;
    layer0_outputs(12231) <= a or b;
    layer0_outputs(12232) <= not (a xor b);
    layer0_outputs(12233) <= not b or a;
    layer0_outputs(12234) <= a or b;
    layer0_outputs(12235) <= a or b;
    layer0_outputs(12236) <= not (a xor b);
    layer0_outputs(12237) <= a or b;
    layer0_outputs(12238) <= a and b;
    layer0_outputs(12239) <= not (a or b);
    layer0_outputs(12240) <= not (a or b);
    layer0_outputs(12241) <= not (a or b);
    layer0_outputs(12242) <= not a or b;
    layer0_outputs(12243) <= a and b;
    layer0_outputs(12244) <= a and not b;
    layer0_outputs(12245) <= a xor b;
    layer0_outputs(12246) <= not a or b;
    layer0_outputs(12247) <= a or b;
    layer0_outputs(12248) <= a or b;
    layer0_outputs(12249) <= b and not a;
    layer0_outputs(12250) <= a and not b;
    layer0_outputs(12251) <= not (a or b);
    layer0_outputs(12252) <= a or b;
    layer0_outputs(12253) <= a and not b;
    layer0_outputs(12254) <= not (a or b);
    layer0_outputs(12255) <= a and not b;
    layer0_outputs(12256) <= not (a and b);
    layer0_outputs(12257) <= a or b;
    layer0_outputs(12258) <= not (a xor b);
    layer0_outputs(12259) <= a and not b;
    layer0_outputs(12260) <= 1'b0;
    layer0_outputs(12261) <= a xor b;
    layer0_outputs(12262) <= not (a or b);
    layer0_outputs(12263) <= a or b;
    layer0_outputs(12264) <= not (a or b);
    layer0_outputs(12265) <= not a;
    layer0_outputs(12266) <= a and not b;
    layer0_outputs(12267) <= a;
    layer0_outputs(12268) <= a or b;
    layer0_outputs(12269) <= not (a xor b);
    layer0_outputs(12270) <= a or b;
    layer0_outputs(12271) <= not a or b;
    layer0_outputs(12272) <= a and b;
    layer0_outputs(12273) <= not (a or b);
    layer0_outputs(12274) <= a xor b;
    layer0_outputs(12275) <= b and not a;
    layer0_outputs(12276) <= not (a or b);
    layer0_outputs(12277) <= a or b;
    layer0_outputs(12278) <= a and not b;
    layer0_outputs(12279) <= a or b;
    layer0_outputs(12280) <= not (a or b);
    layer0_outputs(12281) <= a xor b;
    layer0_outputs(12282) <= not a or b;
    layer0_outputs(12283) <= a or b;
    layer0_outputs(12284) <= not a;
    layer0_outputs(12285) <= a xor b;
    layer0_outputs(12286) <= not a;
    layer0_outputs(12287) <= not a;
    layer0_outputs(12288) <= b;
    layer0_outputs(12289) <= a;
    layer0_outputs(12290) <= a xor b;
    layer0_outputs(12291) <= not (a or b);
    layer0_outputs(12292) <= b and not a;
    layer0_outputs(12293) <= not (a or b);
    layer0_outputs(12294) <= b and not a;
    layer0_outputs(12295) <= a or b;
    layer0_outputs(12296) <= not a;
    layer0_outputs(12297) <= a or b;
    layer0_outputs(12298) <= not (a or b);
    layer0_outputs(12299) <= a or b;
    layer0_outputs(12300) <= a xor b;
    layer0_outputs(12301) <= not a;
    layer0_outputs(12302) <= a xor b;
    layer0_outputs(12303) <= a and b;
    layer0_outputs(12304) <= a or b;
    layer0_outputs(12305) <= 1'b1;
    layer0_outputs(12306) <= a xor b;
    layer0_outputs(12307) <= not (a or b);
    layer0_outputs(12308) <= a;
    layer0_outputs(12309) <= not (a or b);
    layer0_outputs(12310) <= not a;
    layer0_outputs(12311) <= a xor b;
    layer0_outputs(12312) <= not (a xor b);
    layer0_outputs(12313) <= not (a or b);
    layer0_outputs(12314) <= not a;
    layer0_outputs(12315) <= b;
    layer0_outputs(12316) <= not (a xor b);
    layer0_outputs(12317) <= a or b;
    layer0_outputs(12318) <= not (a or b);
    layer0_outputs(12319) <= b;
    layer0_outputs(12320) <= not a;
    layer0_outputs(12321) <= a xor b;
    layer0_outputs(12322) <= 1'b1;
    layer0_outputs(12323) <= not b;
    layer0_outputs(12324) <= not a;
    layer0_outputs(12325) <= a xor b;
    layer0_outputs(12326) <= a or b;
    layer0_outputs(12327) <= a;
    layer0_outputs(12328) <= b and not a;
    layer0_outputs(12329) <= a or b;
    layer0_outputs(12330) <= not b or a;
    layer0_outputs(12331) <= b and not a;
    layer0_outputs(12332) <= not (a or b);
    layer0_outputs(12333) <= a or b;
    layer0_outputs(12334) <= b;
    layer0_outputs(12335) <= not b or a;
    layer0_outputs(12336) <= not a;
    layer0_outputs(12337) <= a or b;
    layer0_outputs(12338) <= a and not b;
    layer0_outputs(12339) <= not a or b;
    layer0_outputs(12340) <= a or b;
    layer0_outputs(12341) <= b;
    layer0_outputs(12342) <= a or b;
    layer0_outputs(12343) <= a and b;
    layer0_outputs(12344) <= a and not b;
    layer0_outputs(12345) <= not b or a;
    layer0_outputs(12346) <= not (a or b);
    layer0_outputs(12347) <= not b or a;
    layer0_outputs(12348) <= a or b;
    layer0_outputs(12349) <= b and not a;
    layer0_outputs(12350) <= not b;
    layer0_outputs(12351) <= not (a xor b);
    layer0_outputs(12352) <= 1'b0;
    layer0_outputs(12353) <= not a or b;
    layer0_outputs(12354) <= not a;
    layer0_outputs(12355) <= not (a xor b);
    layer0_outputs(12356) <= a xor b;
    layer0_outputs(12357) <= not a;
    layer0_outputs(12358) <= not (a or b);
    layer0_outputs(12359) <= not b;
    layer0_outputs(12360) <= not (a or b);
    layer0_outputs(12361) <= a;
    layer0_outputs(12362) <= a;
    layer0_outputs(12363) <= not (a or b);
    layer0_outputs(12364) <= a or b;
    layer0_outputs(12365) <= 1'b0;
    layer0_outputs(12366) <= not (a xor b);
    layer0_outputs(12367) <= b and not a;
    layer0_outputs(12368) <= not (a xor b);
    layer0_outputs(12369) <= not b;
    layer0_outputs(12370) <= a and not b;
    layer0_outputs(12371) <= not (a or b);
    layer0_outputs(12372) <= not b;
    layer0_outputs(12373) <= not b or a;
    layer0_outputs(12374) <= b;
    layer0_outputs(12375) <= a xor b;
    layer0_outputs(12376) <= a or b;
    layer0_outputs(12377) <= not a or b;
    layer0_outputs(12378) <= a;
    layer0_outputs(12379) <= not (a or b);
    layer0_outputs(12380) <= a and not b;
    layer0_outputs(12381) <= not (a or b);
    layer0_outputs(12382) <= b and not a;
    layer0_outputs(12383) <= a or b;
    layer0_outputs(12384) <= not a or b;
    layer0_outputs(12385) <= not (a or b);
    layer0_outputs(12386) <= b;
    layer0_outputs(12387) <= a;
    layer0_outputs(12388) <= a xor b;
    layer0_outputs(12389) <= not b;
    layer0_outputs(12390) <= a or b;
    layer0_outputs(12391) <= b;
    layer0_outputs(12392) <= 1'b1;
    layer0_outputs(12393) <= not (a xor b);
    layer0_outputs(12394) <= not (a xor b);
    layer0_outputs(12395) <= not b;
    layer0_outputs(12396) <= not b;
    layer0_outputs(12397) <= a;
    layer0_outputs(12398) <= a or b;
    layer0_outputs(12399) <= b and not a;
    layer0_outputs(12400) <= not b;
    layer0_outputs(12401) <= a xor b;
    layer0_outputs(12402) <= not (a or b);
    layer0_outputs(12403) <= not a;
    layer0_outputs(12404) <= a or b;
    layer0_outputs(12405) <= not (a xor b);
    layer0_outputs(12406) <= a or b;
    layer0_outputs(12407) <= not b or a;
    layer0_outputs(12408) <= a or b;
    layer0_outputs(12409) <= a;
    layer0_outputs(12410) <= not (a or b);
    layer0_outputs(12411) <= not a;
    layer0_outputs(12412) <= a and not b;
    layer0_outputs(12413) <= a xor b;
    layer0_outputs(12414) <= a xor b;
    layer0_outputs(12415) <= not a or b;
    layer0_outputs(12416) <= not b;
    layer0_outputs(12417) <= a and not b;
    layer0_outputs(12418) <= not b;
    layer0_outputs(12419) <= a and not b;
    layer0_outputs(12420) <= b;
    layer0_outputs(12421) <= not a or b;
    layer0_outputs(12422) <= b and not a;
    layer0_outputs(12423) <= b and not a;
    layer0_outputs(12424) <= a or b;
    layer0_outputs(12425) <= not (a xor b);
    layer0_outputs(12426) <= a xor b;
    layer0_outputs(12427) <= not (a and b);
    layer0_outputs(12428) <= not a;
    layer0_outputs(12429) <= b and not a;
    layer0_outputs(12430) <= b;
    layer0_outputs(12431) <= not b;
    layer0_outputs(12432) <= a;
    layer0_outputs(12433) <= a or b;
    layer0_outputs(12434) <= not a;
    layer0_outputs(12435) <= a xor b;
    layer0_outputs(12436) <= 1'b0;
    layer0_outputs(12437) <= a xor b;
    layer0_outputs(12438) <= not a;
    layer0_outputs(12439) <= b and not a;
    layer0_outputs(12440) <= not a;
    layer0_outputs(12441) <= not a;
    layer0_outputs(12442) <= not (a xor b);
    layer0_outputs(12443) <= a;
    layer0_outputs(12444) <= a xor b;
    layer0_outputs(12445) <= not (a xor b);
    layer0_outputs(12446) <= a;
    layer0_outputs(12447) <= not (a xor b);
    layer0_outputs(12448) <= not b or a;
    layer0_outputs(12449) <= not (a xor b);
    layer0_outputs(12450) <= not a or b;
    layer0_outputs(12451) <= b and not a;
    layer0_outputs(12452) <= not (a or b);
    layer0_outputs(12453) <= not b;
    layer0_outputs(12454) <= a xor b;
    layer0_outputs(12455) <= not (a or b);
    layer0_outputs(12456) <= a xor b;
    layer0_outputs(12457) <= b;
    layer0_outputs(12458) <= a and not b;
    layer0_outputs(12459) <= a xor b;
    layer0_outputs(12460) <= a;
    layer0_outputs(12461) <= not a or b;
    layer0_outputs(12462) <= not b or a;
    layer0_outputs(12463) <= a;
    layer0_outputs(12464) <= not b or a;
    layer0_outputs(12465) <= b;
    layer0_outputs(12466) <= a xor b;
    layer0_outputs(12467) <= a or b;
    layer0_outputs(12468) <= not a;
    layer0_outputs(12469) <= a or b;
    layer0_outputs(12470) <= b;
    layer0_outputs(12471) <= a or b;
    layer0_outputs(12472) <= not (a or b);
    layer0_outputs(12473) <= a or b;
    layer0_outputs(12474) <= not (a xor b);
    layer0_outputs(12475) <= not (a or b);
    layer0_outputs(12476) <= a;
    layer0_outputs(12477) <= 1'b1;
    layer0_outputs(12478) <= b;
    layer0_outputs(12479) <= not (a xor b);
    layer0_outputs(12480) <= a or b;
    layer0_outputs(12481) <= a and b;
    layer0_outputs(12482) <= not b;
    layer0_outputs(12483) <= not b or a;
    layer0_outputs(12484) <= not b;
    layer0_outputs(12485) <= b and not a;
    layer0_outputs(12486) <= a and not b;
    layer0_outputs(12487) <= not a;
    layer0_outputs(12488) <= a and not b;
    layer0_outputs(12489) <= not (a or b);
    layer0_outputs(12490) <= not (a xor b);
    layer0_outputs(12491) <= not a or b;
    layer0_outputs(12492) <= a and not b;
    layer0_outputs(12493) <= a or b;
    layer0_outputs(12494) <= b;
    layer0_outputs(12495) <= not a;
    layer0_outputs(12496) <= a or b;
    layer0_outputs(12497) <= a or b;
    layer0_outputs(12498) <= b;
    layer0_outputs(12499) <= a;
    layer0_outputs(12500) <= not (a or b);
    layer0_outputs(12501) <= not (a xor b);
    layer0_outputs(12502) <= b and not a;
    layer0_outputs(12503) <= not (a xor b);
    layer0_outputs(12504) <= not (a xor b);
    layer0_outputs(12505) <= a xor b;
    layer0_outputs(12506) <= a or b;
    layer0_outputs(12507) <= b;
    layer0_outputs(12508) <= not (a or b);
    layer0_outputs(12509) <= a or b;
    layer0_outputs(12510) <= not a or b;
    layer0_outputs(12511) <= a and not b;
    layer0_outputs(12512) <= a;
    layer0_outputs(12513) <= not a or b;
    layer0_outputs(12514) <= not a or b;
    layer0_outputs(12515) <= a or b;
    layer0_outputs(12516) <= a or b;
    layer0_outputs(12517) <= not (a or b);
    layer0_outputs(12518) <= 1'b1;
    layer0_outputs(12519) <= not (a or b);
    layer0_outputs(12520) <= a xor b;
    layer0_outputs(12521) <= not (a xor b);
    layer0_outputs(12522) <= a and b;
    layer0_outputs(12523) <= 1'b0;
    layer0_outputs(12524) <= not (a or b);
    layer0_outputs(12525) <= a or b;
    layer0_outputs(12526) <= not (a xor b);
    layer0_outputs(12527) <= a and b;
    layer0_outputs(12528) <= a;
    layer0_outputs(12529) <= a xor b;
    layer0_outputs(12530) <= a and b;
    layer0_outputs(12531) <= a or b;
    layer0_outputs(12532) <= a;
    layer0_outputs(12533) <= not (a or b);
    layer0_outputs(12534) <= not (a xor b);
    layer0_outputs(12535) <= not a;
    layer0_outputs(12536) <= a and not b;
    layer0_outputs(12537) <= a or b;
    layer0_outputs(12538) <= not a or b;
    layer0_outputs(12539) <= a xor b;
    layer0_outputs(12540) <= a xor b;
    layer0_outputs(12541) <= b;
    layer0_outputs(12542) <= a and not b;
    layer0_outputs(12543) <= b and not a;
    layer0_outputs(12544) <= a or b;
    layer0_outputs(12545) <= a and not b;
    layer0_outputs(12546) <= not (a xor b);
    layer0_outputs(12547) <= a or b;
    layer0_outputs(12548) <= not (a or b);
    layer0_outputs(12549) <= not (a or b);
    layer0_outputs(12550) <= a;
    layer0_outputs(12551) <= a xor b;
    layer0_outputs(12552) <= not (a or b);
    layer0_outputs(12553) <= a or b;
    layer0_outputs(12554) <= not a;
    layer0_outputs(12555) <= 1'b1;
    layer0_outputs(12556) <= a;
    layer0_outputs(12557) <= not (a xor b);
    layer0_outputs(12558) <= a;
    layer0_outputs(12559) <= a or b;
    layer0_outputs(12560) <= a xor b;
    layer0_outputs(12561) <= not (a or b);
    layer0_outputs(12562) <= not b;
    layer0_outputs(12563) <= not (a or b);
    layer0_outputs(12564) <= a;
    layer0_outputs(12565) <= not a;
    layer0_outputs(12566) <= a and not b;
    layer0_outputs(12567) <= a or b;
    layer0_outputs(12568) <= a;
    layer0_outputs(12569) <= not b;
    layer0_outputs(12570) <= not a or b;
    layer0_outputs(12571) <= not b or a;
    layer0_outputs(12572) <= a or b;
    layer0_outputs(12573) <= a and not b;
    layer0_outputs(12574) <= not (a or b);
    layer0_outputs(12575) <= a xor b;
    layer0_outputs(12576) <= not a;
    layer0_outputs(12577) <= not b;
    layer0_outputs(12578) <= not a;
    layer0_outputs(12579) <= b;
    layer0_outputs(12580) <= not a;
    layer0_outputs(12581) <= b;
    layer0_outputs(12582) <= not (a or b);
    layer0_outputs(12583) <= a and not b;
    layer0_outputs(12584) <= b and not a;
    layer0_outputs(12585) <= a or b;
    layer0_outputs(12586) <= not (a or b);
    layer0_outputs(12587) <= a or b;
    layer0_outputs(12588) <= not (a or b);
    layer0_outputs(12589) <= not b or a;
    layer0_outputs(12590) <= not a or b;
    layer0_outputs(12591) <= a;
    layer0_outputs(12592) <= not b;
    layer0_outputs(12593) <= not a or b;
    layer0_outputs(12594) <= not b or a;
    layer0_outputs(12595) <= b and not a;
    layer0_outputs(12596) <= a;
    layer0_outputs(12597) <= a and not b;
    layer0_outputs(12598) <= not a;
    layer0_outputs(12599) <= not (a or b);
    layer0_outputs(12600) <= not (a or b);
    layer0_outputs(12601) <= a xor b;
    layer0_outputs(12602) <= a or b;
    layer0_outputs(12603) <= not b;
    layer0_outputs(12604) <= b;
    layer0_outputs(12605) <= not a;
    layer0_outputs(12606) <= b;
    layer0_outputs(12607) <= not b or a;
    layer0_outputs(12608) <= not b;
    layer0_outputs(12609) <= a or b;
    layer0_outputs(12610) <= a xor b;
    layer0_outputs(12611) <= not a or b;
    layer0_outputs(12612) <= a xor b;
    layer0_outputs(12613) <= not (a or b);
    layer0_outputs(12614) <= a or b;
    layer0_outputs(12615) <= a;
    layer0_outputs(12616) <= not (a xor b);
    layer0_outputs(12617) <= not a or b;
    layer0_outputs(12618) <= not (a or b);
    layer0_outputs(12619) <= a;
    layer0_outputs(12620) <= a and not b;
    layer0_outputs(12621) <= b and not a;
    layer0_outputs(12622) <= not (a xor b);
    layer0_outputs(12623) <= 1'b0;
    layer0_outputs(12624) <= not (a xor b);
    layer0_outputs(12625) <= a;
    layer0_outputs(12626) <= a and b;
    layer0_outputs(12627) <= not a or b;
    layer0_outputs(12628) <= a;
    layer0_outputs(12629) <= a;
    layer0_outputs(12630) <= not b or a;
    layer0_outputs(12631) <= not (a or b);
    layer0_outputs(12632) <= a or b;
    layer0_outputs(12633) <= not b or a;
    layer0_outputs(12634) <= not (a or b);
    layer0_outputs(12635) <= not (a or b);
    layer0_outputs(12636) <= not (a or b);
    layer0_outputs(12637) <= a or b;
    layer0_outputs(12638) <= a;
    layer0_outputs(12639) <= a and not b;
    layer0_outputs(12640) <= not (a xor b);
    layer0_outputs(12641) <= not (a xor b);
    layer0_outputs(12642) <= not (a and b);
    layer0_outputs(12643) <= not b or a;
    layer0_outputs(12644) <= b;
    layer0_outputs(12645) <= not a or b;
    layer0_outputs(12646) <= a xor b;
    layer0_outputs(12647) <= not b or a;
    layer0_outputs(12648) <= not a;
    layer0_outputs(12649) <= a xor b;
    layer0_outputs(12650) <= not (a or b);
    layer0_outputs(12651) <= not b or a;
    layer0_outputs(12652) <= not a;
    layer0_outputs(12653) <= not (a xor b);
    layer0_outputs(12654) <= 1'b0;
    layer0_outputs(12655) <= a or b;
    layer0_outputs(12656) <= not (a or b);
    layer0_outputs(12657) <= b and not a;
    layer0_outputs(12658) <= a;
    layer0_outputs(12659) <= not a;
    layer0_outputs(12660) <= a;
    layer0_outputs(12661) <= not b;
    layer0_outputs(12662) <= not a or b;
    layer0_outputs(12663) <= a;
    layer0_outputs(12664) <= not a or b;
    layer0_outputs(12665) <= not (a xor b);
    layer0_outputs(12666) <= not (a xor b);
    layer0_outputs(12667) <= not (a or b);
    layer0_outputs(12668) <= not (a or b);
    layer0_outputs(12669) <= not (a or b);
    layer0_outputs(12670) <= not a;
    layer0_outputs(12671) <= not b or a;
    layer0_outputs(12672) <= a xor b;
    layer0_outputs(12673) <= not (a xor b);
    layer0_outputs(12674) <= a xor b;
    layer0_outputs(12675) <= 1'b1;
    layer0_outputs(12676) <= not a or b;
    layer0_outputs(12677) <= not b;
    layer0_outputs(12678) <= a xor b;
    layer0_outputs(12679) <= not a or b;
    layer0_outputs(12680) <= a or b;
    layer0_outputs(12681) <= 1'b1;
    layer0_outputs(12682) <= a xor b;
    layer0_outputs(12683) <= not (a xor b);
    layer0_outputs(12684) <= a or b;
    layer0_outputs(12685) <= not b;
    layer0_outputs(12686) <= a and b;
    layer0_outputs(12687) <= b;
    layer0_outputs(12688) <= a xor b;
    layer0_outputs(12689) <= a and not b;
    layer0_outputs(12690) <= a or b;
    layer0_outputs(12691) <= not (a xor b);
    layer0_outputs(12692) <= a and not b;
    layer0_outputs(12693) <= not (a or b);
    layer0_outputs(12694) <= a xor b;
    layer0_outputs(12695) <= a xor b;
    layer0_outputs(12696) <= not (a or b);
    layer0_outputs(12697) <= not b;
    layer0_outputs(12698) <= not a or b;
    layer0_outputs(12699) <= a or b;
    layer0_outputs(12700) <= not b;
    layer0_outputs(12701) <= not (a or b);
    layer0_outputs(12702) <= a and not b;
    layer0_outputs(12703) <= not (a xor b);
    layer0_outputs(12704) <= not b;
    layer0_outputs(12705) <= a xor b;
    layer0_outputs(12706) <= not b or a;
    layer0_outputs(12707) <= not b;
    layer0_outputs(12708) <= b and not a;
    layer0_outputs(12709) <= b;
    layer0_outputs(12710) <= not (a xor b);
    layer0_outputs(12711) <= a xor b;
    layer0_outputs(12712) <= b;
    layer0_outputs(12713) <= not b;
    layer0_outputs(12714) <= not (a or b);
    layer0_outputs(12715) <= not (a or b);
    layer0_outputs(12716) <= not (a and b);
    layer0_outputs(12717) <= not b or a;
    layer0_outputs(12718) <= a xor b;
    layer0_outputs(12719) <= b and not a;
    layer0_outputs(12720) <= a and not b;
    layer0_outputs(12721) <= a and not b;
    layer0_outputs(12722) <= a;
    layer0_outputs(12723) <= not (a or b);
    layer0_outputs(12724) <= a or b;
    layer0_outputs(12725) <= 1'b0;
    layer0_outputs(12726) <= a and not b;
    layer0_outputs(12727) <= a;
    layer0_outputs(12728) <= not (a or b);
    layer0_outputs(12729) <= a xor b;
    layer0_outputs(12730) <= not a or b;
    layer0_outputs(12731) <= a;
    layer0_outputs(12732) <= a and not b;
    layer0_outputs(12733) <= not a or b;
    layer0_outputs(12734) <= a;
    layer0_outputs(12735) <= a xor b;
    layer0_outputs(12736) <= a xor b;
    layer0_outputs(12737) <= a or b;
    layer0_outputs(12738) <= a and not b;
    layer0_outputs(12739) <= not (a xor b);
    layer0_outputs(12740) <= not a;
    layer0_outputs(12741) <= 1'b0;
    layer0_outputs(12742) <= not (a and b);
    layer0_outputs(12743) <= a;
    layer0_outputs(12744) <= a xor b;
    layer0_outputs(12745) <= a or b;
    layer0_outputs(12746) <= b and not a;
    layer0_outputs(12747) <= a xor b;
    layer0_outputs(12748) <= a or b;
    layer0_outputs(12749) <= not b;
    layer0_outputs(12750) <= a and not b;
    layer0_outputs(12751) <= b and not a;
    layer0_outputs(12752) <= not (a or b);
    layer0_outputs(12753) <= not a or b;
    layer0_outputs(12754) <= not a or b;
    layer0_outputs(12755) <= not (a xor b);
    layer0_outputs(12756) <= not a;
    layer0_outputs(12757) <= a and not b;
    layer0_outputs(12758) <= b;
    layer0_outputs(12759) <= a and not b;
    layer0_outputs(12760) <= a or b;
    layer0_outputs(12761) <= not b;
    layer0_outputs(12762) <= a xor b;
    layer0_outputs(12763) <= not (a or b);
    layer0_outputs(12764) <= not a;
    layer0_outputs(12765) <= a and not b;
    layer0_outputs(12766) <= a or b;
    layer0_outputs(12767) <= a;
    layer0_outputs(12768) <= a or b;
    layer0_outputs(12769) <= not b or a;
    layer0_outputs(12770) <= not b or a;
    layer0_outputs(12771) <= not a;
    layer0_outputs(12772) <= not (a or b);
    layer0_outputs(12773) <= b;
    layer0_outputs(12774) <= not (a xor b);
    layer0_outputs(12775) <= b;
    layer0_outputs(12776) <= a or b;
    layer0_outputs(12777) <= a xor b;
    layer0_outputs(12778) <= a xor b;
    layer0_outputs(12779) <= not a or b;
    layer0_outputs(12780) <= not b;
    layer0_outputs(12781) <= a or b;
    layer0_outputs(12782) <= a;
    layer0_outputs(12783) <= 1'b1;
    layer0_outputs(12784) <= b and not a;
    layer0_outputs(12785) <= 1'b1;
    layer0_outputs(12786) <= not a;
    layer0_outputs(12787) <= not b;
    layer0_outputs(12788) <= b;
    layer0_outputs(12789) <= b;
    layer0_outputs(12790) <= not (a or b);
    layer0_outputs(12791) <= a xor b;
    layer0_outputs(12792) <= not (a or b);
    layer0_outputs(12793) <= not (a or b);
    layer0_outputs(12794) <= a and not b;
    layer0_outputs(12795) <= not a or b;
    layer0_outputs(12796) <= not a;
    layer0_outputs(12797) <= a xor b;
    layer0_outputs(12798) <= a xor b;
    layer0_outputs(12799) <= not (a xor b);
    outputs(0) <= a xor b;
    outputs(1) <= not a;
    outputs(2) <= a xor b;
    outputs(3) <= not a;
    outputs(4) <= a xor b;
    outputs(5) <= not (a xor b);
    outputs(6) <= a xor b;
    outputs(7) <= not (a xor b);
    outputs(8) <= not a;
    outputs(9) <= b;
    outputs(10) <= not a or b;
    outputs(11) <= a;
    outputs(12) <= not (a xor b);
    outputs(13) <= b;
    outputs(14) <= not b;
    outputs(15) <= not (a or b);
    outputs(16) <= not (a or b);
    outputs(17) <= a xor b;
    outputs(18) <= b and not a;
    outputs(19) <= b and not a;
    outputs(20) <= not b;
    outputs(21) <= not (a xor b);
    outputs(22) <= a;
    outputs(23) <= b and not a;
    outputs(24) <= b and not a;
    outputs(25) <= not a;
    outputs(26) <= not (a xor b);
    outputs(27) <= not b or a;
    outputs(28) <= a;
    outputs(29) <= a and b;
    outputs(30) <= not a;
    outputs(31) <= not b or a;
    outputs(32) <= b;
    outputs(33) <= not (a xor b);
    outputs(34) <= not b;
    outputs(35) <= a xor b;
    outputs(36) <= a xor b;
    outputs(37) <= not b;
    outputs(38) <= not a;
    outputs(39) <= a and b;
    outputs(40) <= not b;
    outputs(41) <= b;
    outputs(42) <= b;
    outputs(43) <= not b;
    outputs(44) <= a xor b;
    outputs(45) <= a;
    outputs(46) <= not (a xor b);
    outputs(47) <= b;
    outputs(48) <= not b;
    outputs(49) <= a or b;
    outputs(50) <= a xor b;
    outputs(51) <= not a;
    outputs(52) <= a xor b;
    outputs(53) <= a xor b;
    outputs(54) <= a;
    outputs(55) <= b and not a;
    outputs(56) <= not b;
    outputs(57) <= b;
    outputs(58) <= not (a xor b);
    outputs(59) <= a xor b;
    outputs(60) <= not (a xor b);
    outputs(61) <= a;
    outputs(62) <= a xor b;
    outputs(63) <= a or b;
    outputs(64) <= not (a xor b);
    outputs(65) <= not a;
    outputs(66) <= b;
    outputs(67) <= a xor b;
    outputs(68) <= not (a or b);
    outputs(69) <= b;
    outputs(70) <= not a;
    outputs(71) <= not a or b;
    outputs(72) <= a;
    outputs(73) <= not b;
    outputs(74) <= a and b;
    outputs(75) <= a xor b;
    outputs(76) <= not (a xor b);
    outputs(77) <= a;
    outputs(78) <= a and not b;
    outputs(79) <= a xor b;
    outputs(80) <= not b;
    outputs(81) <= b;
    outputs(82) <= not b;
    outputs(83) <= a xor b;
    outputs(84) <= a and not b;
    outputs(85) <= b;
    outputs(86) <= a and not b;
    outputs(87) <= not b;
    outputs(88) <= a and not b;
    outputs(89) <= not b;
    outputs(90) <= a xor b;
    outputs(91) <= a xor b;
    outputs(92) <= b;
    outputs(93) <= not b;
    outputs(94) <= not b or a;
    outputs(95) <= not a;
    outputs(96) <= a xor b;
    outputs(97) <= a;
    outputs(98) <= not (a xor b);
    outputs(99) <= not a;
    outputs(100) <= a xor b;
    outputs(101) <= not b;
    outputs(102) <= not a;
    outputs(103) <= not (a and b);
    outputs(104) <= a xor b;
    outputs(105) <= b and not a;
    outputs(106) <= not b;
    outputs(107) <= not a;
    outputs(108) <= a and b;
    outputs(109) <= a and not b;
    outputs(110) <= b;
    outputs(111) <= b and not a;
    outputs(112) <= a xor b;
    outputs(113) <= not a;
    outputs(114) <= not a;
    outputs(115) <= a xor b;
    outputs(116) <= not a;
    outputs(117) <= not (a xor b);
    outputs(118) <= a xor b;
    outputs(119) <= not (a xor b);
    outputs(120) <= a xor b;
    outputs(121) <= not (a or b);
    outputs(122) <= not b;
    outputs(123) <= not a;
    outputs(124) <= not b;
    outputs(125) <= a xor b;
    outputs(126) <= not a;
    outputs(127) <= not (a xor b);
    outputs(128) <= not a;
    outputs(129) <= a xor b;
    outputs(130) <= not b;
    outputs(131) <= not b;
    outputs(132) <= not (a or b);
    outputs(133) <= a xor b;
    outputs(134) <= a and b;
    outputs(135) <= not (a and b);
    outputs(136) <= b;
    outputs(137) <= not (a or b);
    outputs(138) <= a and b;
    outputs(139) <= b;
    outputs(140) <= not (a xor b);
    outputs(141) <= b;
    outputs(142) <= a xor b;
    outputs(143) <= not (a xor b);
    outputs(144) <= not a;
    outputs(145) <= not (a or b);
    outputs(146) <= a and not b;
    outputs(147) <= not b;
    outputs(148) <= a;
    outputs(149) <= not (a xor b);
    outputs(150) <= not b;
    outputs(151) <= not a;
    outputs(152) <= a or b;
    outputs(153) <= not (a and b);
    outputs(154) <= a or b;
    outputs(155) <= not (a xor b);
    outputs(156) <= not a or b;
    outputs(157) <= a xor b;
    outputs(158) <= a and b;
    outputs(159) <= not b;
    outputs(160) <= not (a xor b);
    outputs(161) <= a and not b;
    outputs(162) <= a xor b;
    outputs(163) <= not b;
    outputs(164) <= a;
    outputs(165) <= not b;
    outputs(166) <= a xor b;
    outputs(167) <= a and not b;
    outputs(168) <= not b;
    outputs(169) <= a and not b;
    outputs(170) <= b and not a;
    outputs(171) <= b and not a;
    outputs(172) <= a xor b;
    outputs(173) <= a and not b;
    outputs(174) <= b;
    outputs(175) <= a;
    outputs(176) <= not b;
    outputs(177) <= not (a xor b);
    outputs(178) <= not a;
    outputs(179) <= a;
    outputs(180) <= a xor b;
    outputs(181) <= b;
    outputs(182) <= not b;
    outputs(183) <= not (a xor b);
    outputs(184) <= a or b;
    outputs(185) <= a and b;
    outputs(186) <= a;
    outputs(187) <= not (a xor b);
    outputs(188) <= a and b;
    outputs(189) <= not a;
    outputs(190) <= not a or b;
    outputs(191) <= not a;
    outputs(192) <= not a;
    outputs(193) <= not (a and b);
    outputs(194) <= not (a and b);
    outputs(195) <= a and b;
    outputs(196) <= a xor b;
    outputs(197) <= not (a or b);
    outputs(198) <= not b or a;
    outputs(199) <= a;
    outputs(200) <= b;
    outputs(201) <= a xor b;
    outputs(202) <= a xor b;
    outputs(203) <= not b;
    outputs(204) <= b;
    outputs(205) <= not (a xor b);
    outputs(206) <= a and b;
    outputs(207) <= a and not b;
    outputs(208) <= a xor b;
    outputs(209) <= a and b;
    outputs(210) <= a or b;
    outputs(211) <= a and b;
    outputs(212) <= b;
    outputs(213) <= not (a or b);
    outputs(214) <= not a;
    outputs(215) <= a and not b;
    outputs(216) <= a and b;
    outputs(217) <= not (a and b);
    outputs(218) <= not a;
    outputs(219) <= b;
    outputs(220) <= b;
    outputs(221) <= not (a xor b);
    outputs(222) <= a or b;
    outputs(223) <= a;
    outputs(224) <= not (a and b);
    outputs(225) <= a;
    outputs(226) <= a;
    outputs(227) <= a xor b;
    outputs(228) <= b and not a;
    outputs(229) <= a;
    outputs(230) <= b and not a;
    outputs(231) <= not (a xor b);
    outputs(232) <= not b;
    outputs(233) <= a or b;
    outputs(234) <= a xor b;
    outputs(235) <= a;
    outputs(236) <= a xor b;
    outputs(237) <= not a;
    outputs(238) <= a;
    outputs(239) <= b;
    outputs(240) <= not (a xor b);
    outputs(241) <= b;
    outputs(242) <= b and not a;
    outputs(243) <= a xor b;
    outputs(244) <= not (a xor b);
    outputs(245) <= a xor b;
    outputs(246) <= not a;
    outputs(247) <= a xor b;
    outputs(248) <= a;
    outputs(249) <= b;
    outputs(250) <= not (a or b);
    outputs(251) <= not (a and b);
    outputs(252) <= not (a xor b);
    outputs(253) <= not (a or b);
    outputs(254) <= a and not b;
    outputs(255) <= a;
    outputs(256) <= a;
    outputs(257) <= a;
    outputs(258) <= a xor b;
    outputs(259) <= not b;
    outputs(260) <= not a or b;
    outputs(261) <= a;
    outputs(262) <= not (a and b);
    outputs(263) <= a xor b;
    outputs(264) <= a;
    outputs(265) <= b;
    outputs(266) <= not (a xor b);
    outputs(267) <= not a or b;
    outputs(268) <= a xor b;
    outputs(269) <= a and not b;
    outputs(270) <= not b;
    outputs(271) <= not a;
    outputs(272) <= not a;
    outputs(273) <= not b;
    outputs(274) <= a xor b;
    outputs(275) <= not (a xor b);
    outputs(276) <= b and not a;
    outputs(277) <= a;
    outputs(278) <= a;
    outputs(279) <= a or b;
    outputs(280) <= not (a and b);
    outputs(281) <= a and not b;
    outputs(282) <= a and not b;
    outputs(283) <= a xor b;
    outputs(284) <= a xor b;
    outputs(285) <= not a;
    outputs(286) <= not b;
    outputs(287) <= not (a xor b);
    outputs(288) <= b;
    outputs(289) <= a xor b;
    outputs(290) <= a or b;
    outputs(291) <= not (a xor b);
    outputs(292) <= a or b;
    outputs(293) <= not b;
    outputs(294) <= a and b;
    outputs(295) <= b;
    outputs(296) <= a and b;
    outputs(297) <= not b or a;
    outputs(298) <= not a;
    outputs(299) <= a or b;
    outputs(300) <= a;
    outputs(301) <= not b or a;
    outputs(302) <= not b;
    outputs(303) <= b;
    outputs(304) <= not a;
    outputs(305) <= not b;
    outputs(306) <= not b;
    outputs(307) <= not a;
    outputs(308) <= b;
    outputs(309) <= a or b;
    outputs(310) <= not (a or b);
    outputs(311) <= a;
    outputs(312) <= a xor b;
    outputs(313) <= not a;
    outputs(314) <= a;
    outputs(315) <= a xor b;
    outputs(316) <= a and b;
    outputs(317) <= a;
    outputs(318) <= not a or b;
    outputs(319) <= not (a xor b);
    outputs(320) <= not (a or b);
    outputs(321) <= a and not b;
    outputs(322) <= not (a xor b);
    outputs(323) <= not b;
    outputs(324) <= not a;
    outputs(325) <= not a;
    outputs(326) <= not b;
    outputs(327) <= b;
    outputs(328) <= not a;
    outputs(329) <= a and b;
    outputs(330) <= not b;
    outputs(331) <= not a;
    outputs(332) <= not (a xor b);
    outputs(333) <= a;
    outputs(334) <= b;
    outputs(335) <= not b;
    outputs(336) <= a and b;
    outputs(337) <= a;
    outputs(338) <= a xor b;
    outputs(339) <= a xor b;
    outputs(340) <= not (a or b);
    outputs(341) <= b and not a;
    outputs(342) <= not (a xor b);
    outputs(343) <= not a;
    outputs(344) <= a or b;
    outputs(345) <= a and b;
    outputs(346) <= a and b;
    outputs(347) <= b;
    outputs(348) <= a and not b;
    outputs(349) <= not (a or b);
    outputs(350) <= b;
    outputs(351) <= not (a and b);
    outputs(352) <= a and b;
    outputs(353) <= not a;
    outputs(354) <= not (a or b);
    outputs(355) <= a and not b;
    outputs(356) <= a xor b;
    outputs(357) <= a;
    outputs(358) <= a and b;
    outputs(359) <= not (a xor b);
    outputs(360) <= not (a xor b);
    outputs(361) <= a xor b;
    outputs(362) <= b and not a;
    outputs(363) <= a xor b;
    outputs(364) <= not b;
    outputs(365) <= a and b;
    outputs(366) <= a and b;
    outputs(367) <= b;
    outputs(368) <= not (a or b);
    outputs(369) <= b and not a;
    outputs(370) <= a xor b;
    outputs(371) <= b;
    outputs(372) <= not (a xor b);
    outputs(373) <= not a;
    outputs(374) <= not (a or b);
    outputs(375) <= not (a xor b);
    outputs(376) <= not (a xor b);
    outputs(377) <= a xor b;
    outputs(378) <= not b;
    outputs(379) <= 1'b0;
    outputs(380) <= not b;
    outputs(381) <= not a;
    outputs(382) <= not b;
    outputs(383) <= b;
    outputs(384) <= not (a xor b);
    outputs(385) <= a and not b;
    outputs(386) <= not b;
    outputs(387) <= not b;
    outputs(388) <= a or b;
    outputs(389) <= a;
    outputs(390) <= not b;
    outputs(391) <= not b or a;
    outputs(392) <= not b;
    outputs(393) <= a xor b;
    outputs(394) <= b;
    outputs(395) <= a xor b;
    outputs(396) <= not a;
    outputs(397) <= a;
    outputs(398) <= a and not b;
    outputs(399) <= b;
    outputs(400) <= not b or a;
    outputs(401) <= a and b;
    outputs(402) <= not (a xor b);
    outputs(403) <= not b or a;
    outputs(404) <= a;
    outputs(405) <= not (a or b);
    outputs(406) <= not (a xor b);
    outputs(407) <= not a;
    outputs(408) <= a xor b;
    outputs(409) <= b and not a;
    outputs(410) <= a;
    outputs(411) <= a and b;
    outputs(412) <= not (a xor b);
    outputs(413) <= a;
    outputs(414) <= a and not b;
    outputs(415) <= a xor b;
    outputs(416) <= b;
    outputs(417) <= not b;
    outputs(418) <= a xor b;
    outputs(419) <= a xor b;
    outputs(420) <= a xor b;
    outputs(421) <= not (a xor b);
    outputs(422) <= not a;
    outputs(423) <= b;
    outputs(424) <= not a or b;
    outputs(425) <= a;
    outputs(426) <= b;
    outputs(427) <= not (a or b);
    outputs(428) <= not b or a;
    outputs(429) <= b;
    outputs(430) <= not (a xor b);
    outputs(431) <= a and not b;
    outputs(432) <= b;
    outputs(433) <= a and not b;
    outputs(434) <= not a;
    outputs(435) <= not (a or b);
    outputs(436) <= not a or b;
    outputs(437) <= a;
    outputs(438) <= b and not a;
    outputs(439) <= not a;
    outputs(440) <= not b;
    outputs(441) <= not (a xor b);
    outputs(442) <= b and not a;
    outputs(443) <= not b;
    outputs(444) <= a;
    outputs(445) <= a and not b;
    outputs(446) <= not a;
    outputs(447) <= not a;
    outputs(448) <= a xor b;
    outputs(449) <= a xor b;
    outputs(450) <= a and not b;
    outputs(451) <= not (a xor b);
    outputs(452) <= a xor b;
    outputs(453) <= not a;
    outputs(454) <= not b;
    outputs(455) <= not a;
    outputs(456) <= not a;
    outputs(457) <= b and not a;
    outputs(458) <= not (a and b);
    outputs(459) <= not a;
    outputs(460) <= b;
    outputs(461) <= a;
    outputs(462) <= b;
    outputs(463) <= a xor b;
    outputs(464) <= a xor b;
    outputs(465) <= a and not b;
    outputs(466) <= a xor b;
    outputs(467) <= not (a xor b);
    outputs(468) <= b and not a;
    outputs(469) <= not (a xor b);
    outputs(470) <= b;
    outputs(471) <= not b;
    outputs(472) <= a xor b;
    outputs(473) <= not a;
    outputs(474) <= a;
    outputs(475) <= not a;
    outputs(476) <= not a;
    outputs(477) <= a xor b;
    outputs(478) <= a xor b;
    outputs(479) <= a and not b;
    outputs(480) <= not b or a;
    outputs(481) <= b;
    outputs(482) <= not (a xor b);
    outputs(483) <= b;
    outputs(484) <= b;
    outputs(485) <= not (a xor b);
    outputs(486) <= not b;
    outputs(487) <= not (a xor b);
    outputs(488) <= a and b;
    outputs(489) <= not a;
    outputs(490) <= b;
    outputs(491) <= a or b;
    outputs(492) <= not a;
    outputs(493) <= not a;
    outputs(494) <= not b;
    outputs(495) <= b;
    outputs(496) <= a xor b;
    outputs(497) <= b;
    outputs(498) <= not a;
    outputs(499) <= a or b;
    outputs(500) <= a and b;
    outputs(501) <= not a;
    outputs(502) <= not b;
    outputs(503) <= a and not b;
    outputs(504) <= not a;
    outputs(505) <= b;
    outputs(506) <= not (a and b);
    outputs(507) <= a;
    outputs(508) <= a;
    outputs(509) <= a xor b;
    outputs(510) <= b and not a;
    outputs(511) <= a and not b;
    outputs(512) <= a and b;
    outputs(513) <= not (a xor b);
    outputs(514) <= not b;
    outputs(515) <= b and not a;
    outputs(516) <= a xor b;
    outputs(517) <= a and not b;
    outputs(518) <= not (a or b);
    outputs(519) <= a xor b;
    outputs(520) <= not (a xor b);
    outputs(521) <= b;
    outputs(522) <= a xor b;
    outputs(523) <= not a;
    outputs(524) <= not (a xor b);
    outputs(525) <= not a;
    outputs(526) <= a xor b;
    outputs(527) <= b;
    outputs(528) <= a;
    outputs(529) <= not b;
    outputs(530) <= a and not b;
    outputs(531) <= not b;
    outputs(532) <= not a or b;
    outputs(533) <= b;
    outputs(534) <= not a;
    outputs(535) <= not a;
    outputs(536) <= a and b;
    outputs(537) <= not b;
    outputs(538) <= not (a and b);
    outputs(539) <= not a;
    outputs(540) <= not (a xor b);
    outputs(541) <= not b;
    outputs(542) <= a;
    outputs(543) <= not (a xor b);
    outputs(544) <= not (a xor b);
    outputs(545) <= not b or a;
    outputs(546) <= a and b;
    outputs(547) <= a and b;
    outputs(548) <= not (a xor b);
    outputs(549) <= not b;
    outputs(550) <= not a or b;
    outputs(551) <= a;
    outputs(552) <= a and not b;
    outputs(553) <= b;
    outputs(554) <= a xor b;
    outputs(555) <= b and not a;
    outputs(556) <= b and not a;
    outputs(557) <= a xor b;
    outputs(558) <= b;
    outputs(559) <= not (a and b);
    outputs(560) <= not (a xor b);
    outputs(561) <= a and not b;
    outputs(562) <= not (a or b);
    outputs(563) <= not (a and b);
    outputs(564) <= not (a xor b);
    outputs(565) <= not a;
    outputs(566) <= a xor b;
    outputs(567) <= a;
    outputs(568) <= not b;
    outputs(569) <= not a;
    outputs(570) <= a;
    outputs(571) <= not (a or b);
    outputs(572) <= a;
    outputs(573) <= b;
    outputs(574) <= not a;
    outputs(575) <= not (a xor b);
    outputs(576) <= b and not a;
    outputs(577) <= a;
    outputs(578) <= not a;
    outputs(579) <= not (a xor b);
    outputs(580) <= a;
    outputs(581) <= a xor b;
    outputs(582) <= a;
    outputs(583) <= b and not a;
    outputs(584) <= a and b;
    outputs(585) <= not b;
    outputs(586) <= not a;
    outputs(587) <= a xor b;
    outputs(588) <= a and b;
    outputs(589) <= a xor b;
    outputs(590) <= a;
    outputs(591) <= a and not b;
    outputs(592) <= not b;
    outputs(593) <= not a;
    outputs(594) <= not a;
    outputs(595) <= not a or b;
    outputs(596) <= b;
    outputs(597) <= not (a or b);
    outputs(598) <= a;
    outputs(599) <= a xor b;
    outputs(600) <= a;
    outputs(601) <= b;
    outputs(602) <= a and not b;
    outputs(603) <= not b;
    outputs(604) <= a;
    outputs(605) <= b;
    outputs(606) <= not (a xor b);
    outputs(607) <= a and b;
    outputs(608) <= a and not b;
    outputs(609) <= a;
    outputs(610) <= b;
    outputs(611) <= not b or a;
    outputs(612) <= not a or b;
    outputs(613) <= a xor b;
    outputs(614) <= not (a xor b);
    outputs(615) <= a xor b;
    outputs(616) <= a xor b;
    outputs(617) <= a xor b;
    outputs(618) <= not a;
    outputs(619) <= a;
    outputs(620) <= b and not a;
    outputs(621) <= not a or b;
    outputs(622) <= a;
    outputs(623) <= b;
    outputs(624) <= not b;
    outputs(625) <= a xor b;
    outputs(626) <= not b or a;
    outputs(627) <= a;
    outputs(628) <= not (a xor b);
    outputs(629) <= a or b;
    outputs(630) <= b;
    outputs(631) <= a and b;
    outputs(632) <= not (a or b);
    outputs(633) <= a and not b;
    outputs(634) <= a xor b;
    outputs(635) <= a;
    outputs(636) <= b;
    outputs(637) <= a;
    outputs(638) <= b;
    outputs(639) <= b and not a;
    outputs(640) <= b;
    outputs(641) <= b;
    outputs(642) <= not b;
    outputs(643) <= not (a xor b);
    outputs(644) <= a xor b;
    outputs(645) <= not (a xor b);
    outputs(646) <= b;
    outputs(647) <= not (a xor b);
    outputs(648) <= a or b;
    outputs(649) <= not b;
    outputs(650) <= not b;
    outputs(651) <= a;
    outputs(652) <= not a or b;
    outputs(653) <= not a or b;
    outputs(654) <= not (a xor b);
    outputs(655) <= not a;
    outputs(656) <= not b;
    outputs(657) <= not a;
    outputs(658) <= a or b;
    outputs(659) <= b;
    outputs(660) <= not (a xor b);
    outputs(661) <= not (a or b);
    outputs(662) <= a;
    outputs(663) <= a;
    outputs(664) <= b;
    outputs(665) <= b;
    outputs(666) <= not a;
    outputs(667) <= not (a xor b);
    outputs(668) <= b;
    outputs(669) <= b;
    outputs(670) <= a xor b;
    outputs(671) <= a and not b;
    outputs(672) <= b and not a;
    outputs(673) <= not (a xor b);
    outputs(674) <= a;
    outputs(675) <= b;
    outputs(676) <= a xor b;
    outputs(677) <= not b;
    outputs(678) <= a xor b;
    outputs(679) <= not a or b;
    outputs(680) <= a;
    outputs(681) <= not a;
    outputs(682) <= not (a xor b);
    outputs(683) <= not (a xor b);
    outputs(684) <= a xor b;
    outputs(685) <= a and not b;
    outputs(686) <= not b;
    outputs(687) <= not a or b;
    outputs(688) <= not (a xor b);
    outputs(689) <= a xor b;
    outputs(690) <= a;
    outputs(691) <= not (a xor b);
    outputs(692) <= not (a and b);
    outputs(693) <= a xor b;
    outputs(694) <= a and b;
    outputs(695) <= a xor b;
    outputs(696) <= not a;
    outputs(697) <= a;
    outputs(698) <= a xor b;
    outputs(699) <= not (a or b);
    outputs(700) <= a xor b;
    outputs(701) <= a xor b;
    outputs(702) <= b;
    outputs(703) <= a;
    outputs(704) <= not b;
    outputs(705) <= b;
    outputs(706) <= not a or b;
    outputs(707) <= not a;
    outputs(708) <= a;
    outputs(709) <= a and not b;
    outputs(710) <= not a;
    outputs(711) <= a xor b;
    outputs(712) <= a xor b;
    outputs(713) <= not b;
    outputs(714) <= not a or b;
    outputs(715) <= a and b;
    outputs(716) <= not b or a;
    outputs(717) <= a and not b;
    outputs(718) <= a and not b;
    outputs(719) <= a and not b;
    outputs(720) <= a;
    outputs(721) <= not a or b;
    outputs(722) <= b;
    outputs(723) <= not a;
    outputs(724) <= not b;
    outputs(725) <= a xor b;
    outputs(726) <= not b;
    outputs(727) <= a or b;
    outputs(728) <= a xor b;
    outputs(729) <= not (a xor b);
    outputs(730) <= b and not a;
    outputs(731) <= not (a or b);
    outputs(732) <= a;
    outputs(733) <= not (a or b);
    outputs(734) <= a;
    outputs(735) <= a;
    outputs(736) <= a and not b;
    outputs(737) <= b;
    outputs(738) <= a xor b;
    outputs(739) <= b;
    outputs(740) <= a and not b;
    outputs(741) <= a;
    outputs(742) <= a and not b;
    outputs(743) <= not a;
    outputs(744) <= not a;
    outputs(745) <= a or b;
    outputs(746) <= not a;
    outputs(747) <= a;
    outputs(748) <= a or b;
    outputs(749) <= a and not b;
    outputs(750) <= a xor b;
    outputs(751) <= a or b;
    outputs(752) <= a or b;
    outputs(753) <= not a;
    outputs(754) <= not a or b;
    outputs(755) <= a;
    outputs(756) <= b;
    outputs(757) <= not a;
    outputs(758) <= not a;
    outputs(759) <= a xor b;
    outputs(760) <= not b;
    outputs(761) <= a xor b;
    outputs(762) <= not (a and b);
    outputs(763) <= not b;
    outputs(764) <= a;
    outputs(765) <= b and not a;
    outputs(766) <= not b;
    outputs(767) <= not a;
    outputs(768) <= not a;
    outputs(769) <= a xor b;
    outputs(770) <= a;
    outputs(771) <= a xor b;
    outputs(772) <= a and b;
    outputs(773) <= b and not a;
    outputs(774) <= a;
    outputs(775) <= a xor b;
    outputs(776) <= a xor b;
    outputs(777) <= not a;
    outputs(778) <= a;
    outputs(779) <= not (a xor b);
    outputs(780) <= not (a and b);
    outputs(781) <= a and not b;
    outputs(782) <= a and not b;
    outputs(783) <= not b;
    outputs(784) <= not b;
    outputs(785) <= not (a xor b);
    outputs(786) <= a;
    outputs(787) <= not a;
    outputs(788) <= not (a xor b);
    outputs(789) <= not b;
    outputs(790) <= a and not b;
    outputs(791) <= not (a xor b);
    outputs(792) <= not b;
    outputs(793) <= not (a xor b);
    outputs(794) <= a;
    outputs(795) <= not (a xor b);
    outputs(796) <= not (a xor b);
    outputs(797) <= not b;
    outputs(798) <= b and not a;
    outputs(799) <= not b or a;
    outputs(800) <= not b or a;
    outputs(801) <= not b;
    outputs(802) <= not (a xor b);
    outputs(803) <= not (a xor b);
    outputs(804) <= a xor b;
    outputs(805) <= not a;
    outputs(806) <= a or b;
    outputs(807) <= not a or b;
    outputs(808) <= b and not a;
    outputs(809) <= a xor b;
    outputs(810) <= a xor b;
    outputs(811) <= a xor b;
    outputs(812) <= not a;
    outputs(813) <= a and not b;
    outputs(814) <= not a;
    outputs(815) <= a;
    outputs(816) <= not a;
    outputs(817) <= not (a xor b);
    outputs(818) <= not a;
    outputs(819) <= not b;
    outputs(820) <= not a;
    outputs(821) <= a xor b;
    outputs(822) <= not a;
    outputs(823) <= not (a xor b);
    outputs(824) <= not a;
    outputs(825) <= a and not b;
    outputs(826) <= a;
    outputs(827) <= a;
    outputs(828) <= not a;
    outputs(829) <= not (a or b);
    outputs(830) <= not a;
    outputs(831) <= not a;
    outputs(832) <= not (a xor b);
    outputs(833) <= not b;
    outputs(834) <= b;
    outputs(835) <= a and b;
    outputs(836) <= b;
    outputs(837) <= a xor b;
    outputs(838) <= not (a xor b);
    outputs(839) <= a;
    outputs(840) <= b;
    outputs(841) <= a xor b;
    outputs(842) <= b;
    outputs(843) <= a and not b;
    outputs(844) <= not a;
    outputs(845) <= a;
    outputs(846) <= not (a or b);
    outputs(847) <= b and not a;
    outputs(848) <= not b;
    outputs(849) <= not a;
    outputs(850) <= not (a and b);
    outputs(851) <= not b;
    outputs(852) <= not (a xor b);
    outputs(853) <= not b or a;
    outputs(854) <= b;
    outputs(855) <= b;
    outputs(856) <= not b;
    outputs(857) <= not (a xor b);
    outputs(858) <= a;
    outputs(859) <= not a;
    outputs(860) <= not b;
    outputs(861) <= not (a or b);
    outputs(862) <= b;
    outputs(863) <= not (a xor b);
    outputs(864) <= b;
    outputs(865) <= a;
    outputs(866) <= a;
    outputs(867) <= a;
    outputs(868) <= not (a xor b);
    outputs(869) <= not (a xor b);
    outputs(870) <= not (a xor b);
    outputs(871) <= b;
    outputs(872) <= a and b;
    outputs(873) <= b and not a;
    outputs(874) <= not (a xor b);
    outputs(875) <= b;
    outputs(876) <= a and b;
    outputs(877) <= a;
    outputs(878) <= b;
    outputs(879) <= not b;
    outputs(880) <= not (a or b);
    outputs(881) <= not b;
    outputs(882) <= not (a or b);
    outputs(883) <= b;
    outputs(884) <= b;
    outputs(885) <= a and b;
    outputs(886) <= not b or a;
    outputs(887) <= not b or a;
    outputs(888) <= not b or a;
    outputs(889) <= b;
    outputs(890) <= a xor b;
    outputs(891) <= b and not a;
    outputs(892) <= b;
    outputs(893) <= a;
    outputs(894) <= not (a or b);
    outputs(895) <= a;
    outputs(896) <= not b;
    outputs(897) <= a and not b;
    outputs(898) <= a;
    outputs(899) <= a and b;
    outputs(900) <= not (a xor b);
    outputs(901) <= not (a or b);
    outputs(902) <= not (a xor b);
    outputs(903) <= a;
    outputs(904) <= not (a or b);
    outputs(905) <= a xor b;
    outputs(906) <= not (a xor b);
    outputs(907) <= a;
    outputs(908) <= b;
    outputs(909) <= b and not a;
    outputs(910) <= b;
    outputs(911) <= not b;
    outputs(912) <= a or b;
    outputs(913) <= a xor b;
    outputs(914) <= not (a xor b);
    outputs(915) <= not b;
    outputs(916) <= a and not b;
    outputs(917) <= 1'b1;
    outputs(918) <= a and not b;
    outputs(919) <= not b;
    outputs(920) <= not (a or b);
    outputs(921) <= a;
    outputs(922) <= not a;
    outputs(923) <= not (a xor b);
    outputs(924) <= a;
    outputs(925) <= not (a or b);
    outputs(926) <= not a;
    outputs(927) <= not b;
    outputs(928) <= a xor b;
    outputs(929) <= b;
    outputs(930) <= a;
    outputs(931) <= not b;
    outputs(932) <= a xor b;
    outputs(933) <= not (a and b);
    outputs(934) <= not b;
    outputs(935) <= a and not b;
    outputs(936) <= a or b;
    outputs(937) <= not (a or b);
    outputs(938) <= a and b;
    outputs(939) <= b and not a;
    outputs(940) <= a;
    outputs(941) <= a or b;
    outputs(942) <= not b or a;
    outputs(943) <= b;
    outputs(944) <= a xor b;
    outputs(945) <= a and not b;
    outputs(946) <= a and b;
    outputs(947) <= a xor b;
    outputs(948) <= not a;
    outputs(949) <= b and not a;
    outputs(950) <= not (a xor b);
    outputs(951) <= not a or b;
    outputs(952) <= not b;
    outputs(953) <= not b;
    outputs(954) <= a xor b;
    outputs(955) <= a and not b;
    outputs(956) <= not (a and b);
    outputs(957) <= not (a xor b);
    outputs(958) <= a;
    outputs(959) <= not (a xor b);
    outputs(960) <= not a;
    outputs(961) <= b;
    outputs(962) <= not (a xor b);
    outputs(963) <= a xor b;
    outputs(964) <= a;
    outputs(965) <= b and not a;
    outputs(966) <= b;
    outputs(967) <= not (a xor b);
    outputs(968) <= a xor b;
    outputs(969) <= not b or a;
    outputs(970) <= not b;
    outputs(971) <= b;
    outputs(972) <= a xor b;
    outputs(973) <= a;
    outputs(974) <= b;
    outputs(975) <= a xor b;
    outputs(976) <= b;
    outputs(977) <= not a;
    outputs(978) <= b;
    outputs(979) <= a;
    outputs(980) <= not a;
    outputs(981) <= b and not a;
    outputs(982) <= b and not a;
    outputs(983) <= a xor b;
    outputs(984) <= a xor b;
    outputs(985) <= a;
    outputs(986) <= a and not b;
    outputs(987) <= b;
    outputs(988) <= a;
    outputs(989) <= b;
    outputs(990) <= a;
    outputs(991) <= not (a xor b);
    outputs(992) <= not a;
    outputs(993) <= b;
    outputs(994) <= b;
    outputs(995) <= a or b;
    outputs(996) <= b and not a;
    outputs(997) <= not b or a;
    outputs(998) <= a and not b;
    outputs(999) <= b;
    outputs(1000) <= not b;
    outputs(1001) <= b;
    outputs(1002) <= not (a or b);
    outputs(1003) <= a;
    outputs(1004) <= a xor b;
    outputs(1005) <= a;
    outputs(1006) <= not (a or b);
    outputs(1007) <= not (a xor b);
    outputs(1008) <= not (a xor b);
    outputs(1009) <= b;
    outputs(1010) <= b;
    outputs(1011) <= not a;
    outputs(1012) <= not b;
    outputs(1013) <= not (a xor b);
    outputs(1014) <= not (a xor b);
    outputs(1015) <= b and not a;
    outputs(1016) <= not (a xor b);
    outputs(1017) <= not b or a;
    outputs(1018) <= a xor b;
    outputs(1019) <= not (a xor b);
    outputs(1020) <= a;
    outputs(1021) <= a;
    outputs(1022) <= not (a or b);
    outputs(1023) <= a;
    outputs(1024) <= not a or b;
    outputs(1025) <= b;
    outputs(1026) <= not (a xor b);
    outputs(1027) <= b and not a;
    outputs(1028) <= b;
    outputs(1029) <= not b;
    outputs(1030) <= a;
    outputs(1031) <= not (a xor b);
    outputs(1032) <= b;
    outputs(1033) <= not (a xor b);
    outputs(1034) <= not a;
    outputs(1035) <= a xor b;
    outputs(1036) <= a;
    outputs(1037) <= not b or a;
    outputs(1038) <= not a;
    outputs(1039) <= not (a xor b);
    outputs(1040) <= b;
    outputs(1041) <= a and not b;
    outputs(1042) <= a;
    outputs(1043) <= not b;
    outputs(1044) <= a and not b;
    outputs(1045) <= not a or b;
    outputs(1046) <= a xor b;
    outputs(1047) <= not b;
    outputs(1048) <= not a;
    outputs(1049) <= not a;
    outputs(1050) <= not (a or b);
    outputs(1051) <= b;
    outputs(1052) <= a;
    outputs(1053) <= not b;
    outputs(1054) <= a and not b;
    outputs(1055) <= not a;
    outputs(1056) <= not a;
    outputs(1057) <= a xor b;
    outputs(1058) <= a and not b;
    outputs(1059) <= b;
    outputs(1060) <= not (a or b);
    outputs(1061) <= a xor b;
    outputs(1062) <= b and not a;
    outputs(1063) <= not a;
    outputs(1064) <= b;
    outputs(1065) <= a xor b;
    outputs(1066) <= b;
    outputs(1067) <= not a;
    outputs(1068) <= not (a and b);
    outputs(1069) <= a and b;
    outputs(1070) <= b;
    outputs(1071) <= a or b;
    outputs(1072) <= a and b;
    outputs(1073) <= not a;
    outputs(1074) <= not (a and b);
    outputs(1075) <= b;
    outputs(1076) <= a xor b;
    outputs(1077) <= b;
    outputs(1078) <= a;
    outputs(1079) <= b and not a;
    outputs(1080) <= a and not b;
    outputs(1081) <= b;
    outputs(1082) <= a xor b;
    outputs(1083) <= not a;
    outputs(1084) <= a xor b;
    outputs(1085) <= not b;
    outputs(1086) <= b;
    outputs(1087) <= a and not b;
    outputs(1088) <= not b or a;
    outputs(1089) <= not a;
    outputs(1090) <= not (a xor b);
    outputs(1091) <= not a;
    outputs(1092) <= a;
    outputs(1093) <= a xor b;
    outputs(1094) <= not (a xor b);
    outputs(1095) <= not (a xor b);
    outputs(1096) <= a xor b;
    outputs(1097) <= not a;
    outputs(1098) <= a;
    outputs(1099) <= b and not a;
    outputs(1100) <= not a;
    outputs(1101) <= not (a xor b);
    outputs(1102) <= b;
    outputs(1103) <= not (a xor b);
    outputs(1104) <= a and b;
    outputs(1105) <= not b or a;
    outputs(1106) <= a xor b;
    outputs(1107) <= b;
    outputs(1108) <= a and not b;
    outputs(1109) <= a xor b;
    outputs(1110) <= not (a xor b);
    outputs(1111) <= not (a and b);
    outputs(1112) <= not (a xor b);
    outputs(1113) <= not b;
    outputs(1114) <= a and b;
    outputs(1115) <= a;
    outputs(1116) <= a xor b;
    outputs(1117) <= not (a or b);
    outputs(1118) <= a xor b;
    outputs(1119) <= a xor b;
    outputs(1120) <= not (a xor b);
    outputs(1121) <= not a or b;
    outputs(1122) <= not a;
    outputs(1123) <= not (a and b);
    outputs(1124) <= not b;
    outputs(1125) <= not a;
    outputs(1126) <= not a or b;
    outputs(1127) <= a or b;
    outputs(1128) <= b;
    outputs(1129) <= not (a and b);
    outputs(1130) <= a and b;
    outputs(1131) <= not (a or b);
    outputs(1132) <= a xor b;
    outputs(1133) <= b;
    outputs(1134) <= a xor b;
    outputs(1135) <= a xor b;
    outputs(1136) <= not b;
    outputs(1137) <= not (a xor b);
    outputs(1138) <= not a;
    outputs(1139) <= a and b;
    outputs(1140) <= b;
    outputs(1141) <= not (a and b);
    outputs(1142) <= a;
    outputs(1143) <= a xor b;
    outputs(1144) <= a or b;
    outputs(1145) <= a;
    outputs(1146) <= b;
    outputs(1147) <= b and not a;
    outputs(1148) <= a;
    outputs(1149) <= a xor b;
    outputs(1150) <= b;
    outputs(1151) <= a and not b;
    outputs(1152) <= not (a xor b);
    outputs(1153) <= b;
    outputs(1154) <= not (a or b);
    outputs(1155) <= b;
    outputs(1156) <= not (a or b);
    outputs(1157) <= not (a or b);
    outputs(1158) <= a;
    outputs(1159) <= a or b;
    outputs(1160) <= not (a xor b);
    outputs(1161) <= not a or b;
    outputs(1162) <= a or b;
    outputs(1163) <= not b;
    outputs(1164) <= not a or b;
    outputs(1165) <= not (a and b);
    outputs(1166) <= not a;
    outputs(1167) <= not (a and b);
    outputs(1168) <= a;
    outputs(1169) <= a xor b;
    outputs(1170) <= b and not a;
    outputs(1171) <= a;
    outputs(1172) <= a or b;
    outputs(1173) <= a;
    outputs(1174) <= a;
    outputs(1175) <= not a;
    outputs(1176) <= not a;
    outputs(1177) <= a;
    outputs(1178) <= b;
    outputs(1179) <= not a;
    outputs(1180) <= a;
    outputs(1181) <= a and not b;
    outputs(1182) <= a xor b;
    outputs(1183) <= not a;
    outputs(1184) <= a xor b;
    outputs(1185) <= a xor b;
    outputs(1186) <= not a;
    outputs(1187) <= a xor b;
    outputs(1188) <= not b;
    outputs(1189) <= a;
    outputs(1190) <= not a;
    outputs(1191) <= not b;
    outputs(1192) <= a;
    outputs(1193) <= a xor b;
    outputs(1194) <= a xor b;
    outputs(1195) <= not (a or b);
    outputs(1196) <= a or b;
    outputs(1197) <= b;
    outputs(1198) <= a xor b;
    outputs(1199) <= a or b;
    outputs(1200) <= b;
    outputs(1201) <= a xor b;
    outputs(1202) <= not (a xor b);
    outputs(1203) <= not (a and b);
    outputs(1204) <= not a;
    outputs(1205) <= not (a xor b);
    outputs(1206) <= not (a xor b);
    outputs(1207) <= a xor b;
    outputs(1208) <= not (a and b);
    outputs(1209) <= a xor b;
    outputs(1210) <= not (a xor b);
    outputs(1211) <= not a or b;
    outputs(1212) <= not a;
    outputs(1213) <= a xor b;
    outputs(1214) <= b;
    outputs(1215) <= not b;
    outputs(1216) <= a xor b;
    outputs(1217) <= a;
    outputs(1218) <= b;
    outputs(1219) <= not a;
    outputs(1220) <= not b;
    outputs(1221) <= a xor b;
    outputs(1222) <= b;
    outputs(1223) <= not b;
    outputs(1224) <= not a;
    outputs(1225) <= a or b;
    outputs(1226) <= not a;
    outputs(1227) <= not a;
    outputs(1228) <= not b;
    outputs(1229) <= a;
    outputs(1230) <= b;
    outputs(1231) <= not (a and b);
    outputs(1232) <= not (a xor b);
    outputs(1233) <= a;
    outputs(1234) <= a and b;
    outputs(1235) <= a and b;
    outputs(1236) <= a xor b;
    outputs(1237) <= not b or a;
    outputs(1238) <= a xor b;
    outputs(1239) <= not b;
    outputs(1240) <= not a;
    outputs(1241) <= a xor b;
    outputs(1242) <= not (a or b);
    outputs(1243) <= not a;
    outputs(1244) <= not b;
    outputs(1245) <= not a;
    outputs(1246) <= a and b;
    outputs(1247) <= not b;
    outputs(1248) <= a xor b;
    outputs(1249) <= a xor b;
    outputs(1250) <= not (a or b);
    outputs(1251) <= not a;
    outputs(1252) <= not (a and b);
    outputs(1253) <= a;
    outputs(1254) <= not a;
    outputs(1255) <= not (a xor b);
    outputs(1256) <= not a;
    outputs(1257) <= b and not a;
    outputs(1258) <= not (a xor b);
    outputs(1259) <= a xor b;
    outputs(1260) <= a and not b;
    outputs(1261) <= a;
    outputs(1262) <= b and not a;
    outputs(1263) <= not a;
    outputs(1264) <= a xor b;
    outputs(1265) <= not a;
    outputs(1266) <= not a;
    outputs(1267) <= a and b;
    outputs(1268) <= not a;
    outputs(1269) <= b;
    outputs(1270) <= not (a xor b);
    outputs(1271) <= a;
    outputs(1272) <= b;
    outputs(1273) <= not b or a;
    outputs(1274) <= not a;
    outputs(1275) <= b and not a;
    outputs(1276) <= not a;
    outputs(1277) <= a xor b;
    outputs(1278) <= a;
    outputs(1279) <= not a or b;
    outputs(1280) <= not b;
    outputs(1281) <= not (a xor b);
    outputs(1282) <= a and not b;
    outputs(1283) <= a;
    outputs(1284) <= a xor b;
    outputs(1285) <= a xor b;
    outputs(1286) <= not (a or b);
    outputs(1287) <= not (a xor b);
    outputs(1288) <= a or b;
    outputs(1289) <= not (a or b);
    outputs(1290) <= not b;
    outputs(1291) <= b and not a;
    outputs(1292) <= a and b;
    outputs(1293) <= not (a and b);
    outputs(1294) <= not (a or b);
    outputs(1295) <= a;
    outputs(1296) <= not (a or b);
    outputs(1297) <= a;
    outputs(1298) <= b;
    outputs(1299) <= a xor b;
    outputs(1300) <= b and not a;
    outputs(1301) <= not (a or b);
    outputs(1302) <= b;
    outputs(1303) <= a and b;
    outputs(1304) <= not (a xor b);
    outputs(1305) <= a and not b;
    outputs(1306) <= not a;
    outputs(1307) <= b;
    outputs(1308) <= b;
    outputs(1309) <= b;
    outputs(1310) <= a xor b;
    outputs(1311) <= b and not a;
    outputs(1312) <= a xor b;
    outputs(1313) <= b and not a;
    outputs(1314) <= a xor b;
    outputs(1315) <= a and not b;
    outputs(1316) <= not (a xor b);
    outputs(1317) <= not b;
    outputs(1318) <= a xor b;
    outputs(1319) <= not (a xor b);
    outputs(1320) <= b;
    outputs(1321) <= a and b;
    outputs(1322) <= a and b;
    outputs(1323) <= a xor b;
    outputs(1324) <= b and not a;
    outputs(1325) <= a and b;
    outputs(1326) <= a xor b;
    outputs(1327) <= not (a xor b);
    outputs(1328) <= a;
    outputs(1329) <= a xor b;
    outputs(1330) <= a;
    outputs(1331) <= not b;
    outputs(1332) <= a;
    outputs(1333) <= b and not a;
    outputs(1334) <= not (a xor b);
    outputs(1335) <= not (a xor b);
    outputs(1336) <= not (a xor b);
    outputs(1337) <= not a;
    outputs(1338) <= a and b;
    outputs(1339) <= a and b;
    outputs(1340) <= b and not a;
    outputs(1341) <= b and not a;
    outputs(1342) <= a xor b;
    outputs(1343) <= not (a or b);
    outputs(1344) <= not (a xor b);
    outputs(1345) <= 1'b0;
    outputs(1346) <= not a;
    outputs(1347) <= not b;
    outputs(1348) <= a xor b;
    outputs(1349) <= a and not b;
    outputs(1350) <= b and not a;
    outputs(1351) <= not (a or b);
    outputs(1352) <= a and b;
    outputs(1353) <= not (a xor b);
    outputs(1354) <= b and not a;
    outputs(1355) <= a;
    outputs(1356) <= not (a or b);
    outputs(1357) <= a xor b;
    outputs(1358) <= a and b;
    outputs(1359) <= a;
    outputs(1360) <= a xor b;
    outputs(1361) <= a and not b;
    outputs(1362) <= not (a xor b);
    outputs(1363) <= b and not a;
    outputs(1364) <= a;
    outputs(1365) <= a xor b;
    outputs(1366) <= a xor b;
    outputs(1367) <= not a;
    outputs(1368) <= a and b;
    outputs(1369) <= not (a or b);
    outputs(1370) <= not b;
    outputs(1371) <= b and not a;
    outputs(1372) <= not b;
    outputs(1373) <= not b;
    outputs(1374) <= a;
    outputs(1375) <= a xor b;
    outputs(1376) <= b;
    outputs(1377) <= a and b;
    outputs(1378) <= a and b;
    outputs(1379) <= b;
    outputs(1380) <= a and not b;
    outputs(1381) <= a and b;
    outputs(1382) <= a and b;
    outputs(1383) <= a xor b;
    outputs(1384) <= a xor b;
    outputs(1385) <= not a;
    outputs(1386) <= a;
    outputs(1387) <= a and b;
    outputs(1388) <= not (a xor b);
    outputs(1389) <= not (a or b);
    outputs(1390) <= a or b;
    outputs(1391) <= not (a xor b);
    outputs(1392) <= a and not b;
    outputs(1393) <= b and not a;
    outputs(1394) <= b and not a;
    outputs(1395) <= a xor b;
    outputs(1396) <= b;
    outputs(1397) <= not a;
    outputs(1398) <= not (a or b);
    outputs(1399) <= a;
    outputs(1400) <= not (a or b);
    outputs(1401) <= a and b;
    outputs(1402) <= a xor b;
    outputs(1403) <= a and b;
    outputs(1404) <= not (a or b);
    outputs(1405) <= a;
    outputs(1406) <= a and not b;
    outputs(1407) <= a xor b;
    outputs(1408) <= not b;
    outputs(1409) <= b;
    outputs(1410) <= a xor b;
    outputs(1411) <= not a;
    outputs(1412) <= a and b;
    outputs(1413) <= b and not a;
    outputs(1414) <= b;
    outputs(1415) <= a xor b;
    outputs(1416) <= not (a or b);
    outputs(1417) <= not (a xor b);
    outputs(1418) <= not b;
    outputs(1419) <= not a;
    outputs(1420) <= not a;
    outputs(1421) <= b and not a;
    outputs(1422) <= a xor b;
    outputs(1423) <= not b;
    outputs(1424) <= not a;
    outputs(1425) <= b and not a;
    outputs(1426) <= a and not b;
    outputs(1427) <= not (a or b);
    outputs(1428) <= a and b;
    outputs(1429) <= not a;
    outputs(1430) <= a;
    outputs(1431) <= not a or b;
    outputs(1432) <= not (a or b);
    outputs(1433) <= b and not a;
    outputs(1434) <= b;
    outputs(1435) <= b and not a;
    outputs(1436) <= not (a or b);
    outputs(1437) <= b;
    outputs(1438) <= a xor b;
    outputs(1439) <= a xor b;
    outputs(1440) <= a and not b;
    outputs(1441) <= a xor b;
    outputs(1442) <= not (a or b);
    outputs(1443) <= a and not b;
    outputs(1444) <= not b;
    outputs(1445) <= b and not a;
    outputs(1446) <= b and not a;
    outputs(1447) <= not a;
    outputs(1448) <= a;
    outputs(1449) <= b;
    outputs(1450) <= a;
    outputs(1451) <= b;
    outputs(1452) <= a and b;
    outputs(1453) <= not b;
    outputs(1454) <= not (a xor b);
    outputs(1455) <= a xor b;
    outputs(1456) <= a and b;
    outputs(1457) <= not (a xor b);
    outputs(1458) <= a xor b;
    outputs(1459) <= a;
    outputs(1460) <= a and b;
    outputs(1461) <= b;
    outputs(1462) <= not (a xor b);
    outputs(1463) <= not b;
    outputs(1464) <= b and not a;
    outputs(1465) <= not (a xor b);
    outputs(1466) <= 1'b0;
    outputs(1467) <= b and not a;
    outputs(1468) <= not (a xor b);
    outputs(1469) <= not (a or b);
    outputs(1470) <= a xor b;
    outputs(1471) <= not (a or b);
    outputs(1472) <= not a;
    outputs(1473) <= not a;
    outputs(1474) <= a xor b;
    outputs(1475) <= a;
    outputs(1476) <= a xor b;
    outputs(1477) <= a and b;
    outputs(1478) <= a;
    outputs(1479) <= not (a or b);
    outputs(1480) <= a and not b;
    outputs(1481) <= a and not b;
    outputs(1482) <= not (a xor b);
    outputs(1483) <= a and not b;
    outputs(1484) <= b and not a;
    outputs(1485) <= not a;
    outputs(1486) <= not (a or b);
    outputs(1487) <= not (a xor b);
    outputs(1488) <= b;
    outputs(1489) <= not (a xor b);
    outputs(1490) <= not (a or b);
    outputs(1491) <= not b;
    outputs(1492) <= b and not a;
    outputs(1493) <= 1'b0;
    outputs(1494) <= a;
    outputs(1495) <= a and b;
    outputs(1496) <= b and not a;
    outputs(1497) <= a xor b;
    outputs(1498) <= 1'b0;
    outputs(1499) <= a xor b;
    outputs(1500) <= a xor b;
    outputs(1501) <= b and not a;
    outputs(1502) <= not (a or b);
    outputs(1503) <= not a;
    outputs(1504) <= not b;
    outputs(1505) <= not (a xor b);
    outputs(1506) <= a xor b;
    outputs(1507) <= not (a xor b);
    outputs(1508) <= b and not a;
    outputs(1509) <= 1'b0;
    outputs(1510) <= a and b;
    outputs(1511) <= not (a xor b);
    outputs(1512) <= not a;
    outputs(1513) <= not b;
    outputs(1514) <= b and not a;
    outputs(1515) <= a and not b;
    outputs(1516) <= a and not b;
    outputs(1517) <= a xor b;
    outputs(1518) <= not (a xor b);
    outputs(1519) <= not (a xor b);
    outputs(1520) <= not b;
    outputs(1521) <= b;
    outputs(1522) <= a;
    outputs(1523) <= a xor b;
    outputs(1524) <= a xor b;
    outputs(1525) <= a xor b;
    outputs(1526) <= b and not a;
    outputs(1527) <= b;
    outputs(1528) <= b and not a;
    outputs(1529) <= b;
    outputs(1530) <= a and b;
    outputs(1531) <= not (a xor b);
    outputs(1532) <= not b;
    outputs(1533) <= b and not a;
    outputs(1534) <= not (a xor b);
    outputs(1535) <= not (a xor b);
    outputs(1536) <= b and not a;
    outputs(1537) <= b;
    outputs(1538) <= not (a or b);
    outputs(1539) <= not (a xor b);
    outputs(1540) <= a and not b;
    outputs(1541) <= not b or a;
    outputs(1542) <= b;
    outputs(1543) <= a and not b;
    outputs(1544) <= not (a xor b);
    outputs(1545) <= b and not a;
    outputs(1546) <= not b;
    outputs(1547) <= a and not b;
    outputs(1548) <= b and not a;
    outputs(1549) <= b and not a;
    outputs(1550) <= a and b;
    outputs(1551) <= b and not a;
    outputs(1552) <= not (a xor b);
    outputs(1553) <= not (a xor b);
    outputs(1554) <= a and b;
    outputs(1555) <= a xor b;
    outputs(1556) <= b and not a;
    outputs(1557) <= a;
    outputs(1558) <= a xor b;
    outputs(1559) <= not b;
    outputs(1560) <= b and not a;
    outputs(1561) <= a and b;
    outputs(1562) <= b and not a;
    outputs(1563) <= b;
    outputs(1564) <= 1'b1;
    outputs(1565) <= not (a xor b);
    outputs(1566) <= not (a xor b);
    outputs(1567) <= a xor b;
    outputs(1568) <= b and not a;
    outputs(1569) <= not (a or b);
    outputs(1570) <= a and not b;
    outputs(1571) <= a xor b;
    outputs(1572) <= not (a xor b);
    outputs(1573) <= a and not b;
    outputs(1574) <= a and b;
    outputs(1575) <= b and not a;
    outputs(1576) <= a and b;
    outputs(1577) <= b and not a;
    outputs(1578) <= a and not b;
    outputs(1579) <= not (a or b);
    outputs(1580) <= not (a xor b);
    outputs(1581) <= a xor b;
    outputs(1582) <= a and b;
    outputs(1583) <= not b;
    outputs(1584) <= not a;
    outputs(1585) <= not (a xor b);
    outputs(1586) <= a and b;
    outputs(1587) <= not a;
    outputs(1588) <= a xor b;
    outputs(1589) <= not (a and b);
    outputs(1590) <= not a;
    outputs(1591) <= not a or b;
    outputs(1592) <= b and not a;
    outputs(1593) <= not a;
    outputs(1594) <= not (a xor b);
    outputs(1595) <= not b;
    outputs(1596) <= not (a xor b);
    outputs(1597) <= a and not b;
    outputs(1598) <= not b;
    outputs(1599) <= a and b;
    outputs(1600) <= b;
    outputs(1601) <= b and not a;
    outputs(1602) <= not a;
    outputs(1603) <= b and not a;
    outputs(1604) <= a xor b;
    outputs(1605) <= a and not b;
    outputs(1606) <= not (a xor b);
    outputs(1607) <= not (a xor b);
    outputs(1608) <= b and not a;
    outputs(1609) <= a xor b;
    outputs(1610) <= b and not a;
    outputs(1611) <= not (a or b);
    outputs(1612) <= b and not a;
    outputs(1613) <= b;
    outputs(1614) <= b;
    outputs(1615) <= b and not a;
    outputs(1616) <= not b;
    outputs(1617) <= a xor b;
    outputs(1618) <= b;
    outputs(1619) <= a and not b;
    outputs(1620) <= not a;
    outputs(1621) <= not a;
    outputs(1622) <= not a;
    outputs(1623) <= b;
    outputs(1624) <= a xor b;
    outputs(1625) <= a;
    outputs(1626) <= not b;
    outputs(1627) <= not (a or b);
    outputs(1628) <= a;
    outputs(1629) <= b and not a;
    outputs(1630) <= b and not a;
    outputs(1631) <= not (a xor b);
    outputs(1632) <= b;
    outputs(1633) <= a;
    outputs(1634) <= a and b;
    outputs(1635) <= a xor b;
    outputs(1636) <= b;
    outputs(1637) <= a xor b;
    outputs(1638) <= a xor b;
    outputs(1639) <= not a;
    outputs(1640) <= not (a or b);
    outputs(1641) <= b;
    outputs(1642) <= a and b;
    outputs(1643) <= not (a or b);
    outputs(1644) <= a and b;
    outputs(1645) <= not a;
    outputs(1646) <= not (a or b);
    outputs(1647) <= a xor b;
    outputs(1648) <= not (a or b);
    outputs(1649) <= a;
    outputs(1650) <= not (a or b);
    outputs(1651) <= not b;
    outputs(1652) <= a and b;
    outputs(1653) <= b and not a;
    outputs(1654) <= b;
    outputs(1655) <= 1'b0;
    outputs(1656) <= a xor b;
    outputs(1657) <= a;
    outputs(1658) <= a and b;
    outputs(1659) <= a and b;
    outputs(1660) <= a xor b;
    outputs(1661) <= b;
    outputs(1662) <= a and b;
    outputs(1663) <= not (a or b);
    outputs(1664) <= b;
    outputs(1665) <= not (a xor b);
    outputs(1666) <= b and not a;
    outputs(1667) <= not (a xor b);
    outputs(1668) <= a xor b;
    outputs(1669) <= not (a xor b);
    outputs(1670) <= a and b;
    outputs(1671) <= not b;
    outputs(1672) <= a and not b;
    outputs(1673) <= not b or a;
    outputs(1674) <= not (a xor b);
    outputs(1675) <= a xor b;
    outputs(1676) <= not (a or b);
    outputs(1677) <= not a;
    outputs(1678) <= not (a or b);
    outputs(1679) <= not a;
    outputs(1680) <= not a;
    outputs(1681) <= a and b;
    outputs(1682) <= a xor b;
    outputs(1683) <= b;
    outputs(1684) <= a xor b;
    outputs(1685) <= not a;
    outputs(1686) <= a;
    outputs(1687) <= not (a or b);
    outputs(1688) <= a and not b;
    outputs(1689) <= not a;
    outputs(1690) <= not (a or b);
    outputs(1691) <= not a;
    outputs(1692) <= b;
    outputs(1693) <= not (a or b);
    outputs(1694) <= a;
    outputs(1695) <= a and b;
    outputs(1696) <= not b;
    outputs(1697) <= b;
    outputs(1698) <= a and b;
    outputs(1699) <= a and b;
    outputs(1700) <= b and not a;
    outputs(1701) <= not b;
    outputs(1702) <= not a or b;
    outputs(1703) <= b and not a;
    outputs(1704) <= not b;
    outputs(1705) <= not (a xor b);
    outputs(1706) <= a xor b;
    outputs(1707) <= not a;
    outputs(1708) <= not (a xor b);
    outputs(1709) <= not a;
    outputs(1710) <= a and b;
    outputs(1711) <= not (a or b);
    outputs(1712) <= a;
    outputs(1713) <= a and b;
    outputs(1714) <= not b;
    outputs(1715) <= b and not a;
    outputs(1716) <= a and not b;
    outputs(1717) <= b and not a;
    outputs(1718) <= 1'b0;
    outputs(1719) <= not b or a;
    outputs(1720) <= not (a or b);
    outputs(1721) <= not (a xor b);
    outputs(1722) <= not (a or b);
    outputs(1723) <= a xor b;
    outputs(1724) <= 1'b0;
    outputs(1725) <= a xor b;
    outputs(1726) <= b and not a;
    outputs(1727) <= a and not b;
    outputs(1728) <= a xor b;
    outputs(1729) <= not (a or b);
    outputs(1730) <= not (a or b);
    outputs(1731) <= a and not b;
    outputs(1732) <= a and not b;
    outputs(1733) <= not (a xor b);
    outputs(1734) <= a and not b;
    outputs(1735) <= not (a or b);
    outputs(1736) <= not (a xor b);
    outputs(1737) <= b and not a;
    outputs(1738) <= b and not a;
    outputs(1739) <= a xor b;
    outputs(1740) <= 1'b0;
    outputs(1741) <= not (a xor b);
    outputs(1742) <= b and not a;
    outputs(1743) <= a xor b;
    outputs(1744) <= not b;
    outputs(1745) <= not (a xor b);
    outputs(1746) <= not b;
    outputs(1747) <= a and not b;
    outputs(1748) <= a and b;
    outputs(1749) <= b and not a;
    outputs(1750) <= a xor b;
    outputs(1751) <= not a;
    outputs(1752) <= not (a xor b);
    outputs(1753) <= a and not b;
    outputs(1754) <= not (a xor b);
    outputs(1755) <= 1'b0;
    outputs(1756) <= a and b;
    outputs(1757) <= a and not b;
    outputs(1758) <= a xor b;
    outputs(1759) <= b;
    outputs(1760) <= a and not b;
    outputs(1761) <= not b or a;
    outputs(1762) <= not b;
    outputs(1763) <= not b;
    outputs(1764) <= a xor b;
    outputs(1765) <= b and not a;
    outputs(1766) <= not (a xor b);
    outputs(1767) <= a xor b;
    outputs(1768) <= b;
    outputs(1769) <= a xor b;
    outputs(1770) <= not (a or b);
    outputs(1771) <= a and not b;
    outputs(1772) <= not b;
    outputs(1773) <= not (a xor b);
    outputs(1774) <= not (a xor b);
    outputs(1775) <= not a or b;
    outputs(1776) <= not (a xor b);
    outputs(1777) <= a xor b;
    outputs(1778) <= not a;
    outputs(1779) <= a;
    outputs(1780) <= not (a or b);
    outputs(1781) <= 1'b0;
    outputs(1782) <= not a;
    outputs(1783) <= not (a or b);
    outputs(1784) <= a;
    outputs(1785) <= not (a or b);
    outputs(1786) <= not (a xor b);
    outputs(1787) <= not (a xor b);
    outputs(1788) <= a;
    outputs(1789) <= a xor b;
    outputs(1790) <= b and not a;
    outputs(1791) <= not b;
    outputs(1792) <= a or b;
    outputs(1793) <= b and not a;
    outputs(1794) <= a and not b;
    outputs(1795) <= not (a xor b);
    outputs(1796) <= a and b;
    outputs(1797) <= a and b;
    outputs(1798) <= b and not a;
    outputs(1799) <= not b;
    outputs(1800) <= not (a xor b);
    outputs(1801) <= a xor b;
    outputs(1802) <= a xor b;
    outputs(1803) <= not a;
    outputs(1804) <= a xor b;
    outputs(1805) <= not (a or b);
    outputs(1806) <= a and not b;
    outputs(1807) <= a xor b;
    outputs(1808) <= a;
    outputs(1809) <= a xor b;
    outputs(1810) <= not (a xor b);
    outputs(1811) <= a xor b;
    outputs(1812) <= a xor b;
    outputs(1813) <= a and not b;
    outputs(1814) <= not (a or b);
    outputs(1815) <= not b;
    outputs(1816) <= a and b;
    outputs(1817) <= not a;
    outputs(1818) <= a and not b;
    outputs(1819) <= a xor b;
    outputs(1820) <= b and not a;
    outputs(1821) <= b and not a;
    outputs(1822) <= b;
    outputs(1823) <= not (a or b);
    outputs(1824) <= a and b;
    outputs(1825) <= not b;
    outputs(1826) <= a xor b;
    outputs(1827) <= not b;
    outputs(1828) <= not (a xor b);
    outputs(1829) <= b and not a;
    outputs(1830) <= b;
    outputs(1831) <= not (a or b);
    outputs(1832) <= not a;
    outputs(1833) <= not b;
    outputs(1834) <= a xor b;
    outputs(1835) <= a;
    outputs(1836) <= a and b;
    outputs(1837) <= a;
    outputs(1838) <= a or b;
    outputs(1839) <= not (a or b);
    outputs(1840) <= a;
    outputs(1841) <= not (a or b);
    outputs(1842) <= not (a or b);
    outputs(1843) <= a;
    outputs(1844) <= a and b;
    outputs(1845) <= a and b;
    outputs(1846) <= b and not a;
    outputs(1847) <= not (a or b);
    outputs(1848) <= b;
    outputs(1849) <= a and not b;
    outputs(1850) <= a xor b;
    outputs(1851) <= b and not a;
    outputs(1852) <= a;
    outputs(1853) <= not b;
    outputs(1854) <= not b;
    outputs(1855) <= not a;
    outputs(1856) <= a xor b;
    outputs(1857) <= not (a xor b);
    outputs(1858) <= a and b;
    outputs(1859) <= a xor b;
    outputs(1860) <= a xor b;
    outputs(1861) <= not b;
    outputs(1862) <= not b;
    outputs(1863) <= not a;
    outputs(1864) <= not a;
    outputs(1865) <= b;
    outputs(1866) <= not (a xor b);
    outputs(1867) <= a and b;
    outputs(1868) <= not b;
    outputs(1869) <= b and not a;
    outputs(1870) <= b and not a;
    outputs(1871) <= b;
    outputs(1872) <= b and not a;
    outputs(1873) <= a xor b;
    outputs(1874) <= a and not b;
    outputs(1875) <= not (a xor b);
    outputs(1876) <= not (a or b);
    outputs(1877) <= a and b;
    outputs(1878) <= not b;
    outputs(1879) <= a;
    outputs(1880) <= not (a or b);
    outputs(1881) <= not (a xor b);
    outputs(1882) <= not (a xor b);
    outputs(1883) <= b and not a;
    outputs(1884) <= b and not a;
    outputs(1885) <= a xor b;
    outputs(1886) <= a;
    outputs(1887) <= a xor b;
    outputs(1888) <= a and b;
    outputs(1889) <= a and b;
    outputs(1890) <= 1'b0;
    outputs(1891) <= not (a xor b);
    outputs(1892) <= not (a or b);
    outputs(1893) <= not (a or b);
    outputs(1894) <= a and not b;
    outputs(1895) <= a and not b;
    outputs(1896) <= a and not b;
    outputs(1897) <= b and not a;
    outputs(1898) <= not (a or b);
    outputs(1899) <= b and not a;
    outputs(1900) <= b and not a;
    outputs(1901) <= not a;
    outputs(1902) <= a;
    outputs(1903) <= not (a xor b);
    outputs(1904) <= b and not a;
    outputs(1905) <= a xor b;
    outputs(1906) <= not b;
    outputs(1907) <= a and not b;
    outputs(1908) <= a xor b;
    outputs(1909) <= not a;
    outputs(1910) <= not (a or b);
    outputs(1911) <= a xor b;
    outputs(1912) <= not a;
    outputs(1913) <= a;
    outputs(1914) <= a xor b;
    outputs(1915) <= not b;
    outputs(1916) <= not a;
    outputs(1917) <= b and not a;
    outputs(1918) <= b and not a;
    outputs(1919) <= not a;
    outputs(1920) <= not (a xor b);
    outputs(1921) <= not b;
    outputs(1922) <= not b;
    outputs(1923) <= not a or b;
    outputs(1924) <= not (a or b);
    outputs(1925) <= b and not a;
    outputs(1926) <= b and not a;
    outputs(1927) <= a and not b;
    outputs(1928) <= not (a xor b);
    outputs(1929) <= a;
    outputs(1930) <= 1'b0;
    outputs(1931) <= not a;
    outputs(1932) <= a and b;
    outputs(1933) <= a;
    outputs(1934) <= b and not a;
    outputs(1935) <= a and not b;
    outputs(1936) <= a and b;
    outputs(1937) <= a xor b;
    outputs(1938) <= not b;
    outputs(1939) <= a xor b;
    outputs(1940) <= a xor b;
    outputs(1941) <= not (a or b);
    outputs(1942) <= not (a or b);
    outputs(1943) <= not b;
    outputs(1944) <= a;
    outputs(1945) <= a and b;
    outputs(1946) <= b and not a;
    outputs(1947) <= a xor b;
    outputs(1948) <= not (a or b);
    outputs(1949) <= not a;
    outputs(1950) <= not a;
    outputs(1951) <= b and not a;
    outputs(1952) <= not (a or b);
    outputs(1953) <= a;
    outputs(1954) <= b and not a;
    outputs(1955) <= a and not b;
    outputs(1956) <= not (a or b);
    outputs(1957) <= a;
    outputs(1958) <= not (a or b);
    outputs(1959) <= not (a and b);
    outputs(1960) <= a xor b;
    outputs(1961) <= a and b;
    outputs(1962) <= a and b;
    outputs(1963) <= not (a xor b);
    outputs(1964) <= a or b;
    outputs(1965) <= not (a or b);
    outputs(1966) <= a and b;
    outputs(1967) <= a;
    outputs(1968) <= a xor b;
    outputs(1969) <= not a;
    outputs(1970) <= a and not b;
    outputs(1971) <= a and not b;
    outputs(1972) <= b;
    outputs(1973) <= not a;
    outputs(1974) <= b and not a;
    outputs(1975) <= b and not a;
    outputs(1976) <= b and not a;
    outputs(1977) <= a xor b;
    outputs(1978) <= 1'b0;
    outputs(1979) <= a and b;
    outputs(1980) <= b and not a;
    outputs(1981) <= not b;
    outputs(1982) <= a and not b;
    outputs(1983) <= b and not a;
    outputs(1984) <= not a;
    outputs(1985) <= not a;
    outputs(1986) <= a and b;
    outputs(1987) <= a and b;
    outputs(1988) <= a and b;
    outputs(1989) <= a and b;
    outputs(1990) <= a xor b;
    outputs(1991) <= a;
    outputs(1992) <= b and not a;
    outputs(1993) <= not (a or b);
    outputs(1994) <= not b;
    outputs(1995) <= a and b;
    outputs(1996) <= b;
    outputs(1997) <= a and b;
    outputs(1998) <= not (a and b);
    outputs(1999) <= not (a or b);
    outputs(2000) <= not a;
    outputs(2001) <= a and b;
    outputs(2002) <= not a;
    outputs(2003) <= not (a xor b);
    outputs(2004) <= a xor b;
    outputs(2005) <= not (a xor b);
    outputs(2006) <= a xor b;
    outputs(2007) <= not b;
    outputs(2008) <= b;
    outputs(2009) <= not (a or b);
    outputs(2010) <= not (a xor b);
    outputs(2011) <= b and not a;
    outputs(2012) <= a and not b;
    outputs(2013) <= not (a xor b);
    outputs(2014) <= not (a xor b);
    outputs(2015) <= b and not a;
    outputs(2016) <= not a;
    outputs(2017) <= not b;
    outputs(2018) <= not a;
    outputs(2019) <= not (a xor b);
    outputs(2020) <= a and b;
    outputs(2021) <= a and b;
    outputs(2022) <= a;
    outputs(2023) <= a and b;
    outputs(2024) <= 1'b0;
    outputs(2025) <= a;
    outputs(2026) <= a xor b;
    outputs(2027) <= not (a or b);
    outputs(2028) <= not b;
    outputs(2029) <= a and b;
    outputs(2030) <= a xor b;
    outputs(2031) <= a xor b;
    outputs(2032) <= not (a or b);
    outputs(2033) <= not (a and b);
    outputs(2034) <= not b;
    outputs(2035) <= not (a or b);
    outputs(2036) <= b;
    outputs(2037) <= not (a or b);
    outputs(2038) <= a and b;
    outputs(2039) <= a and b;
    outputs(2040) <= not b;
    outputs(2041) <= a and not b;
    outputs(2042) <= a and not b;
    outputs(2043) <= a and b;
    outputs(2044) <= a;
    outputs(2045) <= a xor b;
    outputs(2046) <= a xor b;
    outputs(2047) <= b and not a;
    outputs(2048) <= a and not b;
    outputs(2049) <= not (a or b);
    outputs(2050) <= b;
    outputs(2051) <= not a or b;
    outputs(2052) <= a xor b;
    outputs(2053) <= not a;
    outputs(2054) <= a;
    outputs(2055) <= not a;
    outputs(2056) <= not (a xor b);
    outputs(2057) <= a and b;
    outputs(2058) <= a xor b;
    outputs(2059) <= a and b;
    outputs(2060) <= not (a or b);
    outputs(2061) <= not a;
    outputs(2062) <= a and b;
    outputs(2063) <= a and b;
    outputs(2064) <= a;
    outputs(2065) <= a;
    outputs(2066) <= a;
    outputs(2067) <= a;
    outputs(2068) <= not (a xor b);
    outputs(2069) <= not a;
    outputs(2070) <= a xor b;
    outputs(2071) <= a;
    outputs(2072) <= a xor b;
    outputs(2073) <= not (a xor b);
    outputs(2074) <= a and not b;
    outputs(2075) <= not a or b;
    outputs(2076) <= b and not a;
    outputs(2077) <= not (a xor b);
    outputs(2078) <= a and b;
    outputs(2079) <= b;
    outputs(2080) <= not a;
    outputs(2081) <= not b;
    outputs(2082) <= not a or b;
    outputs(2083) <= a xor b;
    outputs(2084) <= a;
    outputs(2085) <= a and b;
    outputs(2086) <= a xor b;
    outputs(2087) <= not b;
    outputs(2088) <= a xor b;
    outputs(2089) <= not a;
    outputs(2090) <= b and not a;
    outputs(2091) <= not a;
    outputs(2092) <= not (a or b);
    outputs(2093) <= a and not b;
    outputs(2094) <= a;
    outputs(2095) <= not a;
    outputs(2096) <= b;
    outputs(2097) <= b and not a;
    outputs(2098) <= not a;
    outputs(2099) <= a xor b;
    outputs(2100) <= a xor b;
    outputs(2101) <= a xor b;
    outputs(2102) <= a and b;
    outputs(2103) <= a;
    outputs(2104) <= not (a or b);
    outputs(2105) <= a;
    outputs(2106) <= a and b;
    outputs(2107) <= not (a or b);
    outputs(2108) <= a and not b;
    outputs(2109) <= not (a xor b);
    outputs(2110) <= not (a or b);
    outputs(2111) <= not a;
    outputs(2112) <= not (a xor b);
    outputs(2113) <= a and not b;
    outputs(2114) <= a xor b;
    outputs(2115) <= b;
    outputs(2116) <= a and not b;
    outputs(2117) <= a and not b;
    outputs(2118) <= not a;
    outputs(2119) <= a and not b;
    outputs(2120) <= not (a xor b);
    outputs(2121) <= a;
    outputs(2122) <= not (a or b);
    outputs(2123) <= a and b;
    outputs(2124) <= b and not a;
    outputs(2125) <= not (a xor b);
    outputs(2126) <= not (a xor b);
    outputs(2127) <= b;
    outputs(2128) <= a and b;
    outputs(2129) <= a;
    outputs(2130) <= b and not a;
    outputs(2131) <= b and not a;
    outputs(2132) <= not a;
    outputs(2133) <= not (a xor b);
    outputs(2134) <= a xor b;
    outputs(2135) <= a and b;
    outputs(2136) <= a and b;
    outputs(2137) <= not (a xor b);
    outputs(2138) <= b and not a;
    outputs(2139) <= a and b;
    outputs(2140) <= not (a xor b);
    outputs(2141) <= a and b;
    outputs(2142) <= a xor b;
    outputs(2143) <= a and b;
    outputs(2144) <= not (a xor b);
    outputs(2145) <= not (a xor b);
    outputs(2146) <= a and b;
    outputs(2147) <= not b;
    outputs(2148) <= a;
    outputs(2149) <= not b;
    outputs(2150) <= not (a xor b);
    outputs(2151) <= b;
    outputs(2152) <= b;
    outputs(2153) <= not (a xor b);
    outputs(2154) <= a xor b;
    outputs(2155) <= a and not b;
    outputs(2156) <= not b or a;
    outputs(2157) <= a and not b;
    outputs(2158) <= b;
    outputs(2159) <= not a;
    outputs(2160) <= not (a or b);
    outputs(2161) <= not (a xor b);
    outputs(2162) <= a and b;
    outputs(2163) <= a and b;
    outputs(2164) <= a and not b;
    outputs(2165) <= a and not b;
    outputs(2166) <= b and not a;
    outputs(2167) <= a xor b;
    outputs(2168) <= not (a xor b);
    outputs(2169) <= b;
    outputs(2170) <= a and b;
    outputs(2171) <= b and not a;
    outputs(2172) <= not b;
    outputs(2173) <= not a;
    outputs(2174) <= not a;
    outputs(2175) <= a;
    outputs(2176) <= a and b;
    outputs(2177) <= b and not a;
    outputs(2178) <= b;
    outputs(2179) <= a and not b;
    outputs(2180) <= a and not b;
    outputs(2181) <= not (a and b);
    outputs(2182) <= not (a xor b);
    outputs(2183) <= not (a or b);
    outputs(2184) <= a;
    outputs(2185) <= a;
    outputs(2186) <= not b or a;
    outputs(2187) <= not (a or b);
    outputs(2188) <= not a;
    outputs(2189) <= a and not b;
    outputs(2190) <= not (a xor b);
    outputs(2191) <= a and b;
    outputs(2192) <= a xor b;
    outputs(2193) <= a and b;
    outputs(2194) <= b;
    outputs(2195) <= not (a or b);
    outputs(2196) <= a and not b;
    outputs(2197) <= a and b;
    outputs(2198) <= not a;
    outputs(2199) <= a xor b;
    outputs(2200) <= a or b;
    outputs(2201) <= a and not b;
    outputs(2202) <= not b;
    outputs(2203) <= not (a or b);
    outputs(2204) <= a;
    outputs(2205) <= b and not a;
    outputs(2206) <= 1'b0;
    outputs(2207) <= b and not a;
    outputs(2208) <= not (a xor b);
    outputs(2209) <= a;
    outputs(2210) <= not (a xor b);
    outputs(2211) <= not (a xor b);
    outputs(2212) <= not a;
    outputs(2213) <= not (a or b);
    outputs(2214) <= a and not b;
    outputs(2215) <= b and not a;
    outputs(2216) <= a and b;
    outputs(2217) <= 1'b0;
    outputs(2218) <= a and not b;
    outputs(2219) <= a and b;
    outputs(2220) <= b and not a;
    outputs(2221) <= not (a or b);
    outputs(2222) <= a and not b;
    outputs(2223) <= not a;
    outputs(2224) <= a and not b;
    outputs(2225) <= not (a xor b);
    outputs(2226) <= not b;
    outputs(2227) <= 1'b0;
    outputs(2228) <= a xor b;
    outputs(2229) <= a and not b;
    outputs(2230) <= b and not a;
    outputs(2231) <= not (a xor b);
    outputs(2232) <= not (a or b);
    outputs(2233) <= a and not b;
    outputs(2234) <= a xor b;
    outputs(2235) <= a and not b;
    outputs(2236) <= a xor b;
    outputs(2237) <= a and b;
    outputs(2238) <= 1'b0;
    outputs(2239) <= a xor b;
    outputs(2240) <= not (a xor b);
    outputs(2241) <= 1'b0;
    outputs(2242) <= not (a or b);
    outputs(2243) <= not (a xor b);
    outputs(2244) <= a and b;
    outputs(2245) <= b;
    outputs(2246) <= a and not b;
    outputs(2247) <= not b;
    outputs(2248) <= a and not b;
    outputs(2249) <= b and not a;
    outputs(2250) <= b and not a;
    outputs(2251) <= a xor b;
    outputs(2252) <= a and b;
    outputs(2253) <= a and b;
    outputs(2254) <= not b;
    outputs(2255) <= not b;
    outputs(2256) <= a and not b;
    outputs(2257) <= b and not a;
    outputs(2258) <= a and b;
    outputs(2259) <= not (a xor b);
    outputs(2260) <= not (a or b);
    outputs(2261) <= a and not b;
    outputs(2262) <= b;
    outputs(2263) <= a xor b;
    outputs(2264) <= b;
    outputs(2265) <= a xor b;
    outputs(2266) <= not a;
    outputs(2267) <= not b;
    outputs(2268) <= a and not b;
    outputs(2269) <= not a;
    outputs(2270) <= a and b;
    outputs(2271) <= a and not b;
    outputs(2272) <= a and b;
    outputs(2273) <= not (a or b);
    outputs(2274) <= b and not a;
    outputs(2275) <= b and not a;
    outputs(2276) <= not a;
    outputs(2277) <= b;
    outputs(2278) <= b and not a;
    outputs(2279) <= not b;
    outputs(2280) <= not (a xor b);
    outputs(2281) <= b;
    outputs(2282) <= b and not a;
    outputs(2283) <= not (a xor b);
    outputs(2284) <= a xor b;
    outputs(2285) <= a and not b;
    outputs(2286) <= a and b;
    outputs(2287) <= b and not a;
    outputs(2288) <= a and b;
    outputs(2289) <= a and not b;
    outputs(2290) <= not a;
    outputs(2291) <= b and not a;
    outputs(2292) <= a;
    outputs(2293) <= not (a or b);
    outputs(2294) <= not (a xor b);
    outputs(2295) <= a and not b;
    outputs(2296) <= not a;
    outputs(2297) <= not (a xor b);
    outputs(2298) <= b and not a;
    outputs(2299) <= not (a or b);
    outputs(2300) <= not (a xor b);
    outputs(2301) <= a and b;
    outputs(2302) <= a;
    outputs(2303) <= a and b;
    outputs(2304) <= not b;
    outputs(2305) <= not (a xor b);
    outputs(2306) <= not b;
    outputs(2307) <= a and b;
    outputs(2308) <= a and b;
    outputs(2309) <= not a;
    outputs(2310) <= not (a xor b);
    outputs(2311) <= not (a or b);
    outputs(2312) <= b;
    outputs(2313) <= b;
    outputs(2314) <= a;
    outputs(2315) <= a and b;
    outputs(2316) <= b;
    outputs(2317) <= not a;
    outputs(2318) <= a and not b;
    outputs(2319) <= 1'b0;
    outputs(2320) <= b;
    outputs(2321) <= b and not a;
    outputs(2322) <= not (a xor b);
    outputs(2323) <= b and not a;
    outputs(2324) <= not b;
    outputs(2325) <= not b;
    outputs(2326) <= a xor b;
    outputs(2327) <= a and b;
    outputs(2328) <= a and b;
    outputs(2329) <= a and not b;
    outputs(2330) <= b;
    outputs(2331) <= a and not b;
    outputs(2332) <= a xor b;
    outputs(2333) <= a;
    outputs(2334) <= b;
    outputs(2335) <= not (a xor b);
    outputs(2336) <= a and b;
    outputs(2337) <= a and not b;
    outputs(2338) <= a and b;
    outputs(2339) <= not a;
    outputs(2340) <= b and not a;
    outputs(2341) <= b and not a;
    outputs(2342) <= not (a xor b);
    outputs(2343) <= not (a or b);
    outputs(2344) <= b;
    outputs(2345) <= not (a or b);
    outputs(2346) <= not (a xor b);
    outputs(2347) <= b and not a;
    outputs(2348) <= b and not a;
    outputs(2349) <= not (a xor b);
    outputs(2350) <= not b;
    outputs(2351) <= not (a or b);
    outputs(2352) <= not b;
    outputs(2353) <= not (a xor b);
    outputs(2354) <= a;
    outputs(2355) <= a and not b;
    outputs(2356) <= not (a xor b);
    outputs(2357) <= a and b;
    outputs(2358) <= a;
    outputs(2359) <= a;
    outputs(2360) <= a and not b;
    outputs(2361) <= a;
    outputs(2362) <= a xor b;
    outputs(2363) <= b;
    outputs(2364) <= not (a or b);
    outputs(2365) <= not (a or b);
    outputs(2366) <= not a;
    outputs(2367) <= a or b;
    outputs(2368) <= a xor b;
    outputs(2369) <= a and b;
    outputs(2370) <= a;
    outputs(2371) <= a xor b;
    outputs(2372) <= not (a xor b);
    outputs(2373) <= b and not a;
    outputs(2374) <= a xor b;
    outputs(2375) <= a xor b;
    outputs(2376) <= a and b;
    outputs(2377) <= b and not a;
    outputs(2378) <= b and not a;
    outputs(2379) <= not b;
    outputs(2380) <= not (a or b);
    outputs(2381) <= a and not b;
    outputs(2382) <= not b;
    outputs(2383) <= not (a xor b);
    outputs(2384) <= not a;
    outputs(2385) <= not (a or b);
    outputs(2386) <= b;
    outputs(2387) <= a;
    outputs(2388) <= a and b;
    outputs(2389) <= not (a or b);
    outputs(2390) <= a and not b;
    outputs(2391) <= not (a or b);
    outputs(2392) <= a and not b;
    outputs(2393) <= not (a or b);
    outputs(2394) <= a and b;
    outputs(2395) <= a and not b;
    outputs(2396) <= a and not b;
    outputs(2397) <= a xor b;
    outputs(2398) <= a;
    outputs(2399) <= not a;
    outputs(2400) <= b and not a;
    outputs(2401) <= not (a xor b);
    outputs(2402) <= a;
    outputs(2403) <= b and not a;
    outputs(2404) <= a and b;
    outputs(2405) <= not (a xor b);
    outputs(2406) <= a xor b;
    outputs(2407) <= a and not b;
    outputs(2408) <= b and not a;
    outputs(2409) <= a and b;
    outputs(2410) <= b and not a;
    outputs(2411) <= b;
    outputs(2412) <= a xor b;
    outputs(2413) <= a and b;
    outputs(2414) <= not (a or b);
    outputs(2415) <= a xor b;
    outputs(2416) <= not (a or b);
    outputs(2417) <= b;
    outputs(2418) <= b;
    outputs(2419) <= b and not a;
    outputs(2420) <= not a;
    outputs(2421) <= a;
    outputs(2422) <= b;
    outputs(2423) <= a;
    outputs(2424) <= a and b;
    outputs(2425) <= a xor b;
    outputs(2426) <= a and not b;
    outputs(2427) <= b and not a;
    outputs(2428) <= a xor b;
    outputs(2429) <= not (a or b);
    outputs(2430) <= not a;
    outputs(2431) <= not (a xor b);
    outputs(2432) <= not (a xor b);
    outputs(2433) <= not b;
    outputs(2434) <= a and b;
    outputs(2435) <= not b;
    outputs(2436) <= a and not b;
    outputs(2437) <= a and b;
    outputs(2438) <= not (a xor b);
    outputs(2439) <= not (a xor b);
    outputs(2440) <= b and not a;
    outputs(2441) <= a xor b;
    outputs(2442) <= not (a or b);
    outputs(2443) <= b;
    outputs(2444) <= a and not b;
    outputs(2445) <= b and not a;
    outputs(2446) <= a and b;
    outputs(2447) <= b and not a;
    outputs(2448) <= b and not a;
    outputs(2449) <= a xor b;
    outputs(2450) <= not b;
    outputs(2451) <= b;
    outputs(2452) <= not (a or b);
    outputs(2453) <= a and not b;
    outputs(2454) <= 1'b0;
    outputs(2455) <= not (a or b);
    outputs(2456) <= a and not b;
    outputs(2457) <= a and b;
    outputs(2458) <= not (a xor b);
    outputs(2459) <= a xor b;
    outputs(2460) <= not a;
    outputs(2461) <= b and not a;
    outputs(2462) <= a xor b;
    outputs(2463) <= not (a or b);
    outputs(2464) <= not (a xor b);
    outputs(2465) <= b and not a;
    outputs(2466) <= b and not a;
    outputs(2467) <= not (a or b);
    outputs(2468) <= not (a xor b);
    outputs(2469) <= a and b;
    outputs(2470) <= b;
    outputs(2471) <= 1'b0;
    outputs(2472) <= a and b;
    outputs(2473) <= not (a or b);
    outputs(2474) <= a xor b;
    outputs(2475) <= not (a xor b);
    outputs(2476) <= not a;
    outputs(2477) <= not (a or b);
    outputs(2478) <= a and not b;
    outputs(2479) <= not (a xor b);
    outputs(2480) <= a and b;
    outputs(2481) <= not (a or b);
    outputs(2482) <= not (a xor b);
    outputs(2483) <= a and not b;
    outputs(2484) <= a xor b;
    outputs(2485) <= b and not a;
    outputs(2486) <= not (a xor b);
    outputs(2487) <= a xor b;
    outputs(2488) <= not b;
    outputs(2489) <= not (a xor b);
    outputs(2490) <= b;
    outputs(2491) <= b and not a;
    outputs(2492) <= not (a xor b);
    outputs(2493) <= a xor b;
    outputs(2494) <= not (a or b);
    outputs(2495) <= not (a or b);
    outputs(2496) <= b and not a;
    outputs(2497) <= b;
    outputs(2498) <= a;
    outputs(2499) <= a xor b;
    outputs(2500) <= b;
    outputs(2501) <= not a;
    outputs(2502) <= not a;
    outputs(2503) <= a and b;
    outputs(2504) <= a and b;
    outputs(2505) <= not (a xor b);
    outputs(2506) <= a;
    outputs(2507) <= b and not a;
    outputs(2508) <= a xor b;
    outputs(2509) <= not (a or b);
    outputs(2510) <= b;
    outputs(2511) <= a and not b;
    outputs(2512) <= a and not b;
    outputs(2513) <= not (a xor b);
    outputs(2514) <= b;
    outputs(2515) <= not (a xor b);
    outputs(2516) <= b and not a;
    outputs(2517) <= not a;
    outputs(2518) <= not (a xor b);
    outputs(2519) <= a;
    outputs(2520) <= not (a or b);
    outputs(2521) <= a xor b;
    outputs(2522) <= not (a or b);
    outputs(2523) <= a and not b;
    outputs(2524) <= b and not a;
    outputs(2525) <= a xor b;
    outputs(2526) <= not (a xor b);
    outputs(2527) <= not a;
    outputs(2528) <= b and not a;
    outputs(2529) <= a and b;
    outputs(2530) <= b and not a;
    outputs(2531) <= b;
    outputs(2532) <= a xor b;
    outputs(2533) <= b;
    outputs(2534) <= not a;
    outputs(2535) <= a;
    outputs(2536) <= not b;
    outputs(2537) <= not b;
    outputs(2538) <= b and not a;
    outputs(2539) <= not (a or b);
    outputs(2540) <= not b;
    outputs(2541) <= a and not b;
    outputs(2542) <= a and not b;
    outputs(2543) <= b;
    outputs(2544) <= a and b;
    outputs(2545) <= not b;
    outputs(2546) <= a and b;
    outputs(2547) <= a and b;
    outputs(2548) <= 1'b0;
    outputs(2549) <= a and not b;
    outputs(2550) <= b;
    outputs(2551) <= not (a xor b);
    outputs(2552) <= a or b;
    outputs(2553) <= a and b;
    outputs(2554) <= not (a xor b);
    outputs(2555) <= a;
    outputs(2556) <= a and not b;
    outputs(2557) <= not a or b;
    outputs(2558) <= a and b;
    outputs(2559) <= not (a or b);
    outputs(2560) <= a;
    outputs(2561) <= not (a and b);
    outputs(2562) <= not (a xor b);
    outputs(2563) <= not a or b;
    outputs(2564) <= a and not b;
    outputs(2565) <= b and not a;
    outputs(2566) <= b;
    outputs(2567) <= a and not b;
    outputs(2568) <= not (a and b);
    outputs(2569) <= a or b;
    outputs(2570) <= a xor b;
    outputs(2571) <= not a;
    outputs(2572) <= b;
    outputs(2573) <= b and not a;
    outputs(2574) <= a;
    outputs(2575) <= not b;
    outputs(2576) <= a or b;
    outputs(2577) <= a;
    outputs(2578) <= not a;
    outputs(2579) <= not (a and b);
    outputs(2580) <= not b or a;
    outputs(2581) <= not (a xor b);
    outputs(2582) <= not a;
    outputs(2583) <= not (a xor b);
    outputs(2584) <= b and not a;
    outputs(2585) <= a;
    outputs(2586) <= a or b;
    outputs(2587) <= a xor b;
    outputs(2588) <= a;
    outputs(2589) <= a;
    outputs(2590) <= a and not b;
    outputs(2591) <= a xor b;
    outputs(2592) <= b;
    outputs(2593) <= b;
    outputs(2594) <= not (a and b);
    outputs(2595) <= not a;
    outputs(2596) <= a xor b;
    outputs(2597) <= not (a or b);
    outputs(2598) <= not b;
    outputs(2599) <= not (a and b);
    outputs(2600) <= not (a xor b);
    outputs(2601) <= b and not a;
    outputs(2602) <= a xor b;
    outputs(2603) <= b and not a;
    outputs(2604) <= not a or b;
    outputs(2605) <= a or b;
    outputs(2606) <= a xor b;
    outputs(2607) <= not (a xor b);
    outputs(2608) <= a;
    outputs(2609) <= a;
    outputs(2610) <= not a;
    outputs(2611) <= not (a or b);
    outputs(2612) <= not a;
    outputs(2613) <= a xor b;
    outputs(2614) <= a xor b;
    outputs(2615) <= 1'b1;
    outputs(2616) <= not (a and b);
    outputs(2617) <= not (a xor b);
    outputs(2618) <= not (a xor b);
    outputs(2619) <= b;
    outputs(2620) <= not (a xor b);
    outputs(2621) <= not (a or b);
    outputs(2622) <= not a;
    outputs(2623) <= a xor b;
    outputs(2624) <= a xor b;
    outputs(2625) <= not (a xor b);
    outputs(2626) <= not a or b;
    outputs(2627) <= not a;
    outputs(2628) <= b;
    outputs(2629) <= not (a xor b);
    outputs(2630) <= not b or a;
    outputs(2631) <= a or b;
    outputs(2632) <= b;
    outputs(2633) <= not b or a;
    outputs(2634) <= not a or b;
    outputs(2635) <= a xor b;
    outputs(2636) <= not b;
    outputs(2637) <= not (a or b);
    outputs(2638) <= b;
    outputs(2639) <= not a or b;
    outputs(2640) <= not b or a;
    outputs(2641) <= b;
    outputs(2642) <= not a;
    outputs(2643) <= not (a xor b);
    outputs(2644) <= not a or b;
    outputs(2645) <= not b;
    outputs(2646) <= a xor b;
    outputs(2647) <= not (a and b);
    outputs(2648) <= a;
    outputs(2649) <= b;
    outputs(2650) <= a xor b;
    outputs(2651) <= not (a xor b);
    outputs(2652) <= a xor b;
    outputs(2653) <= not b;
    outputs(2654) <= not a or b;
    outputs(2655) <= not (a xor b);
    outputs(2656) <= not b;
    outputs(2657) <= not b or a;
    outputs(2658) <= a and not b;
    outputs(2659) <= a and not b;
    outputs(2660) <= a or b;
    outputs(2661) <= a xor b;
    outputs(2662) <= not a;
    outputs(2663) <= not b or a;
    outputs(2664) <= not a;
    outputs(2665) <= not (a xor b);
    outputs(2666) <= a or b;
    outputs(2667) <= not (a xor b);
    outputs(2668) <= not (a xor b);
    outputs(2669) <= a and b;
    outputs(2670) <= not b or a;
    outputs(2671) <= not a or b;
    outputs(2672) <= a or b;
    outputs(2673) <= not b;
    outputs(2674) <= a xor b;
    outputs(2675) <= b;
    outputs(2676) <= a;
    outputs(2677) <= not a;
    outputs(2678) <= a xor b;
    outputs(2679) <= 1'b1;
    outputs(2680) <= a;
    outputs(2681) <= b and not a;
    outputs(2682) <= not b;
    outputs(2683) <= b;
    outputs(2684) <= not (a xor b);
    outputs(2685) <= not a or b;
    outputs(2686) <= not b;
    outputs(2687) <= b;
    outputs(2688) <= not (a xor b);
    outputs(2689) <= a and not b;
    outputs(2690) <= not (a xor b);
    outputs(2691) <= not b;
    outputs(2692) <= a xor b;
    outputs(2693) <= b;
    outputs(2694) <= not (a or b);
    outputs(2695) <= not (a and b);
    outputs(2696) <= b;
    outputs(2697) <= b;
    outputs(2698) <= not b or a;
    outputs(2699) <= not (a xor b);
    outputs(2700) <= not (a or b);
    outputs(2701) <= not b;
    outputs(2702) <= not b or a;
    outputs(2703) <= a and b;
    outputs(2704) <= not b or a;
    outputs(2705) <= b;
    outputs(2706) <= a xor b;
    outputs(2707) <= not a;
    outputs(2708) <= not (a xor b);
    outputs(2709) <= a;
    outputs(2710) <= not (a or b);
    outputs(2711) <= a;
    outputs(2712) <= not b;
    outputs(2713) <= a;
    outputs(2714) <= not a;
    outputs(2715) <= b;
    outputs(2716) <= not (a and b);
    outputs(2717) <= b and not a;
    outputs(2718) <= not a or b;
    outputs(2719) <= a or b;
    outputs(2720) <= not (a and b);
    outputs(2721) <= a or b;
    outputs(2722) <= not a;
    outputs(2723) <= b;
    outputs(2724) <= not a or b;
    outputs(2725) <= not (a xor b);
    outputs(2726) <= b and not a;
    outputs(2727) <= a and b;
    outputs(2728) <= not b or a;
    outputs(2729) <= a or b;
    outputs(2730) <= b;
    outputs(2731) <= not b;
    outputs(2732) <= not a or b;
    outputs(2733) <= b and not a;
    outputs(2734) <= a xor b;
    outputs(2735) <= not b or a;
    outputs(2736) <= not (a xor b);
    outputs(2737) <= a and b;
    outputs(2738) <= a or b;
    outputs(2739) <= a;
    outputs(2740) <= not b or a;
    outputs(2741) <= not (a and b);
    outputs(2742) <= a and not b;
    outputs(2743) <= not (a and b);
    outputs(2744) <= b;
    outputs(2745) <= not a or b;
    outputs(2746) <= not b;
    outputs(2747) <= a and b;
    outputs(2748) <= not (a xor b);
    outputs(2749) <= a or b;
    outputs(2750) <= not b;
    outputs(2751) <= not (a xor b);
    outputs(2752) <= not b or a;
    outputs(2753) <= a;
    outputs(2754) <= not a or b;
    outputs(2755) <= a xor b;
    outputs(2756) <= not a;
    outputs(2757) <= b;
    outputs(2758) <= a and b;
    outputs(2759) <= a;
    outputs(2760) <= not (a and b);
    outputs(2761) <= a;
    outputs(2762) <= a and b;
    outputs(2763) <= not (a xor b);
    outputs(2764) <= b;
    outputs(2765) <= not (a or b);
    outputs(2766) <= not a;
    outputs(2767) <= not (a xor b);
    outputs(2768) <= not a;
    outputs(2769) <= a;
    outputs(2770) <= a xor b;
    outputs(2771) <= not b;
    outputs(2772) <= a;
    outputs(2773) <= not a;
    outputs(2774) <= a;
    outputs(2775) <= b;
    outputs(2776) <= a and not b;
    outputs(2777) <= a xor b;
    outputs(2778) <= not a or b;
    outputs(2779) <= not (a and b);
    outputs(2780) <= not (a xor b);
    outputs(2781) <= a;
    outputs(2782) <= not (a or b);
    outputs(2783) <= a xor b;
    outputs(2784) <= not a;
    outputs(2785) <= not (a xor b);
    outputs(2786) <= not b;
    outputs(2787) <= not (a and b);
    outputs(2788) <= not (a xor b);
    outputs(2789) <= not (a or b);
    outputs(2790) <= not b or a;
    outputs(2791) <= a;
    outputs(2792) <= not b;
    outputs(2793) <= a xor b;
    outputs(2794) <= a;
    outputs(2795) <= b;
    outputs(2796) <= a and b;
    outputs(2797) <= a;
    outputs(2798) <= a xor b;
    outputs(2799) <= a;
    outputs(2800) <= not (a and b);
    outputs(2801) <= b and not a;
    outputs(2802) <= not a or b;
    outputs(2803) <= a;
    outputs(2804) <= b and not a;
    outputs(2805) <= not a or b;
    outputs(2806) <= not (a xor b);
    outputs(2807) <= not (a xor b);
    outputs(2808) <= not (a xor b);
    outputs(2809) <= a xor b;
    outputs(2810) <= not (a and b);
    outputs(2811) <= b;
    outputs(2812) <= a;
    outputs(2813) <= not (a xor b);
    outputs(2814) <= a xor b;
    outputs(2815) <= a or b;
    outputs(2816) <= not b or a;
    outputs(2817) <= not b;
    outputs(2818) <= not a;
    outputs(2819) <= not a or b;
    outputs(2820) <= a or b;
    outputs(2821) <= not (a xor b);
    outputs(2822) <= b and not a;
    outputs(2823) <= a or b;
    outputs(2824) <= not a;
    outputs(2825) <= a and not b;
    outputs(2826) <= a and b;
    outputs(2827) <= b;
    outputs(2828) <= a or b;
    outputs(2829) <= a or b;
    outputs(2830) <= b;
    outputs(2831) <= not a;
    outputs(2832) <= b;
    outputs(2833) <= not b;
    outputs(2834) <= not b;
    outputs(2835) <= not b;
    outputs(2836) <= a;
    outputs(2837) <= a or b;
    outputs(2838) <= not (a xor b);
    outputs(2839) <= not a;
    outputs(2840) <= a xor b;
    outputs(2841) <= b;
    outputs(2842) <= a or b;
    outputs(2843) <= not b or a;
    outputs(2844) <= not (a xor b);
    outputs(2845) <= not b;
    outputs(2846) <= not (a xor b);
    outputs(2847) <= a xor b;
    outputs(2848) <= a xor b;
    outputs(2849) <= a or b;
    outputs(2850) <= not a;
    outputs(2851) <= not a or b;
    outputs(2852) <= not b or a;
    outputs(2853) <= a or b;
    outputs(2854) <= b;
    outputs(2855) <= a or b;
    outputs(2856) <= a and not b;
    outputs(2857) <= a xor b;
    outputs(2858) <= a xor b;
    outputs(2859) <= a or b;
    outputs(2860) <= a xor b;
    outputs(2861) <= not a or b;
    outputs(2862) <= not a or b;
    outputs(2863) <= not b;
    outputs(2864) <= a xor b;
    outputs(2865) <= a and not b;
    outputs(2866) <= not (a and b);
    outputs(2867) <= not a;
    outputs(2868) <= a and b;
    outputs(2869) <= not b;
    outputs(2870) <= b;
    outputs(2871) <= not b or a;
    outputs(2872) <= not (a xor b);
    outputs(2873) <= not (a xor b);
    outputs(2874) <= not (a xor b);
    outputs(2875) <= a xor b;
    outputs(2876) <= a and not b;
    outputs(2877) <= a xor b;
    outputs(2878) <= 1'b1;
    outputs(2879) <= not (a xor b);
    outputs(2880) <= a xor b;
    outputs(2881) <= a;
    outputs(2882) <= b and not a;
    outputs(2883) <= not b or a;
    outputs(2884) <= not (a or b);
    outputs(2885) <= a;
    outputs(2886) <= a xor b;
    outputs(2887) <= a or b;
    outputs(2888) <= a or b;
    outputs(2889) <= not b or a;
    outputs(2890) <= not a;
    outputs(2891) <= not a;
    outputs(2892) <= a;
    outputs(2893) <= not (a xor b);
    outputs(2894) <= not (a xor b);
    outputs(2895) <= a or b;
    outputs(2896) <= a;
    outputs(2897) <= not a or b;
    outputs(2898) <= b;
    outputs(2899) <= not a;
    outputs(2900) <= not (a xor b);
    outputs(2901) <= b and not a;
    outputs(2902) <= not (a and b);
    outputs(2903) <= not b;
    outputs(2904) <= b;
    outputs(2905) <= a xor b;
    outputs(2906) <= a;
    outputs(2907) <= not b or a;
    outputs(2908) <= not b;
    outputs(2909) <= not (a xor b);
    outputs(2910) <= a;
    outputs(2911) <= not a or b;
    outputs(2912) <= not a or b;
    outputs(2913) <= not a;
    outputs(2914) <= a or b;
    outputs(2915) <= not b or a;
    outputs(2916) <= b;
    outputs(2917) <= a xor b;
    outputs(2918) <= not (a and b);
    outputs(2919) <= not (a xor b);
    outputs(2920) <= a and not b;
    outputs(2921) <= not a;
    outputs(2922) <= not a or b;
    outputs(2923) <= not (a xor b);
    outputs(2924) <= not b;
    outputs(2925) <= not (a xor b);
    outputs(2926) <= not (a or b);
    outputs(2927) <= a xor b;
    outputs(2928) <= not (a xor b);
    outputs(2929) <= a and not b;
    outputs(2930) <= not b;
    outputs(2931) <= not b;
    outputs(2932) <= a;
    outputs(2933) <= b;
    outputs(2934) <= not a or b;
    outputs(2935) <= not a;
    outputs(2936) <= not (a xor b);
    outputs(2937) <= b;
    outputs(2938) <= not (a and b);
    outputs(2939) <= a;
    outputs(2940) <= not b or a;
    outputs(2941) <= not (a xor b);
    outputs(2942) <= a and not b;
    outputs(2943) <= a or b;
    outputs(2944) <= a and not b;
    outputs(2945) <= not b or a;
    outputs(2946) <= not a;
    outputs(2947) <= not b;
    outputs(2948) <= b;
    outputs(2949) <= b and not a;
    outputs(2950) <= not a;
    outputs(2951) <= a and not b;
    outputs(2952) <= a;
    outputs(2953) <= not (a and b);
    outputs(2954) <= a or b;
    outputs(2955) <= a or b;
    outputs(2956) <= not b;
    outputs(2957) <= a;
    outputs(2958) <= b;
    outputs(2959) <= a;
    outputs(2960) <= a and not b;
    outputs(2961) <= a or b;
    outputs(2962) <= a and b;
    outputs(2963) <= not (a xor b);
    outputs(2964) <= a xor b;
    outputs(2965) <= not (a xor b);
    outputs(2966) <= not b or a;
    outputs(2967) <= not a;
    outputs(2968) <= not a or b;
    outputs(2969) <= a xor b;
    outputs(2970) <= a or b;
    outputs(2971) <= not b or a;
    outputs(2972) <= not (a and b);
    outputs(2973) <= a or b;
    outputs(2974) <= a and not b;
    outputs(2975) <= not a or b;
    outputs(2976) <= not (a xor b);
    outputs(2977) <= not (a xor b);
    outputs(2978) <= not b;
    outputs(2979) <= a xor b;
    outputs(2980) <= a xor b;
    outputs(2981) <= a xor b;
    outputs(2982) <= a and b;
    outputs(2983) <= a xor b;
    outputs(2984) <= a;
    outputs(2985) <= a xor b;
    outputs(2986) <= not b or a;
    outputs(2987) <= not a;
    outputs(2988) <= a;
    outputs(2989) <= b;
    outputs(2990) <= not b;
    outputs(2991) <= not (a and b);
    outputs(2992) <= a;
    outputs(2993) <= not (a xor b);
    outputs(2994) <= not (a and b);
    outputs(2995) <= not b;
    outputs(2996) <= a;
    outputs(2997) <= not (a and b);
    outputs(2998) <= a xor b;
    outputs(2999) <= a xor b;
    outputs(3000) <= not a;
    outputs(3001) <= a;
    outputs(3002) <= a xor b;
    outputs(3003) <= not (a xor b);
    outputs(3004) <= a or b;
    outputs(3005) <= not b;
    outputs(3006) <= a xor b;
    outputs(3007) <= not (a xor b);
    outputs(3008) <= a;
    outputs(3009) <= not a;
    outputs(3010) <= not (a and b);
    outputs(3011) <= a xor b;
    outputs(3012) <= not (a xor b);
    outputs(3013) <= not a or b;
    outputs(3014) <= not b or a;
    outputs(3015) <= not a or b;
    outputs(3016) <= not a;
    outputs(3017) <= not a or b;
    outputs(3018) <= not a;
    outputs(3019) <= a or b;
    outputs(3020) <= not (a and b);
    outputs(3021) <= not a;
    outputs(3022) <= not (a xor b);
    outputs(3023) <= not (a and b);
    outputs(3024) <= a or b;
    outputs(3025) <= b and not a;
    outputs(3026) <= not (a xor b);
    outputs(3027) <= a;
    outputs(3028) <= a;
    outputs(3029) <= a and b;
    outputs(3030) <= not a;
    outputs(3031) <= b;
    outputs(3032) <= a or b;
    outputs(3033) <= a xor b;
    outputs(3034) <= not (a and b);
    outputs(3035) <= a;
    outputs(3036) <= not a or b;
    outputs(3037) <= not (a and b);
    outputs(3038) <= a xor b;
    outputs(3039) <= a;
    outputs(3040) <= a xor b;
    outputs(3041) <= not a or b;
    outputs(3042) <= a xor b;
    outputs(3043) <= a and b;
    outputs(3044) <= not (a xor b);
    outputs(3045) <= not (a or b);
    outputs(3046) <= a xor b;
    outputs(3047) <= a xor b;
    outputs(3048) <= not b;
    outputs(3049) <= a;
    outputs(3050) <= not b or a;
    outputs(3051) <= a or b;
    outputs(3052) <= not b or a;
    outputs(3053) <= not a;
    outputs(3054) <= not (a xor b);
    outputs(3055) <= not (a or b);
    outputs(3056) <= not (a or b);
    outputs(3057) <= a and b;
    outputs(3058) <= a xor b;
    outputs(3059) <= a and b;
    outputs(3060) <= not a;
    outputs(3061) <= not b;
    outputs(3062) <= a;
    outputs(3063) <= not (a xor b);
    outputs(3064) <= not (a xor b);
    outputs(3065) <= not a or b;
    outputs(3066) <= a or b;
    outputs(3067) <= not (a or b);
    outputs(3068) <= a xor b;
    outputs(3069) <= b;
    outputs(3070) <= a and not b;
    outputs(3071) <= not (a xor b);
    outputs(3072) <= a and not b;
    outputs(3073) <= a xor b;
    outputs(3074) <= not a or b;
    outputs(3075) <= not (a and b);
    outputs(3076) <= not a;
    outputs(3077) <= a xor b;
    outputs(3078) <= not b;
    outputs(3079) <= not (a xor b);
    outputs(3080) <= a;
    outputs(3081) <= not (a and b);
    outputs(3082) <= not b or a;
    outputs(3083) <= not a;
    outputs(3084) <= not (a xor b);
    outputs(3085) <= a;
    outputs(3086) <= not (a xor b);
    outputs(3087) <= not a;
    outputs(3088) <= b and not a;
    outputs(3089) <= not (a and b);
    outputs(3090) <= not a;
    outputs(3091) <= not a;
    outputs(3092) <= a;
    outputs(3093) <= a and b;
    outputs(3094) <= a and not b;
    outputs(3095) <= a xor b;
    outputs(3096) <= not a;
    outputs(3097) <= not (a or b);
    outputs(3098) <= not b or a;
    outputs(3099) <= not (a and b);
    outputs(3100) <= not b;
    outputs(3101) <= a and not b;
    outputs(3102) <= a xor b;
    outputs(3103) <= not b or a;
    outputs(3104) <= not a;
    outputs(3105) <= a xor b;
    outputs(3106) <= a xor b;
    outputs(3107) <= a;
    outputs(3108) <= not a;
    outputs(3109) <= a or b;
    outputs(3110) <= a;
    outputs(3111) <= a;
    outputs(3112) <= not (a or b);
    outputs(3113) <= not (a xor b);
    outputs(3114) <= not a;
    outputs(3115) <= a xor b;
    outputs(3116) <= not (a xor b);
    outputs(3117) <= a or b;
    outputs(3118) <= a xor b;
    outputs(3119) <= not a;
    outputs(3120) <= a xor b;
    outputs(3121) <= a;
    outputs(3122) <= not a;
    outputs(3123) <= a or b;
    outputs(3124) <= b;
    outputs(3125) <= a or b;
    outputs(3126) <= not (a or b);
    outputs(3127) <= a and b;
    outputs(3128) <= not a;
    outputs(3129) <= a and not b;
    outputs(3130) <= not (a and b);
    outputs(3131) <= b;
    outputs(3132) <= not a;
    outputs(3133) <= a and not b;
    outputs(3134) <= not (a or b);
    outputs(3135) <= not a or b;
    outputs(3136) <= a;
    outputs(3137) <= a;
    outputs(3138) <= not b;
    outputs(3139) <= not b or a;
    outputs(3140) <= not a;
    outputs(3141) <= not b;
    outputs(3142) <= not b or a;
    outputs(3143) <= b;
    outputs(3144) <= not b;
    outputs(3145) <= a;
    outputs(3146) <= a xor b;
    outputs(3147) <= not b or a;
    outputs(3148) <= a xor b;
    outputs(3149) <= not b;
    outputs(3150) <= a and b;
    outputs(3151) <= not b;
    outputs(3152) <= not b or a;
    outputs(3153) <= not b or a;
    outputs(3154) <= not a;
    outputs(3155) <= not (a or b);
    outputs(3156) <= not b;
    outputs(3157) <= not b or a;
    outputs(3158) <= a and not b;
    outputs(3159) <= a or b;
    outputs(3160) <= not a or b;
    outputs(3161) <= a xor b;
    outputs(3162) <= not a or b;
    outputs(3163) <= not (a xor b);
    outputs(3164) <= b;
    outputs(3165) <= not b or a;
    outputs(3166) <= not b or a;
    outputs(3167) <= not (a and b);
    outputs(3168) <= not (a xor b);
    outputs(3169) <= a xor b;
    outputs(3170) <= a xor b;
    outputs(3171) <= a or b;
    outputs(3172) <= b and not a;
    outputs(3173) <= a xor b;
    outputs(3174) <= not (a and b);
    outputs(3175) <= not b;
    outputs(3176) <= not (a xor b);
    outputs(3177) <= not a;
    outputs(3178) <= b;
    outputs(3179) <= not b;
    outputs(3180) <= not a or b;
    outputs(3181) <= b;
    outputs(3182) <= b;
    outputs(3183) <= a xor b;
    outputs(3184) <= a xor b;
    outputs(3185) <= not b;
    outputs(3186) <= not b;
    outputs(3187) <= a xor b;
    outputs(3188) <= a and not b;
    outputs(3189) <= a xor b;
    outputs(3190) <= b;
    outputs(3191) <= not a or b;
    outputs(3192) <= b;
    outputs(3193) <= not (a or b);
    outputs(3194) <= not (a xor b);
    outputs(3195) <= b;
    outputs(3196) <= not (a or b);
    outputs(3197) <= not a;
    outputs(3198) <= not a;
    outputs(3199) <= not (a or b);
    outputs(3200) <= not b;
    outputs(3201) <= not a;
    outputs(3202) <= a;
    outputs(3203) <= not a or b;
    outputs(3204) <= a or b;
    outputs(3205) <= not a or b;
    outputs(3206) <= a xor b;
    outputs(3207) <= not b;
    outputs(3208) <= a;
    outputs(3209) <= a or b;
    outputs(3210) <= not (a and b);
    outputs(3211) <= b and not a;
    outputs(3212) <= a xor b;
    outputs(3213) <= not a or b;
    outputs(3214) <= a and not b;
    outputs(3215) <= not a;
    outputs(3216) <= not (a xor b);
    outputs(3217) <= a and not b;
    outputs(3218) <= not b;
    outputs(3219) <= b and not a;
    outputs(3220) <= not a or b;
    outputs(3221) <= a xor b;
    outputs(3222) <= not b or a;
    outputs(3223) <= a xor b;
    outputs(3224) <= not (a xor b);
    outputs(3225) <= a and b;
    outputs(3226) <= not a;
    outputs(3227) <= a;
    outputs(3228) <= a or b;
    outputs(3229) <= a or b;
    outputs(3230) <= not a;
    outputs(3231) <= not (a and b);
    outputs(3232) <= not (a xor b);
    outputs(3233) <= not (a and b);
    outputs(3234) <= not (a or b);
    outputs(3235) <= not a;
    outputs(3236) <= a and not b;
    outputs(3237) <= 1'b0;
    outputs(3238) <= a;
    outputs(3239) <= not (a and b);
    outputs(3240) <= not a;
    outputs(3241) <= a and not b;
    outputs(3242) <= not (a xor b);
    outputs(3243) <= a or b;
    outputs(3244) <= a or b;
    outputs(3245) <= b and not a;
    outputs(3246) <= b;
    outputs(3247) <= not b;
    outputs(3248) <= not (a xor b);
    outputs(3249) <= a;
    outputs(3250) <= b;
    outputs(3251) <= a or b;
    outputs(3252) <= not a or b;
    outputs(3253) <= not b or a;
    outputs(3254) <= a;
    outputs(3255) <= not (a xor b);
    outputs(3256) <= a;
    outputs(3257) <= a;
    outputs(3258) <= not (a xor b);
    outputs(3259) <= not a or b;
    outputs(3260) <= not (a or b);
    outputs(3261) <= not b or a;
    outputs(3262) <= not (a or b);
    outputs(3263) <= a xor b;
    outputs(3264) <= a and b;
    outputs(3265) <= not b or a;
    outputs(3266) <= a or b;
    outputs(3267) <= not (a xor b);
    outputs(3268) <= a xor b;
    outputs(3269) <= not (a and b);
    outputs(3270) <= not (a and b);
    outputs(3271) <= not b;
    outputs(3272) <= a;
    outputs(3273) <= a;
    outputs(3274) <= not b;
    outputs(3275) <= not (a xor b);
    outputs(3276) <= a xor b;
    outputs(3277) <= a and not b;
    outputs(3278) <= not (a xor b);
    outputs(3279) <= b;
    outputs(3280) <= not a;
    outputs(3281) <= b and not a;
    outputs(3282) <= b;
    outputs(3283) <= a;
    outputs(3284) <= not b or a;
    outputs(3285) <= a;
    outputs(3286) <= a;
    outputs(3287) <= a and b;
    outputs(3288) <= not b;
    outputs(3289) <= a xor b;
    outputs(3290) <= not b;
    outputs(3291) <= not (a or b);
    outputs(3292) <= b;
    outputs(3293) <= not (a xor b);
    outputs(3294) <= not b;
    outputs(3295) <= not (a and b);
    outputs(3296) <= not (a xor b);
    outputs(3297) <= not b;
    outputs(3298) <= a xor b;
    outputs(3299) <= not b;
    outputs(3300) <= not a;
    outputs(3301) <= not (a xor b);
    outputs(3302) <= b;
    outputs(3303) <= not (a and b);
    outputs(3304) <= b and not a;
    outputs(3305) <= not a;
    outputs(3306) <= b;
    outputs(3307) <= a xor b;
    outputs(3308) <= not b;
    outputs(3309) <= not (a or b);
    outputs(3310) <= a;
    outputs(3311) <= not (a xor b);
    outputs(3312) <= a and not b;
    outputs(3313) <= not b;
    outputs(3314) <= not (a xor b);
    outputs(3315) <= a xor b;
    outputs(3316) <= a xor b;
    outputs(3317) <= not b;
    outputs(3318) <= not (a and b);
    outputs(3319) <= not a;
    outputs(3320) <= b;
    outputs(3321) <= not b;
    outputs(3322) <= not (a xor b);
    outputs(3323) <= not (a and b);
    outputs(3324) <= b;
    outputs(3325) <= not (a xor b);
    outputs(3326) <= not (a xor b);
    outputs(3327) <= a or b;
    outputs(3328) <= not b;
    outputs(3329) <= not a;
    outputs(3330) <= a;
    outputs(3331) <= not b;
    outputs(3332) <= not b or a;
    outputs(3333) <= a or b;
    outputs(3334) <= 1'b1;
    outputs(3335) <= b;
    outputs(3336) <= not b;
    outputs(3337) <= not b;
    outputs(3338) <= b;
    outputs(3339) <= a xor b;
    outputs(3340) <= not b or a;
    outputs(3341) <= a or b;
    outputs(3342) <= b;
    outputs(3343) <= not (a xor b);
    outputs(3344) <= not a or b;
    outputs(3345) <= a xor b;
    outputs(3346) <= not (a xor b);
    outputs(3347) <= not (a and b);
    outputs(3348) <= a;
    outputs(3349) <= not b;
    outputs(3350) <= not (a xor b);
    outputs(3351) <= b;
    outputs(3352) <= not a;
    outputs(3353) <= a xor b;
    outputs(3354) <= a or b;
    outputs(3355) <= not a;
    outputs(3356) <= not (a or b);
    outputs(3357) <= not (a xor b);
    outputs(3358) <= a or b;
    outputs(3359) <= b;
    outputs(3360) <= a;
    outputs(3361) <= a xor b;
    outputs(3362) <= a and b;
    outputs(3363) <= b;
    outputs(3364) <= a xor b;
    outputs(3365) <= b;
    outputs(3366) <= not b;
    outputs(3367) <= not b;
    outputs(3368) <= not (a xor b);
    outputs(3369) <= not (a or b);
    outputs(3370) <= not (a xor b);
    outputs(3371) <= not (a xor b);
    outputs(3372) <= not (a xor b);
    outputs(3373) <= a xor b;
    outputs(3374) <= not (a or b);
    outputs(3375) <= not a or b;
    outputs(3376) <= a and b;
    outputs(3377) <= not b;
    outputs(3378) <= a and not b;
    outputs(3379) <= a xor b;
    outputs(3380) <= not (a and b);
    outputs(3381) <= not b;
    outputs(3382) <= b and not a;
    outputs(3383) <= a and b;
    outputs(3384) <= not b;
    outputs(3385) <= not b;
    outputs(3386) <= not a;
    outputs(3387) <= not a or b;
    outputs(3388) <= not (a xor b);
    outputs(3389) <= a;
    outputs(3390) <= a;
    outputs(3391) <= a;
    outputs(3392) <= a;
    outputs(3393) <= not a or b;
    outputs(3394) <= not a;
    outputs(3395) <= not (a and b);
    outputs(3396) <= not a;
    outputs(3397) <= not b;
    outputs(3398) <= a;
    outputs(3399) <= a xor b;
    outputs(3400) <= not b or a;
    outputs(3401) <= not b;
    outputs(3402) <= not a;
    outputs(3403) <= not a;
    outputs(3404) <= a and b;
    outputs(3405) <= not (a or b);
    outputs(3406) <= a or b;
    outputs(3407) <= not (a xor b);
    outputs(3408) <= not (a xor b);
    outputs(3409) <= a and not b;
    outputs(3410) <= a xor b;
    outputs(3411) <= a;
    outputs(3412) <= not a;
    outputs(3413) <= not (a xor b);
    outputs(3414) <= not b;
    outputs(3415) <= not b;
    outputs(3416) <= a xor b;
    outputs(3417) <= a xor b;
    outputs(3418) <= a;
    outputs(3419) <= not b or a;
    outputs(3420) <= not (a xor b);
    outputs(3421) <= not a or b;
    outputs(3422) <= not a;
    outputs(3423) <= b;
    outputs(3424) <= not a or b;
    outputs(3425) <= b;
    outputs(3426) <= not a or b;
    outputs(3427) <= a;
    outputs(3428) <= a xor b;
    outputs(3429) <= not a;
    outputs(3430) <= not b or a;
    outputs(3431) <= a xor b;
    outputs(3432) <= a;
    outputs(3433) <= not (a and b);
    outputs(3434) <= not (a xor b);
    outputs(3435) <= b;
    outputs(3436) <= not (a xor b);
    outputs(3437) <= a and b;
    outputs(3438) <= not b;
    outputs(3439) <= not b;
    outputs(3440) <= not a;
    outputs(3441) <= a;
    outputs(3442) <= b;
    outputs(3443) <= a or b;
    outputs(3444) <= a or b;
    outputs(3445) <= a xor b;
    outputs(3446) <= not (a xor b);
    outputs(3447) <= not a;
    outputs(3448) <= not a;
    outputs(3449) <= a or b;
    outputs(3450) <= not a;
    outputs(3451) <= not (a and b);
    outputs(3452) <= not a or b;
    outputs(3453) <= not b;
    outputs(3454) <= a;
    outputs(3455) <= a and not b;
    outputs(3456) <= not (a xor b);
    outputs(3457) <= not b or a;
    outputs(3458) <= b;
    outputs(3459) <= not a;
    outputs(3460) <= not (a xor b);
    outputs(3461) <= a and not b;
    outputs(3462) <= not (a and b);
    outputs(3463) <= b and not a;
    outputs(3464) <= a;
    outputs(3465) <= not a;
    outputs(3466) <= not a;
    outputs(3467) <= not (a and b);
    outputs(3468) <= not a;
    outputs(3469) <= a or b;
    outputs(3470) <= not a or b;
    outputs(3471) <= a;
    outputs(3472) <= a;
    outputs(3473) <= b;
    outputs(3474) <= a and not b;
    outputs(3475) <= a;
    outputs(3476) <= a xor b;
    outputs(3477) <= a xor b;
    outputs(3478) <= b;
    outputs(3479) <= a xor b;
    outputs(3480) <= not a;
    outputs(3481) <= a xor b;
    outputs(3482) <= a xor b;
    outputs(3483) <= not a;
    outputs(3484) <= not b or a;
    outputs(3485) <= a xor b;
    outputs(3486) <= a or b;
    outputs(3487) <= not a or b;
    outputs(3488) <= a xor b;
    outputs(3489) <= not a;
    outputs(3490) <= not a;
    outputs(3491) <= not a;
    outputs(3492) <= not a or b;
    outputs(3493) <= not (a and b);
    outputs(3494) <= a xor b;
    outputs(3495) <= not b;
    outputs(3496) <= a xor b;
    outputs(3497) <= not (a xor b);
    outputs(3498) <= not a or b;
    outputs(3499) <= not b;
    outputs(3500) <= not (a and b);
    outputs(3501) <= not a;
    outputs(3502) <= not (a xor b);
    outputs(3503) <= a or b;
    outputs(3504) <= not b or a;
    outputs(3505) <= a xor b;
    outputs(3506) <= b;
    outputs(3507) <= not b or a;
    outputs(3508) <= b;
    outputs(3509) <= not b or a;
    outputs(3510) <= a xor b;
    outputs(3511) <= b and not a;
    outputs(3512) <= b;
    outputs(3513) <= a xor b;
    outputs(3514) <= not (a or b);
    outputs(3515) <= a or b;
    outputs(3516) <= not (a xor b);
    outputs(3517) <= not b;
    outputs(3518) <= a;
    outputs(3519) <= not (a xor b);
    outputs(3520) <= not (a and b);
    outputs(3521) <= a or b;
    outputs(3522) <= not (a or b);
    outputs(3523) <= not (a xor b);
    outputs(3524) <= not b or a;
    outputs(3525) <= a xor b;
    outputs(3526) <= b;
    outputs(3527) <= a and b;
    outputs(3528) <= not b or a;
    outputs(3529) <= a xor b;
    outputs(3530) <= not b or a;
    outputs(3531) <= a xor b;
    outputs(3532) <= not (a and b);
    outputs(3533) <= b;
    outputs(3534) <= a;
    outputs(3535) <= a;
    outputs(3536) <= not a;
    outputs(3537) <= a;
    outputs(3538) <= not a;
    outputs(3539) <= not (a xor b);
    outputs(3540) <= b and not a;
    outputs(3541) <= b;
    outputs(3542) <= a xor b;
    outputs(3543) <= not (a xor b);
    outputs(3544) <= b;
    outputs(3545) <= a xor b;
    outputs(3546) <= a xor b;
    outputs(3547) <= b;
    outputs(3548) <= a;
    outputs(3549) <= a;
    outputs(3550) <= a xor b;
    outputs(3551) <= not b;
    outputs(3552) <= not (a and b);
    outputs(3553) <= a xor b;
    outputs(3554) <= not b or a;
    outputs(3555) <= b;
    outputs(3556) <= not b or a;
    outputs(3557) <= not (a and b);
    outputs(3558) <= a xor b;
    outputs(3559) <= not (a xor b);
    outputs(3560) <= b;
    outputs(3561) <= not a;
    outputs(3562) <= a or b;
    outputs(3563) <= a and b;
    outputs(3564) <= not (a and b);
    outputs(3565) <= a;
    outputs(3566) <= not (a xor b);
    outputs(3567) <= a xor b;
    outputs(3568) <= not (a xor b);
    outputs(3569) <= not (a and b);
    outputs(3570) <= a;
    outputs(3571) <= not b;
    outputs(3572) <= not b;
    outputs(3573) <= b;
    outputs(3574) <= a xor b;
    outputs(3575) <= a or b;
    outputs(3576) <= a xor b;
    outputs(3577) <= not b or a;
    outputs(3578) <= a xor b;
    outputs(3579) <= not a;
    outputs(3580) <= a;
    outputs(3581) <= b;
    outputs(3582) <= not b;
    outputs(3583) <= not a;
    outputs(3584) <= not a;
    outputs(3585) <= not (a xor b);
    outputs(3586) <= not b or a;
    outputs(3587) <= not (a xor b);
    outputs(3588) <= not a;
    outputs(3589) <= not (a and b);
    outputs(3590) <= not a;
    outputs(3591) <= b;
    outputs(3592) <= b;
    outputs(3593) <= a and not b;
    outputs(3594) <= 1'b1;
    outputs(3595) <= a and not b;
    outputs(3596) <= a xor b;
    outputs(3597) <= not (a and b);
    outputs(3598) <= not (a and b);
    outputs(3599) <= not a or b;
    outputs(3600) <= not a or b;
    outputs(3601) <= b and not a;
    outputs(3602) <= not (a xor b);
    outputs(3603) <= a and b;
    outputs(3604) <= a and not b;
    outputs(3605) <= not b;
    outputs(3606) <= a xor b;
    outputs(3607) <= a or b;
    outputs(3608) <= not a or b;
    outputs(3609) <= not a or b;
    outputs(3610) <= not (a xor b);
    outputs(3611) <= a xor b;
    outputs(3612) <= a;
    outputs(3613) <= b and not a;
    outputs(3614) <= not b;
    outputs(3615) <= not (a xor b);
    outputs(3616) <= not b or a;
    outputs(3617) <= not (a xor b);
    outputs(3618) <= not (a or b);
    outputs(3619) <= not b or a;
    outputs(3620) <= not b or a;
    outputs(3621) <= b;
    outputs(3622) <= b;
    outputs(3623) <= b and not a;
    outputs(3624) <= a and not b;
    outputs(3625) <= not b or a;
    outputs(3626) <= a xor b;
    outputs(3627) <= not a or b;
    outputs(3628) <= not (a and b);
    outputs(3629) <= a;
    outputs(3630) <= not a;
    outputs(3631) <= b and not a;
    outputs(3632) <= not (a xor b);
    outputs(3633) <= a xor b;
    outputs(3634) <= not a or b;
    outputs(3635) <= a xor b;
    outputs(3636) <= not (a xor b);
    outputs(3637) <= not (a xor b);
    outputs(3638) <= b and not a;
    outputs(3639) <= a and b;
    outputs(3640) <= a or b;
    outputs(3641) <= a and not b;
    outputs(3642) <= b;
    outputs(3643) <= a;
    outputs(3644) <= a;
    outputs(3645) <= a or b;
    outputs(3646) <= not a;
    outputs(3647) <= a xor b;
    outputs(3648) <= not (a xor b);
    outputs(3649) <= not b or a;
    outputs(3650) <= a xor b;
    outputs(3651) <= a or b;
    outputs(3652) <= not b;
    outputs(3653) <= a or b;
    outputs(3654) <= not b;
    outputs(3655) <= a xor b;
    outputs(3656) <= a xor b;
    outputs(3657) <= not a;
    outputs(3658) <= not b;
    outputs(3659) <= not b;
    outputs(3660) <= a xor b;
    outputs(3661) <= a xor b;
    outputs(3662) <= a or b;
    outputs(3663) <= a and not b;
    outputs(3664) <= a xor b;
    outputs(3665) <= not (a and b);
    outputs(3666) <= not b or a;
    outputs(3667) <= not b;
    outputs(3668) <= a xor b;
    outputs(3669) <= not b;
    outputs(3670) <= a;
    outputs(3671) <= not b or a;
    outputs(3672) <= a xor b;
    outputs(3673) <= a;
    outputs(3674) <= not (a and b);
    outputs(3675) <= not (a or b);
    outputs(3676) <= a xor b;
    outputs(3677) <= not b;
    outputs(3678) <= not (a xor b);
    outputs(3679) <= not a;
    outputs(3680) <= b;
    outputs(3681) <= b;
    outputs(3682) <= not (a xor b);
    outputs(3683) <= not (a and b);
    outputs(3684) <= a xor b;
    outputs(3685) <= not b or a;
    outputs(3686) <= not b;
    outputs(3687) <= a or b;
    outputs(3688) <= a and b;
    outputs(3689) <= not (a xor b);
    outputs(3690) <= not b;
    outputs(3691) <= not (a or b);
    outputs(3692) <= a xor b;
    outputs(3693) <= not (a and b);
    outputs(3694) <= a and not b;
    outputs(3695) <= a xor b;
    outputs(3696) <= not (a xor b);
    outputs(3697) <= not (a and b);
    outputs(3698) <= a and b;
    outputs(3699) <= not b;
    outputs(3700) <= a xor b;
    outputs(3701) <= not b;
    outputs(3702) <= not (a xor b);
    outputs(3703) <= b;
    outputs(3704) <= not a or b;
    outputs(3705) <= b;
    outputs(3706) <= not (a xor b);
    outputs(3707) <= a xor b;
    outputs(3708) <= not b;
    outputs(3709) <= a xor b;
    outputs(3710) <= a or b;
    outputs(3711) <= a;
    outputs(3712) <= a xor b;
    outputs(3713) <= a or b;
    outputs(3714) <= not (a xor b);
    outputs(3715) <= not b;
    outputs(3716) <= a xor b;
    outputs(3717) <= not (a xor b);
    outputs(3718) <= not a;
    outputs(3719) <= b and not a;
    outputs(3720) <= not a or b;
    outputs(3721) <= b;
    outputs(3722) <= a and b;
    outputs(3723) <= not b;
    outputs(3724) <= not (a xor b);
    outputs(3725) <= a or b;
    outputs(3726) <= a;
    outputs(3727) <= not (a xor b);
    outputs(3728) <= b;
    outputs(3729) <= not (a xor b);
    outputs(3730) <= not (a xor b);
    outputs(3731) <= not a or b;
    outputs(3732) <= b and not a;
    outputs(3733) <= a;
    outputs(3734) <= not (a xor b);
    outputs(3735) <= a or b;
    outputs(3736) <= not (a xor b);
    outputs(3737) <= not (a xor b);
    outputs(3738) <= a xor b;
    outputs(3739) <= a xor b;
    outputs(3740) <= not a;
    outputs(3741) <= not a or b;
    outputs(3742) <= not a or b;
    outputs(3743) <= not b or a;
    outputs(3744) <= a xor b;
    outputs(3745) <= a xor b;
    outputs(3746) <= a or b;
    outputs(3747) <= not b;
    outputs(3748) <= a;
    outputs(3749) <= a xor b;
    outputs(3750) <= not a;
    outputs(3751) <= a and not b;
    outputs(3752) <= a;
    outputs(3753) <= not b;
    outputs(3754) <= not a;
    outputs(3755) <= not (a and b);
    outputs(3756) <= a xor b;
    outputs(3757) <= not b;
    outputs(3758) <= not b;
    outputs(3759) <= not (a or b);
    outputs(3760) <= not (a xor b);
    outputs(3761) <= not (a or b);
    outputs(3762) <= not a or b;
    outputs(3763) <= a or b;
    outputs(3764) <= a xor b;
    outputs(3765) <= not a;
    outputs(3766) <= not b or a;
    outputs(3767) <= a;
    outputs(3768) <= not (a xor b);
    outputs(3769) <= not (a and b);
    outputs(3770) <= b and not a;
    outputs(3771) <= a;
    outputs(3772) <= a or b;
    outputs(3773) <= b;
    outputs(3774) <= not (a xor b);
    outputs(3775) <= a;
    outputs(3776) <= b;
    outputs(3777) <= a or b;
    outputs(3778) <= a or b;
    outputs(3779) <= a;
    outputs(3780) <= a;
    outputs(3781) <= b;
    outputs(3782) <= not a or b;
    outputs(3783) <= not a or b;
    outputs(3784) <= a;
    outputs(3785) <= b;
    outputs(3786) <= a xor b;
    outputs(3787) <= not b or a;
    outputs(3788) <= a xor b;
    outputs(3789) <= not (a xor b);
    outputs(3790) <= not a;
    outputs(3791) <= not b;
    outputs(3792) <= b;
    outputs(3793) <= not b;
    outputs(3794) <= a xor b;
    outputs(3795) <= a xor b;
    outputs(3796) <= not (a xor b);
    outputs(3797) <= not b or a;
    outputs(3798) <= not b or a;
    outputs(3799) <= a or b;
    outputs(3800) <= not a or b;
    outputs(3801) <= b and not a;
    outputs(3802) <= not a;
    outputs(3803) <= not a;
    outputs(3804) <= not a or b;
    outputs(3805) <= not b;
    outputs(3806) <= a;
    outputs(3807) <= b;
    outputs(3808) <= b and not a;
    outputs(3809) <= b and not a;
    outputs(3810) <= a xor b;
    outputs(3811) <= not (a xor b);
    outputs(3812) <= b;
    outputs(3813) <= not (a and b);
    outputs(3814) <= b;
    outputs(3815) <= a;
    outputs(3816) <= not (a and b);
    outputs(3817) <= not (a and b);
    outputs(3818) <= b and not a;
    outputs(3819) <= not (a and b);
    outputs(3820) <= b and not a;
    outputs(3821) <= a;
    outputs(3822) <= a or b;
    outputs(3823) <= not a or b;
    outputs(3824) <= not a or b;
    outputs(3825) <= a xor b;
    outputs(3826) <= b;
    outputs(3827) <= a and not b;
    outputs(3828) <= not (a and b);
    outputs(3829) <= a xor b;
    outputs(3830) <= not b;
    outputs(3831) <= a and not b;
    outputs(3832) <= not a or b;
    outputs(3833) <= a xor b;
    outputs(3834) <= not a;
    outputs(3835) <= not (a xor b);
    outputs(3836) <= b and not a;
    outputs(3837) <= a xor b;
    outputs(3838) <= b and not a;
    outputs(3839) <= a;
    outputs(3840) <= b;
    outputs(3841) <= not (a xor b);
    outputs(3842) <= b and not a;
    outputs(3843) <= not (a or b);
    outputs(3844) <= not a or b;
    outputs(3845) <= not (a xor b);
    outputs(3846) <= not (a xor b);
    outputs(3847) <= not (a xor b);
    outputs(3848) <= not a;
    outputs(3849) <= a;
    outputs(3850) <= not (a or b);
    outputs(3851) <= not (a xor b);
    outputs(3852) <= not a;
    outputs(3853) <= a xor b;
    outputs(3854) <= not (a xor b);
    outputs(3855) <= a or b;
    outputs(3856) <= not (a xor b);
    outputs(3857) <= b and not a;
    outputs(3858) <= not (a and b);
    outputs(3859) <= not b;
    outputs(3860) <= b;
    outputs(3861) <= b;
    outputs(3862) <= not b;
    outputs(3863) <= a;
    outputs(3864) <= not a;
    outputs(3865) <= a xor b;
    outputs(3866) <= not (a xor b);
    outputs(3867) <= not b;
    outputs(3868) <= not b;
    outputs(3869) <= not (a xor b);
    outputs(3870) <= a and b;
    outputs(3871) <= not (a xor b);
    outputs(3872) <= a xor b;
    outputs(3873) <= a or b;
    outputs(3874) <= a or b;
    outputs(3875) <= not b;
    outputs(3876) <= a or b;
    outputs(3877) <= b and not a;
    outputs(3878) <= not (a xor b);
    outputs(3879) <= not b or a;
    outputs(3880) <= not a;
    outputs(3881) <= a;
    outputs(3882) <= a;
    outputs(3883) <= not (a xor b);
    outputs(3884) <= b;
    outputs(3885) <= not a or b;
    outputs(3886) <= a or b;
    outputs(3887) <= not (a and b);
    outputs(3888) <= not (a or b);
    outputs(3889) <= b and not a;
    outputs(3890) <= b and not a;
    outputs(3891) <= a xor b;
    outputs(3892) <= not (a xor b);
    outputs(3893) <= a xor b;
    outputs(3894) <= b;
    outputs(3895) <= a xor b;
    outputs(3896) <= not b or a;
    outputs(3897) <= not (a and b);
    outputs(3898) <= a xor b;
    outputs(3899) <= b;
    outputs(3900) <= not a or b;
    outputs(3901) <= not (a xor b);
    outputs(3902) <= a xor b;
    outputs(3903) <= not b or a;
    outputs(3904) <= a xor b;
    outputs(3905) <= not (a xor b);
    outputs(3906) <= not (a xor b);
    outputs(3907) <= not a or b;
    outputs(3908) <= b;
    outputs(3909) <= not a;
    outputs(3910) <= not a or b;
    outputs(3911) <= not b;
    outputs(3912) <= a and b;
    outputs(3913) <= a xor b;
    outputs(3914) <= b;
    outputs(3915) <= b;
    outputs(3916) <= a;
    outputs(3917) <= not (a and b);
    outputs(3918) <= not (a or b);
    outputs(3919) <= b and not a;
    outputs(3920) <= a xor b;
    outputs(3921) <= not (a and b);
    outputs(3922) <= b;
    outputs(3923) <= not (a xor b);
    outputs(3924) <= not (a or b);
    outputs(3925) <= not a or b;
    outputs(3926) <= not b;
    outputs(3927) <= not (a and b);
    outputs(3928) <= a and b;
    outputs(3929) <= b;
    outputs(3930) <= a xor b;
    outputs(3931) <= a xor b;
    outputs(3932) <= not b;
    outputs(3933) <= not a or b;
    outputs(3934) <= not b;
    outputs(3935) <= not a or b;
    outputs(3936) <= not (a and b);
    outputs(3937) <= a xor b;
    outputs(3938) <= a and b;
    outputs(3939) <= a;
    outputs(3940) <= a and b;
    outputs(3941) <= not b;
    outputs(3942) <= a;
    outputs(3943) <= not a or b;
    outputs(3944) <= not a or b;
    outputs(3945) <= a;
    outputs(3946) <= a xor b;
    outputs(3947) <= a;
    outputs(3948) <= not (a and b);
    outputs(3949) <= not (a and b);
    outputs(3950) <= b and not a;
    outputs(3951) <= not a or b;
    outputs(3952) <= a xor b;
    outputs(3953) <= not a;
    outputs(3954) <= b;
    outputs(3955) <= b;
    outputs(3956) <= a;
    outputs(3957) <= a;
    outputs(3958) <= a;
    outputs(3959) <= a or b;
    outputs(3960) <= a and not b;
    outputs(3961) <= not a;
    outputs(3962) <= not (a xor b);
    outputs(3963) <= a xor b;
    outputs(3964) <= not a or b;
    outputs(3965) <= not (a xor b);
    outputs(3966) <= not b;
    outputs(3967) <= not (a and b);
    outputs(3968) <= not (a or b);
    outputs(3969) <= b;
    outputs(3970) <= a or b;
    outputs(3971) <= not b;
    outputs(3972) <= a and b;
    outputs(3973) <= a xor b;
    outputs(3974) <= b;
    outputs(3975) <= a;
    outputs(3976) <= not (a xor b);
    outputs(3977) <= not b or a;
    outputs(3978) <= a and b;
    outputs(3979) <= not (a and b);
    outputs(3980) <= not a or b;
    outputs(3981) <= not (a and b);
    outputs(3982) <= not (a or b);
    outputs(3983) <= not (a or b);
    outputs(3984) <= not (a xor b);
    outputs(3985) <= b;
    outputs(3986) <= b;
    outputs(3987) <= b and not a;
    outputs(3988) <= not a;
    outputs(3989) <= a xor b;
    outputs(3990) <= a xor b;
    outputs(3991) <= not b;
    outputs(3992) <= not b or a;
    outputs(3993) <= a xor b;
    outputs(3994) <= not a or b;
    outputs(3995) <= a and b;
    outputs(3996) <= not (a xor b);
    outputs(3997) <= not a;
    outputs(3998) <= not a;
    outputs(3999) <= b;
    outputs(4000) <= a xor b;
    outputs(4001) <= a xor b;
    outputs(4002) <= a and not b;
    outputs(4003) <= not (a or b);
    outputs(4004) <= a xor b;
    outputs(4005) <= not b;
    outputs(4006) <= b;
    outputs(4007) <= a xor b;
    outputs(4008) <= b and not a;
    outputs(4009) <= a xor b;
    outputs(4010) <= a;
    outputs(4011) <= a;
    outputs(4012) <= a and b;
    outputs(4013) <= a and not b;
    outputs(4014) <= a or b;
    outputs(4015) <= b;
    outputs(4016) <= not (a xor b);
    outputs(4017) <= not b or a;
    outputs(4018) <= a and not b;
    outputs(4019) <= not (a xor b);
    outputs(4020) <= not a or b;
    outputs(4021) <= not a;
    outputs(4022) <= a and not b;
    outputs(4023) <= not a or b;
    outputs(4024) <= not b;
    outputs(4025) <= a and not b;
    outputs(4026) <= not (a or b);
    outputs(4027) <= not a or b;
    outputs(4028) <= a xor b;
    outputs(4029) <= not b;
    outputs(4030) <= not (a xor b);
    outputs(4031) <= b;
    outputs(4032) <= not (a xor b);
    outputs(4033) <= a xor b;
    outputs(4034) <= not a;
    outputs(4035) <= a xor b;
    outputs(4036) <= not a;
    outputs(4037) <= not b;
    outputs(4038) <= a xor b;
    outputs(4039) <= not (a and b);
    outputs(4040) <= not (a xor b);
    outputs(4041) <= not b or a;
    outputs(4042) <= not a;
    outputs(4043) <= a xor b;
    outputs(4044) <= a and b;
    outputs(4045) <= a;
    outputs(4046) <= a;
    outputs(4047) <= a xor b;
    outputs(4048) <= a and b;
    outputs(4049) <= not b or a;
    outputs(4050) <= a xor b;
    outputs(4051) <= a and b;
    outputs(4052) <= not b;
    outputs(4053) <= not (a and b);
    outputs(4054) <= not (a xor b);
    outputs(4055) <= not (a xor b);
    outputs(4056) <= not b;
    outputs(4057) <= not a;
    outputs(4058) <= a;
    outputs(4059) <= b and not a;
    outputs(4060) <= a and not b;
    outputs(4061) <= a and b;
    outputs(4062) <= not a or b;
    outputs(4063) <= not a;
    outputs(4064) <= not a or b;
    outputs(4065) <= a xor b;
    outputs(4066) <= b and not a;
    outputs(4067) <= a;
    outputs(4068) <= a xor b;
    outputs(4069) <= a xor b;
    outputs(4070) <= a and b;
    outputs(4071) <= not (a or b);
    outputs(4072) <= not (a xor b);
    outputs(4073) <= a xor b;
    outputs(4074) <= a;
    outputs(4075) <= not a or b;
    outputs(4076) <= a;
    outputs(4077) <= b and not a;
    outputs(4078) <= not (a xor b);
    outputs(4079) <= not (a xor b);
    outputs(4080) <= a xor b;
    outputs(4081) <= a or b;
    outputs(4082) <= not (a xor b);
    outputs(4083) <= a xor b;
    outputs(4084) <= not (a xor b);
    outputs(4085) <= a xor b;
    outputs(4086) <= not (a and b);
    outputs(4087) <= not b;
    outputs(4088) <= a xor b;
    outputs(4089) <= a and not b;
    outputs(4090) <= not (a xor b);
    outputs(4091) <= not a;
    outputs(4092) <= not (a xor b);
    outputs(4093) <= b;
    outputs(4094) <= not b;
    outputs(4095) <= not (a xor b);
    outputs(4096) <= not (a xor b);
    outputs(4097) <= b and not a;
    outputs(4098) <= b and not a;
    outputs(4099) <= a;
    outputs(4100) <= b;
    outputs(4101) <= a xor b;
    outputs(4102) <= b and not a;
    outputs(4103) <= not (a and b);
    outputs(4104) <= not b or a;
    outputs(4105) <= not a;
    outputs(4106) <= a;
    outputs(4107) <= a xor b;
    outputs(4108) <= a and not b;
    outputs(4109) <= not (a xor b);
    outputs(4110) <= not b or a;
    outputs(4111) <= not a;
    outputs(4112) <= not (a xor b);
    outputs(4113) <= a;
    outputs(4114) <= a or b;
    outputs(4115) <= not a;
    outputs(4116) <= not b;
    outputs(4117) <= not a;
    outputs(4118) <= a;
    outputs(4119) <= a;
    outputs(4120) <= not (a xor b);
    outputs(4121) <= not (a and b);
    outputs(4122) <= b;
    outputs(4123) <= a and b;
    outputs(4124) <= b;
    outputs(4125) <= a and not b;
    outputs(4126) <= not (a and b);
    outputs(4127) <= not b or a;
    outputs(4128) <= a and b;
    outputs(4129) <= not (a and b);
    outputs(4130) <= a xor b;
    outputs(4131) <= not b;
    outputs(4132) <= not (a xor b);
    outputs(4133) <= not b;
    outputs(4134) <= a or b;
    outputs(4135) <= not a or b;
    outputs(4136) <= a or b;
    outputs(4137) <= not b or a;
    outputs(4138) <= not a;
    outputs(4139) <= not (a xor b);
    outputs(4140) <= not (a xor b);
    outputs(4141) <= not (a xor b);
    outputs(4142) <= a and not b;
    outputs(4143) <= not (a xor b);
    outputs(4144) <= 1'b1;
    outputs(4145) <= not b;
    outputs(4146) <= not (a xor b);
    outputs(4147) <= not (a xor b);
    outputs(4148) <= not (a xor b);
    outputs(4149) <= a and not b;
    outputs(4150) <= not a;
    outputs(4151) <= a xor b;
    outputs(4152) <= not (a or b);
    outputs(4153) <= not b;
    outputs(4154) <= a xor b;
    outputs(4155) <= not b;
    outputs(4156) <= a and b;
    outputs(4157) <= not (a xor b);
    outputs(4158) <= not b;
    outputs(4159) <= a or b;
    outputs(4160) <= a xor b;
    outputs(4161) <= not b;
    outputs(4162) <= b and not a;
    outputs(4163) <= not (a or b);
    outputs(4164) <= not b or a;
    outputs(4165) <= not (a and b);
    outputs(4166) <= not a or b;
    outputs(4167) <= a xor b;
    outputs(4168) <= a and b;
    outputs(4169) <= not a or b;
    outputs(4170) <= not (a xor b);
    outputs(4171) <= not (a or b);
    outputs(4172) <= not a;
    outputs(4173) <= a and not b;
    outputs(4174) <= not b;
    outputs(4175) <= not (a xor b);
    outputs(4176) <= b;
    outputs(4177) <= not a;
    outputs(4178) <= not (a xor b);
    outputs(4179) <= not (a or b);
    outputs(4180) <= a xor b;
    outputs(4181) <= a xor b;
    outputs(4182) <= a and b;
    outputs(4183) <= a xor b;
    outputs(4184) <= not (a and b);
    outputs(4185) <= not a or b;
    outputs(4186) <= not a;
    outputs(4187) <= a xor b;
    outputs(4188) <= not (a and b);
    outputs(4189) <= a xor b;
    outputs(4190) <= a xor b;
    outputs(4191) <= a;
    outputs(4192) <= a;
    outputs(4193) <= a xor b;
    outputs(4194) <= not (a and b);
    outputs(4195) <= not (a xor b);
    outputs(4196) <= b and not a;
    outputs(4197) <= a and not b;
    outputs(4198) <= not b;
    outputs(4199) <= b and not a;
    outputs(4200) <= not (a xor b);
    outputs(4201) <= not (a xor b);
    outputs(4202) <= not (a or b);
    outputs(4203) <= not (a and b);
    outputs(4204) <= not b;
    outputs(4205) <= a xor b;
    outputs(4206) <= b;
    outputs(4207) <= b;
    outputs(4208) <= not a;
    outputs(4209) <= a xor b;
    outputs(4210) <= not (a or b);
    outputs(4211) <= not a or b;
    outputs(4212) <= not a;
    outputs(4213) <= not a;
    outputs(4214) <= not a;
    outputs(4215) <= not a;
    outputs(4216) <= not b;
    outputs(4217) <= a xor b;
    outputs(4218) <= b;
    outputs(4219) <= not (a or b);
    outputs(4220) <= not (a xor b);
    outputs(4221) <= a xor b;
    outputs(4222) <= not b;
    outputs(4223) <= b;
    outputs(4224) <= a or b;
    outputs(4225) <= not (a xor b);
    outputs(4226) <= a xor b;
    outputs(4227) <= not (a xor b);
    outputs(4228) <= not (a or b);
    outputs(4229) <= not b;
    outputs(4230) <= a;
    outputs(4231) <= not a or b;
    outputs(4232) <= b;
    outputs(4233) <= a xor b;
    outputs(4234) <= not b or a;
    outputs(4235) <= not (a xor b);
    outputs(4236) <= not a or b;
    outputs(4237) <= not (a xor b);
    outputs(4238) <= not (a xor b);
    outputs(4239) <= a;
    outputs(4240) <= a;
    outputs(4241) <= not (a or b);
    outputs(4242) <= b;
    outputs(4243) <= a;
    outputs(4244) <= not b or a;
    outputs(4245) <= not b;
    outputs(4246) <= not b;
    outputs(4247) <= not b;
    outputs(4248) <= not (a xor b);
    outputs(4249) <= not b;
    outputs(4250) <= not b;
    outputs(4251) <= not b;
    outputs(4252) <= a xor b;
    outputs(4253) <= b;
    outputs(4254) <= a and b;
    outputs(4255) <= a and not b;
    outputs(4256) <= not a;
    outputs(4257) <= not b or a;
    outputs(4258) <= not a;
    outputs(4259) <= a or b;
    outputs(4260) <= not (a or b);
    outputs(4261) <= not (a or b);
    outputs(4262) <= not b or a;
    outputs(4263) <= not b or a;
    outputs(4264) <= not b;
    outputs(4265) <= not (a and b);
    outputs(4266) <= a or b;
    outputs(4267) <= a or b;
    outputs(4268) <= not b;
    outputs(4269) <= not (a and b);
    outputs(4270) <= not (a or b);
    outputs(4271) <= not a;
    outputs(4272) <= not a or b;
    outputs(4273) <= not b or a;
    outputs(4274) <= not b;
    outputs(4275) <= a xor b;
    outputs(4276) <= b;
    outputs(4277) <= b and not a;
    outputs(4278) <= a xor b;
    outputs(4279) <= a xor b;
    outputs(4280) <= b and not a;
    outputs(4281) <= not b or a;
    outputs(4282) <= not (a xor b);
    outputs(4283) <= not (a or b);
    outputs(4284) <= not (a xor b);
    outputs(4285) <= a and b;
    outputs(4286) <= b;
    outputs(4287) <= a;
    outputs(4288) <= a or b;
    outputs(4289) <= a and not b;
    outputs(4290) <= a and not b;
    outputs(4291) <= a;
    outputs(4292) <= not a;
    outputs(4293) <= not (a xor b);
    outputs(4294) <= a xor b;
    outputs(4295) <= a xor b;
    outputs(4296) <= a xor b;
    outputs(4297) <= not a or b;
    outputs(4298) <= a;
    outputs(4299) <= not b or a;
    outputs(4300) <= a or b;
    outputs(4301) <= a xor b;
    outputs(4302) <= not a or b;
    outputs(4303) <= a and not b;
    outputs(4304) <= a;
    outputs(4305) <= a;
    outputs(4306) <= not (a and b);
    outputs(4307) <= not (a and b);
    outputs(4308) <= not b;
    outputs(4309) <= not (a xor b);
    outputs(4310) <= not a;
    outputs(4311) <= a xor b;
    outputs(4312) <= not b or a;
    outputs(4313) <= not a or b;
    outputs(4314) <= a;
    outputs(4315) <= not a or b;
    outputs(4316) <= a;
    outputs(4317) <= not (a xor b);
    outputs(4318) <= a;
    outputs(4319) <= a;
    outputs(4320) <= a or b;
    outputs(4321) <= a and b;
    outputs(4322) <= a or b;
    outputs(4323) <= a xor b;
    outputs(4324) <= not a;
    outputs(4325) <= a and b;
    outputs(4326) <= not (a xor b);
    outputs(4327) <= not (a xor b);
    outputs(4328) <= not (a xor b);
    outputs(4329) <= not a;
    outputs(4330) <= not a;
    outputs(4331) <= not (a xor b);
    outputs(4332) <= b;
    outputs(4333) <= not (a or b);
    outputs(4334) <= not (a or b);
    outputs(4335) <= not b;
    outputs(4336) <= a xor b;
    outputs(4337) <= b;
    outputs(4338) <= a and b;
    outputs(4339) <= a xor b;
    outputs(4340) <= a xor b;
    outputs(4341) <= a xor b;
    outputs(4342) <= b and not a;
    outputs(4343) <= not (a xor b);
    outputs(4344) <= not (a xor b);
    outputs(4345) <= not b;
    outputs(4346) <= a or b;
    outputs(4347) <= b and not a;
    outputs(4348) <= a or b;
    outputs(4349) <= not (a or b);
    outputs(4350) <= b and not a;
    outputs(4351) <= not (a xor b);
    outputs(4352) <= a and b;
    outputs(4353) <= not b or a;
    outputs(4354) <= not b or a;
    outputs(4355) <= not (a xor b);
    outputs(4356) <= b;
    outputs(4357) <= a;
    outputs(4358) <= a and not b;
    outputs(4359) <= a or b;
    outputs(4360) <= not a or b;
    outputs(4361) <= not b;
    outputs(4362) <= not b or a;
    outputs(4363) <= not (a and b);
    outputs(4364) <= not (a xor b);
    outputs(4365) <= not (a xor b);
    outputs(4366) <= a or b;
    outputs(4367) <= not a;
    outputs(4368) <= not (a xor b);
    outputs(4369) <= a or b;
    outputs(4370) <= b;
    outputs(4371) <= not (a or b);
    outputs(4372) <= not (a xor b);
    outputs(4373) <= a;
    outputs(4374) <= not a or b;
    outputs(4375) <= a xor b;
    outputs(4376) <= not a;
    outputs(4377) <= a xor b;
    outputs(4378) <= not (a xor b);
    outputs(4379) <= a or b;
    outputs(4380) <= a xor b;
    outputs(4381) <= a xor b;
    outputs(4382) <= not b;
    outputs(4383) <= not (a and b);
    outputs(4384) <= b;
    outputs(4385) <= a xor b;
    outputs(4386) <= not (a and b);
    outputs(4387) <= b;
    outputs(4388) <= a;
    outputs(4389) <= not b or a;
    outputs(4390) <= not b;
    outputs(4391) <= a or b;
    outputs(4392) <= not b;
    outputs(4393) <= not b;
    outputs(4394) <= a and b;
    outputs(4395) <= b;
    outputs(4396) <= not b;
    outputs(4397) <= 1'b1;
    outputs(4398) <= not a;
    outputs(4399) <= not b;
    outputs(4400) <= a or b;
    outputs(4401) <= not a;
    outputs(4402) <= not a;
    outputs(4403) <= not a or b;
    outputs(4404) <= not (a xor b);
    outputs(4405) <= not b or a;
    outputs(4406) <= not b;
    outputs(4407) <= a or b;
    outputs(4408) <= not a or b;
    outputs(4409) <= not (a xor b);
    outputs(4410) <= b;
    outputs(4411) <= b;
    outputs(4412) <= not (a or b);
    outputs(4413) <= not (a xor b);
    outputs(4414) <= a or b;
    outputs(4415) <= a xor b;
    outputs(4416) <= a xor b;
    outputs(4417) <= not a or b;
    outputs(4418) <= a or b;
    outputs(4419) <= a xor b;
    outputs(4420) <= not (a and b);
    outputs(4421) <= a;
    outputs(4422) <= not (a xor b);
    outputs(4423) <= not b;
    outputs(4424) <= not (a and b);
    outputs(4425) <= not (a xor b);
    outputs(4426) <= a xor b;
    outputs(4427) <= not a or b;
    outputs(4428) <= not b or a;
    outputs(4429) <= not (a and b);
    outputs(4430) <= a or b;
    outputs(4431) <= a xor b;
    outputs(4432) <= a and b;
    outputs(4433) <= not b;
    outputs(4434) <= not a;
    outputs(4435) <= not (a and b);
    outputs(4436) <= not (a xor b);
    outputs(4437) <= not (a and b);
    outputs(4438) <= not (a xor b);
    outputs(4439) <= a or b;
    outputs(4440) <= a and b;
    outputs(4441) <= not a;
    outputs(4442) <= not (a xor b);
    outputs(4443) <= not (a xor b);
    outputs(4444) <= not b or a;
    outputs(4445) <= a and b;
    outputs(4446) <= not (a and b);
    outputs(4447) <= not b or a;
    outputs(4448) <= a xor b;
    outputs(4449) <= not (a xor b);
    outputs(4450) <= not b or a;
    outputs(4451) <= not b;
    outputs(4452) <= b;
    outputs(4453) <= not a;
    outputs(4454) <= a and b;
    outputs(4455) <= b;
    outputs(4456) <= b;
    outputs(4457) <= not (a and b);
    outputs(4458) <= not a or b;
    outputs(4459) <= b;
    outputs(4460) <= a xor b;
    outputs(4461) <= not a;
    outputs(4462) <= a xor b;
    outputs(4463) <= a;
    outputs(4464) <= not (a and b);
    outputs(4465) <= not b;
    outputs(4466) <= a;
    outputs(4467) <= not b;
    outputs(4468) <= not (a and b);
    outputs(4469) <= b and not a;
    outputs(4470) <= not (a xor b);
    outputs(4471) <= not (a xor b);
    outputs(4472) <= not (a xor b);
    outputs(4473) <= a;
    outputs(4474) <= not (a xor b);
    outputs(4475) <= a xor b;
    outputs(4476) <= a;
    outputs(4477) <= not (a and b);
    outputs(4478) <= not a;
    outputs(4479) <= not (a xor b);
    outputs(4480) <= not a;
    outputs(4481) <= not (a and b);
    outputs(4482) <= not (a and b);
    outputs(4483) <= b and not a;
    outputs(4484) <= not (a xor b);
    outputs(4485) <= a xor b;
    outputs(4486) <= a or b;
    outputs(4487) <= not (a or b);
    outputs(4488) <= a xor b;
    outputs(4489) <= not b or a;
    outputs(4490) <= not b or a;
    outputs(4491) <= a xor b;
    outputs(4492) <= a xor b;
    outputs(4493) <= not b or a;
    outputs(4494) <= a or b;
    outputs(4495) <= not b or a;
    outputs(4496) <= not b;
    outputs(4497) <= not a;
    outputs(4498) <= not (a and b);
    outputs(4499) <= not (a xor b);
    outputs(4500) <= not (a and b);
    outputs(4501) <= not b;
    outputs(4502) <= not (a xor b);
    outputs(4503) <= a or b;
    outputs(4504) <= b and not a;
    outputs(4505) <= not b or a;
    outputs(4506) <= a xor b;
    outputs(4507) <= b;
    outputs(4508) <= b;
    outputs(4509) <= not a;
    outputs(4510) <= b;
    outputs(4511) <= not b or a;
    outputs(4512) <= a;
    outputs(4513) <= a;
    outputs(4514) <= not a;
    outputs(4515) <= not (a or b);
    outputs(4516) <= not (a or b);
    outputs(4517) <= not b;
    outputs(4518) <= a xor b;
    outputs(4519) <= not a or b;
    outputs(4520) <= not b;
    outputs(4521) <= not a;
    outputs(4522) <= not b;
    outputs(4523) <= not (a xor b);
    outputs(4524) <= a xor b;
    outputs(4525) <= not b or a;
    outputs(4526) <= not (a xor b);
    outputs(4527) <= not b or a;
    outputs(4528) <= b;
    outputs(4529) <= b;
    outputs(4530) <= not a;
    outputs(4531) <= not b;
    outputs(4532) <= a xor b;
    outputs(4533) <= a;
    outputs(4534) <= not (a xor b);
    outputs(4535) <= not (a and b);
    outputs(4536) <= not (a xor b);
    outputs(4537) <= a;
    outputs(4538) <= b;
    outputs(4539) <= b and not a;
    outputs(4540) <= not (a xor b);
    outputs(4541) <= a xor b;
    outputs(4542) <= not b or a;
    outputs(4543) <= not a;
    outputs(4544) <= not b or a;
    outputs(4545) <= a xor b;
    outputs(4546) <= a and not b;
    outputs(4547) <= not (a xor b);
    outputs(4548) <= b and not a;
    outputs(4549) <= a;
    outputs(4550) <= not a or b;
    outputs(4551) <= not (a or b);
    outputs(4552) <= not b or a;
    outputs(4553) <= not (a or b);
    outputs(4554) <= not a or b;
    outputs(4555) <= a;
    outputs(4556) <= b;
    outputs(4557) <= not (a and b);
    outputs(4558) <= not (a xor b);
    outputs(4559) <= a xor b;
    outputs(4560) <= not b;
    outputs(4561) <= a or b;
    outputs(4562) <= not (a or b);
    outputs(4563) <= a and b;
    outputs(4564) <= not b;
    outputs(4565) <= b;
    outputs(4566) <= a;
    outputs(4567) <= not (a xor b);
    outputs(4568) <= a or b;
    outputs(4569) <= b;
    outputs(4570) <= not a or b;
    outputs(4571) <= not a;
    outputs(4572) <= a or b;
    outputs(4573) <= b and not a;
    outputs(4574) <= not (a xor b);
    outputs(4575) <= not (a and b);
    outputs(4576) <= not (a or b);
    outputs(4577) <= a;
    outputs(4578) <= not b or a;
    outputs(4579) <= not (a xor b);
    outputs(4580) <= not a or b;
    outputs(4581) <= a and b;
    outputs(4582) <= a xor b;
    outputs(4583) <= not (a and b);
    outputs(4584) <= not a;
    outputs(4585) <= b;
    outputs(4586) <= a xor b;
    outputs(4587) <= a and not b;
    outputs(4588) <= a or b;
    outputs(4589) <= not (a and b);
    outputs(4590) <= not b;
    outputs(4591) <= a xor b;
    outputs(4592) <= not b or a;
    outputs(4593) <= a xor b;
    outputs(4594) <= a or b;
    outputs(4595) <= a xor b;
    outputs(4596) <= not a;
    outputs(4597) <= a and b;
    outputs(4598) <= a xor b;
    outputs(4599) <= not (a or b);
    outputs(4600) <= not b;
    outputs(4601) <= b;
    outputs(4602) <= not a;
    outputs(4603) <= b and not a;
    outputs(4604) <= not (a xor b);
    outputs(4605) <= not b;
    outputs(4606) <= a xor b;
    outputs(4607) <= b and not a;
    outputs(4608) <= a and not b;
    outputs(4609) <= not (a xor b);
    outputs(4610) <= not a;
    outputs(4611) <= a or b;
    outputs(4612) <= b and not a;
    outputs(4613) <= not b;
    outputs(4614) <= not (a xor b);
    outputs(4615) <= b;
    outputs(4616) <= a and not b;
    outputs(4617) <= a xor b;
    outputs(4618) <= a or b;
    outputs(4619) <= not a;
    outputs(4620) <= not (a xor b);
    outputs(4621) <= not (a xor b);
    outputs(4622) <= a;
    outputs(4623) <= not (a and b);
    outputs(4624) <= a xor b;
    outputs(4625) <= not (a xor b);
    outputs(4626) <= not b or a;
    outputs(4627) <= not (a and b);
    outputs(4628) <= not b or a;
    outputs(4629) <= not a;
    outputs(4630) <= b;
    outputs(4631) <= not (a xor b);
    outputs(4632) <= not b;
    outputs(4633) <= b;
    outputs(4634) <= not a or b;
    outputs(4635) <= a and b;
    outputs(4636) <= b and not a;
    outputs(4637) <= not (a xor b);
    outputs(4638) <= a or b;
    outputs(4639) <= not b or a;
    outputs(4640) <= b;
    outputs(4641) <= b and not a;
    outputs(4642) <= not b or a;
    outputs(4643) <= b and not a;
    outputs(4644) <= a xor b;
    outputs(4645) <= a;
    outputs(4646) <= b;
    outputs(4647) <= not a;
    outputs(4648) <= a or b;
    outputs(4649) <= not a;
    outputs(4650) <= a or b;
    outputs(4651) <= not b;
    outputs(4652) <= not (a xor b);
    outputs(4653) <= not (a and b);
    outputs(4654) <= not a;
    outputs(4655) <= not b or a;
    outputs(4656) <= b;
    outputs(4657) <= not (a or b);
    outputs(4658) <= a and b;
    outputs(4659) <= not a;
    outputs(4660) <= not b;
    outputs(4661) <= not b;
    outputs(4662) <= a and b;
    outputs(4663) <= b;
    outputs(4664) <= a;
    outputs(4665) <= a xor b;
    outputs(4666) <= not (a xor b);
    outputs(4667) <= a xor b;
    outputs(4668) <= not (a or b);
    outputs(4669) <= not b;
    outputs(4670) <= a;
    outputs(4671) <= not b or a;
    outputs(4672) <= not a or b;
    outputs(4673) <= not a;
    outputs(4674) <= a;
    outputs(4675) <= not (a xor b);
    outputs(4676) <= a;
    outputs(4677) <= not (a and b);
    outputs(4678) <= b;
    outputs(4679) <= a xor b;
    outputs(4680) <= not a;
    outputs(4681) <= not a;
    outputs(4682) <= a;
    outputs(4683) <= not a;
    outputs(4684) <= b;
    outputs(4685) <= a xor b;
    outputs(4686) <= a and not b;
    outputs(4687) <= not (a and b);
    outputs(4688) <= not (a xor b);
    outputs(4689) <= a or b;
    outputs(4690) <= b;
    outputs(4691) <= b;
    outputs(4692) <= b;
    outputs(4693) <= not a;
    outputs(4694) <= not (a xor b);
    outputs(4695) <= not (a or b);
    outputs(4696) <= not (a xor b);
    outputs(4697) <= a;
    outputs(4698) <= not (a xor b);
    outputs(4699) <= b;
    outputs(4700) <= a and b;
    outputs(4701) <= b;
    outputs(4702) <= not (a xor b);
    outputs(4703) <= not (a xor b);
    outputs(4704) <= a or b;
    outputs(4705) <= a;
    outputs(4706) <= not (a xor b);
    outputs(4707) <= b;
    outputs(4708) <= not b or a;
    outputs(4709) <= a and not b;
    outputs(4710) <= not b;
    outputs(4711) <= not (a xor b);
    outputs(4712) <= a xor b;
    outputs(4713) <= a;
    outputs(4714) <= a xor b;
    outputs(4715) <= not b;
    outputs(4716) <= a and b;
    outputs(4717) <= not (a xor b);
    outputs(4718) <= not b or a;
    outputs(4719) <= not (a xor b);
    outputs(4720) <= b;
    outputs(4721) <= a xor b;
    outputs(4722) <= a xor b;
    outputs(4723) <= not a or b;
    outputs(4724) <= b;
    outputs(4725) <= a;
    outputs(4726) <= not a;
    outputs(4727) <= not b or a;
    outputs(4728) <= a or b;
    outputs(4729) <= not (a or b);
    outputs(4730) <= a xor b;
    outputs(4731) <= b;
    outputs(4732) <= not (a xor b);
    outputs(4733) <= not a;
    outputs(4734) <= not (a xor b);
    outputs(4735) <= a or b;
    outputs(4736) <= b and not a;
    outputs(4737) <= not b or a;
    outputs(4738) <= not (a xor b);
    outputs(4739) <= not b or a;
    outputs(4740) <= a;
    outputs(4741) <= not (a and b);
    outputs(4742) <= b;
    outputs(4743) <= not b;
    outputs(4744) <= a xor b;
    outputs(4745) <= a and b;
    outputs(4746) <= b;
    outputs(4747) <= a xor b;
    outputs(4748) <= not b;
    outputs(4749) <= b;
    outputs(4750) <= not a or b;
    outputs(4751) <= not (a and b);
    outputs(4752) <= b;
    outputs(4753) <= a;
    outputs(4754) <= a xor b;
    outputs(4755) <= a;
    outputs(4756) <= not a or b;
    outputs(4757) <= a and not b;
    outputs(4758) <= b;
    outputs(4759) <= a;
    outputs(4760) <= not (a and b);
    outputs(4761) <= not b or a;
    outputs(4762) <= a and not b;
    outputs(4763) <= a xor b;
    outputs(4764) <= not (a and b);
    outputs(4765) <= not b or a;
    outputs(4766) <= not (a xor b);
    outputs(4767) <= not (a xor b);
    outputs(4768) <= a xor b;
    outputs(4769) <= not a;
    outputs(4770) <= not (a and b);
    outputs(4771) <= not (a and b);
    outputs(4772) <= a xor b;
    outputs(4773) <= not b;
    outputs(4774) <= not a;
    outputs(4775) <= not (a xor b);
    outputs(4776) <= not b or a;
    outputs(4777) <= b;
    outputs(4778) <= not (a and b);
    outputs(4779) <= not b;
    outputs(4780) <= not a;
    outputs(4781) <= not (a xor b);
    outputs(4782) <= not (a xor b);
    outputs(4783) <= not b;
    outputs(4784) <= not b;
    outputs(4785) <= not (a xor b);
    outputs(4786) <= not (a xor b);
    outputs(4787) <= a;
    outputs(4788) <= not a;
    outputs(4789) <= not a;
    outputs(4790) <= a and b;
    outputs(4791) <= a;
    outputs(4792) <= not a or b;
    outputs(4793) <= not (a and b);
    outputs(4794) <= b;
    outputs(4795) <= b;
    outputs(4796) <= not b or a;
    outputs(4797) <= a;
    outputs(4798) <= b and not a;
    outputs(4799) <= a xor b;
    outputs(4800) <= not b;
    outputs(4801) <= not b;
    outputs(4802) <= not (a xor b);
    outputs(4803) <= a or b;
    outputs(4804) <= a and not b;
    outputs(4805) <= a and not b;
    outputs(4806) <= a xor b;
    outputs(4807) <= not (a or b);
    outputs(4808) <= b;
    outputs(4809) <= b;
    outputs(4810) <= not b;
    outputs(4811) <= not (a xor b);
    outputs(4812) <= b;
    outputs(4813) <= a or b;
    outputs(4814) <= a xor b;
    outputs(4815) <= not b;
    outputs(4816) <= b and not a;
    outputs(4817) <= not a;
    outputs(4818) <= not a or b;
    outputs(4819) <= not a;
    outputs(4820) <= not b or a;
    outputs(4821) <= not a or b;
    outputs(4822) <= not (a or b);
    outputs(4823) <= a;
    outputs(4824) <= a;
    outputs(4825) <= b;
    outputs(4826) <= not b or a;
    outputs(4827) <= a xor b;
    outputs(4828) <= not b or a;
    outputs(4829) <= a xor b;
    outputs(4830) <= not b;
    outputs(4831) <= a and b;
    outputs(4832) <= a xor b;
    outputs(4833) <= not (a xor b);
    outputs(4834) <= a or b;
    outputs(4835) <= not (a xor b);
    outputs(4836) <= a xor b;
    outputs(4837) <= not b;
    outputs(4838) <= a;
    outputs(4839) <= a;
    outputs(4840) <= a xor b;
    outputs(4841) <= a;
    outputs(4842) <= b;
    outputs(4843) <= not b;
    outputs(4844) <= not (a xor b);
    outputs(4845) <= not b or a;
    outputs(4846) <= a;
    outputs(4847) <= a or b;
    outputs(4848) <= b;
    outputs(4849) <= not a or b;
    outputs(4850) <= not b;
    outputs(4851) <= not (a xor b);
    outputs(4852) <= a;
    outputs(4853) <= a and not b;
    outputs(4854) <= not (a xor b);
    outputs(4855) <= a xor b;
    outputs(4856) <= not a;
    outputs(4857) <= not (a xor b);
    outputs(4858) <= not a;
    outputs(4859) <= not (a xor b);
    outputs(4860) <= a and not b;
    outputs(4861) <= a and b;
    outputs(4862) <= not (a and b);
    outputs(4863) <= b;
    outputs(4864) <= not a;
    outputs(4865) <= not (a xor b);
    outputs(4866) <= a xor b;
    outputs(4867) <= a xor b;
    outputs(4868) <= not a;
    outputs(4869) <= not (a or b);
    outputs(4870) <= not (a or b);
    outputs(4871) <= a xor b;
    outputs(4872) <= a and not b;
    outputs(4873) <= a xor b;
    outputs(4874) <= a;
    outputs(4875) <= not b;
    outputs(4876) <= a;
    outputs(4877) <= b;
    outputs(4878) <= a xor b;
    outputs(4879) <= not (a and b);
    outputs(4880) <= not a;
    outputs(4881) <= not (a xor b);
    outputs(4882) <= b and not a;
    outputs(4883) <= not b;
    outputs(4884) <= a xor b;
    outputs(4885) <= b;
    outputs(4886) <= not b or a;
    outputs(4887) <= b;
    outputs(4888) <= not (a or b);
    outputs(4889) <= not (a xor b);
    outputs(4890) <= not a or b;
    outputs(4891) <= a;
    outputs(4892) <= not (a xor b);
    outputs(4893) <= not a or b;
    outputs(4894) <= not a or b;
    outputs(4895) <= a xor b;
    outputs(4896) <= not (a xor b);
    outputs(4897) <= not a;
    outputs(4898) <= a and not b;
    outputs(4899) <= a;
    outputs(4900) <= a xor b;
    outputs(4901) <= not (a or b);
    outputs(4902) <= b;
    outputs(4903) <= a or b;
    outputs(4904) <= a;
    outputs(4905) <= not (a and b);
    outputs(4906) <= not b or a;
    outputs(4907) <= b;
    outputs(4908) <= not (a xor b);
    outputs(4909) <= a;
    outputs(4910) <= not (a xor b);
    outputs(4911) <= not b;
    outputs(4912) <= b and not a;
    outputs(4913) <= b and not a;
    outputs(4914) <= not (a xor b);
    outputs(4915) <= a xor b;
    outputs(4916) <= not (a and b);
    outputs(4917) <= not (a xor b);
    outputs(4918) <= not a or b;
    outputs(4919) <= a xor b;
    outputs(4920) <= not a;
    outputs(4921) <= not b;
    outputs(4922) <= not b;
    outputs(4923) <= a;
    outputs(4924) <= a and b;
    outputs(4925) <= not a;
    outputs(4926) <= not a;
    outputs(4927) <= b and not a;
    outputs(4928) <= b;
    outputs(4929) <= not (a xor b);
    outputs(4930) <= a xor b;
    outputs(4931) <= b;
    outputs(4932) <= a;
    outputs(4933) <= a and not b;
    outputs(4934) <= not (a or b);
    outputs(4935) <= a and not b;
    outputs(4936) <= not (a xor b);
    outputs(4937) <= not (a xor b);
    outputs(4938) <= not b or a;
    outputs(4939) <= a xor b;
    outputs(4940) <= not a or b;
    outputs(4941) <= not b;
    outputs(4942) <= not a;
    outputs(4943) <= a;
    outputs(4944) <= b;
    outputs(4945) <= a and not b;
    outputs(4946) <= b;
    outputs(4947) <= b;
    outputs(4948) <= a or b;
    outputs(4949) <= a xor b;
    outputs(4950) <= not (a xor b);
    outputs(4951) <= a or b;
    outputs(4952) <= not a;
    outputs(4953) <= not (a or b);
    outputs(4954) <= not (a xor b);
    outputs(4955) <= b;
    outputs(4956) <= a xor b;
    outputs(4957) <= a;
    outputs(4958) <= not b or a;
    outputs(4959) <= not (a or b);
    outputs(4960) <= not (a xor b);
    outputs(4961) <= not (a xor b);
    outputs(4962) <= not (a and b);
    outputs(4963) <= a;
    outputs(4964) <= not b or a;
    outputs(4965) <= not a;
    outputs(4966) <= a;
    outputs(4967) <= a;
    outputs(4968) <= not (a or b);
    outputs(4969) <= a and b;
    outputs(4970) <= not b;
    outputs(4971) <= a or b;
    outputs(4972) <= b;
    outputs(4973) <= a xor b;
    outputs(4974) <= not (a and b);
    outputs(4975) <= not a;
    outputs(4976) <= not (a and b);
    outputs(4977) <= not (a xor b);
    outputs(4978) <= a xor b;
    outputs(4979) <= a or b;
    outputs(4980) <= not (a or b);
    outputs(4981) <= not (a xor b);
    outputs(4982) <= a and not b;
    outputs(4983) <= a xor b;
    outputs(4984) <= not b or a;
    outputs(4985) <= a;
    outputs(4986) <= a or b;
    outputs(4987) <= not a;
    outputs(4988) <= a;
    outputs(4989) <= a;
    outputs(4990) <= a xor b;
    outputs(4991) <= not (a xor b);
    outputs(4992) <= not b;
    outputs(4993) <= not b;
    outputs(4994) <= b;
    outputs(4995) <= not (a xor b);
    outputs(4996) <= a or b;
    outputs(4997) <= a xor b;
    outputs(4998) <= not b;
    outputs(4999) <= not a;
    outputs(5000) <= b;
    outputs(5001) <= not (a or b);
    outputs(5002) <= not a or b;
    outputs(5003) <= b;
    outputs(5004) <= not a or b;
    outputs(5005) <= not (a and b);
    outputs(5006) <= not (a xor b);
    outputs(5007) <= not a;
    outputs(5008) <= a and not b;
    outputs(5009) <= b;
    outputs(5010) <= not b or a;
    outputs(5011) <= not a;
    outputs(5012) <= not a;
    outputs(5013) <= b and not a;
    outputs(5014) <= a;
    outputs(5015) <= not a;
    outputs(5016) <= b and not a;
    outputs(5017) <= a and not b;
    outputs(5018) <= a or b;
    outputs(5019) <= b and not a;
    outputs(5020) <= not b;
    outputs(5021) <= not (a xor b);
    outputs(5022) <= b and not a;
    outputs(5023) <= a xor b;
    outputs(5024) <= not (a xor b);
    outputs(5025) <= not b;
    outputs(5026) <= not (a and b);
    outputs(5027) <= not a;
    outputs(5028) <= not (a xor b);
    outputs(5029) <= a xor b;
    outputs(5030) <= not (a or b);
    outputs(5031) <= a or b;
    outputs(5032) <= a;
    outputs(5033) <= a xor b;
    outputs(5034) <= not a;
    outputs(5035) <= a;
    outputs(5036) <= a or b;
    outputs(5037) <= not a;
    outputs(5038) <= not a;
    outputs(5039) <= b;
    outputs(5040) <= not (a xor b);
    outputs(5041) <= a xor b;
    outputs(5042) <= a;
    outputs(5043) <= not b;
    outputs(5044) <= not a;
    outputs(5045) <= a xor b;
    outputs(5046) <= not a;
    outputs(5047) <= not b or a;
    outputs(5048) <= a or b;
    outputs(5049) <= a xor b;
    outputs(5050) <= a xor b;
    outputs(5051) <= not b;
    outputs(5052) <= not (a xor b);
    outputs(5053) <= not a;
    outputs(5054) <= not (a or b);
    outputs(5055) <= not b or a;
    outputs(5056) <= a;
    outputs(5057) <= not (a and b);
    outputs(5058) <= a;
    outputs(5059) <= not a;
    outputs(5060) <= a and b;
    outputs(5061) <= not b;
    outputs(5062) <= b and not a;
    outputs(5063) <= not b;
    outputs(5064) <= a and not b;
    outputs(5065) <= not a;
    outputs(5066) <= b and not a;
    outputs(5067) <= a or b;
    outputs(5068) <= not b or a;
    outputs(5069) <= b;
    outputs(5070) <= not a;
    outputs(5071) <= not a or b;
    outputs(5072) <= not (a and b);
    outputs(5073) <= b;
    outputs(5074) <= a or b;
    outputs(5075) <= not (a xor b);
    outputs(5076) <= b;
    outputs(5077) <= not (a xor b);
    outputs(5078) <= not (a and b);
    outputs(5079) <= not (a xor b);
    outputs(5080) <= b and not a;
    outputs(5081) <= not (a xor b);
    outputs(5082) <= not (a xor b);
    outputs(5083) <= not b or a;
    outputs(5084) <= not b or a;
    outputs(5085) <= not (a xor b);
    outputs(5086) <= not a;
    outputs(5087) <= a xor b;
    outputs(5088) <= not b;
    outputs(5089) <= a xor b;
    outputs(5090) <= a xor b;
    outputs(5091) <= not (a xor b);
    outputs(5092) <= not b;
    outputs(5093) <= b;
    outputs(5094) <= a xor b;
    outputs(5095) <= a or b;
    outputs(5096) <= not b;
    outputs(5097) <= not (a xor b);
    outputs(5098) <= not b or a;
    outputs(5099) <= not (a xor b);
    outputs(5100) <= a xor b;
    outputs(5101) <= not (a and b);
    outputs(5102) <= not b or a;
    outputs(5103) <= not b;
    outputs(5104) <= a xor b;
    outputs(5105) <= a xor b;
    outputs(5106) <= a xor b;
    outputs(5107) <= a and not b;
    outputs(5108) <= not b;
    outputs(5109) <= not a;
    outputs(5110) <= a xor b;
    outputs(5111) <= b and not a;
    outputs(5112) <= not (a or b);
    outputs(5113) <= a xor b;
    outputs(5114) <= a xor b;
    outputs(5115) <= b;
    outputs(5116) <= b;
    outputs(5117) <= not b;
    outputs(5118) <= a xor b;
    outputs(5119) <= not b or a;
    outputs(5120) <= a and b;
    outputs(5121) <= not (a or b);
    outputs(5122) <= not a;
    outputs(5123) <= not (a or b);
    outputs(5124) <= not (a or b);
    outputs(5125) <= not (a or b);
    outputs(5126) <= not (a or b);
    outputs(5127) <= b;
    outputs(5128) <= b;
    outputs(5129) <= a;
    outputs(5130) <= not (a or b);
    outputs(5131) <= a;
    outputs(5132) <= not (a xor b);
    outputs(5133) <= not b;
    outputs(5134) <= a and b;
    outputs(5135) <= a xor b;
    outputs(5136) <= not (a xor b);
    outputs(5137) <= b and not a;
    outputs(5138) <= not a or b;
    outputs(5139) <= a;
    outputs(5140) <= a;
    outputs(5141) <= a xor b;
    outputs(5142) <= not (a xor b);
    outputs(5143) <= not b;
    outputs(5144) <= a xor b;
    outputs(5145) <= not (a xor b);
    outputs(5146) <= b and not a;
    outputs(5147) <= not b;
    outputs(5148) <= not (a or b);
    outputs(5149) <= a xor b;
    outputs(5150) <= b;
    outputs(5151) <= a;
    outputs(5152) <= not (a and b);
    outputs(5153) <= a xor b;
    outputs(5154) <= a and b;
    outputs(5155) <= b and not a;
    outputs(5156) <= not (a xor b);
    outputs(5157) <= a xor b;
    outputs(5158) <= a;
    outputs(5159) <= not (a xor b);
    outputs(5160) <= not b or a;
    outputs(5161) <= a or b;
    outputs(5162) <= not a;
    outputs(5163) <= not (a xor b);
    outputs(5164) <= b;
    outputs(5165) <= a xor b;
    outputs(5166) <= a and b;
    outputs(5167) <= a;
    outputs(5168) <= not a or b;
    outputs(5169) <= b;
    outputs(5170) <= b and not a;
    outputs(5171) <= not (a xor b);
    outputs(5172) <= b;
    outputs(5173) <= b and not a;
    outputs(5174) <= a;
    outputs(5175) <= not b;
    outputs(5176) <= not b;
    outputs(5177) <= not b;
    outputs(5178) <= b and not a;
    outputs(5179) <= b;
    outputs(5180) <= a and not b;
    outputs(5181) <= not a or b;
    outputs(5182) <= not (a or b);
    outputs(5183) <= b and not a;
    outputs(5184) <= not b;
    outputs(5185) <= a xor b;
    outputs(5186) <= b;
    outputs(5187) <= not (a xor b);
    outputs(5188) <= b and not a;
    outputs(5189) <= b and not a;
    outputs(5190) <= b and not a;
    outputs(5191) <= a and b;
    outputs(5192) <= a;
    outputs(5193) <= not a;
    outputs(5194) <= a and not b;
    outputs(5195) <= a and not b;
    outputs(5196) <= a xor b;
    outputs(5197) <= not (a xor b);
    outputs(5198) <= a;
    outputs(5199) <= not (a xor b);
    outputs(5200) <= not (a xor b);
    outputs(5201) <= not a;
    outputs(5202) <= a and b;
    outputs(5203) <= 1'b0;
    outputs(5204) <= b;
    outputs(5205) <= a xor b;
    outputs(5206) <= a and not b;
    outputs(5207) <= a xor b;
    outputs(5208) <= not (a xor b);
    outputs(5209) <= not b;
    outputs(5210) <= b;
    outputs(5211) <= b and not a;
    outputs(5212) <= a and b;
    outputs(5213) <= a and not b;
    outputs(5214) <= not b;
    outputs(5215) <= b;
    outputs(5216) <= not (a or b);
    outputs(5217) <= a and not b;
    outputs(5218) <= not (a xor b);
    outputs(5219) <= not a;
    outputs(5220) <= not a;
    outputs(5221) <= a;
    outputs(5222) <= not (a or b);
    outputs(5223) <= not (a xor b);
    outputs(5224) <= a;
    outputs(5225) <= a;
    outputs(5226) <= a and b;
    outputs(5227) <= a xor b;
    outputs(5228) <= not b;
    outputs(5229) <= not a;
    outputs(5230) <= a or b;
    outputs(5231) <= a and not b;
    outputs(5232) <= a xor b;
    outputs(5233) <= not b;
    outputs(5234) <= 1'b0;
    outputs(5235) <= a;
    outputs(5236) <= a and b;
    outputs(5237) <= not a or b;
    outputs(5238) <= b;
    outputs(5239) <= not (a xor b);
    outputs(5240) <= a and b;
    outputs(5241) <= not a;
    outputs(5242) <= b;
    outputs(5243) <= not b;
    outputs(5244) <= not a or b;
    outputs(5245) <= not b;
    outputs(5246) <= not (a or b);
    outputs(5247) <= not (a xor b);
    outputs(5248) <= a and b;
    outputs(5249) <= a and not b;
    outputs(5250) <= a;
    outputs(5251) <= not b;
    outputs(5252) <= a and not b;
    outputs(5253) <= not (a or b);
    outputs(5254) <= not (a xor b);
    outputs(5255) <= a xor b;
    outputs(5256) <= a and b;
    outputs(5257) <= a xor b;
    outputs(5258) <= a and b;
    outputs(5259) <= b and not a;
    outputs(5260) <= b;
    outputs(5261) <= b and not a;
    outputs(5262) <= a and b;
    outputs(5263) <= a and not b;
    outputs(5264) <= not b;
    outputs(5265) <= not a;
    outputs(5266) <= a or b;
    outputs(5267) <= a;
    outputs(5268) <= not b;
    outputs(5269) <= not (a xor b);
    outputs(5270) <= b;
    outputs(5271) <= not (a xor b);
    outputs(5272) <= b and not a;
    outputs(5273) <= a and b;
    outputs(5274) <= a and not b;
    outputs(5275) <= a and not b;
    outputs(5276) <= not b;
    outputs(5277) <= b;
    outputs(5278) <= not a;
    outputs(5279) <= not b;
    outputs(5280) <= not a;
    outputs(5281) <= b and not a;
    outputs(5282) <= a xor b;
    outputs(5283) <= b and not a;
    outputs(5284) <= not (a or b);
    outputs(5285) <= a and not b;
    outputs(5286) <= b and not a;
    outputs(5287) <= a;
    outputs(5288) <= not (a xor b);
    outputs(5289) <= not a;
    outputs(5290) <= b;
    outputs(5291) <= a;
    outputs(5292) <= a and b;
    outputs(5293) <= a xor b;
    outputs(5294) <= a and b;
    outputs(5295) <= a xor b;
    outputs(5296) <= not a;
    outputs(5297) <= not (a xor b);
    outputs(5298) <= not (a and b);
    outputs(5299) <= a;
    outputs(5300) <= not a or b;
    outputs(5301) <= b;
    outputs(5302) <= a;
    outputs(5303) <= a;
    outputs(5304) <= a;
    outputs(5305) <= a or b;
    outputs(5306) <= b and not a;
    outputs(5307) <= not a;
    outputs(5308) <= a xor b;
    outputs(5309) <= not a;
    outputs(5310) <= not (a or b);
    outputs(5311) <= not (a or b);
    outputs(5312) <= not (a xor b);
    outputs(5313) <= not a;
    outputs(5314) <= not (a or b);
    outputs(5315) <= a xor b;
    outputs(5316) <= a;
    outputs(5317) <= a xor b;
    outputs(5318) <= a and b;
    outputs(5319) <= a and not b;
    outputs(5320) <= not (a xor b);
    outputs(5321) <= a and b;
    outputs(5322) <= b and not a;
    outputs(5323) <= a xor b;
    outputs(5324) <= not a;
    outputs(5325) <= not b;
    outputs(5326) <= b and not a;
    outputs(5327) <= b;
    outputs(5328) <= not b;
    outputs(5329) <= b;
    outputs(5330) <= a;
    outputs(5331) <= not (a xor b);
    outputs(5332) <= not (a or b);
    outputs(5333) <= not a;
    outputs(5334) <= a and b;
    outputs(5335) <= b and not a;
    outputs(5336) <= a and not b;
    outputs(5337) <= not a;
    outputs(5338) <= b;
    outputs(5339) <= not a;
    outputs(5340) <= not a;
    outputs(5341) <= not b;
    outputs(5342) <= 1'b0;
    outputs(5343) <= a and b;
    outputs(5344) <= not b;
    outputs(5345) <= a;
    outputs(5346) <= not (a xor b);
    outputs(5347) <= a and not b;
    outputs(5348) <= a and not b;
    outputs(5349) <= not b or a;
    outputs(5350) <= a and not b;
    outputs(5351) <= a and not b;
    outputs(5352) <= a xor b;
    outputs(5353) <= not b;
    outputs(5354) <= a and not b;
    outputs(5355) <= b;
    outputs(5356) <= b;
    outputs(5357) <= a xor b;
    outputs(5358) <= not (a or b);
    outputs(5359) <= not b or a;
    outputs(5360) <= a xor b;
    outputs(5361) <= a and b;
    outputs(5362) <= not (a or b);
    outputs(5363) <= not a;
    outputs(5364) <= not (a and b);
    outputs(5365) <= a;
    outputs(5366) <= a and not b;
    outputs(5367) <= b and not a;
    outputs(5368) <= a and not b;
    outputs(5369) <= b and not a;
    outputs(5370) <= not b;
    outputs(5371) <= not a;
    outputs(5372) <= a and b;
    outputs(5373) <= a and b;
    outputs(5374) <= not a;
    outputs(5375) <= a and not b;
    outputs(5376) <= a and b;
    outputs(5377) <= a;
    outputs(5378) <= a;
    outputs(5379) <= not a or b;
    outputs(5380) <= not (a xor b);
    outputs(5381) <= a xor b;
    outputs(5382) <= a and not b;
    outputs(5383) <= not b;
    outputs(5384) <= not (a xor b);
    outputs(5385) <= a xor b;
    outputs(5386) <= b;
    outputs(5387) <= not b;
    outputs(5388) <= a;
    outputs(5389) <= not (a or b);
    outputs(5390) <= not a or b;
    outputs(5391) <= a and b;
    outputs(5392) <= a;
    outputs(5393) <= a and not b;
    outputs(5394) <= not (a xor b);
    outputs(5395) <= not (a xor b);
    outputs(5396) <= a and not b;
    outputs(5397) <= a or b;
    outputs(5398) <= not (a xor b);
    outputs(5399) <= a xor b;
    outputs(5400) <= b and not a;
    outputs(5401) <= not b;
    outputs(5402) <= not b;
    outputs(5403) <= not (a xor b);
    outputs(5404) <= a and b;
    outputs(5405) <= a;
    outputs(5406) <= a xor b;
    outputs(5407) <= not b;
    outputs(5408) <= a xor b;
    outputs(5409) <= a xor b;
    outputs(5410) <= a and b;
    outputs(5411) <= a;
    outputs(5412) <= not (a xor b);
    outputs(5413) <= a and not b;
    outputs(5414) <= not (a or b);
    outputs(5415) <= b and not a;
    outputs(5416) <= a xor b;
    outputs(5417) <= a;
    outputs(5418) <= not a;
    outputs(5419) <= not b or a;
    outputs(5420) <= a;
    outputs(5421) <= not (a xor b);
    outputs(5422) <= a and b;
    outputs(5423) <= a and not b;
    outputs(5424) <= a;
    outputs(5425) <= not a;
    outputs(5426) <= not b;
    outputs(5427) <= not (a xor b);
    outputs(5428) <= not b;
    outputs(5429) <= a;
    outputs(5430) <= b and not a;
    outputs(5431) <= a or b;
    outputs(5432) <= a or b;
    outputs(5433) <= b;
    outputs(5434) <= a;
    outputs(5435) <= a and b;
    outputs(5436) <= a xor b;
    outputs(5437) <= b and not a;
    outputs(5438) <= not a;
    outputs(5439) <= a;
    outputs(5440) <= not (a xor b);
    outputs(5441) <= not (a xor b);
    outputs(5442) <= b and not a;
    outputs(5443) <= not (a xor b);
    outputs(5444) <= a and b;
    outputs(5445) <= a;
    outputs(5446) <= not (a or b);
    outputs(5447) <= a and not b;
    outputs(5448) <= a and not b;
    outputs(5449) <= not (a or b);
    outputs(5450) <= b and not a;
    outputs(5451) <= not a;
    outputs(5452) <= not b;
    outputs(5453) <= a xor b;
    outputs(5454) <= not b;
    outputs(5455) <= not (a xor b);
    outputs(5456) <= not (a xor b);
    outputs(5457) <= a xor b;
    outputs(5458) <= b;
    outputs(5459) <= not (a xor b);
    outputs(5460) <= a xor b;
    outputs(5461) <= a;
    outputs(5462) <= not a or b;
    outputs(5463) <= a xor b;
    outputs(5464) <= a and not b;
    outputs(5465) <= not (a xor b);
    outputs(5466) <= a and not b;
    outputs(5467) <= not b;
    outputs(5468) <= b;
    outputs(5469) <= b and not a;
    outputs(5470) <= a and not b;
    outputs(5471) <= not (a xor b);
    outputs(5472) <= a;
    outputs(5473) <= not b;
    outputs(5474) <= a and not b;
    outputs(5475) <= a;
    outputs(5476) <= a and b;
    outputs(5477) <= 1'b0;
    outputs(5478) <= a;
    outputs(5479) <= a xor b;
    outputs(5480) <= b;
    outputs(5481) <= a xor b;
    outputs(5482) <= a xor b;
    outputs(5483) <= a xor b;
    outputs(5484) <= not a or b;
    outputs(5485) <= b;
    outputs(5486) <= a xor b;
    outputs(5487) <= a;
    outputs(5488) <= not a;
    outputs(5489) <= not (a or b);
    outputs(5490) <= a and not b;
    outputs(5491) <= a and b;
    outputs(5492) <= a and not b;
    outputs(5493) <= not (a or b);
    outputs(5494) <= b;
    outputs(5495) <= not (a and b);
    outputs(5496) <= not (a or b);
    outputs(5497) <= a xor b;
    outputs(5498) <= a and not b;
    outputs(5499) <= not a;
    outputs(5500) <= not (a xor b);
    outputs(5501) <= not a;
    outputs(5502) <= a;
    outputs(5503) <= not (a and b);
    outputs(5504) <= a and b;
    outputs(5505) <= b and not a;
    outputs(5506) <= a and not b;
    outputs(5507) <= a and not b;
    outputs(5508) <= not (a xor b);
    outputs(5509) <= not (a or b);
    outputs(5510) <= a and b;
    outputs(5511) <= not (a xor b);
    outputs(5512) <= not (a or b);
    outputs(5513) <= a;
    outputs(5514) <= not (a or b);
    outputs(5515) <= not b or a;
    outputs(5516) <= not a;
    outputs(5517) <= b and not a;
    outputs(5518) <= a;
    outputs(5519) <= not (a xor b);
    outputs(5520) <= not a;
    outputs(5521) <= a xor b;
    outputs(5522) <= not (a or b);
    outputs(5523) <= not b;
    outputs(5524) <= b;
    outputs(5525) <= a or b;
    outputs(5526) <= a xor b;
    outputs(5527) <= a and not b;
    outputs(5528) <= not b;
    outputs(5529) <= not (a xor b);
    outputs(5530) <= a and not b;
    outputs(5531) <= not a;
    outputs(5532) <= a;
    outputs(5533) <= b and not a;
    outputs(5534) <= a;
    outputs(5535) <= not (a and b);
    outputs(5536) <= b;
    outputs(5537) <= not b;
    outputs(5538) <= a and not b;
    outputs(5539) <= b;
    outputs(5540) <= a xor b;
    outputs(5541) <= a and b;
    outputs(5542) <= a and b;
    outputs(5543) <= not b;
    outputs(5544) <= a;
    outputs(5545) <= a and b;
    outputs(5546) <= not (a or b);
    outputs(5547) <= b and not a;
    outputs(5548) <= not (a and b);
    outputs(5549) <= not (a xor b);
    outputs(5550) <= a;
    outputs(5551) <= a xor b;
    outputs(5552) <= not (a xor b);
    outputs(5553) <= a and b;
    outputs(5554) <= a;
    outputs(5555) <= not a;
    outputs(5556) <= not (a or b);
    outputs(5557) <= a and not b;
    outputs(5558) <= a and b;
    outputs(5559) <= a xor b;
    outputs(5560) <= not b;
    outputs(5561) <= not (a xor b);
    outputs(5562) <= b and not a;
    outputs(5563) <= not (a xor b);
    outputs(5564) <= a and not b;
    outputs(5565) <= b;
    outputs(5566) <= not (a xor b);
    outputs(5567) <= not (a or b);
    outputs(5568) <= not a or b;
    outputs(5569) <= a and not b;
    outputs(5570) <= b;
    outputs(5571) <= b and not a;
    outputs(5572) <= b and not a;
    outputs(5573) <= not a;
    outputs(5574) <= not (a or b);
    outputs(5575) <= not a or b;
    outputs(5576) <= not b;
    outputs(5577) <= a xor b;
    outputs(5578) <= not (a xor b);
    outputs(5579) <= a and not b;
    outputs(5580) <= not b;
    outputs(5581) <= not (a xor b);
    outputs(5582) <= not a;
    outputs(5583) <= not b or a;
    outputs(5584) <= a and not b;
    outputs(5585) <= a and b;
    outputs(5586) <= a;
    outputs(5587) <= a or b;
    outputs(5588) <= a and b;
    outputs(5589) <= a xor b;
    outputs(5590) <= b and not a;
    outputs(5591) <= not a;
    outputs(5592) <= not a;
    outputs(5593) <= a and b;
    outputs(5594) <= a xor b;
    outputs(5595) <= b;
    outputs(5596) <= b;
    outputs(5597) <= not b;
    outputs(5598) <= not b;
    outputs(5599) <= a xor b;
    outputs(5600) <= not b;
    outputs(5601) <= not a;
    outputs(5602) <= a and b;
    outputs(5603) <= not a;
    outputs(5604) <= a;
    outputs(5605) <= a and not b;
    outputs(5606) <= not b;
    outputs(5607) <= a and not b;
    outputs(5608) <= not a;
    outputs(5609) <= a;
    outputs(5610) <= a and b;
    outputs(5611) <= b;
    outputs(5612) <= not a;
    outputs(5613) <= not b;
    outputs(5614) <= not (a xor b);
    outputs(5615) <= a xor b;
    outputs(5616) <= b;
    outputs(5617) <= a;
    outputs(5618) <= a xor b;
    outputs(5619) <= not (a xor b);
    outputs(5620) <= not (a xor b);
    outputs(5621) <= a xor b;
    outputs(5622) <= not (a or b);
    outputs(5623) <= a and b;
    outputs(5624) <= a and not b;
    outputs(5625) <= not (a xor b);
    outputs(5626) <= b;
    outputs(5627) <= a and not b;
    outputs(5628) <= not a;
    outputs(5629) <= not (a xor b);
    outputs(5630) <= b and not a;
    outputs(5631) <= b;
    outputs(5632) <= a or b;
    outputs(5633) <= not (a and b);
    outputs(5634) <= not (a or b);
    outputs(5635) <= a and not b;
    outputs(5636) <= not b or a;
    outputs(5637) <= not a;
    outputs(5638) <= not (a xor b);
    outputs(5639) <= a xor b;
    outputs(5640) <= b and not a;
    outputs(5641) <= b and not a;
    outputs(5642) <= a xor b;
    outputs(5643) <= not b or a;
    outputs(5644) <= a and b;
    outputs(5645) <= not b;
    outputs(5646) <= not b;
    outputs(5647) <= a xor b;
    outputs(5648) <= a;
    outputs(5649) <= a;
    outputs(5650) <= a xor b;
    outputs(5651) <= a;
    outputs(5652) <= not a;
    outputs(5653) <= b and not a;
    outputs(5654) <= a;
    outputs(5655) <= a;
    outputs(5656) <= a and not b;
    outputs(5657) <= not (a and b);
    outputs(5658) <= not b;
    outputs(5659) <= not b;
    outputs(5660) <= b and not a;
    outputs(5661) <= b and not a;
    outputs(5662) <= a and not b;
    outputs(5663) <= a and b;
    outputs(5664) <= a xor b;
    outputs(5665) <= not (a xor b);
    outputs(5666) <= 1'b0;
    outputs(5667) <= not b;
    outputs(5668) <= a xor b;
    outputs(5669) <= not (a or b);
    outputs(5670) <= a;
    outputs(5671) <= not (a or b);
    outputs(5672) <= a and b;
    outputs(5673) <= a and not b;
    outputs(5674) <= b and not a;
    outputs(5675) <= b and not a;
    outputs(5676) <= not (a or b);
    outputs(5677) <= not a;
    outputs(5678) <= not (a or b);
    outputs(5679) <= a and b;
    outputs(5680) <= not (a xor b);
    outputs(5681) <= a and b;
    outputs(5682) <= a xor b;
    outputs(5683) <= not b;
    outputs(5684) <= a and b;
    outputs(5685) <= not (a xor b);
    outputs(5686) <= not (a xor b);
    outputs(5687) <= not (a or b);
    outputs(5688) <= not a;
    outputs(5689) <= not (a or b);
    outputs(5690) <= a and not b;
    outputs(5691) <= a and b;
    outputs(5692) <= not a;
    outputs(5693) <= a xor b;
    outputs(5694) <= b;
    outputs(5695) <= b;
    outputs(5696) <= a and not b;
    outputs(5697) <= a and b;
    outputs(5698) <= b and not a;
    outputs(5699) <= b and not a;
    outputs(5700) <= a xor b;
    outputs(5701) <= a xor b;
    outputs(5702) <= not (a xor b);
    outputs(5703) <= a or b;
    outputs(5704) <= b and not a;
    outputs(5705) <= not a;
    outputs(5706) <= not (a and b);
    outputs(5707) <= a and b;
    outputs(5708) <= a and b;
    outputs(5709) <= a xor b;
    outputs(5710) <= a and not b;
    outputs(5711) <= b and not a;
    outputs(5712) <= not (a or b);
    outputs(5713) <= a xor b;
    outputs(5714) <= not b;
    outputs(5715) <= b;
    outputs(5716) <= a xor b;
    outputs(5717) <= a and not b;
    outputs(5718) <= not b;
    outputs(5719) <= not (a or b);
    outputs(5720) <= not b;
    outputs(5721) <= a xor b;
    outputs(5722) <= b;
    outputs(5723) <= b and not a;
    outputs(5724) <= b and not a;
    outputs(5725) <= a;
    outputs(5726) <= b;
    outputs(5727) <= a xor b;
    outputs(5728) <= a and b;
    outputs(5729) <= b;
    outputs(5730) <= a;
    outputs(5731) <= b and not a;
    outputs(5732) <= a;
    outputs(5733) <= not (a xor b);
    outputs(5734) <= a and b;
    outputs(5735) <= a xor b;
    outputs(5736) <= b and not a;
    outputs(5737) <= a xor b;
    outputs(5738) <= not (a or b);
    outputs(5739) <= not (a and b);
    outputs(5740) <= not a;
    outputs(5741) <= b and not a;
    outputs(5742) <= a and b;
    outputs(5743) <= not (a or b);
    outputs(5744) <= a xor b;
    outputs(5745) <= a and not b;
    outputs(5746) <= not a;
    outputs(5747) <= a and b;
    outputs(5748) <= a and b;
    outputs(5749) <= a and not b;
    outputs(5750) <= not a;
    outputs(5751) <= a xor b;
    outputs(5752) <= not a;
    outputs(5753) <= a and b;
    outputs(5754) <= a xor b;
    outputs(5755) <= not (a or b);
    outputs(5756) <= not b;
    outputs(5757) <= b;
    outputs(5758) <= not a;
    outputs(5759) <= not a;
    outputs(5760) <= a xor b;
    outputs(5761) <= not b;
    outputs(5762) <= b;
    outputs(5763) <= not (a xor b);
    outputs(5764) <= not b or a;
    outputs(5765) <= b;
    outputs(5766) <= not (a xor b);
    outputs(5767) <= a and b;
    outputs(5768) <= b;
    outputs(5769) <= a and not b;
    outputs(5770) <= b;
    outputs(5771) <= not a;
    outputs(5772) <= a and not b;
    outputs(5773) <= 1'b0;
    outputs(5774) <= not a or b;
    outputs(5775) <= a;
    outputs(5776) <= b;
    outputs(5777) <= b;
    outputs(5778) <= not (a xor b);
    outputs(5779) <= b and not a;
    outputs(5780) <= not (a xor b);
    outputs(5781) <= not b;
    outputs(5782) <= 1'b0;
    outputs(5783) <= not a;
    outputs(5784) <= a xor b;
    outputs(5785) <= not b;
    outputs(5786) <= not b or a;
    outputs(5787) <= a and not b;
    outputs(5788) <= a xor b;
    outputs(5789) <= b and not a;
    outputs(5790) <= not b;
    outputs(5791) <= not (a xor b);
    outputs(5792) <= a xor b;
    outputs(5793) <= a and not b;
    outputs(5794) <= a and not b;
    outputs(5795) <= not b;
    outputs(5796) <= a xor b;
    outputs(5797) <= not (a or b);
    outputs(5798) <= not (a xor b);
    outputs(5799) <= not a;
    outputs(5800) <= b;
    outputs(5801) <= not a;
    outputs(5802) <= not b or a;
    outputs(5803) <= not b;
    outputs(5804) <= a and b;
    outputs(5805) <= a xor b;
    outputs(5806) <= not (a xor b);
    outputs(5807) <= a;
    outputs(5808) <= not (a or b);
    outputs(5809) <= b and not a;
    outputs(5810) <= not a or b;
    outputs(5811) <= a;
    outputs(5812) <= a;
    outputs(5813) <= a xor b;
    outputs(5814) <= not b;
    outputs(5815) <= a xor b;
    outputs(5816) <= not (a or b);
    outputs(5817) <= a and b;
    outputs(5818) <= b and not a;
    outputs(5819) <= not a;
    outputs(5820) <= a and not b;
    outputs(5821) <= b and not a;
    outputs(5822) <= not (a xor b);
    outputs(5823) <= a;
    outputs(5824) <= a and b;
    outputs(5825) <= a and not b;
    outputs(5826) <= not b;
    outputs(5827) <= a;
    outputs(5828) <= not b;
    outputs(5829) <= not (a xor b);
    outputs(5830) <= not a;
    outputs(5831) <= a;
    outputs(5832) <= b;
    outputs(5833) <= not (a xor b);
    outputs(5834) <= b and not a;
    outputs(5835) <= a and not b;
    outputs(5836) <= not (a xor b);
    outputs(5837) <= a;
    outputs(5838) <= a and not b;
    outputs(5839) <= not b;
    outputs(5840) <= not a or b;
    outputs(5841) <= a xor b;
    outputs(5842) <= not (a or b);
    outputs(5843) <= a or b;
    outputs(5844) <= not a;
    outputs(5845) <= b;
    outputs(5846) <= not a;
    outputs(5847) <= a;
    outputs(5848) <= not b or a;
    outputs(5849) <= a;
    outputs(5850) <= b and not a;
    outputs(5851) <= a and not b;
    outputs(5852) <= a and not b;
    outputs(5853) <= not (a or b);
    outputs(5854) <= a xor b;
    outputs(5855) <= a and not b;
    outputs(5856) <= not a;
    outputs(5857) <= b;
    outputs(5858) <= a or b;
    outputs(5859) <= a and not b;
    outputs(5860) <= a and not b;
    outputs(5861) <= not a;
    outputs(5862) <= a and b;
    outputs(5863) <= a and not b;
    outputs(5864) <= not b;
    outputs(5865) <= not (a xor b);
    outputs(5866) <= a and b;
    outputs(5867) <= a and not b;
    outputs(5868) <= not b;
    outputs(5869) <= not a or b;
    outputs(5870) <= b and not a;
    outputs(5871) <= not (a or b);
    outputs(5872) <= not b;
    outputs(5873) <= b;
    outputs(5874) <= not (a or b);
    outputs(5875) <= a and b;
    outputs(5876) <= a xor b;
    outputs(5877) <= a xor b;
    outputs(5878) <= a or b;
    outputs(5879) <= a xor b;
    outputs(5880) <= not (a or b);
    outputs(5881) <= not a or b;
    outputs(5882) <= not (a xor b);
    outputs(5883) <= 1'b0;
    outputs(5884) <= b and not a;
    outputs(5885) <= not b;
    outputs(5886) <= b and not a;
    outputs(5887) <= a;
    outputs(5888) <= b and not a;
    outputs(5889) <= not (a xor b);
    outputs(5890) <= not b;
    outputs(5891) <= b and not a;
    outputs(5892) <= not a;
    outputs(5893) <= not b;
    outputs(5894) <= not (a xor b);
    outputs(5895) <= not a;
    outputs(5896) <= a xor b;
    outputs(5897) <= a;
    outputs(5898) <= not b;
    outputs(5899) <= not (a or b);
    outputs(5900) <= b;
    outputs(5901) <= not (a xor b);
    outputs(5902) <= not b;
    outputs(5903) <= not (a xor b);
    outputs(5904) <= not a;
    outputs(5905) <= not b;
    outputs(5906) <= a and b;
    outputs(5907) <= not (a xor b);
    outputs(5908) <= a;
    outputs(5909) <= not (a xor b);
    outputs(5910) <= not a;
    outputs(5911) <= b and not a;
    outputs(5912) <= b;
    outputs(5913) <= a and b;
    outputs(5914) <= a;
    outputs(5915) <= not (a or b);
    outputs(5916) <= a;
    outputs(5917) <= a and b;
    outputs(5918) <= not (a or b);
    outputs(5919) <= a xor b;
    outputs(5920) <= a and not b;
    outputs(5921) <= not a;
    outputs(5922) <= a xor b;
    outputs(5923) <= not (a or b);
    outputs(5924) <= not (a xor b);
    outputs(5925) <= a xor b;
    outputs(5926) <= a and b;
    outputs(5927) <= a and not b;
    outputs(5928) <= not (a xor b);
    outputs(5929) <= not (a xor b);
    outputs(5930) <= not b;
    outputs(5931) <= a xor b;
    outputs(5932) <= b;
    outputs(5933) <= not a;
    outputs(5934) <= a and b;
    outputs(5935) <= not (a or b);
    outputs(5936) <= not (a or b);
    outputs(5937) <= a xor b;
    outputs(5938) <= not a;
    outputs(5939) <= not (a xor b);
    outputs(5940) <= not a;
    outputs(5941) <= not b;
    outputs(5942) <= b and not a;
    outputs(5943) <= a and not b;
    outputs(5944) <= a xor b;
    outputs(5945) <= not a;
    outputs(5946) <= a xor b;
    outputs(5947) <= a and b;
    outputs(5948) <= not a;
    outputs(5949) <= not b or a;
    outputs(5950) <= not (a xor b);
    outputs(5951) <= a and not b;
    outputs(5952) <= a xor b;
    outputs(5953) <= a and not b;
    outputs(5954) <= not (a xor b);
    outputs(5955) <= not (a or b);
    outputs(5956) <= a and b;
    outputs(5957) <= not (a xor b);
    outputs(5958) <= b and not a;
    outputs(5959) <= not b;
    outputs(5960) <= a xor b;
    outputs(5961) <= not (a xor b);
    outputs(5962) <= a xor b;
    outputs(5963) <= not b;
    outputs(5964) <= a;
    outputs(5965) <= not b;
    outputs(5966) <= b and not a;
    outputs(5967) <= not (a xor b);
    outputs(5968) <= b;
    outputs(5969) <= not b or a;
    outputs(5970) <= a and not b;
    outputs(5971) <= a and not b;
    outputs(5972) <= not b;
    outputs(5973) <= a and not b;
    outputs(5974) <= a xor b;
    outputs(5975) <= not b;
    outputs(5976) <= b and not a;
    outputs(5977) <= not (a and b);
    outputs(5978) <= not (a xor b);
    outputs(5979) <= a xor b;
    outputs(5980) <= not (a or b);
    outputs(5981) <= a xor b;
    outputs(5982) <= b;
    outputs(5983) <= b;
    outputs(5984) <= not (a or b);
    outputs(5985) <= not (a xor b);
    outputs(5986) <= not (a xor b);
    outputs(5987) <= a and b;
    outputs(5988) <= a or b;
    outputs(5989) <= a and not b;
    outputs(5990) <= a and b;
    outputs(5991) <= not (a or b);
    outputs(5992) <= not (a or b);
    outputs(5993) <= a;
    outputs(5994) <= a and not b;
    outputs(5995) <= not a;
    outputs(5996) <= a and not b;
    outputs(5997) <= a xor b;
    outputs(5998) <= a and b;
    outputs(5999) <= not b;
    outputs(6000) <= a and b;
    outputs(6001) <= b and not a;
    outputs(6002) <= b and not a;
    outputs(6003) <= not b;
    outputs(6004) <= a;
    outputs(6005) <= a;
    outputs(6006) <= not (a xor b);
    outputs(6007) <= not (a or b);
    outputs(6008) <= a and b;
    outputs(6009) <= not a;
    outputs(6010) <= a;
    outputs(6011) <= b;
    outputs(6012) <= b;
    outputs(6013) <= not (a xor b);
    outputs(6014) <= not (a or b);
    outputs(6015) <= not (a xor b);
    outputs(6016) <= a;
    outputs(6017) <= a;
    outputs(6018) <= not b;
    outputs(6019) <= not b;
    outputs(6020) <= b;
    outputs(6021) <= a;
    outputs(6022) <= b and not a;
    outputs(6023) <= not a;
    outputs(6024) <= a and b;
    outputs(6025) <= a;
    outputs(6026) <= a;
    outputs(6027) <= not b;
    outputs(6028) <= b and not a;
    outputs(6029) <= not a;
    outputs(6030) <= a xor b;
    outputs(6031) <= not b;
    outputs(6032) <= a or b;
    outputs(6033) <= a and b;
    outputs(6034) <= not (a xor b);
    outputs(6035) <= a and b;
    outputs(6036) <= a or b;
    outputs(6037) <= not (a or b);
    outputs(6038) <= b;
    outputs(6039) <= b and not a;
    outputs(6040) <= not (a xor b);
    outputs(6041) <= a;
    outputs(6042) <= b and not a;
    outputs(6043) <= a and b;
    outputs(6044) <= b;
    outputs(6045) <= a and not b;
    outputs(6046) <= b;
    outputs(6047) <= b and not a;
    outputs(6048) <= a or b;
    outputs(6049) <= not b;
    outputs(6050) <= a;
    outputs(6051) <= a;
    outputs(6052) <= not b;
    outputs(6053) <= a xor b;
    outputs(6054) <= a;
    outputs(6055) <= not b;
    outputs(6056) <= not a;
    outputs(6057) <= a and b;
    outputs(6058) <= not (a or b);
    outputs(6059) <= not a;
    outputs(6060) <= not a or b;
    outputs(6061) <= a or b;
    outputs(6062) <= a;
    outputs(6063) <= a and not b;
    outputs(6064) <= b;
    outputs(6065) <= not b;
    outputs(6066) <= a and not b;
    outputs(6067) <= a xor b;
    outputs(6068) <= not a or b;
    outputs(6069) <= not (a xor b);
    outputs(6070) <= not a;
    outputs(6071) <= a xor b;
    outputs(6072) <= a;
    outputs(6073) <= not b or a;
    outputs(6074) <= not a;
    outputs(6075) <= not (a xor b);
    outputs(6076) <= not (a or b);
    outputs(6077) <= not b or a;
    outputs(6078) <= a;
    outputs(6079) <= not (a xor b);
    outputs(6080) <= a and not b;
    outputs(6081) <= a xor b;
    outputs(6082) <= a xor b;
    outputs(6083) <= not b or a;
    outputs(6084) <= a and b;
    outputs(6085) <= b and not a;
    outputs(6086) <= a or b;
    outputs(6087) <= not (a or b);
    outputs(6088) <= not (a xor b);
    outputs(6089) <= a and b;
    outputs(6090) <= b and not a;
    outputs(6091) <= a xor b;
    outputs(6092) <= not (a xor b);
    outputs(6093) <= not a;
    outputs(6094) <= b and not a;
    outputs(6095) <= not (a xor b);
    outputs(6096) <= b and not a;
    outputs(6097) <= not a;
    outputs(6098) <= a and b;
    outputs(6099) <= 1'b0;
    outputs(6100) <= not b;
    outputs(6101) <= not a;
    outputs(6102) <= not (a or b);
    outputs(6103) <= a xor b;
    outputs(6104) <= b;
    outputs(6105) <= a and b;
    outputs(6106) <= a;
    outputs(6107) <= not a;
    outputs(6108) <= b and not a;
    outputs(6109) <= a xor b;
    outputs(6110) <= a and b;
    outputs(6111) <= not (a and b);
    outputs(6112) <= a and b;
    outputs(6113) <= a and not b;
    outputs(6114) <= not (a or b);
    outputs(6115) <= not (a xor b);
    outputs(6116) <= not a;
    outputs(6117) <= a;
    outputs(6118) <= not b;
    outputs(6119) <= not b;
    outputs(6120) <= a and not b;
    outputs(6121) <= not a;
    outputs(6122) <= not (a xor b);
    outputs(6123) <= a and b;
    outputs(6124) <= a and b;
    outputs(6125) <= not (a xor b);
    outputs(6126) <= not (a or b);
    outputs(6127) <= a and b;
    outputs(6128) <= not (a xor b);
    outputs(6129) <= a and b;
    outputs(6130) <= not a;
    outputs(6131) <= not (a xor b);
    outputs(6132) <= not a;
    outputs(6133) <= a;
    outputs(6134) <= not (a xor b);
    outputs(6135) <= a or b;
    outputs(6136) <= not a;
    outputs(6137) <= b;
    outputs(6138) <= b;
    outputs(6139) <= a and not b;
    outputs(6140) <= a xor b;
    outputs(6141) <= not (a xor b);
    outputs(6142) <= not (a xor b);
    outputs(6143) <= not (a xor b);
    outputs(6144) <= not (a xor b);
    outputs(6145) <= a and not b;
    outputs(6146) <= a and b;
    outputs(6147) <= a xor b;
    outputs(6148) <= a and b;
    outputs(6149) <= not (a or b);
    outputs(6150) <= b;
    outputs(6151) <= a;
    outputs(6152) <= a and not b;
    outputs(6153) <= not (a or b);
    outputs(6154) <= a and b;
    outputs(6155) <= a;
    outputs(6156) <= a and b;
    outputs(6157) <= a;
    outputs(6158) <= a and not b;
    outputs(6159) <= b and not a;
    outputs(6160) <= not b;
    outputs(6161) <= a;
    outputs(6162) <= not a;
    outputs(6163) <= not (a xor b);
    outputs(6164) <= not (a xor b);
    outputs(6165) <= not a or b;
    outputs(6166) <= not a;
    outputs(6167) <= a and b;
    outputs(6168) <= not (a xor b);
    outputs(6169) <= not a;
    outputs(6170) <= a and not b;
    outputs(6171) <= a;
    outputs(6172) <= not (a or b);
    outputs(6173) <= b and not a;
    outputs(6174) <= not b or a;
    outputs(6175) <= not (a xor b);
    outputs(6176) <= a;
    outputs(6177) <= not a;
    outputs(6178) <= not (a xor b);
    outputs(6179) <= a;
    outputs(6180) <= b;
    outputs(6181) <= a xor b;
    outputs(6182) <= not b or a;
    outputs(6183) <= not (a xor b);
    outputs(6184) <= a and not b;
    outputs(6185) <= a and not b;
    outputs(6186) <= a xor b;
    outputs(6187) <= a and not b;
    outputs(6188) <= b;
    outputs(6189) <= b and not a;
    outputs(6190) <= a;
    outputs(6191) <= b;
    outputs(6192) <= a and not b;
    outputs(6193) <= a xor b;
    outputs(6194) <= a xor b;
    outputs(6195) <= not (a or b);
    outputs(6196) <= a xor b;
    outputs(6197) <= a and not b;
    outputs(6198) <= a xor b;
    outputs(6199) <= a and b;
    outputs(6200) <= a and not b;
    outputs(6201) <= not b;
    outputs(6202) <= a and not b;
    outputs(6203) <= a and not b;
    outputs(6204) <= not (a or b);
    outputs(6205) <= not b;
    outputs(6206) <= a and b;
    outputs(6207) <= a and b;
    outputs(6208) <= a xor b;
    outputs(6209) <= a and not b;
    outputs(6210) <= a xor b;
    outputs(6211) <= b;
    outputs(6212) <= a and b;
    outputs(6213) <= b;
    outputs(6214) <= b;
    outputs(6215) <= a and b;
    outputs(6216) <= not (a xor b);
    outputs(6217) <= not a;
    outputs(6218) <= a xor b;
    outputs(6219) <= not a or b;
    outputs(6220) <= a and b;
    outputs(6221) <= a xor b;
    outputs(6222) <= b;
    outputs(6223) <= a and b;
    outputs(6224) <= not a;
    outputs(6225) <= a xor b;
    outputs(6226) <= not b;
    outputs(6227) <= not (a xor b);
    outputs(6228) <= b;
    outputs(6229) <= not a;
    outputs(6230) <= a;
    outputs(6231) <= not (a xor b);
    outputs(6232) <= not (a and b);
    outputs(6233) <= not (a xor b);
    outputs(6234) <= b;
    outputs(6235) <= not a;
    outputs(6236) <= a xor b;
    outputs(6237) <= a;
    outputs(6238) <= not (a or b);
    outputs(6239) <= a;
    outputs(6240) <= a and b;
    outputs(6241) <= b and not a;
    outputs(6242) <= a xor b;
    outputs(6243) <= b;
    outputs(6244) <= not b;
    outputs(6245) <= not b;
    outputs(6246) <= b;
    outputs(6247) <= not a;
    outputs(6248) <= a;
    outputs(6249) <= a and not b;
    outputs(6250) <= a and b;
    outputs(6251) <= b and not a;
    outputs(6252) <= not (a xor b);
    outputs(6253) <= a and b;
    outputs(6254) <= a and not b;
    outputs(6255) <= not a or b;
    outputs(6256) <= b and not a;
    outputs(6257) <= not (a or b);
    outputs(6258) <= not (a or b);
    outputs(6259) <= a and not b;
    outputs(6260) <= b and not a;
    outputs(6261) <= not (a xor b);
    outputs(6262) <= b;
    outputs(6263) <= not b or a;
    outputs(6264) <= a;
    outputs(6265) <= a and b;
    outputs(6266) <= a;
    outputs(6267) <= not (a xor b);
    outputs(6268) <= not (a xor b);
    outputs(6269) <= a xor b;
    outputs(6270) <= not (a or b);
    outputs(6271) <= b and not a;
    outputs(6272) <= a and b;
    outputs(6273) <= a;
    outputs(6274) <= b;
    outputs(6275) <= not (a xor b);
    outputs(6276) <= a;
    outputs(6277) <= not b or a;
    outputs(6278) <= a and not b;
    outputs(6279) <= b;
    outputs(6280) <= a and not b;
    outputs(6281) <= b and not a;
    outputs(6282) <= a xor b;
    outputs(6283) <= b and not a;
    outputs(6284) <= b;
    outputs(6285) <= not b;
    outputs(6286) <= not (a xor b);
    outputs(6287) <= a;
    outputs(6288) <= not (a xor b);
    outputs(6289) <= not a or b;
    outputs(6290) <= not (a xor b);
    outputs(6291) <= b;
    outputs(6292) <= not (a xor b);
    outputs(6293) <= a and not b;
    outputs(6294) <= not (a or b);
    outputs(6295) <= b;
    outputs(6296) <= a and not b;
    outputs(6297) <= a and b;
    outputs(6298) <= b and not a;
    outputs(6299) <= b;
    outputs(6300) <= not a;
    outputs(6301) <= not (a xor b);
    outputs(6302) <= b and not a;
    outputs(6303) <= not a or b;
    outputs(6304) <= not b;
    outputs(6305) <= a;
    outputs(6306) <= b and not a;
    outputs(6307) <= a xor b;
    outputs(6308) <= a and b;
    outputs(6309) <= not b;
    outputs(6310) <= not b;
    outputs(6311) <= a and b;
    outputs(6312) <= not (a or b);
    outputs(6313) <= a and not b;
    outputs(6314) <= not (a xor b);
    outputs(6315) <= b;
    outputs(6316) <= not (a xor b);
    outputs(6317) <= not (a or b);
    outputs(6318) <= not (a xor b);
    outputs(6319) <= a xor b;
    outputs(6320) <= b;
    outputs(6321) <= b and not a;
    outputs(6322) <= a and not b;
    outputs(6323) <= not b;
    outputs(6324) <= a and not b;
    outputs(6325) <= b and not a;
    outputs(6326) <= b;
    outputs(6327) <= a and b;
    outputs(6328) <= not b;
    outputs(6329) <= a;
    outputs(6330) <= a and not b;
    outputs(6331) <= not (a xor b);
    outputs(6332) <= b and not a;
    outputs(6333) <= a and not b;
    outputs(6334) <= b;
    outputs(6335) <= b;
    outputs(6336) <= not (a or b);
    outputs(6337) <= not a;
    outputs(6338) <= not (a or b);
    outputs(6339) <= b;
    outputs(6340) <= not a or b;
    outputs(6341) <= not a;
    outputs(6342) <= not (a or b);
    outputs(6343) <= b and not a;
    outputs(6344) <= b and not a;
    outputs(6345) <= a xor b;
    outputs(6346) <= not b;
    outputs(6347) <= not (a or b);
    outputs(6348) <= b and not a;
    outputs(6349) <= not (a xor b);
    outputs(6350) <= a and not b;
    outputs(6351) <= not (a xor b);
    outputs(6352) <= a xor b;
    outputs(6353) <= a and b;
    outputs(6354) <= a xor b;
    outputs(6355) <= not a;
    outputs(6356) <= a and not b;
    outputs(6357) <= not b;
    outputs(6358) <= b and not a;
    outputs(6359) <= b;
    outputs(6360) <= a and not b;
    outputs(6361) <= b;
    outputs(6362) <= not a;
    outputs(6363) <= a;
    outputs(6364) <= a;
    outputs(6365) <= not (a xor b);
    outputs(6366) <= a and b;
    outputs(6367) <= not (a or b);
    outputs(6368) <= not b or a;
    outputs(6369) <= a and not b;
    outputs(6370) <= not a;
    outputs(6371) <= b;
    outputs(6372) <= not (a or b);
    outputs(6373) <= not a;
    outputs(6374) <= b and not a;
    outputs(6375) <= b and not a;
    outputs(6376) <= a xor b;
    outputs(6377) <= not b;
    outputs(6378) <= a xor b;
    outputs(6379) <= not b;
    outputs(6380) <= a and not b;
    outputs(6381) <= a;
    outputs(6382) <= not (a xor b);
    outputs(6383) <= a and b;
    outputs(6384) <= b and not a;
    outputs(6385) <= not (a xor b);
    outputs(6386) <= not a or b;
    outputs(6387) <= not (a xor b);
    outputs(6388) <= not (a xor b);
    outputs(6389) <= not a;
    outputs(6390) <= b;
    outputs(6391) <= not a;
    outputs(6392) <= a and not b;
    outputs(6393) <= a and not b;
    outputs(6394) <= not (a xor b);
    outputs(6395) <= not (a xor b);
    outputs(6396) <= not a;
    outputs(6397) <= b;
    outputs(6398) <= not b;
    outputs(6399) <= a and b;
    outputs(6400) <= a and not b;
    outputs(6401) <= not (a xor b);
    outputs(6402) <= b;
    outputs(6403) <= a;
    outputs(6404) <= a;
    outputs(6405) <= not (a xor b);
    outputs(6406) <= not a or b;
    outputs(6407) <= b and not a;
    outputs(6408) <= not a or b;
    outputs(6409) <= b;
    outputs(6410) <= a xor b;
    outputs(6411) <= a xor b;
    outputs(6412) <= a xor b;
    outputs(6413) <= not b;
    outputs(6414) <= not a or b;
    outputs(6415) <= b;
    outputs(6416) <= not (a and b);
    outputs(6417) <= not a or b;
    outputs(6418) <= a xor b;
    outputs(6419) <= not b;
    outputs(6420) <= b;
    outputs(6421) <= a xor b;
    outputs(6422) <= not a;
    outputs(6423) <= not (a xor b);
    outputs(6424) <= a and b;
    outputs(6425) <= a xor b;
    outputs(6426) <= a xor b;
    outputs(6427) <= a xor b;
    outputs(6428) <= a xor b;
    outputs(6429) <= not b;
    outputs(6430) <= b and not a;
    outputs(6431) <= not (a and b);
    outputs(6432) <= not (a or b);
    outputs(6433) <= not (a xor b);
    outputs(6434) <= not b or a;
    outputs(6435) <= a xor b;
    outputs(6436) <= not (a xor b);
    outputs(6437) <= a xor b;
    outputs(6438) <= not a or b;
    outputs(6439) <= a xor b;
    outputs(6440) <= a and not b;
    outputs(6441) <= not (a xor b);
    outputs(6442) <= a xor b;
    outputs(6443) <= b and not a;
    outputs(6444) <= not (a xor b);
    outputs(6445) <= a xor b;
    outputs(6446) <= not b;
    outputs(6447) <= a;
    outputs(6448) <= not (a xor b);
    outputs(6449) <= not b;
    outputs(6450) <= a or b;
    outputs(6451) <= a xor b;
    outputs(6452) <= b and not a;
    outputs(6453) <= a xor b;
    outputs(6454) <= not (a or b);
    outputs(6455) <= not b;
    outputs(6456) <= a or b;
    outputs(6457) <= not a or b;
    outputs(6458) <= a;
    outputs(6459) <= b and not a;
    outputs(6460) <= a and b;
    outputs(6461) <= a xor b;
    outputs(6462) <= a xor b;
    outputs(6463) <= not a;
    outputs(6464) <= not a or b;
    outputs(6465) <= a;
    outputs(6466) <= not (a xor b);
    outputs(6467) <= a;
    outputs(6468) <= a;
    outputs(6469) <= not (a or b);
    outputs(6470) <= a xor b;
    outputs(6471) <= b;
    outputs(6472) <= not b;
    outputs(6473) <= b;
    outputs(6474) <= a xor b;
    outputs(6475) <= a xor b;
    outputs(6476) <= not a;
    outputs(6477) <= not b or a;
    outputs(6478) <= a or b;
    outputs(6479) <= a and b;
    outputs(6480) <= b;
    outputs(6481) <= a xor b;
    outputs(6482) <= not b;
    outputs(6483) <= a xor b;
    outputs(6484) <= a and b;
    outputs(6485) <= not b;
    outputs(6486) <= not (a and b);
    outputs(6487) <= b and not a;
    outputs(6488) <= b;
    outputs(6489) <= a and not b;
    outputs(6490) <= not (a and b);
    outputs(6491) <= not (a xor b);
    outputs(6492) <= a or b;
    outputs(6493) <= a and not b;
    outputs(6494) <= not (a xor b);
    outputs(6495) <= a;
    outputs(6496) <= not a or b;
    outputs(6497) <= not (a xor b);
    outputs(6498) <= not (a xor b);
    outputs(6499) <= not b or a;
    outputs(6500) <= b;
    outputs(6501) <= not (a xor b);
    outputs(6502) <= not (a xor b);
    outputs(6503) <= b and not a;
    outputs(6504) <= b and not a;
    outputs(6505) <= a or b;
    outputs(6506) <= a;
    outputs(6507) <= a;
    outputs(6508) <= a xor b;
    outputs(6509) <= a xor b;
    outputs(6510) <= b;
    outputs(6511) <= a;
    outputs(6512) <= a;
    outputs(6513) <= not a or b;
    outputs(6514) <= not a or b;
    outputs(6515) <= a xor b;
    outputs(6516) <= a xor b;
    outputs(6517) <= a xor b;
    outputs(6518) <= not (a xor b);
    outputs(6519) <= b;
    outputs(6520) <= a xor b;
    outputs(6521) <= not (a and b);
    outputs(6522) <= not a;
    outputs(6523) <= a xor b;
    outputs(6524) <= not a or b;
    outputs(6525) <= a xor b;
    outputs(6526) <= not (a xor b);
    outputs(6527) <= b;
    outputs(6528) <= not b;
    outputs(6529) <= b;
    outputs(6530) <= not a or b;
    outputs(6531) <= a xor b;
    outputs(6532) <= not (a or b);
    outputs(6533) <= a;
    outputs(6534) <= a and not b;
    outputs(6535) <= a;
    outputs(6536) <= not (a xor b);
    outputs(6537) <= b;
    outputs(6538) <= a xor b;
    outputs(6539) <= a xor b;
    outputs(6540) <= a and b;
    outputs(6541) <= a and b;
    outputs(6542) <= a xor b;
    outputs(6543) <= 1'b1;
    outputs(6544) <= not a or b;
    outputs(6545) <= not b or a;
    outputs(6546) <= b and not a;
    outputs(6547) <= not b;
    outputs(6548) <= a;
    outputs(6549) <= a;
    outputs(6550) <= not (a xor b);
    outputs(6551) <= b;
    outputs(6552) <= not (a xor b);
    outputs(6553) <= b;
    outputs(6554) <= not (a xor b);
    outputs(6555) <= a xor b;
    outputs(6556) <= a xor b;
    outputs(6557) <= b;
    outputs(6558) <= b;
    outputs(6559) <= not (a and b);
    outputs(6560) <= a xor b;
    outputs(6561) <= not b or a;
    outputs(6562) <= a xor b;
    outputs(6563) <= b and not a;
    outputs(6564) <= not (a xor b);
    outputs(6565) <= not a;
    outputs(6566) <= not (a xor b);
    outputs(6567) <= b;
    outputs(6568) <= b;
    outputs(6569) <= not (a and b);
    outputs(6570) <= not a or b;
    outputs(6571) <= not b;
    outputs(6572) <= not a or b;
    outputs(6573) <= not (a xor b);
    outputs(6574) <= not a;
    outputs(6575) <= b and not a;
    outputs(6576) <= not b;
    outputs(6577) <= not (a xor b);
    outputs(6578) <= not (a xor b);
    outputs(6579) <= b and not a;
    outputs(6580) <= not a or b;
    outputs(6581) <= a or b;
    outputs(6582) <= not (a xor b);
    outputs(6583) <= b and not a;
    outputs(6584) <= not b;
    outputs(6585) <= not (a or b);
    outputs(6586) <= not a;
    outputs(6587) <= not a or b;
    outputs(6588) <= b;
    outputs(6589) <= not a or b;
    outputs(6590) <= not (a and b);
    outputs(6591) <= a and b;
    outputs(6592) <= a;
    outputs(6593) <= a;
    outputs(6594) <= not (a xor b);
    outputs(6595) <= not (a xor b);
    outputs(6596) <= a and b;
    outputs(6597) <= a;
    outputs(6598) <= not (a and b);
    outputs(6599) <= a xor b;
    outputs(6600) <= not (a and b);
    outputs(6601) <= not a;
    outputs(6602) <= b and not a;
    outputs(6603) <= a xor b;
    outputs(6604) <= not (a xor b);
    outputs(6605) <= not (a xor b);
    outputs(6606) <= not (a xor b);
    outputs(6607) <= not (a xor b);
    outputs(6608) <= a and not b;
    outputs(6609) <= a xor b;
    outputs(6610) <= not (a xor b);
    outputs(6611) <= a xor b;
    outputs(6612) <= not (a xor b);
    outputs(6613) <= not a;
    outputs(6614) <= a or b;
    outputs(6615) <= not (a or b);
    outputs(6616) <= b;
    outputs(6617) <= b;
    outputs(6618) <= not b;
    outputs(6619) <= not (a xor b);
    outputs(6620) <= not (a and b);
    outputs(6621) <= not (a xor b);
    outputs(6622) <= a xor b;
    outputs(6623) <= not b;
    outputs(6624) <= not b;
    outputs(6625) <= not a;
    outputs(6626) <= a;
    outputs(6627) <= a xor b;
    outputs(6628) <= a xor b;
    outputs(6629) <= not b or a;
    outputs(6630) <= a;
    outputs(6631) <= not (a xor b);
    outputs(6632) <= a xor b;
    outputs(6633) <= b and not a;
    outputs(6634) <= not a;
    outputs(6635) <= not a;
    outputs(6636) <= not (a xor b);
    outputs(6637) <= a and b;
    outputs(6638) <= not a or b;
    outputs(6639) <= b;
    outputs(6640) <= not (a and b);
    outputs(6641) <= a and b;
    outputs(6642) <= not (a or b);
    outputs(6643) <= a or b;
    outputs(6644) <= a;
    outputs(6645) <= a xor b;
    outputs(6646) <= b;
    outputs(6647) <= not b or a;
    outputs(6648) <= not a;
    outputs(6649) <= not (a xor b);
    outputs(6650) <= a or b;
    outputs(6651) <= not (a xor b);
    outputs(6652) <= not a;
    outputs(6653) <= not (a xor b);
    outputs(6654) <= not (a xor b);
    outputs(6655) <= not a;
    outputs(6656) <= a or b;
    outputs(6657) <= not a;
    outputs(6658) <= a;
    outputs(6659) <= a xor b;
    outputs(6660) <= not (a xor b);
    outputs(6661) <= a xor b;
    outputs(6662) <= b;
    outputs(6663) <= not b or a;
    outputs(6664) <= not (a xor b);
    outputs(6665) <= b;
    outputs(6666) <= a xor b;
    outputs(6667) <= a or b;
    outputs(6668) <= a xor b;
    outputs(6669) <= b;
    outputs(6670) <= a;
    outputs(6671) <= a xor b;
    outputs(6672) <= a xor b;
    outputs(6673) <= a xor b;
    outputs(6674) <= not b or a;
    outputs(6675) <= a;
    outputs(6676) <= not (a xor b);
    outputs(6677) <= not (a xor b);
    outputs(6678) <= a xor b;
    outputs(6679) <= not (a xor b);
    outputs(6680) <= not (a and b);
    outputs(6681) <= a and b;
    outputs(6682) <= not (a or b);
    outputs(6683) <= a;
    outputs(6684) <= a or b;
    outputs(6685) <= b;
    outputs(6686) <= b and not a;
    outputs(6687) <= a xor b;
    outputs(6688) <= b and not a;
    outputs(6689) <= a xor b;
    outputs(6690) <= a xor b;
    outputs(6691) <= not b;
    outputs(6692) <= not b;
    outputs(6693) <= not (a or b);
    outputs(6694) <= not (a xor b);
    outputs(6695) <= not (a xor b);
    outputs(6696) <= not (a and b);
    outputs(6697) <= b;
    outputs(6698) <= a and b;
    outputs(6699) <= a xor b;
    outputs(6700) <= not (a and b);
    outputs(6701) <= not b;
    outputs(6702) <= a or b;
    outputs(6703) <= b and not a;
    outputs(6704) <= a;
    outputs(6705) <= a;
    outputs(6706) <= b and not a;
    outputs(6707) <= b;
    outputs(6708) <= not a;
    outputs(6709) <= a and b;
    outputs(6710) <= not (a and b);
    outputs(6711) <= a xor b;
    outputs(6712) <= a;
    outputs(6713) <= a xor b;
    outputs(6714) <= not a or b;
    outputs(6715) <= not (a and b);
    outputs(6716) <= not (a xor b);
    outputs(6717) <= not a;
    outputs(6718) <= not b or a;
    outputs(6719) <= b;
    outputs(6720) <= not b or a;
    outputs(6721) <= not (a or b);
    outputs(6722) <= not (a and b);
    outputs(6723) <= a xor b;
    outputs(6724) <= a xor b;
    outputs(6725) <= a or b;
    outputs(6726) <= not a or b;
    outputs(6727) <= not b or a;
    outputs(6728) <= b;
    outputs(6729) <= not (a xor b);
    outputs(6730) <= a xor b;
    outputs(6731) <= a and not b;
    outputs(6732) <= a xor b;
    outputs(6733) <= not a or b;
    outputs(6734) <= b;
    outputs(6735) <= a and not b;
    outputs(6736) <= not a;
    outputs(6737) <= not (a and b);
    outputs(6738) <= b and not a;
    outputs(6739) <= b;
    outputs(6740) <= b;
    outputs(6741) <= not a or b;
    outputs(6742) <= not b;
    outputs(6743) <= not b or a;
    outputs(6744) <= a;
    outputs(6745) <= not b;
    outputs(6746) <= not (a xor b);
    outputs(6747) <= not (a xor b);
    outputs(6748) <= not b;
    outputs(6749) <= not b;
    outputs(6750) <= not (a xor b);
    outputs(6751) <= not (a xor b);
    outputs(6752) <= not (a xor b);
    outputs(6753) <= not b or a;
    outputs(6754) <= a and b;
    outputs(6755) <= not a or b;
    outputs(6756) <= not (a xor b);
    outputs(6757) <= a or b;
    outputs(6758) <= not (a and b);
    outputs(6759) <= not a;
    outputs(6760) <= a and not b;
    outputs(6761) <= a xor b;
    outputs(6762) <= a and b;
    outputs(6763) <= not a;
    outputs(6764) <= not b;
    outputs(6765) <= a;
    outputs(6766) <= a xor b;
    outputs(6767) <= not a;
    outputs(6768) <= a;
    outputs(6769) <= a xor b;
    outputs(6770) <= not b;
    outputs(6771) <= a and b;
    outputs(6772) <= a xor b;
    outputs(6773) <= a;
    outputs(6774) <= a xor b;
    outputs(6775) <= a xor b;
    outputs(6776) <= not b;
    outputs(6777) <= a xor b;
    outputs(6778) <= b and not a;
    outputs(6779) <= not a;
    outputs(6780) <= b;
    outputs(6781) <= a xor b;
    outputs(6782) <= a xor b;
    outputs(6783) <= not a;
    outputs(6784) <= a;
    outputs(6785) <= not b;
    outputs(6786) <= a xor b;
    outputs(6787) <= a xor b;
    outputs(6788) <= not (a xor b);
    outputs(6789) <= not (a or b);
    outputs(6790) <= not (a xor b);
    outputs(6791) <= b;
    outputs(6792) <= not a;
    outputs(6793) <= a xor b;
    outputs(6794) <= not b;
    outputs(6795) <= not a;
    outputs(6796) <= not (a and b);
    outputs(6797) <= not (a xor b);
    outputs(6798) <= a;
    outputs(6799) <= a xor b;
    outputs(6800) <= not (a xor b);
    outputs(6801) <= not (a xor b);
    outputs(6802) <= not a;
    outputs(6803) <= not b;
    outputs(6804) <= b;
    outputs(6805) <= a and b;
    outputs(6806) <= a and b;
    outputs(6807) <= not a;
    outputs(6808) <= not b;
    outputs(6809) <= b;
    outputs(6810) <= a and b;
    outputs(6811) <= b;
    outputs(6812) <= not b;
    outputs(6813) <= b;
    outputs(6814) <= a xor b;
    outputs(6815) <= b;
    outputs(6816) <= not (a xor b);
    outputs(6817) <= b and not a;
    outputs(6818) <= b and not a;
    outputs(6819) <= not b or a;
    outputs(6820) <= not (a xor b);
    outputs(6821) <= not (a xor b);
    outputs(6822) <= not (a and b);
    outputs(6823) <= a xor b;
    outputs(6824) <= not b or a;
    outputs(6825) <= not (a and b);
    outputs(6826) <= a and b;
    outputs(6827) <= b and not a;
    outputs(6828) <= not b;
    outputs(6829) <= a or b;
    outputs(6830) <= not (a xor b);
    outputs(6831) <= not (a xor b);
    outputs(6832) <= a and b;
    outputs(6833) <= not (a xor b);
    outputs(6834) <= a or b;
    outputs(6835) <= not (a xor b);
    outputs(6836) <= a xor b;
    outputs(6837) <= a xor b;
    outputs(6838) <= not (a and b);
    outputs(6839) <= not b or a;
    outputs(6840) <= not a or b;
    outputs(6841) <= not b or a;
    outputs(6842) <= not a;
    outputs(6843) <= a and b;
    outputs(6844) <= a and b;
    outputs(6845) <= a xor b;
    outputs(6846) <= a;
    outputs(6847) <= b;
    outputs(6848) <= a and b;
    outputs(6849) <= a or b;
    outputs(6850) <= a;
    outputs(6851) <= not (a xor b);
    outputs(6852) <= a and b;
    outputs(6853) <= not b;
    outputs(6854) <= not a;
    outputs(6855) <= a;
    outputs(6856) <= a;
    outputs(6857) <= a and not b;
    outputs(6858) <= not a;
    outputs(6859) <= a xor b;
    outputs(6860) <= not (a and b);
    outputs(6861) <= a xor b;
    outputs(6862) <= not b or a;
    outputs(6863) <= not (a xor b);
    outputs(6864) <= a and not b;
    outputs(6865) <= not b;
    outputs(6866) <= a or b;
    outputs(6867) <= a xor b;
    outputs(6868) <= not b;
    outputs(6869) <= a and b;
    outputs(6870) <= b and not a;
    outputs(6871) <= not (a xor b);
    outputs(6872) <= not (a or b);
    outputs(6873) <= not a;
    outputs(6874) <= not (a xor b);
    outputs(6875) <= not a;
    outputs(6876) <= not (a and b);
    outputs(6877) <= not b;
    outputs(6878) <= not (a xor b);
    outputs(6879) <= not (a xor b);
    outputs(6880) <= not a;
    outputs(6881) <= not b or a;
    outputs(6882) <= a and not b;
    outputs(6883) <= not (a xor b);
    outputs(6884) <= not (a xor b);
    outputs(6885) <= not b;
    outputs(6886) <= not b;
    outputs(6887) <= a xor b;
    outputs(6888) <= a xor b;
    outputs(6889) <= a xor b;
    outputs(6890) <= a and b;
    outputs(6891) <= a or b;
    outputs(6892) <= a and b;
    outputs(6893) <= not a or b;
    outputs(6894) <= a;
    outputs(6895) <= not a or b;
    outputs(6896) <= not a;
    outputs(6897) <= a xor b;
    outputs(6898) <= not (a xor b);
    outputs(6899) <= not b;
    outputs(6900) <= not (a and b);
    outputs(6901) <= not a or b;
    outputs(6902) <= a xor b;
    outputs(6903) <= not a or b;
    outputs(6904) <= b;
    outputs(6905) <= not (a xor b);
    outputs(6906) <= not (a xor b);
    outputs(6907) <= a xor b;
    outputs(6908) <= a xor b;
    outputs(6909) <= b;
    outputs(6910) <= a;
    outputs(6911) <= not b;
    outputs(6912) <= not a;
    outputs(6913) <= not (a xor b);
    outputs(6914) <= not b;
    outputs(6915) <= b;
    outputs(6916) <= a xor b;
    outputs(6917) <= a or b;
    outputs(6918) <= not b or a;
    outputs(6919) <= not b or a;
    outputs(6920) <= b;
    outputs(6921) <= a xor b;
    outputs(6922) <= not a;
    outputs(6923) <= not b;
    outputs(6924) <= a xor b;
    outputs(6925) <= b;
    outputs(6926) <= not (a xor b);
    outputs(6927) <= b;
    outputs(6928) <= a xor b;
    outputs(6929) <= a and b;
    outputs(6930) <= b;
    outputs(6931) <= b;
    outputs(6932) <= a or b;
    outputs(6933) <= not (a or b);
    outputs(6934) <= a and not b;
    outputs(6935) <= not (a xor b);
    outputs(6936) <= not (a and b);
    outputs(6937) <= a and not b;
    outputs(6938) <= not (a or b);
    outputs(6939) <= a xor b;
    outputs(6940) <= not a;
    outputs(6941) <= not a;
    outputs(6942) <= a xor b;
    outputs(6943) <= not (a or b);
    outputs(6944) <= not (a xor b);
    outputs(6945) <= not b;
    outputs(6946) <= not a or b;
    outputs(6947) <= a xor b;
    outputs(6948) <= not (a xor b);
    outputs(6949) <= not b or a;
    outputs(6950) <= a xor b;
    outputs(6951) <= b and not a;
    outputs(6952) <= not b or a;
    outputs(6953) <= not (a xor b);
    outputs(6954) <= 1'b0;
    outputs(6955) <= not b;
    outputs(6956) <= not b;
    outputs(6957) <= b;
    outputs(6958) <= b and not a;
    outputs(6959) <= not a or b;
    outputs(6960) <= a xor b;
    outputs(6961) <= b;
    outputs(6962) <= not a;
    outputs(6963) <= not b;
    outputs(6964) <= not a or b;
    outputs(6965) <= a;
    outputs(6966) <= a or b;
    outputs(6967) <= not b or a;
    outputs(6968) <= not b;
    outputs(6969) <= not (a and b);
    outputs(6970) <= not (a xor b);
    outputs(6971) <= b;
    outputs(6972) <= not b or a;
    outputs(6973) <= a or b;
    outputs(6974) <= a;
    outputs(6975) <= b and not a;
    outputs(6976) <= not b;
    outputs(6977) <= not (a and b);
    outputs(6978) <= a xor b;
    outputs(6979) <= 1'b1;
    outputs(6980) <= not (a and b);
    outputs(6981) <= a xor b;
    outputs(6982) <= b and not a;
    outputs(6983) <= a;
    outputs(6984) <= a;
    outputs(6985) <= a or b;
    outputs(6986) <= not (a and b);
    outputs(6987) <= a and b;
    outputs(6988) <= not a;
    outputs(6989) <= a and b;
    outputs(6990) <= b;
    outputs(6991) <= b;
    outputs(6992) <= b;
    outputs(6993) <= b and not a;
    outputs(6994) <= not (a xor b);
    outputs(6995) <= not b;
    outputs(6996) <= not b;
    outputs(6997) <= a xor b;
    outputs(6998) <= a xor b;
    outputs(6999) <= a;
    outputs(7000) <= not (a xor b);
    outputs(7001) <= 1'b0;
    outputs(7002) <= not a;
    outputs(7003) <= not a;
    outputs(7004) <= not b;
    outputs(7005) <= not a or b;
    outputs(7006) <= not b;
    outputs(7007) <= a or b;
    outputs(7008) <= b and not a;
    outputs(7009) <= not (a xor b);
    outputs(7010) <= not (a xor b);
    outputs(7011) <= not (a xor b);
    outputs(7012) <= not a;
    outputs(7013) <= not (a or b);
    outputs(7014) <= not (a xor b);
    outputs(7015) <= a;
    outputs(7016) <= a xor b;
    outputs(7017) <= not (a xor b);
    outputs(7018) <= not b or a;
    outputs(7019) <= not (a or b);
    outputs(7020) <= not (a xor b);
    outputs(7021) <= a and b;
    outputs(7022) <= a xor b;
    outputs(7023) <= a;
    outputs(7024) <= not a or b;
    outputs(7025) <= a and b;
    outputs(7026) <= not (a xor b);
    outputs(7027) <= a;
    outputs(7028) <= a;
    outputs(7029) <= a;
    outputs(7030) <= b;
    outputs(7031) <= not (a xor b);
    outputs(7032) <= b;
    outputs(7033) <= not (a xor b);
    outputs(7034) <= not (a xor b);
    outputs(7035) <= a xor b;
    outputs(7036) <= not (a xor b);
    outputs(7037) <= a;
    outputs(7038) <= b;
    outputs(7039) <= b;
    outputs(7040) <= a xor b;
    outputs(7041) <= not (a xor b);
    outputs(7042) <= not (a xor b);
    outputs(7043) <= not a or b;
    outputs(7044) <= a xor b;
    outputs(7045) <= not (a and b);
    outputs(7046) <= not (a xor b);
    outputs(7047) <= a or b;
    outputs(7048) <= a or b;
    outputs(7049) <= a and b;
    outputs(7050) <= not (a and b);
    outputs(7051) <= not b;
    outputs(7052) <= not (a xor b);
    outputs(7053) <= not b;
    outputs(7054) <= a xor b;
    outputs(7055) <= a or b;
    outputs(7056) <= not b or a;
    outputs(7057) <= not (a and b);
    outputs(7058) <= not b;
    outputs(7059) <= not (a and b);
    outputs(7060) <= not (a and b);
    outputs(7061) <= not b;
    outputs(7062) <= a xor b;
    outputs(7063) <= not b;
    outputs(7064) <= not (a xor b);
    outputs(7065) <= not (a xor b);
    outputs(7066) <= not b;
    outputs(7067) <= not b;
    outputs(7068) <= not (a and b);
    outputs(7069) <= not (a xor b);
    outputs(7070) <= a;
    outputs(7071) <= not b;
    outputs(7072) <= not a;
    outputs(7073) <= not (a and b);
    outputs(7074) <= a or b;
    outputs(7075) <= a xor b;
    outputs(7076) <= b;
    outputs(7077) <= a;
    outputs(7078) <= a;
    outputs(7079) <= a;
    outputs(7080) <= a xor b;
    outputs(7081) <= a xor b;
    outputs(7082) <= b and not a;
    outputs(7083) <= not b or a;
    outputs(7084) <= a xor b;
    outputs(7085) <= not (a xor b);
    outputs(7086) <= a xor b;
    outputs(7087) <= not b or a;
    outputs(7088) <= b;
    outputs(7089) <= not b;
    outputs(7090) <= not a;
    outputs(7091) <= not a;
    outputs(7092) <= not a;
    outputs(7093) <= a xor b;
    outputs(7094) <= a and not b;
    outputs(7095) <= a xor b;
    outputs(7096) <= not (a xor b);
    outputs(7097) <= not a;
    outputs(7098) <= not (a xor b);
    outputs(7099) <= a;
    outputs(7100) <= a;
    outputs(7101) <= a xor b;
    outputs(7102) <= not a or b;
    outputs(7103) <= not (a and b);
    outputs(7104) <= not b;
    outputs(7105) <= a and b;
    outputs(7106) <= a xor b;
    outputs(7107) <= a xor b;
    outputs(7108) <= not (a or b);
    outputs(7109) <= not (a xor b);
    outputs(7110) <= a and not b;
    outputs(7111) <= a;
    outputs(7112) <= a and b;
    outputs(7113) <= not b;
    outputs(7114) <= a xor b;
    outputs(7115) <= not a;
    outputs(7116) <= not (a xor b);
    outputs(7117) <= not (a xor b);
    outputs(7118) <= a xor b;
    outputs(7119) <= b;
    outputs(7120) <= not a;
    outputs(7121) <= not (a xor b);
    outputs(7122) <= not (a xor b);
    outputs(7123) <= not (a or b);
    outputs(7124) <= b;
    outputs(7125) <= not b or a;
    outputs(7126) <= not (a xor b);
    outputs(7127) <= not b or a;
    outputs(7128) <= not (a and b);
    outputs(7129) <= a xor b;
    outputs(7130) <= not a;
    outputs(7131) <= a xor b;
    outputs(7132) <= a xor b;
    outputs(7133) <= a;
    outputs(7134) <= not a;
    outputs(7135) <= b;
    outputs(7136) <= not (a xor b);
    outputs(7137) <= not a;
    outputs(7138) <= a or b;
    outputs(7139) <= not (a xor b);
    outputs(7140) <= not (a and b);
    outputs(7141) <= not (a xor b);
    outputs(7142) <= a;
    outputs(7143) <= not (a xor b);
    outputs(7144) <= b;
    outputs(7145) <= a xor b;
    outputs(7146) <= not b;
    outputs(7147) <= not (a xor b);
    outputs(7148) <= a xor b;
    outputs(7149) <= not a or b;
    outputs(7150) <= a xor b;
    outputs(7151) <= a;
    outputs(7152) <= a or b;
    outputs(7153) <= a xor b;
    outputs(7154) <= b;
    outputs(7155) <= not (a xor b);
    outputs(7156) <= not b or a;
    outputs(7157) <= not (a xor b);
    outputs(7158) <= a xor b;
    outputs(7159) <= not (a or b);
    outputs(7160) <= not (a xor b);
    outputs(7161) <= not (a xor b);
    outputs(7162) <= not a;
    outputs(7163) <= not b;
    outputs(7164) <= b and not a;
    outputs(7165) <= b;
    outputs(7166) <= not (a xor b);
    outputs(7167) <= not (a and b);
    outputs(7168) <= not a or b;
    outputs(7169) <= not a or b;
    outputs(7170) <= a xor b;
    outputs(7171) <= not (a or b);
    outputs(7172) <= a xor b;
    outputs(7173) <= not (a xor b);
    outputs(7174) <= b;
    outputs(7175) <= not (a and b);
    outputs(7176) <= a and b;
    outputs(7177) <= not (a xor b);
    outputs(7178) <= not b;
    outputs(7179) <= not a or b;
    outputs(7180) <= b;
    outputs(7181) <= a or b;
    outputs(7182) <= not (a xor b);
    outputs(7183) <= not (a xor b);
    outputs(7184) <= not (a xor b);
    outputs(7185) <= b;
    outputs(7186) <= not (a xor b);
    outputs(7187) <= a xor b;
    outputs(7188) <= not a;
    outputs(7189) <= a and b;
    outputs(7190) <= a xor b;
    outputs(7191) <= not a;
    outputs(7192) <= b;
    outputs(7193) <= not (a xor b);
    outputs(7194) <= a;
    outputs(7195) <= not b or a;
    outputs(7196) <= a xor b;
    outputs(7197) <= a xor b;
    outputs(7198) <= b;
    outputs(7199) <= not (a xor b);
    outputs(7200) <= not (a xor b);
    outputs(7201) <= not b or a;
    outputs(7202) <= a or b;
    outputs(7203) <= not (a xor b);
    outputs(7204) <= not (a xor b);
    outputs(7205) <= not (a and b);
    outputs(7206) <= a;
    outputs(7207) <= not b;
    outputs(7208) <= a;
    outputs(7209) <= not (a and b);
    outputs(7210) <= a and b;
    outputs(7211) <= a;
    outputs(7212) <= not (a xor b);
    outputs(7213) <= a xor b;
    outputs(7214) <= not b;
    outputs(7215) <= a;
    outputs(7216) <= not (a and b);
    outputs(7217) <= not b or a;
    outputs(7218) <= not (a xor b);
    outputs(7219) <= a and not b;
    outputs(7220) <= not (a xor b);
    outputs(7221) <= a or b;
    outputs(7222) <= b and not a;
    outputs(7223) <= not a or b;
    outputs(7224) <= a xor b;
    outputs(7225) <= not b or a;
    outputs(7226) <= b;
    outputs(7227) <= not b;
    outputs(7228) <= not a or b;
    outputs(7229) <= not a or b;
    outputs(7230) <= a;
    outputs(7231) <= b and not a;
    outputs(7232) <= a or b;
    outputs(7233) <= not b or a;
    outputs(7234) <= a xor b;
    outputs(7235) <= not (a xor b);
    outputs(7236) <= not b or a;
    outputs(7237) <= not (a xor b);
    outputs(7238) <= not (a xor b);
    outputs(7239) <= a;
    outputs(7240) <= a or b;
    outputs(7241) <= a xor b;
    outputs(7242) <= not (a xor b);
    outputs(7243) <= not b or a;
    outputs(7244) <= a or b;
    outputs(7245) <= not b;
    outputs(7246) <= a;
    outputs(7247) <= not (a or b);
    outputs(7248) <= a xor b;
    outputs(7249) <= b and not a;
    outputs(7250) <= a;
    outputs(7251) <= not b or a;
    outputs(7252) <= not b;
    outputs(7253) <= not (a xor b);
    outputs(7254) <= a xor b;
    outputs(7255) <= a and b;
    outputs(7256) <= a xor b;
    outputs(7257) <= not a;
    outputs(7258) <= a and not b;
    outputs(7259) <= not (a xor b);
    outputs(7260) <= not (a and b);
    outputs(7261) <= a;
    outputs(7262) <= not (a xor b);
    outputs(7263) <= a xor b;
    outputs(7264) <= not (a xor b);
    outputs(7265) <= a or b;
    outputs(7266) <= a;
    outputs(7267) <= not a or b;
    outputs(7268) <= a;
    outputs(7269) <= b;
    outputs(7270) <= a xor b;
    outputs(7271) <= not a or b;
    outputs(7272) <= a xor b;
    outputs(7273) <= a and not b;
    outputs(7274) <= a xor b;
    outputs(7275) <= a;
    outputs(7276) <= not (a and b);
    outputs(7277) <= not (a xor b);
    outputs(7278) <= a or b;
    outputs(7279) <= a xor b;
    outputs(7280) <= a or b;
    outputs(7281) <= not (a and b);
    outputs(7282) <= a xor b;
    outputs(7283) <= a xor b;
    outputs(7284) <= b;
    outputs(7285) <= a;
    outputs(7286) <= not a;
    outputs(7287) <= a xor b;
    outputs(7288) <= not b;
    outputs(7289) <= a and b;
    outputs(7290) <= not (a xor b);
    outputs(7291) <= b and not a;
    outputs(7292) <= a xor b;
    outputs(7293) <= not a;
    outputs(7294) <= not (a and b);
    outputs(7295) <= not a or b;
    outputs(7296) <= not (a xor b);
    outputs(7297) <= not (a xor b);
    outputs(7298) <= not b or a;
    outputs(7299) <= a xor b;
    outputs(7300) <= not b;
    outputs(7301) <= b;
    outputs(7302) <= a or b;
    outputs(7303) <= a xor b;
    outputs(7304) <= a or b;
    outputs(7305) <= not a;
    outputs(7306) <= a xor b;
    outputs(7307) <= a xor b;
    outputs(7308) <= a;
    outputs(7309) <= a and b;
    outputs(7310) <= a xor b;
    outputs(7311) <= not (a or b);
    outputs(7312) <= a or b;
    outputs(7313) <= a xor b;
    outputs(7314) <= not a or b;
    outputs(7315) <= a xor b;
    outputs(7316) <= not (a xor b);
    outputs(7317) <= not a or b;
    outputs(7318) <= a;
    outputs(7319) <= a or b;
    outputs(7320) <= b;
    outputs(7321) <= not (a or b);
    outputs(7322) <= not (a and b);
    outputs(7323) <= not b;
    outputs(7324) <= a;
    outputs(7325) <= a and not b;
    outputs(7326) <= a or b;
    outputs(7327) <= a xor b;
    outputs(7328) <= a and not b;
    outputs(7329) <= a xor b;
    outputs(7330) <= b;
    outputs(7331) <= not a;
    outputs(7332) <= a and not b;
    outputs(7333) <= b;
    outputs(7334) <= not a;
    outputs(7335) <= not (a xor b);
    outputs(7336) <= a and not b;
    outputs(7337) <= a xor b;
    outputs(7338) <= a;
    outputs(7339) <= b;
    outputs(7340) <= a xor b;
    outputs(7341) <= not (a or b);
    outputs(7342) <= b;
    outputs(7343) <= not (a xor b);
    outputs(7344) <= not (a or b);
    outputs(7345) <= not (a xor b);
    outputs(7346) <= a;
    outputs(7347) <= b;
    outputs(7348) <= not a or b;
    outputs(7349) <= not b;
    outputs(7350) <= a xor b;
    outputs(7351) <= not a;
    outputs(7352) <= a;
    outputs(7353) <= not (a or b);
    outputs(7354) <= a xor b;
    outputs(7355) <= not a or b;
    outputs(7356) <= not (a xor b);
    outputs(7357) <= a and b;
    outputs(7358) <= not (a xor b);
    outputs(7359) <= a and b;
    outputs(7360) <= not b;
    outputs(7361) <= not b or a;
    outputs(7362) <= not a or b;
    outputs(7363) <= a xor b;
    outputs(7364) <= b and not a;
    outputs(7365) <= not (a xor b);
    outputs(7366) <= not b;
    outputs(7367) <= not (a xor b);
    outputs(7368) <= b;
    outputs(7369) <= a xor b;
    outputs(7370) <= a;
    outputs(7371) <= a;
    outputs(7372) <= a or b;
    outputs(7373) <= not b;
    outputs(7374) <= not b;
    outputs(7375) <= not (a xor b);
    outputs(7376) <= b;
    outputs(7377) <= not (a and b);
    outputs(7378) <= b;
    outputs(7379) <= not a;
    outputs(7380) <= not (a or b);
    outputs(7381) <= a and not b;
    outputs(7382) <= b;
    outputs(7383) <= a and not b;
    outputs(7384) <= not (a xor b);
    outputs(7385) <= a xor b;
    outputs(7386) <= a and b;
    outputs(7387) <= a;
    outputs(7388) <= a and not b;
    outputs(7389) <= a or b;
    outputs(7390) <= a or b;
    outputs(7391) <= not (a or b);
    outputs(7392) <= not b;
    outputs(7393) <= a xor b;
    outputs(7394) <= not a;
    outputs(7395) <= not b;
    outputs(7396) <= not a or b;
    outputs(7397) <= a;
    outputs(7398) <= a xor b;
    outputs(7399) <= b;
    outputs(7400) <= a xor b;
    outputs(7401) <= a;
    outputs(7402) <= a xor b;
    outputs(7403) <= b;
    outputs(7404) <= a xor b;
    outputs(7405) <= not (a xor b);
    outputs(7406) <= b and not a;
    outputs(7407) <= not b;
    outputs(7408) <= a xor b;
    outputs(7409) <= not b or a;
    outputs(7410) <= a or b;
    outputs(7411) <= a and not b;
    outputs(7412) <= a or b;
    outputs(7413) <= a xor b;
    outputs(7414) <= a or b;
    outputs(7415) <= a xor b;
    outputs(7416) <= a xor b;
    outputs(7417) <= a xor b;
    outputs(7418) <= not b;
    outputs(7419) <= a xor b;
    outputs(7420) <= a xor b;
    outputs(7421) <= a xor b;
    outputs(7422) <= a;
    outputs(7423) <= a xor b;
    outputs(7424) <= not a or b;
    outputs(7425) <= b and not a;
    outputs(7426) <= not (a xor b);
    outputs(7427) <= not (a xor b);
    outputs(7428) <= a xor b;
    outputs(7429) <= a xor b;
    outputs(7430) <= not a;
    outputs(7431) <= a and not b;
    outputs(7432) <= not b;
    outputs(7433) <= a xor b;
    outputs(7434) <= a and not b;
    outputs(7435) <= not a;
    outputs(7436) <= not b;
    outputs(7437) <= b and not a;
    outputs(7438) <= a xor b;
    outputs(7439) <= not a;
    outputs(7440) <= a;
    outputs(7441) <= not (a and b);
    outputs(7442) <= a;
    outputs(7443) <= not (a xor b);
    outputs(7444) <= a xor b;
    outputs(7445) <= not a or b;
    outputs(7446) <= a xor b;
    outputs(7447) <= not (a xor b);
    outputs(7448) <= not (a xor b);
    outputs(7449) <= a xor b;
    outputs(7450) <= a;
    outputs(7451) <= not a;
    outputs(7452) <= not b or a;
    outputs(7453) <= not (a and b);
    outputs(7454) <= not a;
    outputs(7455) <= not b;
    outputs(7456) <= a and b;
    outputs(7457) <= not (a xor b);
    outputs(7458) <= a and b;
    outputs(7459) <= not (a and b);
    outputs(7460) <= a xor b;
    outputs(7461) <= not b;
    outputs(7462) <= not a;
    outputs(7463) <= a xor b;
    outputs(7464) <= a and not b;
    outputs(7465) <= not a;
    outputs(7466) <= not (a and b);
    outputs(7467) <= not (a xor b);
    outputs(7468) <= a xor b;
    outputs(7469) <= not (a xor b);
    outputs(7470) <= a and b;
    outputs(7471) <= a xor b;
    outputs(7472) <= b;
    outputs(7473) <= a;
    outputs(7474) <= not a;
    outputs(7475) <= a xor b;
    outputs(7476) <= a xor b;
    outputs(7477) <= not a;
    outputs(7478) <= not (a and b);
    outputs(7479) <= not (a xor b);
    outputs(7480) <= not a or b;
    outputs(7481) <= b and not a;
    outputs(7482) <= b and not a;
    outputs(7483) <= not b;
    outputs(7484) <= a xor b;
    outputs(7485) <= not (a or b);
    outputs(7486) <= a or b;
    outputs(7487) <= a xor b;
    outputs(7488) <= not (a or b);
    outputs(7489) <= a;
    outputs(7490) <= not (a and b);
    outputs(7491) <= a and b;
    outputs(7492) <= not (a xor b);
    outputs(7493) <= not a;
    outputs(7494) <= a xor b;
    outputs(7495) <= a;
    outputs(7496) <= not (a xor b);
    outputs(7497) <= not (a xor b);
    outputs(7498) <= not a;
    outputs(7499) <= not a;
    outputs(7500) <= not (a xor b);
    outputs(7501) <= b and not a;
    outputs(7502) <= not a;
    outputs(7503) <= a xor b;
    outputs(7504) <= not (a xor b);
    outputs(7505) <= not a or b;
    outputs(7506) <= not a;
    outputs(7507) <= not a;
    outputs(7508) <= b and not a;
    outputs(7509) <= b and not a;
    outputs(7510) <= not (a and b);
    outputs(7511) <= a and not b;
    outputs(7512) <= a or b;
    outputs(7513) <= a xor b;
    outputs(7514) <= b;
    outputs(7515) <= a or b;
    outputs(7516) <= not (a or b);
    outputs(7517) <= a xor b;
    outputs(7518) <= not (a xor b);
    outputs(7519) <= a and not b;
    outputs(7520) <= not a;
    outputs(7521) <= not (a xor b);
    outputs(7522) <= b;
    outputs(7523) <= not a or b;
    outputs(7524) <= not (a xor b);
    outputs(7525) <= not (a and b);
    outputs(7526) <= not (a xor b);
    outputs(7527) <= not b;
    outputs(7528) <= b;
    outputs(7529) <= not b;
    outputs(7530) <= a;
    outputs(7531) <= not b;
    outputs(7532) <= a or b;
    outputs(7533) <= not (a xor b);
    outputs(7534) <= not (a xor b);
    outputs(7535) <= not (a or b);
    outputs(7536) <= not a;
    outputs(7537) <= a xor b;
    outputs(7538) <= not a;
    outputs(7539) <= not a or b;
    outputs(7540) <= b;
    outputs(7541) <= not (a and b);
    outputs(7542) <= a and not b;
    outputs(7543) <= not a;
    outputs(7544) <= not b or a;
    outputs(7545) <= not b or a;
    outputs(7546) <= not a;
    outputs(7547) <= not (a xor b);
    outputs(7548) <= not (a and b);
    outputs(7549) <= b and not a;
    outputs(7550) <= a xor b;
    outputs(7551) <= a;
    outputs(7552) <= not b;
    outputs(7553) <= not (a xor b);
    outputs(7554) <= not a;
    outputs(7555) <= not b or a;
    outputs(7556) <= a or b;
    outputs(7557) <= not a or b;
    outputs(7558) <= not a;
    outputs(7559) <= a;
    outputs(7560) <= a and b;
    outputs(7561) <= not b;
    outputs(7562) <= b and not a;
    outputs(7563) <= not (a or b);
    outputs(7564) <= a and not b;
    outputs(7565) <= a xor b;
    outputs(7566) <= not (a xor b);
    outputs(7567) <= a and not b;
    outputs(7568) <= a;
    outputs(7569) <= a and b;
    outputs(7570) <= not (a xor b);
    outputs(7571) <= a;
    outputs(7572) <= not b;
    outputs(7573) <= not a;
    outputs(7574) <= not a;
    outputs(7575) <= not (a xor b);
    outputs(7576) <= a xor b;
    outputs(7577) <= not b;
    outputs(7578) <= not a;
    outputs(7579) <= not (a xor b);
    outputs(7580) <= a xor b;
    outputs(7581) <= not a;
    outputs(7582) <= a xor b;
    outputs(7583) <= not b or a;
    outputs(7584) <= not b;
    outputs(7585) <= not a or b;
    outputs(7586) <= not b;
    outputs(7587) <= b;
    outputs(7588) <= not (a xor b);
    outputs(7589) <= b;
    outputs(7590) <= b and not a;
    outputs(7591) <= a or b;
    outputs(7592) <= not b;
    outputs(7593) <= not b or a;
    outputs(7594) <= not (a xor b);
    outputs(7595) <= a and b;
    outputs(7596) <= not (a or b);
    outputs(7597) <= a xor b;
    outputs(7598) <= 1'b1;
    outputs(7599) <= not (a and b);
    outputs(7600) <= a;
    outputs(7601) <= not (a xor b);
    outputs(7602) <= a or b;
    outputs(7603) <= b;
    outputs(7604) <= 1'b1;
    outputs(7605) <= not (a xor b);
    outputs(7606) <= a;
    outputs(7607) <= not a or b;
    outputs(7608) <= not a;
    outputs(7609) <= not (a xor b);
    outputs(7610) <= a or b;
    outputs(7611) <= not (a xor b);
    outputs(7612) <= not a;
    outputs(7613) <= not a;
    outputs(7614) <= a xor b;
    outputs(7615) <= a xor b;
    outputs(7616) <= a and b;
    outputs(7617) <= a xor b;
    outputs(7618) <= not (a xor b);
    outputs(7619) <= a;
    outputs(7620) <= not (a xor b);
    outputs(7621) <= b;
    outputs(7622) <= not (a xor b);
    outputs(7623) <= b;
    outputs(7624) <= b;
    outputs(7625) <= not a or b;
    outputs(7626) <= b;
    outputs(7627) <= a;
    outputs(7628) <= not (a xor b);
    outputs(7629) <= a xor b;
    outputs(7630) <= not a;
    outputs(7631) <= a;
    outputs(7632) <= not (a xor b);
    outputs(7633) <= not a or b;
    outputs(7634) <= a;
    outputs(7635) <= not b or a;
    outputs(7636) <= a xor b;
    outputs(7637) <= a xor b;
    outputs(7638) <= a xor b;
    outputs(7639) <= a xor b;
    outputs(7640) <= not a;
    outputs(7641) <= not b;
    outputs(7642) <= not (a xor b);
    outputs(7643) <= a or b;
    outputs(7644) <= not b or a;
    outputs(7645) <= a;
    outputs(7646) <= a xor b;
    outputs(7647) <= b;
    outputs(7648) <= not (a xor b);
    outputs(7649) <= not (a or b);
    outputs(7650) <= not b;
    outputs(7651) <= not (a and b);
    outputs(7652) <= not b;
    outputs(7653) <= a and not b;
    outputs(7654) <= not (a and b);
    outputs(7655) <= not a or b;
    outputs(7656) <= a or b;
    outputs(7657) <= a xor b;
    outputs(7658) <= not b;
    outputs(7659) <= a xor b;
    outputs(7660) <= not (a xor b);
    outputs(7661) <= 1'b1;
    outputs(7662) <= a xor b;
    outputs(7663) <= not (a and b);
    outputs(7664) <= not (a xor b);
    outputs(7665) <= a or b;
    outputs(7666) <= a or b;
    outputs(7667) <= 1'b1;
    outputs(7668) <= not a;
    outputs(7669) <= b;
    outputs(7670) <= b;
    outputs(7671) <= not (a and b);
    outputs(7672) <= a;
    outputs(7673) <= a xor b;
    outputs(7674) <= b and not a;
    outputs(7675) <= b and not a;
    outputs(7676) <= a;
    outputs(7677) <= b;
    outputs(7678) <= not a;
    outputs(7679) <= not (a xor b);
    outputs(7680) <= a;
    outputs(7681) <= not (a xor b);
    outputs(7682) <= a;
    outputs(7683) <= a and b;
    outputs(7684) <= not (a xor b);
    outputs(7685) <= a;
    outputs(7686) <= not b;
    outputs(7687) <= a and b;
    outputs(7688) <= a and b;
    outputs(7689) <= a xor b;
    outputs(7690) <= not (a or b);
    outputs(7691) <= not (a xor b);
    outputs(7692) <= a;
    outputs(7693) <= a;
    outputs(7694) <= a xor b;
    outputs(7695) <= not a;
    outputs(7696) <= not a;
    outputs(7697) <= not (a xor b);
    outputs(7698) <= not a or b;
    outputs(7699) <= a;
    outputs(7700) <= not (a xor b);
    outputs(7701) <= a xor b;
    outputs(7702) <= not b;
    outputs(7703) <= not b;
    outputs(7704) <= not (a xor b);
    outputs(7705) <= a xor b;
    outputs(7706) <= a xor b;
    outputs(7707) <= not a;
    outputs(7708) <= a xor b;
    outputs(7709) <= a xor b;
    outputs(7710) <= b;
    outputs(7711) <= b;
    outputs(7712) <= b and not a;
    outputs(7713) <= not a;
    outputs(7714) <= a xor b;
    outputs(7715) <= b;
    outputs(7716) <= b and not a;
    outputs(7717) <= b;
    outputs(7718) <= a xor b;
    outputs(7719) <= a xor b;
    outputs(7720) <= b;
    outputs(7721) <= b and not a;
    outputs(7722) <= not (a xor b);
    outputs(7723) <= a;
    outputs(7724) <= a;
    outputs(7725) <= a;
    outputs(7726) <= b;
    outputs(7727) <= a xor b;
    outputs(7728) <= not (a and b);
    outputs(7729) <= not b;
    outputs(7730) <= not a;
    outputs(7731) <= b and not a;
    outputs(7732) <= b;
    outputs(7733) <= not (a xor b);
    outputs(7734) <= not b;
    outputs(7735) <= a xor b;
    outputs(7736) <= a xor b;
    outputs(7737) <= b and not a;
    outputs(7738) <= a xor b;
    outputs(7739) <= not (a or b);
    outputs(7740) <= a xor b;
    outputs(7741) <= not a;
    outputs(7742) <= not (a xor b);
    outputs(7743) <= a and b;
    outputs(7744) <= b and not a;
    outputs(7745) <= not b;
    outputs(7746) <= a xor b;
    outputs(7747) <= a xor b;
    outputs(7748) <= a;
    outputs(7749) <= a xor b;
    outputs(7750) <= not (a xor b);
    outputs(7751) <= a and not b;
    outputs(7752) <= b and not a;
    outputs(7753) <= not (a xor b);
    outputs(7754) <= b;
    outputs(7755) <= not a;
    outputs(7756) <= b;
    outputs(7757) <= b;
    outputs(7758) <= a xor b;
    outputs(7759) <= not (a xor b);
    outputs(7760) <= b;
    outputs(7761) <= not (a xor b);
    outputs(7762) <= a and b;
    outputs(7763) <= a xor b;
    outputs(7764) <= not (a xor b);
    outputs(7765) <= not a;
    outputs(7766) <= not (a and b);
    outputs(7767) <= a xor b;
    outputs(7768) <= not b;
    outputs(7769) <= a and not b;
    outputs(7770) <= a;
    outputs(7771) <= a xor b;
    outputs(7772) <= a and not b;
    outputs(7773) <= not (a and b);
    outputs(7774) <= a;
    outputs(7775) <= not b;
    outputs(7776) <= not (a or b);
    outputs(7777) <= not (a xor b);
    outputs(7778) <= a;
    outputs(7779) <= not a;
    outputs(7780) <= not b;
    outputs(7781) <= b and not a;
    outputs(7782) <= not (a xor b);
    outputs(7783) <= a xor b;
    outputs(7784) <= a xor b;
    outputs(7785) <= a xor b;
    outputs(7786) <= b;
    outputs(7787) <= not (a xor b);
    outputs(7788) <= not b;
    outputs(7789) <= not b;
    outputs(7790) <= a;
    outputs(7791) <= not (a xor b);
    outputs(7792) <= a;
    outputs(7793) <= a xor b;
    outputs(7794) <= not b or a;
    outputs(7795) <= b and not a;
    outputs(7796) <= b and not a;
    outputs(7797) <= a xor b;
    outputs(7798) <= not (a or b);
    outputs(7799) <= a and b;
    outputs(7800) <= a xor b;
    outputs(7801) <= not a;
    outputs(7802) <= not b;
    outputs(7803) <= not a;
    outputs(7804) <= not (a xor b);
    outputs(7805) <= a xor b;
    outputs(7806) <= not a;
    outputs(7807) <= not (a or b);
    outputs(7808) <= a and b;
    outputs(7809) <= a xor b;
    outputs(7810) <= not b;
    outputs(7811) <= a;
    outputs(7812) <= b;
    outputs(7813) <= not a;
    outputs(7814) <= not b;
    outputs(7815) <= a;
    outputs(7816) <= not (a xor b);
    outputs(7817) <= not (a or b);
    outputs(7818) <= b;
    outputs(7819) <= b and not a;
    outputs(7820) <= a;
    outputs(7821) <= not (a xor b);
    outputs(7822) <= a or b;
    outputs(7823) <= not b;
    outputs(7824) <= a xor b;
    outputs(7825) <= not (a xor b);
    outputs(7826) <= a xor b;
    outputs(7827) <= a and b;
    outputs(7828) <= not (a xor b);
    outputs(7829) <= not (a xor b);
    outputs(7830) <= a and not b;
    outputs(7831) <= not b;
    outputs(7832) <= a xor b;
    outputs(7833) <= not (a xor b);
    outputs(7834) <= b;
    outputs(7835) <= a and b;
    outputs(7836) <= a;
    outputs(7837) <= a xor b;
    outputs(7838) <= not b;
    outputs(7839) <= not a;
    outputs(7840) <= not a;
    outputs(7841) <= b;
    outputs(7842) <= b;
    outputs(7843) <= b;
    outputs(7844) <= a;
    outputs(7845) <= not (a or b);
    outputs(7846) <= b;
    outputs(7847) <= a;
    outputs(7848) <= a;
    outputs(7849) <= a xor b;
    outputs(7850) <= not (a xor b);
    outputs(7851) <= a and not b;
    outputs(7852) <= a and not b;
    outputs(7853) <= a;
    outputs(7854) <= not (a or b);
    outputs(7855) <= a xor b;
    outputs(7856) <= not a;
    outputs(7857) <= a;
    outputs(7858) <= a xor b;
    outputs(7859) <= a xor b;
    outputs(7860) <= a or b;
    outputs(7861) <= b;
    outputs(7862) <= b and not a;
    outputs(7863) <= a xor b;
    outputs(7864) <= a;
    outputs(7865) <= not (a xor b);
    outputs(7866) <= a xor b;
    outputs(7867) <= not a;
    outputs(7868) <= not (a or b);
    outputs(7869) <= not b;
    outputs(7870) <= not (a xor b);
    outputs(7871) <= a and not b;
    outputs(7872) <= not a;
    outputs(7873) <= b and not a;
    outputs(7874) <= a;
    outputs(7875) <= b;
    outputs(7876) <= a or b;
    outputs(7877) <= a;
    outputs(7878) <= b;
    outputs(7879) <= not (a xor b);
    outputs(7880) <= not a;
    outputs(7881) <= not a;
    outputs(7882) <= a xor b;
    outputs(7883) <= not (a xor b);
    outputs(7884) <= not a;
    outputs(7885) <= not b;
    outputs(7886) <= b;
    outputs(7887) <= a;
    outputs(7888) <= not a;
    outputs(7889) <= not b;
    outputs(7890) <= a xor b;
    outputs(7891) <= a xor b;
    outputs(7892) <= not a or b;
    outputs(7893) <= a xor b;
    outputs(7894) <= a xor b;
    outputs(7895) <= a and not b;
    outputs(7896) <= b;
    outputs(7897) <= a;
    outputs(7898) <= a;
    outputs(7899) <= not b;
    outputs(7900) <= not a;
    outputs(7901) <= not a;
    outputs(7902) <= not (a and b);
    outputs(7903) <= not b;
    outputs(7904) <= not b;
    outputs(7905) <= a xor b;
    outputs(7906) <= b;
    outputs(7907) <= not (a xor b);
    outputs(7908) <= a;
    outputs(7909) <= not a or b;
    outputs(7910) <= a xor b;
    outputs(7911) <= a and not b;
    outputs(7912) <= a and b;
    outputs(7913) <= not (a or b);
    outputs(7914) <= a and b;
    outputs(7915) <= b and not a;
    outputs(7916) <= not b or a;
    outputs(7917) <= not (a xor b);
    outputs(7918) <= a xor b;
    outputs(7919) <= a;
    outputs(7920) <= not (a xor b);
    outputs(7921) <= not a;
    outputs(7922) <= not (a xor b);
    outputs(7923) <= not a;
    outputs(7924) <= a;
    outputs(7925) <= a or b;
    outputs(7926) <= not a;
    outputs(7927) <= not b;
    outputs(7928) <= a;
    outputs(7929) <= not (a xor b);
    outputs(7930) <= a xor b;
    outputs(7931) <= not (a or b);
    outputs(7932) <= b;
    outputs(7933) <= not a;
    outputs(7934) <= a;
    outputs(7935) <= not b;
    outputs(7936) <= not b;
    outputs(7937) <= a xor b;
    outputs(7938) <= a;
    outputs(7939) <= not a;
    outputs(7940) <= not a;
    outputs(7941) <= a;
    outputs(7942) <= a and b;
    outputs(7943) <= not (a xor b);
    outputs(7944) <= not (a xor b);
    outputs(7945) <= b;
    outputs(7946) <= a xor b;
    outputs(7947) <= a xor b;
    outputs(7948) <= not b;
    outputs(7949) <= not (a xor b);
    outputs(7950) <= not (a and b);
    outputs(7951) <= not (a xor b);
    outputs(7952) <= not (a or b);
    outputs(7953) <= a xor b;
    outputs(7954) <= not (a xor b);
    outputs(7955) <= a;
    outputs(7956) <= not (a xor b);
    outputs(7957) <= a xor b;
    outputs(7958) <= a xor b;
    outputs(7959) <= not (a xor b);
    outputs(7960) <= not b or a;
    outputs(7961) <= not (a xor b);
    outputs(7962) <= b;
    outputs(7963) <= b;
    outputs(7964) <= a;
    outputs(7965) <= b;
    outputs(7966) <= a xor b;
    outputs(7967) <= a and not b;
    outputs(7968) <= not (a xor b);
    outputs(7969) <= not b;
    outputs(7970) <= a and not b;
    outputs(7971) <= not a;
    outputs(7972) <= not (a xor b);
    outputs(7973) <= a xor b;
    outputs(7974) <= not b;
    outputs(7975) <= not b;
    outputs(7976) <= a and not b;
    outputs(7977) <= a xor b;
    outputs(7978) <= a and b;
    outputs(7979) <= a xor b;
    outputs(7980) <= a or b;
    outputs(7981) <= not (a or b);
    outputs(7982) <= a xor b;
    outputs(7983) <= not a;
    outputs(7984) <= not a;
    outputs(7985) <= a xor b;
    outputs(7986) <= a xor b;
    outputs(7987) <= a xor b;
    outputs(7988) <= not a;
    outputs(7989) <= a;
    outputs(7990) <= b;
    outputs(7991) <= a or b;
    outputs(7992) <= b and not a;
    outputs(7993) <= b;
    outputs(7994) <= not (a and b);
    outputs(7995) <= not b or a;
    outputs(7996) <= not (a and b);
    outputs(7997) <= b;
    outputs(7998) <= b;
    outputs(7999) <= not (a xor b);
    outputs(8000) <= not (a and b);
    outputs(8001) <= a xor b;
    outputs(8002) <= not b;
    outputs(8003) <= a and b;
    outputs(8004) <= a xor b;
    outputs(8005) <= a;
    outputs(8006) <= a;
    outputs(8007) <= not b;
    outputs(8008) <= a;
    outputs(8009) <= a and b;
    outputs(8010) <= not (a xor b);
    outputs(8011) <= a xor b;
    outputs(8012) <= not b;
    outputs(8013) <= a xor b;
    outputs(8014) <= not (a or b);
    outputs(8015) <= a xor b;
    outputs(8016) <= not (a xor b);
    outputs(8017) <= not b;
    outputs(8018) <= not a;
    outputs(8019) <= not (a or b);
    outputs(8020) <= b;
    outputs(8021) <= a;
    outputs(8022) <= a and b;
    outputs(8023) <= a;
    outputs(8024) <= not (a or b);
    outputs(8025) <= a xor b;
    outputs(8026) <= not (a and b);
    outputs(8027) <= not a;
    outputs(8028) <= a xor b;
    outputs(8029) <= not b;
    outputs(8030) <= not (a xor b);
    outputs(8031) <= a xor b;
    outputs(8032) <= b;
    outputs(8033) <= not b;
    outputs(8034) <= a xor b;
    outputs(8035) <= a and not b;
    outputs(8036) <= b and not a;
    outputs(8037) <= not b;
    outputs(8038) <= a xor b;
    outputs(8039) <= b;
    outputs(8040) <= not a or b;
    outputs(8041) <= not (a xor b);
    outputs(8042) <= a xor b;
    outputs(8043) <= not (a or b);
    outputs(8044) <= b;
    outputs(8045) <= a and b;
    outputs(8046) <= a and b;
    outputs(8047) <= a xor b;
    outputs(8048) <= not b;
    outputs(8049) <= not (a xor b);
    outputs(8050) <= not a;
    outputs(8051) <= a and b;
    outputs(8052) <= not b;
    outputs(8053) <= b;
    outputs(8054) <= not (a xor b);
    outputs(8055) <= a and not b;
    outputs(8056) <= a and not b;
    outputs(8057) <= a xor b;
    outputs(8058) <= not (a xor b);
    outputs(8059) <= b and not a;
    outputs(8060) <= b;
    outputs(8061) <= not (a or b);
    outputs(8062) <= a xor b;
    outputs(8063) <= b;
    outputs(8064) <= b;
    outputs(8065) <= not (a xor b);
    outputs(8066) <= not b;
    outputs(8067) <= not (a xor b);
    outputs(8068) <= a;
    outputs(8069) <= b;
    outputs(8070) <= a;
    outputs(8071) <= not b;
    outputs(8072) <= not a or b;
    outputs(8073) <= b;
    outputs(8074) <= a xor b;
    outputs(8075) <= a xor b;
    outputs(8076) <= b;
    outputs(8077) <= a xor b;
    outputs(8078) <= a;
    outputs(8079) <= not (a xor b);
    outputs(8080) <= not (a xor b);
    outputs(8081) <= not (a xor b);
    outputs(8082) <= a and not b;
    outputs(8083) <= a;
    outputs(8084) <= not b;
    outputs(8085) <= not b;
    outputs(8086) <= a;
    outputs(8087) <= a or b;
    outputs(8088) <= a;
    outputs(8089) <= not a or b;
    outputs(8090) <= a;
    outputs(8091) <= b;
    outputs(8092) <= not (a xor b);
    outputs(8093) <= not b;
    outputs(8094) <= b;
    outputs(8095) <= a;
    outputs(8096) <= a xor b;
    outputs(8097) <= a xor b;
    outputs(8098) <= not b;
    outputs(8099) <= not a;
    outputs(8100) <= a;
    outputs(8101) <= b;
    outputs(8102) <= a;
    outputs(8103) <= a;
    outputs(8104) <= not (a and b);
    outputs(8105) <= a or b;
    outputs(8106) <= not (a xor b);
    outputs(8107) <= a xor b;
    outputs(8108) <= not (a xor b);
    outputs(8109) <= a xor b;
    outputs(8110) <= b;
    outputs(8111) <= a;
    outputs(8112) <= a and b;
    outputs(8113) <= b;
    outputs(8114) <= not (a or b);
    outputs(8115) <= not (a xor b);
    outputs(8116) <= b;
    outputs(8117) <= not (a and b);
    outputs(8118) <= not (a or b);
    outputs(8119) <= not (a xor b);
    outputs(8120) <= a;
    outputs(8121) <= not a;
    outputs(8122) <= not (a xor b);
    outputs(8123) <= not a or b;
    outputs(8124) <= a or b;
    outputs(8125) <= b;
    outputs(8126) <= not a or b;
    outputs(8127) <= b;
    outputs(8128) <= a xor b;
    outputs(8129) <= not (a xor b);
    outputs(8130) <= not b;
    outputs(8131) <= a;
    outputs(8132) <= a and not b;
    outputs(8133) <= a xor b;
    outputs(8134) <= not b;
    outputs(8135) <= not (a xor b);
    outputs(8136) <= a xor b;
    outputs(8137) <= not b;
    outputs(8138) <= a and not b;
    outputs(8139) <= not b;
    outputs(8140) <= not a;
    outputs(8141) <= not (a xor b);
    outputs(8142) <= a;
    outputs(8143) <= a xor b;
    outputs(8144) <= a;
    outputs(8145) <= not b;
    outputs(8146) <= b;
    outputs(8147) <= b;
    outputs(8148) <= not (a xor b);
    outputs(8149) <= a xor b;
    outputs(8150) <= not (a xor b);
    outputs(8151) <= not (a xor b);
    outputs(8152) <= not b;
    outputs(8153) <= not (a xor b);
    outputs(8154) <= not (a xor b);
    outputs(8155) <= a;
    outputs(8156) <= b;
    outputs(8157) <= a and not b;
    outputs(8158) <= not (a and b);
    outputs(8159) <= not b;
    outputs(8160) <= b;
    outputs(8161) <= not b;
    outputs(8162) <= not (a xor b);
    outputs(8163) <= not (a or b);
    outputs(8164) <= a;
    outputs(8165) <= not b;
    outputs(8166) <= a and b;
    outputs(8167) <= not a;
    outputs(8168) <= a;
    outputs(8169) <= a xor b;
    outputs(8170) <= not a;
    outputs(8171) <= not b;
    outputs(8172) <= a xor b;
    outputs(8173) <= a xor b;
    outputs(8174) <= not (a or b);
    outputs(8175) <= not (a xor b);
    outputs(8176) <= a and not b;
    outputs(8177) <= a and not b;
    outputs(8178) <= b;
    outputs(8179) <= a and not b;
    outputs(8180) <= not (a xor b);
    outputs(8181) <= b;
    outputs(8182) <= not (a xor b);
    outputs(8183) <= not b;
    outputs(8184) <= not b;
    outputs(8185) <= a;
    outputs(8186) <= not b;
    outputs(8187) <= not b or a;
    outputs(8188) <= not a or b;
    outputs(8189) <= not a;
    outputs(8190) <= b;
    outputs(8191) <= not (a xor b);
    outputs(8192) <= b and not a;
    outputs(8193) <= a or b;
    outputs(8194) <= b;
    outputs(8195) <= b;
    outputs(8196) <= not b or a;
    outputs(8197) <= a;
    outputs(8198) <= not a or b;
    outputs(8199) <= not a;
    outputs(8200) <= not b;
    outputs(8201) <= not (a xor b);
    outputs(8202) <= not a;
    outputs(8203) <= not (a or b);
    outputs(8204) <= not b;
    outputs(8205) <= not (a or b);
    outputs(8206) <= not b;
    outputs(8207) <= not (a and b);
    outputs(8208) <= b and not a;
    outputs(8209) <= a;
    outputs(8210) <= a xor b;
    outputs(8211) <= a xor b;
    outputs(8212) <= not b or a;
    outputs(8213) <= b;
    outputs(8214) <= not (a xor b);
    outputs(8215) <= not b or a;
    outputs(8216) <= a xor b;
    outputs(8217) <= not (a xor b);
    outputs(8218) <= a;
    outputs(8219) <= a xor b;
    outputs(8220) <= a;
    outputs(8221) <= not (a or b);
    outputs(8222) <= not a;
    outputs(8223) <= a or b;
    outputs(8224) <= not (a xor b);
    outputs(8225) <= not a;
    outputs(8226) <= a xor b;
    outputs(8227) <= a xor b;
    outputs(8228) <= not a or b;
    outputs(8229) <= a;
    outputs(8230) <= not (a or b);
    outputs(8231) <= b;
    outputs(8232) <= a xor b;
    outputs(8233) <= a;
    outputs(8234) <= not (a and b);
    outputs(8235) <= a xor b;
    outputs(8236) <= b;
    outputs(8237) <= not (a and b);
    outputs(8238) <= b;
    outputs(8239) <= not b;
    outputs(8240) <= a and b;
    outputs(8241) <= a xor b;
    outputs(8242) <= a xor b;
    outputs(8243) <= not b;
    outputs(8244) <= 1'b0;
    outputs(8245) <= not (a xor b);
    outputs(8246) <= not (a xor b);
    outputs(8247) <= not (a and b);
    outputs(8248) <= not b;
    outputs(8249) <= not (a or b);
    outputs(8250) <= a or b;
    outputs(8251) <= b and not a;
    outputs(8252) <= b;
    outputs(8253) <= a xor b;
    outputs(8254) <= not b;
    outputs(8255) <= not (a xor b);
    outputs(8256) <= not b;
    outputs(8257) <= b;
    outputs(8258) <= not b;
    outputs(8259) <= not (a and b);
    outputs(8260) <= a and b;
    outputs(8261) <= a xor b;
    outputs(8262) <= a xor b;
    outputs(8263) <= not (a or b);
    outputs(8264) <= not (a xor b);
    outputs(8265) <= a;
    outputs(8266) <= a;
    outputs(8267) <= b;
    outputs(8268) <= not b;
    outputs(8269) <= not b;
    outputs(8270) <= not (a xor b);
    outputs(8271) <= a xor b;
    outputs(8272) <= not b;
    outputs(8273) <= not (a or b);
    outputs(8274) <= not b or a;
    outputs(8275) <= a;
    outputs(8276) <= not a or b;
    outputs(8277) <= not (a or b);
    outputs(8278) <= a xor b;
    outputs(8279) <= not (a or b);
    outputs(8280) <= not b;
    outputs(8281) <= a xor b;
    outputs(8282) <= a and b;
    outputs(8283) <= not (a xor b);
    outputs(8284) <= a;
    outputs(8285) <= not a;
    outputs(8286) <= not b or a;
    outputs(8287) <= a and not b;
    outputs(8288) <= a and b;
    outputs(8289) <= a;
    outputs(8290) <= not b;
    outputs(8291) <= not (a xor b);
    outputs(8292) <= a xor b;
    outputs(8293) <= not (a xor b);
    outputs(8294) <= not (a and b);
    outputs(8295) <= not (a xor b);
    outputs(8296) <= not b or a;
    outputs(8297) <= not b;
    outputs(8298) <= not (a xor b);
    outputs(8299) <= a and b;
    outputs(8300) <= a and not b;
    outputs(8301) <= a and b;
    outputs(8302) <= not a or b;
    outputs(8303) <= not (a or b);
    outputs(8304) <= not b or a;
    outputs(8305) <= not (a xor b);
    outputs(8306) <= not (a or b);
    outputs(8307) <= b;
    outputs(8308) <= a xor b;
    outputs(8309) <= not (a xor b);
    outputs(8310) <= not b or a;
    outputs(8311) <= a xor b;
    outputs(8312) <= a and b;
    outputs(8313) <= not a or b;
    outputs(8314) <= a xor b;
    outputs(8315) <= a and not b;
    outputs(8316) <= not a;
    outputs(8317) <= not b or a;
    outputs(8318) <= b and not a;
    outputs(8319) <= a xor b;
    outputs(8320) <= a xor b;
    outputs(8321) <= a;
    outputs(8322) <= not (a xor b);
    outputs(8323) <= a xor b;
    outputs(8324) <= not (a xor b);
    outputs(8325) <= b;
    outputs(8326) <= a xor b;
    outputs(8327) <= a and not b;
    outputs(8328) <= not b;
    outputs(8329) <= not (a xor b);
    outputs(8330) <= a xor b;
    outputs(8331) <= b;
    outputs(8332) <= not a;
    outputs(8333) <= b;
    outputs(8334) <= not (a xor b);
    outputs(8335) <= not a;
    outputs(8336) <= b;
    outputs(8337) <= not (a xor b);
    outputs(8338) <= not a;
    outputs(8339) <= a;
    outputs(8340) <= not b;
    outputs(8341) <= not b or a;
    outputs(8342) <= a;
    outputs(8343) <= a xor b;
    outputs(8344) <= b and not a;
    outputs(8345) <= not a;
    outputs(8346) <= not b or a;
    outputs(8347) <= b;
    outputs(8348) <= b;
    outputs(8349) <= not (a xor b);
    outputs(8350) <= not b or a;
    outputs(8351) <= a xor b;
    outputs(8352) <= a and not b;
    outputs(8353) <= a xor b;
    outputs(8354) <= a xor b;
    outputs(8355) <= not (a xor b);
    outputs(8356) <= b;
    outputs(8357) <= a or b;
    outputs(8358) <= not (a or b);
    outputs(8359) <= a and not b;
    outputs(8360) <= not a;
    outputs(8361) <= not (a xor b);
    outputs(8362) <= a xor b;
    outputs(8363) <= not b;
    outputs(8364) <= not b;
    outputs(8365) <= a xor b;
    outputs(8366) <= a xor b;
    outputs(8367) <= not a;
    outputs(8368) <= not (a xor b);
    outputs(8369) <= a xor b;
    outputs(8370) <= a xor b;
    outputs(8371) <= a xor b;
    outputs(8372) <= a xor b;
    outputs(8373) <= not a;
    outputs(8374) <= a xor b;
    outputs(8375) <= a and b;
    outputs(8376) <= not (a xor b);
    outputs(8377) <= a or b;
    outputs(8378) <= a xor b;
    outputs(8379) <= a xor b;
    outputs(8380) <= not b;
    outputs(8381) <= not a;
    outputs(8382) <= b;
    outputs(8383) <= not b;
    outputs(8384) <= b;
    outputs(8385) <= not (a xor b);
    outputs(8386) <= not (a or b);
    outputs(8387) <= not (a or b);
    outputs(8388) <= a xor b;
    outputs(8389) <= a and not b;
    outputs(8390) <= not a or b;
    outputs(8391) <= not (a xor b);
    outputs(8392) <= not a;
    outputs(8393) <= a xor b;
    outputs(8394) <= b;
    outputs(8395) <= not a;
    outputs(8396) <= not a;
    outputs(8397) <= b;
    outputs(8398) <= a xor b;
    outputs(8399) <= not b;
    outputs(8400) <= not (a xor b);
    outputs(8401) <= not (a or b);
    outputs(8402) <= a xor b;
    outputs(8403) <= b;
    outputs(8404) <= a;
    outputs(8405) <= not (a xor b);
    outputs(8406) <= a and not b;
    outputs(8407) <= a;
    outputs(8408) <= a xor b;
    outputs(8409) <= not b;
    outputs(8410) <= not b;
    outputs(8411) <= not b;
    outputs(8412) <= a or b;
    outputs(8413) <= not (a xor b);
    outputs(8414) <= not b;
    outputs(8415) <= a;
    outputs(8416) <= not (a xor b);
    outputs(8417) <= b and not a;
    outputs(8418) <= a and b;
    outputs(8419) <= b;
    outputs(8420) <= a or b;
    outputs(8421) <= not (a xor b);
    outputs(8422) <= not b;
    outputs(8423) <= a;
    outputs(8424) <= not (a xor b);
    outputs(8425) <= a;
    outputs(8426) <= not b;
    outputs(8427) <= a xor b;
    outputs(8428) <= not a;
    outputs(8429) <= a and not b;
    outputs(8430) <= a and not b;
    outputs(8431) <= a xor b;
    outputs(8432) <= not (a xor b);
    outputs(8433) <= not (a xor b);
    outputs(8434) <= a xor b;
    outputs(8435) <= a xor b;
    outputs(8436) <= a or b;
    outputs(8437) <= not (a or b);
    outputs(8438) <= a and b;
    outputs(8439) <= a xor b;
    outputs(8440) <= a;
    outputs(8441) <= not (a xor b);
    outputs(8442) <= a;
    outputs(8443) <= a;
    outputs(8444) <= not a or b;
    outputs(8445) <= not a or b;
    outputs(8446) <= a xor b;
    outputs(8447) <= not b;
    outputs(8448) <= a;
    outputs(8449) <= not (a or b);
    outputs(8450) <= not (a xor b);
    outputs(8451) <= a xor b;
    outputs(8452) <= not b or a;
    outputs(8453) <= not (a and b);
    outputs(8454) <= not b or a;
    outputs(8455) <= not a;
    outputs(8456) <= not a;
    outputs(8457) <= a xor b;
    outputs(8458) <= not (a or b);
    outputs(8459) <= not b;
    outputs(8460) <= not b;
    outputs(8461) <= not (a xor b);
    outputs(8462) <= not (a and b);
    outputs(8463) <= a xor b;
    outputs(8464) <= not a;
    outputs(8465) <= a xor b;
    outputs(8466) <= not b or a;
    outputs(8467) <= b;
    outputs(8468) <= a;
    outputs(8469) <= b;
    outputs(8470) <= not (a xor b);
    outputs(8471) <= not (a xor b);
    outputs(8472) <= not (a or b);
    outputs(8473) <= b and not a;
    outputs(8474) <= a xor b;
    outputs(8475) <= a or b;
    outputs(8476) <= not (a xor b);
    outputs(8477) <= a xor b;
    outputs(8478) <= a and b;
    outputs(8479) <= not (a or b);
    outputs(8480) <= a;
    outputs(8481) <= not a or b;
    outputs(8482) <= not b or a;
    outputs(8483) <= a xor b;
    outputs(8484) <= not (a xor b);
    outputs(8485) <= a xor b;
    outputs(8486) <= b;
    outputs(8487) <= a and not b;
    outputs(8488) <= b;
    outputs(8489) <= not a;
    outputs(8490) <= not a;
    outputs(8491) <= a and not b;
    outputs(8492) <= not (a xor b);
    outputs(8493) <= not (a xor b);
    outputs(8494) <= not b;
    outputs(8495) <= not b;
    outputs(8496) <= a xor b;
    outputs(8497) <= b;
    outputs(8498) <= a;
    outputs(8499) <= b;
    outputs(8500) <= not (a or b);
    outputs(8501) <= b;
    outputs(8502) <= b;
    outputs(8503) <= b;
    outputs(8504) <= not (a or b);
    outputs(8505) <= b;
    outputs(8506) <= not (a xor b);
    outputs(8507) <= a xor b;
    outputs(8508) <= not (a xor b);
    outputs(8509) <= b;
    outputs(8510) <= a and not b;
    outputs(8511) <= a or b;
    outputs(8512) <= b;
    outputs(8513) <= a xor b;
    outputs(8514) <= not (a or b);
    outputs(8515) <= a xor b;
    outputs(8516) <= not b or a;
    outputs(8517) <= a xor b;
    outputs(8518) <= b;
    outputs(8519) <= not a;
    outputs(8520) <= a and not b;
    outputs(8521) <= not a;
    outputs(8522) <= not a;
    outputs(8523) <= b and not a;
    outputs(8524) <= not b or a;
    outputs(8525) <= not a;
    outputs(8526) <= not b;
    outputs(8527) <= a and b;
    outputs(8528) <= a and not b;
    outputs(8529) <= b;
    outputs(8530) <= not (a xor b);
    outputs(8531) <= not b;
    outputs(8532) <= a and not b;
    outputs(8533) <= b and not a;
    outputs(8534) <= a xor b;
    outputs(8535) <= a xor b;
    outputs(8536) <= b;
    outputs(8537) <= 1'b0;
    outputs(8538) <= a;
    outputs(8539) <= a;
    outputs(8540) <= not a;
    outputs(8541) <= a xor b;
    outputs(8542) <= a xor b;
    outputs(8543) <= a xor b;
    outputs(8544) <= not (a or b);
    outputs(8545) <= not (a xor b);
    outputs(8546) <= b;
    outputs(8547) <= a and not b;
    outputs(8548) <= a and not b;
    outputs(8549) <= a xor b;
    outputs(8550) <= not a;
    outputs(8551) <= b and not a;
    outputs(8552) <= not (a xor b);
    outputs(8553) <= not b or a;
    outputs(8554) <= not a;
    outputs(8555) <= not a;
    outputs(8556) <= b and not a;
    outputs(8557) <= a xor b;
    outputs(8558) <= not b;
    outputs(8559) <= b;
    outputs(8560) <= not b;
    outputs(8561) <= a xor b;
    outputs(8562) <= not (a xor b);
    outputs(8563) <= not (a xor b);
    outputs(8564) <= not b;
    outputs(8565) <= a or b;
    outputs(8566) <= b and not a;
    outputs(8567) <= a and b;
    outputs(8568) <= not a;
    outputs(8569) <= a;
    outputs(8570) <= b;
    outputs(8571) <= not (a or b);
    outputs(8572) <= a and b;
    outputs(8573) <= not (a or b);
    outputs(8574) <= a;
    outputs(8575) <= not a or b;
    outputs(8576) <= a xor b;
    outputs(8577) <= not (a xor b);
    outputs(8578) <= not b or a;
    outputs(8579) <= not a or b;
    outputs(8580) <= not a;
    outputs(8581) <= not a;
    outputs(8582) <= not a;
    outputs(8583) <= a xor b;
    outputs(8584) <= b;
    outputs(8585) <= a xor b;
    outputs(8586) <= not b or a;
    outputs(8587) <= not b;
    outputs(8588) <= b and not a;
    outputs(8589) <= not a;
    outputs(8590) <= not a;
    outputs(8591) <= not a or b;
    outputs(8592) <= a;
    outputs(8593) <= a or b;
    outputs(8594) <= not (a xor b);
    outputs(8595) <= not b;
    outputs(8596) <= a xor b;
    outputs(8597) <= not b;
    outputs(8598) <= not a or b;
    outputs(8599) <= b;
    outputs(8600) <= not (a and b);
    outputs(8601) <= not b or a;
    outputs(8602) <= not a;
    outputs(8603) <= not (a xor b);
    outputs(8604) <= b;
    outputs(8605) <= a and not b;
    outputs(8606) <= not a;
    outputs(8607) <= b;
    outputs(8608) <= a or b;
    outputs(8609) <= a;
    outputs(8610) <= not (a xor b);
    outputs(8611) <= a xor b;
    outputs(8612) <= a and not b;
    outputs(8613) <= a xor b;
    outputs(8614) <= a xor b;
    outputs(8615) <= a and b;
    outputs(8616) <= b;
    outputs(8617) <= a;
    outputs(8618) <= a xor b;
    outputs(8619) <= not b;
    outputs(8620) <= not b;
    outputs(8621) <= not (a xor b);
    outputs(8622) <= a and not b;
    outputs(8623) <= not a;
    outputs(8624) <= not a or b;
    outputs(8625) <= a xor b;
    outputs(8626) <= a or b;
    outputs(8627) <= not (a and b);
    outputs(8628) <= a;
    outputs(8629) <= b and not a;
    outputs(8630) <= a xor b;
    outputs(8631) <= not b or a;
    outputs(8632) <= not a;
    outputs(8633) <= not (a xor b);
    outputs(8634) <= a and b;
    outputs(8635) <= not (a xor b);
    outputs(8636) <= a xor b;
    outputs(8637) <= not (a and b);
    outputs(8638) <= a;
    outputs(8639) <= b;
    outputs(8640) <= a xor b;
    outputs(8641) <= b;
    outputs(8642) <= a xor b;
    outputs(8643) <= not (a or b);
    outputs(8644) <= not (a xor b);
    outputs(8645) <= a xor b;
    outputs(8646) <= not (a or b);
    outputs(8647) <= not a;
    outputs(8648) <= not a;
    outputs(8649) <= a xor b;
    outputs(8650) <= not (a or b);
    outputs(8651) <= not (a or b);
    outputs(8652) <= not b;
    outputs(8653) <= a xor b;
    outputs(8654) <= b and not a;
    outputs(8655) <= not (a xor b);
    outputs(8656) <= a and not b;
    outputs(8657) <= a or b;
    outputs(8658) <= b;
    outputs(8659) <= a xor b;
    outputs(8660) <= not b;
    outputs(8661) <= not b;
    outputs(8662) <= a xor b;
    outputs(8663) <= a xor b;
    outputs(8664) <= a and b;
    outputs(8665) <= a xor b;
    outputs(8666) <= not (a xor b);
    outputs(8667) <= a xor b;
    outputs(8668) <= not b or a;
    outputs(8669) <= not a;
    outputs(8670) <= not a;
    outputs(8671) <= a and b;
    outputs(8672) <= b and not a;
    outputs(8673) <= a and b;
    outputs(8674) <= not (a xor b);
    outputs(8675) <= a or b;
    outputs(8676) <= a and not b;
    outputs(8677) <= b;
    outputs(8678) <= a and not b;
    outputs(8679) <= b and not a;
    outputs(8680) <= a xor b;
    outputs(8681) <= a;
    outputs(8682) <= not b;
    outputs(8683) <= b;
    outputs(8684) <= a xor b;
    outputs(8685) <= not (a xor b);
    outputs(8686) <= a xor b;
    outputs(8687) <= not (a xor b);
    outputs(8688) <= b;
    outputs(8689) <= a or b;
    outputs(8690) <= not a or b;
    outputs(8691) <= not a;
    outputs(8692) <= not (a xor b);
    outputs(8693) <= b;
    outputs(8694) <= a;
    outputs(8695) <= not b;
    outputs(8696) <= not (a xor b);
    outputs(8697) <= b;
    outputs(8698) <= not (a xor b);
    outputs(8699) <= b;
    outputs(8700) <= a xor b;
    outputs(8701) <= a xor b;
    outputs(8702) <= a;
    outputs(8703) <= not b;
    outputs(8704) <= not a or b;
    outputs(8705) <= a xor b;
    outputs(8706) <= not (a or b);
    outputs(8707) <= not b;
    outputs(8708) <= b;
    outputs(8709) <= not a or b;
    outputs(8710) <= not (a or b);
    outputs(8711) <= a xor b;
    outputs(8712) <= not (a or b);
    outputs(8713) <= not b;
    outputs(8714) <= not b or a;
    outputs(8715) <= not a;
    outputs(8716) <= not b;
    outputs(8717) <= not b;
    outputs(8718) <= b;
    outputs(8719) <= not (a xor b);
    outputs(8720) <= a and b;
    outputs(8721) <= b;
    outputs(8722) <= not b;
    outputs(8723) <= a xor b;
    outputs(8724) <= not (a xor b);
    outputs(8725) <= not (a xor b);
    outputs(8726) <= not (a xor b);
    outputs(8727) <= a;
    outputs(8728) <= a or b;
    outputs(8729) <= not b or a;
    outputs(8730) <= a and b;
    outputs(8731) <= not (a or b);
    outputs(8732) <= not (a xor b);
    outputs(8733) <= b;
    outputs(8734) <= a xor b;
    outputs(8735) <= not (a xor b);
    outputs(8736) <= not (a or b);
    outputs(8737) <= b;
    outputs(8738) <= a and b;
    outputs(8739) <= not (a or b);
    outputs(8740) <= not a;
    outputs(8741) <= a;
    outputs(8742) <= not (a xor b);
    outputs(8743) <= not (a xor b);
    outputs(8744) <= not (a xor b);
    outputs(8745) <= not (a xor b);
    outputs(8746) <= a xor b;
    outputs(8747) <= not a;
    outputs(8748) <= b;
    outputs(8749) <= not b;
    outputs(8750) <= not (a or b);
    outputs(8751) <= not a;
    outputs(8752) <= not a;
    outputs(8753) <= a xor b;
    outputs(8754) <= a xor b;
    outputs(8755) <= a xor b;
    outputs(8756) <= a or b;
    outputs(8757) <= not b;
    outputs(8758) <= not (a xor b);
    outputs(8759) <= not (a xor b);
    outputs(8760) <= a or b;
    outputs(8761) <= b;
    outputs(8762) <= not a;
    outputs(8763) <= b;
    outputs(8764) <= a xor b;
    outputs(8765) <= not b;
    outputs(8766) <= b and not a;
    outputs(8767) <= b and not a;
    outputs(8768) <= a xor b;
    outputs(8769) <= b;
    outputs(8770) <= not (a xor b);
    outputs(8771) <= not (a xor b);
    outputs(8772) <= not b;
    outputs(8773) <= a xor b;
    outputs(8774) <= a;
    outputs(8775) <= a xor b;
    outputs(8776) <= not (a xor b);
    outputs(8777) <= a;
    outputs(8778) <= not a;
    outputs(8779) <= a;
    outputs(8780) <= b;
    outputs(8781) <= b and not a;
    outputs(8782) <= not b;
    outputs(8783) <= not (a xor b);
    outputs(8784) <= not b or a;
    outputs(8785) <= a xor b;
    outputs(8786) <= a;
    outputs(8787) <= not (a xor b);
    outputs(8788) <= not (a or b);
    outputs(8789) <= a xor b;
    outputs(8790) <= b and not a;
    outputs(8791) <= not b or a;
    outputs(8792) <= b and not a;
    outputs(8793) <= not a or b;
    outputs(8794) <= a and b;
    outputs(8795) <= not a or b;
    outputs(8796) <= not b;
    outputs(8797) <= not a;
    outputs(8798) <= b;
    outputs(8799) <= not (a xor b);
    outputs(8800) <= b;
    outputs(8801) <= a xor b;
    outputs(8802) <= a;
    outputs(8803) <= a;
    outputs(8804) <= a xor b;
    outputs(8805) <= b;
    outputs(8806) <= not b;
    outputs(8807) <= not a;
    outputs(8808) <= not (a xor b);
    outputs(8809) <= b;
    outputs(8810) <= b;
    outputs(8811) <= not (a or b);
    outputs(8812) <= a;
    outputs(8813) <= not (a xor b);
    outputs(8814) <= a;
    outputs(8815) <= a and not b;
    outputs(8816) <= b;
    outputs(8817) <= a and b;
    outputs(8818) <= not b;
    outputs(8819) <= not (a xor b);
    outputs(8820) <= b;
    outputs(8821) <= a;
    outputs(8822) <= not b or a;
    outputs(8823) <= b and not a;
    outputs(8824) <= not (a xor b);
    outputs(8825) <= b;
    outputs(8826) <= not (a xor b);
    outputs(8827) <= not b;
    outputs(8828) <= a;
    outputs(8829) <= not (a xor b);
    outputs(8830) <= not a;
    outputs(8831) <= a or b;
    outputs(8832) <= not (a or b);
    outputs(8833) <= not a;
    outputs(8834) <= b;
    outputs(8835) <= a xor b;
    outputs(8836) <= not b or a;
    outputs(8837) <= not (a xor b);
    outputs(8838) <= not b;
    outputs(8839) <= b;
    outputs(8840) <= a;
    outputs(8841) <= a xor b;
    outputs(8842) <= a;
    outputs(8843) <= a xor b;
    outputs(8844) <= a xor b;
    outputs(8845) <= not (a xor b);
    outputs(8846) <= not b or a;
    outputs(8847) <= not a or b;
    outputs(8848) <= b;
    outputs(8849) <= a xor b;
    outputs(8850) <= not (a xor b);
    outputs(8851) <= a xor b;
    outputs(8852) <= a xor b;
    outputs(8853) <= b;
    outputs(8854) <= a xor b;
    outputs(8855) <= b and not a;
    outputs(8856) <= a xor b;
    outputs(8857) <= not (a and b);
    outputs(8858) <= a and b;
    outputs(8859) <= a or b;
    outputs(8860) <= not a;
    outputs(8861) <= not (a and b);
    outputs(8862) <= not (a and b);
    outputs(8863) <= b;
    outputs(8864) <= b;
    outputs(8865) <= a xor b;
    outputs(8866) <= a xor b;
    outputs(8867) <= not (a xor b);
    outputs(8868) <= b;
    outputs(8869) <= not b;
    outputs(8870) <= b;
    outputs(8871) <= not b or a;
    outputs(8872) <= a xor b;
    outputs(8873) <= not a or b;
    outputs(8874) <= a xor b;
    outputs(8875) <= a xor b;
    outputs(8876) <= a;
    outputs(8877) <= a and b;
    outputs(8878) <= b;
    outputs(8879) <= not (a or b);
    outputs(8880) <= not b or a;
    outputs(8881) <= a and b;
    outputs(8882) <= not a;
    outputs(8883) <= a xor b;
    outputs(8884) <= not (a or b);
    outputs(8885) <= b;
    outputs(8886) <= a xor b;
    outputs(8887) <= not (a or b);
    outputs(8888) <= a xor b;
    outputs(8889) <= a xor b;
    outputs(8890) <= a xor b;
    outputs(8891) <= not b;
    outputs(8892) <= not a;
    outputs(8893) <= not b;
    outputs(8894) <= not a;
    outputs(8895) <= not (a and b);
    outputs(8896) <= not a or b;
    outputs(8897) <= b and not a;
    outputs(8898) <= a;
    outputs(8899) <= b;
    outputs(8900) <= b;
    outputs(8901) <= not a;
    outputs(8902) <= not (a xor b);
    outputs(8903) <= not b or a;
    outputs(8904) <= a;
    outputs(8905) <= not (a xor b);
    outputs(8906) <= not a;
    outputs(8907) <= not (a or b);
    outputs(8908) <= a xor b;
    outputs(8909) <= a or b;
    outputs(8910) <= a;
    outputs(8911) <= a and not b;
    outputs(8912) <= a;
    outputs(8913) <= not (a xor b);
    outputs(8914) <= a and not b;
    outputs(8915) <= a xor b;
    outputs(8916) <= not (a and b);
    outputs(8917) <= not b or a;
    outputs(8918) <= a xor b;
    outputs(8919) <= b and not a;
    outputs(8920) <= not a;
    outputs(8921) <= a and not b;
    outputs(8922) <= a;
    outputs(8923) <= not b;
    outputs(8924) <= a;
    outputs(8925) <= b and not a;
    outputs(8926) <= a;
    outputs(8927) <= not (a xor b);
    outputs(8928) <= not (a or b);
    outputs(8929) <= a xor b;
    outputs(8930) <= not a;
    outputs(8931) <= a xor b;
    outputs(8932) <= not a;
    outputs(8933) <= b;
    outputs(8934) <= not (a xor b);
    outputs(8935) <= not (a xor b);
    outputs(8936) <= not (a xor b);
    outputs(8937) <= a xor b;
    outputs(8938) <= a or b;
    outputs(8939) <= not (a xor b);
    outputs(8940) <= a;
    outputs(8941) <= not (a xor b);
    outputs(8942) <= a or b;
    outputs(8943) <= a xor b;
    outputs(8944) <= not b;
    outputs(8945) <= a xor b;
    outputs(8946) <= a and b;
    outputs(8947) <= not b;
    outputs(8948) <= not b;
    outputs(8949) <= b;
    outputs(8950) <= b;
    outputs(8951) <= b;
    outputs(8952) <= not (a or b);
    outputs(8953) <= a xor b;
    outputs(8954) <= b;
    outputs(8955) <= a and b;
    outputs(8956) <= a and b;
    outputs(8957) <= a xor b;
    outputs(8958) <= not b;
    outputs(8959) <= not (a xor b);
    outputs(8960) <= not a;
    outputs(8961) <= not b;
    outputs(8962) <= a;
    outputs(8963) <= not (a xor b);
    outputs(8964) <= not (a and b);
    outputs(8965) <= a xor b;
    outputs(8966) <= not a;
    outputs(8967) <= a xor b;
    outputs(8968) <= a xor b;
    outputs(8969) <= a and b;
    outputs(8970) <= b;
    outputs(8971) <= not (a or b);
    outputs(8972) <= not (a xor b);
    outputs(8973) <= not b;
    outputs(8974) <= not b;
    outputs(8975) <= not b;
    outputs(8976) <= a;
    outputs(8977) <= b and not a;
    outputs(8978) <= not b;
    outputs(8979) <= b and not a;
    outputs(8980) <= a xor b;
    outputs(8981) <= a xor b;
    outputs(8982) <= a;
    outputs(8983) <= not b;
    outputs(8984) <= a xor b;
    outputs(8985) <= not b;
    outputs(8986) <= not (a and b);
    outputs(8987) <= not a;
    outputs(8988) <= 1'b0;
    outputs(8989) <= not b;
    outputs(8990) <= a and not b;
    outputs(8991) <= not (a xor b);
    outputs(8992) <= not a or b;
    outputs(8993) <= a and b;
    outputs(8994) <= b;
    outputs(8995) <= not a;
    outputs(8996) <= a;
    outputs(8997) <= a;
    outputs(8998) <= not (a xor b);
    outputs(8999) <= not (a and b);
    outputs(9000) <= not (a xor b);
    outputs(9001) <= not (a and b);
    outputs(9002) <= a xor b;
    outputs(9003) <= a xor b;
    outputs(9004) <= a xor b;
    outputs(9005) <= not (a xor b);
    outputs(9006) <= not (a or b);
    outputs(9007) <= not (a and b);
    outputs(9008) <= not (a xor b);
    outputs(9009) <= not (a xor b);
    outputs(9010) <= a and not b;
    outputs(9011) <= not b or a;
    outputs(9012) <= not a or b;
    outputs(9013) <= not a;
    outputs(9014) <= a and not b;
    outputs(9015) <= not a;
    outputs(9016) <= a xor b;
    outputs(9017) <= not (a xor b);
    outputs(9018) <= a and not b;
    outputs(9019) <= not b;
    outputs(9020) <= b and not a;
    outputs(9021) <= b and not a;
    outputs(9022) <= b and not a;
    outputs(9023) <= a xor b;
    outputs(9024) <= b and not a;
    outputs(9025) <= not b;
    outputs(9026) <= a and not b;
    outputs(9027) <= not (a xor b);
    outputs(9028) <= not (a xor b);
    outputs(9029) <= not a;
    outputs(9030) <= a and b;
    outputs(9031) <= a and b;
    outputs(9032) <= a;
    outputs(9033) <= not b;
    outputs(9034) <= a;
    outputs(9035) <= a and not b;
    outputs(9036) <= not a;
    outputs(9037) <= a and not b;
    outputs(9038) <= a and b;
    outputs(9039) <= not a;
    outputs(9040) <= a xor b;
    outputs(9041) <= not (a or b);
    outputs(9042) <= a and not b;
    outputs(9043) <= not (a xor b);
    outputs(9044) <= a or b;
    outputs(9045) <= not a;
    outputs(9046) <= a and b;
    outputs(9047) <= not (a and b);
    outputs(9048) <= not b;
    outputs(9049) <= not (a xor b);
    outputs(9050) <= a xor b;
    outputs(9051) <= a xor b;
    outputs(9052) <= a xor b;
    outputs(9053) <= not b;
    outputs(9054) <= not a;
    outputs(9055) <= not b;
    outputs(9056) <= not a;
    outputs(9057) <= not a;
    outputs(9058) <= b;
    outputs(9059) <= not b;
    outputs(9060) <= not a;
    outputs(9061) <= not (a or b);
    outputs(9062) <= a and not b;
    outputs(9063) <= not b;
    outputs(9064) <= a;
    outputs(9065) <= not a or b;
    outputs(9066) <= b;
    outputs(9067) <= b;
    outputs(9068) <= a;
    outputs(9069) <= a xor b;
    outputs(9070) <= not (a xor b);
    outputs(9071) <= a and not b;
    outputs(9072) <= a and b;
    outputs(9073) <= b;
    outputs(9074) <= b;
    outputs(9075) <= a and not b;
    outputs(9076) <= not a;
    outputs(9077) <= a and b;
    outputs(9078) <= a and b;
    outputs(9079) <= not a;
    outputs(9080) <= a and not b;
    outputs(9081) <= not (a xor b);
    outputs(9082) <= not (a or b);
    outputs(9083) <= not (a xor b);
    outputs(9084) <= b;
    outputs(9085) <= not a;
    outputs(9086) <= not (a or b);
    outputs(9087) <= a or b;
    outputs(9088) <= not a;
    outputs(9089) <= a and not b;
    outputs(9090) <= not a or b;
    outputs(9091) <= a and not b;
    outputs(9092) <= not b;
    outputs(9093) <= not a or b;
    outputs(9094) <= not b;
    outputs(9095) <= b and not a;
    outputs(9096) <= a xor b;
    outputs(9097) <= a;
    outputs(9098) <= not (a or b);
    outputs(9099) <= not (a xor b);
    outputs(9100) <= a xor b;
    outputs(9101) <= a;
    outputs(9102) <= not (a or b);
    outputs(9103) <= not (a xor b);
    outputs(9104) <= a xor b;
    outputs(9105) <= not b or a;
    outputs(9106) <= b and not a;
    outputs(9107) <= not (a xor b);
    outputs(9108) <= not (a xor b);
    outputs(9109) <= not b;
    outputs(9110) <= not b;
    outputs(9111) <= not a;
    outputs(9112) <= b;
    outputs(9113) <= not a or b;
    outputs(9114) <= not b;
    outputs(9115) <= b and not a;
    outputs(9116) <= b and not a;
    outputs(9117) <= not (a xor b);
    outputs(9118) <= a and not b;
    outputs(9119) <= a xor b;
    outputs(9120) <= not (a xor b);
    outputs(9121) <= a and not b;
    outputs(9122) <= not a;
    outputs(9123) <= a and not b;
    outputs(9124) <= a xor b;
    outputs(9125) <= a xor b;
    outputs(9126) <= not a;
    outputs(9127) <= not a or b;
    outputs(9128) <= not b;
    outputs(9129) <= not (a xor b);
    outputs(9130) <= a;
    outputs(9131) <= not (a xor b);
    outputs(9132) <= a xor b;
    outputs(9133) <= not a;
    outputs(9134) <= not a;
    outputs(9135) <= a xor b;
    outputs(9136) <= not (a and b);
    outputs(9137) <= not (a xor b);
    outputs(9138) <= a;
    outputs(9139) <= not b;
    outputs(9140) <= not a;
    outputs(9141) <= not (a xor b);
    outputs(9142) <= not a;
    outputs(9143) <= not (a xor b);
    outputs(9144) <= not (a and b);
    outputs(9145) <= a and b;
    outputs(9146) <= a xor b;
    outputs(9147) <= not b or a;
    outputs(9148) <= a and not b;
    outputs(9149) <= b;
    outputs(9150) <= a and not b;
    outputs(9151) <= not (a xor b);
    outputs(9152) <= not b;
    outputs(9153) <= not b;
    outputs(9154) <= a xor b;
    outputs(9155) <= b and not a;
    outputs(9156) <= b;
    outputs(9157) <= not (a xor b);
    outputs(9158) <= a xor b;
    outputs(9159) <= not (a xor b);
    outputs(9160) <= a xor b;
    outputs(9161) <= a and b;
    outputs(9162) <= not (a and b);
    outputs(9163) <= a or b;
    outputs(9164) <= b and not a;
    outputs(9165) <= a and not b;
    outputs(9166) <= not (a and b);
    outputs(9167) <= not a;
    outputs(9168) <= a xor b;
    outputs(9169) <= b and not a;
    outputs(9170) <= b and not a;
    outputs(9171) <= not b or a;
    outputs(9172) <= not (a or b);
    outputs(9173) <= a and not b;
    outputs(9174) <= a and b;
    outputs(9175) <= a or b;
    outputs(9176) <= a;
    outputs(9177) <= a xor b;
    outputs(9178) <= not (a and b);
    outputs(9179) <= not b;
    outputs(9180) <= not b or a;
    outputs(9181) <= b;
    outputs(9182) <= b;
    outputs(9183) <= not (a or b);
    outputs(9184) <= b and not a;
    outputs(9185) <= not (a xor b);
    outputs(9186) <= b;
    outputs(9187) <= not a;
    outputs(9188) <= b;
    outputs(9189) <= not b;
    outputs(9190) <= not b or a;
    outputs(9191) <= not b or a;
    outputs(9192) <= a and b;
    outputs(9193) <= not (a or b);
    outputs(9194) <= not (a and b);
    outputs(9195) <= not a;
    outputs(9196) <= a xor b;
    outputs(9197) <= a;
    outputs(9198) <= a;
    outputs(9199) <= b and not a;
    outputs(9200) <= a and not b;
    outputs(9201) <= not (a or b);
    outputs(9202) <= not (a xor b);
    outputs(9203) <= not a or b;
    outputs(9204) <= a and b;
    outputs(9205) <= not (a or b);
    outputs(9206) <= a and b;
    outputs(9207) <= not (a xor b);
    outputs(9208) <= a xor b;
    outputs(9209) <= not a;
    outputs(9210) <= not (a or b);
    outputs(9211) <= a and b;
    outputs(9212) <= b and not a;
    outputs(9213) <= not (a xor b);
    outputs(9214) <= a;
    outputs(9215) <= a and b;
    outputs(9216) <= not (a xor b);
    outputs(9217) <= not (a xor b);
    outputs(9218) <= not (a or b);
    outputs(9219) <= 1'b0;
    outputs(9220) <= not (a xor b);
    outputs(9221) <= not (a xor b);
    outputs(9222) <= not (a xor b);
    outputs(9223) <= a;
    outputs(9224) <= a xor b;
    outputs(9225) <= a xor b;
    outputs(9226) <= not b;
    outputs(9227) <= a;
    outputs(9228) <= not a;
    outputs(9229) <= b;
    outputs(9230) <= a and b;
    outputs(9231) <= not (a xor b);
    outputs(9232) <= a and b;
    outputs(9233) <= a and b;
    outputs(9234) <= not b;
    outputs(9235) <= a and not b;
    outputs(9236) <= b;
    outputs(9237) <= a xor b;
    outputs(9238) <= not (a xor b);
    outputs(9239) <= not a;
    outputs(9240) <= b;
    outputs(9241) <= b;
    outputs(9242) <= not (a xor b);
    outputs(9243) <= a or b;
    outputs(9244) <= not b;
    outputs(9245) <= not (a xor b);
    outputs(9246) <= not (a or b);
    outputs(9247) <= not a;
    outputs(9248) <= not b;
    outputs(9249) <= not b;
    outputs(9250) <= not (a or b);
    outputs(9251) <= a and not b;
    outputs(9252) <= not (a xor b);
    outputs(9253) <= a xor b;
    outputs(9254) <= a and not b;
    outputs(9255) <= a and not b;
    outputs(9256) <= not b;
    outputs(9257) <= a xor b;
    outputs(9258) <= a or b;
    outputs(9259) <= a;
    outputs(9260) <= not (a xor b);
    outputs(9261) <= not b;
    outputs(9262) <= not (a and b);
    outputs(9263) <= not a;
    outputs(9264) <= a and b;
    outputs(9265) <= a and not b;
    outputs(9266) <= not a;
    outputs(9267) <= not (a or b);
    outputs(9268) <= a or b;
    outputs(9269) <= not b;
    outputs(9270) <= not a;
    outputs(9271) <= b;
    outputs(9272) <= a xor b;
    outputs(9273) <= not (a xor b);
    outputs(9274) <= b;
    outputs(9275) <= not a;
    outputs(9276) <= not a;
    outputs(9277) <= not (a xor b);
    outputs(9278) <= not a;
    outputs(9279) <= b;
    outputs(9280) <= a and not b;
    outputs(9281) <= not a;
    outputs(9282) <= not b or a;
    outputs(9283) <= a and not b;
    outputs(9284) <= not a;
    outputs(9285) <= not a;
    outputs(9286) <= not (a xor b);
    outputs(9287) <= a;
    outputs(9288) <= not (a xor b);
    outputs(9289) <= a;
    outputs(9290) <= not (a xor b);
    outputs(9291) <= a xor b;
    outputs(9292) <= not a;
    outputs(9293) <= a and b;
    outputs(9294) <= a xor b;
    outputs(9295) <= not b or a;
    outputs(9296) <= not a;
    outputs(9297) <= not (a or b);
    outputs(9298) <= a and not b;
    outputs(9299) <= a and not b;
    outputs(9300) <= not (a xor b);
    outputs(9301) <= not a or b;
    outputs(9302) <= a;
    outputs(9303) <= a and b;
    outputs(9304) <= not (a or b);
    outputs(9305) <= a and not b;
    outputs(9306) <= a and not b;
    outputs(9307) <= a xor b;
    outputs(9308) <= not a;
    outputs(9309) <= a;
    outputs(9310) <= not (a xor b);
    outputs(9311) <= not a;
    outputs(9312) <= b and not a;
    outputs(9313) <= not (a xor b);
    outputs(9314) <= not (a xor b);
    outputs(9315) <= b;
    outputs(9316) <= not a;
    outputs(9317) <= not a;
    outputs(9318) <= a xor b;
    outputs(9319) <= a;
    outputs(9320) <= not b;
    outputs(9321) <= a xor b;
    outputs(9322) <= not a;
    outputs(9323) <= not b or a;
    outputs(9324) <= not b;
    outputs(9325) <= not (a and b);
    outputs(9326) <= a xor b;
    outputs(9327) <= b;
    outputs(9328) <= not (a xor b);
    outputs(9329) <= a;
    outputs(9330) <= a and not b;
    outputs(9331) <= not (a and b);
    outputs(9332) <= not b;
    outputs(9333) <= not b;
    outputs(9334) <= b and not a;
    outputs(9335) <= b;
    outputs(9336) <= a and b;
    outputs(9337) <= not (a or b);
    outputs(9338) <= a;
    outputs(9339) <= not b;
    outputs(9340) <= not b;
    outputs(9341) <= not b;
    outputs(9342) <= a xor b;
    outputs(9343) <= not a;
    outputs(9344) <= a and not b;
    outputs(9345) <= a xor b;
    outputs(9346) <= not a;
    outputs(9347) <= a xor b;
    outputs(9348) <= not a;
    outputs(9349) <= b and not a;
    outputs(9350) <= a and b;
    outputs(9351) <= a xor b;
    outputs(9352) <= a xor b;
    outputs(9353) <= a and not b;
    outputs(9354) <= a;
    outputs(9355) <= b and not a;
    outputs(9356) <= a;
    outputs(9357) <= not (a or b);
    outputs(9358) <= not b;
    outputs(9359) <= a xor b;
    outputs(9360) <= a;
    outputs(9361) <= not a;
    outputs(9362) <= a xor b;
    outputs(9363) <= a xor b;
    outputs(9364) <= a;
    outputs(9365) <= not b or a;
    outputs(9366) <= b and not a;
    outputs(9367) <= not b;
    outputs(9368) <= not a or b;
    outputs(9369) <= not b;
    outputs(9370) <= not (a and b);
    outputs(9371) <= a xor b;
    outputs(9372) <= a xor b;
    outputs(9373) <= b;
    outputs(9374) <= not b or a;
    outputs(9375) <= b;
    outputs(9376) <= not b or a;
    outputs(9377) <= not b;
    outputs(9378) <= b;
    outputs(9379) <= b and not a;
    outputs(9380) <= not (a xor b);
    outputs(9381) <= not (a and b);
    outputs(9382) <= a;
    outputs(9383) <= b and not a;
    outputs(9384) <= b;
    outputs(9385) <= a;
    outputs(9386) <= not b;
    outputs(9387) <= a xor b;
    outputs(9388) <= not a or b;
    outputs(9389) <= not (a xor b);
    outputs(9390) <= not (a xor b);
    outputs(9391) <= a and b;
    outputs(9392) <= a;
    outputs(9393) <= not b or a;
    outputs(9394) <= b;
    outputs(9395) <= a;
    outputs(9396) <= not a;
    outputs(9397) <= b and not a;
    outputs(9398) <= a xor b;
    outputs(9399) <= a xor b;
    outputs(9400) <= b and not a;
    outputs(9401) <= not (a xor b);
    outputs(9402) <= not a;
    outputs(9403) <= not b;
    outputs(9404) <= a and not b;
    outputs(9405) <= not (a and b);
    outputs(9406) <= not a;
    outputs(9407) <= not a;
    outputs(9408) <= b;
    outputs(9409) <= a xor b;
    outputs(9410) <= b and not a;
    outputs(9411) <= a xor b;
    outputs(9412) <= a or b;
    outputs(9413) <= a and not b;
    outputs(9414) <= a and b;
    outputs(9415) <= not (a or b);
    outputs(9416) <= not (a xor b);
    outputs(9417) <= not a;
    outputs(9418) <= not b;
    outputs(9419) <= a xor b;
    outputs(9420) <= a;
    outputs(9421) <= not (a or b);
    outputs(9422) <= not b;
    outputs(9423) <= not b;
    outputs(9424) <= a xor b;
    outputs(9425) <= not a;
    outputs(9426) <= a and not b;
    outputs(9427) <= not a;
    outputs(9428) <= not b;
    outputs(9429) <= a and b;
    outputs(9430) <= a xor b;
    outputs(9431) <= not (a xor b);
    outputs(9432) <= not (a and b);
    outputs(9433) <= not (a xor b);
    outputs(9434) <= not (a xor b);
    outputs(9435) <= not a;
    outputs(9436) <= not a;
    outputs(9437) <= a;
    outputs(9438) <= a or b;
    outputs(9439) <= not (a xor b);
    outputs(9440) <= a;
    outputs(9441) <= b;
    outputs(9442) <= a xor b;
    outputs(9443) <= a and b;
    outputs(9444) <= a xor b;
    outputs(9445) <= not b;
    outputs(9446) <= b;
    outputs(9447) <= not (a xor b);
    outputs(9448) <= a;
    outputs(9449) <= a;
    outputs(9450) <= b;
    outputs(9451) <= not (a and b);
    outputs(9452) <= not (a xor b);
    outputs(9453) <= not (a or b);
    outputs(9454) <= a and not b;
    outputs(9455) <= not b or a;
    outputs(9456) <= a;
    outputs(9457) <= b;
    outputs(9458) <= not (a xor b);
    outputs(9459) <= a xor b;
    outputs(9460) <= b and not a;
    outputs(9461) <= a;
    outputs(9462) <= b and not a;
    outputs(9463) <= b and not a;
    outputs(9464) <= not a;
    outputs(9465) <= not (a xor b);
    outputs(9466) <= a xor b;
    outputs(9467) <= not b or a;
    outputs(9468) <= not a;
    outputs(9469) <= a;
    outputs(9470) <= not (a xor b);
    outputs(9471) <= a xor b;
    outputs(9472) <= not (a and b);
    outputs(9473) <= not b;
    outputs(9474) <= not (a xor b);
    outputs(9475) <= a xor b;
    outputs(9476) <= not b or a;
    outputs(9477) <= a and not b;
    outputs(9478) <= a or b;
    outputs(9479) <= b;
    outputs(9480) <= not a;
    outputs(9481) <= b;
    outputs(9482) <= not (a or b);
    outputs(9483) <= a xor b;
    outputs(9484) <= b;
    outputs(9485) <= b;
    outputs(9486) <= not a;
    outputs(9487) <= not (a or b);
    outputs(9488) <= not (a or b);
    outputs(9489) <= a or b;
    outputs(9490) <= a or b;
    outputs(9491) <= not b;
    outputs(9492) <= a;
    outputs(9493) <= b and not a;
    outputs(9494) <= not b;
    outputs(9495) <= b;
    outputs(9496) <= a and not b;
    outputs(9497) <= a and not b;
    outputs(9498) <= a xor b;
    outputs(9499) <= not (a xor b);
    outputs(9500) <= a;
    outputs(9501) <= b;
    outputs(9502) <= not a;
    outputs(9503) <= not a;
    outputs(9504) <= a xor b;
    outputs(9505) <= a and b;
    outputs(9506) <= not a;
    outputs(9507) <= not a;
    outputs(9508) <= not (a or b);
    outputs(9509) <= not b or a;
    outputs(9510) <= not (a xor b);
    outputs(9511) <= b;
    outputs(9512) <= not b;
    outputs(9513) <= b and not a;
    outputs(9514) <= a and not b;
    outputs(9515) <= not (a xor b);
    outputs(9516) <= b and not a;
    outputs(9517) <= not a;
    outputs(9518) <= not (a xor b);
    outputs(9519) <= a and not b;
    outputs(9520) <= not (a xor b);
    outputs(9521) <= b and not a;
    outputs(9522) <= a and b;
    outputs(9523) <= not (a xor b);
    outputs(9524) <= not (a xor b);
    outputs(9525) <= not (a xor b);
    outputs(9526) <= a xor b;
    outputs(9527) <= b;
    outputs(9528) <= not a;
    outputs(9529) <= a xor b;
    outputs(9530) <= a;
    outputs(9531) <= not b or a;
    outputs(9532) <= b and not a;
    outputs(9533) <= not a;
    outputs(9534) <= not (a xor b);
    outputs(9535) <= not a;
    outputs(9536) <= b;
    outputs(9537) <= not (a or b);
    outputs(9538) <= a;
    outputs(9539) <= a xor b;
    outputs(9540) <= not a;
    outputs(9541) <= a and b;
    outputs(9542) <= not (a or b);
    outputs(9543) <= a and b;
    outputs(9544) <= b and not a;
    outputs(9545) <= a;
    outputs(9546) <= a;
    outputs(9547) <= not (a and b);
    outputs(9548) <= a and not b;
    outputs(9549) <= not a;
    outputs(9550) <= a;
    outputs(9551) <= not a;
    outputs(9552) <= a and not b;
    outputs(9553) <= a xor b;
    outputs(9554) <= a xor b;
    outputs(9555) <= a xor b;
    outputs(9556) <= not b;
    outputs(9557) <= a and not b;
    outputs(9558) <= not (a xor b);
    outputs(9559) <= a;
    outputs(9560) <= not (a and b);
    outputs(9561) <= a and b;
    outputs(9562) <= b;
    outputs(9563) <= not (a xor b);
    outputs(9564) <= not a;
    outputs(9565) <= a and not b;
    outputs(9566) <= b and not a;
    outputs(9567) <= b;
    outputs(9568) <= b and not a;
    outputs(9569) <= not (a xor b);
    outputs(9570) <= not a;
    outputs(9571) <= not a;
    outputs(9572) <= not b;
    outputs(9573) <= not a;
    outputs(9574) <= not (a xor b);
    outputs(9575) <= not (a or b);
    outputs(9576) <= b and not a;
    outputs(9577) <= b and not a;
    outputs(9578) <= not a;
    outputs(9579) <= a xor b;
    outputs(9580) <= a xor b;
    outputs(9581) <= not a or b;
    outputs(9582) <= b;
    outputs(9583) <= not (a xor b);
    outputs(9584) <= b and not a;
    outputs(9585) <= b;
    outputs(9586) <= a xor b;
    outputs(9587) <= a;
    outputs(9588) <= not b;
    outputs(9589) <= not (a xor b);
    outputs(9590) <= b and not a;
    outputs(9591) <= not (a xor b);
    outputs(9592) <= not (a xor b);
    outputs(9593) <= a;
    outputs(9594) <= a;
    outputs(9595) <= not a;
    outputs(9596) <= a xor b;
    outputs(9597) <= b and not a;
    outputs(9598) <= a and not b;
    outputs(9599) <= b;
    outputs(9600) <= b;
    outputs(9601) <= not (a or b);
    outputs(9602) <= not a;
    outputs(9603) <= not (a xor b);
    outputs(9604) <= a xor b;
    outputs(9605) <= not a or b;
    outputs(9606) <= not b or a;
    outputs(9607) <= not (a xor b);
    outputs(9608) <= a and b;
    outputs(9609) <= not (a or b);
    outputs(9610) <= not (a xor b);
    outputs(9611) <= not a or b;
    outputs(9612) <= not (a xor b);
    outputs(9613) <= b and not a;
    outputs(9614) <= not b or a;
    outputs(9615) <= not b;
    outputs(9616) <= not a or b;
    outputs(9617) <= a xor b;
    outputs(9618) <= not (a xor b);
    outputs(9619) <= not a;
    outputs(9620) <= not (a and b);
    outputs(9621) <= not (a xor b);
    outputs(9622) <= a xor b;
    outputs(9623) <= not (a or b);
    outputs(9624) <= not (a or b);
    outputs(9625) <= not (a or b);
    outputs(9626) <= not b;
    outputs(9627) <= a;
    outputs(9628) <= not b;
    outputs(9629) <= not (a xor b);
    outputs(9630) <= not b or a;
    outputs(9631) <= a xor b;
    outputs(9632) <= a and not b;
    outputs(9633) <= a and b;
    outputs(9634) <= not (a or b);
    outputs(9635) <= not (a or b);
    outputs(9636) <= a and b;
    outputs(9637) <= not b;
    outputs(9638) <= not a;
    outputs(9639) <= not a;
    outputs(9640) <= b and not a;
    outputs(9641) <= b;
    outputs(9642) <= b;
    outputs(9643) <= b;
    outputs(9644) <= a xor b;
    outputs(9645) <= a xor b;
    outputs(9646) <= not b or a;
    outputs(9647) <= not (a xor b);
    outputs(9648) <= b and not a;
    outputs(9649) <= b;
    outputs(9650) <= not a;
    outputs(9651) <= not a or b;
    outputs(9652) <= a xor b;
    outputs(9653) <= a and not b;
    outputs(9654) <= not (a xor b);
    outputs(9655) <= not (a xor b);
    outputs(9656) <= not b;
    outputs(9657) <= not b;
    outputs(9658) <= not (a xor b);
    outputs(9659) <= not b;
    outputs(9660) <= a;
    outputs(9661) <= not (a xor b);
    outputs(9662) <= b and not a;
    outputs(9663) <= a xor b;
    outputs(9664) <= not (a xor b);
    outputs(9665) <= not (a or b);
    outputs(9666) <= b and not a;
    outputs(9667) <= not a;
    outputs(9668) <= b;
    outputs(9669) <= a xor b;
    outputs(9670) <= not (a or b);
    outputs(9671) <= not (a or b);
    outputs(9672) <= a and b;
    outputs(9673) <= b;
    outputs(9674) <= not (a xor b);
    outputs(9675) <= a xor b;
    outputs(9676) <= b and not a;
    outputs(9677) <= not (a xor b);
    outputs(9678) <= a xor b;
    outputs(9679) <= not a or b;
    outputs(9680) <= not (a xor b);
    outputs(9681) <= a xor b;
    outputs(9682) <= a and not b;
    outputs(9683) <= a and b;
    outputs(9684) <= not (a xor b);
    outputs(9685) <= not a or b;
    outputs(9686) <= a xor b;
    outputs(9687) <= not (a or b);
    outputs(9688) <= a xor b;
    outputs(9689) <= a;
    outputs(9690) <= not (a xor b);
    outputs(9691) <= a;
    outputs(9692) <= not (a and b);
    outputs(9693) <= a and not b;
    outputs(9694) <= not (a xor b);
    outputs(9695) <= a and not b;
    outputs(9696) <= b;
    outputs(9697) <= not (a or b);
    outputs(9698) <= a;
    outputs(9699) <= b;
    outputs(9700) <= not (a or b);
    outputs(9701) <= a xor b;
    outputs(9702) <= a and not b;
    outputs(9703) <= not b;
    outputs(9704) <= a;
    outputs(9705) <= not a;
    outputs(9706) <= not b;
    outputs(9707) <= not b;
    outputs(9708) <= not (a xor b);
    outputs(9709) <= a and not b;
    outputs(9710) <= a or b;
    outputs(9711) <= a and b;
    outputs(9712) <= not (a or b);
    outputs(9713) <= not (a xor b);
    outputs(9714) <= not b;
    outputs(9715) <= a xor b;
    outputs(9716) <= a xor b;
    outputs(9717) <= not (a or b);
    outputs(9718) <= not (a xor b);
    outputs(9719) <= b;
    outputs(9720) <= b;
    outputs(9721) <= b;
    outputs(9722) <= a and not b;
    outputs(9723) <= a xor b;
    outputs(9724) <= a and b;
    outputs(9725) <= b;
    outputs(9726) <= a xor b;
    outputs(9727) <= b and not a;
    outputs(9728) <= not (a and b);
    outputs(9729) <= a xor b;
    outputs(9730) <= a and b;
    outputs(9731) <= not b;
    outputs(9732) <= not b;
    outputs(9733) <= a and not b;
    outputs(9734) <= a and b;
    outputs(9735) <= not a;
    outputs(9736) <= a and not b;
    outputs(9737) <= a and not b;
    outputs(9738) <= not (a or b);
    outputs(9739) <= not (a xor b);
    outputs(9740) <= not (a or b);
    outputs(9741) <= a and b;
    outputs(9742) <= b;
    outputs(9743) <= a;
    outputs(9744) <= b;
    outputs(9745) <= a and not b;
    outputs(9746) <= not a or b;
    outputs(9747) <= not b;
    outputs(9748) <= b and not a;
    outputs(9749) <= a xor b;
    outputs(9750) <= not (a xor b);
    outputs(9751) <= a;
    outputs(9752) <= a xor b;
    outputs(9753) <= b;
    outputs(9754) <= a xor b;
    outputs(9755) <= a xor b;
    outputs(9756) <= not a;
    outputs(9757) <= a and b;
    outputs(9758) <= not a;
    outputs(9759) <= not b;
    outputs(9760) <= a xor b;
    outputs(9761) <= not (a or b);
    outputs(9762) <= not a;
    outputs(9763) <= not (a xor b);
    outputs(9764) <= b;
    outputs(9765) <= a and not b;
    outputs(9766) <= not b;
    outputs(9767) <= not b or a;
    outputs(9768) <= not (a or b);
    outputs(9769) <= a or b;
    outputs(9770) <= a xor b;
    outputs(9771) <= not a;
    outputs(9772) <= not a;
    outputs(9773) <= not (a or b);
    outputs(9774) <= a xor b;
    outputs(9775) <= b;
    outputs(9776) <= not a;
    outputs(9777) <= not b;
    outputs(9778) <= not b;
    outputs(9779) <= a and b;
    outputs(9780) <= not b;
    outputs(9781) <= not b;
    outputs(9782) <= b;
    outputs(9783) <= a xor b;
    outputs(9784) <= b and not a;
    outputs(9785) <= not b;
    outputs(9786) <= b and not a;
    outputs(9787) <= not b or a;
    outputs(9788) <= b;
    outputs(9789) <= a and b;
    outputs(9790) <= not (a xor b);
    outputs(9791) <= a and not b;
    outputs(9792) <= not (a xor b);
    outputs(9793) <= b;
    outputs(9794) <= a xor b;
    outputs(9795) <= a;
    outputs(9796) <= a;
    outputs(9797) <= a and b;
    outputs(9798) <= not (a xor b);
    outputs(9799) <= not a;
    outputs(9800) <= a xor b;
    outputs(9801) <= a and b;
    outputs(9802) <= a and not b;
    outputs(9803) <= not a;
    outputs(9804) <= not b;
    outputs(9805) <= not b;
    outputs(9806) <= a and b;
    outputs(9807) <= a and not b;
    outputs(9808) <= b and not a;
    outputs(9809) <= not (a xor b);
    outputs(9810) <= a;
    outputs(9811) <= not b;
    outputs(9812) <= not b;
    outputs(9813) <= not (a xor b);
    outputs(9814) <= not b;
    outputs(9815) <= b;
    outputs(9816) <= not (a or b);
    outputs(9817) <= b and not a;
    outputs(9818) <= not (a or b);
    outputs(9819) <= a;
    outputs(9820) <= a xor b;
    outputs(9821) <= a and not b;
    outputs(9822) <= b;
    outputs(9823) <= not b;
    outputs(9824) <= not b or a;
    outputs(9825) <= not b or a;
    outputs(9826) <= a xor b;
    outputs(9827) <= not a;
    outputs(9828) <= b;
    outputs(9829) <= a;
    outputs(9830) <= a;
    outputs(9831) <= not a;
    outputs(9832) <= a xor b;
    outputs(9833) <= not b;
    outputs(9834) <= a;
    outputs(9835) <= a and not b;
    outputs(9836) <= not (a xor b);
    outputs(9837) <= not a;
    outputs(9838) <= a and not b;
    outputs(9839) <= a and b;
    outputs(9840) <= a xor b;
    outputs(9841) <= a and not b;
    outputs(9842) <= not a;
    outputs(9843) <= not (a xor b);
    outputs(9844) <= not (a xor b);
    outputs(9845) <= not (a xor b);
    outputs(9846) <= not (a xor b);
    outputs(9847) <= b;
    outputs(9848) <= b;
    outputs(9849) <= a and not b;
    outputs(9850) <= a xor b;
    outputs(9851) <= a and b;
    outputs(9852) <= b;
    outputs(9853) <= b;
    outputs(9854) <= a and not b;
    outputs(9855) <= not b;
    outputs(9856) <= not a or b;
    outputs(9857) <= not b;
    outputs(9858) <= b and not a;
    outputs(9859) <= a and not b;
    outputs(9860) <= b;
    outputs(9861) <= a and b;
    outputs(9862) <= not a;
    outputs(9863) <= a;
    outputs(9864) <= a and b;
    outputs(9865) <= b and not a;
    outputs(9866) <= a;
    outputs(9867) <= a and not b;
    outputs(9868) <= a and not b;
    outputs(9869) <= a xor b;
    outputs(9870) <= a xor b;
    outputs(9871) <= b;
    outputs(9872) <= b and not a;
    outputs(9873) <= a xor b;
    outputs(9874) <= a xor b;
    outputs(9875) <= a xor b;
    outputs(9876) <= a xor b;
    outputs(9877) <= not (a or b);
    outputs(9878) <= b;
    outputs(9879) <= not (a xor b);
    outputs(9880) <= not (a xor b);
    outputs(9881) <= a and b;
    outputs(9882) <= a xor b;
    outputs(9883) <= b;
    outputs(9884) <= not a;
    outputs(9885) <= a;
    outputs(9886) <= not b or a;
    outputs(9887) <= a or b;
    outputs(9888) <= a and not b;
    outputs(9889) <= not a;
    outputs(9890) <= a and not b;
    outputs(9891) <= b and not a;
    outputs(9892) <= not b;
    outputs(9893) <= a or b;
    outputs(9894) <= a xor b;
    outputs(9895) <= a xor b;
    outputs(9896) <= not (a xor b);
    outputs(9897) <= not (a or b);
    outputs(9898) <= not (a xor b);
    outputs(9899) <= a and not b;
    outputs(9900) <= not a;
    outputs(9901) <= not a;
    outputs(9902) <= a xor b;
    outputs(9903) <= not (a or b);
    outputs(9904) <= not a;
    outputs(9905) <= not b;
    outputs(9906) <= not (a xor b);
    outputs(9907) <= b and not a;
    outputs(9908) <= not a;
    outputs(9909) <= not (a xor b);
    outputs(9910) <= a and not b;
    outputs(9911) <= b;
    outputs(9912) <= b;
    outputs(9913) <= a xor b;
    outputs(9914) <= not b;
    outputs(9915) <= not (a xor b);
    outputs(9916) <= not b;
    outputs(9917) <= not (a or b);
    outputs(9918) <= not a;
    outputs(9919) <= a;
    outputs(9920) <= a xor b;
    outputs(9921) <= a xor b;
    outputs(9922) <= not a or b;
    outputs(9923) <= a xor b;
    outputs(9924) <= not (a and b);
    outputs(9925) <= b and not a;
    outputs(9926) <= a xor b;
    outputs(9927) <= a and b;
    outputs(9928) <= a and b;
    outputs(9929) <= a and b;
    outputs(9930) <= not (a xor b);
    outputs(9931) <= not (a xor b);
    outputs(9932) <= a xor b;
    outputs(9933) <= not (a xor b);
    outputs(9934) <= a;
    outputs(9935) <= not (a or b);
    outputs(9936) <= b;
    outputs(9937) <= a xor b;
    outputs(9938) <= not (a xor b);
    outputs(9939) <= a;
    outputs(9940) <= not b;
    outputs(9941) <= a and not b;
    outputs(9942) <= b and not a;
    outputs(9943) <= b and not a;
    outputs(9944) <= 1'b0;
    outputs(9945) <= not (a xor b);
    outputs(9946) <= not (a or b);
    outputs(9947) <= not b or a;
    outputs(9948) <= a xor b;
    outputs(9949) <= not (a xor b);
    outputs(9950) <= a xor b;
    outputs(9951) <= b and not a;
    outputs(9952) <= not b;
    outputs(9953) <= not (a xor b);
    outputs(9954) <= not (a or b);
    outputs(9955) <= not (a xor b);
    outputs(9956) <= a or b;
    outputs(9957) <= not b;
    outputs(9958) <= a xor b;
    outputs(9959) <= a xor b;
    outputs(9960) <= not (a and b);
    outputs(9961) <= not (a xor b);
    outputs(9962) <= not a;
    outputs(9963) <= a or b;
    outputs(9964) <= a xor b;
    outputs(9965) <= not a;
    outputs(9966) <= a;
    outputs(9967) <= a xor b;
    outputs(9968) <= a and b;
    outputs(9969) <= not b;
    outputs(9970) <= b;
    outputs(9971) <= a;
    outputs(9972) <= b and not a;
    outputs(9973) <= not a;
    outputs(9974) <= a and b;
    outputs(9975) <= a and b;
    outputs(9976) <= b;
    outputs(9977) <= not a;
    outputs(9978) <= a and not b;
    outputs(9979) <= not (a and b);
    outputs(9980) <= a and not b;
    outputs(9981) <= not (a or b);
    outputs(9982) <= not b;
    outputs(9983) <= a and b;
    outputs(9984) <= not (a xor b);
    outputs(9985) <= b;
    outputs(9986) <= a;
    outputs(9987) <= not b or a;
    outputs(9988) <= a xor b;
    outputs(9989) <= a and not b;
    outputs(9990) <= a and not b;
    outputs(9991) <= a and not b;
    outputs(9992) <= not (a xor b);
    outputs(9993) <= a and b;
    outputs(9994) <= a and not b;
    outputs(9995) <= not (a and b);
    outputs(9996) <= b and not a;
    outputs(9997) <= a and b;
    outputs(9998) <= a xor b;
    outputs(9999) <= not a;
    outputs(10000) <= a xor b;
    outputs(10001) <= not (a xor b);
    outputs(10002) <= a xor b;
    outputs(10003) <= not (a xor b);
    outputs(10004) <= a xor b;
    outputs(10005) <= a or b;
    outputs(10006) <= not (a xor b);
    outputs(10007) <= not a;
    outputs(10008) <= not (a xor b);
    outputs(10009) <= b and not a;
    outputs(10010) <= not (a xor b);
    outputs(10011) <= a;
    outputs(10012) <= a;
    outputs(10013) <= b;
    outputs(10014) <= a and not b;
    outputs(10015) <= not (a xor b);
    outputs(10016) <= not (a and b);
    outputs(10017) <= b;
    outputs(10018) <= b;
    outputs(10019) <= a or b;
    outputs(10020) <= not b;
    outputs(10021) <= a and b;
    outputs(10022) <= a;
    outputs(10023) <= not a;
    outputs(10024) <= b;
    outputs(10025) <= b and not a;
    outputs(10026) <= not (a xor b);
    outputs(10027) <= not (a xor b);
    outputs(10028) <= a;
    outputs(10029) <= b;
    outputs(10030) <= a xor b;
    outputs(10031) <= not a;
    outputs(10032) <= not b or a;
    outputs(10033) <= not b or a;
    outputs(10034) <= not b;
    outputs(10035) <= a xor b;
    outputs(10036) <= not (a xor b);
    outputs(10037) <= a or b;
    outputs(10038) <= b and not a;
    outputs(10039) <= a xor b;
    outputs(10040) <= a;
    outputs(10041) <= a xor b;
    outputs(10042) <= not a;
    outputs(10043) <= not b;
    outputs(10044) <= not b;
    outputs(10045) <= not (a or b);
    outputs(10046) <= not b;
    outputs(10047) <= not (a xor b);
    outputs(10048) <= b and not a;
    outputs(10049) <= b;
    outputs(10050) <= not (a or b);
    outputs(10051) <= not (a or b);
    outputs(10052) <= not b;
    outputs(10053) <= not b;
    outputs(10054) <= not b;
    outputs(10055) <= a and not b;
    outputs(10056) <= a;
    outputs(10057) <= not (a xor b);
    outputs(10058) <= not (a xor b);
    outputs(10059) <= not b;
    outputs(10060) <= a;
    outputs(10061) <= a xor b;
    outputs(10062) <= a and b;
    outputs(10063) <= not a;
    outputs(10064) <= a xor b;
    outputs(10065) <= not a;
    outputs(10066) <= b;
    outputs(10067) <= b;
    outputs(10068) <= not a or b;
    outputs(10069) <= not b;
    outputs(10070) <= not (a xor b);
    outputs(10071) <= not a or b;
    outputs(10072) <= b;
    outputs(10073) <= a xor b;
    outputs(10074) <= not b;
    outputs(10075) <= not (a xor b);
    outputs(10076) <= 1'b0;
    outputs(10077) <= not a;
    outputs(10078) <= a xor b;
    outputs(10079) <= not (a xor b);
    outputs(10080) <= not a;
    outputs(10081) <= a and not b;
    outputs(10082) <= not b;
    outputs(10083) <= a;
    outputs(10084) <= b;
    outputs(10085) <= not a;
    outputs(10086) <= not (a and b);
    outputs(10087) <= a and b;
    outputs(10088) <= a xor b;
    outputs(10089) <= a and not b;
    outputs(10090) <= not a;
    outputs(10091) <= a;
    outputs(10092) <= not b;
    outputs(10093) <= b;
    outputs(10094) <= a xor b;
    outputs(10095) <= a xor b;
    outputs(10096) <= not (a xor b);
    outputs(10097) <= a xor b;
    outputs(10098) <= b and not a;
    outputs(10099) <= a xor b;
    outputs(10100) <= a and not b;
    outputs(10101) <= not b;
    outputs(10102) <= a;
    outputs(10103) <= not a;
    outputs(10104) <= a;
    outputs(10105) <= not a;
    outputs(10106) <= not (a or b);
    outputs(10107) <= not (a xor b);
    outputs(10108) <= b and not a;
    outputs(10109) <= not a;
    outputs(10110) <= not b;
    outputs(10111) <= a and b;
    outputs(10112) <= not b or a;
    outputs(10113) <= not (a xor b);
    outputs(10114) <= not (a xor b);
    outputs(10115) <= a;
    outputs(10116) <= b;
    outputs(10117) <= not a;
    outputs(10118) <= a;
    outputs(10119) <= a xor b;
    outputs(10120) <= a xor b;
    outputs(10121) <= a and not b;
    outputs(10122) <= not (a xor b);
    outputs(10123) <= not (a and b);
    outputs(10124) <= not (a and b);
    outputs(10125) <= b and not a;
    outputs(10126) <= not b or a;
    outputs(10127) <= a and b;
    outputs(10128) <= not (a xor b);
    outputs(10129) <= not b;
    outputs(10130) <= a xor b;
    outputs(10131) <= not (a and b);
    outputs(10132) <= b and not a;
    outputs(10133) <= not b;
    outputs(10134) <= not (a or b);
    outputs(10135) <= b and not a;
    outputs(10136) <= a and not b;
    outputs(10137) <= b and not a;
    outputs(10138) <= not (a or b);
    outputs(10139) <= b;
    outputs(10140) <= a;
    outputs(10141) <= b;
    outputs(10142) <= a and b;
    outputs(10143) <= not (a and b);
    outputs(10144) <= a and b;
    outputs(10145) <= not (a xor b);
    outputs(10146) <= not (a xor b);
    outputs(10147) <= a and not b;
    outputs(10148) <= not (a or b);
    outputs(10149) <= b and not a;
    outputs(10150) <= not (a xor b);
    outputs(10151) <= b;
    outputs(10152) <= a;
    outputs(10153) <= a xor b;
    outputs(10154) <= b;
    outputs(10155) <= b;
    outputs(10156) <= not b;
    outputs(10157) <= not b;
    outputs(10158) <= b and not a;
    outputs(10159) <= not (a or b);
    outputs(10160) <= a and not b;
    outputs(10161) <= b;
    outputs(10162) <= not (a xor b);
    outputs(10163) <= a;
    outputs(10164) <= a xor b;
    outputs(10165) <= a xor b;
    outputs(10166) <= not (a xor b);
    outputs(10167) <= a;
    outputs(10168) <= b and not a;
    outputs(10169) <= b and not a;
    outputs(10170) <= not b or a;
    outputs(10171) <= not b;
    outputs(10172) <= a;
    outputs(10173) <= a;
    outputs(10174) <= not (a xor b);
    outputs(10175) <= not (a xor b);
    outputs(10176) <= a and b;
    outputs(10177) <= a xor b;
    outputs(10178) <= b and not a;
    outputs(10179) <= b;
    outputs(10180) <= not (a or b);
    outputs(10181) <= not a;
    outputs(10182) <= b;
    outputs(10183) <= a;
    outputs(10184) <= not a;
    outputs(10185) <= a or b;
    outputs(10186) <= not a;
    outputs(10187) <= not a;
    outputs(10188) <= a and not b;
    outputs(10189) <= a and not b;
    outputs(10190) <= a;
    outputs(10191) <= not b;
    outputs(10192) <= not (a and b);
    outputs(10193) <= not (a and b);
    outputs(10194) <= not (a xor b);
    outputs(10195) <= a xor b;
    outputs(10196) <= not a;
    outputs(10197) <= not (a xor b);
    outputs(10198) <= not (a xor b);
    outputs(10199) <= not (a or b);
    outputs(10200) <= a and not b;
    outputs(10201) <= not (a xor b);
    outputs(10202) <= a and b;
    outputs(10203) <= not b;
    outputs(10204) <= b;
    outputs(10205) <= a xor b;
    outputs(10206) <= a;
    outputs(10207) <= not b;
    outputs(10208) <= not (a xor b);
    outputs(10209) <= not b;
    outputs(10210) <= not (a xor b);
    outputs(10211) <= a and not b;
    outputs(10212) <= b and not a;
    outputs(10213) <= a xor b;
    outputs(10214) <= not b;
    outputs(10215) <= not (a or b);
    outputs(10216) <= not (a or b);
    outputs(10217) <= a and b;
    outputs(10218) <= a xor b;
    outputs(10219) <= a and not b;
    outputs(10220) <= not (a or b);
    outputs(10221) <= a or b;
    outputs(10222) <= not b;
    outputs(10223) <= a;
    outputs(10224) <= not a;
    outputs(10225) <= not (a xor b);
    outputs(10226) <= not (a xor b);
    outputs(10227) <= b;
    outputs(10228) <= not (a or b);
    outputs(10229) <= b;
    outputs(10230) <= b and not a;
    outputs(10231) <= b;
    outputs(10232) <= not b;
    outputs(10233) <= a and not b;
    outputs(10234) <= not (a xor b);
    outputs(10235) <= a xor b;
    outputs(10236) <= b;
    outputs(10237) <= a xor b;
    outputs(10238) <= not a;
    outputs(10239) <= a xor b;
    outputs(10240) <= a xor b;
    outputs(10241) <= a;
    outputs(10242) <= a;
    outputs(10243) <= not b or a;
    outputs(10244) <= not b;
    outputs(10245) <= a xor b;
    outputs(10246) <= not b or a;
    outputs(10247) <= b;
    outputs(10248) <= b;
    outputs(10249) <= a xor b;
    outputs(10250) <= not (a xor b);
    outputs(10251) <= a xor b;
    outputs(10252) <= not (a or b);
    outputs(10253) <= a;
    outputs(10254) <= not (a xor b);
    outputs(10255) <= a xor b;
    outputs(10256) <= not a;
    outputs(10257) <= a or b;
    outputs(10258) <= b;
    outputs(10259) <= not (a xor b);
    outputs(10260) <= not (a xor b);
    outputs(10261) <= a xor b;
    outputs(10262) <= a;
    outputs(10263) <= b;
    outputs(10264) <= not a;
    outputs(10265) <= a xor b;
    outputs(10266) <= a xor b;
    outputs(10267) <= b;
    outputs(10268) <= a or b;
    outputs(10269) <= b;
    outputs(10270) <= not a or b;
    outputs(10271) <= a xor b;
    outputs(10272) <= not (a and b);
    outputs(10273) <= not (a xor b);
    outputs(10274) <= a xor b;
    outputs(10275) <= not b;
    outputs(10276) <= not a;
    outputs(10277) <= a xor b;
    outputs(10278) <= a xor b;
    outputs(10279) <= a and not b;
    outputs(10280) <= a;
    outputs(10281) <= not a;
    outputs(10282) <= a or b;
    outputs(10283) <= not (a and b);
    outputs(10284) <= not b;
    outputs(10285) <= a xor b;
    outputs(10286) <= not (a and b);
    outputs(10287) <= not b;
    outputs(10288) <= not a;
    outputs(10289) <= not (a xor b);
    outputs(10290) <= not (a and b);
    outputs(10291) <= b;
    outputs(10292) <= a;
    outputs(10293) <= not a;
    outputs(10294) <= not a;
    outputs(10295) <= not (a xor b);
    outputs(10296) <= not a;
    outputs(10297) <= not a;
    outputs(10298) <= a xor b;
    outputs(10299) <= not b;
    outputs(10300) <= not a;
    outputs(10301) <= b and not a;
    outputs(10302) <= not (a xor b);
    outputs(10303) <= a xor b;
    outputs(10304) <= a xor b;
    outputs(10305) <= not a;
    outputs(10306) <= not a;
    outputs(10307) <= a xor b;
    outputs(10308) <= b and not a;
    outputs(10309) <= b and not a;
    outputs(10310) <= not (a xor b);
    outputs(10311) <= not (a xor b);
    outputs(10312) <= a xor b;
    outputs(10313) <= a;
    outputs(10314) <= not (a xor b);
    outputs(10315) <= b;
    outputs(10316) <= not b;
    outputs(10317) <= not (a xor b);
    outputs(10318) <= not (a xor b);
    outputs(10319) <= b;
    outputs(10320) <= a;
    outputs(10321) <= not b;
    outputs(10322) <= b and not a;
    outputs(10323) <= not b;
    outputs(10324) <= not (a or b);
    outputs(10325) <= a and not b;
    outputs(10326) <= a or b;
    outputs(10327) <= a and b;
    outputs(10328) <= b;
    outputs(10329) <= not a;
    outputs(10330) <= not (a and b);
    outputs(10331) <= a and b;
    outputs(10332) <= a xor b;
    outputs(10333) <= not (a or b);
    outputs(10334) <= a xor b;
    outputs(10335) <= not (a xor b);
    outputs(10336) <= a and b;
    outputs(10337) <= a xor b;
    outputs(10338) <= not b;
    outputs(10339) <= a xor b;
    outputs(10340) <= not b;
    outputs(10341) <= a xor b;
    outputs(10342) <= a;
    outputs(10343) <= not b;
    outputs(10344) <= a xor b;
    outputs(10345) <= b;
    outputs(10346) <= a and not b;
    outputs(10347) <= a and not b;
    outputs(10348) <= not (a or b);
    outputs(10349) <= not (a and b);
    outputs(10350) <= 1'b1;
    outputs(10351) <= not (a xor b);
    outputs(10352) <= a xor b;
    outputs(10353) <= a xor b;
    outputs(10354) <= a or b;
    outputs(10355) <= b;
    outputs(10356) <= a or b;
    outputs(10357) <= a or b;
    outputs(10358) <= a xor b;
    outputs(10359) <= not (a xor b);
    outputs(10360) <= a xor b;
    outputs(10361) <= a and not b;
    outputs(10362) <= a xor b;
    outputs(10363) <= not a;
    outputs(10364) <= a and b;
    outputs(10365) <= not b;
    outputs(10366) <= b;
    outputs(10367) <= not (a xor b);
    outputs(10368) <= b;
    outputs(10369) <= b;
    outputs(10370) <= not (a and b);
    outputs(10371) <= a xor b;
    outputs(10372) <= a and b;
    outputs(10373) <= a xor b;
    outputs(10374) <= not (a xor b);
    outputs(10375) <= not b;
    outputs(10376) <= not (a xor b);
    outputs(10377) <= not a or b;
    outputs(10378) <= a xor b;
    outputs(10379) <= a;
    outputs(10380) <= not a or b;
    outputs(10381) <= b and not a;
    outputs(10382) <= not (a xor b);
    outputs(10383) <= a xor b;
    outputs(10384) <= not a;
    outputs(10385) <= a xor b;
    outputs(10386) <= a or b;
    outputs(10387) <= not (a xor b);
    outputs(10388) <= a xor b;
    outputs(10389) <= not (a xor b);
    outputs(10390) <= not (a and b);
    outputs(10391) <= a;
    outputs(10392) <= b;
    outputs(10393) <= a xor b;
    outputs(10394) <= a xor b;
    outputs(10395) <= a;
    outputs(10396) <= not b;
    outputs(10397) <= a or b;
    outputs(10398) <= not (a xor b);
    outputs(10399) <= not a or b;
    outputs(10400) <= not a;
    outputs(10401) <= not (a and b);
    outputs(10402) <= b;
    outputs(10403) <= a xor b;
    outputs(10404) <= a;
    outputs(10405) <= not (a xor b);
    outputs(10406) <= not (a xor b);
    outputs(10407) <= not b;
    outputs(10408) <= not (a xor b);
    outputs(10409) <= a;
    outputs(10410) <= a xor b;
    outputs(10411) <= b;
    outputs(10412) <= not a;
    outputs(10413) <= not b or a;
    outputs(10414) <= a xor b;
    outputs(10415) <= b;
    outputs(10416) <= a or b;
    outputs(10417) <= b;
    outputs(10418) <= a and not b;
    outputs(10419) <= not b or a;
    outputs(10420) <= not (a xor b);
    outputs(10421) <= a and not b;
    outputs(10422) <= not a or b;
    outputs(10423) <= a and not b;
    outputs(10424) <= not a;
    outputs(10425) <= not (a and b);
    outputs(10426) <= a or b;
    outputs(10427) <= not (a xor b);
    outputs(10428) <= not (a and b);
    outputs(10429) <= not (a xor b);
    outputs(10430) <= a;
    outputs(10431) <= a and b;
    outputs(10432) <= b;
    outputs(10433) <= a xor b;
    outputs(10434) <= 1'b1;
    outputs(10435) <= not (a and b);
    outputs(10436) <= not a;
    outputs(10437) <= a;
    outputs(10438) <= a or b;
    outputs(10439) <= b;
    outputs(10440) <= not (a xor b);
    outputs(10441) <= a xor b;
    outputs(10442) <= a xor b;
    outputs(10443) <= not (a or b);
    outputs(10444) <= not (a or b);
    outputs(10445) <= not (a xor b);
    outputs(10446) <= a;
    outputs(10447) <= a or b;
    outputs(10448) <= not (a or b);
    outputs(10449) <= not a;
    outputs(10450) <= not (a xor b);
    outputs(10451) <= not (a xor b);
    outputs(10452) <= not a;
    outputs(10453) <= a and not b;
    outputs(10454) <= a;
    outputs(10455) <= b;
    outputs(10456) <= a;
    outputs(10457) <= not a or b;
    outputs(10458) <= not (a xor b);
    outputs(10459) <= a xor b;
    outputs(10460) <= b;
    outputs(10461) <= not (a xor b);
    outputs(10462) <= a xor b;
    outputs(10463) <= a xor b;
    outputs(10464) <= not b or a;
    outputs(10465) <= b;
    outputs(10466) <= a and not b;
    outputs(10467) <= a;
    outputs(10468) <= not a;
    outputs(10469) <= not a;
    outputs(10470) <= a xor b;
    outputs(10471) <= not b or a;
    outputs(10472) <= not a or b;
    outputs(10473) <= not (a xor b);
    outputs(10474) <= not (a and b);
    outputs(10475) <= a xor b;
    outputs(10476) <= not (a xor b);
    outputs(10477) <= not (a xor b);
    outputs(10478) <= a or b;
    outputs(10479) <= b;
    outputs(10480) <= a and not b;
    outputs(10481) <= not b;
    outputs(10482) <= b and not a;
    outputs(10483) <= a xor b;
    outputs(10484) <= a and b;
    outputs(10485) <= b;
    outputs(10486) <= a xor b;
    outputs(10487) <= a xor b;
    outputs(10488) <= a or b;
    outputs(10489) <= not (a and b);
    outputs(10490) <= b;
    outputs(10491) <= a;
    outputs(10492) <= a xor b;
    outputs(10493) <= a and b;
    outputs(10494) <= b;
    outputs(10495) <= a xor b;
    outputs(10496) <= b;
    outputs(10497) <= not (a xor b);
    outputs(10498) <= not (a xor b);
    outputs(10499) <= b;
    outputs(10500) <= a xor b;
    outputs(10501) <= a xor b;
    outputs(10502) <= a and b;
    outputs(10503) <= a;
    outputs(10504) <= not a;
    outputs(10505) <= not a or b;
    outputs(10506) <= not b;
    outputs(10507) <= a or b;
    outputs(10508) <= not (a xor b);
    outputs(10509) <= not b;
    outputs(10510) <= a xor b;
    outputs(10511) <= not (a xor b);
    outputs(10512) <= b and not a;
    outputs(10513) <= not (a and b);
    outputs(10514) <= b;
    outputs(10515) <= a or b;
    outputs(10516) <= a xor b;
    outputs(10517) <= not b or a;
    outputs(10518) <= not b;
    outputs(10519) <= b and not a;
    outputs(10520) <= not b;
    outputs(10521) <= b;
    outputs(10522) <= a xor b;
    outputs(10523) <= a and b;
    outputs(10524) <= not (a xor b);
    outputs(10525) <= a;
    outputs(10526) <= not b;
    outputs(10527) <= a;
    outputs(10528) <= not b;
    outputs(10529) <= a or b;
    outputs(10530) <= not (a xor b);
    outputs(10531) <= a;
    outputs(10532) <= b and not a;
    outputs(10533) <= a;
    outputs(10534) <= b;
    outputs(10535) <= not (a xor b);
    outputs(10536) <= not (a xor b);
    outputs(10537) <= a xor b;
    outputs(10538) <= not a;
    outputs(10539) <= not a or b;
    outputs(10540) <= not a or b;
    outputs(10541) <= not a;
    outputs(10542) <= a xor b;
    outputs(10543) <= not (a xor b);
    outputs(10544) <= a;
    outputs(10545) <= not b;
    outputs(10546) <= a and not b;
    outputs(10547) <= not (a or b);
    outputs(10548) <= not (a xor b);
    outputs(10549) <= b;
    outputs(10550) <= not (a or b);
    outputs(10551) <= not (a xor b);
    outputs(10552) <= not a or b;
    outputs(10553) <= a;
    outputs(10554) <= a xor b;
    outputs(10555) <= not b;
    outputs(10556) <= a xor b;
    outputs(10557) <= b and not a;
    outputs(10558) <= not a;
    outputs(10559) <= b;
    outputs(10560) <= not b or a;
    outputs(10561) <= not a or b;
    outputs(10562) <= not a;
    outputs(10563) <= not (a xor b);
    outputs(10564) <= a xor b;
    outputs(10565) <= a;
    outputs(10566) <= a;
    outputs(10567) <= b;
    outputs(10568) <= b;
    outputs(10569) <= not b;
    outputs(10570) <= not a or b;
    outputs(10571) <= a and b;
    outputs(10572) <= not b;
    outputs(10573) <= not (a xor b);
    outputs(10574) <= a;
    outputs(10575) <= not b or a;
    outputs(10576) <= not (a xor b);
    outputs(10577) <= not (a xor b);
    outputs(10578) <= a or b;
    outputs(10579) <= a;
    outputs(10580) <= b;
    outputs(10581) <= a and b;
    outputs(10582) <= not (a or b);
    outputs(10583) <= a;
    outputs(10584) <= not a or b;
    outputs(10585) <= not b;
    outputs(10586) <= not (a and b);
    outputs(10587) <= not b;
    outputs(10588) <= not (a xor b);
    outputs(10589) <= not (a xor b);
    outputs(10590) <= not (a xor b);
    outputs(10591) <= a and b;
    outputs(10592) <= not (a xor b);
    outputs(10593) <= a and not b;
    outputs(10594) <= not (a xor b);
    outputs(10595) <= not b;
    outputs(10596) <= a xor b;
    outputs(10597) <= a;
    outputs(10598) <= not (a xor b);
    outputs(10599) <= a xor b;
    outputs(10600) <= a xor b;
    outputs(10601) <= b;
    outputs(10602) <= not (a xor b);
    outputs(10603) <= a xor b;
    outputs(10604) <= a xor b;
    outputs(10605) <= not b;
    outputs(10606) <= not (a xor b);
    outputs(10607) <= not b;
    outputs(10608) <= not b or a;
    outputs(10609) <= not b;
    outputs(10610) <= a or b;
    outputs(10611) <= a or b;
    outputs(10612) <= not b;
    outputs(10613) <= b;
    outputs(10614) <= not a or b;
    outputs(10615) <= not b;
    outputs(10616) <= b;
    outputs(10617) <= not (a xor b);
    outputs(10618) <= a xor b;
    outputs(10619) <= a xor b;
    outputs(10620) <= a;
    outputs(10621) <= not a;
    outputs(10622) <= not (a xor b);
    outputs(10623) <= b and not a;
    outputs(10624) <= a xor b;
    outputs(10625) <= b and not a;
    outputs(10626) <= a or b;
    outputs(10627) <= not b;
    outputs(10628) <= not b;
    outputs(10629) <= a xor b;
    outputs(10630) <= b and not a;
    outputs(10631) <= not b or a;
    outputs(10632) <= a and not b;
    outputs(10633) <= not (a or b);
    outputs(10634) <= not a or b;
    outputs(10635) <= b;
    outputs(10636) <= b;
    outputs(10637) <= not (a and b);
    outputs(10638) <= a xor b;
    outputs(10639) <= b and not a;
    outputs(10640) <= b and not a;
    outputs(10641) <= a xor b;
    outputs(10642) <= a xor b;
    outputs(10643) <= not (a or b);
    outputs(10644) <= a xor b;
    outputs(10645) <= b;
    outputs(10646) <= a;
    outputs(10647) <= not b;
    outputs(10648) <= not (a xor b);
    outputs(10649) <= b;
    outputs(10650) <= a xor b;
    outputs(10651) <= not (a xor b);
    outputs(10652) <= a;
    outputs(10653) <= not b;
    outputs(10654) <= not b or a;
    outputs(10655) <= b;
    outputs(10656) <= a or b;
    outputs(10657) <= not a or b;
    outputs(10658) <= a and not b;
    outputs(10659) <= b;
    outputs(10660) <= b;
    outputs(10661) <= not a or b;
    outputs(10662) <= a;
    outputs(10663) <= not (a xor b);
    outputs(10664) <= b and not a;
    outputs(10665) <= b;
    outputs(10666) <= not a;
    outputs(10667) <= not (a and b);
    outputs(10668) <= not (a xor b);
    outputs(10669) <= not (a xor b);
    outputs(10670) <= a;
    outputs(10671) <= not (a and b);
    outputs(10672) <= not (a xor b);
    outputs(10673) <= not (a xor b);
    outputs(10674) <= a and b;
    outputs(10675) <= not (a xor b);
    outputs(10676) <= b and not a;
    outputs(10677) <= a;
    outputs(10678) <= not (a xor b);
    outputs(10679) <= a xor b;
    outputs(10680) <= not (a or b);
    outputs(10681) <= not (a xor b);
    outputs(10682) <= not (a and b);
    outputs(10683) <= not (a xor b);
    outputs(10684) <= b and not a;
    outputs(10685) <= not b;
    outputs(10686) <= a xor b;
    outputs(10687) <= not b;
    outputs(10688) <= b and not a;
    outputs(10689) <= not (a xor b);
    outputs(10690) <= a xor b;
    outputs(10691) <= not a or b;
    outputs(10692) <= b;
    outputs(10693) <= b;
    outputs(10694) <= a;
    outputs(10695) <= a;
    outputs(10696) <= not a;
    outputs(10697) <= not b or a;
    outputs(10698) <= not (a xor b);
    outputs(10699) <= not b;
    outputs(10700) <= not (a xor b);
    outputs(10701) <= a xor b;
    outputs(10702) <= a;
    outputs(10703) <= a xor b;
    outputs(10704) <= not (a and b);
    outputs(10705) <= not a or b;
    outputs(10706) <= a and not b;
    outputs(10707) <= b and not a;
    outputs(10708) <= not (a xor b);
    outputs(10709) <= a xor b;
    outputs(10710) <= a xor b;
    outputs(10711) <= a xor b;
    outputs(10712) <= a xor b;
    outputs(10713) <= not b;
    outputs(10714) <= b;
    outputs(10715) <= a;
    outputs(10716) <= not b or a;
    outputs(10717) <= not (a xor b);
    outputs(10718) <= 1'b1;
    outputs(10719) <= not a;
    outputs(10720) <= b;
    outputs(10721) <= a xor b;
    outputs(10722) <= a and b;
    outputs(10723) <= b;
    outputs(10724) <= not b;
    outputs(10725) <= a xor b;
    outputs(10726) <= not (a xor b);
    outputs(10727) <= not a;
    outputs(10728) <= not a;
    outputs(10729) <= b;
    outputs(10730) <= a;
    outputs(10731) <= a xor b;
    outputs(10732) <= b;
    outputs(10733) <= a or b;
    outputs(10734) <= not a or b;
    outputs(10735) <= not (a xor b);
    outputs(10736) <= not b;
    outputs(10737) <= a xor b;
    outputs(10738) <= not (a xor b);
    outputs(10739) <= b;
    outputs(10740) <= a;
    outputs(10741) <= a xor b;
    outputs(10742) <= a;
    outputs(10743) <= not (a or b);
    outputs(10744) <= not b or a;
    outputs(10745) <= a xor b;
    outputs(10746) <= not b or a;
    outputs(10747) <= not b;
    outputs(10748) <= not b;
    outputs(10749) <= not (a xor b);
    outputs(10750) <= a;
    outputs(10751) <= b;
    outputs(10752) <= a;
    outputs(10753) <= b and not a;
    outputs(10754) <= a xor b;
    outputs(10755) <= not b;
    outputs(10756) <= a xor b;
    outputs(10757) <= not a;
    outputs(10758) <= not (a xor b);
    outputs(10759) <= not b;
    outputs(10760) <= a xor b;
    outputs(10761) <= a xor b;
    outputs(10762) <= b;
    outputs(10763) <= b;
    outputs(10764) <= a xor b;
    outputs(10765) <= not (a xor b);
    outputs(10766) <= b and not a;
    outputs(10767) <= a xor b;
    outputs(10768) <= not b;
    outputs(10769) <= b and not a;
    outputs(10770) <= a;
    outputs(10771) <= b;
    outputs(10772) <= not (a and b);
    outputs(10773) <= b and not a;
    outputs(10774) <= a xor b;
    outputs(10775) <= not b;
    outputs(10776) <= not b or a;
    outputs(10777) <= a;
    outputs(10778) <= a;
    outputs(10779) <= a xor b;
    outputs(10780) <= not (a and b);
    outputs(10781) <= not (a xor b);
    outputs(10782) <= not (a xor b);
    outputs(10783) <= a and b;
    outputs(10784) <= not b;
    outputs(10785) <= a xor b;
    outputs(10786) <= not a;
    outputs(10787) <= a xor b;
    outputs(10788) <= b;
    outputs(10789) <= b and not a;
    outputs(10790) <= a xor b;
    outputs(10791) <= a and b;
    outputs(10792) <= not a;
    outputs(10793) <= a xor b;
    outputs(10794) <= not (a xor b);
    outputs(10795) <= b;
    outputs(10796) <= a xor b;
    outputs(10797) <= not b;
    outputs(10798) <= a;
    outputs(10799) <= a xor b;
    outputs(10800) <= a;
    outputs(10801) <= not (a xor b);
    outputs(10802) <= a xor b;
    outputs(10803) <= b;
    outputs(10804) <= a and not b;
    outputs(10805) <= a;
    outputs(10806) <= a;
    outputs(10807) <= a and b;
    outputs(10808) <= b;
    outputs(10809) <= a xor b;
    outputs(10810) <= not (a xor b);
    outputs(10811) <= b;
    outputs(10812) <= not a or b;
    outputs(10813) <= not (a xor b);
    outputs(10814) <= a xor b;
    outputs(10815) <= not (a xor b);
    outputs(10816) <= not (a and b);
    outputs(10817) <= b and not a;
    outputs(10818) <= not a;
    outputs(10819) <= a;
    outputs(10820) <= not (a xor b);
    outputs(10821) <= a xor b;
    outputs(10822) <= a or b;
    outputs(10823) <= b;
    outputs(10824) <= not (a xor b);
    outputs(10825) <= b;
    outputs(10826) <= not b;
    outputs(10827) <= not b;
    outputs(10828) <= a;
    outputs(10829) <= not a;
    outputs(10830) <= a and not b;
    outputs(10831) <= not (a xor b);
    outputs(10832) <= not (a xor b);
    outputs(10833) <= not b or a;
    outputs(10834) <= a;
    outputs(10835) <= not b or a;
    outputs(10836) <= not (a or b);
    outputs(10837) <= not (a xor b);
    outputs(10838) <= not b or a;
    outputs(10839) <= not (a xor b);
    outputs(10840) <= a;
    outputs(10841) <= a xor b;
    outputs(10842) <= a;
    outputs(10843) <= a xor b;
    outputs(10844) <= a xor b;
    outputs(10845) <= not (a xor b);
    outputs(10846) <= not (a xor b);
    outputs(10847) <= not (a xor b);
    outputs(10848) <= not (a and b);
    outputs(10849) <= a xor b;
    outputs(10850) <= b;
    outputs(10851) <= not a or b;
    outputs(10852) <= a and b;
    outputs(10853) <= a xor b;
    outputs(10854) <= a and b;
    outputs(10855) <= not a;
    outputs(10856) <= not a or b;
    outputs(10857) <= not b or a;
    outputs(10858) <= a or b;
    outputs(10859) <= b;
    outputs(10860) <= b;
    outputs(10861) <= not (a or b);
    outputs(10862) <= not b or a;
    outputs(10863) <= a or b;
    outputs(10864) <= not (a xor b);
    outputs(10865) <= not (a and b);
    outputs(10866) <= not (a xor b);
    outputs(10867) <= not a or b;
    outputs(10868) <= a;
    outputs(10869) <= not (a and b);
    outputs(10870) <= not (a xor b);
    outputs(10871) <= not (a xor b);
    outputs(10872) <= not a;
    outputs(10873) <= not (a xor b);
    outputs(10874) <= a xor b;
    outputs(10875) <= a xor b;
    outputs(10876) <= not (a xor b);
    outputs(10877) <= not a or b;
    outputs(10878) <= a;
    outputs(10879) <= not (a and b);
    outputs(10880) <= not b;
    outputs(10881) <= b;
    outputs(10882) <= a xor b;
    outputs(10883) <= not (a xor b);
    outputs(10884) <= not (a xor b);
    outputs(10885) <= not b or a;
    outputs(10886) <= b and not a;
    outputs(10887) <= not a or b;
    outputs(10888) <= not (a xor b);
    outputs(10889) <= not (a xor b);
    outputs(10890) <= not b or a;
    outputs(10891) <= not a;
    outputs(10892) <= a xor b;
    outputs(10893) <= not a;
    outputs(10894) <= not b or a;
    outputs(10895) <= a xor b;
    outputs(10896) <= a;
    outputs(10897) <= not b;
    outputs(10898) <= b;
    outputs(10899) <= a;
    outputs(10900) <= a xor b;
    outputs(10901) <= not b;
    outputs(10902) <= a and b;
    outputs(10903) <= b;
    outputs(10904) <= a and b;
    outputs(10905) <= not (a xor b);
    outputs(10906) <= not (a or b);
    outputs(10907) <= b;
    outputs(10908) <= not (a xor b);
    outputs(10909) <= not a;
    outputs(10910) <= not (a xor b);
    outputs(10911) <= not (a xor b);
    outputs(10912) <= not (a xor b);
    outputs(10913) <= not b;
    outputs(10914) <= a xor b;
    outputs(10915) <= a xor b;
    outputs(10916) <= a or b;
    outputs(10917) <= a xor b;
    outputs(10918) <= not (a xor b);
    outputs(10919) <= a and not b;
    outputs(10920) <= not (a xor b);
    outputs(10921) <= not a;
    outputs(10922) <= a and not b;
    outputs(10923) <= b;
    outputs(10924) <= a xor b;
    outputs(10925) <= not b;
    outputs(10926) <= a and not b;
    outputs(10927) <= a;
    outputs(10928) <= not a;
    outputs(10929) <= not a or b;
    outputs(10930) <= a xor b;
    outputs(10931) <= b;
    outputs(10932) <= not (a xor b);
    outputs(10933) <= not b;
    outputs(10934) <= not a;
    outputs(10935) <= a or b;
    outputs(10936) <= not (a and b);
    outputs(10937) <= not (a xor b);
    outputs(10938) <= a;
    outputs(10939) <= not a;
    outputs(10940) <= not (a xor b);
    outputs(10941) <= not (a xor b);
    outputs(10942) <= not a;
    outputs(10943) <= not a or b;
    outputs(10944) <= b;
    outputs(10945) <= not (a xor b);
    outputs(10946) <= a;
    outputs(10947) <= a xor b;
    outputs(10948) <= a and not b;
    outputs(10949) <= a;
    outputs(10950) <= not (a xor b);
    outputs(10951) <= not b;
    outputs(10952) <= a;
    outputs(10953) <= 1'b1;
    outputs(10954) <= not a;
    outputs(10955) <= not (a xor b);
    outputs(10956) <= not (a xor b);
    outputs(10957) <= a and b;
    outputs(10958) <= a xor b;
    outputs(10959) <= not (a xor b);
    outputs(10960) <= not a or b;
    outputs(10961) <= a xor b;
    outputs(10962) <= a xor b;
    outputs(10963) <= a xor b;
    outputs(10964) <= not a;
    outputs(10965) <= a xor b;
    outputs(10966) <= not (a or b);
    outputs(10967) <= a xor b;
    outputs(10968) <= not (a xor b);
    outputs(10969) <= not a;
    outputs(10970) <= a;
    outputs(10971) <= b;
    outputs(10972) <= not (a xor b);
    outputs(10973) <= not (a xor b);
    outputs(10974) <= b;
    outputs(10975) <= a and not b;
    outputs(10976) <= not b;
    outputs(10977) <= not (a and b);
    outputs(10978) <= not b;
    outputs(10979) <= not a or b;
    outputs(10980) <= a xor b;
    outputs(10981) <= b;
    outputs(10982) <= not b;
    outputs(10983) <= not b;
    outputs(10984) <= not a;
    outputs(10985) <= a xor b;
    outputs(10986) <= not a;
    outputs(10987) <= not a;
    outputs(10988) <= not a;
    outputs(10989) <= b;
    outputs(10990) <= not (a xor b);
    outputs(10991) <= not a or b;
    outputs(10992) <= not (a xor b);
    outputs(10993) <= not b;
    outputs(10994) <= a and not b;
    outputs(10995) <= not (a and b);
    outputs(10996) <= a xor b;
    outputs(10997) <= not (a xor b);
    outputs(10998) <= not b;
    outputs(10999) <= not a or b;
    outputs(11000) <= not (a and b);
    outputs(11001) <= a and b;
    outputs(11002) <= b;
    outputs(11003) <= not (a xor b);
    outputs(11004) <= not a or b;
    outputs(11005) <= not (a xor b);
    outputs(11006) <= a or b;
    outputs(11007) <= b and not a;
    outputs(11008) <= b and not a;
    outputs(11009) <= a xor b;
    outputs(11010) <= a;
    outputs(11011) <= b;
    outputs(11012) <= a xor b;
    outputs(11013) <= a or b;
    outputs(11014) <= not (a and b);
    outputs(11015) <= not a;
    outputs(11016) <= a xor b;
    outputs(11017) <= not (a xor b);
    outputs(11018) <= not (a or b);
    outputs(11019) <= not a;
    outputs(11020) <= not a or b;
    outputs(11021) <= a xor b;
    outputs(11022) <= a or b;
    outputs(11023) <= not (a and b);
    outputs(11024) <= not (a xor b);
    outputs(11025) <= a;
    outputs(11026) <= not (a and b);
    outputs(11027) <= not a or b;
    outputs(11028) <= a and not b;
    outputs(11029) <= a xor b;
    outputs(11030) <= a xor b;
    outputs(11031) <= not (a xor b);
    outputs(11032) <= not a;
    outputs(11033) <= not (a xor b);
    outputs(11034) <= not (a and b);
    outputs(11035) <= not (a or b);
    outputs(11036) <= not a;
    outputs(11037) <= a xor b;
    outputs(11038) <= not a or b;
    outputs(11039) <= not (a xor b);
    outputs(11040) <= a and not b;
    outputs(11041) <= not a;
    outputs(11042) <= not b or a;
    outputs(11043) <= a or b;
    outputs(11044) <= a and not b;
    outputs(11045) <= not b;
    outputs(11046) <= not (a xor b);
    outputs(11047) <= not b;
    outputs(11048) <= not b or a;
    outputs(11049) <= a;
    outputs(11050) <= a or b;
    outputs(11051) <= a or b;
    outputs(11052) <= b and not a;
    outputs(11053) <= a or b;
    outputs(11054) <= a or b;
    outputs(11055) <= a and b;
    outputs(11056) <= a;
    outputs(11057) <= not b;
    outputs(11058) <= not a;
    outputs(11059) <= not (a xor b);
    outputs(11060) <= not (a and b);
    outputs(11061) <= not (a and b);
    outputs(11062) <= not b;
    outputs(11063) <= a xor b;
    outputs(11064) <= a;
    outputs(11065) <= a xor b;
    outputs(11066) <= not b or a;
    outputs(11067) <= a or b;
    outputs(11068) <= b;
    outputs(11069) <= a;
    outputs(11070) <= not (a or b);
    outputs(11071) <= not (a and b);
    outputs(11072) <= a xor b;
    outputs(11073) <= a or b;
    outputs(11074) <= not a;
    outputs(11075) <= a;
    outputs(11076) <= not (a and b);
    outputs(11077) <= not (a xor b);
    outputs(11078) <= not a;
    outputs(11079) <= b;
    outputs(11080) <= not b;
    outputs(11081) <= a xor b;
    outputs(11082) <= not (a xor b);
    outputs(11083) <= a xor b;
    outputs(11084) <= not (a xor b);
    outputs(11085) <= a xor b;
    outputs(11086) <= a;
    outputs(11087) <= a xor b;
    outputs(11088) <= not a or b;
    outputs(11089) <= b;
    outputs(11090) <= not (a xor b);
    outputs(11091) <= a xor b;
    outputs(11092) <= a;
    outputs(11093) <= a and b;
    outputs(11094) <= a;
    outputs(11095) <= not (a xor b);
    outputs(11096) <= a and b;
    outputs(11097) <= not a or b;
    outputs(11098) <= b;
    outputs(11099) <= a or b;
    outputs(11100) <= a xor b;
    outputs(11101) <= not (a or b);
    outputs(11102) <= b;
    outputs(11103) <= b;
    outputs(11104) <= b;
    outputs(11105) <= a;
    outputs(11106) <= b;
    outputs(11107) <= not a;
    outputs(11108) <= a;
    outputs(11109) <= a xor b;
    outputs(11110) <= not a or b;
    outputs(11111) <= b and not a;
    outputs(11112) <= not a;
    outputs(11113) <= not b or a;
    outputs(11114) <= not (a and b);
    outputs(11115) <= a or b;
    outputs(11116) <= not a or b;
    outputs(11117) <= b and not a;
    outputs(11118) <= a;
    outputs(11119) <= a;
    outputs(11120) <= not b;
    outputs(11121) <= a;
    outputs(11122) <= not (a and b);
    outputs(11123) <= not b;
    outputs(11124) <= a xor b;
    outputs(11125) <= not (a xor b);
    outputs(11126) <= a;
    outputs(11127) <= not (a xor b);
    outputs(11128) <= b and not a;
    outputs(11129) <= not (a and b);
    outputs(11130) <= a xor b;
    outputs(11131) <= b;
    outputs(11132) <= a xor b;
    outputs(11133) <= not (a xor b);
    outputs(11134) <= a xor b;
    outputs(11135) <= not (a xor b);
    outputs(11136) <= not (a xor b);
    outputs(11137) <= a or b;
    outputs(11138) <= a and not b;
    outputs(11139) <= a;
    outputs(11140) <= not (a and b);
    outputs(11141) <= not a or b;
    outputs(11142) <= not a or b;
    outputs(11143) <= b and not a;
    outputs(11144) <= a xor b;
    outputs(11145) <= not a or b;
    outputs(11146) <= a or b;
    outputs(11147) <= not a;
    outputs(11148) <= a and b;
    outputs(11149) <= a or b;
    outputs(11150) <= a;
    outputs(11151) <= not a;
    outputs(11152) <= not (a xor b);
    outputs(11153) <= a or b;
    outputs(11154) <= not a;
    outputs(11155) <= not a;
    outputs(11156) <= a xor b;
    outputs(11157) <= a and not b;
    outputs(11158) <= not (a xor b);
    outputs(11159) <= not (a xor b);
    outputs(11160) <= a xor b;
    outputs(11161) <= a and not b;
    outputs(11162) <= a and not b;
    outputs(11163) <= a xor b;
    outputs(11164) <= a or b;
    outputs(11165) <= not a or b;
    outputs(11166) <= not b;
    outputs(11167) <= a and b;
    outputs(11168) <= not (a xor b);
    outputs(11169) <= a and b;
    outputs(11170) <= not (a xor b);
    outputs(11171) <= not a or b;
    outputs(11172) <= not b;
    outputs(11173) <= a;
    outputs(11174) <= b and not a;
    outputs(11175) <= a and b;
    outputs(11176) <= not a;
    outputs(11177) <= not (a xor b);
    outputs(11178) <= a or b;
    outputs(11179) <= a xor b;
    outputs(11180) <= a and not b;
    outputs(11181) <= not (a xor b);
    outputs(11182) <= not (a or b);
    outputs(11183) <= a xor b;
    outputs(11184) <= not b;
    outputs(11185) <= not (a xor b);
    outputs(11186) <= a;
    outputs(11187) <= a xor b;
    outputs(11188) <= a and b;
    outputs(11189) <= b;
    outputs(11190) <= not (a xor b);
    outputs(11191) <= not a;
    outputs(11192) <= not a or b;
    outputs(11193) <= a;
    outputs(11194) <= not a;
    outputs(11195) <= not (a xor b);
    outputs(11196) <= a xor b;
    outputs(11197) <= a and not b;
    outputs(11198) <= not a;
    outputs(11199) <= a;
    outputs(11200) <= not (a xor b);
    outputs(11201) <= not a or b;
    outputs(11202) <= a xor b;
    outputs(11203) <= a;
    outputs(11204) <= not a;
    outputs(11205) <= a xor b;
    outputs(11206) <= a xor b;
    outputs(11207) <= b;
    outputs(11208) <= b and not a;
    outputs(11209) <= a and b;
    outputs(11210) <= b and not a;
    outputs(11211) <= a and not b;
    outputs(11212) <= a or b;
    outputs(11213) <= not (a xor b);
    outputs(11214) <= a;
    outputs(11215) <= a;
    outputs(11216) <= not b;
    outputs(11217) <= a;
    outputs(11218) <= not b or a;
    outputs(11219) <= a or b;
    outputs(11220) <= b;
    outputs(11221) <= not (a xor b);
    outputs(11222) <= not b;
    outputs(11223) <= not b;
    outputs(11224) <= not (a xor b);
    outputs(11225) <= not (a and b);
    outputs(11226) <= a and not b;
    outputs(11227) <= not b;
    outputs(11228) <= a xor b;
    outputs(11229) <= a and b;
    outputs(11230) <= b;
    outputs(11231) <= not a or b;
    outputs(11232) <= not (a xor b);
    outputs(11233) <= b;
    outputs(11234) <= b;
    outputs(11235) <= not b;
    outputs(11236) <= not (a xor b);
    outputs(11237) <= not (a or b);
    outputs(11238) <= not (a xor b);
    outputs(11239) <= a and not b;
    outputs(11240) <= a xor b;
    outputs(11241) <= not a;
    outputs(11242) <= a;
    outputs(11243) <= not b;
    outputs(11244) <= not b or a;
    outputs(11245) <= not b;
    outputs(11246) <= not a;
    outputs(11247) <= not b;
    outputs(11248) <= not (a xor b);
    outputs(11249) <= a xor b;
    outputs(11250) <= not (a or b);
    outputs(11251) <= not a;
    outputs(11252) <= a and b;
    outputs(11253) <= a xor b;
    outputs(11254) <= a;
    outputs(11255) <= a or b;
    outputs(11256) <= a and b;
    outputs(11257) <= not a;
    outputs(11258) <= not (a xor b);
    outputs(11259) <= not (a xor b);
    outputs(11260) <= not (a xor b);
    outputs(11261) <= a;
    outputs(11262) <= not a;
    outputs(11263) <= a;
    outputs(11264) <= b;
    outputs(11265) <= b;
    outputs(11266) <= a xor b;
    outputs(11267) <= not (a xor b);
    outputs(11268) <= not a;
    outputs(11269) <= a xor b;
    outputs(11270) <= a or b;
    outputs(11271) <= not (a xor b);
    outputs(11272) <= not b or a;
    outputs(11273) <= not (a xor b);
    outputs(11274) <= not a;
    outputs(11275) <= a;
    outputs(11276) <= b;
    outputs(11277) <= not a;
    outputs(11278) <= not a;
    outputs(11279) <= not b or a;
    outputs(11280) <= a;
    outputs(11281) <= a xor b;
    outputs(11282) <= b;
    outputs(11283) <= a xor b;
    outputs(11284) <= not a;
    outputs(11285) <= b;
    outputs(11286) <= not (a and b);
    outputs(11287) <= a or b;
    outputs(11288) <= a and b;
    outputs(11289) <= a;
    outputs(11290) <= not (a xor b);
    outputs(11291) <= a xor b;
    outputs(11292) <= not b;
    outputs(11293) <= not (a xor b);
    outputs(11294) <= a xor b;
    outputs(11295) <= not b;
    outputs(11296) <= a and not b;
    outputs(11297) <= a xor b;
    outputs(11298) <= not (a xor b);
    outputs(11299) <= not b or a;
    outputs(11300) <= not a;
    outputs(11301) <= not (a xor b);
    outputs(11302) <= not b or a;
    outputs(11303) <= not b;
    outputs(11304) <= a xor b;
    outputs(11305) <= not (a xor b);
    outputs(11306) <= a or b;
    outputs(11307) <= a xor b;
    outputs(11308) <= b and not a;
    outputs(11309) <= not a;
    outputs(11310) <= a and b;
    outputs(11311) <= not b;
    outputs(11312) <= b;
    outputs(11313) <= not (a xor b);
    outputs(11314) <= a and not b;
    outputs(11315) <= not (a and b);
    outputs(11316) <= not b or a;
    outputs(11317) <= not (a or b);
    outputs(11318) <= not (a and b);
    outputs(11319) <= a;
    outputs(11320) <= b;
    outputs(11321) <= not (a xor b);
    outputs(11322) <= not b;
    outputs(11323) <= a xor b;
    outputs(11324) <= not b;
    outputs(11325) <= a xor b;
    outputs(11326) <= a;
    outputs(11327) <= not (a xor b);
    outputs(11328) <= not b;
    outputs(11329) <= a xor b;
    outputs(11330) <= a and not b;
    outputs(11331) <= a and not b;
    outputs(11332) <= a and b;
    outputs(11333) <= not (a and b);
    outputs(11334) <= not b;
    outputs(11335) <= a xor b;
    outputs(11336) <= b;
    outputs(11337) <= not (a and b);
    outputs(11338) <= b;
    outputs(11339) <= a and not b;
    outputs(11340) <= not a;
    outputs(11341) <= not a;
    outputs(11342) <= b and not a;
    outputs(11343) <= not (a xor b);
    outputs(11344) <= b;
    outputs(11345) <= not (a and b);
    outputs(11346) <= a;
    outputs(11347) <= a xor b;
    outputs(11348) <= not a;
    outputs(11349) <= not (a xor b);
    outputs(11350) <= not (a or b);
    outputs(11351) <= a;
    outputs(11352) <= not (a xor b);
    outputs(11353) <= a or b;
    outputs(11354) <= a xor b;
    outputs(11355) <= not (a and b);
    outputs(11356) <= not (a xor b);
    outputs(11357) <= a;
    outputs(11358) <= a xor b;
    outputs(11359) <= not a;
    outputs(11360) <= not a;
    outputs(11361) <= 1'b1;
    outputs(11362) <= not (a xor b);
    outputs(11363) <= a;
    outputs(11364) <= b and not a;
    outputs(11365) <= a;
    outputs(11366) <= not a;
    outputs(11367) <= not b;
    outputs(11368) <= not b;
    outputs(11369) <= not b;
    outputs(11370) <= not a;
    outputs(11371) <= not a or b;
    outputs(11372) <= a;
    outputs(11373) <= a xor b;
    outputs(11374) <= b and not a;
    outputs(11375) <= a xor b;
    outputs(11376) <= not a;
    outputs(11377) <= not (a or b);
    outputs(11378) <= a xor b;
    outputs(11379) <= a;
    outputs(11380) <= a and not b;
    outputs(11381) <= a xor b;
    outputs(11382) <= b;
    outputs(11383) <= not (a and b);
    outputs(11384) <= b and not a;
    outputs(11385) <= not (a xor b);
    outputs(11386) <= a xor b;
    outputs(11387) <= not (a xor b);
    outputs(11388) <= not (a xor b);
    outputs(11389) <= b;
    outputs(11390) <= a xor b;
    outputs(11391) <= a or b;
    outputs(11392) <= not b;
    outputs(11393) <= a xor b;
    outputs(11394) <= not a;
    outputs(11395) <= a;
    outputs(11396) <= not a;
    outputs(11397) <= not b;
    outputs(11398) <= not (a xor b);
    outputs(11399) <= not a;
    outputs(11400) <= a and b;
    outputs(11401) <= a;
    outputs(11402) <= a;
    outputs(11403) <= a xor b;
    outputs(11404) <= a;
    outputs(11405) <= not a or b;
    outputs(11406) <= a xor b;
    outputs(11407) <= not (a xor b);
    outputs(11408) <= not (a or b);
    outputs(11409) <= a;
    outputs(11410) <= not b or a;
    outputs(11411) <= not b;
    outputs(11412) <= not b or a;
    outputs(11413) <= b and not a;
    outputs(11414) <= not (a xor b);
    outputs(11415) <= a xor b;
    outputs(11416) <= a xor b;
    outputs(11417) <= not (a or b);
    outputs(11418) <= a xor b;
    outputs(11419) <= b and not a;
    outputs(11420) <= not (a or b);
    outputs(11421) <= a or b;
    outputs(11422) <= a;
    outputs(11423) <= not (a xor b);
    outputs(11424) <= a and b;
    outputs(11425) <= a and b;
    outputs(11426) <= a;
    outputs(11427) <= a and not b;
    outputs(11428) <= a xor b;
    outputs(11429) <= not a or b;
    outputs(11430) <= b;
    outputs(11431) <= not a or b;
    outputs(11432) <= not b;
    outputs(11433) <= a;
    outputs(11434) <= not (a xor b);
    outputs(11435) <= not (a xor b);
    outputs(11436) <= a;
    outputs(11437) <= not (a xor b);
    outputs(11438) <= not b;
    outputs(11439) <= b and not a;
    outputs(11440) <= a;
    outputs(11441) <= not (a xor b);
    outputs(11442) <= not b;
    outputs(11443) <= not (a xor b);
    outputs(11444) <= a and b;
    outputs(11445) <= a or b;
    outputs(11446) <= b and not a;
    outputs(11447) <= not b or a;
    outputs(11448) <= a and not b;
    outputs(11449) <= a;
    outputs(11450) <= not (a xor b);
    outputs(11451) <= a or b;
    outputs(11452) <= not a or b;
    outputs(11453) <= a and b;
    outputs(11454) <= not (a xor b);
    outputs(11455) <= a;
    outputs(11456) <= not (a xor b);
    outputs(11457) <= not b or a;
    outputs(11458) <= a xor b;
    outputs(11459) <= a xor b;
    outputs(11460) <= b;
    outputs(11461) <= a xor b;
    outputs(11462) <= a or b;
    outputs(11463) <= not b;
    outputs(11464) <= not b or a;
    outputs(11465) <= not (a xor b);
    outputs(11466) <= not (a xor b);
    outputs(11467) <= b;
    outputs(11468) <= a xor b;
    outputs(11469) <= not (a xor b);
    outputs(11470) <= a and not b;
    outputs(11471) <= not (a and b);
    outputs(11472) <= a xor b;
    outputs(11473) <= not a;
    outputs(11474) <= not b;
    outputs(11475) <= not (a xor b);
    outputs(11476) <= not (a xor b);
    outputs(11477) <= not (a xor b);
    outputs(11478) <= not b;
    outputs(11479) <= not a;
    outputs(11480) <= b;
    outputs(11481) <= not (a and b);
    outputs(11482) <= not b;
    outputs(11483) <= not (a xor b);
    outputs(11484) <= not b;
    outputs(11485) <= b and not a;
    outputs(11486) <= a;
    outputs(11487) <= a xor b;
    outputs(11488) <= a xor b;
    outputs(11489) <= a;
    outputs(11490) <= a;
    outputs(11491) <= not (a and b);
    outputs(11492) <= not (a xor b);
    outputs(11493) <= not (a xor b);
    outputs(11494) <= not b;
    outputs(11495) <= not b;
    outputs(11496) <= a xor b;
    outputs(11497) <= not (a xor b);
    outputs(11498) <= not (a xor b);
    outputs(11499) <= a or b;
    outputs(11500) <= b and not a;
    outputs(11501) <= b;
    outputs(11502) <= b and not a;
    outputs(11503) <= not b;
    outputs(11504) <= a xor b;
    outputs(11505) <= a xor b;
    outputs(11506) <= a xor b;
    outputs(11507) <= a xor b;
    outputs(11508) <= not a or b;
    outputs(11509) <= not b or a;
    outputs(11510) <= not b;
    outputs(11511) <= not a or b;
    outputs(11512) <= a and not b;
    outputs(11513) <= a xor b;
    outputs(11514) <= b and not a;
    outputs(11515) <= not (a xor b);
    outputs(11516) <= a or b;
    outputs(11517) <= not (a xor b);
    outputs(11518) <= not (a xor b);
    outputs(11519) <= not a or b;
    outputs(11520) <= a or b;
    outputs(11521) <= a and b;
    outputs(11522) <= a;
    outputs(11523) <= a and not b;
    outputs(11524) <= a or b;
    outputs(11525) <= not b;
    outputs(11526) <= not a;
    outputs(11527) <= a and b;
    outputs(11528) <= a;
    outputs(11529) <= not (a or b);
    outputs(11530) <= not a;
    outputs(11531) <= a or b;
    outputs(11532) <= a xor b;
    outputs(11533) <= not (a and b);
    outputs(11534) <= a or b;
    outputs(11535) <= b and not a;
    outputs(11536) <= a;
    outputs(11537) <= b and not a;
    outputs(11538) <= not a;
    outputs(11539) <= not b;
    outputs(11540) <= not a or b;
    outputs(11541) <= not b or a;
    outputs(11542) <= not b;
    outputs(11543) <= not (a or b);
    outputs(11544) <= not (a xor b);
    outputs(11545) <= a and not b;
    outputs(11546) <= b and not a;
    outputs(11547) <= not (a or b);
    outputs(11548) <= a and b;
    outputs(11549) <= a xor b;
    outputs(11550) <= not b;
    outputs(11551) <= a xor b;
    outputs(11552) <= not a;
    outputs(11553) <= b;
    outputs(11554) <= not b or a;
    outputs(11555) <= not a;
    outputs(11556) <= a and not b;
    outputs(11557) <= a xor b;
    outputs(11558) <= not a;
    outputs(11559) <= not a;
    outputs(11560) <= not (a xor b);
    outputs(11561) <= a xor b;
    outputs(11562) <= a and b;
    outputs(11563) <= not a;
    outputs(11564) <= a and not b;
    outputs(11565) <= not (a and b);
    outputs(11566) <= not a;
    outputs(11567) <= not a;
    outputs(11568) <= a;
    outputs(11569) <= a;
    outputs(11570) <= a xor b;
    outputs(11571) <= 1'b0;
    outputs(11572) <= not a or b;
    outputs(11573) <= not (a xor b);
    outputs(11574) <= not a;
    outputs(11575) <= a or b;
    outputs(11576) <= a xor b;
    outputs(11577) <= a and b;
    outputs(11578) <= b;
    outputs(11579) <= a xor b;
    outputs(11580) <= not b;
    outputs(11581) <= a;
    outputs(11582) <= not a;
    outputs(11583) <= b and not a;
    outputs(11584) <= not (a or b);
    outputs(11585) <= not b or a;
    outputs(11586) <= a and not b;
    outputs(11587) <= b;
    outputs(11588) <= a xor b;
    outputs(11589) <= a;
    outputs(11590) <= not a;
    outputs(11591) <= not (a or b);
    outputs(11592) <= a xor b;
    outputs(11593) <= a or b;
    outputs(11594) <= not a;
    outputs(11595) <= b and not a;
    outputs(11596) <= not b or a;
    outputs(11597) <= a and b;
    outputs(11598) <= not b;
    outputs(11599) <= not (a or b);
    outputs(11600) <= not b;
    outputs(11601) <= a xor b;
    outputs(11602) <= not b;
    outputs(11603) <= not (a and b);
    outputs(11604) <= a;
    outputs(11605) <= not (a xor b);
    outputs(11606) <= not a or b;
    outputs(11607) <= a xor b;
    outputs(11608) <= a;
    outputs(11609) <= b;
    outputs(11610) <= not a;
    outputs(11611) <= a and b;
    outputs(11612) <= b;
    outputs(11613) <= b;
    outputs(11614) <= a xor b;
    outputs(11615) <= a xor b;
    outputs(11616) <= not a;
    outputs(11617) <= a and b;
    outputs(11618) <= b;
    outputs(11619) <= b and not a;
    outputs(11620) <= b and not a;
    outputs(11621) <= a and not b;
    outputs(11622) <= a and not b;
    outputs(11623) <= a and b;
    outputs(11624) <= not (a and b);
    outputs(11625) <= a;
    outputs(11626) <= b;
    outputs(11627) <= a and not b;
    outputs(11628) <= a xor b;
    outputs(11629) <= a and not b;
    outputs(11630) <= a and b;
    outputs(11631) <= a and not b;
    outputs(11632) <= not (a xor b);
    outputs(11633) <= not b;
    outputs(11634) <= a xor b;
    outputs(11635) <= not b;
    outputs(11636) <= b;
    outputs(11637) <= a xor b;
    outputs(11638) <= not (a or b);
    outputs(11639) <= not b or a;
    outputs(11640) <= a xor b;
    outputs(11641) <= not b or a;
    outputs(11642) <= not (a or b);
    outputs(11643) <= a;
    outputs(11644) <= b;
    outputs(11645) <= a xor b;
    outputs(11646) <= a and b;
    outputs(11647) <= a xor b;
    outputs(11648) <= a and b;
    outputs(11649) <= a xor b;
    outputs(11650) <= a and b;
    outputs(11651) <= not a;
    outputs(11652) <= not a or b;
    outputs(11653) <= a and b;
    outputs(11654) <= not a;
    outputs(11655) <= not b or a;
    outputs(11656) <= b;
    outputs(11657) <= not b or a;
    outputs(11658) <= a xor b;
    outputs(11659) <= b and not a;
    outputs(11660) <= not a;
    outputs(11661) <= not (a xor b);
    outputs(11662) <= not b or a;
    outputs(11663) <= not (a xor b);
    outputs(11664) <= b and not a;
    outputs(11665) <= not (a xor b);
    outputs(11666) <= a and not b;
    outputs(11667) <= b;
    outputs(11668) <= a xor b;
    outputs(11669) <= not (a xor b);
    outputs(11670) <= not a;
    outputs(11671) <= not (a or b);
    outputs(11672) <= not b;
    outputs(11673) <= a and b;
    outputs(11674) <= a xor b;
    outputs(11675) <= not (a xor b);
    outputs(11676) <= a;
    outputs(11677) <= b;
    outputs(11678) <= b;
    outputs(11679) <= a xor b;
    outputs(11680) <= not (a xor b);
    outputs(11681) <= not a;
    outputs(11682) <= a xor b;
    outputs(11683) <= b and not a;
    outputs(11684) <= not b;
    outputs(11685) <= b and not a;
    outputs(11686) <= b;
    outputs(11687) <= a xor b;
    outputs(11688) <= not b or a;
    outputs(11689) <= a;
    outputs(11690) <= a or b;
    outputs(11691) <= a xor b;
    outputs(11692) <= a or b;
    outputs(11693) <= not (a or b);
    outputs(11694) <= not a;
    outputs(11695) <= a;
    outputs(11696) <= a xor b;
    outputs(11697) <= a and not b;
    outputs(11698) <= not b;
    outputs(11699) <= a and not b;
    outputs(11700) <= a;
    outputs(11701) <= not b;
    outputs(11702) <= a xor b;
    outputs(11703) <= a and not b;
    outputs(11704) <= a and b;
    outputs(11705) <= not (a xor b);
    outputs(11706) <= not (a xor b);
    outputs(11707) <= a and not b;
    outputs(11708) <= not b;
    outputs(11709) <= a xor b;
    outputs(11710) <= b;
    outputs(11711) <= b and not a;
    outputs(11712) <= a xor b;
    outputs(11713) <= not a;
    outputs(11714) <= a;
    outputs(11715) <= not (a xor b);
    outputs(11716) <= not (a xor b);
    outputs(11717) <= not (a and b);
    outputs(11718) <= not (a or b);
    outputs(11719) <= not b;
    outputs(11720) <= a and not b;
    outputs(11721) <= a xor b;
    outputs(11722) <= b and not a;
    outputs(11723) <= not (a or b);
    outputs(11724) <= not (a xor b);
    outputs(11725) <= b;
    outputs(11726) <= a xor b;
    outputs(11727) <= b;
    outputs(11728) <= a;
    outputs(11729) <= b and not a;
    outputs(11730) <= b and not a;
    outputs(11731) <= not (a or b);
    outputs(11732) <= b and not a;
    outputs(11733) <= a and not b;
    outputs(11734) <= b;
    outputs(11735) <= a and not b;
    outputs(11736) <= a or b;
    outputs(11737) <= a xor b;
    outputs(11738) <= a xor b;
    outputs(11739) <= b;
    outputs(11740) <= not a;
    outputs(11741) <= not (a or b);
    outputs(11742) <= b and not a;
    outputs(11743) <= a and b;
    outputs(11744) <= a or b;
    outputs(11745) <= not b or a;
    outputs(11746) <= not (a xor b);
    outputs(11747) <= b;
    outputs(11748) <= a;
    outputs(11749) <= b and not a;
    outputs(11750) <= not b;
    outputs(11751) <= a or b;
    outputs(11752) <= not (a xor b);
    outputs(11753) <= a;
    outputs(11754) <= b and not a;
    outputs(11755) <= b;
    outputs(11756) <= a and not b;
    outputs(11757) <= not (a or b);
    outputs(11758) <= not b;
    outputs(11759) <= b and not a;
    outputs(11760) <= a xor b;
    outputs(11761) <= not b or a;
    outputs(11762) <= a xor b;
    outputs(11763) <= not a;
    outputs(11764) <= not a;
    outputs(11765) <= b and not a;
    outputs(11766) <= not b or a;
    outputs(11767) <= a and b;
    outputs(11768) <= not (a xor b);
    outputs(11769) <= not (a xor b);
    outputs(11770) <= not b;
    outputs(11771) <= a and b;
    outputs(11772) <= not (a and b);
    outputs(11773) <= not (a xor b);
    outputs(11774) <= not a;
    outputs(11775) <= not (a and b);
    outputs(11776) <= not (a and b);
    outputs(11777) <= not (a or b);
    outputs(11778) <= not (a or b);
    outputs(11779) <= a xor b;
    outputs(11780) <= a and not b;
    outputs(11781) <= a;
    outputs(11782) <= a;
    outputs(11783) <= not b;
    outputs(11784) <= a xor b;
    outputs(11785) <= not a or b;
    outputs(11786) <= a xor b;
    outputs(11787) <= not (a xor b);
    outputs(11788) <= not (a or b);
    outputs(11789) <= not (a xor b);
    outputs(11790) <= a xor b;
    outputs(11791) <= a;
    outputs(11792) <= not (a xor b);
    outputs(11793) <= a xor b;
    outputs(11794) <= not (a xor b);
    outputs(11795) <= not b or a;
    outputs(11796) <= a xor b;
    outputs(11797) <= a;
    outputs(11798) <= a;
    outputs(11799) <= not (a xor b);
    outputs(11800) <= not a;
    outputs(11801) <= a;
    outputs(11802) <= not b;
    outputs(11803) <= a and b;
    outputs(11804) <= not (a or b);
    outputs(11805) <= not (a or b);
    outputs(11806) <= not b;
    outputs(11807) <= a and not b;
    outputs(11808) <= not b;
    outputs(11809) <= a;
    outputs(11810) <= a and not b;
    outputs(11811) <= not (a or b);
    outputs(11812) <= a xor b;
    outputs(11813) <= not (a or b);
    outputs(11814) <= not b or a;
    outputs(11815) <= not (a xor b);
    outputs(11816) <= a xor b;
    outputs(11817) <= not b;
    outputs(11818) <= a and b;
    outputs(11819) <= a xor b;
    outputs(11820) <= not (a or b);
    outputs(11821) <= not (a xor b);
    outputs(11822) <= not (a xor b);
    outputs(11823) <= a and not b;
    outputs(11824) <= a;
    outputs(11825) <= a xor b;
    outputs(11826) <= b and not a;
    outputs(11827) <= b and not a;
    outputs(11828) <= a and not b;
    outputs(11829) <= not a;
    outputs(11830) <= a xor b;
    outputs(11831) <= a and b;
    outputs(11832) <= b;
    outputs(11833) <= a and b;
    outputs(11834) <= not b;
    outputs(11835) <= b and not a;
    outputs(11836) <= b;
    outputs(11837) <= not b or a;
    outputs(11838) <= b;
    outputs(11839) <= b and not a;
    outputs(11840) <= b;
    outputs(11841) <= a;
    outputs(11842) <= not a;
    outputs(11843) <= not b;
    outputs(11844) <= a;
    outputs(11845) <= not (a xor b);
    outputs(11846) <= a xor b;
    outputs(11847) <= not b;
    outputs(11848) <= a and b;
    outputs(11849) <= not a or b;
    outputs(11850) <= not b;
    outputs(11851) <= a and b;
    outputs(11852) <= not (a xor b);
    outputs(11853) <= a xor b;
    outputs(11854) <= a and b;
    outputs(11855) <= not (a or b);
    outputs(11856) <= a or b;
    outputs(11857) <= a and b;
    outputs(11858) <= a or b;
    outputs(11859) <= not (a xor b);
    outputs(11860) <= a and b;
    outputs(11861) <= not (a xor b);
    outputs(11862) <= not (a or b);
    outputs(11863) <= a;
    outputs(11864) <= not (a and b);
    outputs(11865) <= not b;
    outputs(11866) <= not a or b;
    outputs(11867) <= not (a or b);
    outputs(11868) <= not (a xor b);
    outputs(11869) <= a xor b;
    outputs(11870) <= not (a xor b);
    outputs(11871) <= not (a xor b);
    outputs(11872) <= a and b;
    outputs(11873) <= b;
    outputs(11874) <= not a;
    outputs(11875) <= a xor b;
    outputs(11876) <= a xor b;
    outputs(11877) <= a and b;
    outputs(11878) <= not (a xor b);
    outputs(11879) <= not (a xor b);
    outputs(11880) <= b;
    outputs(11881) <= a xor b;
    outputs(11882) <= not (a xor b);
    outputs(11883) <= a xor b;
    outputs(11884) <= not b or a;
    outputs(11885) <= a xor b;
    outputs(11886) <= b;
    outputs(11887) <= not (a or b);
    outputs(11888) <= a;
    outputs(11889) <= a xor b;
    outputs(11890) <= a;
    outputs(11891) <= a xor b;
    outputs(11892) <= not (a xor b);
    outputs(11893) <= not b;
    outputs(11894) <= b;
    outputs(11895) <= not (a xor b);
    outputs(11896) <= a xor b;
    outputs(11897) <= not a;
    outputs(11898) <= not b;
    outputs(11899) <= not b;
    outputs(11900) <= a;
    outputs(11901) <= a and b;
    outputs(11902) <= b;
    outputs(11903) <= not b;
    outputs(11904) <= a and not b;
    outputs(11905) <= a xor b;
    outputs(11906) <= not b;
    outputs(11907) <= 1'b0;
    outputs(11908) <= b and not a;
    outputs(11909) <= not b;
    outputs(11910) <= a or b;
    outputs(11911) <= not a or b;
    outputs(11912) <= not (a and b);
    outputs(11913) <= a and not b;
    outputs(11914) <= not b or a;
    outputs(11915) <= a xor b;
    outputs(11916) <= not a;
    outputs(11917) <= not a;
    outputs(11918) <= not (a xor b);
    outputs(11919) <= not b;
    outputs(11920) <= a xor b;
    outputs(11921) <= b;
    outputs(11922) <= not (a xor b);
    outputs(11923) <= a xor b;
    outputs(11924) <= b and not a;
    outputs(11925) <= a;
    outputs(11926) <= not (a or b);
    outputs(11927) <= not b;
    outputs(11928) <= not (a xor b);
    outputs(11929) <= a and not b;
    outputs(11930) <= a;
    outputs(11931) <= not b;
    outputs(11932) <= a or b;
    outputs(11933) <= b and not a;
    outputs(11934) <= a and not b;
    outputs(11935) <= a xor b;
    outputs(11936) <= not (a xor b);
    outputs(11937) <= a xor b;
    outputs(11938) <= b;
    outputs(11939) <= a and not b;
    outputs(11940) <= a and b;
    outputs(11941) <= b;
    outputs(11942) <= a xor b;
    outputs(11943) <= not (a xor b);
    outputs(11944) <= not a;
    outputs(11945) <= not (a xor b);
    outputs(11946) <= b;
    outputs(11947) <= a xor b;
    outputs(11948) <= a xor b;
    outputs(11949) <= not (a xor b);
    outputs(11950) <= not b or a;
    outputs(11951) <= not a;
    outputs(11952) <= a xor b;
    outputs(11953) <= b and not a;
    outputs(11954) <= not (a xor b);
    outputs(11955) <= not (a xor b);
    outputs(11956) <= a and not b;
    outputs(11957) <= a or b;
    outputs(11958) <= not b;
    outputs(11959) <= b and not a;
    outputs(11960) <= a and b;
    outputs(11961) <= not b or a;
    outputs(11962) <= not a;
    outputs(11963) <= a and b;
    outputs(11964) <= not (a or b);
    outputs(11965) <= a xor b;
    outputs(11966) <= not (a xor b);
    outputs(11967) <= not b or a;
    outputs(11968) <= a xor b;
    outputs(11969) <= not (a xor b);
    outputs(11970) <= a xor b;
    outputs(11971) <= not (a or b);
    outputs(11972) <= b;
    outputs(11973) <= a and b;
    outputs(11974) <= not b or a;
    outputs(11975) <= a and b;
    outputs(11976) <= a xor b;
    outputs(11977) <= not (a xor b);
    outputs(11978) <= a;
    outputs(11979) <= not (a or b);
    outputs(11980) <= a xor b;
    outputs(11981) <= not a;
    outputs(11982) <= not b;
    outputs(11983) <= not (a xor b);
    outputs(11984) <= not b or a;
    outputs(11985) <= not (a xor b);
    outputs(11986) <= not (a xor b);
    outputs(11987) <= a xor b;
    outputs(11988) <= a;
    outputs(11989) <= not a;
    outputs(11990) <= not a;
    outputs(11991) <= a xor b;
    outputs(11992) <= a and b;
    outputs(11993) <= a and not b;
    outputs(11994) <= not (a or b);
    outputs(11995) <= not (a xor b);
    outputs(11996) <= not (a and b);
    outputs(11997) <= not a;
    outputs(11998) <= not a;
    outputs(11999) <= a and b;
    outputs(12000) <= b and not a;
    outputs(12001) <= a and not b;
    outputs(12002) <= a xor b;
    outputs(12003) <= not a;
    outputs(12004) <= a xor b;
    outputs(12005) <= a xor b;
    outputs(12006) <= b;
    outputs(12007) <= not a;
    outputs(12008) <= not a;
    outputs(12009) <= a xor b;
    outputs(12010) <= b;
    outputs(12011) <= a or b;
    outputs(12012) <= not a;
    outputs(12013) <= not (a xor b);
    outputs(12014) <= not (a or b);
    outputs(12015) <= b and not a;
    outputs(12016) <= not b;
    outputs(12017) <= not (a xor b);
    outputs(12018) <= not (a xor b);
    outputs(12019) <= b and not a;
    outputs(12020) <= not (a or b);
    outputs(12021) <= not a;
    outputs(12022) <= not (a or b);
    outputs(12023) <= not a;
    outputs(12024) <= not (a and b);
    outputs(12025) <= not b;
    outputs(12026) <= not a;
    outputs(12027) <= a xor b;
    outputs(12028) <= not a or b;
    outputs(12029) <= a;
    outputs(12030) <= not (a xor b);
    outputs(12031) <= a and not b;
    outputs(12032) <= a xor b;
    outputs(12033) <= not b or a;
    outputs(12034) <= not (a xor b);
    outputs(12035) <= b and not a;
    outputs(12036) <= not b;
    outputs(12037) <= a and not b;
    outputs(12038) <= not (a or b);
    outputs(12039) <= a;
    outputs(12040) <= not b;
    outputs(12041) <= not a;
    outputs(12042) <= b;
    outputs(12043) <= a and not b;
    outputs(12044) <= not b;
    outputs(12045) <= a xor b;
    outputs(12046) <= not (a or b);
    outputs(12047) <= a and not b;
    outputs(12048) <= not (a or b);
    outputs(12049) <= not (a or b);
    outputs(12050) <= a;
    outputs(12051) <= a and b;
    outputs(12052) <= not a;
    outputs(12053) <= not (a or b);
    outputs(12054) <= a xor b;
    outputs(12055) <= not a or b;
    outputs(12056) <= a;
    outputs(12057) <= not (a xor b);
    outputs(12058) <= a xor b;
    outputs(12059) <= a and not b;
    outputs(12060) <= a;
    outputs(12061) <= not a;
    outputs(12062) <= not a or b;
    outputs(12063) <= not b or a;
    outputs(12064) <= a and not b;
    outputs(12065) <= b;
    outputs(12066) <= not (a xor b);
    outputs(12067) <= a and b;
    outputs(12068) <= a xor b;
    outputs(12069) <= b;
    outputs(12070) <= a xor b;
    outputs(12071) <= a and b;
    outputs(12072) <= b and not a;
    outputs(12073) <= b;
    outputs(12074) <= a;
    outputs(12075) <= not b or a;
    outputs(12076) <= not b;
    outputs(12077) <= not a;
    outputs(12078) <= a and not b;
    outputs(12079) <= not a or b;
    outputs(12080) <= a and not b;
    outputs(12081) <= not a;
    outputs(12082) <= not b;
    outputs(12083) <= not (a and b);
    outputs(12084) <= not (a xor b);
    outputs(12085) <= not b;
    outputs(12086) <= a and b;
    outputs(12087) <= not a;
    outputs(12088) <= not (a xor b);
    outputs(12089) <= not a;
    outputs(12090) <= not (a xor b);
    outputs(12091) <= not a;
    outputs(12092) <= a and b;
    outputs(12093) <= a xor b;
    outputs(12094) <= not (a xor b);
    outputs(12095) <= not (a xor b);
    outputs(12096) <= a and not b;
    outputs(12097) <= a xor b;
    outputs(12098) <= a xor b;
    outputs(12099) <= a xor b;
    outputs(12100) <= not b;
    outputs(12101) <= a xor b;
    outputs(12102) <= b and not a;
    outputs(12103) <= a xor b;
    outputs(12104) <= not a;
    outputs(12105) <= not b;
    outputs(12106) <= not (a xor b);
    outputs(12107) <= a xor b;
    outputs(12108) <= a and not b;
    outputs(12109) <= a and not b;
    outputs(12110) <= not b;
    outputs(12111) <= not (a or b);
    outputs(12112) <= a and b;
    outputs(12113) <= not a or b;
    outputs(12114) <= a and not b;
    outputs(12115) <= a xor b;
    outputs(12116) <= a;
    outputs(12117) <= a and not b;
    outputs(12118) <= b;
    outputs(12119) <= a xor b;
    outputs(12120) <= 1'b0;
    outputs(12121) <= b and not a;
    outputs(12122) <= a;
    outputs(12123) <= not b or a;
    outputs(12124) <= b and not a;
    outputs(12125) <= b and not a;
    outputs(12126) <= b and not a;
    outputs(12127) <= a xor b;
    outputs(12128) <= not (a or b);
    outputs(12129) <= b;
    outputs(12130) <= not a;
    outputs(12131) <= not b;
    outputs(12132) <= a;
    outputs(12133) <= b and not a;
    outputs(12134) <= not (a xor b);
    outputs(12135) <= b;
    outputs(12136) <= a and b;
    outputs(12137) <= a and b;
    outputs(12138) <= b and not a;
    outputs(12139) <= not a or b;
    outputs(12140) <= not (a or b);
    outputs(12141) <= not (a xor b);
    outputs(12142) <= a and not b;
    outputs(12143) <= a;
    outputs(12144) <= not (a xor b);
    outputs(12145) <= a and b;
    outputs(12146) <= a;
    outputs(12147) <= a xor b;
    outputs(12148) <= not (a xor b);
    outputs(12149) <= b;
    outputs(12150) <= a or b;
    outputs(12151) <= not b;
    outputs(12152) <= a and not b;
    outputs(12153) <= a and not b;
    outputs(12154) <= not (a xor b);
    outputs(12155) <= a xor b;
    outputs(12156) <= not (a xor b);
    outputs(12157) <= not a;
    outputs(12158) <= b;
    outputs(12159) <= a;
    outputs(12160) <= not (a or b);
    outputs(12161) <= b and not a;
    outputs(12162) <= a xor b;
    outputs(12163) <= a xor b;
    outputs(12164) <= a and b;
    outputs(12165) <= b;
    outputs(12166) <= b;
    outputs(12167) <= a xor b;
    outputs(12168) <= not (a or b);
    outputs(12169) <= a and b;
    outputs(12170) <= not b or a;
    outputs(12171) <= not a;
    outputs(12172) <= not a;
    outputs(12173) <= a and not b;
    outputs(12174) <= not (a xor b);
    outputs(12175) <= a and b;
    outputs(12176) <= a or b;
    outputs(12177) <= not (a xor b);
    outputs(12178) <= a;
    outputs(12179) <= not (a xor b);
    outputs(12180) <= b;
    outputs(12181) <= not (a xor b);
    outputs(12182) <= not (a xor b);
    outputs(12183) <= not a or b;
    outputs(12184) <= a xor b;
    outputs(12185) <= not (a xor b);
    outputs(12186) <= b;
    outputs(12187) <= a;
    outputs(12188) <= a and not b;
    outputs(12189) <= a xor b;
    outputs(12190) <= a;
    outputs(12191) <= b;
    outputs(12192) <= not (a xor b);
    outputs(12193) <= not a or b;
    outputs(12194) <= not (a xor b);
    outputs(12195) <= a xor b;
    outputs(12196) <= not b;
    outputs(12197) <= a and not b;
    outputs(12198) <= not (a xor b);
    outputs(12199) <= not (a or b);
    outputs(12200) <= not b or a;
    outputs(12201) <= not b;
    outputs(12202) <= not (a and b);
    outputs(12203) <= not a;
    outputs(12204) <= a and not b;
    outputs(12205) <= not b;
    outputs(12206) <= not (a xor b);
    outputs(12207) <= a xor b;
    outputs(12208) <= not a;
    outputs(12209) <= not b;
    outputs(12210) <= b and not a;
    outputs(12211) <= b and not a;
    outputs(12212) <= a and b;
    outputs(12213) <= a and not b;
    outputs(12214) <= a and b;
    outputs(12215) <= b;
    outputs(12216) <= a xor b;
    outputs(12217) <= a xor b;
    outputs(12218) <= a and b;
    outputs(12219) <= b;
    outputs(12220) <= a xor b;
    outputs(12221) <= a and b;
    outputs(12222) <= b and not a;
    outputs(12223) <= not (a xor b);
    outputs(12224) <= a xor b;
    outputs(12225) <= b and not a;
    outputs(12226) <= b;
    outputs(12227) <= not b;
    outputs(12228) <= not (a and b);
    outputs(12229) <= a xor b;
    outputs(12230) <= not b or a;
    outputs(12231) <= b and not a;
    outputs(12232) <= not a;
    outputs(12233) <= not a;
    outputs(12234) <= a;
    outputs(12235) <= a and b;
    outputs(12236) <= not (a or b);
    outputs(12237) <= not (a or b);
    outputs(12238) <= a xor b;
    outputs(12239) <= a and not b;
    outputs(12240) <= a or b;
    outputs(12241) <= not (a or b);
    outputs(12242) <= a xor b;
    outputs(12243) <= a;
    outputs(12244) <= not a or b;
    outputs(12245) <= b and not a;
    outputs(12246) <= a;
    outputs(12247) <= a and not b;
    outputs(12248) <= a and b;
    outputs(12249) <= not (a xor b);
    outputs(12250) <= a and not b;
    outputs(12251) <= a xor b;
    outputs(12252) <= not (a xor b);
    outputs(12253) <= a or b;
    outputs(12254) <= a xor b;
    outputs(12255) <= b;
    outputs(12256) <= b;
    outputs(12257) <= a xor b;
    outputs(12258) <= b and not a;
    outputs(12259) <= not a;
    outputs(12260) <= a xor b;
    outputs(12261) <= not (a and b);
    outputs(12262) <= a and not b;
    outputs(12263) <= a xor b;
    outputs(12264) <= not (a or b);
    outputs(12265) <= not (a xor b);
    outputs(12266) <= not (a xor b);
    outputs(12267) <= a xor b;
    outputs(12268) <= not (a xor b);
    outputs(12269) <= not (a xor b);
    outputs(12270) <= a and not b;
    outputs(12271) <= b and not a;
    outputs(12272) <= a xor b;
    outputs(12273) <= b and not a;
    outputs(12274) <= a xor b;
    outputs(12275) <= not b;
    outputs(12276) <= a;
    outputs(12277) <= not a;
    outputs(12278) <= a;
    outputs(12279) <= not b or a;
    outputs(12280) <= b;
    outputs(12281) <= a xor b;
    outputs(12282) <= a and not b;
    outputs(12283) <= a xor b;
    outputs(12284) <= not (a xor b);
    outputs(12285) <= a xor b;
    outputs(12286) <= not (a or b);
    outputs(12287) <= b;
    outputs(12288) <= a;
    outputs(12289) <= a;
    outputs(12290) <= a xor b;
    outputs(12291) <= not (a and b);
    outputs(12292) <= b;
    outputs(12293) <= not a;
    outputs(12294) <= b and not a;
    outputs(12295) <= not a;
    outputs(12296) <= b and not a;
    outputs(12297) <= a;
    outputs(12298) <= not b;
    outputs(12299) <= not (a xor b);
    outputs(12300) <= a and b;
    outputs(12301) <= b;
    outputs(12302) <= b and not a;
    outputs(12303) <= a xor b;
    outputs(12304) <= not a;
    outputs(12305) <= a;
    outputs(12306) <= not (a xor b);
    outputs(12307) <= a xor b;
    outputs(12308) <= not a;
    outputs(12309) <= not (a or b);
    outputs(12310) <= not (a or b);
    outputs(12311) <= not a or b;
    outputs(12312) <= not (a xor b);
    outputs(12313) <= not a;
    outputs(12314) <= not (a xor b);
    outputs(12315) <= b and not a;
    outputs(12316) <= not (a xor b);
    outputs(12317) <= b and not a;
    outputs(12318) <= a xor b;
    outputs(12319) <= b and not a;
    outputs(12320) <= not (a and b);
    outputs(12321) <= not (a or b);
    outputs(12322) <= not (a or b);
    outputs(12323) <= not (a xor b);
    outputs(12324) <= a xor b;
    outputs(12325) <= not a or b;
    outputs(12326) <= not (a xor b);
    outputs(12327) <= a;
    outputs(12328) <= a xor b;
    outputs(12329) <= a;
    outputs(12330) <= a xor b;
    outputs(12331) <= a xor b;
    outputs(12332) <= a;
    outputs(12333) <= not b;
    outputs(12334) <= not b or a;
    outputs(12335) <= not (a xor b);
    outputs(12336) <= not (a or b);
    outputs(12337) <= b and not a;
    outputs(12338) <= a xor b;
    outputs(12339) <= a xor b;
    outputs(12340) <= a and b;
    outputs(12341) <= not (a or b);
    outputs(12342) <= not a or b;
    outputs(12343) <= a and not b;
    outputs(12344) <= not b;
    outputs(12345) <= a;
    outputs(12346) <= a and b;
    outputs(12347) <= not b;
    outputs(12348) <= not (a xor b);
    outputs(12349) <= a;
    outputs(12350) <= b and not a;
    outputs(12351) <= not b;
    outputs(12352) <= b;
    outputs(12353) <= a xor b;
    outputs(12354) <= not (a xor b);
    outputs(12355) <= a and not b;
    outputs(12356) <= not (a and b);
    outputs(12357) <= a and not b;
    outputs(12358) <= a xor b;
    outputs(12359) <= a;
    outputs(12360) <= not (a xor b);
    outputs(12361) <= a and not b;
    outputs(12362) <= a and b;
    outputs(12363) <= a and not b;
    outputs(12364) <= a xor b;
    outputs(12365) <= not b;
    outputs(12366) <= not (a or b);
    outputs(12367) <= not (a xor b);
    outputs(12368) <= a;
    outputs(12369) <= a or b;
    outputs(12370) <= not (a or b);
    outputs(12371) <= not b;
    outputs(12372) <= not (a xor b);
    outputs(12373) <= b and not a;
    outputs(12374) <= a and not b;
    outputs(12375) <= not (a xor b);
    outputs(12376) <= b;
    outputs(12377) <= a xor b;
    outputs(12378) <= b;
    outputs(12379) <= not a;
    outputs(12380) <= not a;
    outputs(12381) <= b;
    outputs(12382) <= b;
    outputs(12383) <= a xor b;
    outputs(12384) <= a xor b;
    outputs(12385) <= a or b;
    outputs(12386) <= not (a xor b);
    outputs(12387) <= b and not a;
    outputs(12388) <= a xor b;
    outputs(12389) <= not (a or b);
    outputs(12390) <= not (a xor b);
    outputs(12391) <= not a;
    outputs(12392) <= a and not b;
    outputs(12393) <= a xor b;
    outputs(12394) <= not b;
    outputs(12395) <= not a;
    outputs(12396) <= not (a or b);
    outputs(12397) <= a;
    outputs(12398) <= not (a or b);
    outputs(12399) <= a and b;
    outputs(12400) <= a and not b;
    outputs(12401) <= a;
    outputs(12402) <= b and not a;
    outputs(12403) <= not b;
    outputs(12404) <= not (a xor b);
    outputs(12405) <= not b;
    outputs(12406) <= a;
    outputs(12407) <= a;
    outputs(12408) <= a xor b;
    outputs(12409) <= not (a xor b);
    outputs(12410) <= not (a xor b);
    outputs(12411) <= not b;
    outputs(12412) <= b;
    outputs(12413) <= a and b;
    outputs(12414) <= b and not a;
    outputs(12415) <= a xor b;
    outputs(12416) <= not b;
    outputs(12417) <= b and not a;
    outputs(12418) <= a xor b;
    outputs(12419) <= a and b;
    outputs(12420) <= not (a and b);
    outputs(12421) <= a xor b;
    outputs(12422) <= a;
    outputs(12423) <= a;
    outputs(12424) <= not a;
    outputs(12425) <= not (a xor b);
    outputs(12426) <= not a;
    outputs(12427) <= a and not b;
    outputs(12428) <= a xor b;
    outputs(12429) <= not (a or b);
    outputs(12430) <= a xor b;
    outputs(12431) <= not b;
    outputs(12432) <= a and not b;
    outputs(12433) <= b;
    outputs(12434) <= a and b;
    outputs(12435) <= not (a xor b);
    outputs(12436) <= not a or b;
    outputs(12437) <= not (a xor b);
    outputs(12438) <= not a or b;
    outputs(12439) <= not a;
    outputs(12440) <= not a;
    outputs(12441) <= not b;
    outputs(12442) <= not (a or b);
    outputs(12443) <= b;
    outputs(12444) <= not b or a;
    outputs(12445) <= not a;
    outputs(12446) <= b and not a;
    outputs(12447) <= not b;
    outputs(12448) <= not (a xor b);
    outputs(12449) <= not a;
    outputs(12450) <= not (a or b);
    outputs(12451) <= not a;
    outputs(12452) <= a;
    outputs(12453) <= not a;
    outputs(12454) <= a;
    outputs(12455) <= not (a xor b);
    outputs(12456) <= not (a xor b);
    outputs(12457) <= a and not b;
    outputs(12458) <= b and not a;
    outputs(12459) <= a and b;
    outputs(12460) <= a;
    outputs(12461) <= a xor b;
    outputs(12462) <= b and not a;
    outputs(12463) <= not b;
    outputs(12464) <= b and not a;
    outputs(12465) <= not b or a;
    outputs(12466) <= a xor b;
    outputs(12467) <= not (a xor b);
    outputs(12468) <= b and not a;
    outputs(12469) <= a and b;
    outputs(12470) <= a;
    outputs(12471) <= a xor b;
    outputs(12472) <= a and b;
    outputs(12473) <= a xor b;
    outputs(12474) <= not (a or b);
    outputs(12475) <= not (a or b);
    outputs(12476) <= a xor b;
    outputs(12477) <= a and not b;
    outputs(12478) <= not (a and b);
    outputs(12479) <= not (a xor b);
    outputs(12480) <= not (a xor b);
    outputs(12481) <= not (a and b);
    outputs(12482) <= not a;
    outputs(12483) <= b;
    outputs(12484) <= not a;
    outputs(12485) <= a and b;
    outputs(12486) <= not b;
    outputs(12487) <= a and b;
    outputs(12488) <= b and not a;
    outputs(12489) <= not b;
    outputs(12490) <= a;
    outputs(12491) <= not (a xor b);
    outputs(12492) <= a xor b;
    outputs(12493) <= not b;
    outputs(12494) <= b;
    outputs(12495) <= not a;
    outputs(12496) <= not b;
    outputs(12497) <= a and not b;
    outputs(12498) <= not a;
    outputs(12499) <= not b or a;
    outputs(12500) <= a and b;
    outputs(12501) <= not (a or b);
    outputs(12502) <= a and b;
    outputs(12503) <= not (a and b);
    outputs(12504) <= a and b;
    outputs(12505) <= not (a xor b);
    outputs(12506) <= a xor b;
    outputs(12507) <= b;
    outputs(12508) <= not a or b;
    outputs(12509) <= not (a xor b);
    outputs(12510) <= b;
    outputs(12511) <= not (a xor b);
    outputs(12512) <= not b;
    outputs(12513) <= not b;
    outputs(12514) <= a xor b;
    outputs(12515) <= not (a or b);
    outputs(12516) <= not (a xor b);
    outputs(12517) <= not (a xor b);
    outputs(12518) <= a and b;
    outputs(12519) <= not (a xor b);
    outputs(12520) <= a xor b;
    outputs(12521) <= not (a xor b);
    outputs(12522) <= not (a xor b);
    outputs(12523) <= a;
    outputs(12524) <= not a;
    outputs(12525) <= not (a xor b);
    outputs(12526) <= b;
    outputs(12527) <= b and not a;
    outputs(12528) <= a xor b;
    outputs(12529) <= not (a or b);
    outputs(12530) <= a xor b;
    outputs(12531) <= a and b;
    outputs(12532) <= a xor b;
    outputs(12533) <= a and not b;
    outputs(12534) <= not (a xor b);
    outputs(12535) <= a or b;
    outputs(12536) <= not a;
    outputs(12537) <= not b;
    outputs(12538) <= not a;
    outputs(12539) <= a xor b;
    outputs(12540) <= not a;
    outputs(12541) <= b;
    outputs(12542) <= not (a or b);
    outputs(12543) <= b and not a;
    outputs(12544) <= a;
    outputs(12545) <= a xor b;
    outputs(12546) <= a xor b;
    outputs(12547) <= not a;
    outputs(12548) <= b and not a;
    outputs(12549) <= a or b;
    outputs(12550) <= b and not a;
    outputs(12551) <= not a;
    outputs(12552) <= not (a xor b);
    outputs(12553) <= b and not a;
    outputs(12554) <= not (a xor b);
    outputs(12555) <= a xor b;
    outputs(12556) <= a and not b;
    outputs(12557) <= a and b;
    outputs(12558) <= a and not b;
    outputs(12559) <= not a or b;
    outputs(12560) <= not b;
    outputs(12561) <= not (a xor b);
    outputs(12562) <= not (a xor b);
    outputs(12563) <= not (a xor b);
    outputs(12564) <= a xor b;
    outputs(12565) <= a and b;
    outputs(12566) <= not (a or b);
    outputs(12567) <= a and b;
    outputs(12568) <= not a;
    outputs(12569) <= a and b;
    outputs(12570) <= not a;
    outputs(12571) <= not (a or b);
    outputs(12572) <= a;
    outputs(12573) <= a xor b;
    outputs(12574) <= a and b;
    outputs(12575) <= not a;
    outputs(12576) <= a;
    outputs(12577) <= a or b;
    outputs(12578) <= a xor b;
    outputs(12579) <= not b;
    outputs(12580) <= a;
    outputs(12581) <= not a;
    outputs(12582) <= a;
    outputs(12583) <= b;
    outputs(12584) <= b and not a;
    outputs(12585) <= a and b;
    outputs(12586) <= not b or a;
    outputs(12587) <= not (a xor b);
    outputs(12588) <= b;
    outputs(12589) <= not (a xor b);
    outputs(12590) <= not a or b;
    outputs(12591) <= not (a or b);
    outputs(12592) <= a and not b;
    outputs(12593) <= not (a xor b);
    outputs(12594) <= not (a and b);
    outputs(12595) <= not (a or b);
    outputs(12596) <= a and b;
    outputs(12597) <= not (a xor b);
    outputs(12598) <= b;
    outputs(12599) <= a;
    outputs(12600) <= b and not a;
    outputs(12601) <= not b;
    outputs(12602) <= a xor b;
    outputs(12603) <= a and b;
    outputs(12604) <= a and b;
    outputs(12605) <= not (a and b);
    outputs(12606) <= not (a xor b);
    outputs(12607) <= not (a or b);
    outputs(12608) <= not (a and b);
    outputs(12609) <= not (a or b);
    outputs(12610) <= not a;
    outputs(12611) <= a xor b;
    outputs(12612) <= not (a xor b);
    outputs(12613) <= not b;
    outputs(12614) <= not a;
    outputs(12615) <= not (a xor b);
    outputs(12616) <= not (a xor b);
    outputs(12617) <= a and b;
    outputs(12618) <= a and not b;
    outputs(12619) <= a;
    outputs(12620) <= a;
    outputs(12621) <= not (a or b);
    outputs(12622) <= not a;
    outputs(12623) <= not b or a;
    outputs(12624) <= not (a and b);
    outputs(12625) <= b;
    outputs(12626) <= a and b;
    outputs(12627) <= b;
    outputs(12628) <= not a;
    outputs(12629) <= not (a xor b);
    outputs(12630) <= not a or b;
    outputs(12631) <= not (a xor b);
    outputs(12632) <= not (a xor b);
    outputs(12633) <= not b;
    outputs(12634) <= a xor b;
    outputs(12635) <= not a;
    outputs(12636) <= not (a xor b);
    outputs(12637) <= a xor b;
    outputs(12638) <= a and b;
    outputs(12639) <= not (a xor b);
    outputs(12640) <= not (a or b);
    outputs(12641) <= not b;
    outputs(12642) <= a;
    outputs(12643) <= b and not a;
    outputs(12644) <= not (a xor b);
    outputs(12645) <= not (a or b);
    outputs(12646) <= not a;
    outputs(12647) <= not a or b;
    outputs(12648) <= not (a xor b);
    outputs(12649) <= b;
    outputs(12650) <= not (a xor b);
    outputs(12651) <= b and not a;
    outputs(12652) <= b and not a;
    outputs(12653) <= b and not a;
    outputs(12654) <= not a or b;
    outputs(12655) <= not (a or b);
    outputs(12656) <= not a;
    outputs(12657) <= a xor b;
    outputs(12658) <= not b;
    outputs(12659) <= not a;
    outputs(12660) <= a xor b;
    outputs(12661) <= a xor b;
    outputs(12662) <= a xor b;
    outputs(12663) <= b and not a;
    outputs(12664) <= a xor b;
    outputs(12665) <= not a;
    outputs(12666) <= b;
    outputs(12667) <= a xor b;
    outputs(12668) <= a and not b;
    outputs(12669) <= not a;
    outputs(12670) <= a;
    outputs(12671) <= a xor b;
    outputs(12672) <= b and not a;
    outputs(12673) <= not a;
    outputs(12674) <= not b;
    outputs(12675) <= not a or b;
    outputs(12676) <= not a;
    outputs(12677) <= not a;
    outputs(12678) <= b and not a;
    outputs(12679) <= not (a xor b);
    outputs(12680) <= not b;
    outputs(12681) <= not (a xor b);
    outputs(12682) <= a or b;
    outputs(12683) <= a and b;
    outputs(12684) <= b and not a;
    outputs(12685) <= a and b;
    outputs(12686) <= not (a xor b);
    outputs(12687) <= not (a xor b);
    outputs(12688) <= a or b;
    outputs(12689) <= not (a xor b);
    outputs(12690) <= not (a xor b);
    outputs(12691) <= a xor b;
    outputs(12692) <= not b or a;
    outputs(12693) <= a;
    outputs(12694) <= not (a and b);
    outputs(12695) <= b;
    outputs(12696) <= not b;
    outputs(12697) <= not (a xor b);
    outputs(12698) <= a;
    outputs(12699) <= a;
    outputs(12700) <= not a or b;
    outputs(12701) <= not (a xor b);
    outputs(12702) <= not (a xor b);
    outputs(12703) <= not (a xor b);
    outputs(12704) <= not (a xor b);
    outputs(12705) <= a xor b;
    outputs(12706) <= a and b;
    outputs(12707) <= a;
    outputs(12708) <= b;
    outputs(12709) <= not (a xor b);
    outputs(12710) <= not b;
    outputs(12711) <= not (a xor b);
    outputs(12712) <= not a;
    outputs(12713) <= b;
    outputs(12714) <= not (a xor b);
    outputs(12715) <= a and b;
    outputs(12716) <= not a;
    outputs(12717) <= b and not a;
    outputs(12718) <= b and not a;
    outputs(12719) <= b and not a;
    outputs(12720) <= a;
    outputs(12721) <= a xor b;
    outputs(12722) <= not (a xor b);
    outputs(12723) <= not b;
    outputs(12724) <= not (a xor b);
    outputs(12725) <= not a;
    outputs(12726) <= b;
    outputs(12727) <= a and not b;
    outputs(12728) <= a or b;
    outputs(12729) <= not (a xor b);
    outputs(12730) <= a;
    outputs(12731) <= a xor b;
    outputs(12732) <= b;
    outputs(12733) <= b and not a;
    outputs(12734) <= b;
    outputs(12735) <= not (a xor b);
    outputs(12736) <= not (a or b);
    outputs(12737) <= a xor b;
    outputs(12738) <= a or b;
    outputs(12739) <= a;
    outputs(12740) <= not b;
    outputs(12741) <= not (a and b);
    outputs(12742) <= a and b;
    outputs(12743) <= b;
    outputs(12744) <= not b;
    outputs(12745) <= not b;
    outputs(12746) <= not b;
    outputs(12747) <= a or b;
    outputs(12748) <= a;
    outputs(12749) <= a or b;
    outputs(12750) <= not b;
    outputs(12751) <= a and b;
    outputs(12752) <= a xor b;
    outputs(12753) <= not a;
    outputs(12754) <= a xor b;
    outputs(12755) <= a;
    outputs(12756) <= not (a or b);
    outputs(12757) <= not (a or b);
    outputs(12758) <= a;
    outputs(12759) <= not a;
    outputs(12760) <= not b;
    outputs(12761) <= a xor b;
    outputs(12762) <= b;
    outputs(12763) <= not a or b;
    outputs(12764) <= a xor b;
    outputs(12765) <= a xor b;
    outputs(12766) <= not (a xor b);
    outputs(12767) <= not a;
    outputs(12768) <= not b;
    outputs(12769) <= b and not a;
    outputs(12770) <= a and b;
    outputs(12771) <= not (a and b);
    outputs(12772) <= a and b;
    outputs(12773) <= a and b;
    outputs(12774) <= a;
    outputs(12775) <= a xor b;
    outputs(12776) <= not b or a;
    outputs(12777) <= a and not b;
    outputs(12778) <= not (a xor b);
    outputs(12779) <= b and not a;
    outputs(12780) <= a;
    outputs(12781) <= b;
    outputs(12782) <= not (a xor b);
    outputs(12783) <= not (a and b);
    outputs(12784) <= not (a xor b);
    outputs(12785) <= not (a xor b);
    outputs(12786) <= b and not a;
    outputs(12787) <= not a;
    outputs(12788) <= a xor b;
    outputs(12789) <= not (a or b);
    outputs(12790) <= not (a or b);
    outputs(12791) <= not b or a;
    outputs(12792) <= a and not b;
    outputs(12793) <= not a;
    outputs(12794) <= a and not b;
    outputs(12795) <= a xor b;
    outputs(12796) <= a xor b;
    outputs(12797) <= not a;
    outputs(12798) <= a xor b;
    outputs(12799) <= not (a xor b);
end Behavioral;
